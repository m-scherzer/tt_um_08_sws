VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_08_sws
  CLASS BLOCK ;
  FOREIGN tt_um_08_sws ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 200.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNADIFFAREA 394.109192 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 10.655 206.170 10.825 206.360 ;
        RECT 12.090 206.220 12.210 206.330 ;
        RECT 13.875 206.170 14.045 206.360 ;
        RECT 19.395 206.170 19.565 206.360 ;
        RECT 24.915 206.170 25.085 206.360 ;
        RECT 26.755 206.170 26.925 206.360 ;
        RECT 32.275 206.170 32.445 206.360 ;
        RECT 37.795 206.170 37.965 206.360 ;
        RECT 39.635 206.170 39.805 206.360 ;
        RECT 45.155 206.170 45.325 206.360 ;
        RECT 50.675 206.170 50.845 206.360 ;
        RECT 52.515 206.170 52.685 206.360 ;
        RECT 58.035 206.170 58.205 206.360 ;
        RECT 63.555 206.170 63.725 206.360 ;
        RECT 65.855 206.170 66.025 206.360 ;
        RECT 66.315 206.170 66.485 206.360 ;
        RECT 70.915 206.170 71.085 206.360 ;
        RECT 76.435 206.170 76.605 206.360 ;
        RECT 78.275 206.170 78.445 206.360 ;
        RECT 83.795 206.170 83.965 206.360 ;
        RECT 89.315 206.170 89.485 206.360 ;
        RECT 91.155 206.170 91.325 206.360 ;
        RECT 96.675 206.170 96.845 206.360 ;
        RECT 102.195 206.170 102.365 206.360 ;
        RECT 103.170 206.220 103.290 206.330 ;
        RECT 108.635 206.170 108.805 206.360 ;
        RECT 114.155 206.170 114.325 206.360 ;
        RECT 115.535 206.170 115.705 206.360 ;
        RECT 10.515 205.360 11.885 206.170 ;
        RECT 12.365 205.300 12.795 206.085 ;
        RECT 12.815 205.360 14.185 206.170 ;
        RECT 14.195 205.360 19.705 206.170 ;
        RECT 19.715 205.360 25.225 206.170 ;
        RECT 25.245 205.300 25.675 206.085 ;
        RECT 25.695 205.360 27.065 206.170 ;
        RECT 27.075 205.360 32.585 206.170 ;
        RECT 32.595 205.360 38.105 206.170 ;
        RECT 38.125 205.300 38.555 206.085 ;
        RECT 38.575 205.360 39.945 206.170 ;
        RECT 39.955 205.360 45.465 206.170 ;
        RECT 45.475 205.360 50.985 206.170 ;
        RECT 51.005 205.300 51.435 206.085 ;
        RECT 51.455 205.360 52.825 206.170 ;
        RECT 52.835 205.360 58.345 206.170 ;
        RECT 58.355 205.360 63.865 206.170 ;
        RECT 63.885 205.300 64.315 206.085 ;
        RECT 64.335 205.360 66.165 206.170 ;
        RECT 66.185 205.260 67.535 206.170 ;
        RECT 67.555 205.360 71.225 206.170 ;
        RECT 71.235 205.360 76.745 206.170 ;
        RECT 76.765 205.300 77.195 206.085 ;
        RECT 77.215 205.360 78.585 206.170 ;
        RECT 78.595 205.360 84.105 206.170 ;
        RECT 84.115 205.360 89.625 206.170 ;
        RECT 89.645 205.300 90.075 206.085 ;
        RECT 90.095 205.360 91.465 206.170 ;
        RECT 91.475 205.360 96.985 206.170 ;
        RECT 96.995 205.360 102.505 206.170 ;
        RECT 102.525 205.300 102.955 206.085 ;
        RECT 103.435 205.360 108.945 206.170 ;
        RECT 108.955 205.360 114.465 206.170 ;
        RECT 114.475 205.360 115.845 206.170 ;
      LAYER nwell ;
        RECT 10.320 202.140 116.040 204.970 ;
      LAYER pwell ;
        RECT 10.515 200.940 11.885 201.750 ;
        RECT 12.365 201.025 12.795 201.810 ;
        RECT 13.275 200.940 16.025 201.750 ;
        RECT 16.035 200.940 21.545 201.750 ;
        RECT 21.555 200.940 27.065 201.750 ;
        RECT 27.075 200.940 32.585 201.750 ;
        RECT 32.595 200.940 38.105 201.750 ;
        RECT 38.125 201.025 38.555 201.810 ;
        RECT 39.495 200.940 45.005 201.750 ;
        RECT 45.015 200.940 50.525 201.750 ;
        RECT 50.535 200.940 56.045 201.750 ;
        RECT 56.065 200.940 57.415 201.850 ;
        RECT 57.435 200.940 60.185 201.750 ;
        RECT 60.195 200.940 61.565 201.720 ;
        RECT 61.575 201.620 62.495 201.850 ;
        RECT 61.575 200.940 63.865 201.620 ;
        RECT 63.885 201.025 64.315 201.810 ;
        RECT 64.335 201.620 65.255 201.850 ;
        RECT 68.085 201.620 69.015 201.840 ;
        RECT 64.335 200.940 73.525 201.620 ;
        RECT 73.995 200.940 75.825 201.750 ;
        RECT 75.835 200.940 77.205 201.720 ;
        RECT 77.215 200.940 78.585 201.750 ;
        RECT 78.595 200.940 84.105 201.750 ;
        RECT 84.115 200.940 89.625 201.750 ;
        RECT 89.645 201.025 90.075 201.810 ;
        RECT 90.555 200.940 92.385 201.750 ;
        RECT 92.395 200.940 97.905 201.750 ;
        RECT 97.915 200.940 103.425 201.750 ;
        RECT 103.435 200.940 108.945 201.750 ;
        RECT 108.955 200.940 114.465 201.750 ;
        RECT 114.475 200.940 115.845 201.750 ;
        RECT 10.655 200.730 10.825 200.940 ;
        RECT 12.090 200.780 12.210 200.890 ;
        RECT 13.010 200.780 13.130 200.890 ;
        RECT 13.875 200.730 14.045 200.920 ;
        RECT 15.715 200.750 15.885 200.940 ;
        RECT 19.395 200.730 19.565 200.920 ;
        RECT 21.235 200.750 21.405 200.940 ;
        RECT 24.915 200.730 25.085 200.920 ;
        RECT 25.890 200.780 26.010 200.890 ;
        RECT 26.755 200.750 26.925 200.940 ;
        RECT 28.595 200.730 28.765 200.920 ;
        RECT 32.275 200.750 32.445 200.940 ;
        RECT 34.115 200.730 34.285 200.920 ;
        RECT 37.795 200.750 37.965 200.940 ;
        RECT 39.175 200.785 39.335 200.895 ;
        RECT 39.635 200.730 39.805 200.920 ;
        RECT 44.695 200.750 44.865 200.940 ;
        RECT 45.155 200.730 45.325 200.920 ;
        RECT 50.215 200.750 50.385 200.940 ;
        RECT 50.675 200.730 50.845 200.920 ;
        RECT 55.735 200.750 55.905 200.940 ;
        RECT 57.115 200.750 57.285 200.940 ;
        RECT 59.875 200.750 60.045 200.940 ;
        RECT 61.255 200.750 61.425 200.940 ;
        RECT 61.715 200.730 61.885 200.920 ;
        RECT 62.230 200.780 62.350 200.890 ;
        RECT 10.515 199.920 11.885 200.730 ;
        RECT 12.355 199.920 14.185 200.730 ;
        RECT 14.195 199.920 19.705 200.730 ;
        RECT 19.715 199.920 25.225 200.730 ;
        RECT 25.245 199.860 25.675 200.645 ;
        RECT 26.155 199.920 28.905 200.730 ;
        RECT 28.915 199.920 34.425 200.730 ;
        RECT 34.435 199.920 39.945 200.730 ;
        RECT 39.955 199.920 45.465 200.730 ;
        RECT 45.475 199.920 50.985 200.730 ;
        RECT 51.005 199.860 51.435 200.645 ;
        RECT 51.655 200.050 62.025 200.730 ;
        RECT 62.635 200.700 62.805 200.920 ;
        RECT 63.555 200.750 63.725 200.940 ;
        RECT 65.855 200.730 66.025 200.920 ;
        RECT 73.215 200.750 73.385 200.940 ;
        RECT 73.730 200.780 73.850 200.890 ;
        RECT 75.515 200.750 75.685 200.940 ;
        RECT 76.435 200.730 76.605 200.920 ;
        RECT 76.895 200.750 77.065 200.940 ;
        RECT 78.275 200.730 78.445 200.940 ;
        RECT 80.115 200.730 80.285 200.920 ;
        RECT 83.795 200.750 83.965 200.940 ;
        RECT 85.635 200.730 85.805 200.920 ;
        RECT 89.315 200.750 89.485 200.940 ;
        RECT 90.290 200.780 90.410 200.890 ;
        RECT 91.155 200.730 91.325 200.920 ;
        RECT 92.075 200.750 92.245 200.940 ;
        RECT 96.675 200.730 96.845 200.920 ;
        RECT 97.595 200.750 97.765 200.940 ;
        RECT 102.195 200.730 102.365 200.920 ;
        RECT 103.115 200.890 103.285 200.940 ;
        RECT 103.115 200.780 103.290 200.890 ;
        RECT 103.115 200.750 103.285 200.780 ;
        RECT 108.635 200.730 108.805 200.940 ;
        RECT 114.155 200.730 114.325 200.940 ;
        RECT 115.535 200.730 115.705 200.940 ;
        RECT 64.760 200.700 65.705 200.730 ;
        RECT 62.635 200.500 65.705 200.700 ;
        RECT 51.655 199.820 53.865 200.050 ;
        RECT 56.585 199.830 57.515 200.050 ;
        RECT 62.495 200.020 65.705 200.500 ;
        RECT 65.715 200.050 67.545 200.730 ;
        RECT 62.495 199.820 63.425 200.020 ;
        RECT 64.760 199.820 65.705 200.020 ;
        RECT 66.200 199.820 67.545 200.050 ;
        RECT 67.555 200.050 76.745 200.730 ;
        RECT 67.555 199.820 68.475 200.050 ;
        RECT 71.305 199.830 72.235 200.050 ;
        RECT 76.765 199.860 77.195 200.645 ;
        RECT 77.225 199.820 78.575 200.730 ;
        RECT 78.595 199.920 80.425 200.730 ;
        RECT 80.435 199.920 85.945 200.730 ;
        RECT 85.955 199.920 91.465 200.730 ;
        RECT 91.475 199.920 96.985 200.730 ;
        RECT 96.995 199.920 102.505 200.730 ;
        RECT 102.525 199.860 102.955 200.645 ;
        RECT 103.435 199.920 108.945 200.730 ;
        RECT 108.955 199.920 114.465 200.730 ;
        RECT 114.475 199.920 115.845 200.730 ;
      LAYER nwell ;
        RECT 10.320 196.700 116.040 199.530 ;
      LAYER pwell ;
        RECT 10.515 195.500 11.885 196.310 ;
        RECT 12.365 195.585 12.795 196.370 ;
        RECT 13.275 195.500 16.025 196.310 ;
        RECT 16.035 195.500 21.545 196.310 ;
        RECT 21.555 195.500 27.065 196.310 ;
        RECT 27.075 195.500 32.585 196.310 ;
        RECT 32.595 195.500 38.105 196.310 ;
        RECT 38.125 195.585 38.555 196.370 ;
        RECT 38.575 195.500 44.085 196.310 ;
        RECT 44.095 195.500 49.605 196.310 ;
        RECT 54.125 196.180 55.055 196.400 ;
        RECT 57.885 196.180 59.225 196.410 ;
        RECT 49.615 195.500 59.225 196.180 ;
        RECT 59.275 195.500 62.385 196.410 ;
        RECT 62.515 195.500 63.865 196.410 ;
        RECT 63.885 195.585 64.315 196.370 ;
        RECT 64.335 195.500 67.255 196.410 ;
        RECT 68.575 195.500 71.685 196.410 ;
        RECT 71.695 196.180 72.615 196.410 ;
        RECT 75.445 196.180 76.375 196.400 ;
        RECT 71.695 195.500 80.885 196.180 ;
        RECT 81.355 195.500 84.105 196.310 ;
        RECT 84.115 195.500 89.625 196.310 ;
        RECT 89.645 195.585 90.075 196.370 ;
        RECT 90.555 195.500 92.385 196.310 ;
        RECT 92.395 195.500 97.905 196.310 ;
        RECT 97.915 195.500 103.425 196.310 ;
        RECT 103.435 195.500 108.945 196.310 ;
        RECT 108.955 195.500 114.465 196.310 ;
        RECT 114.475 195.500 115.845 196.310 ;
        RECT 10.655 195.290 10.825 195.500 ;
        RECT 12.090 195.340 12.210 195.450 ;
        RECT 13.010 195.340 13.130 195.450 ;
        RECT 13.875 195.290 14.045 195.480 ;
        RECT 15.715 195.310 15.885 195.500 ;
        RECT 19.395 195.290 19.565 195.480 ;
        RECT 21.235 195.310 21.405 195.500 ;
        RECT 24.915 195.290 25.085 195.480 ;
        RECT 26.755 195.310 26.925 195.500 ;
        RECT 30.895 195.290 31.065 195.480 ;
        RECT 32.275 195.310 32.445 195.500 ;
        RECT 36.415 195.290 36.585 195.480 ;
        RECT 37.795 195.310 37.965 195.500 ;
        RECT 41.935 195.290 42.105 195.480 ;
        RECT 42.395 195.290 42.565 195.480 ;
        RECT 43.775 195.310 43.945 195.500 ;
        RECT 45.155 195.290 45.325 195.480 ;
        RECT 49.295 195.310 49.465 195.500 ;
        RECT 49.755 195.310 49.925 195.500 ;
        RECT 50.675 195.290 50.845 195.480 ;
        RECT 53.895 195.290 54.065 195.480 ;
        RECT 55.275 195.290 55.445 195.480 ;
        RECT 55.790 195.340 55.910 195.450 ;
        RECT 56.195 195.290 56.365 195.480 ;
        RECT 60.795 195.290 60.965 195.480 ;
        RECT 10.515 194.480 11.885 195.290 ;
        RECT 12.355 194.480 14.185 195.290 ;
        RECT 14.195 194.480 19.705 195.290 ;
        RECT 19.715 194.480 25.225 195.290 ;
        RECT 25.245 194.420 25.675 195.205 ;
        RECT 25.695 194.480 31.205 195.290 ;
        RECT 31.215 194.480 36.725 195.290 ;
        RECT 36.735 194.480 42.245 195.290 ;
        RECT 42.265 194.380 43.615 195.290 ;
        RECT 43.635 194.480 45.465 195.290 ;
        RECT 45.475 194.480 50.985 195.290 ;
        RECT 51.005 194.420 51.435 195.205 ;
        RECT 51.455 194.480 54.205 195.290 ;
        RECT 54.225 194.380 55.575 195.290 ;
        RECT 56.165 194.610 59.630 195.290 ;
        RECT 58.710 194.380 59.630 194.610 ;
        RECT 59.735 194.480 61.105 195.290 ;
        RECT 61.255 195.260 61.425 195.480 ;
        RECT 62.175 195.310 62.345 195.500 ;
        RECT 62.630 195.310 62.800 195.500 ;
        RECT 64.480 195.310 64.650 195.500 ;
        RECT 67.695 195.290 67.865 195.480 ;
        RECT 68.155 195.345 68.315 195.455 ;
        RECT 68.615 195.310 68.785 195.500 ;
        RECT 69.075 195.310 69.245 195.480 ;
        RECT 69.080 195.290 69.245 195.310 ;
        RECT 71.375 195.290 71.545 195.480 ;
        RECT 73.730 195.340 73.850 195.450 ;
        RECT 74.135 195.290 74.305 195.480 ;
        RECT 75.515 195.290 75.685 195.480 ;
        RECT 77.815 195.335 77.975 195.445 ;
        RECT 80.575 195.310 80.745 195.500 ;
        RECT 81.090 195.340 81.210 195.450 ;
        RECT 81.495 195.290 81.665 195.480 ;
        RECT 83.795 195.310 83.965 195.500 ;
        RECT 87.015 195.290 87.185 195.480 ;
        RECT 87.475 195.290 87.645 195.480 ;
        RECT 89.315 195.310 89.485 195.500 ;
        RECT 90.290 195.340 90.410 195.450 ;
        RECT 92.075 195.310 92.245 195.500 ;
        RECT 97.135 195.335 97.295 195.445 ;
        RECT 97.595 195.310 97.765 195.500 ;
        RECT 100.815 195.290 100.985 195.480 ;
        RECT 102.195 195.290 102.365 195.480 ;
        RECT 103.115 195.310 103.285 195.500 ;
        RECT 103.575 195.335 103.735 195.445 ;
        RECT 104.035 195.290 104.205 195.480 ;
        RECT 108.635 195.290 108.805 195.500 ;
        RECT 114.155 195.290 114.325 195.500 ;
        RECT 115.535 195.290 115.705 195.500 ;
        RECT 63.380 195.260 64.325 195.290 ;
        RECT 61.255 195.060 64.325 195.260 ;
        RECT 61.115 194.580 64.325 195.060 ;
        RECT 61.115 194.380 62.045 194.580 ;
        RECT 63.380 194.380 64.325 194.580 ;
        RECT 64.335 194.610 68.005 195.290 ;
        RECT 69.080 194.610 70.915 195.290 ;
        RECT 71.235 194.610 73.525 195.290 ;
        RECT 64.335 194.380 65.265 194.610 ;
        RECT 69.985 194.380 70.915 194.610 ;
        RECT 72.605 194.380 73.525 194.610 ;
        RECT 74.005 194.380 75.355 195.290 ;
        RECT 75.385 194.380 76.735 195.290 ;
        RECT 76.765 194.420 77.195 195.205 ;
        RECT 78.135 194.480 81.805 195.290 ;
        RECT 81.815 194.480 87.325 195.290 ;
        RECT 87.335 194.610 96.525 195.290 ;
        RECT 91.845 194.390 92.775 194.610 ;
        RECT 95.605 194.380 96.525 194.610 ;
        RECT 97.455 194.480 101.125 195.290 ;
        RECT 101.145 194.380 102.495 195.290 ;
        RECT 102.525 194.420 102.955 195.205 ;
        RECT 103.895 194.510 105.265 195.290 ;
        RECT 105.275 194.480 108.945 195.290 ;
        RECT 108.955 194.480 114.465 195.290 ;
        RECT 114.475 194.480 115.845 195.290 ;
      LAYER nwell ;
        RECT 10.320 191.260 116.040 194.090 ;
      LAYER pwell ;
        RECT 10.515 190.060 11.885 190.870 ;
        RECT 12.365 190.145 12.795 190.930 ;
        RECT 13.735 190.060 17.405 190.870 ;
        RECT 17.415 190.060 22.925 190.870 ;
        RECT 23.305 190.860 24.225 190.970 ;
        RECT 23.305 190.740 25.640 190.860 ;
        RECT 30.305 190.740 31.225 190.960 ;
        RECT 23.305 190.060 32.585 190.740 ;
        RECT 32.595 190.060 38.105 190.870 ;
        RECT 38.125 190.145 38.555 190.930 ;
        RECT 39.505 190.060 40.855 190.970 ;
        RECT 43.530 190.740 44.450 190.970 ;
        RECT 40.985 190.060 44.450 190.740 ;
        RECT 45.475 190.060 46.845 190.840 ;
        RECT 47.775 190.060 53.285 190.870 ;
        RECT 53.295 190.060 58.805 190.870 ;
        RECT 58.815 190.060 61.105 190.970 ;
        RECT 61.115 190.060 63.865 190.870 ;
        RECT 63.885 190.145 64.315 190.930 ;
        RECT 65.265 190.740 68.265 190.970 ;
        RECT 69.950 190.740 70.870 190.970 ;
        RECT 65.265 190.650 69.845 190.740 ;
        RECT 65.255 190.290 69.845 190.650 ;
        RECT 65.255 190.100 66.185 190.290 ;
        RECT 65.265 190.060 66.185 190.100 ;
        RECT 68.275 190.060 69.845 190.290 ;
        RECT 69.950 190.060 73.415 190.740 ;
        RECT 73.535 190.060 74.905 190.870 ;
        RECT 74.915 190.060 80.425 190.870 ;
        RECT 80.445 190.060 81.795 190.970 ;
        RECT 81.815 190.060 83.185 190.840 ;
        RECT 83.195 190.060 84.565 190.870 ;
        RECT 84.575 190.060 88.245 190.870 ;
        RECT 88.265 190.060 89.615 190.970 ;
        RECT 89.645 190.145 90.075 190.930 ;
        RECT 90.190 190.740 91.110 190.970 ;
        RECT 97.350 190.740 98.270 190.970 ;
        RECT 90.190 190.060 93.655 190.740 ;
        RECT 94.805 190.060 98.270 190.740 ;
        RECT 98.375 190.740 99.295 190.970 ;
        RECT 102.125 190.740 103.055 190.960 ;
        RECT 98.375 190.060 107.565 190.740 ;
        RECT 107.575 190.060 109.405 190.870 ;
        RECT 109.415 190.060 110.785 190.840 ;
        RECT 110.795 190.060 114.465 190.870 ;
        RECT 114.475 190.060 115.845 190.870 ;
        RECT 10.655 189.850 10.825 190.060 ;
        RECT 12.090 189.900 12.210 190.010 ;
        RECT 12.495 189.895 12.655 190.005 ;
        RECT 13.415 189.905 13.575 190.015 ;
        RECT 17.095 189.870 17.265 190.060 ;
        RECT 18.015 189.850 18.185 190.040 ;
        RECT 22.615 189.870 22.785 190.060 ;
        RECT 23.535 189.850 23.705 190.040 ;
        RECT 23.995 189.850 24.165 190.040 ;
        RECT 26.295 189.895 26.455 190.005 ;
        RECT 30.160 189.850 30.330 190.040 ;
        RECT 30.950 189.900 31.070 190.010 ;
        RECT 31.355 189.850 31.525 190.040 ;
        RECT 32.275 189.870 32.445 190.060 ;
        RECT 35.955 189.850 36.125 190.040 ;
        RECT 36.690 189.850 36.860 190.040 ;
        RECT 37.795 189.870 37.965 190.060 ;
        RECT 39.175 189.905 39.335 190.015 ;
        RECT 40.555 189.870 40.725 190.060 ;
        RECT 41.015 189.870 41.185 190.060 ;
        RECT 45.155 189.905 45.315 190.015 ;
        RECT 45.615 189.870 45.785 190.060 ;
        RECT 47.455 189.905 47.615 190.015 ;
        RECT 49.295 189.850 49.465 190.040 ;
        RECT 50.675 189.850 50.845 190.040 ;
        RECT 51.650 189.900 51.770 190.010 ;
        RECT 52.975 189.870 53.145 190.060 ;
        RECT 54.355 189.850 54.525 190.040 ;
        RECT 54.815 189.850 54.985 190.040 ;
        RECT 57.115 189.850 57.285 190.040 ;
        RECT 58.495 189.870 58.665 190.060 ;
        RECT 58.960 189.870 59.130 190.060 ;
        RECT 60.795 189.850 60.965 190.040 ;
        RECT 63.555 189.870 63.725 190.060 ;
        RECT 64.935 189.905 65.095 190.015 ;
        RECT 66.315 189.850 66.485 190.040 ;
        RECT 66.775 189.850 66.945 190.040 ;
        RECT 69.535 189.850 69.705 190.060 ;
        RECT 69.995 189.850 70.165 190.040 ;
        RECT 72.295 189.895 72.455 190.005 ;
        RECT 73.215 189.870 73.385 190.060 ;
        RECT 74.595 189.870 74.765 190.060 ;
        RECT 76.160 189.850 76.330 190.040 ;
        RECT 80.115 189.870 80.285 190.060 ;
        RECT 80.575 189.870 80.745 190.060 ;
        RECT 81.955 189.870 82.125 190.060 ;
        RECT 84.255 189.870 84.425 190.060 ;
        RECT 86.555 189.850 86.725 190.040 ;
        RECT 87.935 189.850 88.105 190.060 ;
        RECT 88.395 189.870 88.565 190.060 ;
        RECT 91.800 189.850 91.970 190.040 ;
        RECT 93.455 189.850 93.625 190.060 ;
        RECT 94.375 189.895 94.535 190.015 ;
        RECT 94.835 189.850 95.005 190.060 ;
        RECT 101.920 189.850 102.090 190.040 ;
        RECT 103.170 189.900 103.290 190.010 ;
        RECT 103.575 189.850 103.745 190.040 ;
        RECT 107.255 189.870 107.425 190.060 ;
        RECT 109.095 189.870 109.265 190.060 ;
        RECT 109.555 189.870 109.725 190.060 ;
        RECT 113.695 189.850 113.865 190.040 ;
        RECT 114.155 190.010 114.325 190.060 ;
        RECT 114.155 189.900 114.330 190.010 ;
        RECT 114.155 189.870 114.325 189.900 ;
        RECT 115.535 189.850 115.705 190.060 ;
        RECT 10.515 189.040 11.885 189.850 ;
        RECT 12.815 189.040 18.325 189.850 ;
        RECT 18.335 189.040 23.845 189.850 ;
        RECT 23.865 188.940 25.215 189.850 ;
        RECT 25.245 188.980 25.675 189.765 ;
        RECT 26.845 189.170 30.745 189.850 ;
        RECT 29.815 188.940 30.745 189.170 ;
        RECT 31.225 188.940 32.575 189.850 ;
        RECT 32.690 189.170 36.155 189.850 ;
        RECT 36.275 189.170 40.175 189.850 ;
        RECT 40.415 189.170 49.605 189.850 ;
        RECT 32.690 188.940 33.610 189.170 ;
        RECT 36.275 188.940 37.205 189.170 ;
        RECT 40.415 188.940 41.335 189.170 ;
        RECT 44.165 188.950 45.095 189.170 ;
        RECT 49.615 189.070 50.985 189.850 ;
        RECT 51.005 188.980 51.435 189.765 ;
        RECT 51.915 189.040 54.665 189.850 ;
        RECT 54.675 189.070 56.045 189.850 ;
        RECT 56.055 189.040 57.425 189.850 ;
        RECT 57.435 189.040 61.105 189.850 ;
        RECT 61.115 189.040 66.625 189.850 ;
        RECT 66.635 189.170 68.465 189.850 ;
        RECT 68.475 189.040 69.845 189.850 ;
        RECT 69.855 189.170 71.685 189.850 ;
        RECT 72.845 189.170 76.745 189.850 ;
        RECT 75.815 188.940 76.745 189.170 ;
        RECT 76.765 188.980 77.195 189.765 ;
        RECT 77.585 189.170 86.865 189.850 ;
        RECT 77.585 189.050 79.920 189.170 ;
        RECT 77.585 188.940 78.505 189.050 ;
        RECT 84.585 188.950 85.505 189.170 ;
        RECT 86.875 189.040 88.245 189.850 ;
        RECT 88.485 189.170 92.385 189.850 ;
        RECT 91.455 188.940 92.385 189.170 ;
        RECT 92.395 189.070 93.765 189.850 ;
        RECT 94.805 189.170 98.270 189.850 ;
        RECT 98.605 189.170 102.505 189.850 ;
        RECT 97.350 188.940 98.270 189.170 ;
        RECT 101.575 188.940 102.505 189.170 ;
        RECT 102.525 188.980 102.955 189.765 ;
        RECT 103.445 188.940 104.795 189.850 ;
        RECT 104.815 189.170 114.005 189.850 ;
        RECT 104.815 188.940 105.735 189.170 ;
        RECT 108.565 188.950 109.495 189.170 ;
        RECT 114.475 189.040 115.845 189.850 ;
      LAYER nwell ;
        RECT 10.320 185.820 116.040 188.650 ;
      LAYER pwell ;
        RECT 10.515 184.620 11.885 185.430 ;
        RECT 12.365 184.705 12.795 185.490 ;
        RECT 12.815 184.620 14.185 185.430 ;
        RECT 14.195 184.620 19.705 185.430 ;
        RECT 19.715 185.300 20.635 185.530 ;
        RECT 23.465 185.300 24.395 185.520 ;
        RECT 28.915 185.300 29.835 185.530 ;
        RECT 32.665 185.300 33.595 185.520 ;
        RECT 19.715 184.620 28.905 185.300 ;
        RECT 28.915 184.620 38.105 185.300 ;
        RECT 38.125 184.705 38.555 185.490 ;
        RECT 39.035 185.300 39.955 185.530 ;
        RECT 42.785 185.300 43.715 185.520 ;
        RECT 39.035 184.620 48.225 185.300 ;
        RECT 48.245 184.620 49.595 185.530 ;
        RECT 49.615 185.300 50.535 185.530 ;
        RECT 53.365 185.300 54.295 185.520 ;
        RECT 49.615 184.620 58.805 185.300 ;
        RECT 58.815 184.620 60.645 185.430 ;
        RECT 60.895 184.850 63.650 185.530 ;
        RECT 60.895 184.620 63.165 184.850 ;
        RECT 63.885 184.705 64.315 185.490 ;
        RECT 64.335 184.620 66.165 185.430 ;
        RECT 66.175 184.620 71.685 185.430 ;
        RECT 71.705 184.620 73.055 185.530 ;
        RECT 73.445 185.420 74.365 185.530 ;
        RECT 73.445 185.300 75.780 185.420 ;
        RECT 80.445 185.300 81.365 185.520 ;
        RECT 73.445 184.620 82.725 185.300 ;
        RECT 82.735 184.620 88.245 185.430 ;
        RECT 88.265 184.620 89.615 185.530 ;
        RECT 89.645 184.705 90.075 185.490 ;
        RECT 94.605 185.300 95.535 185.520 ;
        RECT 98.365 185.300 99.285 185.530 ;
        RECT 90.095 184.620 99.285 185.300 ;
        RECT 99.295 184.620 101.125 185.430 ;
        RECT 101.135 184.620 102.505 185.400 ;
        RECT 105.715 185.300 106.645 185.530 ;
        RECT 102.745 184.620 106.645 185.300 ;
        RECT 106.750 185.300 107.670 185.530 ;
        RECT 106.750 184.620 110.215 185.300 ;
        RECT 110.795 184.620 114.465 185.430 ;
        RECT 114.475 184.620 115.845 185.430 ;
        RECT 10.655 184.410 10.825 184.620 ;
        RECT 12.090 184.460 12.210 184.570 ;
        RECT 13.875 184.410 14.045 184.620 ;
        RECT 19.395 184.410 19.565 184.620 ;
        RECT 24.915 184.410 25.085 184.600 ;
        RECT 26.755 184.410 26.925 184.600 ;
        RECT 28.135 184.410 28.305 184.600 ;
        RECT 28.595 184.410 28.765 184.620 ;
        RECT 30.895 184.410 31.065 184.600 ;
        RECT 32.735 184.410 32.905 184.600 ;
        RECT 33.195 184.410 33.365 184.600 ;
        RECT 34.575 184.410 34.745 184.600 ;
        RECT 37.795 184.430 37.965 184.620 ;
        RECT 38.770 184.460 38.890 184.570 ;
        RECT 41.660 184.410 41.830 184.600 ;
        RECT 45.800 184.410 45.970 184.600 ;
        RECT 46.590 184.460 46.710 184.570 ;
        RECT 47.915 184.430 48.085 184.620 ;
        RECT 48.375 184.430 48.545 184.620 ;
        RECT 50.400 184.410 50.570 184.600 ;
        RECT 51.595 184.410 51.765 184.600 ;
        RECT 53.435 184.455 53.595 184.565 ;
        RECT 57.115 184.410 57.285 184.600 ;
        RECT 57.575 184.430 57.745 184.600 ;
        RECT 58.495 184.430 58.665 184.620 ;
        RECT 60.335 184.430 60.505 184.620 ;
        RECT 60.895 184.600 60.965 184.620 ;
        RECT 60.795 184.430 60.965 184.600 ;
        RECT 57.675 184.410 57.745 184.430 ;
        RECT 65.855 184.410 66.025 184.620 ;
        RECT 70.455 184.410 70.625 184.600 ;
        RECT 71.375 184.430 71.545 184.620 ;
        RECT 72.295 184.410 72.465 184.600 ;
        RECT 72.755 184.430 72.925 184.620 ;
        RECT 76.160 184.410 76.330 184.600 ;
        RECT 77.360 184.410 77.530 184.600 ;
        RECT 80.115 184.410 80.285 184.600 ;
        RECT 82.415 184.430 82.585 184.620 ;
        RECT 83.795 184.410 83.965 184.600 ;
        RECT 87.935 184.430 88.105 184.620 ;
        RECT 88.395 184.430 88.565 184.620 ;
        RECT 90.235 184.430 90.405 184.620 ;
        RECT 92.995 184.410 93.165 184.600 ;
        RECT 96.860 184.410 97.030 184.600 ;
        RECT 98.055 184.455 98.215 184.565 ;
        RECT 100.815 184.430 100.985 184.620 ;
        RECT 101.275 184.430 101.445 184.620 ;
        RECT 101.920 184.410 102.090 184.600 ;
        RECT 104.035 184.410 104.205 184.600 ;
        RECT 104.955 184.455 105.115 184.565 ;
        RECT 106.060 184.430 106.230 184.620 ;
        RECT 110.015 184.430 110.185 184.620 ;
        RECT 110.530 184.460 110.650 184.570 ;
        RECT 114.155 184.410 114.325 184.620 ;
        RECT 115.535 184.410 115.705 184.620 ;
        RECT 10.515 183.600 11.885 184.410 ;
        RECT 12.355 183.600 14.185 184.410 ;
        RECT 14.195 183.600 19.705 184.410 ;
        RECT 19.715 183.600 25.225 184.410 ;
        RECT 25.245 183.540 25.675 184.325 ;
        RECT 25.705 183.500 27.055 184.410 ;
        RECT 27.075 183.600 28.445 184.410 ;
        RECT 28.455 183.630 29.825 184.410 ;
        RECT 29.835 183.630 31.205 184.410 ;
        RECT 31.215 183.600 33.045 184.410 ;
        RECT 33.055 183.630 34.425 184.410 ;
        RECT 34.545 183.730 38.010 184.410 ;
        RECT 38.345 183.730 42.245 184.410 ;
        RECT 42.485 183.730 46.385 184.410 ;
        RECT 47.085 183.730 50.985 184.410 ;
        RECT 37.090 183.500 38.010 183.730 ;
        RECT 41.315 183.500 42.245 183.730 ;
        RECT 45.455 183.500 46.385 183.730 ;
        RECT 50.055 183.500 50.985 183.730 ;
        RECT 51.005 183.540 51.435 184.325 ;
        RECT 51.455 183.630 52.825 184.410 ;
        RECT 53.755 183.600 57.425 184.410 ;
        RECT 57.675 184.180 59.945 184.410 ;
        RECT 61.740 184.180 66.165 184.410 ;
        RECT 66.185 184.370 67.105 184.410 ;
        RECT 57.675 183.500 60.430 184.180 ;
        RECT 60.800 183.500 66.165 184.180 ;
        RECT 66.175 184.180 67.105 184.370 ;
        RECT 69.195 184.180 70.765 184.410 ;
        RECT 66.175 183.820 70.765 184.180 ;
        RECT 66.185 183.730 70.765 183.820 ;
        RECT 66.185 183.500 69.185 183.730 ;
        RECT 70.775 183.600 72.605 184.410 ;
        RECT 72.845 183.730 76.745 184.410 ;
        RECT 75.815 183.500 76.745 183.730 ;
        RECT 76.765 183.540 77.195 184.325 ;
        RECT 77.215 183.500 79.825 184.410 ;
        RECT 79.975 183.630 81.345 184.410 ;
        RECT 81.365 183.730 84.105 184.410 ;
        RECT 84.115 183.730 93.305 184.410 ;
        RECT 93.545 183.730 97.445 184.410 ;
        RECT 98.605 183.730 102.505 184.410 ;
        RECT 84.115 183.500 85.035 183.730 ;
        RECT 87.865 183.510 88.795 183.730 ;
        RECT 96.515 183.500 97.445 183.730 ;
        RECT 101.575 183.500 102.505 183.730 ;
        RECT 102.525 183.540 102.955 184.325 ;
        RECT 102.985 183.500 104.335 184.410 ;
        RECT 105.275 183.730 114.465 184.410 ;
        RECT 105.275 183.500 106.195 183.730 ;
        RECT 109.025 183.510 109.955 183.730 ;
        RECT 114.475 183.600 115.845 184.410 ;
      LAYER nwell ;
        RECT 10.320 180.380 116.040 183.210 ;
      LAYER pwell ;
        RECT 10.515 179.180 11.885 179.990 ;
        RECT 12.365 179.265 12.795 180.050 ;
        RECT 12.815 179.180 14.185 179.990 ;
        RECT 14.195 179.180 19.705 179.990 ;
        RECT 22.370 179.860 23.290 180.090 ;
        RECT 26.050 179.860 26.970 180.090 ;
        RECT 30.275 179.860 31.205 180.090 ;
        RECT 19.825 179.180 23.290 179.860 ;
        RECT 23.505 179.180 26.970 179.860 ;
        RECT 27.305 179.180 31.205 179.860 ;
        RECT 31.215 179.180 32.585 179.960 ;
        RECT 32.595 179.180 34.425 179.990 ;
        RECT 34.630 179.180 38.105 180.090 ;
        RECT 38.125 179.265 38.555 180.050 ;
        RECT 38.575 179.180 39.945 179.990 ;
        RECT 39.965 179.180 41.315 180.090 ;
        RECT 43.990 179.860 44.910 180.090 ;
        RECT 41.445 179.180 44.910 179.860 ;
        RECT 45.475 179.860 46.395 180.090 ;
        RECT 49.225 179.860 50.155 180.080 ;
        RECT 45.475 179.180 54.665 179.860 ;
        RECT 55.595 179.180 59.265 179.990 ;
        RECT 59.285 179.180 60.635 180.090 ;
        RECT 60.870 179.410 63.625 180.090 ;
        RECT 61.355 179.180 63.625 179.410 ;
        RECT 63.885 179.265 64.315 180.050 ;
        RECT 64.335 179.180 65.705 179.990 ;
        RECT 65.715 179.180 69.385 179.990 ;
        RECT 69.395 179.180 72.135 179.860 ;
        RECT 72.615 179.180 74.445 179.990 ;
        RECT 74.455 179.860 75.375 180.090 ;
        RECT 78.205 179.860 79.135 180.080 ;
        RECT 74.455 179.180 83.645 179.860 ;
        RECT 83.655 179.180 85.025 179.960 ;
        RECT 86.050 179.860 86.970 180.090 ;
        RECT 86.050 179.180 89.515 179.860 ;
        RECT 89.645 179.265 90.075 180.050 ;
        RECT 90.105 179.180 91.455 180.090 ;
        RECT 91.475 179.180 92.845 179.960 ;
        RECT 92.950 179.860 93.870 180.090 ;
        RECT 92.950 179.180 96.415 179.860 ;
        RECT 96.995 179.180 98.825 179.990 ;
        RECT 98.835 179.860 99.755 180.090 ;
        RECT 102.585 179.860 103.515 180.080 ;
        RECT 98.835 179.180 108.025 179.860 ;
        RECT 108.045 179.180 109.395 180.090 ;
        RECT 110.335 179.180 111.705 179.960 ;
        RECT 111.715 179.180 114.465 179.990 ;
        RECT 114.475 179.180 115.845 179.990 ;
        RECT 10.655 178.970 10.825 179.180 ;
        RECT 12.090 179.020 12.210 179.130 ;
        RECT 13.875 178.990 14.045 179.180 ;
        RECT 15.255 178.970 15.425 179.160 ;
        RECT 15.715 178.970 15.885 179.160 ;
        RECT 19.395 179.130 19.565 179.180 ;
        RECT 19.395 179.020 19.570 179.130 ;
        RECT 19.395 178.990 19.565 179.020 ;
        RECT 19.855 178.990 20.025 179.180 ;
        RECT 20.775 178.970 20.945 179.160 ;
        RECT 23.535 178.990 23.705 179.180 ;
        RECT 30.620 179.160 30.790 179.180 ;
        RECT 24.640 178.970 24.810 179.160 ;
        RECT 26.295 179.015 26.455 179.125 ;
        RECT 29.970 178.970 30.140 179.160 ;
        RECT 30.620 178.990 30.880 179.160 ;
        RECT 31.355 178.990 31.525 179.180 ;
        RECT 34.115 178.990 34.285 179.180 ;
        RECT 30.710 178.970 30.880 178.990 ;
        RECT 35.495 178.970 35.665 179.160 ;
        RECT 37.790 178.990 37.960 179.180 ;
        RECT 39.170 178.970 39.340 179.160 ;
        RECT 39.635 178.990 39.805 179.180 ;
        RECT 41.015 178.990 41.185 179.180 ;
        RECT 41.475 178.990 41.645 179.180 ;
        RECT 42.850 178.970 43.020 179.160 ;
        RECT 43.315 178.970 43.485 179.160 ;
        RECT 45.210 179.020 45.330 179.130 ;
        RECT 50.400 178.970 50.570 179.160 ;
        RECT 54.355 178.990 54.525 179.180 ;
        RECT 54.815 178.970 54.985 179.160 ;
        RECT 55.275 179.025 55.435 179.135 ;
        RECT 57.575 178.970 57.745 179.160 ;
        RECT 58.040 178.970 58.210 179.160 ;
        RECT 58.955 178.990 59.125 179.180 ;
        RECT 59.415 178.990 59.585 179.180 ;
        RECT 63.555 179.160 63.625 179.180 ;
        RECT 60.795 178.970 60.965 179.160 ;
        RECT 62.635 178.970 62.805 179.160 ;
        RECT 63.555 178.990 63.725 179.160 ;
        RECT 64.475 178.970 64.645 179.160 ;
        RECT 65.395 178.990 65.565 179.180 ;
        RECT 67.235 178.970 67.405 179.160 ;
        RECT 69.075 178.970 69.245 179.180 ;
        RECT 69.535 178.990 69.705 179.180 ;
        RECT 72.350 179.020 72.470 179.130 ;
        RECT 74.135 178.990 74.305 179.180 ;
        RECT 76.160 178.970 76.330 179.160 ;
        RECT 77.355 178.970 77.525 179.160 ;
        RECT 81.955 178.970 82.125 179.160 ;
        RECT 82.875 179.015 83.035 179.125 ;
        RECT 83.335 178.970 83.505 179.180 ;
        RECT 84.715 178.990 84.885 179.180 ;
        RECT 85.635 179.025 85.795 179.135 ;
        RECT 87.290 178.970 87.460 179.160 ;
        RECT 89.315 178.990 89.485 179.180 ;
        RECT 91.155 178.970 91.325 179.180 ;
        RECT 92.535 178.990 92.705 179.180 ;
        RECT 94.840 178.970 95.010 179.160 ;
        RECT 96.215 178.990 96.385 179.180 ;
        RECT 98.515 179.160 98.685 179.180 ;
        RECT 96.730 179.020 96.850 179.130 ;
        RECT 98.515 178.990 98.690 179.160 ;
        RECT 102.250 179.020 102.370 179.130 ;
        RECT 103.575 179.015 103.735 179.125 ;
        RECT 98.520 178.970 98.690 178.990 ;
        RECT 107.440 178.970 107.610 179.160 ;
        RECT 107.715 178.990 107.885 179.180 ;
        RECT 108.175 178.970 108.345 179.180 ;
        RECT 110.015 179.025 110.175 179.135 ;
        RECT 110.475 178.990 110.645 179.180 ;
        RECT 114.155 178.970 114.325 179.180 ;
        RECT 115.535 178.970 115.705 179.180 ;
        RECT 10.515 178.160 11.885 178.970 ;
        RECT 11.895 178.160 15.565 178.970 ;
        RECT 15.685 178.290 19.150 178.970 ;
        RECT 18.230 178.060 19.150 178.290 ;
        RECT 19.725 178.060 21.075 178.970 ;
        RECT 21.325 178.290 25.225 178.970 ;
        RECT 24.295 178.060 25.225 178.290 ;
        RECT 25.245 178.100 25.675 178.885 ;
        RECT 26.810 178.060 30.285 178.970 ;
        RECT 30.295 178.290 34.195 178.970 ;
        RECT 30.295 178.060 31.225 178.290 ;
        RECT 34.435 178.160 35.805 178.970 ;
        RECT 36.010 178.060 39.485 178.970 ;
        RECT 39.690 178.060 43.165 178.970 ;
        RECT 43.285 178.290 46.750 178.970 ;
        RECT 47.085 178.290 50.985 178.970 ;
        RECT 45.830 178.060 46.750 178.290 ;
        RECT 50.055 178.060 50.985 178.290 ;
        RECT 51.005 178.100 51.435 178.885 ;
        RECT 51.550 178.290 55.015 178.970 ;
        RECT 55.145 178.290 57.885 178.970 ;
        RECT 51.550 178.060 52.470 178.290 ;
        RECT 57.895 178.060 60.505 178.970 ;
        RECT 60.655 178.290 62.485 178.970 ;
        RECT 62.495 178.290 64.325 178.970 ;
        RECT 61.140 178.060 62.485 178.290 ;
        RECT 62.980 178.060 64.325 178.290 ;
        RECT 64.335 178.060 67.055 178.970 ;
        RECT 67.095 178.290 68.925 178.970 ;
        RECT 69.045 178.290 72.510 178.970 ;
        RECT 72.845 178.290 76.745 178.970 ;
        RECT 67.580 178.060 68.925 178.290 ;
        RECT 71.590 178.060 72.510 178.290 ;
        RECT 75.815 178.060 76.745 178.290 ;
        RECT 76.765 178.100 77.195 178.885 ;
        RECT 77.325 178.290 80.790 178.970 ;
        RECT 79.870 178.060 80.790 178.290 ;
        RECT 80.905 178.060 82.255 178.970 ;
        RECT 83.305 178.290 86.770 178.970 ;
        RECT 85.850 178.060 86.770 178.290 ;
        RECT 86.875 178.290 90.775 178.970 ;
        RECT 91.125 178.290 94.590 178.970 ;
        RECT 86.875 178.060 87.805 178.290 ;
        RECT 93.670 178.060 94.590 178.290 ;
        RECT 94.695 178.060 98.170 178.970 ;
        RECT 98.375 178.060 101.850 178.970 ;
        RECT 102.525 178.100 102.955 178.885 ;
        RECT 104.125 178.290 108.025 178.970 ;
        RECT 108.145 178.290 111.610 178.970 ;
        RECT 107.095 178.060 108.025 178.290 ;
        RECT 110.690 178.060 111.610 178.290 ;
        RECT 111.715 178.160 114.465 178.970 ;
        RECT 114.475 178.160 115.845 178.970 ;
      LAYER nwell ;
        RECT 10.320 174.940 116.040 177.770 ;
      LAYER pwell ;
        RECT 10.515 173.740 11.885 174.550 ;
        RECT 12.365 173.825 12.795 174.610 ;
        RECT 13.275 173.740 15.105 174.550 ;
        RECT 15.115 174.420 16.035 174.650 ;
        RECT 18.865 174.420 19.795 174.640 ;
        RECT 24.315 174.420 25.235 174.650 ;
        RECT 28.065 174.420 28.995 174.640 ;
        RECT 15.115 173.740 24.305 174.420 ;
        RECT 24.315 173.740 33.505 174.420 ;
        RECT 34.630 173.740 38.105 174.650 ;
        RECT 38.125 173.825 38.555 174.610 ;
        RECT 39.230 173.740 42.705 174.650 ;
        RECT 42.715 173.740 46.190 174.650 ;
        RECT 49.050 174.420 49.970 174.650 ;
        RECT 54.195 174.420 55.125 174.650 ;
        RECT 46.505 173.740 49.970 174.420 ;
        RECT 51.225 173.740 55.125 174.420 ;
        RECT 55.145 173.740 56.495 174.650 ;
        RECT 56.515 173.740 57.885 174.520 ;
        RECT 58.355 173.740 60.185 174.550 ;
        RECT 60.195 174.420 61.540 174.650 ;
        RECT 62.035 174.420 63.380 174.650 ;
        RECT 60.195 173.740 62.025 174.420 ;
        RECT 62.035 173.740 63.865 174.420 ;
        RECT 63.885 173.825 64.315 174.610 ;
        RECT 64.335 173.740 66.165 174.550 ;
        RECT 66.175 173.740 69.650 174.650 ;
        RECT 69.855 173.740 73.330 174.650 ;
        RECT 73.535 173.740 77.010 174.650 ;
        RECT 78.135 173.740 87.240 174.420 ;
        RECT 88.255 173.740 89.625 174.520 ;
        RECT 89.645 173.825 90.075 174.610 ;
        RECT 90.095 173.740 93.570 174.650 ;
        RECT 94.890 173.740 98.365 174.650 ;
        RECT 98.375 173.740 101.125 174.550 ;
        RECT 103.790 174.420 104.710 174.650 ;
        RECT 101.245 173.740 104.710 174.420 ;
        RECT 104.815 173.740 108.290 174.650 ;
        RECT 108.690 173.740 112.165 174.650 ;
        RECT 112.175 173.740 113.545 174.520 ;
        RECT 114.475 173.740 115.845 174.550 ;
        RECT 10.655 173.530 10.825 173.740 ;
        RECT 12.090 173.580 12.210 173.690 ;
        RECT 13.010 173.580 13.130 173.690 ;
        RECT 14.335 173.530 14.505 173.720 ;
        RECT 14.795 173.550 14.965 173.740 ;
        RECT 19.855 173.530 20.025 173.720 ;
        RECT 21.235 173.530 21.405 173.720 ;
        RECT 23.995 173.550 24.165 173.740 ;
        RECT 24.915 173.530 25.085 173.720 ;
        RECT 26.755 173.530 26.925 173.720 ;
        RECT 28.135 173.530 28.305 173.720 ;
        RECT 28.650 173.580 28.770 173.690 ;
        RECT 32.270 173.530 32.440 173.720 ;
        RECT 32.740 173.530 32.910 173.720 ;
        RECT 33.195 173.550 33.365 173.740 ;
        RECT 37.790 173.720 37.960 173.740 ;
        RECT 34.115 173.585 34.275 173.695 ;
        RECT 37.335 173.530 37.505 173.720 ;
        RECT 37.790 173.550 37.970 173.720 ;
        RECT 38.770 173.580 38.890 173.690 ;
        RECT 42.390 173.550 42.560 173.740 ;
        RECT 42.860 173.550 43.030 173.740 ;
        RECT 46.535 173.550 46.705 173.740 ;
        RECT 37.800 173.530 37.970 173.550 ;
        RECT 50.215 173.530 50.385 173.720 ;
        RECT 50.675 173.690 50.835 173.695 ;
        RECT 50.675 173.585 50.850 173.690 ;
        RECT 50.730 173.580 50.850 173.585 ;
        RECT 54.540 173.550 54.710 173.740 ;
        RECT 56.195 173.550 56.365 173.740 ;
        RECT 56.655 173.550 56.825 173.740 ;
        RECT 58.090 173.580 58.210 173.690 ;
        RECT 59.875 173.550 60.045 173.740 ;
        RECT 60.335 173.530 60.505 173.720 ;
        RECT 61.255 173.575 61.415 173.685 ;
        RECT 61.715 173.550 61.885 173.740 ;
        RECT 63.555 173.550 63.725 173.740 ;
        RECT 64.935 173.530 65.105 173.720 ;
        RECT 65.855 173.550 66.025 173.740 ;
        RECT 66.320 173.550 66.490 173.740 ;
        RECT 70.000 173.550 70.170 173.740 ;
        RECT 70.455 173.530 70.625 173.720 ;
        RECT 70.920 173.530 71.090 173.720 ;
        RECT 73.680 173.550 73.850 173.740 ;
        RECT 74.650 173.580 74.770 173.690 ;
        RECT 76.435 173.530 76.605 173.720 ;
        RECT 77.410 173.580 77.530 173.690 ;
        RECT 77.815 173.585 77.975 173.695 ;
        RECT 78.275 173.550 78.445 173.740 ;
        RECT 81.035 173.530 81.205 173.720 ;
        RECT 81.495 173.530 81.665 173.720 ;
        RECT 82.875 173.530 83.045 173.720 ;
        RECT 87.935 173.585 88.095 173.695 ;
        RECT 88.395 173.550 88.565 173.740 ;
        RECT 90.240 173.550 90.410 173.740 ;
        RECT 98.050 173.720 98.220 173.740 ;
        RECT 94.375 173.585 94.535 173.695 ;
        RECT 95.295 173.530 95.465 173.720 ;
        RECT 98.050 173.550 98.225 173.720 ;
        RECT 100.815 173.550 100.985 173.740 ;
        RECT 101.275 173.550 101.445 173.740 ;
        RECT 98.055 173.530 98.225 173.550 ;
        RECT 101.920 173.530 102.090 173.720 ;
        RECT 103.115 173.530 103.285 173.720 ;
        RECT 104.960 173.550 105.130 173.740 ;
        RECT 111.850 173.550 112.020 173.740 ;
        RECT 113.235 173.530 113.405 173.740 ;
        RECT 114.155 173.575 114.315 173.695 ;
        RECT 115.535 173.530 115.705 173.740 ;
        RECT 10.515 172.720 11.885 173.530 ;
        RECT 11.895 172.720 14.645 173.530 ;
        RECT 14.655 172.720 20.165 173.530 ;
        RECT 20.185 172.620 21.535 173.530 ;
        RECT 21.650 172.850 25.115 173.530 ;
        RECT 21.650 172.620 22.570 172.850 ;
        RECT 25.245 172.660 25.675 173.445 ;
        RECT 25.695 172.720 27.065 173.530 ;
        RECT 27.075 172.750 28.445 173.530 ;
        RECT 29.110 172.620 32.585 173.530 ;
        RECT 32.595 172.620 36.070 173.530 ;
        RECT 36.275 172.720 37.645 173.530 ;
        RECT 37.655 172.620 41.130 173.530 ;
        RECT 41.420 172.850 50.525 173.530 ;
        RECT 51.005 172.660 51.435 173.445 ;
        RECT 51.455 172.850 60.645 173.530 ;
        RECT 51.455 172.620 52.375 172.850 ;
        RECT 55.205 172.630 56.135 172.850 ;
        RECT 61.575 172.720 65.245 173.530 ;
        RECT 65.255 172.720 70.765 173.530 ;
        RECT 70.775 172.620 74.250 173.530 ;
        RECT 74.915 172.720 76.745 173.530 ;
        RECT 76.765 172.660 77.195 173.445 ;
        RECT 77.675 172.720 81.345 173.530 ;
        RECT 81.365 172.620 82.715 173.530 ;
        RECT 82.735 172.850 91.925 173.530 ;
        RECT 87.245 172.630 88.175 172.850 ;
        RECT 91.005 172.620 91.925 172.850 ;
        RECT 92.030 172.850 95.495 173.530 ;
        RECT 92.030 172.620 92.950 172.850 ;
        RECT 95.615 172.720 98.365 173.530 ;
        RECT 98.605 172.850 102.505 173.530 ;
        RECT 101.575 172.620 102.505 172.850 ;
        RECT 102.525 172.660 102.955 173.445 ;
        RECT 102.985 172.620 104.335 173.530 ;
        RECT 104.355 172.850 113.545 173.530 ;
        RECT 104.355 172.620 105.275 172.850 ;
        RECT 108.105 172.630 109.035 172.850 ;
        RECT 114.475 172.720 115.845 173.530 ;
      LAYER nwell ;
        RECT 10.320 169.500 116.040 172.330 ;
      LAYER pwell ;
        RECT 10.515 168.300 11.885 169.110 ;
        RECT 12.365 168.385 12.795 169.170 ;
        RECT 13.275 168.300 16.025 169.110 ;
        RECT 16.035 168.300 21.545 169.110 ;
        RECT 21.640 168.300 30.745 168.980 ;
        RECT 31.685 168.300 33.035 169.210 ;
        RECT 33.515 168.300 36.265 169.110 ;
        RECT 36.285 168.300 37.635 169.210 ;
        RECT 38.125 168.385 38.555 169.170 ;
        RECT 39.035 168.300 41.785 169.110 ;
        RECT 41.890 168.980 42.810 169.210 ;
        RECT 47.315 168.980 48.235 169.210 ;
        RECT 51.065 168.980 51.995 169.200 ;
        RECT 41.890 168.300 45.355 168.980 ;
        RECT 45.475 168.300 46.840 168.980 ;
        RECT 47.315 168.300 56.505 168.980 ;
        RECT 56.515 168.300 60.185 169.110 ;
        RECT 60.195 168.980 61.540 169.210 ;
        RECT 62.035 168.980 63.380 169.210 ;
        RECT 60.195 168.300 62.025 168.980 ;
        RECT 62.035 168.300 63.865 168.980 ;
        RECT 63.885 168.385 64.315 169.170 ;
        RECT 65.255 168.300 70.765 169.110 ;
        RECT 71.145 169.100 72.065 169.210 ;
        RECT 71.145 168.980 73.480 169.100 ;
        RECT 78.145 168.980 79.065 169.200 ;
        RECT 71.145 168.300 80.425 168.980 ;
        RECT 80.435 168.300 83.185 169.110 ;
        RECT 86.395 168.980 87.325 169.210 ;
        RECT 83.425 168.300 87.325 168.980 ;
        RECT 87.795 168.300 89.165 169.080 ;
        RECT 89.645 168.385 90.075 169.170 ;
        RECT 90.095 168.300 92.845 169.110 ;
        RECT 92.865 168.300 94.215 169.210 ;
        RECT 96.890 168.980 97.810 169.210 ;
        RECT 94.345 168.300 97.810 168.980 ;
        RECT 97.915 168.300 107.020 168.980 ;
        RECT 107.775 168.300 109.865 169.110 ;
        RECT 109.875 168.300 111.705 168.980 ;
        RECT 111.715 168.300 114.465 169.110 ;
        RECT 114.475 168.300 115.845 169.110 ;
        RECT 10.655 168.090 10.825 168.300 ;
        RECT 12.090 168.140 12.210 168.250 ;
        RECT 13.010 168.140 13.130 168.250 ;
        RECT 13.875 168.090 14.045 168.280 ;
        RECT 15.715 168.110 15.885 168.300 ;
        RECT 19.395 168.090 19.565 168.280 ;
        RECT 20.775 168.090 20.945 168.280 ;
        RECT 21.235 168.090 21.405 168.300 ;
        RECT 22.615 168.090 22.785 168.280 ;
        RECT 23.995 168.090 24.165 168.280 ;
        RECT 26.295 168.135 26.455 168.245 ;
        RECT 26.755 168.090 26.925 168.280 ;
        RECT 30.435 168.090 30.605 168.300 ;
        RECT 31.355 168.145 31.515 168.255 ;
        RECT 32.735 168.110 32.905 168.300 ;
        RECT 33.250 168.140 33.370 168.250 ;
        RECT 34.115 168.090 34.285 168.280 ;
        RECT 35.955 168.110 36.125 168.300 ;
        RECT 36.415 168.110 36.585 168.300 ;
        RECT 37.850 168.140 37.970 168.250 ;
        RECT 38.770 168.140 38.890 168.250 ;
        RECT 41.475 168.110 41.645 168.300 ;
        RECT 45.155 168.110 45.325 168.300 ;
        RECT 46.535 168.090 46.705 168.280 ;
        RECT 46.995 168.110 47.165 168.280 ;
        RECT 49.295 168.090 49.465 168.280 ;
        RECT 49.755 168.090 49.925 168.280 ;
        RECT 52.975 168.090 53.145 168.280 ;
        RECT 55.730 168.090 55.900 168.280 ;
        RECT 56.195 168.110 56.365 168.300 ;
        RECT 56.655 168.135 56.815 168.245 ;
        RECT 59.875 168.110 60.045 168.300 ;
        RECT 60.335 168.090 60.505 168.280 ;
        RECT 60.795 168.090 60.965 168.280 ;
        RECT 61.715 168.110 61.885 168.300 ;
        RECT 63.555 168.090 63.725 168.300 ;
        RECT 64.935 168.145 65.095 168.255 ;
        RECT 69.720 168.090 69.890 168.280 ;
        RECT 70.455 168.110 70.625 168.300 ;
        RECT 73.860 168.090 74.030 168.280 ;
        RECT 74.650 168.140 74.770 168.250 ;
        RECT 75.975 168.090 76.145 168.280 ;
        RECT 76.490 168.140 76.610 168.250 ;
        RECT 77.355 168.090 77.525 168.280 ;
        RECT 78.790 168.140 78.910 168.250 ;
        RECT 80.115 168.110 80.285 168.300 ;
        RECT 81.495 168.090 81.665 168.280 ;
        RECT 82.875 168.110 83.045 168.300 ;
        RECT 86.740 168.110 86.910 168.300 ;
        RECT 87.015 168.090 87.185 168.280 ;
        RECT 87.475 168.250 87.645 168.280 ;
        RECT 87.475 168.140 87.650 168.250 ;
        RECT 87.475 168.090 87.645 168.140 ;
        RECT 88.855 168.090 89.025 168.300 ;
        RECT 89.370 168.140 89.490 168.250 ;
        RECT 92.535 168.110 92.705 168.300 ;
        RECT 92.995 168.110 93.165 168.300 ;
        RECT 94.375 168.110 94.545 168.300 ;
        RECT 98.055 168.110 98.225 168.300 ;
        RECT 101.275 168.090 101.445 168.280 ;
        RECT 102.195 168.135 102.355 168.245 ;
        RECT 103.170 168.140 103.290 168.250 ;
        RECT 103.575 168.090 103.745 168.280 ;
        RECT 109.555 168.110 109.725 168.300 ;
        RECT 111.395 168.110 111.565 168.300 ;
        RECT 113.695 168.090 113.865 168.280 ;
        RECT 114.155 168.250 114.325 168.300 ;
        RECT 114.155 168.140 114.330 168.250 ;
        RECT 114.155 168.110 114.325 168.140 ;
        RECT 115.535 168.090 115.705 168.300 ;
        RECT 10.515 167.280 11.885 168.090 ;
        RECT 12.355 167.280 14.185 168.090 ;
        RECT 14.195 167.280 19.705 168.090 ;
        RECT 19.725 167.180 21.075 168.090 ;
        RECT 21.095 167.310 22.465 168.090 ;
        RECT 22.485 167.180 23.835 168.090 ;
        RECT 23.855 167.310 25.225 168.090 ;
        RECT 25.245 167.220 25.675 168.005 ;
        RECT 26.725 167.410 30.190 168.090 ;
        RECT 30.405 167.410 33.870 168.090 ;
        RECT 34.085 167.410 37.550 168.090 ;
        RECT 29.270 167.180 30.190 167.410 ;
        RECT 32.950 167.180 33.870 167.410 ;
        RECT 36.630 167.180 37.550 167.410 ;
        RECT 37.655 167.410 46.845 168.090 ;
        RECT 37.655 167.180 38.575 167.410 ;
        RECT 41.405 167.190 42.335 167.410 ;
        RECT 46.855 167.280 49.605 168.090 ;
        RECT 49.625 167.180 50.975 168.090 ;
        RECT 51.005 167.220 51.435 168.005 ;
        RECT 51.455 167.280 53.285 168.090 ;
        RECT 53.435 167.180 56.045 168.090 ;
        RECT 56.975 167.280 60.645 168.090 ;
        RECT 60.655 167.410 63.395 168.090 ;
        RECT 63.415 167.180 66.135 168.090 ;
        RECT 66.405 167.410 70.305 168.090 ;
        RECT 70.545 167.410 74.445 168.090 ;
        RECT 69.375 167.180 70.305 167.410 ;
        RECT 73.515 167.180 74.445 167.410 ;
        RECT 74.925 167.180 76.275 168.090 ;
        RECT 76.765 167.220 77.195 168.005 ;
        RECT 77.215 167.310 78.585 168.090 ;
        RECT 79.055 167.280 81.805 168.090 ;
        RECT 81.815 167.280 87.325 168.090 ;
        RECT 87.345 167.180 88.695 168.090 ;
        RECT 88.825 167.410 92.290 168.090 ;
        RECT 91.370 167.180 92.290 167.410 ;
        RECT 92.395 167.410 101.585 168.090 ;
        RECT 92.395 167.180 93.315 167.410 ;
        RECT 96.145 167.190 97.075 167.410 ;
        RECT 102.525 167.220 102.955 168.005 ;
        RECT 103.445 167.180 104.795 168.090 ;
        RECT 104.815 167.410 114.005 168.090 ;
        RECT 104.815 167.180 105.735 167.410 ;
        RECT 108.565 167.190 109.495 167.410 ;
        RECT 114.475 167.280 115.845 168.090 ;
      LAYER nwell ;
        RECT 10.320 164.060 116.040 166.890 ;
      LAYER pwell ;
        RECT 10.515 162.860 11.885 163.670 ;
        RECT 12.365 162.945 12.795 163.730 ;
        RECT 12.815 162.860 16.485 163.670 ;
        RECT 16.495 163.540 17.415 163.770 ;
        RECT 20.245 163.540 21.175 163.760 ;
        RECT 16.495 162.860 25.685 163.540 ;
        RECT 26.815 162.860 28.905 163.670 ;
        RECT 28.915 163.540 29.835 163.770 ;
        RECT 32.665 163.540 33.595 163.760 ;
        RECT 28.915 162.860 38.105 163.540 ;
        RECT 38.125 162.945 38.555 163.730 ;
        RECT 38.575 162.860 39.945 163.640 ;
        RECT 39.955 162.860 41.785 163.670 ;
        RECT 44.995 163.540 45.925 163.770 ;
        RECT 49.135 163.540 50.065 163.770 ;
        RECT 42.025 162.860 45.925 163.540 ;
        RECT 46.165 162.860 50.065 163.540 ;
        RECT 50.075 162.860 51.905 163.670 ;
        RECT 51.915 162.860 53.285 163.640 ;
        RECT 54.225 162.860 56.965 163.540 ;
        RECT 57.115 162.860 59.725 163.770 ;
        RECT 59.745 162.860 62.485 163.540 ;
        RECT 62.495 162.860 63.865 163.670 ;
        RECT 63.885 162.945 64.315 163.730 ;
        RECT 64.335 162.860 68.005 163.670 ;
        RECT 68.385 163.660 69.305 163.770 ;
        RECT 68.385 163.540 70.720 163.660 ;
        RECT 75.385 163.540 76.305 163.760 ;
        RECT 68.385 162.860 77.665 163.540 ;
        RECT 77.675 162.860 79.045 163.640 ;
        RECT 79.055 162.860 84.565 163.670 ;
        RECT 87.775 163.540 88.705 163.770 ;
        RECT 84.805 162.860 88.705 163.540 ;
        RECT 89.645 162.945 90.075 163.730 ;
        RECT 94.215 163.540 95.145 163.770 ;
        RECT 91.245 162.860 95.145 163.540 ;
        RECT 95.155 162.860 96.525 163.640 ;
        RECT 96.535 163.540 97.465 163.770 ;
        RECT 96.535 162.860 100.435 163.540 ;
        RECT 101.605 162.860 102.955 163.770 ;
        RECT 102.975 163.540 103.895 163.770 ;
        RECT 106.725 163.540 107.655 163.760 ;
        RECT 102.975 162.860 112.165 163.540 ;
        RECT 112.175 162.860 113.545 163.640 ;
        RECT 114.475 162.860 115.845 163.670 ;
        RECT 10.655 162.650 10.825 162.860 ;
        RECT 12.090 162.700 12.210 162.810 ;
        RECT 14.795 162.650 14.965 162.840 ;
        RECT 15.255 162.650 15.425 162.840 ;
        RECT 16.175 162.670 16.345 162.860 ;
        RECT 20.040 162.650 20.210 162.840 ;
        RECT 21.050 162.650 21.220 162.840 ;
        RECT 24.970 162.700 25.090 162.810 ;
        RECT 25.375 162.670 25.545 162.860 ;
        RECT 25.835 162.810 26.005 162.840 ;
        RECT 25.835 162.700 26.010 162.810 ;
        RECT 25.835 162.650 26.005 162.700 ;
        RECT 28.595 162.670 28.765 162.860 ;
        RECT 35.090 162.700 35.210 162.810 ;
        RECT 35.770 162.650 35.940 162.840 ;
        RECT 37.795 162.670 37.965 162.860 ;
        RECT 39.635 162.670 39.805 162.860 ;
        RECT 40.555 162.650 40.725 162.840 ;
        RECT 41.475 162.670 41.645 162.860 ;
        RECT 44.230 162.650 44.400 162.840 ;
        RECT 44.750 162.700 44.870 162.810 ;
        RECT 45.340 162.670 45.510 162.860 ;
        RECT 46.075 162.650 46.245 162.840 ;
        RECT 46.590 162.700 46.710 162.810 ;
        RECT 49.295 162.650 49.465 162.840 ;
        RECT 49.480 162.670 49.650 162.860 ;
        RECT 49.755 162.650 49.925 162.840 ;
        RECT 51.595 162.810 51.765 162.860 ;
        RECT 51.595 162.700 51.770 162.810 ;
        RECT 51.595 162.670 51.765 162.700 ;
        RECT 52.055 162.670 52.225 162.860 ;
        RECT 53.895 162.705 54.055 162.815 ;
        RECT 56.655 162.670 56.825 162.860 ;
        RECT 57.115 162.650 57.285 162.840 ;
        RECT 58.955 162.650 59.125 162.840 ;
        RECT 59.410 162.670 59.580 162.860 ;
        RECT 60.795 162.650 60.965 162.840 ;
        RECT 61.255 162.650 61.425 162.840 ;
        RECT 62.175 162.670 62.345 162.860 ;
        RECT 63.095 162.650 63.265 162.840 ;
        RECT 63.555 162.670 63.725 162.860 ;
        RECT 65.395 162.695 65.555 162.805 ;
        RECT 67.695 162.670 67.865 162.860 ;
        RECT 70.915 162.650 71.085 162.840 ;
        RECT 72.295 162.650 72.465 162.840 ;
        RECT 76.160 162.650 76.330 162.840 ;
        RECT 77.355 162.670 77.525 162.860 ;
        RECT 78.275 162.650 78.445 162.840 ;
        RECT 78.735 162.810 78.905 162.860 ;
        RECT 78.735 162.700 78.910 162.810 ;
        RECT 78.735 162.670 78.905 162.700 ;
        RECT 79.195 162.650 79.365 162.840 ;
        RECT 84.255 162.670 84.425 162.860 ;
        RECT 88.120 162.670 88.290 162.860 ;
        RECT 89.315 162.705 89.475 162.815 ;
        RECT 89.775 162.650 89.945 162.840 ;
        RECT 90.695 162.705 90.855 162.815 ;
        RECT 94.560 162.670 94.730 162.860 ;
        RECT 95.295 162.670 95.465 162.860 ;
        RECT 96.950 162.670 97.120 162.860 ;
        RECT 99.435 162.650 99.605 162.840 ;
        RECT 101.275 162.705 101.435 162.815 ;
        RECT 101.735 162.670 101.905 162.860 ;
        RECT 102.190 162.650 102.360 162.840 ;
        RECT 106.520 162.650 106.690 162.840 ;
        RECT 110.475 162.650 110.645 162.840 ;
        RECT 110.935 162.650 111.105 162.840 ;
        RECT 111.855 162.670 112.025 162.860 ;
        RECT 113.235 162.670 113.405 162.860 ;
        RECT 114.155 162.705 114.315 162.815 ;
        RECT 115.535 162.650 115.705 162.860 ;
        RECT 10.515 161.840 11.885 162.650 ;
        RECT 12.355 161.840 15.105 162.650 ;
        RECT 15.125 161.740 16.475 162.650 ;
        RECT 16.725 161.970 20.625 162.650 ;
        RECT 19.695 161.740 20.625 161.970 ;
        RECT 20.635 161.970 24.535 162.650 ;
        RECT 20.635 161.740 21.565 161.970 ;
        RECT 25.245 161.780 25.675 162.565 ;
        RECT 25.695 161.970 34.885 162.650 ;
        RECT 30.205 161.750 31.135 161.970 ;
        RECT 33.965 161.740 34.885 161.970 ;
        RECT 35.355 161.970 39.255 162.650 ;
        RECT 35.355 161.740 36.285 161.970 ;
        RECT 39.495 161.840 40.865 162.650 ;
        RECT 41.070 161.740 44.545 162.650 ;
        RECT 45.015 161.870 46.385 162.650 ;
        RECT 46.855 161.840 49.605 162.650 ;
        RECT 49.625 161.740 50.975 162.650 ;
        RECT 51.005 161.780 51.435 162.565 ;
        RECT 51.915 161.840 57.425 162.650 ;
        RECT 57.435 161.970 59.265 162.650 ;
        RECT 59.275 161.970 61.105 162.650 ;
        RECT 61.115 161.970 62.945 162.650 ;
        RECT 62.955 161.970 64.785 162.650 ;
        RECT 57.435 161.740 58.780 161.970 ;
        RECT 59.275 161.740 60.620 161.970 ;
        RECT 61.600 161.740 62.945 161.970 ;
        RECT 63.440 161.740 64.785 161.970 ;
        RECT 65.715 161.840 71.225 162.650 ;
        RECT 71.245 161.740 72.595 162.650 ;
        RECT 72.845 161.970 76.745 162.650 ;
        RECT 75.815 161.740 76.745 161.970 ;
        RECT 76.765 161.780 77.195 162.565 ;
        RECT 77.225 161.740 78.575 162.650 ;
        RECT 79.055 161.870 80.425 162.650 ;
        RECT 80.805 161.970 90.085 162.650 ;
        RECT 90.465 161.970 99.745 162.650 ;
        RECT 80.805 161.850 83.140 161.970 ;
        RECT 80.805 161.740 81.725 161.850 ;
        RECT 87.805 161.750 88.725 161.970 ;
        RECT 90.465 161.850 92.800 161.970 ;
        RECT 90.465 161.740 91.385 161.850 ;
        RECT 97.465 161.750 98.385 161.970 ;
        RECT 99.895 161.740 102.505 162.650 ;
        RECT 102.525 161.780 102.955 162.565 ;
        RECT 103.205 161.970 107.105 162.650 ;
        RECT 106.175 161.740 107.105 161.970 ;
        RECT 107.210 161.970 110.675 162.650 ;
        RECT 110.905 161.970 114.370 162.650 ;
        RECT 107.210 161.740 108.130 161.970 ;
        RECT 113.450 161.740 114.370 161.970 ;
        RECT 114.475 161.840 115.845 162.650 ;
      LAYER nwell ;
        RECT 10.320 158.620 116.040 161.450 ;
      LAYER pwell ;
        RECT 10.515 157.420 11.885 158.230 ;
        RECT 12.365 157.505 12.795 158.290 ;
        RECT 13.185 158.220 14.105 158.330 ;
        RECT 13.185 158.100 15.520 158.220 ;
        RECT 20.185 158.100 21.105 158.320 ;
        RECT 13.185 157.420 22.465 158.100 ;
        RECT 22.475 157.420 23.845 158.200 ;
        RECT 23.855 157.420 25.225 158.230 ;
        RECT 27.890 158.100 28.810 158.330 ;
        RECT 25.345 157.420 28.810 158.100 ;
        RECT 28.915 158.100 29.845 158.330 ;
        RECT 28.915 157.420 32.815 158.100 ;
        RECT 33.055 157.420 34.425 158.230 ;
        RECT 34.435 157.420 37.910 158.330 ;
        RECT 38.125 157.505 38.555 158.290 ;
        RECT 38.575 157.420 39.945 158.230 ;
        RECT 40.150 157.420 43.625 158.330 ;
        RECT 43.635 157.420 47.110 158.330 ;
        RECT 47.685 158.220 48.605 158.330 ;
        RECT 47.685 158.100 50.020 158.220 ;
        RECT 54.685 158.100 55.605 158.320 ;
        RECT 47.685 157.420 56.965 158.100 ;
        RECT 57.115 157.420 59.725 158.330 ;
        RECT 60.195 157.420 62.025 158.230 ;
        RECT 62.035 158.100 63.380 158.330 ;
        RECT 62.035 157.420 63.865 158.100 ;
        RECT 63.885 157.505 64.315 158.290 ;
        RECT 64.795 157.420 67.545 158.230 ;
        RECT 67.555 157.420 71.030 158.330 ;
        RECT 71.695 157.420 73.525 158.230 ;
        RECT 73.905 158.220 74.825 158.330 ;
        RECT 73.905 158.100 76.240 158.220 ;
        RECT 80.905 158.100 81.825 158.320 ;
        RECT 73.905 157.420 83.185 158.100 ;
        RECT 84.125 157.420 85.475 158.330 ;
        RECT 86.150 157.420 89.625 158.330 ;
        RECT 89.645 157.505 90.075 158.290 ;
        RECT 90.095 157.420 91.465 158.200 ;
        RECT 92.490 158.100 93.410 158.330 ;
        RECT 92.490 157.420 95.955 158.100 ;
        RECT 96.075 157.420 97.445 158.200 ;
        RECT 97.650 157.420 101.125 158.330 ;
        RECT 101.595 157.420 103.425 158.230 ;
        RECT 106.635 158.100 107.565 158.330 ;
        RECT 103.665 157.420 107.565 158.100 ;
        RECT 108.035 157.420 109.865 158.230 ;
        RECT 109.875 157.420 111.245 158.200 ;
        RECT 111.715 157.420 114.465 158.230 ;
        RECT 114.475 157.420 115.845 158.230 ;
        RECT 10.655 157.210 10.825 157.420 ;
        RECT 12.090 157.260 12.210 157.370 ;
        RECT 14.795 157.210 14.965 157.400 ;
        RECT 15.255 157.210 15.425 157.400 ;
        RECT 20.040 157.210 20.210 157.400 ;
        RECT 21.235 157.255 21.395 157.365 ;
        RECT 22.155 157.230 22.325 157.420 ;
        RECT 23.535 157.230 23.705 157.420 ;
        RECT 24.915 157.210 25.085 157.420 ;
        RECT 25.375 157.230 25.545 157.420 ;
        RECT 25.835 157.210 26.005 157.400 ;
        RECT 29.330 157.230 29.500 157.420 ;
        RECT 29.520 157.210 29.690 157.400 ;
        RECT 33.250 157.260 33.370 157.370 ;
        RECT 34.115 157.230 34.285 157.420 ;
        RECT 34.580 157.230 34.750 157.420 ;
        RECT 36.870 157.210 37.040 157.400 ;
        RECT 39.635 157.230 39.805 157.420 ;
        RECT 40.550 157.210 40.720 157.400 ;
        RECT 41.070 157.260 41.190 157.370 ;
        RECT 43.310 157.230 43.480 157.420 ;
        RECT 43.780 157.400 43.950 157.420 ;
        RECT 43.775 157.230 43.950 157.400 ;
        RECT 43.775 157.210 43.945 157.230 ;
        RECT 49.295 157.210 49.465 157.400 ;
        RECT 49.755 157.210 49.925 157.400 ;
        RECT 56.655 157.230 56.825 157.420 ;
        RECT 59.410 157.230 59.580 157.420 ;
        RECT 59.930 157.260 60.050 157.370 ;
        RECT 60.795 157.210 60.965 157.400 ;
        RECT 61.715 157.230 61.885 157.420 ;
        RECT 62.635 157.210 62.805 157.400 ;
        RECT 63.095 157.210 63.265 157.400 ;
        RECT 63.555 157.230 63.725 157.420 ;
        RECT 64.530 157.260 64.650 157.370 ;
        RECT 67.235 157.230 67.405 157.420 ;
        RECT 67.700 157.230 67.870 157.420 ;
        RECT 68.150 157.210 68.320 157.400 ;
        RECT 68.620 157.210 68.790 157.400 ;
        RECT 71.430 157.260 71.550 157.370 ;
        RECT 72.755 157.255 72.915 157.365 ;
        RECT 73.215 157.230 73.385 157.420 ;
        RECT 76.435 157.210 76.605 157.400 ;
        RECT 77.815 157.255 77.975 157.365 ;
        RECT 81.495 157.210 81.665 157.400 ;
        RECT 82.875 157.230 83.045 157.420 ;
        RECT 83.795 157.265 83.955 157.375 ;
        RECT 85.175 157.230 85.345 157.420 ;
        RECT 85.690 157.260 85.810 157.370 ;
        RECT 87.015 157.210 87.185 157.400 ;
        RECT 87.480 157.210 87.650 157.400 ;
        RECT 89.310 157.230 89.480 157.420 ;
        RECT 91.155 157.230 91.325 157.420 ;
        RECT 92.075 157.265 92.235 157.375 ;
        RECT 93.455 157.210 93.625 157.400 ;
        RECT 93.920 157.210 94.090 157.400 ;
        RECT 95.755 157.230 95.925 157.420 ;
        RECT 96.215 157.230 96.385 157.420 ;
        RECT 98.515 157.210 98.685 157.400 ;
        RECT 98.980 157.210 99.150 157.400 ;
        RECT 100.810 157.230 100.980 157.420 ;
        RECT 101.330 157.260 101.450 157.370 ;
        RECT 103.115 157.230 103.285 157.420 ;
        RECT 104.495 157.210 104.665 157.400 ;
        RECT 104.955 157.210 105.125 157.400 ;
        RECT 106.980 157.230 107.150 157.420 ;
        RECT 107.770 157.260 107.890 157.370 ;
        RECT 108.640 157.210 108.810 157.400 ;
        RECT 109.555 157.230 109.725 157.420 ;
        RECT 110.015 157.230 110.185 157.420 ;
        RECT 111.450 157.260 111.570 157.370 ;
        RECT 114.155 157.210 114.325 157.420 ;
        RECT 115.535 157.210 115.705 157.420 ;
        RECT 10.515 156.400 11.885 157.210 ;
        RECT 12.355 156.400 15.105 157.210 ;
        RECT 15.125 156.300 16.475 157.210 ;
        RECT 16.725 156.530 20.625 157.210 ;
        RECT 19.695 156.300 20.625 156.530 ;
        RECT 21.650 156.530 25.115 157.210 ;
        RECT 21.650 156.300 22.570 156.530 ;
        RECT 25.245 156.340 25.675 157.125 ;
        RECT 25.805 156.530 29.270 157.210 ;
        RECT 28.350 156.300 29.270 156.530 ;
        RECT 29.375 156.300 32.850 157.210 ;
        RECT 33.710 156.300 37.185 157.210 ;
        RECT 37.390 156.300 40.865 157.210 ;
        RECT 41.335 156.400 44.085 157.210 ;
        RECT 44.095 156.400 49.605 157.210 ;
        RECT 49.615 156.430 50.985 157.210 ;
        RECT 51.005 156.340 51.435 157.125 ;
        RECT 51.825 156.530 61.105 157.210 ;
        RECT 61.115 156.530 62.945 157.210 ;
        RECT 62.955 156.530 64.785 157.210 ;
        RECT 51.825 156.410 54.160 156.530 ;
        RECT 51.825 156.300 52.745 156.410 ;
        RECT 58.825 156.310 59.745 156.530 ;
        RECT 61.115 156.300 62.460 156.530 ;
        RECT 63.440 156.300 64.785 156.530 ;
        RECT 64.990 156.300 68.465 157.210 ;
        RECT 68.475 156.300 71.950 157.210 ;
        RECT 73.075 156.400 76.745 157.210 ;
        RECT 76.765 156.340 77.195 157.125 ;
        RECT 78.135 156.400 81.805 157.210 ;
        RECT 81.815 156.400 87.325 157.210 ;
        RECT 87.335 156.300 90.810 157.210 ;
        RECT 91.015 156.400 93.765 157.210 ;
        RECT 93.775 156.300 97.250 157.210 ;
        RECT 97.455 156.400 98.825 157.210 ;
        RECT 98.835 156.300 102.310 157.210 ;
        RECT 102.525 156.340 102.955 157.125 ;
        RECT 102.975 156.400 104.805 157.210 ;
        RECT 104.925 156.530 108.390 157.210 ;
        RECT 107.470 156.300 108.390 156.530 ;
        RECT 108.495 156.300 111.105 157.210 ;
        RECT 111.715 156.400 114.465 157.210 ;
        RECT 114.475 156.400 115.845 157.210 ;
      LAYER nwell ;
        RECT 10.320 153.180 116.040 156.010 ;
      LAYER pwell ;
        RECT 10.515 151.980 11.885 152.790 ;
        RECT 12.365 152.065 12.795 152.850 ;
        RECT 13.185 152.780 14.105 152.890 ;
        RECT 13.185 152.660 15.520 152.780 ;
        RECT 20.185 152.660 21.105 152.880 ;
        RECT 13.185 151.980 22.465 152.660 ;
        RECT 22.475 151.980 23.845 152.760 ;
        RECT 24.315 151.980 27.985 152.790 ;
        RECT 27.995 152.660 28.925 152.890 ;
        RECT 27.995 151.980 31.895 152.660 ;
        RECT 32.595 151.980 38.105 152.790 ;
        RECT 38.125 152.065 38.555 152.850 ;
        RECT 39.495 151.980 43.165 152.790 ;
        RECT 43.175 151.980 48.685 152.790 ;
        RECT 48.695 152.660 49.625 152.890 ;
        RECT 52.835 152.660 53.765 152.890 ;
        RECT 48.695 151.980 52.595 152.660 ;
        RECT 52.835 151.980 56.735 152.660 ;
        RECT 57.895 151.980 59.265 152.760 ;
        RECT 59.275 152.660 60.620 152.890 ;
        RECT 61.115 152.660 62.460 152.890 ;
        RECT 59.275 151.980 61.105 152.660 ;
        RECT 61.115 151.980 62.945 152.660 ;
        RECT 63.885 152.065 64.315 152.850 ;
        RECT 64.335 152.660 65.680 152.890 ;
        RECT 64.335 151.980 66.165 152.660 ;
        RECT 66.175 151.980 68.895 152.890 ;
        RECT 68.935 151.980 72.410 152.890 ;
        RECT 73.075 151.980 75.825 152.790 ;
        RECT 75.835 151.980 81.345 152.790 ;
        RECT 81.365 151.980 82.715 152.890 ;
        RECT 82.735 151.980 84.105 152.760 ;
        RECT 84.575 151.980 88.245 152.790 ;
        RECT 88.265 151.980 89.615 152.890 ;
        RECT 89.645 152.065 90.075 152.850 ;
        RECT 90.095 151.980 95.605 152.790 ;
        RECT 95.615 151.980 99.090 152.890 ;
        RECT 102.410 152.660 103.330 152.890 ;
        RECT 106.635 152.660 107.565 152.890 ;
        RECT 99.865 151.980 103.330 152.660 ;
        RECT 103.665 151.980 107.565 152.660 ;
        RECT 107.575 151.980 109.405 152.790 ;
        RECT 109.415 151.980 110.785 152.760 ;
        RECT 110.795 151.980 114.465 152.790 ;
        RECT 114.475 151.980 115.845 152.790 ;
        RECT 10.655 151.770 10.825 151.980 ;
        RECT 12.090 151.820 12.210 151.930 ;
        RECT 12.955 151.770 13.125 151.960 ;
        RECT 16.635 151.770 16.805 151.960 ;
        RECT 20.500 151.770 20.670 151.960 ;
        RECT 22.155 151.790 22.325 151.980 ;
        RECT 23.535 151.770 23.705 151.980 ;
        RECT 23.995 151.930 24.165 151.960 ;
        RECT 23.995 151.820 24.170 151.930 ;
        RECT 23.995 151.770 24.165 151.820 ;
        RECT 27.675 151.790 27.845 151.980 ;
        RECT 28.410 151.790 28.580 151.980 ;
        RECT 32.330 151.820 32.450 151.930 ;
        RECT 35.035 151.770 35.205 151.960 ;
        RECT 35.500 151.770 35.670 151.960 ;
        RECT 37.795 151.790 37.965 151.980 ;
        RECT 39.175 151.825 39.335 151.935 ;
        RECT 40.095 151.770 40.265 151.960 ;
        RECT 10.515 150.960 11.885 151.770 ;
        RECT 11.895 150.960 13.265 151.770 ;
        RECT 13.275 150.960 16.945 151.770 ;
        RECT 17.185 151.090 21.085 151.770 ;
        RECT 20.155 150.860 21.085 151.090 ;
        RECT 21.095 150.960 23.845 151.770 ;
        RECT 23.865 150.860 25.215 151.770 ;
        RECT 25.245 150.900 25.675 151.685 ;
        RECT 26.065 151.090 35.345 151.770 ;
        RECT 26.065 150.970 28.400 151.090 ;
        RECT 26.065 150.860 26.985 150.970 ;
        RECT 33.065 150.870 33.985 151.090 ;
        RECT 35.355 150.860 38.830 151.770 ;
        RECT 39.035 150.960 40.405 151.770 ;
        RECT 40.560 151.740 40.730 151.960 ;
        RECT 42.855 151.790 43.025 151.980 ;
        RECT 42.220 151.740 43.165 151.770 ;
        RECT 40.415 151.060 43.165 151.740 ;
        RECT 42.220 150.860 43.165 151.060 ;
        RECT 43.175 151.740 44.120 151.770 ;
        RECT 45.610 151.740 45.780 151.960 ;
        RECT 46.130 151.820 46.250 151.930 ;
        RECT 46.540 151.770 46.710 151.960 ;
        RECT 48.375 151.790 48.545 151.980 ;
        RECT 49.110 151.790 49.280 151.980 ;
        RECT 50.675 151.815 50.835 151.925 ;
        RECT 51.650 151.820 51.770 151.930 ;
        RECT 52.055 151.770 52.225 151.960 ;
        RECT 53.250 151.790 53.420 151.980 ;
        RECT 53.435 151.770 53.605 151.960 ;
        RECT 57.575 151.825 57.735 151.935 ;
        RECT 58.035 151.790 58.205 151.980 ;
        RECT 60.795 151.790 60.965 151.980 ;
        RECT 62.635 151.790 62.805 151.980 ;
        RECT 63.555 151.770 63.725 151.960 ;
        RECT 65.855 151.790 66.025 151.980 ;
        RECT 66.315 151.770 66.485 151.980 ;
        RECT 67.695 151.770 67.865 151.960 ;
        RECT 69.080 151.790 69.250 151.980 ;
        RECT 43.175 151.060 45.925 151.740 ;
        RECT 43.175 150.860 44.120 151.060 ;
        RECT 46.395 150.860 49.870 151.770 ;
        RECT 51.005 150.900 51.435 151.685 ;
        RECT 51.925 150.860 53.275 151.770 ;
        RECT 53.295 150.990 54.665 151.770 ;
        RECT 54.760 151.090 63.865 151.770 ;
        RECT 63.885 151.090 66.625 151.770 ;
        RECT 66.635 150.960 68.005 151.770 ;
        RECT 68.015 151.740 68.960 151.770 ;
        RECT 70.450 151.740 70.620 151.960 ;
        RECT 70.915 151.770 71.085 151.960 ;
        RECT 72.810 151.820 72.930 151.930 ;
        RECT 73.730 151.820 73.850 151.930 ;
        RECT 75.515 151.790 75.685 151.980 ;
        RECT 76.435 151.770 76.605 151.960 ;
        RECT 81.035 151.790 81.205 151.980 ;
        RECT 82.415 151.790 82.585 151.980 ;
        RECT 82.875 151.790 83.045 151.980 ;
        RECT 84.310 151.820 84.430 151.930 ;
        RECT 86.555 151.770 86.725 151.960 ;
        RECT 87.935 151.790 88.105 151.980 ;
        RECT 88.395 151.790 88.565 151.980 ;
        RECT 95.295 151.790 95.465 151.980 ;
        RECT 95.760 151.960 95.930 151.980 ;
        RECT 95.755 151.790 95.930 151.960 ;
        RECT 95.755 151.770 95.925 151.790 ;
        RECT 68.015 151.060 70.765 151.740 ;
        RECT 70.775 151.090 73.515 151.770 ;
        RECT 68.015 150.860 68.960 151.060 ;
        RECT 73.995 150.960 76.745 151.770 ;
        RECT 76.765 150.900 77.195 151.685 ;
        RECT 77.585 151.090 86.865 151.770 ;
        RECT 86.875 151.090 96.065 151.770 ;
        RECT 96.075 151.740 97.020 151.770 ;
        RECT 98.510 151.740 98.680 151.960 ;
        RECT 98.980 151.770 99.150 151.960 ;
        RECT 99.490 151.820 99.610 151.930 ;
        RECT 99.895 151.790 100.065 151.980 ;
        RECT 103.170 151.820 103.290 151.930 ;
        RECT 103.575 151.770 103.745 151.960 ;
        RECT 106.980 151.790 107.150 151.980 ;
        RECT 109.095 151.790 109.265 151.980 ;
        RECT 109.555 151.790 109.725 151.980 ;
        RECT 113.695 151.770 113.865 151.960 ;
        RECT 114.155 151.930 114.325 151.980 ;
        RECT 114.155 151.820 114.330 151.930 ;
        RECT 114.155 151.790 114.325 151.820 ;
        RECT 115.535 151.770 115.705 151.980 ;
        RECT 77.585 150.970 79.920 151.090 ;
        RECT 77.585 150.860 78.505 150.970 ;
        RECT 84.585 150.870 85.505 151.090 ;
        RECT 86.875 150.860 87.795 151.090 ;
        RECT 90.625 150.870 91.555 151.090 ;
        RECT 96.075 151.060 98.825 151.740 ;
        RECT 96.075 150.860 97.020 151.060 ;
        RECT 98.835 150.860 102.310 151.770 ;
        RECT 102.525 150.900 102.955 151.685 ;
        RECT 103.445 150.860 104.795 151.770 ;
        RECT 104.815 151.090 114.005 151.770 ;
        RECT 104.815 150.860 105.735 151.090 ;
        RECT 108.565 150.870 109.495 151.090 ;
        RECT 114.475 150.960 115.845 151.770 ;
      LAYER nwell ;
        RECT 10.320 147.740 116.040 150.570 ;
      LAYER pwell ;
        RECT 10.515 146.540 11.885 147.350 ;
        RECT 12.365 146.625 12.795 147.410 ;
        RECT 13.185 147.340 14.105 147.450 ;
        RECT 13.185 147.220 15.520 147.340 ;
        RECT 20.185 147.220 21.105 147.440 ;
        RECT 13.185 146.540 22.465 147.220 ;
        RECT 22.475 146.540 23.845 147.350 ;
        RECT 23.855 147.220 24.785 147.450 ;
        RECT 23.855 146.540 27.755 147.220 ;
        RECT 28.915 146.540 30.285 147.320 ;
        RECT 30.490 146.540 33.965 147.450 ;
        RECT 33.975 146.540 36.725 147.350 ;
        RECT 36.745 146.540 38.095 147.450 ;
        RECT 38.125 146.625 38.555 147.410 ;
        RECT 38.575 146.540 41.325 147.350 ;
        RECT 43.140 147.250 44.085 147.450 ;
        RECT 41.335 146.570 44.085 147.250 ;
        RECT 10.655 146.330 10.825 146.540 ;
        RECT 12.090 146.380 12.210 146.490 ;
        RECT 13.875 146.330 14.045 146.520 ;
        RECT 15.255 146.330 15.425 146.520 ;
        RECT 22.155 146.350 22.325 146.540 ;
        RECT 23.535 146.350 23.705 146.540 ;
        RECT 24.270 146.350 24.440 146.540 ;
        RECT 24.915 146.330 25.085 146.520 ;
        RECT 26.755 146.330 26.925 146.520 ;
        RECT 28.595 146.385 28.755 146.495 ;
        RECT 29.055 146.350 29.225 146.540 ;
        RECT 29.515 146.330 29.685 146.520 ;
        RECT 29.980 146.330 30.150 146.520 ;
        RECT 33.650 146.490 33.820 146.540 ;
        RECT 33.650 146.380 33.830 146.490 ;
        RECT 33.650 146.350 33.820 146.380 ;
        RECT 34.115 146.330 34.285 146.520 ;
        RECT 36.415 146.350 36.585 146.540 ;
        RECT 36.875 146.350 37.045 146.540 ;
        RECT 41.015 146.350 41.185 146.540 ;
        RECT 41.480 146.350 41.650 146.570 ;
        RECT 43.140 146.540 44.085 146.570 ;
        RECT 44.095 146.540 47.570 147.450 ;
        RECT 48.695 146.540 52.170 147.450 ;
        RECT 53.665 147.340 54.585 147.450 ;
        RECT 53.665 147.220 56.000 147.340 ;
        RECT 60.665 147.220 61.585 147.440 ;
        RECT 53.665 146.540 62.945 147.220 ;
        RECT 63.885 146.625 64.315 147.410 ;
        RECT 64.335 147.250 65.280 147.450 ;
        RECT 64.335 146.570 67.085 147.250 ;
        RECT 64.335 146.540 65.280 146.570 ;
        RECT 43.830 146.380 43.950 146.490 ;
        RECT 44.240 146.350 44.410 146.540 ;
        RECT 44.510 146.330 44.680 146.520 ;
        RECT 48.375 146.385 48.535 146.495 ;
        RECT 48.840 146.350 49.010 146.540 ;
        RECT 50.675 146.330 50.845 146.520 ;
        RECT 52.975 146.330 53.145 146.520 ;
        RECT 53.435 146.330 53.605 146.520 ;
        RECT 58.220 146.330 58.390 146.520 ;
        RECT 59.875 146.330 60.045 146.520 ;
        RECT 62.635 146.350 62.805 146.540 ;
        RECT 63.555 146.385 63.715 146.495 ;
        RECT 65.395 146.330 65.565 146.520 ;
        RECT 65.855 146.330 66.025 146.520 ;
        RECT 66.770 146.350 66.940 146.570 ;
        RECT 67.290 146.540 70.765 147.450 ;
        RECT 70.775 146.540 74.250 147.450 ;
        RECT 74.455 146.540 75.825 147.320 ;
        RECT 77.195 147.220 78.115 147.440 ;
        RECT 84.195 147.340 85.115 147.450 ;
        RECT 82.780 147.220 85.115 147.340 ;
        RECT 88.695 147.220 89.625 147.450 ;
        RECT 75.835 146.540 85.115 147.220 ;
        RECT 85.725 146.540 89.625 147.220 ;
        RECT 89.645 146.625 90.075 147.410 ;
        RECT 90.095 146.540 91.925 147.350 ;
        RECT 91.935 146.540 93.305 147.320 ;
        RECT 94.235 147.250 95.180 147.450 ;
        RECT 94.235 146.570 96.985 147.250 ;
        RECT 94.235 146.540 95.180 146.570 ;
        RECT 68.615 146.330 68.785 146.520 ;
        RECT 70.450 146.350 70.620 146.540 ;
        RECT 70.920 146.350 71.090 146.540 ;
        RECT 72.295 146.330 72.465 146.520 ;
        RECT 74.595 146.350 74.765 146.540 ;
        RECT 75.975 146.350 76.145 146.540 ;
        RECT 76.160 146.330 76.330 146.520 ;
        RECT 77.410 146.380 77.530 146.490 ;
        RECT 81.220 146.330 81.390 146.520 ;
        RECT 82.875 146.330 83.045 146.520 ;
        RECT 83.390 146.380 83.510 146.490 ;
        RECT 83.795 146.330 83.965 146.520 ;
        RECT 87.530 146.380 87.650 146.490 ;
        RECT 89.040 146.350 89.210 146.540 ;
        RECT 90.235 146.330 90.405 146.520 ;
        RECT 91.615 146.350 91.785 146.540 ;
        RECT 92.075 146.350 92.245 146.540 ;
        RECT 93.915 146.385 94.075 146.495 ;
        RECT 95.755 146.330 95.925 146.520 ;
        RECT 96.670 146.350 96.840 146.570 ;
        RECT 96.995 146.540 100.470 147.450 ;
        RECT 103.875 147.220 104.805 147.450 ;
        RECT 100.905 146.540 104.805 147.220 ;
        RECT 105.185 147.340 106.105 147.450 ;
        RECT 105.185 147.220 107.520 147.340 ;
        RECT 112.185 147.220 113.105 147.440 ;
        RECT 105.185 146.540 114.465 147.220 ;
        RECT 114.475 146.540 115.845 147.350 ;
        RECT 97.140 146.350 97.310 146.540 ;
        RECT 10.515 145.520 11.885 146.330 ;
        RECT 12.355 145.520 14.185 146.330 ;
        RECT 14.205 145.420 15.555 146.330 ;
        RECT 15.945 145.650 25.225 146.330 ;
        RECT 15.945 145.530 18.280 145.650 ;
        RECT 15.945 145.420 16.865 145.530 ;
        RECT 22.945 145.430 23.865 145.650 ;
        RECT 25.245 145.460 25.675 146.245 ;
        RECT 25.695 145.550 27.065 146.330 ;
        RECT 27.075 145.520 29.825 146.330 ;
        RECT 29.835 145.420 33.310 146.330 ;
        RECT 33.975 145.650 43.255 146.330 ;
        RECT 35.335 145.430 36.255 145.650 ;
        RECT 40.920 145.530 43.255 145.650 ;
        RECT 42.335 145.420 43.255 145.530 ;
        RECT 44.095 145.650 47.995 146.330 ;
        RECT 44.095 145.420 45.025 145.650 ;
        RECT 48.235 145.520 50.985 146.330 ;
        RECT 51.005 145.460 51.435 146.245 ;
        RECT 51.455 145.520 53.285 146.330 ;
        RECT 53.305 145.420 54.655 146.330 ;
        RECT 54.905 145.650 58.805 146.330 ;
        RECT 57.875 145.420 58.805 145.650 ;
        RECT 58.815 145.520 60.185 146.330 ;
        RECT 60.195 145.520 65.705 146.330 ;
        RECT 65.715 145.650 67.545 146.330 ;
        RECT 66.200 145.420 67.545 145.650 ;
        RECT 67.555 145.520 68.925 146.330 ;
        RECT 68.935 145.520 72.605 146.330 ;
        RECT 72.845 145.650 76.745 146.330 ;
        RECT 75.815 145.420 76.745 145.650 ;
        RECT 76.765 145.460 77.195 146.245 ;
        RECT 77.905 145.650 81.805 146.330 ;
        RECT 80.875 145.420 81.805 145.650 ;
        RECT 81.825 145.420 83.175 146.330 ;
        RECT 83.765 145.650 87.230 146.330 ;
        RECT 86.310 145.420 87.230 145.650 ;
        RECT 87.795 145.520 90.545 146.330 ;
        RECT 90.555 145.520 96.065 146.330 ;
        RECT 96.075 146.300 97.020 146.330 ;
        RECT 98.510 146.300 98.680 146.520 ;
        RECT 98.980 146.330 99.150 146.520 ;
        RECT 104.035 146.330 104.205 146.520 ;
        RECT 104.220 146.350 104.390 146.540 ;
        RECT 107.715 146.330 107.885 146.520 ;
        RECT 108.175 146.330 108.345 146.520 ;
        RECT 109.610 146.380 109.730 146.490 ;
        RECT 110.015 146.330 110.185 146.520 ;
        RECT 111.450 146.380 111.570 146.490 ;
        RECT 114.155 146.330 114.325 146.540 ;
        RECT 115.535 146.330 115.705 146.540 ;
        RECT 96.075 145.620 98.825 146.300 ;
        RECT 96.075 145.420 97.020 145.620 ;
        RECT 98.835 145.420 102.310 146.330 ;
        RECT 102.525 145.460 102.955 146.245 ;
        RECT 102.975 145.520 104.345 146.330 ;
        RECT 104.355 145.520 108.025 146.330 ;
        RECT 108.045 145.420 109.395 146.330 ;
        RECT 109.875 145.550 111.245 146.330 ;
        RECT 111.715 145.520 114.465 146.330 ;
        RECT 114.475 145.520 115.845 146.330 ;
      LAYER nwell ;
        RECT 10.320 142.300 116.040 145.130 ;
      LAYER pwell ;
        RECT 10.515 141.100 11.885 141.910 ;
        RECT 12.365 141.185 12.795 141.970 ;
        RECT 13.735 141.100 19.245 141.910 ;
        RECT 19.255 141.100 20.625 141.880 ;
        RECT 20.645 141.100 21.995 142.010 ;
        RECT 22.015 141.100 23.385 141.910 ;
        RECT 23.395 141.100 27.065 141.910 ;
        RECT 27.075 141.100 32.585 141.910 ;
        RECT 32.595 141.100 38.105 141.910 ;
        RECT 38.125 141.185 38.555 141.970 ;
        RECT 39.035 141.100 41.785 141.910 ;
        RECT 41.795 141.100 43.165 141.880 ;
        RECT 43.175 141.100 46.650 142.010 ;
        RECT 46.855 141.100 48.225 141.910 ;
        RECT 48.235 141.100 51.710 142.010 ;
        RECT 51.915 141.100 53.285 141.910 ;
        RECT 53.305 141.100 54.655 142.010 ;
        RECT 54.675 141.780 55.595 142.010 ;
        RECT 58.425 141.780 59.355 142.000 ;
        RECT 54.675 141.100 63.865 141.780 ;
        RECT 63.885 141.185 64.315 141.970 ;
        RECT 64.335 141.100 67.085 141.910 ;
        RECT 67.095 141.810 68.040 142.010 ;
        RECT 67.095 141.130 69.845 141.810 ;
        RECT 67.095 141.100 68.040 141.130 ;
        RECT 10.655 140.890 10.825 141.100 ;
        RECT 12.090 140.940 12.210 141.050 ;
        RECT 13.415 140.945 13.575 141.055 ;
        RECT 15.715 140.890 15.885 141.080 ;
        RECT 16.175 140.890 16.345 141.080 ;
        RECT 17.610 140.940 17.730 141.050 ;
        RECT 18.935 140.910 19.105 141.100 ;
        RECT 19.395 140.890 19.565 141.100 ;
        RECT 21.695 140.910 21.865 141.100 ;
        RECT 23.075 140.910 23.245 141.100 ;
        RECT 24.915 140.890 25.085 141.080 ;
        RECT 25.890 140.940 26.010 141.050 ;
        RECT 26.755 140.910 26.925 141.100 ;
        RECT 28.595 140.890 28.765 141.080 ;
        RECT 10.515 140.080 11.885 140.890 ;
        RECT 12.355 140.080 16.025 140.890 ;
        RECT 16.045 139.980 17.395 140.890 ;
        RECT 17.875 140.080 19.705 140.890 ;
        RECT 19.715 140.080 25.225 140.890 ;
        RECT 25.245 140.020 25.675 140.805 ;
        RECT 26.155 140.080 28.905 140.890 ;
        RECT 28.915 140.860 29.860 140.890 ;
        RECT 31.350 140.860 31.520 141.080 ;
        RECT 31.870 140.940 31.990 141.050 ;
        RECT 32.275 140.910 32.445 141.100 ;
        RECT 37.795 141.080 37.965 141.100 ;
        RECT 34.575 140.890 34.745 141.080 ;
        RECT 28.915 140.180 31.665 140.860 ;
        RECT 28.915 139.980 29.860 140.180 ;
        RECT 32.135 140.080 34.885 140.890 ;
        RECT 34.895 140.860 35.840 140.890 ;
        RECT 37.330 140.860 37.500 141.080 ;
        RECT 37.795 140.910 37.970 141.080 ;
        RECT 38.770 140.940 38.890 141.050 ;
        RECT 37.800 140.860 37.970 140.910 ;
        RECT 39.460 140.860 40.405 140.890 ;
        RECT 40.560 140.860 40.730 141.080 ;
        RECT 41.475 140.910 41.645 141.100 ;
        RECT 42.855 140.910 43.025 141.100 ;
        RECT 43.320 140.890 43.490 141.100 ;
        RECT 47.050 140.940 47.170 141.050 ;
        RECT 47.915 140.910 48.085 141.100 ;
        RECT 48.380 140.910 48.550 141.100 ;
        RECT 50.675 140.890 50.845 141.080 ;
        RECT 52.975 140.890 53.145 141.100 ;
        RECT 53.435 140.890 53.605 141.100 ;
        RECT 57.170 140.940 57.290 141.050 ;
        RECT 60.980 140.890 61.150 141.080 ;
        RECT 61.715 140.890 61.885 141.080 ;
        RECT 63.150 140.940 63.270 141.050 ;
        RECT 63.555 140.910 63.725 141.100 ;
        RECT 65.855 140.890 66.025 141.080 ;
        RECT 66.775 140.910 66.945 141.100 ;
        RECT 42.220 140.860 43.165 140.890 ;
        RECT 34.895 140.180 37.645 140.860 ;
        RECT 37.655 140.180 40.405 140.860 ;
        RECT 40.415 140.180 43.165 140.860 ;
        RECT 34.895 139.980 35.840 140.180 ;
        RECT 39.460 139.980 40.405 140.180 ;
        RECT 42.220 139.980 43.165 140.180 ;
        RECT 43.175 139.980 46.650 140.890 ;
        RECT 47.315 140.080 50.985 140.890 ;
        RECT 51.005 140.020 51.435 140.805 ;
        RECT 51.455 140.080 53.285 140.890 ;
        RECT 53.405 140.210 56.870 140.890 ;
        RECT 57.665 140.210 61.565 140.890 ;
        RECT 55.950 139.980 56.870 140.210 ;
        RECT 60.635 139.980 61.565 140.210 ;
        RECT 61.575 140.110 62.945 140.890 ;
        RECT 63.415 140.080 66.165 140.890 ;
        RECT 66.175 140.860 67.120 140.890 ;
        RECT 68.610 140.860 68.780 141.080 ;
        RECT 69.080 140.890 69.250 141.080 ;
        RECT 69.530 140.910 69.700 141.130 ;
        RECT 69.855 141.100 73.330 142.010 ;
        RECT 73.905 141.900 74.825 142.010 ;
        RECT 73.905 141.780 76.240 141.900 ;
        RECT 80.905 141.780 81.825 142.000 ;
        RECT 73.905 141.100 83.185 141.780 ;
        RECT 84.115 141.100 89.625 141.910 ;
        RECT 89.645 141.185 90.075 141.970 ;
        RECT 90.095 141.100 93.765 141.910 ;
        RECT 93.775 141.100 99.285 141.910 ;
        RECT 99.295 141.100 104.805 141.910 ;
        RECT 108.015 141.780 108.945 142.010 ;
        RECT 105.045 141.100 108.945 141.780 ;
        RECT 108.965 141.100 110.315 142.010 ;
        RECT 110.795 141.100 114.465 141.910 ;
        RECT 114.475 141.100 115.845 141.910 ;
        RECT 70.000 140.910 70.170 141.100 ;
        RECT 76.160 140.890 76.330 141.080 ;
        RECT 77.410 140.940 77.530 141.050 ;
        RECT 77.815 140.890 77.985 141.080 ;
        RECT 80.115 140.890 80.285 141.080 ;
        RECT 82.875 140.890 83.045 141.100 ;
        RECT 89.315 141.080 89.485 141.100 ;
        RECT 83.795 140.945 83.955 141.055 ;
        RECT 86.740 140.890 86.910 141.080 ;
        RECT 88.855 140.890 89.025 141.080 ;
        RECT 89.315 140.910 89.490 141.080 ;
        RECT 93.455 140.910 93.625 141.100 ;
        RECT 89.320 140.890 89.490 140.910 ;
        RECT 96.400 140.890 96.570 141.080 ;
        RECT 98.515 140.890 98.685 141.080 ;
        RECT 98.975 140.910 99.145 141.100 ;
        RECT 102.190 140.890 102.360 141.080 ;
        RECT 103.170 140.940 103.290 141.050 ;
        RECT 103.575 140.890 103.745 141.080 ;
        RECT 104.495 140.910 104.665 141.100 ;
        RECT 108.360 140.910 108.530 141.100 ;
        RECT 109.095 140.910 109.265 141.100 ;
        RECT 110.530 140.940 110.650 141.050 ;
        RECT 114.155 140.890 114.325 141.100 ;
        RECT 115.535 140.890 115.705 141.100 ;
        RECT 66.175 140.180 68.925 140.860 ;
        RECT 66.175 139.980 67.120 140.180 ;
        RECT 68.935 139.980 72.410 140.890 ;
        RECT 72.845 140.210 76.745 140.890 ;
        RECT 75.815 139.980 76.745 140.210 ;
        RECT 76.765 140.020 77.195 140.805 ;
        RECT 77.675 140.110 79.045 140.890 ;
        RECT 79.065 139.980 80.415 140.890 ;
        RECT 80.435 140.080 83.185 140.890 ;
        RECT 83.425 140.210 87.325 140.890 ;
        RECT 86.395 139.980 87.325 140.210 ;
        RECT 87.335 140.080 89.165 140.890 ;
        RECT 89.175 139.980 92.650 140.890 ;
        RECT 93.085 140.210 96.985 140.890 ;
        RECT 96.055 139.980 96.985 140.210 ;
        RECT 96.995 140.080 98.825 140.890 ;
        RECT 99.030 139.980 102.505 140.890 ;
        RECT 102.525 140.020 102.955 140.805 ;
        RECT 103.445 139.980 104.795 140.890 ;
        RECT 105.185 140.210 114.465 140.890 ;
        RECT 105.185 140.090 107.520 140.210 ;
        RECT 105.185 139.980 106.105 140.090 ;
        RECT 112.185 139.990 113.105 140.210 ;
        RECT 114.475 140.080 115.845 140.890 ;
      LAYER nwell ;
        RECT 10.320 136.860 116.040 139.690 ;
      LAYER pwell ;
        RECT 10.515 135.660 11.885 136.470 ;
        RECT 12.365 135.745 12.795 136.530 ;
        RECT 14.175 136.340 15.095 136.560 ;
        RECT 21.175 136.460 22.095 136.570 ;
        RECT 28.675 136.480 29.625 136.570 ;
        RECT 19.760 136.340 22.095 136.460 ;
        RECT 12.815 135.660 22.095 136.340 ;
        RECT 22.475 135.660 25.225 136.470 ;
        RECT 25.235 135.660 26.605 136.440 ;
        RECT 27.695 135.660 29.625 136.480 ;
        RECT 29.835 136.370 30.780 136.570 ;
        RECT 33.055 136.370 34.000 136.570 ;
        RECT 29.835 135.690 32.585 136.370 ;
        RECT 33.055 135.690 35.805 136.370 ;
        RECT 29.835 135.660 30.780 135.690 ;
        RECT 10.655 135.450 10.825 135.660 ;
        RECT 12.090 135.500 12.210 135.610 ;
        RECT 12.495 135.495 12.655 135.605 ;
        RECT 12.955 135.450 13.125 135.660 ;
        RECT 14.335 135.450 14.505 135.640 ;
        RECT 24.915 135.450 25.085 135.660 ;
        RECT 26.110 135.450 26.280 135.640 ;
        RECT 26.295 135.470 26.465 135.660 ;
        RECT 27.695 135.640 27.845 135.660 ;
        RECT 27.215 135.505 27.375 135.615 ;
        RECT 27.675 135.470 27.845 135.640 ;
        RECT 31.355 135.450 31.525 135.640 ;
        RECT 32.270 135.470 32.440 135.690 ;
        RECT 33.055 135.660 34.000 135.690 ;
        RECT 32.790 135.500 32.910 135.610 ;
        RECT 10.515 134.640 11.885 135.450 ;
        RECT 12.815 134.670 14.185 135.450 ;
        RECT 14.205 134.540 15.555 135.450 ;
        RECT 15.945 134.770 25.225 135.450 ;
        RECT 15.945 134.650 18.280 134.770 ;
        RECT 15.945 134.540 16.865 134.650 ;
        RECT 22.945 134.550 23.865 134.770 ;
        RECT 25.245 134.580 25.675 135.365 ;
        RECT 25.695 134.770 29.595 135.450 ;
        RECT 25.695 134.540 26.625 134.770 ;
        RECT 29.835 134.640 31.665 135.450 ;
        RECT 31.675 135.420 32.620 135.450 ;
        RECT 34.110 135.420 34.280 135.640 ;
        RECT 34.575 135.470 34.745 135.640 ;
        RECT 35.490 135.470 35.660 135.690 ;
        RECT 36.275 135.660 38.105 136.470 ;
        RECT 38.125 135.745 38.555 136.530 ;
        RECT 38.575 135.660 44.085 136.470 ;
        RECT 44.095 135.660 45.465 136.440 ;
        RECT 45.475 136.340 46.405 136.570 ;
        RECT 45.475 135.660 49.375 136.340 ;
        RECT 49.615 135.660 53.090 136.570 ;
        RECT 53.295 135.660 56.770 136.570 ;
        RECT 56.975 135.660 58.805 136.470 ;
        RECT 58.825 135.660 60.175 136.570 ;
        RECT 60.195 135.660 63.405 136.570 ;
        RECT 63.885 135.745 64.315 136.530 ;
        RECT 64.795 135.660 67.545 136.470 ;
        RECT 67.555 135.660 73.065 136.470 ;
        RECT 73.075 135.660 78.585 136.470 ;
        RECT 78.965 136.460 79.885 136.570 ;
        RECT 78.965 136.340 81.300 136.460 ;
        RECT 85.965 136.340 86.885 136.560 ;
        RECT 78.965 135.660 88.245 136.340 ;
        RECT 88.255 135.660 89.625 136.440 ;
        RECT 89.645 135.745 90.075 136.530 ;
        RECT 90.465 136.460 91.385 136.570 ;
        RECT 90.465 136.340 92.800 136.460 ;
        RECT 97.465 136.340 98.385 136.560 ;
        RECT 102.425 136.460 103.345 136.570 ;
        RECT 90.465 135.660 99.745 136.340 ;
        RECT 99.755 135.660 101.125 136.440 ;
        RECT 102.425 136.340 104.760 136.460 ;
        RECT 109.425 136.340 110.345 136.560 ;
        RECT 102.425 135.660 111.705 136.340 ;
        RECT 111.715 135.660 113.085 136.440 ;
        RECT 113.095 135.660 114.465 136.470 ;
        RECT 114.475 135.660 115.845 136.470 ;
        RECT 36.010 135.500 36.130 135.610 ;
        RECT 37.795 135.470 37.965 135.660 ;
        RECT 43.775 135.640 43.945 135.660 ;
        RECT 34.595 135.450 34.745 135.470 ;
        RECT 40.095 135.450 40.265 135.640 ;
        RECT 40.555 135.470 40.725 135.640 ;
        RECT 43.315 135.495 43.475 135.605 ;
        RECT 43.775 135.470 43.950 135.640 ;
        RECT 45.155 135.470 45.325 135.660 ;
        RECT 45.890 135.470 46.060 135.660 ;
        RECT 40.575 135.450 40.725 135.470 ;
        RECT 43.780 135.450 43.950 135.470 ;
        RECT 47.460 135.450 47.630 135.640 ;
        RECT 49.760 135.470 49.930 135.660 ;
        RECT 53.440 135.640 53.610 135.660 ;
        RECT 52.975 135.450 53.145 135.640 ;
        RECT 53.435 135.470 53.610 135.640 ;
        RECT 58.495 135.470 58.665 135.660 ;
        RECT 58.955 135.470 59.125 135.660 ;
        RECT 60.335 135.470 60.505 135.660 ;
        RECT 63.610 135.500 63.730 135.610 ;
        RECT 64.530 135.500 64.650 135.610 ;
        RECT 53.435 135.450 53.605 135.470 ;
        RECT 66.315 135.450 66.485 135.640 ;
        RECT 67.235 135.470 67.405 135.660 ;
        RECT 67.695 135.450 67.865 135.640 ;
        RECT 68.155 135.470 68.325 135.640 ;
        RECT 68.175 135.450 68.325 135.470 ;
        RECT 72.295 135.470 72.465 135.640 ;
        RECT 72.755 135.610 72.925 135.660 ;
        RECT 72.755 135.500 72.930 135.610 ;
        RECT 72.755 135.470 72.925 135.500 ;
        RECT 72.295 135.450 72.445 135.470 ;
        RECT 76.435 135.450 76.605 135.640 ;
        RECT 78.275 135.450 78.445 135.660 ;
        RECT 81.955 135.450 82.125 135.640 ;
        RECT 83.335 135.450 83.505 135.640 ;
        RECT 87.015 135.450 87.185 135.640 ;
        RECT 31.675 134.740 34.425 135.420 ;
        RECT 31.675 134.540 32.620 134.740 ;
        RECT 34.595 134.630 36.525 135.450 ;
        RECT 36.735 134.640 40.405 135.450 ;
        RECT 40.575 134.630 42.505 135.450 ;
        RECT 35.575 134.540 36.525 134.630 ;
        RECT 41.555 134.540 42.505 134.630 ;
        RECT 43.635 134.540 47.110 135.450 ;
        RECT 47.315 134.540 50.790 135.450 ;
        RECT 51.005 134.580 51.435 135.365 ;
        RECT 51.455 134.640 53.285 135.450 ;
        RECT 53.405 134.770 56.870 135.450 ;
        RECT 55.950 134.540 56.870 134.770 ;
        RECT 57.345 134.770 66.625 135.450 ;
        RECT 57.345 134.650 59.680 134.770 ;
        RECT 57.345 134.540 58.265 134.650 ;
        RECT 64.345 134.550 65.265 134.770 ;
        RECT 66.635 134.640 68.005 135.450 ;
        RECT 68.175 134.630 70.105 135.450 ;
        RECT 69.155 134.540 70.105 134.630 ;
        RECT 70.515 134.630 72.445 135.450 ;
        RECT 73.075 134.640 76.745 135.450 ;
        RECT 70.515 134.540 71.465 134.630 ;
        RECT 76.765 134.580 77.195 135.365 ;
        RECT 77.215 134.640 78.585 135.450 ;
        RECT 78.595 134.640 82.265 135.450 ;
        RECT 82.285 134.540 83.635 135.450 ;
        RECT 83.655 134.640 87.325 135.450 ;
        RECT 87.480 135.420 87.650 135.640 ;
        RECT 87.935 135.470 88.105 135.660 ;
        RECT 89.315 135.470 89.485 135.660 ;
        RECT 90.695 135.495 90.855 135.605 ;
        RECT 91.155 135.450 91.325 135.640 ;
        RECT 92.590 135.500 92.710 135.610 ;
        RECT 89.140 135.420 90.085 135.450 ;
        RECT 87.335 134.740 90.085 135.420 ;
        RECT 89.140 134.540 90.085 134.740 ;
        RECT 91.025 134.540 92.375 135.450 ;
        RECT 93.000 135.420 93.170 135.640 ;
        RECT 95.760 135.450 95.930 135.640 ;
        RECT 99.435 135.470 99.605 135.660 ;
        RECT 100.815 135.470 100.985 135.660 ;
        RECT 94.660 135.420 95.605 135.450 ;
        RECT 92.855 134.740 95.605 135.420 ;
        RECT 94.660 134.540 95.605 134.740 ;
        RECT 95.615 134.540 99.090 135.450 ;
        RECT 99.295 135.420 100.240 135.450 ;
        RECT 101.730 135.420 101.900 135.640 ;
        RECT 102.250 135.500 102.370 135.610 ;
        RECT 106.520 135.450 106.690 135.640 ;
        RECT 107.310 135.500 107.430 135.610 ;
        RECT 107.715 135.450 107.885 135.640 ;
        RECT 111.395 135.470 111.565 135.660 ;
        RECT 111.855 135.470 112.025 135.660 ;
        RECT 114.155 135.450 114.325 135.660 ;
        RECT 115.535 135.450 115.705 135.660 ;
        RECT 99.295 134.740 102.045 135.420 ;
        RECT 99.295 134.540 100.240 134.740 ;
        RECT 102.525 134.580 102.955 135.365 ;
        RECT 103.205 134.770 107.105 135.450 ;
        RECT 106.175 134.540 107.105 134.770 ;
        RECT 107.575 134.670 108.945 135.450 ;
        RECT 108.955 134.640 114.465 135.450 ;
        RECT 114.475 134.640 115.845 135.450 ;
      LAYER nwell ;
        RECT 10.320 131.420 116.040 134.250 ;
      LAYER pwell ;
        RECT 10.515 130.220 11.885 131.030 ;
        RECT 12.365 130.305 12.795 131.090 ;
        RECT 16.015 130.900 16.945 131.130 ;
        RECT 13.045 130.220 16.945 130.900 ;
        RECT 16.955 130.900 17.885 131.130 ;
        RECT 27.755 131.040 28.705 131.130 ;
        RECT 16.955 130.220 20.855 130.900 ;
        RECT 21.095 130.220 26.605 131.030 ;
        RECT 26.775 130.220 28.705 131.040 ;
        RECT 28.915 130.900 29.845 131.130 ;
        RECT 28.915 130.220 32.815 130.900 ;
        RECT 33.055 130.220 34.425 131.030 ;
        RECT 34.435 130.220 38.105 131.030 ;
        RECT 38.125 130.305 38.555 131.090 ;
        RECT 42.015 131.040 42.965 131.130 ;
        RECT 39.035 130.220 40.865 131.030 ;
        RECT 41.035 130.220 42.965 131.040 ;
        RECT 44.535 130.900 45.455 131.120 ;
        RECT 51.535 131.020 52.455 131.130 ;
        RECT 62.715 131.040 63.665 131.130 ;
        RECT 50.120 130.900 52.455 131.020 ;
        RECT 43.175 130.220 52.455 130.900 ;
        RECT 52.835 130.220 54.205 131.030 ;
        RECT 54.215 130.220 59.725 131.030 ;
        RECT 59.735 130.220 61.565 130.900 ;
        RECT 61.735 130.220 63.665 131.040 ;
        RECT 63.885 130.305 64.315 131.090 ;
        RECT 66.375 131.040 67.325 131.130 ;
        RECT 68.675 131.040 69.625 131.130 ;
        RECT 64.335 130.220 66.165 130.900 ;
        RECT 66.375 130.220 68.305 131.040 ;
        RECT 68.675 130.220 70.605 131.040 ;
        RECT 74.895 130.900 75.825 131.130 ;
        RECT 71.925 130.220 75.825 130.900 ;
        RECT 75.835 130.220 78.585 131.030 ;
        RECT 78.595 130.220 84.105 131.030 ;
        RECT 84.115 130.220 89.625 131.030 ;
        RECT 89.645 130.305 90.075 131.090 ;
        RECT 98.135 131.040 99.085 131.130 ;
        RECT 90.095 130.220 91.465 131.030 ;
        RECT 91.475 130.220 96.985 131.030 ;
        RECT 97.155 130.220 99.085 131.040 ;
        RECT 99.495 131.040 100.445 131.130 ;
        RECT 99.495 130.220 101.425 131.040 ;
        RECT 101.595 130.220 103.425 131.030 ;
        RECT 103.435 130.220 108.945 131.030 ;
        RECT 108.955 130.220 114.465 131.030 ;
        RECT 114.475 130.220 115.845 131.030 ;
        RECT 10.655 130.010 10.825 130.220 ;
        RECT 12.090 130.060 12.210 130.170 ;
        RECT 12.495 130.055 12.655 130.165 ;
        RECT 12.955 130.010 13.125 130.200 ;
        RECT 16.360 130.030 16.530 130.220 ;
        RECT 17.370 130.030 17.540 130.220 ;
        RECT 24.915 130.010 25.085 130.200 ;
        RECT 25.835 130.010 26.005 130.200 ;
        RECT 26.295 130.030 26.465 130.220 ;
        RECT 26.775 130.200 26.925 130.220 ;
        RECT 26.755 130.030 26.925 130.200 ;
        RECT 29.330 130.030 29.500 130.220 ;
        RECT 34.115 130.030 34.285 130.220 ;
        RECT 35.550 130.060 35.670 130.170 ;
        RECT 35.955 130.030 36.125 130.200 ;
        RECT 37.795 130.030 37.965 130.220 ;
        RECT 38.770 130.060 38.890 130.170 ;
        RECT 40.095 130.030 40.265 130.200 ;
        RECT 40.555 130.030 40.725 130.220 ;
        RECT 41.035 130.200 41.185 130.220 ;
        RECT 41.015 130.030 41.185 130.200 ;
        RECT 43.315 130.030 43.485 130.220 ;
        RECT 35.975 130.010 36.125 130.030 ;
        RECT 40.095 130.010 40.245 130.030 ;
        RECT 10.515 129.200 11.885 130.010 ;
        RECT 12.815 129.330 22.095 130.010 ;
        RECT 14.175 129.110 15.095 129.330 ;
        RECT 19.760 129.210 22.095 129.330 ;
        RECT 21.175 129.100 22.095 129.210 ;
        RECT 22.475 129.200 25.225 130.010 ;
        RECT 25.245 129.140 25.675 129.925 ;
        RECT 25.695 129.330 34.975 130.010 ;
        RECT 27.055 129.110 27.975 129.330 ;
        RECT 32.640 129.210 34.975 129.330 ;
        RECT 34.055 129.100 34.975 129.210 ;
        RECT 35.975 129.190 37.905 130.010 ;
        RECT 36.955 129.100 37.905 129.190 ;
        RECT 38.315 129.190 40.245 130.010 ;
        RECT 40.575 130.010 40.725 130.030 ;
        RECT 45.155 130.010 45.325 130.200 ;
        RECT 46.535 130.010 46.705 130.200 ;
        RECT 50.400 130.010 50.570 130.200 ;
        RECT 51.650 130.060 51.770 130.170 ;
        RECT 53.435 130.010 53.605 130.200 ;
        RECT 53.895 130.010 54.065 130.220 ;
        RECT 55.330 130.060 55.450 130.170 ;
        RECT 55.735 130.010 55.905 130.200 ;
        RECT 58.495 130.010 58.665 130.200 ;
        RECT 59.415 130.030 59.585 130.220 ;
        RECT 61.255 130.030 61.425 130.220 ;
        RECT 61.735 130.200 61.885 130.220 ;
        RECT 61.715 130.030 61.885 130.200 ;
        RECT 64.015 130.010 64.185 130.200 ;
        RECT 64.475 130.010 64.645 130.220 ;
        RECT 68.155 130.200 68.305 130.220 ;
        RECT 70.455 130.200 70.605 130.220 ;
        RECT 68.155 130.030 68.325 130.200 ;
        RECT 70.455 130.030 70.625 130.200 ;
        RECT 71.375 130.065 71.535 130.175 ;
        RECT 75.240 130.030 75.410 130.220 ;
        RECT 76.435 130.010 76.605 130.200 ;
        RECT 78.275 130.010 78.445 130.220 ;
        RECT 78.790 130.060 78.910 130.170 ;
        RECT 80.575 130.010 80.745 130.200 ;
        RECT 83.795 130.030 83.965 130.220 ;
        RECT 84.440 130.010 84.610 130.200 ;
        RECT 85.230 130.060 85.350 130.170 ;
        RECT 86.555 130.010 86.725 130.200 ;
        RECT 87.015 130.030 87.185 130.200 ;
        RECT 89.315 130.170 89.485 130.220 ;
        RECT 89.315 130.060 89.490 130.170 ;
        RECT 89.315 130.030 89.485 130.060 ;
        RECT 91.155 130.030 91.325 130.220 ;
        RECT 87.035 130.010 87.185 130.030 ;
        RECT 92.995 130.010 93.165 130.200 ;
        RECT 95.295 130.030 95.465 130.200 ;
        RECT 95.810 130.060 95.930 130.170 ;
        RECT 96.675 130.030 96.845 130.220 ;
        RECT 97.155 130.200 97.305 130.220 ;
        RECT 101.275 130.200 101.425 130.220 ;
        RECT 97.135 130.030 97.305 130.200 ;
        RECT 98.055 130.030 98.225 130.200 ;
        RECT 101.275 130.030 101.445 130.200 ;
        RECT 95.295 130.010 95.445 130.030 ;
        RECT 98.055 130.010 98.205 130.030 ;
        RECT 101.920 130.010 102.090 130.200 ;
        RECT 103.115 130.030 103.285 130.220 ;
        RECT 104.955 130.030 105.125 130.200 ;
        RECT 104.955 130.010 105.105 130.030 ;
        RECT 106.335 130.010 106.505 130.200 ;
        RECT 106.795 130.010 106.965 130.200 ;
        RECT 108.230 130.060 108.350 130.170 ;
        RECT 108.635 130.010 108.805 130.220 ;
        RECT 110.475 130.055 110.635 130.165 ;
        RECT 114.155 130.010 114.325 130.220 ;
        RECT 115.535 130.010 115.705 130.220 ;
        RECT 40.575 129.190 42.505 130.010 ;
        RECT 42.725 129.330 45.465 130.010 ;
        RECT 38.315 129.100 39.265 129.190 ;
        RECT 41.555 129.100 42.505 129.190 ;
        RECT 45.485 129.100 46.835 130.010 ;
        RECT 47.085 129.330 50.985 130.010 ;
        RECT 50.055 129.100 50.985 129.330 ;
        RECT 51.005 129.140 51.435 129.925 ;
        RECT 51.915 129.200 53.745 130.010 ;
        RECT 53.765 129.100 55.115 130.010 ;
        RECT 55.595 129.230 56.965 130.010 ;
        RECT 56.975 129.200 58.805 130.010 ;
        RECT 58.815 129.200 64.325 130.010 ;
        RECT 64.335 129.330 67.075 130.010 ;
        RECT 67.465 129.330 76.745 130.010 ;
        RECT 67.465 129.210 69.800 129.330 ;
        RECT 67.465 129.100 68.385 129.210 ;
        RECT 74.465 129.110 75.385 129.330 ;
        RECT 76.765 129.140 77.195 129.925 ;
        RECT 77.215 129.230 78.585 130.010 ;
        RECT 79.055 129.200 80.885 130.010 ;
        RECT 81.125 129.330 85.025 130.010 ;
        RECT 84.095 129.100 85.025 129.330 ;
        RECT 85.495 129.230 86.865 130.010 ;
        RECT 87.035 129.190 88.965 130.010 ;
        RECT 89.635 129.200 93.305 130.010 ;
        RECT 88.015 129.100 88.965 129.190 ;
        RECT 93.515 129.190 95.445 130.010 ;
        RECT 96.275 129.190 98.205 130.010 ;
        RECT 98.605 129.330 102.505 130.010 ;
        RECT 93.515 129.100 94.465 129.190 ;
        RECT 96.275 129.100 97.225 129.190 ;
        RECT 101.575 129.100 102.505 129.330 ;
        RECT 102.525 129.140 102.955 129.925 ;
        RECT 103.175 129.190 105.105 130.010 ;
        RECT 105.275 129.200 106.645 130.010 ;
        RECT 103.175 129.100 104.125 129.190 ;
        RECT 106.665 129.100 108.015 130.010 ;
        RECT 108.495 129.230 109.865 130.010 ;
        RECT 110.795 129.200 114.465 130.010 ;
        RECT 114.475 129.200 115.845 130.010 ;
      LAYER nwell ;
        RECT 10.320 125.980 116.040 128.810 ;
      LAYER pwell ;
        RECT 10.515 124.780 11.885 125.590 ;
        RECT 12.365 124.865 12.795 125.650 ;
        RECT 12.815 124.780 14.645 125.590 ;
        RECT 14.665 124.780 16.015 125.690 ;
        RECT 16.035 124.780 17.405 125.560 ;
        RECT 17.415 125.460 18.345 125.690 ;
        RECT 17.415 124.780 21.315 125.460 ;
        RECT 21.555 124.780 22.925 125.560 ;
        RECT 22.935 124.780 26.605 125.590 ;
        RECT 26.625 124.780 27.975 125.690 ;
        RECT 28.005 124.780 29.355 125.690 ;
        RECT 31.895 125.600 32.845 125.690 ;
        RECT 29.375 124.780 30.745 125.560 ;
        RECT 30.915 124.780 32.845 125.600 ;
        RECT 36.255 125.460 37.185 125.690 ;
        RECT 33.285 124.780 37.185 125.460 ;
        RECT 38.125 124.865 38.555 125.650 ;
        RECT 41.555 125.600 42.505 125.690 ;
        RECT 38.575 124.780 40.405 125.590 ;
        RECT 40.575 124.780 42.505 125.600 ;
        RECT 43.645 124.780 44.995 125.690 ;
        RECT 45.015 124.780 50.525 125.590 ;
        RECT 50.905 125.580 51.825 125.690 ;
        RECT 50.905 125.460 53.240 125.580 ;
        RECT 57.905 125.460 58.825 125.680 ;
        RECT 50.905 124.780 60.185 125.460 ;
        RECT 60.195 124.780 63.865 125.590 ;
        RECT 63.885 124.865 64.315 125.650 ;
        RECT 64.795 124.780 68.465 125.590 ;
        RECT 71.675 125.460 72.605 125.690 ;
        RECT 68.705 124.780 72.605 125.460 ;
        RECT 72.615 124.780 74.445 125.590 ;
        RECT 74.465 124.780 75.815 125.690 ;
        RECT 76.295 124.780 78.125 125.590 ;
        RECT 81.335 125.460 82.255 125.680 ;
        RECT 88.335 125.580 89.255 125.690 ;
        RECT 86.920 125.460 89.255 125.580 ;
        RECT 78.135 124.780 79.500 125.460 ;
        RECT 79.975 124.780 89.255 125.460 ;
        RECT 89.645 124.865 90.075 125.650 ;
        RECT 90.555 124.780 92.385 125.590 ;
        RECT 92.405 124.780 93.755 125.690 ;
        RECT 96.975 125.460 97.905 125.690 ;
        RECT 94.005 124.780 97.905 125.460 ;
        RECT 97.915 124.780 99.745 125.590 ;
        RECT 102.955 125.460 103.885 125.690 ;
        RECT 99.985 124.780 103.885 125.460 ;
        RECT 104.265 125.580 105.185 125.690 ;
        RECT 104.265 125.460 106.600 125.580 ;
        RECT 111.265 125.460 112.185 125.680 ;
        RECT 104.265 124.780 113.545 125.460 ;
        RECT 114.475 124.780 115.845 125.590 ;
        RECT 10.655 124.570 10.825 124.780 ;
        RECT 12.090 124.620 12.210 124.730 ;
        RECT 12.955 124.570 13.125 124.760 ;
        RECT 14.335 124.570 14.505 124.780 ;
        RECT 14.795 124.590 14.965 124.780 ;
        RECT 15.715 124.570 15.885 124.760 ;
        RECT 17.095 124.590 17.265 124.780 ;
        RECT 17.830 124.590 18.000 124.780 ;
        RECT 22.615 124.590 22.785 124.780 ;
        RECT 24.915 124.570 25.085 124.760 ;
        RECT 26.295 124.590 26.465 124.780 ;
        RECT 26.755 124.590 26.925 124.780 ;
        RECT 28.135 124.590 28.305 124.780 ;
        RECT 30.160 124.570 30.330 124.760 ;
        RECT 30.435 124.590 30.605 124.780 ;
        RECT 30.915 124.760 31.065 124.780 ;
        RECT 30.895 124.590 31.065 124.760 ;
        RECT 36.600 124.590 36.770 124.780 ;
        RECT 37.795 124.625 37.955 124.735 ;
        RECT 40.095 124.570 40.265 124.780 ;
        RECT 40.575 124.760 40.725 124.780 ;
        RECT 40.555 124.590 40.725 124.760 ;
        RECT 43.315 124.625 43.475 124.735 ;
        RECT 43.775 124.590 43.945 124.780 ;
        RECT 49.755 124.570 49.925 124.760 ;
        RECT 50.215 124.590 50.385 124.780 ;
        RECT 50.675 124.615 50.835 124.725 ;
        RECT 51.595 124.570 51.765 124.760 ;
        RECT 53.435 124.615 53.595 124.725 ;
        RECT 54.170 124.570 54.340 124.760 ;
        RECT 59.875 124.590 60.045 124.780 ;
        RECT 61.440 124.570 61.610 124.760 ;
        RECT 63.555 124.590 63.725 124.780 ;
        RECT 64.530 124.620 64.650 124.730 ;
        RECT 65.395 124.570 65.565 124.760 ;
        RECT 68.155 124.590 68.325 124.780 ;
        RECT 72.020 124.590 72.190 124.780 ;
        RECT 74.135 124.590 74.305 124.780 ;
        RECT 75.055 124.570 75.225 124.760 ;
        RECT 75.515 124.590 75.685 124.780 ;
        RECT 76.030 124.620 76.150 124.730 ;
        RECT 76.435 124.570 76.605 124.760 ;
        RECT 77.815 124.590 77.985 124.780 ;
        RECT 79.655 124.590 79.825 124.760 ;
        RECT 80.115 124.590 80.285 124.780 ;
        RECT 86.095 124.570 86.265 124.760 ;
        RECT 86.610 124.620 86.730 124.730 ;
        RECT 90.290 124.620 90.410 124.730 ;
        RECT 90.420 124.570 90.590 124.760 ;
        RECT 92.075 124.570 92.245 124.780 ;
        RECT 92.535 124.590 92.705 124.780 ;
        RECT 92.995 124.615 93.155 124.725 ;
        RECT 93.455 124.570 93.625 124.760 ;
        RECT 97.320 124.590 97.490 124.780 ;
        RECT 99.435 124.590 99.605 124.780 ;
        RECT 103.170 124.620 103.290 124.730 ;
        RECT 103.300 124.590 103.470 124.780 ;
        RECT 112.775 124.570 112.945 124.760 ;
        RECT 113.235 124.590 113.405 124.780 ;
        RECT 114.155 124.570 114.325 124.760 ;
        RECT 115.535 124.570 115.705 124.780 ;
        RECT 10.515 123.760 11.885 124.570 ;
        RECT 11.895 123.760 13.265 124.570 ;
        RECT 13.285 123.660 14.635 124.570 ;
        RECT 14.655 123.790 16.025 124.570 ;
        RECT 16.120 123.890 25.225 124.570 ;
        RECT 25.245 123.700 25.675 124.485 ;
        RECT 26.845 123.890 30.745 124.570 ;
        RECT 29.815 123.660 30.745 123.890 ;
        RECT 31.125 123.890 40.405 124.570 ;
        RECT 40.785 123.890 50.065 124.570 ;
        RECT 31.125 123.770 33.460 123.890 ;
        RECT 31.125 123.660 32.045 123.770 ;
        RECT 38.125 123.670 39.045 123.890 ;
        RECT 40.785 123.770 43.120 123.890 ;
        RECT 40.785 123.660 41.705 123.770 ;
        RECT 47.785 123.670 48.705 123.890 ;
        RECT 51.005 123.700 51.435 124.485 ;
        RECT 51.455 123.790 52.825 124.570 ;
        RECT 53.755 123.890 57.655 124.570 ;
        RECT 58.125 123.890 62.025 124.570 ;
        RECT 53.755 123.660 54.685 123.890 ;
        RECT 61.095 123.660 62.025 123.890 ;
        RECT 62.035 123.760 65.705 124.570 ;
        RECT 66.085 123.890 75.365 124.570 ;
        RECT 66.085 123.770 68.420 123.890 ;
        RECT 66.085 123.660 67.005 123.770 ;
        RECT 73.085 123.670 74.005 123.890 ;
        RECT 75.375 123.790 76.745 124.570 ;
        RECT 76.765 123.700 77.195 124.485 ;
        RECT 77.300 123.890 86.405 124.570 ;
        RECT 87.105 123.890 91.005 124.570 ;
        RECT 90.075 123.660 91.005 123.890 ;
        RECT 91.025 123.660 92.375 124.570 ;
        RECT 93.315 123.890 102.420 124.570 ;
        RECT 102.525 123.700 102.955 124.485 ;
        RECT 103.805 123.890 113.085 124.570 ;
        RECT 103.805 123.770 106.140 123.890 ;
        RECT 103.805 123.660 104.725 123.770 ;
        RECT 110.805 123.670 111.725 123.890 ;
        RECT 113.095 123.790 114.465 124.570 ;
        RECT 114.475 123.760 115.845 124.570 ;
      LAYER nwell ;
        RECT 10.320 120.540 116.040 123.370 ;
      LAYER pwell ;
        RECT 10.515 119.340 11.885 120.150 ;
        RECT 12.365 119.425 12.795 120.210 ;
        RECT 14.635 120.020 15.555 120.240 ;
        RECT 21.635 120.140 22.555 120.250 ;
        RECT 20.220 120.020 22.555 120.140 ;
        RECT 13.275 119.340 22.555 120.020 ;
        RECT 22.935 120.020 23.865 120.250 ;
        RECT 27.905 120.140 28.825 120.250 ;
        RECT 27.905 120.020 30.240 120.140 ;
        RECT 34.905 120.020 35.825 120.240 ;
        RECT 22.935 119.340 26.835 120.020 ;
        RECT 27.905 119.340 37.185 120.020 ;
        RECT 38.125 119.425 38.555 120.210 ;
        RECT 39.035 119.340 40.405 120.120 ;
        RECT 40.415 119.340 41.785 120.150 ;
        RECT 41.815 119.340 52.825 120.250 ;
        RECT 52.845 119.340 54.195 120.250 ;
        RECT 54.585 120.140 55.505 120.250 ;
        RECT 54.585 120.020 56.920 120.140 ;
        RECT 61.585 120.020 62.505 120.240 ;
        RECT 54.585 119.340 63.865 120.020 ;
        RECT 63.885 119.425 64.315 120.210 ;
        RECT 64.335 119.340 65.705 120.120 ;
        RECT 65.715 119.340 68.465 120.150 ;
        RECT 68.485 119.340 69.835 120.250 ;
        RECT 73.055 120.020 73.985 120.250 ;
        RECT 70.085 119.340 73.985 120.020 ;
        RECT 73.995 119.340 75.825 120.150 ;
        RECT 79.035 120.020 79.965 120.250 ;
        RECT 76.065 119.340 79.965 120.020 ;
        RECT 80.345 120.140 81.265 120.250 ;
        RECT 80.345 120.020 82.680 120.140 ;
        RECT 87.345 120.020 88.265 120.240 ;
        RECT 80.345 119.340 89.625 120.020 ;
        RECT 89.645 119.425 90.075 120.210 ;
        RECT 90.465 120.140 91.385 120.250 ;
        RECT 90.465 120.020 92.800 120.140 ;
        RECT 97.465 120.020 98.385 120.240 ;
        RECT 100.125 120.140 101.045 120.250 ;
        RECT 100.125 120.020 102.460 120.140 ;
        RECT 107.125 120.020 108.045 120.240 ;
        RECT 90.465 119.340 99.745 120.020 ;
        RECT 100.125 119.340 109.405 120.020 ;
        RECT 109.415 119.340 110.785 120.150 ;
        RECT 110.795 119.340 114.465 120.150 ;
        RECT 114.475 119.340 115.845 120.150 ;
        RECT 10.655 119.130 10.825 119.340 ;
        RECT 12.090 119.180 12.210 119.290 ;
        RECT 13.010 119.180 13.130 119.290 ;
        RECT 13.415 119.130 13.585 119.340 ;
        RECT 13.875 119.130 14.045 119.320 ;
        RECT 23.350 119.150 23.520 119.340 ;
        RECT 24.915 119.130 25.085 119.320 ;
        RECT 27.270 119.180 27.390 119.290 ;
        RECT 35.035 119.130 35.205 119.320 ;
        RECT 36.415 119.130 36.585 119.320 ;
        RECT 36.875 119.150 37.045 119.340 ;
        RECT 37.335 119.175 37.495 119.285 ;
        RECT 37.795 119.185 37.955 119.295 ;
        RECT 38.770 119.180 38.890 119.290 ;
        RECT 40.095 119.150 40.265 119.340 ;
        RECT 41.200 119.130 41.370 119.320 ;
        RECT 41.475 119.150 41.645 119.340 ;
        RECT 52.510 119.320 52.680 119.340 ;
        RECT 41.935 119.130 42.105 119.320 ;
        RECT 52.510 119.150 52.685 119.320 ;
        RECT 52.975 119.290 53.145 119.340 ;
        RECT 52.975 119.180 53.150 119.290 ;
        RECT 52.975 119.150 53.145 119.180 ;
        RECT 52.515 119.130 52.685 119.150 ;
        RECT 53.435 119.130 53.605 119.320 ;
        RECT 63.555 119.150 63.725 119.340 ;
        RECT 65.395 119.130 65.565 119.340 ;
        RECT 68.155 119.150 68.325 119.340 ;
        RECT 68.615 119.150 68.785 119.340 ;
        RECT 73.400 119.150 73.570 119.340 ;
        RECT 75.055 119.130 75.225 119.320 ;
        RECT 75.515 119.130 75.685 119.340 ;
        RECT 79.380 119.150 79.550 119.340 ;
        RECT 86.555 119.130 86.725 119.320 ;
        RECT 87.935 119.130 88.105 119.320 ;
        RECT 88.450 119.180 88.570 119.290 ;
        RECT 89.315 119.150 89.485 119.340 ;
        RECT 89.775 119.130 89.945 119.320 ;
        RECT 90.695 119.175 90.855 119.285 ;
        RECT 94.375 119.130 94.545 119.320 ;
        RECT 94.835 119.130 95.005 119.320 ;
        RECT 96.215 119.130 96.385 119.320 ;
        RECT 98.055 119.175 98.215 119.285 ;
        RECT 99.435 119.150 99.605 119.340 ;
        RECT 101.920 119.130 102.090 119.320 ;
        RECT 104.035 119.150 104.205 119.320 ;
        RECT 105.875 119.130 106.045 119.320 ;
        RECT 106.335 119.130 106.505 119.320 ;
        RECT 108.635 119.130 108.805 119.320 ;
        RECT 109.095 119.150 109.265 119.340 ;
        RECT 110.475 119.150 110.645 119.340 ;
        RECT 114.155 119.130 114.325 119.340 ;
        RECT 115.535 119.130 115.705 119.340 ;
        RECT 10.515 118.320 11.885 119.130 ;
        RECT 11.895 118.320 13.725 119.130 ;
        RECT 13.735 118.450 23.015 119.130 ;
        RECT 15.095 118.230 16.015 118.450 ;
        RECT 20.680 118.330 23.015 118.450 ;
        RECT 22.095 118.220 23.015 118.330 ;
        RECT 23.395 118.320 25.225 119.130 ;
        RECT 25.245 118.260 25.675 119.045 ;
        RECT 26.065 118.450 35.345 119.130 ;
        RECT 26.065 118.330 28.400 118.450 ;
        RECT 26.065 118.220 26.985 118.330 ;
        RECT 33.065 118.230 33.985 118.450 ;
        RECT 35.355 118.350 36.725 119.130 ;
        RECT 37.885 118.450 41.785 119.130 ;
        RECT 41.795 118.450 50.900 119.130 ;
        RECT 40.855 118.220 41.785 118.450 ;
        RECT 51.005 118.260 51.435 119.045 ;
        RECT 51.455 118.350 52.825 119.130 ;
        RECT 53.295 118.450 62.575 119.130 ;
        RECT 54.655 118.230 55.575 118.450 ;
        RECT 60.240 118.330 62.575 118.450 ;
        RECT 61.655 118.220 62.575 118.330 ;
        RECT 62.955 118.320 65.705 119.130 ;
        RECT 66.085 118.450 75.365 119.130 ;
        RECT 66.085 118.330 68.420 118.450 ;
        RECT 66.085 118.220 67.005 118.330 ;
        RECT 73.085 118.230 74.005 118.450 ;
        RECT 75.385 118.220 76.735 119.130 ;
        RECT 76.765 118.260 77.195 119.045 ;
        RECT 77.585 118.450 86.865 119.130 ;
        RECT 77.585 118.330 79.920 118.450 ;
        RECT 77.585 118.220 78.505 118.330 ;
        RECT 84.585 118.230 85.505 118.450 ;
        RECT 86.875 118.350 88.245 119.130 ;
        RECT 88.715 118.350 90.085 119.130 ;
        RECT 91.015 118.320 94.685 119.130 ;
        RECT 94.705 118.220 96.055 119.130 ;
        RECT 96.075 118.350 97.445 119.130 ;
        RECT 98.605 118.450 102.505 119.130 ;
        RECT 101.575 118.220 102.505 118.450 ;
        RECT 102.525 118.260 102.955 119.045 ;
        RECT 102.975 118.450 103.930 119.130 ;
        RECT 104.355 118.320 106.185 119.130 ;
        RECT 106.205 118.220 107.555 119.130 ;
        RECT 107.575 118.320 108.945 119.130 ;
        RECT 108.955 118.320 114.465 119.130 ;
        RECT 114.475 118.320 115.845 119.130 ;
      LAYER nwell ;
        RECT 10.320 115.100 116.040 117.930 ;
      LAYER pwell ;
        RECT 10.515 113.900 11.885 114.710 ;
        RECT 12.365 113.985 12.795 114.770 ;
        RECT 13.735 113.900 17.405 114.710 ;
        RECT 17.425 113.900 18.775 114.810 ;
        RECT 19.715 113.900 23.385 114.710 ;
        RECT 23.395 113.900 28.905 114.710 ;
        RECT 28.925 113.900 30.275 114.810 ;
        RECT 30.295 113.900 32.125 114.710 ;
        RECT 32.135 113.900 33.505 114.680 ;
        RECT 37.175 114.580 38.105 114.810 ;
        RECT 34.205 113.900 38.105 114.580 ;
        RECT 38.125 113.985 38.555 114.770 ;
        RECT 38.575 113.900 41.325 114.710 ;
        RECT 41.345 113.900 42.695 114.810 ;
        RECT 43.175 113.900 45.005 114.710 ;
        RECT 45.155 113.900 47.765 114.810 ;
        RECT 47.775 113.900 51.445 114.710 ;
        RECT 51.455 113.900 56.965 114.710 ;
        RECT 56.985 113.900 58.335 114.810 ;
        RECT 58.355 113.900 63.865 114.710 ;
        RECT 63.885 113.985 64.315 114.770 ;
        RECT 65.255 113.900 68.925 114.710 ;
        RECT 68.945 113.900 70.295 114.810 ;
        RECT 70.775 113.900 72.605 114.710 ;
        RECT 72.615 113.900 73.985 114.680 ;
        RECT 73.995 113.900 75.825 114.710 ;
        RECT 75.835 113.900 81.345 114.710 ;
        RECT 81.365 113.900 82.715 114.810 ;
        RECT 82.735 113.900 84.105 114.710 ;
        RECT 84.115 113.900 89.625 114.710 ;
        RECT 89.645 113.985 90.075 114.770 ;
        RECT 90.095 113.900 95.605 114.710 ;
        RECT 95.615 113.900 101.125 114.710 ;
        RECT 101.135 113.900 102.505 114.680 ;
        RECT 102.975 113.900 106.645 114.710 ;
        RECT 106.655 113.900 108.025 114.680 ;
        RECT 108.045 113.900 109.395 114.810 ;
        RECT 110.335 113.900 111.705 114.680 ;
        RECT 111.715 113.900 114.465 114.710 ;
        RECT 114.475 113.900 115.845 114.710 ;
        RECT 10.655 113.690 10.825 113.900 ;
        RECT 12.090 113.740 12.210 113.850 ;
        RECT 12.955 113.690 13.125 113.880 ;
        RECT 13.415 113.745 13.575 113.855 ;
        RECT 16.635 113.690 16.805 113.880 ;
        RECT 17.095 113.710 17.265 113.900 ;
        RECT 18.475 113.710 18.645 113.900 ;
        RECT 19.395 113.745 19.555 113.855 ;
        RECT 22.155 113.690 22.325 113.880 ;
        RECT 23.075 113.710 23.245 113.900 ;
        RECT 23.535 113.690 23.705 113.880 ;
        RECT 24.915 113.690 25.085 113.880 ;
        RECT 25.890 113.740 26.010 113.850 ;
        RECT 28.595 113.710 28.765 113.900 ;
        RECT 29.055 113.710 29.225 113.900 ;
        RECT 31.355 113.690 31.525 113.880 ;
        RECT 31.815 113.690 31.985 113.900 ;
        RECT 32.275 113.710 32.445 113.900 ;
        RECT 33.250 113.740 33.370 113.850 ;
        RECT 33.710 113.740 33.830 113.850 ;
        RECT 36.875 113.690 37.045 113.880 ;
        RECT 37.520 113.710 37.690 113.900 ;
        RECT 38.255 113.690 38.425 113.880 ;
        RECT 41.015 113.710 41.185 113.900 ;
        RECT 42.395 113.710 42.565 113.900 ;
        RECT 42.910 113.740 43.030 113.850 ;
        RECT 43.775 113.690 43.945 113.880 ;
        RECT 44.695 113.710 44.865 113.900 ;
        RECT 47.450 113.710 47.620 113.900 ;
        RECT 49.295 113.690 49.465 113.880 ;
        RECT 49.755 113.690 49.925 113.880 ;
        RECT 51.135 113.710 51.305 113.900 ;
        RECT 52.515 113.690 52.685 113.880 ;
        RECT 52.980 113.690 53.150 113.880 ;
        RECT 56.655 113.710 56.825 113.900 ;
        RECT 57.115 113.690 57.285 113.900 ;
        RECT 62.635 113.690 62.805 113.880 ;
        RECT 63.555 113.710 63.725 113.900 ;
        RECT 64.935 113.745 65.095 113.855 ;
        RECT 68.155 113.690 68.325 113.880 ;
        RECT 68.615 113.690 68.785 113.900 ;
        RECT 69.075 113.710 69.245 113.900 ;
        RECT 69.995 113.690 70.165 113.880 ;
        RECT 70.510 113.740 70.630 113.850 ;
        RECT 71.380 113.690 71.550 113.880 ;
        RECT 72.295 113.710 72.465 113.900 ;
        RECT 73.675 113.710 73.845 113.900 ;
        RECT 75.515 113.710 75.685 113.900 ;
        RECT 76.435 113.690 76.605 113.880 ;
        RECT 77.410 113.740 77.530 113.850 ;
        RECT 79.195 113.690 79.365 113.880 ;
        RECT 81.035 113.710 81.205 113.900 ;
        RECT 81.495 113.710 81.665 113.900 ;
        RECT 83.795 113.710 83.965 113.900 ;
        RECT 84.715 113.690 84.885 113.880 ;
        RECT 85.175 113.690 85.345 113.880 ;
        RECT 89.315 113.710 89.485 113.900 ;
        RECT 89.775 113.690 89.945 113.880 ;
        RECT 90.235 113.690 90.405 113.880 ;
        RECT 91.670 113.740 91.790 113.850 ;
        RECT 95.295 113.690 95.465 113.900 ;
        RECT 95.755 113.690 95.925 113.880 ;
        RECT 99.435 113.690 99.605 113.880 ;
        RECT 99.895 113.690 100.065 113.880 ;
        RECT 100.815 113.710 100.985 113.900 ;
        RECT 101.275 113.690 101.445 113.900 ;
        RECT 102.710 113.740 102.830 113.850 ;
        RECT 103.575 113.735 103.735 113.845 ;
        RECT 104.035 113.690 104.205 113.880 ;
        RECT 106.335 113.710 106.505 113.900 ;
        RECT 107.715 113.710 107.885 113.900 ;
        RECT 108.175 113.710 108.345 113.900 ;
        RECT 110.015 113.745 110.175 113.855 ;
        RECT 111.395 113.710 111.565 113.900 ;
        RECT 114.155 113.710 114.325 113.900 ;
        RECT 115.535 113.690 115.705 113.900 ;
        RECT 10.515 112.880 11.885 113.690 ;
        RECT 11.895 112.880 13.265 113.690 ;
        RECT 13.275 112.880 16.945 113.690 ;
        RECT 16.955 112.880 22.465 113.690 ;
        RECT 22.475 112.910 23.845 113.690 ;
        RECT 23.855 112.880 25.225 113.690 ;
        RECT 25.245 112.820 25.675 113.605 ;
        RECT 26.155 112.880 31.665 113.690 ;
        RECT 31.675 112.910 33.045 113.690 ;
        RECT 33.515 112.880 37.185 113.690 ;
        RECT 37.195 112.910 38.565 113.690 ;
        RECT 38.575 112.880 44.085 113.690 ;
        RECT 44.095 112.880 49.605 113.690 ;
        RECT 49.615 112.910 50.985 113.690 ;
        RECT 51.005 112.820 51.435 113.605 ;
        RECT 51.455 112.880 52.825 113.690 ;
        RECT 52.835 112.780 55.445 113.690 ;
        RECT 55.595 112.880 57.425 113.690 ;
        RECT 57.435 112.880 62.945 113.690 ;
        RECT 62.955 112.880 68.465 113.690 ;
        RECT 68.475 112.910 69.845 113.690 ;
        RECT 69.855 112.910 71.225 113.690 ;
        RECT 71.235 112.780 73.845 113.690 ;
        RECT 73.995 112.880 76.745 113.690 ;
        RECT 76.765 112.820 77.195 113.605 ;
        RECT 77.675 112.880 79.505 113.690 ;
        RECT 79.515 112.880 85.025 113.690 ;
        RECT 85.035 112.910 86.405 113.690 ;
        RECT 86.415 112.880 90.085 113.690 ;
        RECT 90.095 112.910 91.465 113.690 ;
        RECT 91.935 112.880 95.605 113.690 ;
        RECT 95.615 112.910 96.985 113.690 ;
        RECT 96.995 112.880 99.745 113.690 ;
        RECT 99.755 112.910 101.125 113.690 ;
        RECT 101.135 112.910 102.505 113.690 ;
        RECT 102.525 112.820 102.955 113.605 ;
        RECT 103.895 113.010 114.265 113.690 ;
        RECT 108.405 112.790 109.335 113.010 ;
        RECT 112.055 112.780 114.265 113.010 ;
        RECT 114.475 112.880 115.845 113.690 ;
      LAYER nwell ;
        RECT 10.320 109.660 116.040 112.490 ;
      LAYER pwell ;
        RECT 10.515 108.460 11.885 109.270 ;
        RECT 12.365 108.545 12.795 109.330 ;
        RECT 12.815 108.460 14.185 109.270 ;
        RECT 14.395 109.140 16.605 109.370 ;
        RECT 19.325 109.140 20.255 109.360 ;
        RECT 14.395 108.460 24.765 109.140 ;
        RECT 24.775 108.460 26.145 109.240 ;
        RECT 26.155 108.460 27.525 109.240 ;
        RECT 27.735 109.140 29.945 109.370 ;
        RECT 32.665 109.140 33.595 109.360 ;
        RECT 27.735 108.460 38.105 109.140 ;
        RECT 38.125 108.545 38.555 109.330 ;
        RECT 39.505 108.460 40.855 109.370 ;
        RECT 41.335 108.460 42.705 109.240 ;
        RECT 42.715 108.460 44.545 109.270 ;
        RECT 44.555 108.460 45.925 109.240 ;
        RECT 46.135 109.140 48.345 109.370 ;
        RECT 51.065 109.140 51.995 109.360 ;
        RECT 46.135 108.460 56.505 109.140 ;
        RECT 56.975 108.460 58.345 109.240 ;
        RECT 58.365 108.460 59.715 109.370 ;
        RECT 59.735 108.460 61.105 109.270 ;
        RECT 61.115 108.460 62.485 109.240 ;
        RECT 62.495 108.460 63.865 109.270 ;
        RECT 63.885 108.545 64.315 109.330 ;
        RECT 64.795 108.460 66.165 109.240 ;
        RECT 66.185 108.460 67.535 109.370 ;
        RECT 72.065 109.140 72.995 109.360 ;
        RECT 75.715 109.140 77.925 109.370 ;
        RECT 67.555 108.460 77.925 109.140 ;
        RECT 79.255 109.140 81.465 109.370 ;
        RECT 84.185 109.140 85.115 109.360 ;
        RECT 79.255 108.460 89.625 109.140 ;
        RECT 89.645 108.545 90.075 109.330 ;
        RECT 90.295 109.140 92.505 109.370 ;
        RECT 95.225 109.140 96.155 109.360 ;
        RECT 90.295 108.460 100.665 109.140 ;
        RECT 101.135 108.460 103.885 109.270 ;
        RECT 108.405 109.140 109.335 109.360 ;
        RECT 112.055 109.140 114.265 109.370 ;
        RECT 103.895 108.460 114.265 109.140 ;
        RECT 114.475 108.460 115.845 109.270 ;
        RECT 10.655 108.250 10.825 108.460 ;
        RECT 12.090 108.300 12.210 108.410 ;
        RECT 12.955 108.250 13.125 108.440 ;
        RECT 13.415 108.250 13.585 108.440 ;
        RECT 13.875 108.270 14.045 108.460 ;
        RECT 24.455 108.270 24.625 108.460 ;
        RECT 24.915 108.250 25.085 108.440 ;
        RECT 25.835 108.270 26.005 108.460 ;
        RECT 26.755 108.250 26.925 108.440 ;
        RECT 27.215 108.250 27.385 108.460 ;
        RECT 28.595 108.250 28.765 108.440 ;
        RECT 29.975 108.250 30.145 108.440 ;
        RECT 37.795 108.270 37.965 108.460 ;
        RECT 39.175 108.305 39.335 108.415 ;
        RECT 40.555 108.270 40.725 108.460 ;
        RECT 41.070 108.300 41.190 108.410 ;
        RECT 42.395 108.270 42.565 108.460 ;
        RECT 44.235 108.270 44.405 108.460 ;
        RECT 44.695 108.270 44.865 108.460 ;
        RECT 50.675 108.250 50.845 108.440 ;
        RECT 51.650 108.300 51.770 108.410 ;
        RECT 56.195 108.270 56.365 108.460 ;
        RECT 56.710 108.300 56.830 108.410 ;
        RECT 57.115 108.270 57.285 108.460 ;
        RECT 58.495 108.270 58.665 108.460 ;
        RECT 60.795 108.270 60.965 108.460 ;
        RECT 61.255 108.270 61.425 108.460 ;
        RECT 62.175 108.250 62.345 108.440 ;
        RECT 63.095 108.295 63.255 108.405 ;
        RECT 63.555 108.270 63.725 108.460 ;
        RECT 64.530 108.300 64.650 108.410 ;
        RECT 64.935 108.270 65.105 108.460 ;
        RECT 67.235 108.270 67.405 108.460 ;
        RECT 67.695 108.270 67.865 108.460 ;
        RECT 73.675 108.250 73.845 108.440 ;
        RECT 75.055 108.250 75.225 108.440 ;
        RECT 75.515 108.250 75.685 108.440 ;
        RECT 78.735 108.305 78.895 108.415 ;
        RECT 87.475 108.250 87.645 108.440 ;
        RECT 89.315 108.270 89.485 108.460 ;
        RECT 98.055 108.250 98.225 108.440 ;
        RECT 99.435 108.250 99.605 108.440 ;
        RECT 100.355 108.270 100.525 108.460 ;
        RECT 100.815 108.410 100.985 108.440 ;
        RECT 100.815 108.300 100.990 108.410 ;
        RECT 100.815 108.250 100.985 108.300 ;
        RECT 101.275 108.250 101.445 108.440 ;
        RECT 103.575 108.270 103.745 108.460 ;
        RECT 104.035 108.270 104.205 108.460 ;
        RECT 113.235 108.250 113.405 108.440 ;
        RECT 114.155 108.295 114.315 108.405 ;
        RECT 115.535 108.250 115.705 108.460 ;
        RECT 10.515 107.440 11.885 108.250 ;
        RECT 11.905 107.340 13.255 108.250 ;
        RECT 13.285 107.340 14.635 108.250 ;
        RECT 14.855 107.570 25.225 108.250 ;
        RECT 14.855 107.340 17.065 107.570 ;
        RECT 19.785 107.350 20.715 107.570 ;
        RECT 25.245 107.380 25.675 108.165 ;
        RECT 25.705 107.340 27.055 108.250 ;
        RECT 27.085 107.340 28.435 108.250 ;
        RECT 28.465 107.340 29.815 108.250 ;
        RECT 29.835 107.570 40.205 108.250 ;
        RECT 34.345 107.350 35.275 107.570 ;
        RECT 37.995 107.340 40.205 107.570 ;
        RECT 40.615 107.570 50.985 108.250 ;
        RECT 40.615 107.340 42.825 107.570 ;
        RECT 45.545 107.350 46.475 107.570 ;
        RECT 51.005 107.380 51.435 108.165 ;
        RECT 52.115 107.570 62.485 108.250 ;
        RECT 63.615 107.570 73.985 108.250 ;
        RECT 52.115 107.340 54.325 107.570 ;
        RECT 57.045 107.350 57.975 107.570 ;
        RECT 63.615 107.340 65.825 107.570 ;
        RECT 68.545 107.350 69.475 107.570 ;
        RECT 74.005 107.340 75.355 108.250 ;
        RECT 75.385 107.340 76.735 108.250 ;
        RECT 76.765 107.380 77.195 108.165 ;
        RECT 77.415 107.570 87.785 108.250 ;
        RECT 87.995 107.570 98.365 108.250 ;
        RECT 77.415 107.340 79.625 107.570 ;
        RECT 82.345 107.350 83.275 107.570 ;
        RECT 87.995 107.340 90.205 107.570 ;
        RECT 92.925 107.350 93.855 107.570 ;
        RECT 98.385 107.340 99.735 108.250 ;
        RECT 99.765 107.340 101.115 108.250 ;
        RECT 101.145 107.340 102.495 108.250 ;
        RECT 102.525 107.380 102.955 108.165 ;
        RECT 103.175 107.570 113.545 108.250 ;
        RECT 103.175 107.340 105.385 107.570 ;
        RECT 108.105 107.350 109.035 107.570 ;
        RECT 114.475 107.440 115.845 108.250 ;
      LAYER nwell ;
        RECT 10.320 104.220 116.040 107.050 ;
      LAYER pwell ;
        RECT 10.515 103.020 11.885 103.830 ;
        RECT 12.365 103.105 12.795 103.890 ;
        RECT 13.015 103.700 15.225 103.930 ;
        RECT 17.945 103.700 18.875 103.920 ;
        RECT 13.015 103.020 23.385 103.700 ;
        RECT 23.395 103.020 25.225 103.830 ;
        RECT 25.245 103.105 25.675 103.890 ;
        RECT 25.895 103.700 28.105 103.930 ;
        RECT 30.825 103.700 31.755 103.920 ;
        RECT 25.895 103.020 36.265 103.700 ;
        RECT 36.275 103.020 38.105 103.830 ;
        RECT 38.125 103.105 38.555 103.890 ;
        RECT 39.495 103.020 45.005 103.830 ;
        RECT 45.025 103.020 46.375 103.930 ;
        RECT 46.855 103.020 49.605 103.830 ;
        RECT 49.625 103.020 50.975 103.930 ;
        RECT 51.005 103.105 51.435 103.890 ;
        RECT 51.925 103.020 53.275 103.930 ;
        RECT 53.495 103.700 55.705 103.930 ;
        RECT 58.425 103.700 59.355 103.920 ;
        RECT 53.495 103.020 63.865 103.700 ;
        RECT 63.885 103.105 64.315 103.890 ;
        RECT 64.335 103.020 69.845 103.830 ;
        RECT 69.865 103.020 71.215 103.930 ;
        RECT 71.235 103.020 76.745 103.830 ;
        RECT 76.765 103.105 77.195 103.890 ;
        RECT 78.135 103.020 83.645 103.830 ;
        RECT 83.665 103.020 85.015 103.930 ;
        RECT 85.495 103.020 88.245 103.830 ;
        RECT 88.265 103.020 89.615 103.930 ;
        RECT 89.645 103.105 90.075 103.890 ;
        RECT 90.095 103.020 91.925 103.830 ;
        RECT 92.135 103.700 94.345 103.930 ;
        RECT 97.065 103.700 97.995 103.920 ;
        RECT 92.135 103.020 102.505 103.700 ;
        RECT 102.525 103.105 102.955 103.890 ;
        RECT 102.975 103.020 104.345 103.830 ;
        RECT 104.355 103.020 108.025 103.830 ;
        RECT 108.045 103.020 109.395 103.930 ;
        RECT 109.415 103.020 113.085 103.830 ;
        RECT 113.095 103.020 114.465 103.800 ;
        RECT 114.475 103.020 115.845 103.830 ;
        RECT 10.655 102.830 10.825 103.020 ;
        RECT 12.090 102.860 12.210 102.970 ;
        RECT 23.075 102.830 23.245 103.020 ;
        RECT 24.915 102.830 25.085 103.020 ;
        RECT 35.955 102.830 36.125 103.020 ;
        RECT 37.795 102.830 37.965 103.020 ;
        RECT 39.175 102.865 39.335 102.975 ;
        RECT 44.695 102.830 44.865 103.020 ;
        RECT 46.075 102.830 46.245 103.020 ;
        RECT 46.590 102.860 46.710 102.970 ;
        RECT 49.295 102.830 49.465 103.020 ;
        RECT 49.755 102.830 49.925 103.020 ;
        RECT 51.650 102.860 51.770 102.970 ;
        RECT 52.055 102.830 52.225 103.020 ;
        RECT 63.555 102.830 63.725 103.020 ;
        RECT 69.535 102.830 69.705 103.020 ;
        RECT 70.915 102.830 71.085 103.020 ;
        RECT 76.435 102.830 76.605 103.020 ;
        RECT 77.815 102.865 77.975 102.975 ;
        RECT 83.335 102.830 83.505 103.020 ;
        RECT 84.715 102.830 84.885 103.020 ;
        RECT 85.230 102.860 85.350 102.970 ;
        RECT 87.935 102.830 88.105 103.020 ;
        RECT 88.395 102.830 88.565 103.020 ;
        RECT 91.615 102.830 91.785 103.020 ;
        RECT 102.195 102.830 102.365 103.020 ;
        RECT 104.035 102.830 104.205 103.020 ;
        RECT 107.715 102.830 107.885 103.020 ;
        RECT 108.175 102.830 108.345 103.020 ;
        RECT 112.775 102.830 112.945 103.020 ;
        RECT 114.145 102.830 114.315 103.020 ;
        RECT 115.535 102.830 115.705 103.020 ;
      LAYER nwell ;
        RECT 20.485 54.580 29.875 66.420 ;
        RECT 31.685 54.590 41.075 66.430 ;
        RECT 42.905 54.560 52.295 66.400 ;
        RECT 54.155 54.540 63.545 66.380 ;
        RECT 65.375 54.530 74.765 66.370 ;
        RECT 76.615 54.520 86.005 66.360 ;
        RECT 87.865 54.530 97.255 66.370 ;
        RECT 99.145 54.520 108.535 66.360 ;
        RECT 110.415 54.520 119.805 66.360 ;
        RECT 121.665 54.520 131.055 66.360 ;
        RECT 132.415 54.490 139.375 66.330 ;
        RECT 20.655 49.020 23.115 53.210 ;
      LAYER pwell ;
        RECT 20.555 45.340 22.915 48.340 ;
      LAYER nwell ;
        RECT 24.735 45.940 29.125 53.130 ;
        RECT 31.855 49.030 34.315 53.220 ;
      LAYER pwell ;
        RECT 31.755 45.350 34.115 48.350 ;
      LAYER nwell ;
        RECT 35.935 45.950 40.325 53.140 ;
        RECT 43.075 49.000 45.535 53.190 ;
      LAYER pwell ;
        RECT 42.975 45.320 45.335 48.320 ;
      LAYER nwell ;
        RECT 47.155 45.920 51.545 53.110 ;
        RECT 54.325 48.980 56.785 53.170 ;
      LAYER pwell ;
        RECT 54.225 45.300 56.585 48.300 ;
      LAYER nwell ;
        RECT 58.405 45.900 62.795 53.090 ;
        RECT 65.545 48.970 68.005 53.160 ;
      LAYER pwell ;
        RECT 65.445 45.290 67.805 48.290 ;
      LAYER nwell ;
        RECT 69.625 45.890 74.015 53.080 ;
        RECT 76.785 48.960 79.245 53.150 ;
      LAYER pwell ;
        RECT 76.685 45.280 79.045 48.280 ;
      LAYER nwell ;
        RECT 80.865 45.880 85.255 53.070 ;
        RECT 88.035 48.970 90.495 53.160 ;
      LAYER pwell ;
        RECT 87.935 45.290 90.295 48.290 ;
      LAYER nwell ;
        RECT 92.115 45.890 96.505 53.080 ;
        RECT 99.315 48.960 101.775 53.150 ;
      LAYER pwell ;
        RECT 99.215 45.280 101.575 48.280 ;
      LAYER nwell ;
        RECT 103.395 45.880 107.785 53.070 ;
        RECT 110.585 48.960 113.045 53.150 ;
      LAYER pwell ;
        RECT 110.485 45.280 112.845 48.280 ;
      LAYER nwell ;
        RECT 114.665 45.880 119.055 53.070 ;
        RECT 121.835 48.960 124.295 53.150 ;
      LAYER pwell ;
        RECT 121.735 45.280 124.095 48.280 ;
      LAYER nwell ;
        RECT 125.915 45.880 130.305 53.070 ;
        RECT 19.615 32.280 24.005 39.470 ;
      LAYER pwell ;
        RECT 25.825 37.070 28.185 40.070 ;
      LAYER nwell ;
        RECT 25.625 32.200 28.085 36.390 ;
        RECT 30.895 32.280 35.285 39.470 ;
      LAYER pwell ;
        RECT 37.105 37.070 39.465 40.070 ;
      LAYER nwell ;
        RECT 36.905 32.200 39.365 36.390 ;
        RECT 42.185 32.260 46.575 39.450 ;
      LAYER pwell ;
        RECT 48.395 37.050 50.755 40.050 ;
      LAYER nwell ;
        RECT 48.195 32.180 50.655 36.370 ;
        RECT 53.405 32.260 57.795 39.450 ;
      LAYER pwell ;
        RECT 59.615 37.050 61.975 40.050 ;
      LAYER nwell ;
        RECT 59.415 32.180 61.875 36.370 ;
        RECT 64.605 32.260 68.995 39.450 ;
      LAYER pwell ;
        RECT 70.815 37.050 73.175 40.050 ;
      LAYER nwell ;
        RECT 70.615 32.180 73.075 36.370 ;
        RECT 75.895 32.250 80.285 39.440 ;
      LAYER pwell ;
        RECT 82.105 37.040 84.465 40.040 ;
      LAYER nwell ;
        RECT 81.905 32.170 84.365 36.360 ;
        RECT 87.135 32.270 91.525 39.460 ;
      LAYER pwell ;
        RECT 93.345 37.060 95.705 40.060 ;
      LAYER nwell ;
        RECT 93.145 32.190 95.605 36.380 ;
        RECT 98.345 32.290 102.735 39.480 ;
      LAYER pwell ;
        RECT 104.555 37.080 106.915 40.080 ;
      LAYER nwell ;
        RECT 104.355 32.210 106.815 36.400 ;
        RECT 109.545 32.330 113.935 39.520 ;
      LAYER pwell ;
        RECT 115.755 37.120 118.115 40.120 ;
      LAYER nwell ;
        RECT 115.555 32.250 118.015 36.440 ;
        RECT 120.755 32.350 125.145 39.540 ;
      LAYER pwell ;
        RECT 126.965 37.140 129.325 40.140 ;
      LAYER nwell ;
        RECT 126.765 32.270 129.225 36.460 ;
        RECT 18.865 18.990 28.255 30.830 ;
        RECT 30.145 18.990 39.535 30.830 ;
        RECT 41.435 18.970 50.825 30.810 ;
        RECT 52.655 18.970 62.045 30.810 ;
        RECT 63.855 18.970 73.245 30.810 ;
        RECT 75.145 18.960 84.535 30.800 ;
        RECT 86.385 18.980 95.775 30.820 ;
        RECT 97.595 19.000 106.985 30.840 ;
        RECT 108.795 19.040 118.185 30.880 ;
        RECT 120.005 19.060 129.395 30.900 ;
        RECT 131.725 19.030 138.685 30.870 ;
      LAYER li1 ;
        RECT 10.510 206.190 115.850 206.360 ;
        RECT 10.595 205.440 11.805 206.190 ;
        RECT 12.435 205.465 12.725 206.190 ;
        RECT 12.895 205.440 14.105 206.190 ;
        RECT 14.280 205.645 19.625 206.190 ;
        RECT 19.800 205.645 25.145 206.190 ;
        RECT 10.595 204.900 11.115 205.440 ;
        RECT 11.285 204.730 11.805 205.270 ;
        RECT 10.595 203.640 11.805 204.730 ;
        RECT 12.435 203.640 12.725 204.805 ;
        RECT 12.895 204.730 13.415 205.270 ;
        RECT 13.585 204.900 14.105 205.440 ;
        RECT 12.895 203.640 14.105 204.730 ;
        RECT 15.870 204.075 16.220 205.325 ;
        RECT 17.700 204.815 18.040 205.645 ;
        RECT 21.390 204.075 21.740 205.325 ;
        RECT 23.220 204.815 23.560 205.645 ;
        RECT 25.315 205.465 25.605 206.190 ;
        RECT 25.775 205.440 26.985 206.190 ;
        RECT 27.160 205.645 32.505 206.190 ;
        RECT 32.680 205.645 38.025 206.190 ;
        RECT 14.280 203.640 19.625 204.075 ;
        RECT 19.800 203.640 25.145 204.075 ;
        RECT 25.315 203.640 25.605 204.805 ;
        RECT 25.775 204.730 26.295 205.270 ;
        RECT 26.465 204.900 26.985 205.440 ;
        RECT 25.775 203.640 26.985 204.730 ;
        RECT 28.750 204.075 29.100 205.325 ;
        RECT 30.580 204.815 30.920 205.645 ;
        RECT 34.270 204.075 34.620 205.325 ;
        RECT 36.100 204.815 36.440 205.645 ;
        RECT 38.195 205.465 38.485 206.190 ;
        RECT 38.655 205.440 39.865 206.190 ;
        RECT 40.040 205.645 45.385 206.190 ;
        RECT 45.560 205.645 50.905 206.190 ;
        RECT 27.160 203.640 32.505 204.075 ;
        RECT 32.680 203.640 38.025 204.075 ;
        RECT 38.195 203.640 38.485 204.805 ;
        RECT 38.655 204.730 39.175 205.270 ;
        RECT 39.345 204.900 39.865 205.440 ;
        RECT 38.655 203.640 39.865 204.730 ;
        RECT 41.630 204.075 41.980 205.325 ;
        RECT 43.460 204.815 43.800 205.645 ;
        RECT 47.150 204.075 47.500 205.325 ;
        RECT 48.980 204.815 49.320 205.645 ;
        RECT 51.075 205.465 51.365 206.190 ;
        RECT 51.535 205.440 52.745 206.190 ;
        RECT 52.920 205.645 58.265 206.190 ;
        RECT 58.440 205.645 63.785 206.190 ;
        RECT 40.040 203.640 45.385 204.075 ;
        RECT 45.560 203.640 50.905 204.075 ;
        RECT 51.075 203.640 51.365 204.805 ;
        RECT 51.535 204.730 52.055 205.270 ;
        RECT 52.225 204.900 52.745 205.440 ;
        RECT 51.535 203.640 52.745 204.730 ;
        RECT 54.510 204.075 54.860 205.325 ;
        RECT 56.340 204.815 56.680 205.645 ;
        RECT 60.030 204.075 60.380 205.325 ;
        RECT 61.860 204.815 62.200 205.645 ;
        RECT 63.955 205.465 64.245 206.190 ;
        RECT 64.415 205.420 66.085 206.190 ;
        RECT 52.920 203.640 58.265 204.075 ;
        RECT 58.440 203.640 63.785 204.075 ;
        RECT 63.955 203.640 64.245 204.805 ;
        RECT 64.415 204.730 65.165 205.250 ;
        RECT 65.335 204.900 66.085 205.420 ;
        RECT 66.295 205.370 66.525 206.190 ;
        RECT 66.695 205.390 67.025 206.020 ;
        RECT 66.275 204.950 66.605 205.200 ;
        RECT 66.775 204.790 67.025 205.390 ;
        RECT 67.195 205.370 67.405 206.190 ;
        RECT 67.635 205.420 71.145 206.190 ;
        RECT 71.320 205.645 76.665 206.190 ;
        RECT 64.415 203.640 66.085 204.730 ;
        RECT 66.295 203.640 66.525 204.780 ;
        RECT 66.695 203.810 67.025 204.790 ;
        RECT 67.195 203.640 67.405 204.780 ;
        RECT 67.635 204.730 69.325 205.250 ;
        RECT 69.495 204.900 71.145 205.420 ;
        RECT 67.635 203.640 71.145 204.730 ;
        RECT 72.910 204.075 73.260 205.325 ;
        RECT 74.740 204.815 75.080 205.645 ;
        RECT 76.835 205.465 77.125 206.190 ;
        RECT 77.295 205.440 78.505 206.190 ;
        RECT 78.680 205.645 84.025 206.190 ;
        RECT 84.200 205.645 89.545 206.190 ;
        RECT 71.320 203.640 76.665 204.075 ;
        RECT 76.835 203.640 77.125 204.805 ;
        RECT 77.295 204.730 77.815 205.270 ;
        RECT 77.985 204.900 78.505 205.440 ;
        RECT 77.295 203.640 78.505 204.730 ;
        RECT 80.270 204.075 80.620 205.325 ;
        RECT 82.100 204.815 82.440 205.645 ;
        RECT 85.790 204.075 86.140 205.325 ;
        RECT 87.620 204.815 87.960 205.645 ;
        RECT 89.715 205.465 90.005 206.190 ;
        RECT 90.175 205.440 91.385 206.190 ;
        RECT 91.560 205.645 96.905 206.190 ;
        RECT 97.080 205.645 102.425 206.190 ;
        RECT 78.680 203.640 84.025 204.075 ;
        RECT 84.200 203.640 89.545 204.075 ;
        RECT 89.715 203.640 90.005 204.805 ;
        RECT 90.175 204.730 90.695 205.270 ;
        RECT 90.865 204.900 91.385 205.440 ;
        RECT 90.175 203.640 91.385 204.730 ;
        RECT 93.150 204.075 93.500 205.325 ;
        RECT 94.980 204.815 95.320 205.645 ;
        RECT 98.670 204.075 99.020 205.325 ;
        RECT 100.500 204.815 100.840 205.645 ;
        RECT 102.595 205.465 102.885 206.190 ;
        RECT 103.520 205.645 108.865 206.190 ;
        RECT 109.040 205.645 114.385 206.190 ;
        RECT 91.560 203.640 96.905 204.075 ;
        RECT 97.080 203.640 102.425 204.075 ;
        RECT 102.595 203.640 102.885 204.805 ;
        RECT 105.110 204.075 105.460 205.325 ;
        RECT 106.940 204.815 107.280 205.645 ;
        RECT 110.630 204.075 110.980 205.325 ;
        RECT 112.460 204.815 112.800 205.645 ;
        RECT 114.555 205.440 115.765 206.190 ;
        RECT 114.555 204.730 115.075 205.270 ;
        RECT 115.245 204.900 115.765 205.440 ;
        RECT 103.520 203.640 108.865 204.075 ;
        RECT 109.040 203.640 114.385 204.075 ;
        RECT 114.555 203.640 115.765 204.730 ;
        RECT 10.510 203.470 115.850 203.640 ;
        RECT 10.595 202.380 11.805 203.470 ;
        RECT 10.595 201.670 11.115 202.210 ;
        RECT 11.285 201.840 11.805 202.380 ;
        RECT 12.435 202.305 12.725 203.470 ;
        RECT 13.355 202.380 15.945 203.470 ;
        RECT 16.120 203.035 21.465 203.470 ;
        RECT 21.640 203.035 26.985 203.470 ;
        RECT 27.160 203.035 32.505 203.470 ;
        RECT 32.680 203.035 38.025 203.470 ;
        RECT 13.355 201.860 14.565 202.380 ;
        RECT 14.735 201.690 15.945 202.210 ;
        RECT 17.710 201.785 18.060 203.035 ;
        RECT 10.595 200.920 11.805 201.670 ;
        RECT 12.435 200.920 12.725 201.645 ;
        RECT 13.355 200.920 15.945 201.690 ;
        RECT 19.540 201.465 19.880 202.295 ;
        RECT 23.230 201.785 23.580 203.035 ;
        RECT 25.060 201.465 25.400 202.295 ;
        RECT 28.750 201.785 29.100 203.035 ;
        RECT 30.580 201.465 30.920 202.295 ;
        RECT 34.270 201.785 34.620 203.035 ;
        RECT 38.195 202.305 38.485 203.470 ;
        RECT 39.580 203.035 44.925 203.470 ;
        RECT 45.100 203.035 50.445 203.470 ;
        RECT 50.620 203.035 55.965 203.470 ;
        RECT 36.100 201.465 36.440 202.295 ;
        RECT 41.170 201.785 41.520 203.035 ;
        RECT 16.120 200.920 21.465 201.465 ;
        RECT 21.640 200.920 26.985 201.465 ;
        RECT 27.160 200.920 32.505 201.465 ;
        RECT 32.680 200.920 38.025 201.465 ;
        RECT 38.195 200.920 38.485 201.645 ;
        RECT 43.000 201.465 43.340 202.295 ;
        RECT 46.690 201.785 47.040 203.035 ;
        RECT 48.520 201.465 48.860 202.295 ;
        RECT 52.210 201.785 52.560 203.035 ;
        RECT 56.195 202.330 56.405 203.470 ;
        RECT 56.575 202.320 56.905 203.300 ;
        RECT 57.075 202.330 57.305 203.470 ;
        RECT 57.515 202.380 60.105 203.470 ;
        RECT 60.275 202.395 60.545 203.300 ;
        RECT 60.715 202.710 61.045 203.470 ;
        RECT 61.225 202.540 61.395 203.300 ;
        RECT 54.040 201.465 54.380 202.295 ;
        RECT 39.580 200.920 44.925 201.465 ;
        RECT 45.100 200.920 50.445 201.465 ;
        RECT 50.620 200.920 55.965 201.465 ;
        RECT 56.195 200.920 56.405 201.740 ;
        RECT 56.575 201.720 56.825 202.320 ;
        RECT 56.995 201.910 57.325 202.160 ;
        RECT 57.515 201.860 58.725 202.380 ;
        RECT 56.575 201.090 56.905 201.720 ;
        RECT 57.075 200.920 57.305 201.740 ;
        RECT 58.895 201.690 60.105 202.210 ;
        RECT 57.515 200.920 60.105 201.690 ;
        RECT 60.275 201.595 60.445 202.395 ;
        RECT 60.730 202.370 61.395 202.540 ;
        RECT 61.655 202.600 61.930 203.300 ;
        RECT 62.100 202.925 62.355 203.470 ;
        RECT 62.525 202.960 63.005 203.300 ;
        RECT 63.180 202.915 63.785 203.470 ;
        RECT 63.170 202.815 63.785 202.915 ;
        RECT 63.170 202.790 63.355 202.815 ;
        RECT 60.730 202.225 60.900 202.370 ;
        RECT 60.615 201.895 60.900 202.225 ;
        RECT 60.730 201.640 60.900 201.895 ;
        RECT 61.135 201.820 61.465 202.190 ;
        RECT 60.275 201.090 60.535 201.595 ;
        RECT 60.730 201.470 61.395 201.640 ;
        RECT 60.715 200.920 61.045 201.300 ;
        RECT 61.225 201.090 61.395 201.470 ;
        RECT 61.655 201.570 61.825 202.600 ;
        RECT 62.100 202.470 62.855 202.720 ;
        RECT 63.025 202.545 63.355 202.790 ;
        RECT 62.100 202.435 62.870 202.470 ;
        RECT 62.100 202.425 62.885 202.435 ;
        RECT 61.995 202.410 62.890 202.425 ;
        RECT 61.995 202.395 62.910 202.410 ;
        RECT 61.995 202.385 62.930 202.395 ;
        RECT 61.995 202.375 62.955 202.385 ;
        RECT 61.995 202.345 63.025 202.375 ;
        RECT 61.995 202.315 63.045 202.345 ;
        RECT 61.995 202.285 63.065 202.315 ;
        RECT 61.995 202.260 63.095 202.285 ;
        RECT 61.995 202.225 63.130 202.260 ;
        RECT 61.995 202.220 63.160 202.225 ;
        RECT 61.995 201.825 62.225 202.220 ;
        RECT 62.770 202.215 63.160 202.220 ;
        RECT 62.795 202.205 63.160 202.215 ;
        RECT 62.810 202.200 63.160 202.205 ;
        RECT 62.825 202.195 63.160 202.200 ;
        RECT 63.525 202.195 63.785 202.645 ;
        RECT 63.955 202.305 64.245 203.470 ;
        RECT 62.825 202.190 63.785 202.195 ;
        RECT 62.835 202.180 63.785 202.190 ;
        RECT 62.845 202.175 63.785 202.180 ;
        RECT 62.855 202.165 63.785 202.175 ;
        RECT 62.860 202.155 63.785 202.165 ;
        RECT 62.865 202.150 63.785 202.155 ;
        RECT 62.875 202.135 63.785 202.150 ;
        RECT 62.880 202.120 63.785 202.135 ;
        RECT 62.890 202.095 63.785 202.120 ;
        RECT 62.395 201.625 62.725 202.050 ;
        RECT 61.655 201.090 61.915 201.570 ;
        RECT 62.085 200.920 62.335 201.460 ;
        RECT 62.505 201.140 62.725 201.625 ;
        RECT 62.895 202.025 63.785 202.095 ;
        RECT 64.420 202.280 64.675 203.160 ;
        RECT 64.845 202.330 65.150 203.470 ;
        RECT 65.490 203.090 65.820 203.470 ;
        RECT 66.000 202.920 66.170 203.210 ;
        RECT 66.340 203.010 66.590 203.470 ;
        RECT 65.370 202.750 66.170 202.920 ;
        RECT 66.760 202.960 67.630 203.300 ;
        RECT 62.895 201.300 63.065 202.025 ;
        RECT 63.235 201.470 63.785 201.855 ;
        RECT 62.895 201.130 63.785 201.300 ;
        RECT 63.955 200.920 64.245 201.645 ;
        RECT 64.420 201.630 64.630 202.280 ;
        RECT 65.370 202.160 65.540 202.750 ;
        RECT 66.760 202.580 66.930 202.960 ;
        RECT 67.865 202.840 68.035 203.300 ;
        RECT 68.205 203.010 68.575 203.470 ;
        RECT 68.870 202.870 69.040 203.210 ;
        RECT 69.210 203.040 69.540 203.470 ;
        RECT 69.775 202.870 69.945 203.210 ;
        RECT 65.710 202.410 66.930 202.580 ;
        RECT 67.100 202.500 67.560 202.790 ;
        RECT 67.865 202.670 68.425 202.840 ;
        RECT 68.870 202.700 69.945 202.870 ;
        RECT 70.115 202.970 70.795 203.300 ;
        RECT 71.010 202.970 71.260 203.300 ;
        RECT 71.430 203.010 71.680 203.470 ;
        RECT 68.255 202.530 68.425 202.670 ;
        RECT 67.100 202.490 68.065 202.500 ;
        RECT 66.760 202.320 66.930 202.410 ;
        RECT 67.390 202.330 68.065 202.490 ;
        RECT 64.800 202.130 65.540 202.160 ;
        RECT 64.800 201.830 65.715 202.130 ;
        RECT 65.390 201.655 65.715 201.830 ;
        RECT 64.420 201.100 64.675 201.630 ;
        RECT 64.845 200.920 65.150 201.380 ;
        RECT 65.395 201.300 65.715 201.655 ;
        RECT 65.885 201.870 66.425 202.240 ;
        RECT 66.760 202.150 67.165 202.320 ;
        RECT 65.885 201.470 66.125 201.870 ;
        RECT 66.605 201.700 66.825 201.980 ;
        RECT 66.295 201.530 66.825 201.700 ;
        RECT 66.295 201.300 66.465 201.530 ;
        RECT 66.995 201.370 67.165 202.150 ;
        RECT 67.335 201.540 67.685 202.160 ;
        RECT 67.855 201.540 68.065 202.330 ;
        RECT 68.255 202.360 69.755 202.530 ;
        RECT 68.255 201.670 68.425 202.360 ;
        RECT 70.115 202.190 70.285 202.970 ;
        RECT 71.090 202.840 71.260 202.970 ;
        RECT 68.595 202.020 70.285 202.190 ;
        RECT 70.455 202.410 70.920 202.800 ;
        RECT 71.090 202.670 71.485 202.840 ;
        RECT 68.595 201.840 68.765 202.020 ;
        RECT 65.395 201.130 66.465 201.300 ;
        RECT 66.635 200.920 66.825 201.360 ;
        RECT 66.995 201.090 67.945 201.370 ;
        RECT 68.255 201.280 68.515 201.670 ;
        RECT 68.935 201.600 69.725 201.850 ;
        RECT 68.165 201.110 68.515 201.280 ;
        RECT 68.725 200.920 69.055 201.380 ;
        RECT 69.930 201.310 70.100 202.020 ;
        RECT 70.455 201.820 70.625 202.410 ;
        RECT 70.270 201.600 70.625 201.820 ;
        RECT 70.795 201.600 71.145 202.220 ;
        RECT 71.315 201.310 71.485 202.670 ;
        RECT 71.850 202.500 72.175 203.285 ;
        RECT 71.655 201.450 72.115 202.500 ;
        RECT 69.930 201.140 70.785 201.310 ;
        RECT 70.990 201.140 71.485 201.310 ;
        RECT 71.655 200.920 71.985 201.280 ;
        RECT 72.345 201.180 72.515 203.300 ;
        RECT 72.685 202.970 73.015 203.470 ;
        RECT 73.185 202.800 73.440 203.300 ;
        RECT 72.690 202.630 73.440 202.800 ;
        RECT 72.690 201.640 72.920 202.630 ;
        RECT 73.090 201.810 73.440 202.460 ;
        RECT 74.075 202.380 75.745 203.470 ;
        RECT 75.915 202.395 76.185 203.300 ;
        RECT 76.355 202.710 76.685 203.470 ;
        RECT 76.865 202.540 77.035 203.300 ;
        RECT 74.075 201.860 74.825 202.380 ;
        RECT 74.995 201.690 75.745 202.210 ;
        RECT 72.690 201.470 73.440 201.640 ;
        RECT 72.685 200.920 73.015 201.300 ;
        RECT 73.185 201.180 73.440 201.470 ;
        RECT 74.075 200.920 75.745 201.690 ;
        RECT 75.915 201.595 76.085 202.395 ;
        RECT 76.370 202.370 77.035 202.540 ;
        RECT 77.295 202.380 78.505 203.470 ;
        RECT 78.680 203.035 84.025 203.470 ;
        RECT 84.200 203.035 89.545 203.470 ;
        RECT 76.370 202.225 76.540 202.370 ;
        RECT 76.255 201.895 76.540 202.225 ;
        RECT 76.370 201.640 76.540 201.895 ;
        RECT 76.775 201.820 77.105 202.190 ;
        RECT 77.295 201.840 77.815 202.380 ;
        RECT 77.985 201.670 78.505 202.210 ;
        RECT 80.270 201.785 80.620 203.035 ;
        RECT 75.915 201.090 76.175 201.595 ;
        RECT 76.370 201.470 77.035 201.640 ;
        RECT 76.355 200.920 76.685 201.300 ;
        RECT 76.865 201.090 77.035 201.470 ;
        RECT 77.295 200.920 78.505 201.670 ;
        RECT 82.100 201.465 82.440 202.295 ;
        RECT 85.790 201.785 86.140 203.035 ;
        RECT 89.715 202.305 90.005 203.470 ;
        RECT 90.635 202.380 92.305 203.470 ;
        RECT 92.480 203.035 97.825 203.470 ;
        RECT 98.000 203.035 103.345 203.470 ;
        RECT 103.520 203.035 108.865 203.470 ;
        RECT 109.040 203.035 114.385 203.470 ;
        RECT 87.620 201.465 87.960 202.295 ;
        RECT 90.635 201.860 91.385 202.380 ;
        RECT 91.555 201.690 92.305 202.210 ;
        RECT 94.070 201.785 94.420 203.035 ;
        RECT 78.680 200.920 84.025 201.465 ;
        RECT 84.200 200.920 89.545 201.465 ;
        RECT 89.715 200.920 90.005 201.645 ;
        RECT 90.635 200.920 92.305 201.690 ;
        RECT 95.900 201.465 96.240 202.295 ;
        RECT 99.590 201.785 99.940 203.035 ;
        RECT 101.420 201.465 101.760 202.295 ;
        RECT 105.110 201.785 105.460 203.035 ;
        RECT 106.940 201.465 107.280 202.295 ;
        RECT 110.630 201.785 110.980 203.035 ;
        RECT 114.555 202.380 115.765 203.470 ;
        RECT 112.460 201.465 112.800 202.295 ;
        RECT 114.555 201.840 115.075 202.380 ;
        RECT 115.245 201.670 115.765 202.210 ;
        RECT 92.480 200.920 97.825 201.465 ;
        RECT 98.000 200.920 103.345 201.465 ;
        RECT 103.520 200.920 108.865 201.465 ;
        RECT 109.040 200.920 114.385 201.465 ;
        RECT 114.555 200.920 115.765 201.670 ;
        RECT 10.510 200.750 115.850 200.920 ;
        RECT 10.595 200.000 11.805 200.750 ;
        RECT 10.595 199.460 11.115 200.000 ;
        RECT 12.435 199.980 14.105 200.750 ;
        RECT 14.280 200.205 19.625 200.750 ;
        RECT 19.800 200.205 25.145 200.750 ;
        RECT 11.285 199.290 11.805 199.830 ;
        RECT 10.595 198.200 11.805 199.290 ;
        RECT 12.435 199.290 13.185 199.810 ;
        RECT 13.355 199.460 14.105 199.980 ;
        RECT 12.435 198.200 14.105 199.290 ;
        RECT 15.870 198.635 16.220 199.885 ;
        RECT 17.700 199.375 18.040 200.205 ;
        RECT 21.390 198.635 21.740 199.885 ;
        RECT 23.220 199.375 23.560 200.205 ;
        RECT 25.315 200.025 25.605 200.750 ;
        RECT 26.235 199.980 28.825 200.750 ;
        RECT 29.000 200.205 34.345 200.750 ;
        RECT 34.520 200.205 39.865 200.750 ;
        RECT 40.040 200.205 45.385 200.750 ;
        RECT 45.560 200.205 50.905 200.750 ;
        RECT 14.280 198.200 19.625 198.635 ;
        RECT 19.800 198.200 25.145 198.635 ;
        RECT 25.315 198.200 25.605 199.365 ;
        RECT 26.235 199.290 27.445 199.810 ;
        RECT 27.615 199.460 28.825 199.980 ;
        RECT 26.235 198.200 28.825 199.290 ;
        RECT 30.590 198.635 30.940 199.885 ;
        RECT 32.420 199.375 32.760 200.205 ;
        RECT 36.110 198.635 36.460 199.885 ;
        RECT 37.940 199.375 38.280 200.205 ;
        RECT 41.630 198.635 41.980 199.885 ;
        RECT 43.460 199.375 43.800 200.205 ;
        RECT 47.150 198.635 47.500 199.885 ;
        RECT 48.980 199.375 49.320 200.205 ;
        RECT 51.075 200.025 51.365 200.750 ;
        RECT 51.845 200.280 52.015 200.750 ;
        RECT 52.185 200.100 52.515 200.580 ;
        RECT 52.685 200.280 52.855 200.750 ;
        RECT 53.025 200.100 53.355 200.580 ;
        RECT 51.590 199.930 53.355 200.100 ;
        RECT 53.525 199.940 53.695 200.750 ;
        RECT 53.895 200.370 54.965 200.540 ;
        RECT 53.895 200.015 54.215 200.370 ;
        RECT 51.590 199.380 52.000 199.930 ;
        RECT 53.890 199.760 54.215 200.015 ;
        RECT 52.185 199.550 54.215 199.760 ;
        RECT 53.870 199.540 54.215 199.550 ;
        RECT 54.385 199.800 54.625 200.200 ;
        RECT 54.795 200.140 54.965 200.370 ;
        RECT 55.135 200.310 55.325 200.750 ;
        RECT 55.495 200.300 56.445 200.580 ;
        RECT 56.665 200.390 57.015 200.560 ;
        RECT 54.795 199.970 55.325 200.140 ;
        RECT 29.000 198.200 34.345 198.635 ;
        RECT 34.520 198.200 39.865 198.635 ;
        RECT 40.040 198.200 45.385 198.635 ;
        RECT 45.560 198.200 50.905 198.635 ;
        RECT 51.075 198.200 51.365 199.365 ;
        RECT 51.590 199.210 53.315 199.380 ;
        RECT 51.845 198.200 52.015 199.040 ;
        RECT 52.225 198.370 52.475 199.210 ;
        RECT 52.685 198.200 52.855 199.040 ;
        RECT 53.025 198.370 53.315 199.210 ;
        RECT 53.525 198.200 53.695 199.260 ;
        RECT 53.870 198.920 54.040 199.540 ;
        RECT 54.385 199.430 54.925 199.800 ;
        RECT 55.105 199.690 55.325 199.970 ;
        RECT 55.495 199.520 55.665 200.300 ;
        RECT 55.260 199.350 55.665 199.520 ;
        RECT 55.835 199.510 56.185 200.130 ;
        RECT 55.260 199.260 55.430 199.350 ;
        RECT 56.355 199.340 56.565 200.130 ;
        RECT 54.210 199.090 55.430 199.260 ;
        RECT 55.890 199.180 56.565 199.340 ;
        RECT 53.870 198.750 54.670 198.920 ;
        RECT 53.990 198.200 54.320 198.580 ;
        RECT 54.500 198.460 54.670 198.750 ;
        RECT 55.260 198.710 55.430 199.090 ;
        RECT 55.600 199.170 56.565 199.180 ;
        RECT 56.755 200.000 57.015 200.390 ;
        RECT 57.225 200.290 57.555 200.750 ;
        RECT 58.430 200.360 59.285 200.530 ;
        RECT 59.490 200.360 59.985 200.530 ;
        RECT 60.155 200.390 60.485 200.750 ;
        RECT 56.755 199.310 56.925 200.000 ;
        RECT 57.095 199.650 57.265 199.830 ;
        RECT 57.435 199.820 58.225 200.070 ;
        RECT 58.430 199.650 58.600 200.360 ;
        RECT 58.770 199.850 59.125 200.070 ;
        RECT 57.095 199.480 58.785 199.650 ;
        RECT 55.600 198.880 56.060 199.170 ;
        RECT 56.755 199.140 58.255 199.310 ;
        RECT 56.755 199.000 56.925 199.140 ;
        RECT 56.365 198.830 56.925 199.000 ;
        RECT 54.840 198.200 55.090 198.660 ;
        RECT 55.260 198.370 56.130 198.710 ;
        RECT 56.365 198.370 56.535 198.830 ;
        RECT 57.370 198.800 58.445 198.970 ;
        RECT 56.705 198.200 57.075 198.660 ;
        RECT 57.370 198.460 57.540 198.800 ;
        RECT 57.710 198.200 58.040 198.630 ;
        RECT 58.275 198.460 58.445 198.800 ;
        RECT 58.615 198.700 58.785 199.480 ;
        RECT 58.955 199.260 59.125 199.850 ;
        RECT 59.295 199.450 59.645 200.070 ;
        RECT 58.955 198.870 59.420 199.260 ;
        RECT 59.815 199.000 59.985 200.360 ;
        RECT 60.155 199.170 60.615 200.220 ;
        RECT 59.590 198.830 59.985 199.000 ;
        RECT 59.590 198.700 59.760 198.830 ;
        RECT 58.615 198.370 59.295 198.700 ;
        RECT 59.510 198.370 59.760 198.700 ;
        RECT 59.930 198.200 60.180 198.660 ;
        RECT 60.350 198.385 60.675 199.170 ;
        RECT 60.845 198.370 61.015 200.490 ;
        RECT 61.185 200.370 61.515 200.750 ;
        RECT 61.685 200.200 61.940 200.490 ;
        RECT 61.190 200.030 61.940 200.200 ;
        RECT 61.190 199.040 61.420 200.030 ;
        RECT 62.575 199.930 62.835 200.750 ;
        RECT 63.005 199.930 63.335 200.350 ;
        RECT 63.515 200.180 63.775 200.580 ;
        RECT 63.945 200.350 64.275 200.750 ;
        RECT 64.445 200.180 64.615 200.530 ;
        RECT 64.785 200.350 65.160 200.750 ;
        RECT 63.515 200.010 65.180 200.180 ;
        RECT 65.350 200.075 65.625 200.420 ;
        RECT 61.590 199.210 61.940 199.860 ;
        RECT 63.085 199.840 63.335 199.930 ;
        RECT 65.010 199.840 65.180 200.010 ;
        RECT 62.580 199.510 62.915 199.760 ;
        RECT 63.085 199.510 63.800 199.840 ;
        RECT 64.015 199.510 64.840 199.840 ;
        RECT 65.010 199.510 65.285 199.840 ;
        RECT 61.190 198.870 61.940 199.040 ;
        RECT 61.185 198.200 61.515 198.700 ;
        RECT 61.685 198.370 61.940 198.870 ;
        RECT 62.575 198.200 62.835 199.340 ;
        RECT 63.085 198.950 63.255 199.510 ;
        RECT 63.515 199.050 63.845 199.340 ;
        RECT 64.015 199.220 64.260 199.510 ;
        RECT 65.010 199.340 65.180 199.510 ;
        RECT 65.455 199.340 65.625 200.075 ;
        RECT 65.885 200.200 66.055 200.580 ;
        RECT 66.270 200.370 66.600 200.750 ;
        RECT 65.885 200.030 66.600 200.200 ;
        RECT 65.795 199.480 66.150 199.850 ;
        RECT 66.430 199.840 66.600 200.030 ;
        RECT 66.770 200.005 67.025 200.580 ;
        RECT 66.430 199.510 66.685 199.840 ;
        RECT 64.520 199.170 65.180 199.340 ;
        RECT 64.520 199.050 64.690 199.170 ;
        RECT 63.515 198.880 64.690 199.050 ;
        RECT 63.075 198.380 64.690 198.710 ;
        RECT 64.860 198.200 65.140 199.000 ;
        RECT 65.350 198.370 65.625 199.340 ;
        RECT 66.430 199.300 66.600 199.510 ;
        RECT 65.885 199.130 66.600 199.300 ;
        RECT 66.855 199.275 67.025 200.005 ;
        RECT 67.200 199.910 67.460 200.750 ;
        RECT 67.640 200.040 67.895 200.570 ;
        RECT 68.065 200.290 68.370 200.750 ;
        RECT 68.615 200.370 69.685 200.540 ;
        RECT 67.640 199.390 67.850 200.040 ;
        RECT 68.615 200.015 68.935 200.370 ;
        RECT 68.610 199.840 68.935 200.015 ;
        RECT 68.020 199.540 68.935 199.840 ;
        RECT 69.105 199.800 69.345 200.200 ;
        RECT 69.515 200.140 69.685 200.370 ;
        RECT 69.855 200.310 70.045 200.750 ;
        RECT 70.215 200.300 71.165 200.580 ;
        RECT 71.385 200.390 71.735 200.560 ;
        RECT 69.515 199.970 70.045 200.140 ;
        RECT 68.020 199.510 68.760 199.540 ;
        RECT 65.885 198.370 66.055 199.130 ;
        RECT 66.270 198.200 66.600 198.960 ;
        RECT 66.770 198.370 67.025 199.275 ;
        RECT 67.200 198.200 67.460 199.350 ;
        RECT 67.640 198.510 67.895 199.390 ;
        RECT 68.065 198.200 68.370 199.340 ;
        RECT 68.590 198.920 68.760 199.510 ;
        RECT 69.105 199.430 69.645 199.800 ;
        RECT 69.825 199.690 70.045 199.970 ;
        RECT 70.215 199.520 70.385 200.300 ;
        RECT 69.980 199.350 70.385 199.520 ;
        RECT 70.555 199.510 70.905 200.130 ;
        RECT 69.980 199.260 70.150 199.350 ;
        RECT 71.075 199.340 71.285 200.130 ;
        RECT 68.930 199.090 70.150 199.260 ;
        RECT 70.610 199.180 71.285 199.340 ;
        RECT 68.590 198.750 69.390 198.920 ;
        RECT 68.710 198.200 69.040 198.580 ;
        RECT 69.220 198.460 69.390 198.750 ;
        RECT 69.980 198.710 70.150 199.090 ;
        RECT 70.320 199.170 71.285 199.180 ;
        RECT 71.475 200.000 71.735 200.390 ;
        RECT 71.945 200.290 72.275 200.750 ;
        RECT 73.150 200.360 74.005 200.530 ;
        RECT 74.210 200.360 74.705 200.530 ;
        RECT 74.875 200.390 75.205 200.750 ;
        RECT 71.475 199.310 71.645 200.000 ;
        RECT 71.815 199.650 71.985 199.830 ;
        RECT 72.155 199.820 72.945 200.070 ;
        RECT 73.150 199.650 73.320 200.360 ;
        RECT 73.490 199.850 73.845 200.070 ;
        RECT 71.815 199.480 73.505 199.650 ;
        RECT 70.320 198.880 70.780 199.170 ;
        RECT 71.475 199.140 72.975 199.310 ;
        RECT 71.475 199.000 71.645 199.140 ;
        RECT 71.085 198.830 71.645 199.000 ;
        RECT 69.560 198.200 69.810 198.660 ;
        RECT 69.980 198.370 70.850 198.710 ;
        RECT 71.085 198.370 71.255 198.830 ;
        RECT 72.090 198.800 73.165 198.970 ;
        RECT 71.425 198.200 71.795 198.660 ;
        RECT 72.090 198.460 72.260 198.800 ;
        RECT 72.430 198.200 72.760 198.630 ;
        RECT 72.995 198.460 73.165 198.800 ;
        RECT 73.335 198.700 73.505 199.480 ;
        RECT 73.675 199.260 73.845 199.850 ;
        RECT 74.015 199.450 74.365 200.070 ;
        RECT 73.675 198.870 74.140 199.260 ;
        RECT 74.535 199.000 74.705 200.360 ;
        RECT 74.875 199.170 75.335 200.220 ;
        RECT 74.310 198.830 74.705 199.000 ;
        RECT 74.310 198.700 74.480 198.830 ;
        RECT 73.335 198.370 74.015 198.700 ;
        RECT 74.230 198.370 74.480 198.700 ;
        RECT 74.650 198.200 74.900 198.660 ;
        RECT 75.070 198.385 75.395 199.170 ;
        RECT 75.565 198.370 75.735 200.490 ;
        RECT 75.905 200.370 76.235 200.750 ;
        RECT 76.405 200.200 76.660 200.490 ;
        RECT 75.910 200.030 76.660 200.200 ;
        RECT 75.910 199.040 76.140 200.030 ;
        RECT 76.835 200.025 77.125 200.750 ;
        RECT 77.355 199.930 77.565 200.750 ;
        RECT 77.735 199.950 78.065 200.580 ;
        RECT 76.310 199.210 76.660 199.860 ;
        RECT 75.910 198.870 76.660 199.040 ;
        RECT 75.905 198.200 76.235 198.700 ;
        RECT 76.405 198.370 76.660 198.870 ;
        RECT 76.835 198.200 77.125 199.365 ;
        RECT 77.735 199.350 77.985 199.950 ;
        RECT 78.235 199.930 78.465 200.750 ;
        RECT 78.675 199.980 80.345 200.750 ;
        RECT 80.520 200.205 85.865 200.750 ;
        RECT 86.040 200.205 91.385 200.750 ;
        RECT 91.560 200.205 96.905 200.750 ;
        RECT 97.080 200.205 102.425 200.750 ;
        RECT 78.155 199.510 78.485 199.760 ;
        RECT 77.355 198.200 77.565 199.340 ;
        RECT 77.735 198.370 78.065 199.350 ;
        RECT 78.235 198.200 78.465 199.340 ;
        RECT 78.675 199.290 79.425 199.810 ;
        RECT 79.595 199.460 80.345 199.980 ;
        RECT 78.675 198.200 80.345 199.290 ;
        RECT 82.110 198.635 82.460 199.885 ;
        RECT 83.940 199.375 84.280 200.205 ;
        RECT 87.630 198.635 87.980 199.885 ;
        RECT 89.460 199.375 89.800 200.205 ;
        RECT 93.150 198.635 93.500 199.885 ;
        RECT 94.980 199.375 95.320 200.205 ;
        RECT 98.670 198.635 99.020 199.885 ;
        RECT 100.500 199.375 100.840 200.205 ;
        RECT 102.595 200.025 102.885 200.750 ;
        RECT 103.520 200.205 108.865 200.750 ;
        RECT 109.040 200.205 114.385 200.750 ;
        RECT 80.520 198.200 85.865 198.635 ;
        RECT 86.040 198.200 91.385 198.635 ;
        RECT 91.560 198.200 96.905 198.635 ;
        RECT 97.080 198.200 102.425 198.635 ;
        RECT 102.595 198.200 102.885 199.365 ;
        RECT 105.110 198.635 105.460 199.885 ;
        RECT 106.940 199.375 107.280 200.205 ;
        RECT 110.630 198.635 110.980 199.885 ;
        RECT 112.460 199.375 112.800 200.205 ;
        RECT 114.555 200.000 115.765 200.750 ;
        RECT 114.555 199.290 115.075 199.830 ;
        RECT 115.245 199.460 115.765 200.000 ;
        RECT 103.520 198.200 108.865 198.635 ;
        RECT 109.040 198.200 114.385 198.635 ;
        RECT 114.555 198.200 115.765 199.290 ;
        RECT 10.510 198.030 115.850 198.200 ;
        RECT 10.595 196.940 11.805 198.030 ;
        RECT 10.595 196.230 11.115 196.770 ;
        RECT 11.285 196.400 11.805 196.940 ;
        RECT 12.435 196.865 12.725 198.030 ;
        RECT 13.355 196.940 15.945 198.030 ;
        RECT 16.120 197.595 21.465 198.030 ;
        RECT 21.640 197.595 26.985 198.030 ;
        RECT 27.160 197.595 32.505 198.030 ;
        RECT 32.680 197.595 38.025 198.030 ;
        RECT 13.355 196.420 14.565 196.940 ;
        RECT 14.735 196.250 15.945 196.770 ;
        RECT 17.710 196.345 18.060 197.595 ;
        RECT 10.595 195.480 11.805 196.230 ;
        RECT 12.435 195.480 12.725 196.205 ;
        RECT 13.355 195.480 15.945 196.250 ;
        RECT 19.540 196.025 19.880 196.855 ;
        RECT 23.230 196.345 23.580 197.595 ;
        RECT 25.060 196.025 25.400 196.855 ;
        RECT 28.750 196.345 29.100 197.595 ;
        RECT 30.580 196.025 30.920 196.855 ;
        RECT 34.270 196.345 34.620 197.595 ;
        RECT 38.195 196.865 38.485 198.030 ;
        RECT 38.660 197.595 44.005 198.030 ;
        RECT 44.180 197.595 49.525 198.030 ;
        RECT 36.100 196.025 36.440 196.855 ;
        RECT 40.250 196.345 40.600 197.595 ;
        RECT 16.120 195.480 21.465 196.025 ;
        RECT 21.640 195.480 26.985 196.025 ;
        RECT 27.160 195.480 32.505 196.025 ;
        RECT 32.680 195.480 38.025 196.025 ;
        RECT 38.195 195.480 38.485 196.205 ;
        RECT 42.080 196.025 42.420 196.855 ;
        RECT 45.770 196.345 46.120 197.595 ;
        RECT 49.700 197.360 49.955 197.860 ;
        RECT 50.125 197.530 50.455 198.030 ;
        RECT 49.700 197.190 50.450 197.360 ;
        RECT 47.600 196.025 47.940 196.855 ;
        RECT 49.700 196.370 50.050 197.020 ;
        RECT 50.220 196.200 50.450 197.190 ;
        RECT 49.700 196.030 50.450 196.200 ;
        RECT 38.660 195.480 44.005 196.025 ;
        RECT 44.180 195.480 49.525 196.025 ;
        RECT 49.700 195.740 49.955 196.030 ;
        RECT 50.125 195.480 50.455 195.860 ;
        RECT 50.625 195.740 50.795 197.860 ;
        RECT 50.965 197.060 51.290 197.845 ;
        RECT 51.460 197.570 51.710 198.030 ;
        RECT 51.880 197.530 52.130 197.860 ;
        RECT 52.345 197.530 53.025 197.860 ;
        RECT 51.880 197.400 52.050 197.530 ;
        RECT 51.655 197.230 52.050 197.400 ;
        RECT 51.025 196.010 51.485 197.060 ;
        RECT 51.655 195.870 51.825 197.230 ;
        RECT 52.220 196.970 52.685 197.360 ;
        RECT 51.995 196.160 52.345 196.780 ;
        RECT 52.515 196.380 52.685 196.970 ;
        RECT 52.855 196.750 53.025 197.530 ;
        RECT 53.195 197.430 53.365 197.770 ;
        RECT 53.600 197.600 53.930 198.030 ;
        RECT 54.100 197.430 54.270 197.770 ;
        RECT 54.565 197.570 54.935 198.030 ;
        RECT 53.195 197.260 54.270 197.430 ;
        RECT 55.105 197.400 55.275 197.860 ;
        RECT 55.510 197.520 56.380 197.860 ;
        RECT 56.550 197.570 56.800 198.030 ;
        RECT 54.715 197.230 55.275 197.400 ;
        RECT 54.715 197.090 54.885 197.230 ;
        RECT 53.385 196.920 54.885 197.090 ;
        RECT 55.580 197.060 56.040 197.350 ;
        RECT 52.855 196.580 54.545 196.750 ;
        RECT 52.515 196.160 52.870 196.380 ;
        RECT 53.040 195.870 53.210 196.580 ;
        RECT 53.415 196.160 54.205 196.410 ;
        RECT 54.375 196.400 54.545 196.580 ;
        RECT 54.715 196.230 54.885 196.920 ;
        RECT 51.155 195.480 51.485 195.840 ;
        RECT 51.655 195.700 52.150 195.870 ;
        RECT 52.355 195.700 53.210 195.870 ;
        RECT 54.085 195.480 54.415 195.940 ;
        RECT 54.625 195.840 54.885 196.230 ;
        RECT 55.075 197.050 56.040 197.060 ;
        RECT 56.210 197.140 56.380 197.520 ;
        RECT 56.970 197.480 57.140 197.770 ;
        RECT 57.320 197.650 57.650 198.030 ;
        RECT 56.970 197.310 57.770 197.480 ;
        RECT 55.075 196.890 55.750 197.050 ;
        RECT 56.210 196.970 57.430 197.140 ;
        RECT 55.075 196.100 55.285 196.890 ;
        RECT 56.210 196.880 56.380 196.970 ;
        RECT 55.455 196.100 55.805 196.720 ;
        RECT 55.975 196.710 56.380 196.880 ;
        RECT 55.975 195.930 56.145 196.710 ;
        RECT 56.315 196.260 56.535 196.540 ;
        RECT 56.715 196.430 57.255 196.800 ;
        RECT 57.600 196.720 57.770 197.310 ;
        RECT 57.990 196.890 58.295 198.030 ;
        RECT 58.465 196.840 58.715 197.720 ;
        RECT 58.885 196.890 59.135 198.030 ;
        RECT 59.375 197.520 59.675 198.030 ;
        RECT 59.845 197.520 60.225 197.690 ;
        RECT 60.805 197.520 61.435 198.030 ;
        RECT 59.845 197.350 60.015 197.520 ;
        RECT 61.605 197.350 61.935 197.860 ;
        RECT 62.105 197.520 62.405 198.030 ;
        RECT 59.355 197.150 60.015 197.350 ;
        RECT 60.185 197.180 62.405 197.350 ;
        RECT 57.600 196.690 58.340 196.720 ;
        RECT 56.315 196.090 56.845 196.260 ;
        RECT 54.625 195.670 54.975 195.840 ;
        RECT 55.195 195.650 56.145 195.930 ;
        RECT 56.315 195.480 56.505 195.920 ;
        RECT 56.675 195.860 56.845 196.090 ;
        RECT 57.015 196.030 57.255 196.430 ;
        RECT 57.425 196.390 58.340 196.690 ;
        RECT 57.425 196.215 57.750 196.390 ;
        RECT 57.425 195.860 57.745 196.215 ;
        RECT 58.510 196.190 58.715 196.840 ;
        RECT 56.675 195.690 57.745 195.860 ;
        RECT 57.990 195.480 58.295 195.940 ;
        RECT 58.465 195.660 58.715 196.190 ;
        RECT 58.885 195.480 59.135 196.235 ;
        RECT 59.355 196.220 59.525 197.150 ;
        RECT 60.185 196.980 60.355 197.180 ;
        RECT 59.695 196.810 60.355 196.980 ;
        RECT 60.525 196.840 62.065 197.010 ;
        RECT 59.695 196.390 59.865 196.810 ;
        RECT 60.525 196.640 60.695 196.840 ;
        RECT 60.095 196.470 60.695 196.640 ;
        RECT 60.865 196.470 61.560 196.670 ;
        RECT 61.820 196.390 62.065 196.840 ;
        RECT 60.185 196.220 61.095 196.300 ;
        RECT 59.355 195.740 59.675 196.220 ;
        RECT 59.845 196.130 61.095 196.220 ;
        RECT 59.845 196.050 60.355 196.130 ;
        RECT 59.845 195.650 60.075 196.050 ;
        RECT 60.245 195.480 60.595 195.870 ;
        RECT 60.765 195.650 61.095 196.130 ;
        RECT 61.265 195.480 61.435 196.300 ;
        RECT 62.235 196.220 62.405 197.180 ;
        RECT 62.575 196.890 62.855 198.030 ;
        RECT 63.025 196.880 63.355 197.860 ;
        RECT 63.525 196.890 63.785 198.030 ;
        RECT 62.585 196.450 62.920 196.720 ;
        RECT 63.090 196.280 63.260 196.880 ;
        RECT 63.955 196.865 64.245 198.030 ;
        RECT 64.425 196.970 64.755 197.820 ;
        RECT 63.430 196.470 63.765 196.720 ;
        RECT 61.940 195.675 62.405 196.220 ;
        RECT 62.575 195.480 62.885 196.280 ;
        RECT 63.090 195.650 63.785 196.280 ;
        RECT 64.425 196.205 64.615 196.970 ;
        RECT 64.925 196.890 65.175 198.030 ;
        RECT 65.365 197.390 65.615 197.810 ;
        RECT 65.845 197.560 66.175 198.030 ;
        RECT 66.405 197.390 66.655 197.810 ;
        RECT 65.365 197.220 66.655 197.390 ;
        RECT 66.835 197.390 67.165 197.820 ;
        RECT 68.555 197.520 68.855 198.030 ;
        RECT 66.835 197.220 67.290 197.390 ;
        RECT 69.025 197.350 69.355 197.860 ;
        RECT 69.525 197.520 70.155 198.030 ;
        RECT 70.735 197.520 71.115 197.690 ;
        RECT 71.285 197.520 71.585 198.030 ;
        RECT 70.945 197.350 71.115 197.520 ;
        RECT 65.355 196.720 65.570 197.050 ;
        RECT 64.785 196.390 65.095 196.720 ;
        RECT 65.265 196.390 65.570 196.720 ;
        RECT 65.745 196.390 66.030 197.050 ;
        RECT 66.225 196.390 66.490 197.050 ;
        RECT 66.705 196.390 66.950 197.050 ;
        RECT 64.925 196.220 65.095 196.390 ;
        RECT 67.120 196.220 67.290 197.220 ;
        RECT 63.955 195.480 64.245 196.205 ;
        RECT 64.425 195.695 64.755 196.205 ;
        RECT 64.925 196.050 67.290 196.220 ;
        RECT 68.555 197.180 70.775 197.350 ;
        RECT 68.555 196.220 68.725 197.180 ;
        RECT 68.895 196.840 70.435 197.010 ;
        RECT 68.895 196.390 69.140 196.840 ;
        RECT 69.400 196.470 70.095 196.670 ;
        RECT 70.265 196.640 70.435 196.840 ;
        RECT 70.605 196.980 70.775 197.180 ;
        RECT 70.945 197.150 71.605 197.350 ;
        RECT 70.605 196.810 71.265 196.980 ;
        RECT 70.265 196.470 70.865 196.640 ;
        RECT 71.095 196.390 71.265 196.810 ;
        RECT 64.925 195.480 65.255 195.880 ;
        RECT 66.305 195.710 66.635 196.050 ;
        RECT 66.805 195.480 67.135 195.880 ;
        RECT 68.555 195.675 69.020 196.220 ;
        RECT 69.525 195.480 69.695 196.300 ;
        RECT 69.865 196.220 70.775 196.300 ;
        RECT 71.435 196.220 71.605 197.150 ;
        RECT 69.865 196.130 71.115 196.220 ;
        RECT 69.865 195.650 70.195 196.130 ;
        RECT 70.605 196.050 71.115 196.130 ;
        RECT 70.365 195.480 70.715 195.870 ;
        RECT 70.885 195.650 71.115 196.050 ;
        RECT 71.285 195.740 71.605 196.220 ;
        RECT 71.780 196.840 72.035 197.720 ;
        RECT 72.205 196.890 72.510 198.030 ;
        RECT 72.850 197.650 73.180 198.030 ;
        RECT 73.360 197.480 73.530 197.770 ;
        RECT 73.700 197.570 73.950 198.030 ;
        RECT 72.730 197.310 73.530 197.480 ;
        RECT 74.120 197.520 74.990 197.860 ;
        RECT 71.780 196.190 71.990 196.840 ;
        RECT 72.730 196.720 72.900 197.310 ;
        RECT 74.120 197.140 74.290 197.520 ;
        RECT 75.225 197.400 75.395 197.860 ;
        RECT 75.565 197.570 75.935 198.030 ;
        RECT 76.230 197.430 76.400 197.770 ;
        RECT 76.570 197.600 76.900 198.030 ;
        RECT 77.135 197.430 77.305 197.770 ;
        RECT 73.070 196.970 74.290 197.140 ;
        RECT 74.460 197.060 74.920 197.350 ;
        RECT 75.225 197.230 75.785 197.400 ;
        RECT 76.230 197.260 77.305 197.430 ;
        RECT 77.475 197.530 78.155 197.860 ;
        RECT 78.370 197.530 78.620 197.860 ;
        RECT 78.790 197.570 79.040 198.030 ;
        RECT 75.615 197.090 75.785 197.230 ;
        RECT 74.460 197.050 75.425 197.060 ;
        RECT 74.120 196.880 74.290 196.970 ;
        RECT 74.750 196.890 75.425 197.050 ;
        RECT 72.160 196.690 72.900 196.720 ;
        RECT 72.160 196.390 73.075 196.690 ;
        RECT 72.750 196.215 73.075 196.390 ;
        RECT 71.780 195.660 72.035 196.190 ;
        RECT 72.205 195.480 72.510 195.940 ;
        RECT 72.755 195.860 73.075 196.215 ;
        RECT 73.245 196.430 73.785 196.800 ;
        RECT 74.120 196.710 74.525 196.880 ;
        RECT 73.245 196.030 73.485 196.430 ;
        RECT 73.965 196.260 74.185 196.540 ;
        RECT 73.655 196.090 74.185 196.260 ;
        RECT 73.655 195.860 73.825 196.090 ;
        RECT 74.355 195.930 74.525 196.710 ;
        RECT 74.695 196.100 75.045 196.720 ;
        RECT 75.215 196.100 75.425 196.890 ;
        RECT 75.615 196.920 77.115 197.090 ;
        RECT 75.615 196.230 75.785 196.920 ;
        RECT 77.475 196.750 77.645 197.530 ;
        RECT 78.450 197.400 78.620 197.530 ;
        RECT 75.955 196.580 77.645 196.750 ;
        RECT 77.815 196.970 78.280 197.360 ;
        RECT 78.450 197.230 78.845 197.400 ;
        RECT 75.955 196.400 76.125 196.580 ;
        RECT 72.755 195.690 73.825 195.860 ;
        RECT 73.995 195.480 74.185 195.920 ;
        RECT 74.355 195.650 75.305 195.930 ;
        RECT 75.615 195.840 75.875 196.230 ;
        RECT 76.295 196.160 77.085 196.410 ;
        RECT 75.525 195.670 75.875 195.840 ;
        RECT 76.085 195.480 76.415 195.940 ;
        RECT 77.290 195.870 77.460 196.580 ;
        RECT 77.815 196.380 77.985 196.970 ;
        RECT 77.630 196.160 77.985 196.380 ;
        RECT 78.155 196.160 78.505 196.780 ;
        RECT 78.675 195.870 78.845 197.230 ;
        RECT 79.210 197.060 79.535 197.845 ;
        RECT 79.015 196.010 79.475 197.060 ;
        RECT 77.290 195.700 78.145 195.870 ;
        RECT 78.350 195.700 78.845 195.870 ;
        RECT 79.015 195.480 79.345 195.840 ;
        RECT 79.705 195.740 79.875 197.860 ;
        RECT 80.045 197.530 80.375 198.030 ;
        RECT 80.545 197.360 80.800 197.860 ;
        RECT 80.050 197.190 80.800 197.360 ;
        RECT 80.050 196.200 80.280 197.190 ;
        RECT 80.450 196.370 80.800 197.020 ;
        RECT 81.435 196.940 84.025 198.030 ;
        RECT 84.200 197.595 89.545 198.030 ;
        RECT 81.435 196.420 82.645 196.940 ;
        RECT 82.815 196.250 84.025 196.770 ;
        RECT 85.790 196.345 86.140 197.595 ;
        RECT 89.715 196.865 90.005 198.030 ;
        RECT 90.635 196.940 92.305 198.030 ;
        RECT 92.480 197.595 97.825 198.030 ;
        RECT 98.000 197.595 103.345 198.030 ;
        RECT 103.520 197.595 108.865 198.030 ;
        RECT 109.040 197.595 114.385 198.030 ;
        RECT 80.050 196.030 80.800 196.200 ;
        RECT 80.045 195.480 80.375 195.860 ;
        RECT 80.545 195.740 80.800 196.030 ;
        RECT 81.435 195.480 84.025 196.250 ;
        RECT 87.620 196.025 87.960 196.855 ;
        RECT 90.635 196.420 91.385 196.940 ;
        RECT 91.555 196.250 92.305 196.770 ;
        RECT 94.070 196.345 94.420 197.595 ;
        RECT 84.200 195.480 89.545 196.025 ;
        RECT 89.715 195.480 90.005 196.205 ;
        RECT 90.635 195.480 92.305 196.250 ;
        RECT 95.900 196.025 96.240 196.855 ;
        RECT 99.590 196.345 99.940 197.595 ;
        RECT 101.420 196.025 101.760 196.855 ;
        RECT 105.110 196.345 105.460 197.595 ;
        RECT 106.940 196.025 107.280 196.855 ;
        RECT 110.630 196.345 110.980 197.595 ;
        RECT 114.555 196.940 115.765 198.030 ;
        RECT 112.460 196.025 112.800 196.855 ;
        RECT 114.555 196.400 115.075 196.940 ;
        RECT 115.245 196.230 115.765 196.770 ;
        RECT 92.480 195.480 97.825 196.025 ;
        RECT 98.000 195.480 103.345 196.025 ;
        RECT 103.520 195.480 108.865 196.025 ;
        RECT 109.040 195.480 114.385 196.025 ;
        RECT 114.555 195.480 115.765 196.230 ;
        RECT 10.510 195.310 115.850 195.480 ;
        RECT 10.595 194.560 11.805 195.310 ;
        RECT 10.595 194.020 11.115 194.560 ;
        RECT 12.435 194.540 14.105 195.310 ;
        RECT 14.280 194.765 19.625 195.310 ;
        RECT 19.800 194.765 25.145 195.310 ;
        RECT 11.285 193.850 11.805 194.390 ;
        RECT 10.595 192.760 11.805 193.850 ;
        RECT 12.435 193.850 13.185 194.370 ;
        RECT 13.355 194.020 14.105 194.540 ;
        RECT 12.435 192.760 14.105 193.850 ;
        RECT 15.870 193.195 16.220 194.445 ;
        RECT 17.700 193.935 18.040 194.765 ;
        RECT 21.390 193.195 21.740 194.445 ;
        RECT 23.220 193.935 23.560 194.765 ;
        RECT 25.315 194.585 25.605 195.310 ;
        RECT 25.780 194.765 31.125 195.310 ;
        RECT 31.300 194.765 36.645 195.310 ;
        RECT 36.820 194.765 42.165 195.310 ;
        RECT 14.280 192.760 19.625 193.195 ;
        RECT 19.800 192.760 25.145 193.195 ;
        RECT 25.315 192.760 25.605 193.925 ;
        RECT 27.370 193.195 27.720 194.445 ;
        RECT 29.200 193.935 29.540 194.765 ;
        RECT 32.890 193.195 33.240 194.445 ;
        RECT 34.720 193.935 35.060 194.765 ;
        RECT 38.410 193.195 38.760 194.445 ;
        RECT 40.240 193.935 40.580 194.765 ;
        RECT 42.375 194.490 42.605 195.310 ;
        RECT 42.775 194.510 43.105 195.140 ;
        RECT 42.355 194.070 42.685 194.320 ;
        RECT 42.855 193.910 43.105 194.510 ;
        RECT 43.275 194.490 43.485 195.310 ;
        RECT 43.715 194.540 45.385 195.310 ;
        RECT 45.560 194.765 50.905 195.310 ;
        RECT 25.780 192.760 31.125 193.195 ;
        RECT 31.300 192.760 36.645 193.195 ;
        RECT 36.820 192.760 42.165 193.195 ;
        RECT 42.375 192.760 42.605 193.900 ;
        RECT 42.775 192.930 43.105 193.910 ;
        RECT 43.275 192.760 43.485 193.900 ;
        RECT 43.715 193.850 44.465 194.370 ;
        RECT 44.635 194.020 45.385 194.540 ;
        RECT 43.715 192.760 45.385 193.850 ;
        RECT 47.150 193.195 47.500 194.445 ;
        RECT 48.980 193.935 49.320 194.765 ;
        RECT 51.075 194.585 51.365 195.310 ;
        RECT 51.535 194.540 54.125 195.310 ;
        RECT 45.560 192.760 50.905 193.195 ;
        RECT 51.075 192.760 51.365 193.925 ;
        RECT 51.535 193.850 52.745 194.370 ;
        RECT 52.915 194.020 54.125 194.540 ;
        RECT 54.355 194.490 54.565 195.310 ;
        RECT 54.735 194.510 55.065 195.140 ;
        RECT 54.735 193.910 54.985 194.510 ;
        RECT 55.235 194.490 55.465 195.310 ;
        RECT 56.250 194.680 56.535 195.140 ;
        RECT 56.705 194.850 56.975 195.310 ;
        RECT 56.250 194.510 57.205 194.680 ;
        RECT 55.155 194.070 55.485 194.320 ;
        RECT 51.535 192.760 54.125 193.850 ;
        RECT 54.355 192.760 54.565 193.900 ;
        RECT 54.735 192.930 55.065 193.910 ;
        RECT 55.235 192.760 55.465 193.900 ;
        RECT 56.135 193.780 56.825 194.340 ;
        RECT 56.995 193.610 57.205 194.510 ;
        RECT 56.250 193.390 57.205 193.610 ;
        RECT 57.375 194.340 57.775 195.140 ;
        RECT 57.965 194.680 58.245 195.140 ;
        RECT 58.765 194.850 59.090 195.310 ;
        RECT 57.965 194.510 59.090 194.680 ;
        RECT 59.260 194.570 59.645 195.140 ;
        RECT 58.640 194.400 59.090 194.510 ;
        RECT 57.375 193.780 58.470 194.340 ;
        RECT 58.640 194.070 59.195 194.400 ;
        RECT 56.250 192.930 56.535 193.390 ;
        RECT 56.705 192.760 56.975 193.220 ;
        RECT 57.375 192.930 57.775 193.780 ;
        RECT 58.640 193.610 59.090 194.070 ;
        RECT 59.365 193.900 59.645 194.570 ;
        RECT 59.815 194.560 61.025 195.310 ;
        RECT 57.965 193.390 59.090 193.610 ;
        RECT 57.965 192.930 58.245 193.390 ;
        RECT 58.765 192.760 59.090 193.220 ;
        RECT 59.260 192.930 59.645 193.900 ;
        RECT 59.815 193.850 60.335 194.390 ;
        RECT 60.505 194.020 61.025 194.560 ;
        RECT 61.195 194.490 61.455 195.310 ;
        RECT 61.625 194.490 61.955 194.910 ;
        RECT 62.135 194.740 62.395 195.140 ;
        RECT 62.565 194.910 62.895 195.310 ;
        RECT 63.065 194.740 63.235 195.090 ;
        RECT 63.405 194.910 63.780 195.310 ;
        RECT 64.420 195.055 64.755 195.100 ;
        RECT 62.135 194.570 63.800 194.740 ;
        RECT 63.970 194.635 64.245 194.980 ;
        RECT 61.705 194.400 61.955 194.490 ;
        RECT 63.630 194.400 63.800 194.570 ;
        RECT 61.200 194.070 61.535 194.320 ;
        RECT 61.705 194.070 62.420 194.400 ;
        RECT 62.635 194.070 63.460 194.400 ;
        RECT 63.630 194.070 63.905 194.400 ;
        RECT 59.815 192.760 61.025 193.850 ;
        RECT 61.195 192.760 61.455 193.900 ;
        RECT 61.705 193.510 61.875 194.070 ;
        RECT 62.135 193.610 62.465 193.900 ;
        RECT 62.635 193.780 62.880 194.070 ;
        RECT 63.630 193.900 63.800 194.070 ;
        RECT 64.075 193.900 64.245 194.635 ;
        RECT 63.140 193.730 63.800 193.900 ;
        RECT 63.140 193.610 63.310 193.730 ;
        RECT 62.135 193.440 63.310 193.610 ;
        RECT 61.695 192.940 63.310 193.270 ;
        RECT 63.480 192.760 63.760 193.560 ;
        RECT 63.970 192.930 64.245 193.900 ;
        RECT 64.415 194.590 64.755 195.055 ;
        RECT 64.925 194.930 65.255 195.310 ;
        RECT 64.415 193.900 64.585 194.590 ;
        RECT 64.755 194.070 65.015 194.400 ;
        RECT 64.415 192.930 64.675 193.900 ;
        RECT 64.845 193.520 65.015 194.070 ;
        RECT 65.185 193.700 65.525 194.730 ;
        RECT 65.715 193.950 65.985 194.975 ;
        RECT 65.715 193.780 66.025 193.950 ;
        RECT 65.715 193.700 65.985 193.780 ;
        RECT 66.210 193.700 66.490 194.975 ;
        RECT 66.690 194.810 66.920 195.140 ;
        RECT 67.165 194.930 67.495 195.310 ;
        RECT 66.690 193.520 66.860 194.810 ;
        RECT 67.665 194.740 67.840 195.140 ;
        RECT 69.180 194.800 69.420 195.310 ;
        RECT 69.600 194.800 69.880 195.130 ;
        RECT 70.110 194.800 70.325 195.310 ;
        RECT 67.210 194.570 67.840 194.740 ;
        RECT 67.210 194.400 67.380 194.570 ;
        RECT 67.030 194.070 67.380 194.400 ;
        RECT 64.845 193.350 66.860 193.520 ;
        RECT 67.210 193.550 67.380 194.070 ;
        RECT 67.560 193.720 67.925 194.400 ;
        RECT 69.075 194.070 69.430 194.630 ;
        RECT 69.600 193.900 69.770 194.800 ;
        RECT 69.940 194.070 70.205 194.630 ;
        RECT 70.495 194.570 71.110 195.140 ;
        RECT 71.315 194.930 72.205 195.100 ;
        RECT 70.455 193.900 70.625 194.400 ;
        RECT 69.200 193.730 70.625 193.900 ;
        RECT 69.200 193.555 69.590 193.730 ;
        RECT 67.210 193.380 67.840 193.550 ;
        RECT 64.870 192.760 65.200 193.170 ;
        RECT 65.400 192.930 65.570 193.350 ;
        RECT 65.785 192.760 66.455 193.170 ;
        RECT 66.690 192.930 66.860 193.350 ;
        RECT 67.165 192.760 67.495 193.200 ;
        RECT 67.665 192.930 67.840 193.380 ;
        RECT 70.075 192.760 70.405 193.560 ;
        RECT 70.795 193.550 71.110 194.570 ;
        RECT 71.315 194.375 71.865 194.760 ;
        RECT 72.035 194.205 72.205 194.930 ;
        RECT 71.315 194.135 72.205 194.205 ;
        RECT 72.375 194.605 72.595 195.090 ;
        RECT 72.765 194.770 73.015 195.310 ;
        RECT 73.185 194.660 73.445 195.140 ;
        RECT 72.375 194.180 72.705 194.605 ;
        RECT 71.315 194.110 72.210 194.135 ;
        RECT 71.315 194.095 72.220 194.110 ;
        RECT 71.315 194.080 72.225 194.095 ;
        RECT 71.315 194.075 72.235 194.080 ;
        RECT 71.315 194.065 72.240 194.075 ;
        RECT 71.315 194.055 72.245 194.065 ;
        RECT 71.315 194.050 72.255 194.055 ;
        RECT 71.315 194.040 72.265 194.050 ;
        RECT 71.315 194.035 72.275 194.040 ;
        RECT 71.315 193.585 71.575 194.035 ;
        RECT 71.940 194.030 72.275 194.035 ;
        RECT 71.940 194.025 72.290 194.030 ;
        RECT 71.940 194.015 72.305 194.025 ;
        RECT 71.940 194.010 72.330 194.015 ;
        RECT 72.875 194.010 73.105 194.405 ;
        RECT 71.940 194.005 73.105 194.010 ;
        RECT 71.970 193.970 73.105 194.005 ;
        RECT 72.005 193.945 73.105 193.970 ;
        RECT 72.035 193.915 73.105 193.945 ;
        RECT 72.055 193.885 73.105 193.915 ;
        RECT 72.075 193.855 73.105 193.885 ;
        RECT 72.145 193.845 73.105 193.855 ;
        RECT 72.170 193.835 73.105 193.845 ;
        RECT 72.190 193.820 73.105 193.835 ;
        RECT 72.210 193.805 73.105 193.820 ;
        RECT 72.215 193.795 73.000 193.805 ;
        RECT 72.230 193.760 73.000 193.795 ;
        RECT 70.575 192.930 71.110 193.550 ;
        RECT 71.745 193.440 72.075 193.685 ;
        RECT 72.245 193.510 73.000 193.760 ;
        RECT 73.275 193.630 73.445 194.660 ;
        RECT 74.115 194.490 74.345 195.310 ;
        RECT 74.515 194.510 74.845 195.140 ;
        RECT 74.095 194.070 74.425 194.320 ;
        RECT 74.595 193.910 74.845 194.510 ;
        RECT 75.015 194.490 75.225 195.310 ;
        RECT 75.495 194.490 75.725 195.310 ;
        RECT 75.895 194.510 76.225 195.140 ;
        RECT 75.475 194.070 75.805 194.320 ;
        RECT 75.975 193.910 76.225 194.510 ;
        RECT 76.395 194.490 76.605 195.310 ;
        RECT 76.835 194.585 77.125 195.310 ;
        RECT 78.215 194.540 81.725 195.310 ;
        RECT 81.900 194.765 87.245 195.310 ;
        RECT 71.745 193.415 71.930 193.440 ;
        RECT 71.315 193.315 71.930 193.415 ;
        RECT 71.315 192.760 71.920 193.315 ;
        RECT 72.095 192.930 72.575 193.270 ;
        RECT 72.745 192.760 73.000 193.305 ;
        RECT 73.170 192.930 73.445 193.630 ;
        RECT 74.115 192.760 74.345 193.900 ;
        RECT 74.515 192.930 74.845 193.910 ;
        RECT 75.015 192.760 75.225 193.900 ;
        RECT 75.495 192.760 75.725 193.900 ;
        RECT 75.895 192.930 76.225 193.910 ;
        RECT 76.395 192.760 76.605 193.900 ;
        RECT 76.835 192.760 77.125 193.925 ;
        RECT 78.215 193.850 79.905 194.370 ;
        RECT 80.075 194.020 81.725 194.540 ;
        RECT 78.215 192.760 81.725 193.850 ;
        RECT 83.490 193.195 83.840 194.445 ;
        RECT 85.320 193.935 85.660 194.765 ;
        RECT 87.420 194.760 87.675 195.050 ;
        RECT 87.845 194.930 88.175 195.310 ;
        RECT 87.420 194.590 88.170 194.760 ;
        RECT 87.420 193.770 87.770 194.420 ;
        RECT 87.940 193.600 88.170 194.590 ;
        RECT 87.420 193.430 88.170 193.600 ;
        RECT 81.900 192.760 87.245 193.195 ;
        RECT 87.420 192.930 87.675 193.430 ;
        RECT 87.845 192.760 88.175 193.260 ;
        RECT 88.345 192.930 88.515 195.050 ;
        RECT 88.875 194.950 89.205 195.310 ;
        RECT 89.375 194.920 89.870 195.090 ;
        RECT 90.075 194.920 90.930 195.090 ;
        RECT 88.745 193.730 89.205 194.780 ;
        RECT 88.685 192.945 89.010 193.730 ;
        RECT 89.375 193.560 89.545 194.920 ;
        RECT 89.715 194.010 90.065 194.630 ;
        RECT 90.235 194.410 90.590 194.630 ;
        RECT 90.235 193.820 90.405 194.410 ;
        RECT 90.760 194.210 90.930 194.920 ;
        RECT 91.805 194.850 92.135 195.310 ;
        RECT 92.345 194.950 92.695 195.120 ;
        RECT 91.135 194.380 91.925 194.630 ;
        RECT 92.345 194.560 92.605 194.950 ;
        RECT 92.915 194.860 93.865 195.140 ;
        RECT 94.035 194.870 94.225 195.310 ;
        RECT 94.395 194.930 95.465 195.100 ;
        RECT 92.095 194.210 92.265 194.390 ;
        RECT 89.375 193.390 89.770 193.560 ;
        RECT 89.940 193.430 90.405 193.820 ;
        RECT 90.575 194.040 92.265 194.210 ;
        RECT 89.600 193.260 89.770 193.390 ;
        RECT 90.575 193.260 90.745 194.040 ;
        RECT 92.435 193.870 92.605 194.560 ;
        RECT 91.105 193.700 92.605 193.870 ;
        RECT 92.795 193.900 93.005 194.690 ;
        RECT 93.175 194.070 93.525 194.690 ;
        RECT 93.695 194.080 93.865 194.860 ;
        RECT 94.395 194.700 94.565 194.930 ;
        RECT 94.035 194.530 94.565 194.700 ;
        RECT 94.035 194.250 94.255 194.530 ;
        RECT 94.735 194.360 94.975 194.760 ;
        RECT 93.695 193.910 94.100 194.080 ;
        RECT 94.435 193.990 94.975 194.360 ;
        RECT 95.145 194.575 95.465 194.930 ;
        RECT 95.710 194.850 96.015 195.310 ;
        RECT 96.185 194.600 96.440 195.130 ;
        RECT 95.145 194.400 95.470 194.575 ;
        RECT 95.145 194.100 96.060 194.400 ;
        RECT 95.320 194.070 96.060 194.100 ;
        RECT 92.795 193.740 93.470 193.900 ;
        RECT 93.930 193.820 94.100 193.910 ;
        RECT 92.795 193.730 93.760 193.740 ;
        RECT 92.435 193.560 92.605 193.700 ;
        RECT 89.180 192.760 89.430 193.220 ;
        RECT 89.600 192.930 89.850 193.260 ;
        RECT 90.065 192.930 90.745 193.260 ;
        RECT 90.915 193.360 91.990 193.530 ;
        RECT 92.435 193.390 92.995 193.560 ;
        RECT 93.300 193.440 93.760 193.730 ;
        RECT 93.930 193.650 95.150 193.820 ;
        RECT 90.915 193.020 91.085 193.360 ;
        RECT 91.320 192.760 91.650 193.190 ;
        RECT 91.820 193.020 91.990 193.360 ;
        RECT 92.285 192.760 92.655 193.220 ;
        RECT 92.825 192.930 92.995 193.390 ;
        RECT 93.930 193.270 94.100 193.650 ;
        RECT 95.320 193.480 95.490 194.070 ;
        RECT 96.230 193.950 96.440 194.600 ;
        RECT 97.535 194.540 101.045 195.310 ;
        RECT 93.230 192.930 94.100 193.270 ;
        RECT 94.690 193.310 95.490 193.480 ;
        RECT 94.270 192.760 94.520 193.220 ;
        RECT 94.690 193.020 94.860 193.310 ;
        RECT 95.040 192.760 95.370 193.140 ;
        RECT 95.710 192.760 96.015 193.900 ;
        RECT 96.185 193.070 96.440 193.950 ;
        RECT 97.535 193.850 99.225 194.370 ;
        RECT 99.395 194.020 101.045 194.540 ;
        RECT 101.275 194.490 101.485 195.310 ;
        RECT 101.655 194.510 101.985 195.140 ;
        RECT 101.655 193.910 101.905 194.510 ;
        RECT 102.155 194.490 102.385 195.310 ;
        RECT 102.595 194.585 102.885 195.310 ;
        RECT 104.065 194.760 104.235 195.140 ;
        RECT 104.415 194.930 104.745 195.310 ;
        RECT 104.065 194.590 104.730 194.760 ;
        RECT 104.925 194.635 105.185 195.140 ;
        RECT 102.075 194.070 102.405 194.320 ;
        RECT 103.995 194.040 104.325 194.410 ;
        RECT 104.560 194.335 104.730 194.590 ;
        RECT 104.560 194.005 104.845 194.335 ;
        RECT 97.535 192.760 101.045 193.850 ;
        RECT 101.275 192.760 101.485 193.900 ;
        RECT 101.655 192.930 101.985 193.910 ;
        RECT 102.155 192.760 102.385 193.900 ;
        RECT 102.595 192.760 102.885 193.925 ;
        RECT 104.560 193.860 104.730 194.005 ;
        RECT 104.065 193.690 104.730 193.860 ;
        RECT 105.015 193.835 105.185 194.635 ;
        RECT 105.355 194.540 108.865 195.310 ;
        RECT 109.040 194.765 114.385 195.310 ;
        RECT 104.065 192.930 104.235 193.690 ;
        RECT 104.415 192.760 104.745 193.520 ;
        RECT 104.915 192.930 105.185 193.835 ;
        RECT 105.355 193.850 107.045 194.370 ;
        RECT 107.215 194.020 108.865 194.540 ;
        RECT 105.355 192.760 108.865 193.850 ;
        RECT 110.630 193.195 110.980 194.445 ;
        RECT 112.460 193.935 112.800 194.765 ;
        RECT 114.555 194.560 115.765 195.310 ;
        RECT 114.555 193.850 115.075 194.390 ;
        RECT 115.245 194.020 115.765 194.560 ;
        RECT 109.040 192.760 114.385 193.195 ;
        RECT 114.555 192.760 115.765 193.850 ;
        RECT 10.510 192.590 115.850 192.760 ;
        RECT 10.595 191.500 11.805 192.590 ;
        RECT 10.595 190.790 11.115 191.330 ;
        RECT 11.285 190.960 11.805 191.500 ;
        RECT 12.435 191.425 12.725 192.590 ;
        RECT 13.815 191.500 17.325 192.590 ;
        RECT 17.500 192.155 22.845 192.590 ;
        RECT 13.815 190.980 15.505 191.500 ;
        RECT 15.675 190.810 17.325 191.330 ;
        RECT 19.090 190.905 19.440 192.155 ;
        RECT 23.390 191.610 23.645 192.280 ;
        RECT 23.825 191.790 24.110 192.590 ;
        RECT 24.290 191.870 24.620 192.380 ;
        RECT 10.595 190.040 11.805 190.790 ;
        RECT 12.435 190.040 12.725 190.765 ;
        RECT 13.815 190.040 17.325 190.810 ;
        RECT 20.920 190.585 21.260 191.415 ;
        RECT 23.390 190.750 23.570 191.610 ;
        RECT 24.290 191.280 24.540 191.870 ;
        RECT 24.890 191.720 25.060 192.330 ;
        RECT 25.230 191.900 25.560 192.590 ;
        RECT 25.790 192.040 26.030 192.330 ;
        RECT 26.230 192.210 26.650 192.590 ;
        RECT 26.830 192.120 27.460 192.370 ;
        RECT 27.930 192.210 28.260 192.590 ;
        RECT 26.830 192.040 27.000 192.120 ;
        RECT 28.430 192.040 28.600 192.330 ;
        RECT 28.780 192.210 29.160 192.590 ;
        RECT 29.400 192.205 30.230 192.375 ;
        RECT 25.790 191.870 27.000 192.040 ;
        RECT 23.740 190.950 24.540 191.280 ;
        RECT 17.500 190.040 22.845 190.585 ;
        RECT 23.390 190.550 23.645 190.750 ;
        RECT 23.305 190.380 23.645 190.550 ;
        RECT 23.390 190.220 23.645 190.380 ;
        RECT 23.825 190.040 24.110 190.500 ;
        RECT 24.290 190.300 24.540 190.950 ;
        RECT 24.740 191.700 25.060 191.720 ;
        RECT 24.740 191.530 26.660 191.700 ;
        RECT 24.740 190.635 24.930 191.530 ;
        RECT 26.830 191.360 27.000 191.870 ;
        RECT 27.170 191.610 27.690 191.920 ;
        RECT 25.100 191.190 27.000 191.360 ;
        RECT 25.100 191.130 25.430 191.190 ;
        RECT 25.580 190.960 25.910 191.020 ;
        RECT 25.250 190.690 25.910 190.960 ;
        RECT 24.740 190.305 25.060 190.635 ;
        RECT 25.240 190.040 25.900 190.520 ;
        RECT 26.100 190.430 26.270 191.190 ;
        RECT 27.170 191.020 27.350 191.430 ;
        RECT 26.440 190.850 26.770 190.970 ;
        RECT 27.520 190.850 27.690 191.610 ;
        RECT 26.440 190.680 27.690 190.850 ;
        RECT 27.860 191.790 29.230 192.040 ;
        RECT 27.860 191.020 28.050 191.790 ;
        RECT 28.980 191.530 29.230 191.790 ;
        RECT 28.220 191.360 28.470 191.520 ;
        RECT 29.400 191.360 29.570 192.205 ;
        RECT 30.465 191.920 30.635 192.420 ;
        RECT 30.805 192.090 31.135 192.590 ;
        RECT 29.740 191.530 30.240 191.910 ;
        RECT 30.465 191.750 31.160 191.920 ;
        RECT 28.220 191.190 29.570 191.360 ;
        RECT 29.150 191.150 29.570 191.190 ;
        RECT 27.860 190.680 28.280 191.020 ;
        RECT 28.570 190.690 28.980 191.020 ;
        RECT 26.100 190.260 26.950 190.430 ;
        RECT 27.510 190.040 27.830 190.500 ;
        RECT 28.030 190.250 28.280 190.680 ;
        RECT 28.570 190.040 28.980 190.480 ;
        RECT 29.150 190.420 29.320 191.150 ;
        RECT 29.490 190.600 29.840 190.970 ;
        RECT 30.020 190.660 30.240 191.530 ;
        RECT 30.410 190.960 30.820 191.580 ;
        RECT 30.990 190.780 31.160 191.750 ;
        RECT 30.465 190.590 31.160 190.780 ;
        RECT 29.150 190.220 30.165 190.420 ;
        RECT 30.465 190.260 30.635 190.590 ;
        RECT 30.805 190.040 31.135 190.420 ;
        RECT 31.350 190.300 31.575 192.420 ;
        RECT 31.745 192.090 32.075 192.590 ;
        RECT 32.245 191.920 32.415 192.420 ;
        RECT 32.680 192.155 38.025 192.590 ;
        RECT 31.750 191.750 32.415 191.920 ;
        RECT 31.750 190.760 31.980 191.750 ;
        RECT 32.150 190.930 32.500 191.580 ;
        RECT 34.270 190.905 34.620 192.155 ;
        RECT 38.195 191.425 38.485 192.590 ;
        RECT 39.635 191.450 39.845 192.590 ;
        RECT 40.015 191.440 40.345 192.420 ;
        RECT 40.515 191.450 40.745 192.590 ;
        RECT 41.070 191.960 41.355 192.420 ;
        RECT 41.525 192.130 41.795 192.590 ;
        RECT 41.070 191.740 42.025 191.960 ;
        RECT 31.750 190.590 32.415 190.760 ;
        RECT 31.745 190.040 32.075 190.420 ;
        RECT 32.245 190.300 32.415 190.590 ;
        RECT 36.100 190.585 36.440 191.415 ;
        RECT 32.680 190.040 38.025 190.585 ;
        RECT 38.195 190.040 38.485 190.765 ;
        RECT 39.635 190.040 39.845 190.860 ;
        RECT 40.015 190.840 40.265 191.440 ;
        RECT 40.435 191.030 40.765 191.280 ;
        RECT 40.955 191.010 41.645 191.570 ;
        RECT 40.015 190.210 40.345 190.840 ;
        RECT 40.515 190.040 40.745 190.860 ;
        RECT 41.815 190.840 42.025 191.740 ;
        RECT 41.070 190.670 42.025 190.840 ;
        RECT 42.195 191.570 42.595 192.420 ;
        RECT 42.785 191.960 43.065 192.420 ;
        RECT 43.585 192.130 43.910 192.590 ;
        RECT 42.785 191.740 43.910 191.960 ;
        RECT 42.195 191.010 43.290 191.570 ;
        RECT 43.460 191.280 43.910 191.740 ;
        RECT 44.080 191.450 44.465 192.420 ;
        RECT 45.645 191.660 45.815 192.420 ;
        RECT 45.995 191.830 46.325 192.590 ;
        RECT 45.645 191.490 46.310 191.660 ;
        RECT 46.495 191.515 46.765 192.420 ;
        RECT 47.860 192.155 53.205 192.590 ;
        RECT 53.380 192.155 58.725 192.590 ;
        RECT 41.070 190.210 41.355 190.670 ;
        RECT 41.525 190.040 41.795 190.500 ;
        RECT 42.195 190.210 42.595 191.010 ;
        RECT 43.460 190.950 44.015 191.280 ;
        RECT 43.460 190.840 43.910 190.950 ;
        RECT 42.785 190.670 43.910 190.840 ;
        RECT 44.185 190.780 44.465 191.450 ;
        RECT 46.140 191.345 46.310 191.490 ;
        RECT 45.575 190.940 45.905 191.310 ;
        RECT 46.140 191.015 46.425 191.345 ;
        RECT 42.785 190.210 43.065 190.670 ;
        RECT 43.585 190.040 43.910 190.500 ;
        RECT 44.080 190.210 44.465 190.780 ;
        RECT 46.140 190.760 46.310 191.015 ;
        RECT 45.645 190.590 46.310 190.760 ;
        RECT 46.595 190.715 46.765 191.515 ;
        RECT 49.450 190.905 49.800 192.155 ;
        RECT 45.645 190.210 45.815 190.590 ;
        RECT 45.995 190.040 46.325 190.420 ;
        RECT 46.505 190.210 46.765 190.715 ;
        RECT 51.280 190.585 51.620 191.415 ;
        RECT 54.970 190.905 55.320 192.155 ;
        RECT 58.895 191.450 59.155 192.590 ;
        RECT 59.325 191.620 59.655 192.420 ;
        RECT 59.825 191.790 59.995 192.590 ;
        RECT 60.195 191.620 60.525 192.420 ;
        RECT 60.725 191.790 61.005 192.590 ;
        RECT 59.325 191.450 60.605 191.620 ;
        RECT 56.800 190.585 57.140 191.415 ;
        RECT 58.920 190.950 59.205 191.280 ;
        RECT 59.405 190.950 59.785 191.280 ;
        RECT 59.955 190.950 60.265 191.280 ;
        RECT 47.860 190.040 53.205 190.585 ;
        RECT 53.380 190.040 58.725 190.585 ;
        RECT 58.900 190.040 59.235 190.780 ;
        RECT 59.405 190.255 59.620 190.950 ;
        RECT 59.955 190.780 60.160 190.950 ;
        RECT 60.435 190.780 60.605 191.450 ;
        RECT 60.785 190.950 61.025 191.620 ;
        RECT 61.195 191.500 63.785 192.590 ;
        RECT 61.195 190.980 62.405 191.500 ;
        RECT 63.955 191.425 64.245 192.590 ;
        RECT 62.575 190.810 63.785 191.330 ;
        RECT 59.810 190.255 60.160 190.780 ;
        RECT 60.330 190.210 61.025 190.780 ;
        RECT 61.195 190.040 63.785 190.810 ;
        RECT 63.955 190.040 64.245 190.765 ;
        RECT 65.335 190.210 65.595 192.420 ;
        RECT 65.765 192.210 66.095 192.590 ;
        RECT 66.520 192.040 66.690 192.420 ;
        RECT 66.950 192.210 67.280 192.590 ;
        RECT 67.475 192.040 67.645 192.420 ;
        RECT 67.855 192.210 68.185 192.590 ;
        RECT 68.435 192.040 68.625 192.420 ;
        RECT 68.865 192.210 69.195 192.590 ;
        RECT 69.505 192.090 69.765 192.420 ;
        RECT 65.765 191.870 67.715 192.040 ;
        RECT 65.765 190.950 65.935 191.870 ;
        RECT 66.305 191.280 66.500 191.590 ;
        RECT 66.770 191.280 66.955 191.590 ;
        RECT 66.245 190.950 66.500 191.280 ;
        RECT 66.725 190.950 66.955 191.280 ;
        RECT 65.765 190.040 66.095 190.420 ;
        RECT 66.305 190.375 66.500 190.950 ;
        RECT 66.770 190.370 66.955 190.950 ;
        RECT 67.205 190.380 67.375 191.280 ;
        RECT 67.545 190.880 67.715 191.870 ;
        RECT 67.885 191.870 68.625 192.040 ;
        RECT 67.885 191.360 68.055 191.870 ;
        RECT 68.225 191.530 68.805 191.700 ;
        RECT 69.075 191.580 69.425 191.910 ;
        RECT 68.635 191.410 68.805 191.530 ;
        RECT 69.595 191.410 69.765 192.090 ;
        RECT 67.885 191.190 68.455 191.360 ;
        RECT 68.635 191.240 69.765 191.410 ;
        RECT 67.545 190.550 68.095 190.880 ;
        RECT 68.285 190.710 68.455 191.190 ;
        RECT 68.625 190.900 69.245 191.070 ;
        RECT 69.035 190.720 69.245 190.900 ;
        RECT 68.285 190.380 68.685 190.710 ;
        RECT 69.595 190.540 69.765 191.240 ;
        RECT 67.205 190.210 68.685 190.380 ;
        RECT 68.865 190.040 69.195 190.420 ;
        RECT 69.505 190.210 69.765 190.540 ;
        RECT 69.935 191.450 70.320 192.420 ;
        RECT 70.490 192.130 70.815 192.590 ;
        RECT 71.335 191.960 71.615 192.420 ;
        RECT 70.490 191.740 71.615 191.960 ;
        RECT 69.935 190.780 70.215 191.450 ;
        RECT 70.490 191.280 70.940 191.740 ;
        RECT 71.805 191.570 72.205 192.420 ;
        RECT 72.605 192.130 72.875 192.590 ;
        RECT 73.045 191.960 73.330 192.420 ;
        RECT 70.385 190.950 70.940 191.280 ;
        RECT 71.110 191.010 72.205 191.570 ;
        RECT 70.490 190.840 70.940 190.950 ;
        RECT 69.935 190.210 70.320 190.780 ;
        RECT 70.490 190.670 71.615 190.840 ;
        RECT 70.490 190.040 70.815 190.500 ;
        RECT 71.335 190.210 71.615 190.670 ;
        RECT 71.805 190.210 72.205 191.010 ;
        RECT 72.375 191.740 73.330 191.960 ;
        RECT 72.375 190.840 72.585 191.740 ;
        RECT 72.755 191.010 73.445 191.570 ;
        RECT 73.615 191.500 74.825 192.590 ;
        RECT 75.000 192.155 80.345 192.590 ;
        RECT 73.615 190.960 74.135 191.500 ;
        RECT 72.375 190.670 73.330 190.840 ;
        RECT 74.305 190.790 74.825 191.330 ;
        RECT 76.590 190.905 76.940 192.155 ;
        RECT 80.555 191.450 80.785 192.590 ;
        RECT 80.955 191.440 81.285 192.420 ;
        RECT 81.455 191.450 81.665 192.590 ;
        RECT 81.985 191.660 82.155 192.420 ;
        RECT 82.335 191.830 82.665 192.590 ;
        RECT 81.985 191.490 82.650 191.660 ;
        RECT 82.835 191.515 83.105 192.420 ;
        RECT 72.605 190.040 72.875 190.500 ;
        RECT 73.045 190.210 73.330 190.670 ;
        RECT 73.615 190.040 74.825 190.790 ;
        RECT 78.420 190.585 78.760 191.415 ;
        RECT 80.535 191.030 80.865 191.280 ;
        RECT 75.000 190.040 80.345 190.585 ;
        RECT 80.555 190.040 80.785 190.860 ;
        RECT 81.035 190.840 81.285 191.440 ;
        RECT 82.480 191.345 82.650 191.490 ;
        RECT 81.915 190.940 82.245 191.310 ;
        RECT 82.480 191.015 82.765 191.345 ;
        RECT 80.955 190.210 81.285 190.840 ;
        RECT 81.455 190.040 81.665 190.860 ;
        RECT 82.480 190.760 82.650 191.015 ;
        RECT 81.985 190.590 82.650 190.760 ;
        RECT 82.935 190.715 83.105 191.515 ;
        RECT 83.275 191.500 84.485 192.590 ;
        RECT 84.655 191.500 88.165 192.590 ;
        RECT 83.275 190.960 83.795 191.500 ;
        RECT 83.965 190.790 84.485 191.330 ;
        RECT 84.655 190.980 86.345 191.500 ;
        RECT 88.375 191.450 88.605 192.590 ;
        RECT 88.775 191.440 89.105 192.420 ;
        RECT 89.275 191.450 89.485 192.590 ;
        RECT 86.515 190.810 88.165 191.330 ;
        RECT 88.355 191.030 88.685 191.280 ;
        RECT 81.985 190.210 82.155 190.590 ;
        RECT 82.335 190.040 82.665 190.420 ;
        RECT 82.845 190.210 83.105 190.715 ;
        RECT 83.275 190.040 84.485 190.790 ;
        RECT 84.655 190.040 88.165 190.810 ;
        RECT 88.375 190.040 88.605 190.860 ;
        RECT 88.855 190.840 89.105 191.440 ;
        RECT 89.715 191.425 90.005 192.590 ;
        RECT 90.175 191.450 90.560 192.420 ;
        RECT 90.730 192.130 91.055 192.590 ;
        RECT 91.575 191.960 91.855 192.420 ;
        RECT 90.730 191.740 91.855 191.960 ;
        RECT 88.775 190.210 89.105 190.840 ;
        RECT 89.275 190.040 89.485 190.860 ;
        RECT 90.175 190.780 90.455 191.450 ;
        RECT 90.730 191.280 91.180 191.740 ;
        RECT 92.045 191.570 92.445 192.420 ;
        RECT 92.845 192.130 93.115 192.590 ;
        RECT 93.285 191.960 93.570 192.420 ;
        RECT 90.625 190.950 91.180 191.280 ;
        RECT 91.350 191.010 92.445 191.570 ;
        RECT 90.730 190.840 91.180 190.950 ;
        RECT 89.715 190.040 90.005 190.765 ;
        RECT 90.175 190.210 90.560 190.780 ;
        RECT 90.730 190.670 91.855 190.840 ;
        RECT 90.730 190.040 91.055 190.500 ;
        RECT 91.575 190.210 91.855 190.670 ;
        RECT 92.045 190.210 92.445 191.010 ;
        RECT 92.615 191.740 93.570 191.960 ;
        RECT 94.890 191.960 95.175 192.420 ;
        RECT 95.345 192.130 95.615 192.590 ;
        RECT 94.890 191.740 95.845 191.960 ;
        RECT 92.615 190.840 92.825 191.740 ;
        RECT 92.995 191.010 93.685 191.570 ;
        RECT 94.775 191.010 95.465 191.570 ;
        RECT 95.635 190.840 95.845 191.740 ;
        RECT 92.615 190.670 93.570 190.840 ;
        RECT 92.845 190.040 93.115 190.500 ;
        RECT 93.285 190.210 93.570 190.670 ;
        RECT 94.890 190.670 95.845 190.840 ;
        RECT 96.015 191.570 96.415 192.420 ;
        RECT 96.605 191.960 96.885 192.420 ;
        RECT 97.405 192.130 97.730 192.590 ;
        RECT 96.605 191.740 97.730 191.960 ;
        RECT 96.015 191.010 97.110 191.570 ;
        RECT 97.280 191.280 97.730 191.740 ;
        RECT 97.900 191.450 98.285 192.420 ;
        RECT 94.890 190.210 95.175 190.670 ;
        RECT 95.345 190.040 95.615 190.500 ;
        RECT 96.015 190.210 96.415 191.010 ;
        RECT 97.280 190.950 97.835 191.280 ;
        RECT 97.280 190.840 97.730 190.950 ;
        RECT 96.605 190.670 97.730 190.840 ;
        RECT 98.005 190.780 98.285 191.450 ;
        RECT 96.605 190.210 96.885 190.670 ;
        RECT 97.405 190.040 97.730 190.500 ;
        RECT 97.900 190.210 98.285 190.780 ;
        RECT 98.460 191.400 98.715 192.280 ;
        RECT 98.885 191.450 99.190 192.590 ;
        RECT 99.530 192.210 99.860 192.590 ;
        RECT 100.040 192.040 100.210 192.330 ;
        RECT 100.380 192.130 100.630 192.590 ;
        RECT 99.410 191.870 100.210 192.040 ;
        RECT 100.800 192.080 101.670 192.420 ;
        RECT 98.460 190.750 98.670 191.400 ;
        RECT 99.410 191.280 99.580 191.870 ;
        RECT 100.800 191.700 100.970 192.080 ;
        RECT 101.905 191.960 102.075 192.420 ;
        RECT 102.245 192.130 102.615 192.590 ;
        RECT 102.910 191.990 103.080 192.330 ;
        RECT 103.250 192.160 103.580 192.590 ;
        RECT 103.815 191.990 103.985 192.330 ;
        RECT 99.750 191.530 100.970 191.700 ;
        RECT 101.140 191.620 101.600 191.910 ;
        RECT 101.905 191.790 102.465 191.960 ;
        RECT 102.910 191.820 103.985 191.990 ;
        RECT 104.155 192.090 104.835 192.420 ;
        RECT 105.050 192.090 105.300 192.420 ;
        RECT 105.470 192.130 105.720 192.590 ;
        RECT 102.295 191.650 102.465 191.790 ;
        RECT 101.140 191.610 102.105 191.620 ;
        RECT 100.800 191.440 100.970 191.530 ;
        RECT 101.430 191.450 102.105 191.610 ;
        RECT 98.840 191.250 99.580 191.280 ;
        RECT 98.840 190.950 99.755 191.250 ;
        RECT 99.430 190.775 99.755 190.950 ;
        RECT 98.460 190.220 98.715 190.750 ;
        RECT 98.885 190.040 99.190 190.500 ;
        RECT 99.435 190.420 99.755 190.775 ;
        RECT 99.925 190.990 100.465 191.360 ;
        RECT 100.800 191.270 101.205 191.440 ;
        RECT 99.925 190.590 100.165 190.990 ;
        RECT 100.645 190.820 100.865 191.100 ;
        RECT 100.335 190.650 100.865 190.820 ;
        RECT 100.335 190.420 100.505 190.650 ;
        RECT 101.035 190.490 101.205 191.270 ;
        RECT 101.375 190.660 101.725 191.280 ;
        RECT 101.895 190.660 102.105 191.450 ;
        RECT 102.295 191.480 103.795 191.650 ;
        RECT 102.295 190.790 102.465 191.480 ;
        RECT 104.155 191.310 104.325 192.090 ;
        RECT 105.130 191.960 105.300 192.090 ;
        RECT 102.635 191.140 104.325 191.310 ;
        RECT 104.495 191.530 104.960 191.920 ;
        RECT 105.130 191.790 105.525 191.960 ;
        RECT 102.635 190.960 102.805 191.140 ;
        RECT 99.435 190.250 100.505 190.420 ;
        RECT 100.675 190.040 100.865 190.480 ;
        RECT 101.035 190.210 101.985 190.490 ;
        RECT 102.295 190.400 102.555 190.790 ;
        RECT 102.975 190.720 103.765 190.970 ;
        RECT 102.205 190.230 102.555 190.400 ;
        RECT 102.765 190.040 103.095 190.500 ;
        RECT 103.970 190.430 104.140 191.140 ;
        RECT 104.495 190.940 104.665 191.530 ;
        RECT 104.310 190.720 104.665 190.940 ;
        RECT 104.835 190.720 105.185 191.340 ;
        RECT 105.355 190.430 105.525 191.790 ;
        RECT 105.890 191.620 106.215 192.405 ;
        RECT 105.695 190.570 106.155 191.620 ;
        RECT 103.970 190.260 104.825 190.430 ;
        RECT 105.030 190.260 105.525 190.430 ;
        RECT 105.695 190.040 106.025 190.400 ;
        RECT 106.385 190.300 106.555 192.420 ;
        RECT 106.725 192.090 107.055 192.590 ;
        RECT 107.225 191.920 107.480 192.420 ;
        RECT 106.730 191.750 107.480 191.920 ;
        RECT 106.730 190.760 106.960 191.750 ;
        RECT 107.130 190.930 107.480 191.580 ;
        RECT 107.655 191.500 109.325 192.590 ;
        RECT 109.585 191.660 109.755 192.420 ;
        RECT 109.935 191.830 110.265 192.590 ;
        RECT 107.655 190.980 108.405 191.500 ;
        RECT 109.585 191.490 110.250 191.660 ;
        RECT 110.435 191.515 110.705 192.420 ;
        RECT 110.080 191.345 110.250 191.490 ;
        RECT 108.575 190.810 109.325 191.330 ;
        RECT 109.515 190.940 109.845 191.310 ;
        RECT 110.080 191.015 110.365 191.345 ;
        RECT 106.730 190.590 107.480 190.760 ;
        RECT 106.725 190.040 107.055 190.420 ;
        RECT 107.225 190.300 107.480 190.590 ;
        RECT 107.655 190.040 109.325 190.810 ;
        RECT 110.080 190.760 110.250 191.015 ;
        RECT 109.585 190.590 110.250 190.760 ;
        RECT 110.535 190.715 110.705 191.515 ;
        RECT 110.875 191.500 114.385 192.590 ;
        RECT 114.555 191.500 115.765 192.590 ;
        RECT 110.875 190.980 112.565 191.500 ;
        RECT 112.735 190.810 114.385 191.330 ;
        RECT 114.555 190.960 115.075 191.500 ;
        RECT 109.585 190.210 109.755 190.590 ;
        RECT 109.935 190.040 110.265 190.420 ;
        RECT 110.445 190.210 110.705 190.715 ;
        RECT 110.875 190.040 114.385 190.810 ;
        RECT 115.245 190.790 115.765 191.330 ;
        RECT 114.555 190.040 115.765 190.790 ;
        RECT 10.510 189.870 115.850 190.040 ;
        RECT 10.595 189.120 11.805 189.870 ;
        RECT 12.900 189.325 18.245 189.870 ;
        RECT 18.420 189.325 23.765 189.870 ;
        RECT 10.595 188.580 11.115 189.120 ;
        RECT 11.285 188.410 11.805 188.950 ;
        RECT 10.595 187.320 11.805 188.410 ;
        RECT 14.490 187.755 14.840 189.005 ;
        RECT 16.320 188.495 16.660 189.325 ;
        RECT 20.010 187.755 20.360 189.005 ;
        RECT 21.840 188.495 22.180 189.325 ;
        RECT 23.975 189.050 24.205 189.870 ;
        RECT 24.375 189.070 24.705 189.700 ;
        RECT 23.955 188.630 24.285 188.880 ;
        RECT 24.455 188.470 24.705 189.070 ;
        RECT 24.875 189.050 25.085 189.870 ;
        RECT 25.315 189.145 25.605 189.870 ;
        RECT 26.970 189.060 27.215 189.665 ;
        RECT 27.435 189.335 27.945 189.870 ;
        RECT 26.695 188.890 27.925 189.060 ;
        RECT 12.900 187.320 18.245 187.755 ;
        RECT 18.420 187.320 23.765 187.755 ;
        RECT 23.975 187.320 24.205 188.460 ;
        RECT 24.375 187.490 24.705 188.470 ;
        RECT 24.875 187.320 25.085 188.460 ;
        RECT 25.315 187.320 25.605 188.485 ;
        RECT 26.695 188.080 27.035 188.890 ;
        RECT 27.205 188.325 27.955 188.515 ;
        RECT 26.695 187.670 27.210 188.080 ;
        RECT 27.445 187.320 27.615 188.080 ;
        RECT 27.785 187.660 27.955 188.325 ;
        RECT 28.125 188.340 28.315 189.700 ;
        RECT 28.485 188.850 28.760 189.700 ;
        RECT 28.950 189.335 29.480 189.700 ;
        RECT 29.905 189.470 30.235 189.870 ;
        RECT 29.305 189.300 29.480 189.335 ;
        RECT 28.485 188.680 28.765 188.850 ;
        RECT 28.485 188.540 28.760 188.680 ;
        RECT 28.965 188.340 29.135 189.140 ;
        RECT 28.125 188.170 29.135 188.340 ;
        RECT 29.305 189.130 30.235 189.300 ;
        RECT 30.405 189.130 30.660 189.700 ;
        RECT 29.305 188.000 29.475 189.130 ;
        RECT 30.065 188.960 30.235 189.130 ;
        RECT 28.350 187.830 29.475 188.000 ;
        RECT 29.645 188.630 29.840 188.960 ;
        RECT 30.065 188.630 30.320 188.960 ;
        RECT 29.645 187.660 29.815 188.630 ;
        RECT 30.490 188.460 30.660 189.130 ;
        RECT 31.335 189.050 31.565 189.870 ;
        RECT 31.735 189.070 32.065 189.700 ;
        RECT 31.315 188.630 31.645 188.880 ;
        RECT 31.815 188.470 32.065 189.070 ;
        RECT 32.235 189.050 32.445 189.870 ;
        RECT 32.675 189.130 33.060 189.700 ;
        RECT 33.230 189.410 33.555 189.870 ;
        RECT 34.075 189.240 34.355 189.700 ;
        RECT 27.785 187.490 29.815 187.660 ;
        RECT 29.985 187.320 30.155 188.460 ;
        RECT 30.325 187.490 30.660 188.460 ;
        RECT 31.335 187.320 31.565 188.460 ;
        RECT 31.735 187.490 32.065 188.470 ;
        RECT 32.675 188.460 32.955 189.130 ;
        RECT 33.230 189.070 34.355 189.240 ;
        RECT 33.230 188.960 33.680 189.070 ;
        RECT 33.125 188.630 33.680 188.960 ;
        RECT 34.545 188.900 34.945 189.700 ;
        RECT 35.345 189.410 35.615 189.870 ;
        RECT 35.785 189.240 36.070 189.700 ;
        RECT 32.235 187.320 32.445 188.460 ;
        RECT 32.675 187.490 33.060 188.460 ;
        RECT 33.230 188.170 33.680 188.630 ;
        RECT 33.850 188.340 34.945 188.900 ;
        RECT 33.230 187.950 34.355 188.170 ;
        RECT 33.230 187.320 33.555 187.780 ;
        RECT 34.075 187.490 34.355 187.950 ;
        RECT 34.545 187.490 34.945 188.340 ;
        RECT 35.115 189.070 36.070 189.240 ;
        RECT 36.360 189.130 36.615 189.700 ;
        RECT 36.785 189.470 37.115 189.870 ;
        RECT 37.540 189.335 38.070 189.700 ;
        RECT 37.540 189.300 37.715 189.335 ;
        RECT 36.785 189.130 37.715 189.300 ;
        RECT 35.115 188.170 35.325 189.070 ;
        RECT 35.495 188.340 36.185 188.900 ;
        RECT 36.360 188.460 36.530 189.130 ;
        RECT 36.785 188.960 36.955 189.130 ;
        RECT 36.700 188.630 36.955 188.960 ;
        RECT 37.180 188.630 37.375 188.960 ;
        RECT 35.115 187.950 36.070 188.170 ;
        RECT 35.345 187.320 35.615 187.780 ;
        RECT 35.785 187.490 36.070 187.950 ;
        RECT 36.360 187.490 36.695 188.460 ;
        RECT 36.865 187.320 37.035 188.460 ;
        RECT 37.205 187.660 37.375 188.630 ;
        RECT 37.545 188.000 37.715 189.130 ;
        RECT 37.885 188.340 38.055 189.140 ;
        RECT 38.260 188.850 38.535 189.700 ;
        RECT 38.255 188.680 38.535 188.850 ;
        RECT 38.260 188.540 38.535 188.680 ;
        RECT 38.705 188.340 38.895 189.700 ;
        RECT 39.075 189.335 39.585 189.870 ;
        RECT 39.805 189.060 40.050 189.665 ;
        RECT 40.500 189.160 40.755 189.690 ;
        RECT 40.925 189.410 41.230 189.870 ;
        RECT 41.475 189.490 42.545 189.660 ;
        RECT 39.095 188.890 40.325 189.060 ;
        RECT 37.885 188.170 38.895 188.340 ;
        RECT 39.065 188.325 39.815 188.515 ;
        RECT 37.545 187.830 38.670 188.000 ;
        RECT 39.065 187.660 39.235 188.325 ;
        RECT 39.985 188.080 40.325 188.890 ;
        RECT 37.205 187.490 39.235 187.660 ;
        RECT 39.405 187.320 39.575 188.080 ;
        RECT 39.810 187.670 40.325 188.080 ;
        RECT 40.500 188.510 40.710 189.160 ;
        RECT 41.475 189.135 41.795 189.490 ;
        RECT 41.470 188.960 41.795 189.135 ;
        RECT 40.880 188.660 41.795 188.960 ;
        RECT 41.965 188.920 42.205 189.320 ;
        RECT 42.375 189.260 42.545 189.490 ;
        RECT 42.715 189.430 42.905 189.870 ;
        RECT 43.075 189.420 44.025 189.700 ;
        RECT 44.245 189.510 44.595 189.680 ;
        RECT 42.375 189.090 42.905 189.260 ;
        RECT 40.880 188.630 41.620 188.660 ;
        RECT 40.500 187.630 40.755 188.510 ;
        RECT 40.925 187.320 41.230 188.460 ;
        RECT 41.450 188.040 41.620 188.630 ;
        RECT 41.965 188.550 42.505 188.920 ;
        RECT 42.685 188.810 42.905 189.090 ;
        RECT 43.075 188.640 43.245 189.420 ;
        RECT 42.840 188.470 43.245 188.640 ;
        RECT 43.415 188.630 43.765 189.250 ;
        RECT 42.840 188.380 43.010 188.470 ;
        RECT 43.935 188.460 44.145 189.250 ;
        RECT 41.790 188.210 43.010 188.380 ;
        RECT 43.470 188.300 44.145 188.460 ;
        RECT 41.450 187.870 42.250 188.040 ;
        RECT 41.570 187.320 41.900 187.700 ;
        RECT 42.080 187.580 42.250 187.870 ;
        RECT 42.840 187.830 43.010 188.210 ;
        RECT 43.180 188.290 44.145 188.300 ;
        RECT 44.335 189.120 44.595 189.510 ;
        RECT 44.805 189.410 45.135 189.870 ;
        RECT 46.010 189.480 46.865 189.650 ;
        RECT 47.070 189.480 47.565 189.650 ;
        RECT 47.735 189.510 48.065 189.870 ;
        RECT 44.335 188.430 44.505 189.120 ;
        RECT 44.675 188.770 44.845 188.950 ;
        RECT 45.015 188.940 45.805 189.190 ;
        RECT 46.010 188.770 46.180 189.480 ;
        RECT 46.350 188.970 46.705 189.190 ;
        RECT 44.675 188.600 46.365 188.770 ;
        RECT 43.180 188.000 43.640 188.290 ;
        RECT 44.335 188.260 45.835 188.430 ;
        RECT 44.335 188.120 44.505 188.260 ;
        RECT 43.945 187.950 44.505 188.120 ;
        RECT 42.420 187.320 42.670 187.780 ;
        RECT 42.840 187.490 43.710 187.830 ;
        RECT 43.945 187.490 44.115 187.950 ;
        RECT 44.950 187.920 46.025 188.090 ;
        RECT 44.285 187.320 44.655 187.780 ;
        RECT 44.950 187.580 45.120 187.920 ;
        RECT 45.290 187.320 45.620 187.750 ;
        RECT 45.855 187.580 46.025 187.920 ;
        RECT 46.195 187.820 46.365 188.600 ;
        RECT 46.535 188.380 46.705 188.970 ;
        RECT 46.875 188.570 47.225 189.190 ;
        RECT 46.535 187.990 47.000 188.380 ;
        RECT 47.395 188.120 47.565 189.480 ;
        RECT 47.735 188.290 48.195 189.340 ;
        RECT 47.170 187.950 47.565 188.120 ;
        RECT 47.170 187.820 47.340 187.950 ;
        RECT 46.195 187.490 46.875 187.820 ;
        RECT 47.090 187.490 47.340 187.820 ;
        RECT 47.510 187.320 47.760 187.780 ;
        RECT 47.930 187.505 48.255 188.290 ;
        RECT 48.425 187.490 48.595 189.610 ;
        RECT 48.765 189.490 49.095 189.870 ;
        RECT 49.265 189.320 49.520 189.610 ;
        RECT 48.770 189.150 49.520 189.320 ;
        RECT 49.695 189.195 49.955 189.700 ;
        RECT 50.135 189.490 50.465 189.870 ;
        RECT 50.645 189.320 50.815 189.700 ;
        RECT 48.770 188.160 49.000 189.150 ;
        RECT 49.170 188.330 49.520 188.980 ;
        RECT 49.695 188.395 49.865 189.195 ;
        RECT 50.150 189.150 50.815 189.320 ;
        RECT 50.150 188.895 50.320 189.150 ;
        RECT 51.075 189.145 51.365 189.870 ;
        RECT 51.995 189.100 54.585 189.870 ;
        RECT 54.845 189.320 55.015 189.700 ;
        RECT 55.195 189.490 55.525 189.870 ;
        RECT 54.845 189.150 55.510 189.320 ;
        RECT 55.705 189.195 55.965 189.700 ;
        RECT 50.035 188.565 50.320 188.895 ;
        RECT 50.555 188.600 50.885 188.970 ;
        RECT 50.150 188.420 50.320 188.565 ;
        RECT 48.770 187.990 49.520 188.160 ;
        RECT 48.765 187.320 49.095 187.820 ;
        RECT 49.265 187.490 49.520 187.990 ;
        RECT 49.695 187.490 49.965 188.395 ;
        RECT 50.150 188.250 50.815 188.420 ;
        RECT 50.135 187.320 50.465 188.080 ;
        RECT 50.645 187.490 50.815 188.250 ;
        RECT 51.075 187.320 51.365 188.485 ;
        RECT 51.995 188.410 53.205 188.930 ;
        RECT 53.375 188.580 54.585 189.100 ;
        RECT 54.775 188.600 55.105 188.970 ;
        RECT 55.340 188.895 55.510 189.150 ;
        RECT 55.340 188.565 55.625 188.895 ;
        RECT 55.340 188.420 55.510 188.565 ;
        RECT 51.995 187.320 54.585 188.410 ;
        RECT 54.845 188.250 55.510 188.420 ;
        RECT 55.795 188.395 55.965 189.195 ;
        RECT 56.135 189.120 57.345 189.870 ;
        RECT 54.845 187.490 55.015 188.250 ;
        RECT 55.195 187.320 55.525 188.080 ;
        RECT 55.695 187.490 55.965 188.395 ;
        RECT 56.135 188.410 56.655 188.950 ;
        RECT 56.825 188.580 57.345 189.120 ;
        RECT 57.515 189.100 61.025 189.870 ;
        RECT 61.200 189.325 66.545 189.870 ;
        RECT 66.715 189.370 66.975 189.700 ;
        RECT 67.185 189.390 67.460 189.870 ;
        RECT 57.515 188.410 59.205 188.930 ;
        RECT 59.375 188.580 61.025 189.100 ;
        RECT 56.135 187.320 57.345 188.410 ;
        RECT 57.515 187.320 61.025 188.410 ;
        RECT 62.790 187.755 63.140 189.005 ;
        RECT 64.620 188.495 64.960 189.325 ;
        RECT 66.715 188.460 66.885 189.370 ;
        RECT 67.670 189.300 67.875 189.700 ;
        RECT 68.045 189.470 68.380 189.870 ;
        RECT 67.055 188.630 67.415 189.210 ;
        RECT 67.670 189.130 68.355 189.300 ;
        RECT 67.595 188.460 67.845 188.960 ;
        RECT 66.715 188.290 67.845 188.460 ;
        RECT 61.200 187.320 66.545 187.755 ;
        RECT 66.715 187.520 66.985 188.290 ;
        RECT 68.015 188.100 68.355 189.130 ;
        RECT 68.555 189.120 69.765 189.870 ;
        RECT 67.155 187.320 67.485 188.100 ;
        RECT 67.690 187.925 68.355 188.100 ;
        RECT 68.555 188.410 69.075 188.950 ;
        RECT 69.245 188.580 69.765 189.120 ;
        RECT 69.935 189.370 70.195 189.700 ;
        RECT 70.405 189.390 70.680 189.870 ;
        RECT 69.935 188.460 70.105 189.370 ;
        RECT 70.890 189.300 71.095 189.700 ;
        RECT 71.265 189.470 71.600 189.870 ;
        RECT 70.275 188.630 70.635 189.210 ;
        RECT 70.890 189.130 71.575 189.300 ;
        RECT 70.815 188.460 71.065 188.960 ;
        RECT 67.690 187.520 67.875 187.925 ;
        RECT 68.045 187.320 68.380 187.745 ;
        RECT 68.555 187.320 69.765 188.410 ;
        RECT 69.935 188.290 71.065 188.460 ;
        RECT 69.935 187.520 70.205 188.290 ;
        RECT 71.235 188.100 71.575 189.130 ;
        RECT 72.970 189.060 73.215 189.665 ;
        RECT 73.435 189.335 73.945 189.870 ;
        RECT 70.375 187.320 70.705 188.100 ;
        RECT 70.910 187.925 71.575 188.100 ;
        RECT 72.695 188.890 73.925 189.060 ;
        RECT 72.695 188.080 73.035 188.890 ;
        RECT 73.205 188.325 73.955 188.515 ;
        RECT 70.910 187.520 71.095 187.925 ;
        RECT 71.265 187.320 71.600 187.745 ;
        RECT 72.695 187.670 73.210 188.080 ;
        RECT 73.445 187.320 73.615 188.080 ;
        RECT 73.785 187.660 73.955 188.325 ;
        RECT 74.125 188.340 74.315 189.700 ;
        RECT 74.485 189.190 74.760 189.700 ;
        RECT 74.950 189.335 75.480 189.700 ;
        RECT 75.905 189.470 76.235 189.870 ;
        RECT 75.305 189.300 75.480 189.335 ;
        RECT 74.485 189.020 74.765 189.190 ;
        RECT 74.485 188.540 74.760 189.020 ;
        RECT 74.965 188.340 75.135 189.140 ;
        RECT 74.125 188.170 75.135 188.340 ;
        RECT 75.305 189.130 76.235 189.300 ;
        RECT 76.405 189.130 76.660 189.700 ;
        RECT 76.835 189.145 77.125 189.870 ;
        RECT 77.670 189.160 77.925 189.690 ;
        RECT 78.105 189.410 78.390 189.870 ;
        RECT 75.305 188.000 75.475 189.130 ;
        RECT 76.065 188.960 76.235 189.130 ;
        RECT 74.350 187.830 75.475 188.000 ;
        RECT 75.645 188.630 75.840 188.960 ;
        RECT 76.065 188.630 76.320 188.960 ;
        RECT 75.645 187.660 75.815 188.630 ;
        RECT 76.490 188.460 76.660 189.130 ;
        RECT 73.785 187.490 75.815 187.660 ;
        RECT 75.985 187.320 76.155 188.460 ;
        RECT 76.325 187.490 76.660 188.460 ;
        RECT 76.835 187.320 77.125 188.485 ;
        RECT 77.670 188.300 77.850 189.160 ;
        RECT 78.570 188.960 78.820 189.610 ;
        RECT 78.020 188.630 78.820 188.960 ;
        RECT 77.670 187.830 77.925 188.300 ;
        RECT 77.585 187.660 77.925 187.830 ;
        RECT 77.670 187.630 77.925 187.660 ;
        RECT 78.105 187.320 78.390 188.120 ;
        RECT 78.570 188.040 78.820 188.630 ;
        RECT 79.020 189.275 79.340 189.605 ;
        RECT 79.520 189.390 80.180 189.870 ;
        RECT 80.380 189.480 81.230 189.650 ;
        RECT 79.020 188.380 79.210 189.275 ;
        RECT 79.530 188.950 80.190 189.220 ;
        RECT 79.860 188.890 80.190 188.950 ;
        RECT 79.380 188.720 79.710 188.780 ;
        RECT 80.380 188.720 80.550 189.480 ;
        RECT 81.790 189.410 82.110 189.870 ;
        RECT 82.310 189.230 82.560 189.660 ;
        RECT 82.850 189.430 83.260 189.870 ;
        RECT 83.430 189.490 84.445 189.690 ;
        RECT 80.720 189.060 81.970 189.230 ;
        RECT 80.720 188.940 81.050 189.060 ;
        RECT 79.380 188.550 81.280 188.720 ;
        RECT 79.020 188.210 80.940 188.380 ;
        RECT 79.020 188.190 79.340 188.210 ;
        RECT 78.570 187.530 78.900 188.040 ;
        RECT 79.170 187.580 79.340 188.190 ;
        RECT 81.110 188.040 81.280 188.550 ;
        RECT 81.450 188.480 81.630 188.890 ;
        RECT 81.800 188.300 81.970 189.060 ;
        RECT 79.510 187.320 79.840 188.010 ;
        RECT 80.070 187.870 81.280 188.040 ;
        RECT 81.450 187.990 81.970 188.300 ;
        RECT 82.140 188.890 82.560 189.230 ;
        RECT 82.850 188.890 83.260 189.220 ;
        RECT 82.140 188.120 82.330 188.890 ;
        RECT 83.430 188.760 83.600 189.490 ;
        RECT 84.745 189.320 84.915 189.650 ;
        RECT 85.085 189.490 85.415 189.870 ;
        RECT 83.770 188.940 84.120 189.310 ;
        RECT 83.430 188.720 83.850 188.760 ;
        RECT 82.500 188.550 83.850 188.720 ;
        RECT 82.500 188.390 82.750 188.550 ;
        RECT 83.260 188.120 83.510 188.380 ;
        RECT 82.140 187.870 83.510 188.120 ;
        RECT 80.070 187.580 80.310 187.870 ;
        RECT 81.110 187.790 81.280 187.870 ;
        RECT 80.510 187.320 80.930 187.700 ;
        RECT 81.110 187.540 81.740 187.790 ;
        RECT 82.210 187.320 82.540 187.700 ;
        RECT 82.710 187.580 82.880 187.870 ;
        RECT 83.680 187.705 83.850 188.550 ;
        RECT 84.300 188.380 84.520 189.250 ;
        RECT 84.745 189.130 85.440 189.320 ;
        RECT 84.020 188.000 84.520 188.380 ;
        RECT 84.690 188.330 85.100 188.950 ;
        RECT 85.270 188.160 85.440 189.130 ;
        RECT 84.745 187.990 85.440 188.160 ;
        RECT 83.060 187.320 83.440 187.700 ;
        RECT 83.680 187.535 84.510 187.705 ;
        RECT 84.745 187.490 84.915 187.990 ;
        RECT 85.085 187.320 85.415 187.820 ;
        RECT 85.630 187.490 85.855 189.610 ;
        RECT 86.025 189.490 86.355 189.870 ;
        RECT 86.525 189.320 86.695 189.610 ;
        RECT 86.030 189.150 86.695 189.320 ;
        RECT 86.030 188.160 86.260 189.150 ;
        RECT 86.955 189.120 88.165 189.870 ;
        RECT 86.430 188.330 86.780 188.980 ;
        RECT 86.955 188.410 87.475 188.950 ;
        RECT 87.645 188.580 88.165 189.120 ;
        RECT 88.610 189.060 88.855 189.665 ;
        RECT 89.075 189.335 89.585 189.870 ;
        RECT 88.335 188.890 89.565 189.060 ;
        RECT 86.030 187.990 86.695 188.160 ;
        RECT 86.025 187.320 86.355 187.820 ;
        RECT 86.525 187.490 86.695 187.990 ;
        RECT 86.955 187.320 88.165 188.410 ;
        RECT 88.335 188.080 88.675 188.890 ;
        RECT 88.845 188.325 89.595 188.515 ;
        RECT 88.335 187.670 88.850 188.080 ;
        RECT 89.085 187.320 89.255 188.080 ;
        RECT 89.425 187.660 89.595 188.325 ;
        RECT 89.765 188.340 89.955 189.700 ;
        RECT 90.125 188.850 90.400 189.700 ;
        RECT 90.590 189.335 91.120 189.700 ;
        RECT 91.545 189.470 91.875 189.870 ;
        RECT 90.945 189.300 91.120 189.335 ;
        RECT 90.125 188.680 90.405 188.850 ;
        RECT 90.125 188.540 90.400 188.680 ;
        RECT 90.605 188.340 90.775 189.140 ;
        RECT 89.765 188.170 90.775 188.340 ;
        RECT 90.945 189.130 91.875 189.300 ;
        RECT 92.045 189.130 92.300 189.700 ;
        RECT 90.945 188.000 91.115 189.130 ;
        RECT 91.705 188.960 91.875 189.130 ;
        RECT 89.990 187.830 91.115 188.000 ;
        RECT 91.285 188.630 91.480 188.960 ;
        RECT 91.705 188.630 91.960 188.960 ;
        RECT 91.285 187.660 91.455 188.630 ;
        RECT 92.130 188.460 92.300 189.130 ;
        RECT 89.425 187.490 91.455 187.660 ;
        RECT 91.625 187.320 91.795 188.460 ;
        RECT 91.965 187.490 92.300 188.460 ;
        RECT 92.475 189.195 92.735 189.700 ;
        RECT 92.915 189.490 93.245 189.870 ;
        RECT 93.425 189.320 93.595 189.700 ;
        RECT 92.475 188.395 92.645 189.195 ;
        RECT 92.930 189.150 93.595 189.320 ;
        RECT 94.890 189.240 95.175 189.700 ;
        RECT 95.345 189.410 95.615 189.870 ;
        RECT 92.930 188.895 93.100 189.150 ;
        RECT 94.890 189.070 95.845 189.240 ;
        RECT 92.815 188.565 93.100 188.895 ;
        RECT 93.335 188.600 93.665 188.970 ;
        RECT 92.930 188.420 93.100 188.565 ;
        RECT 92.475 187.490 92.745 188.395 ;
        RECT 92.930 188.250 93.595 188.420 ;
        RECT 94.775 188.340 95.465 188.900 ;
        RECT 92.915 187.320 93.245 188.080 ;
        RECT 93.425 187.490 93.595 188.250 ;
        RECT 95.635 188.170 95.845 189.070 ;
        RECT 94.890 187.950 95.845 188.170 ;
        RECT 96.015 188.900 96.415 189.700 ;
        RECT 96.605 189.240 96.885 189.700 ;
        RECT 97.405 189.410 97.730 189.870 ;
        RECT 96.605 189.070 97.730 189.240 ;
        RECT 97.900 189.130 98.285 189.700 ;
        RECT 97.280 188.960 97.730 189.070 ;
        RECT 96.015 188.340 97.110 188.900 ;
        RECT 97.280 188.630 97.835 188.960 ;
        RECT 94.890 187.490 95.175 187.950 ;
        RECT 95.345 187.320 95.615 187.780 ;
        RECT 96.015 187.490 96.415 188.340 ;
        RECT 97.280 188.170 97.730 188.630 ;
        RECT 98.005 188.460 98.285 189.130 ;
        RECT 98.730 189.060 98.975 189.665 ;
        RECT 99.195 189.335 99.705 189.870 ;
        RECT 96.605 187.950 97.730 188.170 ;
        RECT 96.605 187.490 96.885 187.950 ;
        RECT 97.405 187.320 97.730 187.780 ;
        RECT 97.900 187.490 98.285 188.460 ;
        RECT 98.455 188.890 99.685 189.060 ;
        RECT 98.455 188.080 98.795 188.890 ;
        RECT 98.965 188.325 99.715 188.515 ;
        RECT 98.455 187.670 98.970 188.080 ;
        RECT 99.205 187.320 99.375 188.080 ;
        RECT 99.545 187.660 99.715 188.325 ;
        RECT 99.885 188.340 100.075 189.700 ;
        RECT 100.245 189.190 100.520 189.700 ;
        RECT 100.710 189.335 101.240 189.700 ;
        RECT 101.665 189.470 101.995 189.870 ;
        RECT 101.065 189.300 101.240 189.335 ;
        RECT 100.245 189.020 100.525 189.190 ;
        RECT 100.245 188.540 100.520 189.020 ;
        RECT 100.725 188.340 100.895 189.140 ;
        RECT 99.885 188.170 100.895 188.340 ;
        RECT 101.065 189.130 101.995 189.300 ;
        RECT 102.165 189.130 102.420 189.700 ;
        RECT 102.595 189.145 102.885 189.870 ;
        RECT 101.065 188.000 101.235 189.130 ;
        RECT 101.825 188.960 101.995 189.130 ;
        RECT 100.110 187.830 101.235 188.000 ;
        RECT 101.405 188.630 101.600 188.960 ;
        RECT 101.825 188.630 102.080 188.960 ;
        RECT 101.405 187.660 101.575 188.630 ;
        RECT 102.250 188.460 102.420 189.130 ;
        RECT 103.555 189.050 103.785 189.870 ;
        RECT 103.955 189.070 104.285 189.700 ;
        RECT 103.535 188.630 103.865 188.880 ;
        RECT 99.545 187.490 101.575 187.660 ;
        RECT 101.745 187.320 101.915 188.460 ;
        RECT 102.085 187.490 102.420 188.460 ;
        RECT 102.595 187.320 102.885 188.485 ;
        RECT 104.035 188.470 104.285 189.070 ;
        RECT 104.455 189.050 104.665 189.870 ;
        RECT 104.900 189.160 105.155 189.690 ;
        RECT 105.325 189.410 105.630 189.870 ;
        RECT 105.875 189.490 106.945 189.660 ;
        RECT 103.555 187.320 103.785 188.460 ;
        RECT 103.955 187.490 104.285 188.470 ;
        RECT 104.900 188.510 105.110 189.160 ;
        RECT 105.875 189.135 106.195 189.490 ;
        RECT 105.870 188.960 106.195 189.135 ;
        RECT 105.280 188.660 106.195 188.960 ;
        RECT 106.365 188.920 106.605 189.320 ;
        RECT 106.775 189.260 106.945 189.490 ;
        RECT 107.115 189.430 107.305 189.870 ;
        RECT 107.475 189.420 108.425 189.700 ;
        RECT 108.645 189.510 108.995 189.680 ;
        RECT 106.775 189.090 107.305 189.260 ;
        RECT 105.280 188.630 106.020 188.660 ;
        RECT 104.455 187.320 104.665 188.460 ;
        RECT 104.900 187.630 105.155 188.510 ;
        RECT 105.325 187.320 105.630 188.460 ;
        RECT 105.850 188.040 106.020 188.630 ;
        RECT 106.365 188.550 106.905 188.920 ;
        RECT 107.085 188.810 107.305 189.090 ;
        RECT 107.475 188.640 107.645 189.420 ;
        RECT 107.240 188.470 107.645 188.640 ;
        RECT 107.815 188.630 108.165 189.250 ;
        RECT 107.240 188.380 107.410 188.470 ;
        RECT 108.335 188.460 108.545 189.250 ;
        RECT 106.190 188.210 107.410 188.380 ;
        RECT 107.870 188.300 108.545 188.460 ;
        RECT 105.850 187.870 106.650 188.040 ;
        RECT 105.970 187.320 106.300 187.700 ;
        RECT 106.480 187.580 106.650 187.870 ;
        RECT 107.240 187.830 107.410 188.210 ;
        RECT 107.580 188.290 108.545 188.300 ;
        RECT 108.735 189.120 108.995 189.510 ;
        RECT 109.205 189.410 109.535 189.870 ;
        RECT 110.410 189.480 111.265 189.650 ;
        RECT 111.470 189.480 111.965 189.650 ;
        RECT 112.135 189.510 112.465 189.870 ;
        RECT 108.735 188.430 108.905 189.120 ;
        RECT 109.075 188.770 109.245 188.950 ;
        RECT 109.415 188.940 110.205 189.190 ;
        RECT 110.410 188.770 110.580 189.480 ;
        RECT 110.750 188.970 111.105 189.190 ;
        RECT 109.075 188.600 110.765 188.770 ;
        RECT 107.580 188.000 108.040 188.290 ;
        RECT 108.735 188.260 110.235 188.430 ;
        RECT 108.735 188.120 108.905 188.260 ;
        RECT 108.345 187.950 108.905 188.120 ;
        RECT 106.820 187.320 107.070 187.780 ;
        RECT 107.240 187.490 108.110 187.830 ;
        RECT 108.345 187.490 108.515 187.950 ;
        RECT 109.350 187.920 110.425 188.090 ;
        RECT 108.685 187.320 109.055 187.780 ;
        RECT 109.350 187.580 109.520 187.920 ;
        RECT 109.690 187.320 110.020 187.750 ;
        RECT 110.255 187.580 110.425 187.920 ;
        RECT 110.595 187.820 110.765 188.600 ;
        RECT 110.935 188.380 111.105 188.970 ;
        RECT 111.275 188.570 111.625 189.190 ;
        RECT 110.935 187.990 111.400 188.380 ;
        RECT 111.795 188.120 111.965 189.480 ;
        RECT 112.135 188.290 112.595 189.340 ;
        RECT 111.570 187.950 111.965 188.120 ;
        RECT 111.570 187.820 111.740 187.950 ;
        RECT 110.595 187.490 111.275 187.820 ;
        RECT 111.490 187.490 111.740 187.820 ;
        RECT 111.910 187.320 112.160 187.780 ;
        RECT 112.330 187.505 112.655 188.290 ;
        RECT 112.825 187.490 112.995 189.610 ;
        RECT 113.165 189.490 113.495 189.870 ;
        RECT 113.665 189.320 113.920 189.610 ;
        RECT 113.170 189.150 113.920 189.320 ;
        RECT 113.170 188.160 113.400 189.150 ;
        RECT 114.555 189.120 115.765 189.870 ;
        RECT 113.570 188.330 113.920 188.980 ;
        RECT 114.555 188.410 115.075 188.950 ;
        RECT 115.245 188.580 115.765 189.120 ;
        RECT 113.170 187.990 113.920 188.160 ;
        RECT 113.165 187.320 113.495 187.820 ;
        RECT 113.665 187.490 113.920 187.990 ;
        RECT 114.555 187.320 115.765 188.410 ;
        RECT 10.510 187.150 115.850 187.320 ;
        RECT 10.595 186.060 11.805 187.150 ;
        RECT 10.595 185.350 11.115 185.890 ;
        RECT 11.285 185.520 11.805 186.060 ;
        RECT 12.435 185.985 12.725 187.150 ;
        RECT 12.895 186.060 14.105 187.150 ;
        RECT 14.280 186.715 19.625 187.150 ;
        RECT 12.895 185.520 13.415 186.060 ;
        RECT 13.585 185.350 14.105 185.890 ;
        RECT 15.870 185.465 16.220 186.715 ;
        RECT 10.595 184.600 11.805 185.350 ;
        RECT 12.435 184.600 12.725 185.325 ;
        RECT 12.895 184.600 14.105 185.350 ;
        RECT 17.700 185.145 18.040 185.975 ;
        RECT 19.800 185.960 20.055 186.840 ;
        RECT 20.225 186.010 20.530 187.150 ;
        RECT 20.870 186.770 21.200 187.150 ;
        RECT 21.380 186.600 21.550 186.890 ;
        RECT 21.720 186.690 21.970 187.150 ;
        RECT 20.750 186.430 21.550 186.600 ;
        RECT 22.140 186.640 23.010 186.980 ;
        RECT 19.800 185.310 20.010 185.960 ;
        RECT 20.750 185.840 20.920 186.430 ;
        RECT 22.140 186.260 22.310 186.640 ;
        RECT 23.245 186.520 23.415 186.980 ;
        RECT 23.585 186.690 23.955 187.150 ;
        RECT 24.250 186.550 24.420 186.890 ;
        RECT 24.590 186.720 24.920 187.150 ;
        RECT 25.155 186.550 25.325 186.890 ;
        RECT 21.090 186.090 22.310 186.260 ;
        RECT 22.480 186.180 22.940 186.470 ;
        RECT 23.245 186.350 23.805 186.520 ;
        RECT 24.250 186.380 25.325 186.550 ;
        RECT 25.495 186.650 26.175 186.980 ;
        RECT 26.390 186.650 26.640 186.980 ;
        RECT 26.810 186.690 27.060 187.150 ;
        RECT 23.635 186.210 23.805 186.350 ;
        RECT 22.480 186.170 23.445 186.180 ;
        RECT 22.140 186.000 22.310 186.090 ;
        RECT 22.770 186.010 23.445 186.170 ;
        RECT 20.180 185.810 20.920 185.840 ;
        RECT 20.180 185.510 21.095 185.810 ;
        RECT 20.770 185.335 21.095 185.510 ;
        RECT 14.280 184.600 19.625 185.145 ;
        RECT 19.800 184.780 20.055 185.310 ;
        RECT 20.225 184.600 20.530 185.060 ;
        RECT 20.775 184.980 21.095 185.335 ;
        RECT 21.265 185.550 21.805 185.920 ;
        RECT 22.140 185.830 22.545 186.000 ;
        RECT 21.265 185.150 21.505 185.550 ;
        RECT 21.985 185.380 22.205 185.660 ;
        RECT 21.675 185.210 22.205 185.380 ;
        RECT 21.675 184.980 21.845 185.210 ;
        RECT 22.375 185.050 22.545 185.830 ;
        RECT 22.715 185.220 23.065 185.840 ;
        RECT 23.235 185.220 23.445 186.010 ;
        RECT 23.635 186.040 25.135 186.210 ;
        RECT 23.635 185.350 23.805 186.040 ;
        RECT 25.495 185.870 25.665 186.650 ;
        RECT 26.470 186.520 26.640 186.650 ;
        RECT 23.975 185.700 25.665 185.870 ;
        RECT 25.835 186.090 26.300 186.480 ;
        RECT 26.470 186.350 26.865 186.520 ;
        RECT 23.975 185.520 24.145 185.700 ;
        RECT 20.775 184.810 21.845 184.980 ;
        RECT 22.015 184.600 22.205 185.040 ;
        RECT 22.375 184.770 23.325 185.050 ;
        RECT 23.635 184.960 23.895 185.350 ;
        RECT 24.315 185.280 25.105 185.530 ;
        RECT 23.545 184.790 23.895 184.960 ;
        RECT 24.105 184.600 24.435 185.060 ;
        RECT 25.310 184.990 25.480 185.700 ;
        RECT 25.835 185.500 26.005 186.090 ;
        RECT 25.650 185.280 26.005 185.500 ;
        RECT 26.175 185.280 26.525 185.900 ;
        RECT 26.695 184.990 26.865 186.350 ;
        RECT 27.230 186.180 27.555 186.965 ;
        RECT 27.035 185.130 27.495 186.180 ;
        RECT 25.310 184.820 26.165 184.990 ;
        RECT 26.370 184.820 26.865 184.990 ;
        RECT 27.035 184.600 27.365 184.960 ;
        RECT 27.725 184.860 27.895 186.980 ;
        RECT 28.065 186.650 28.395 187.150 ;
        RECT 28.565 186.480 28.820 186.980 ;
        RECT 28.070 186.310 28.820 186.480 ;
        RECT 28.070 185.320 28.300 186.310 ;
        RECT 28.470 185.490 28.820 186.140 ;
        RECT 29.000 185.960 29.255 186.840 ;
        RECT 29.425 186.010 29.730 187.150 ;
        RECT 30.070 186.770 30.400 187.150 ;
        RECT 30.580 186.600 30.750 186.890 ;
        RECT 30.920 186.690 31.170 187.150 ;
        RECT 29.950 186.430 30.750 186.600 ;
        RECT 31.340 186.640 32.210 186.980 ;
        RECT 28.070 185.150 28.820 185.320 ;
        RECT 28.065 184.600 28.395 184.980 ;
        RECT 28.565 184.860 28.820 185.150 ;
        RECT 29.000 185.310 29.210 185.960 ;
        RECT 29.950 185.840 30.120 186.430 ;
        RECT 31.340 186.260 31.510 186.640 ;
        RECT 32.445 186.520 32.615 186.980 ;
        RECT 32.785 186.690 33.155 187.150 ;
        RECT 33.450 186.550 33.620 186.890 ;
        RECT 33.790 186.720 34.120 187.150 ;
        RECT 34.355 186.550 34.525 186.890 ;
        RECT 30.290 186.090 31.510 186.260 ;
        RECT 31.680 186.180 32.140 186.470 ;
        RECT 32.445 186.350 33.005 186.520 ;
        RECT 33.450 186.380 34.525 186.550 ;
        RECT 34.695 186.650 35.375 186.980 ;
        RECT 35.590 186.650 35.840 186.980 ;
        RECT 36.010 186.690 36.260 187.150 ;
        RECT 32.835 186.210 33.005 186.350 ;
        RECT 31.680 186.170 32.645 186.180 ;
        RECT 31.340 186.000 31.510 186.090 ;
        RECT 31.970 186.010 32.645 186.170 ;
        RECT 29.380 185.810 30.120 185.840 ;
        RECT 29.380 185.510 30.295 185.810 ;
        RECT 29.970 185.335 30.295 185.510 ;
        RECT 29.000 184.780 29.255 185.310 ;
        RECT 29.425 184.600 29.730 185.060 ;
        RECT 29.975 184.980 30.295 185.335 ;
        RECT 30.465 185.550 31.005 185.920 ;
        RECT 31.340 185.830 31.745 186.000 ;
        RECT 30.465 185.150 30.705 185.550 ;
        RECT 31.185 185.380 31.405 185.660 ;
        RECT 30.875 185.210 31.405 185.380 ;
        RECT 30.875 184.980 31.045 185.210 ;
        RECT 31.575 185.050 31.745 185.830 ;
        RECT 31.915 185.220 32.265 185.840 ;
        RECT 32.435 185.220 32.645 186.010 ;
        RECT 32.835 186.040 34.335 186.210 ;
        RECT 32.835 185.350 33.005 186.040 ;
        RECT 34.695 185.870 34.865 186.650 ;
        RECT 35.670 186.520 35.840 186.650 ;
        RECT 33.175 185.700 34.865 185.870 ;
        RECT 35.035 186.090 35.500 186.480 ;
        RECT 35.670 186.350 36.065 186.520 ;
        RECT 33.175 185.520 33.345 185.700 ;
        RECT 29.975 184.810 31.045 184.980 ;
        RECT 31.215 184.600 31.405 185.040 ;
        RECT 31.575 184.770 32.525 185.050 ;
        RECT 32.835 184.960 33.095 185.350 ;
        RECT 33.515 185.280 34.305 185.530 ;
        RECT 32.745 184.790 33.095 184.960 ;
        RECT 33.305 184.600 33.635 185.060 ;
        RECT 34.510 184.990 34.680 185.700 ;
        RECT 35.035 185.500 35.205 186.090 ;
        RECT 34.850 185.280 35.205 185.500 ;
        RECT 35.375 185.280 35.725 185.900 ;
        RECT 35.895 184.990 36.065 186.350 ;
        RECT 36.430 186.180 36.755 186.965 ;
        RECT 36.235 185.130 36.695 186.180 ;
        RECT 34.510 184.820 35.365 184.990 ;
        RECT 35.570 184.820 36.065 184.990 ;
        RECT 36.235 184.600 36.565 184.960 ;
        RECT 36.925 184.860 37.095 186.980 ;
        RECT 37.265 186.650 37.595 187.150 ;
        RECT 37.765 186.480 38.020 186.980 ;
        RECT 37.270 186.310 38.020 186.480 ;
        RECT 37.270 185.320 37.500 186.310 ;
        RECT 37.670 185.490 38.020 186.140 ;
        RECT 38.195 185.985 38.485 187.150 ;
        RECT 39.120 185.960 39.375 186.840 ;
        RECT 39.545 186.010 39.850 187.150 ;
        RECT 40.190 186.770 40.520 187.150 ;
        RECT 40.700 186.600 40.870 186.890 ;
        RECT 41.040 186.690 41.290 187.150 ;
        RECT 40.070 186.430 40.870 186.600 ;
        RECT 41.460 186.640 42.330 186.980 ;
        RECT 37.270 185.150 38.020 185.320 ;
        RECT 37.265 184.600 37.595 184.980 ;
        RECT 37.765 184.860 38.020 185.150 ;
        RECT 38.195 184.600 38.485 185.325 ;
        RECT 39.120 185.310 39.330 185.960 ;
        RECT 40.070 185.840 40.240 186.430 ;
        RECT 41.460 186.260 41.630 186.640 ;
        RECT 42.565 186.520 42.735 186.980 ;
        RECT 42.905 186.690 43.275 187.150 ;
        RECT 43.570 186.550 43.740 186.890 ;
        RECT 43.910 186.720 44.240 187.150 ;
        RECT 44.475 186.550 44.645 186.890 ;
        RECT 40.410 186.090 41.630 186.260 ;
        RECT 41.800 186.180 42.260 186.470 ;
        RECT 42.565 186.350 43.125 186.520 ;
        RECT 43.570 186.380 44.645 186.550 ;
        RECT 44.815 186.650 45.495 186.980 ;
        RECT 45.710 186.650 45.960 186.980 ;
        RECT 46.130 186.690 46.380 187.150 ;
        RECT 42.955 186.210 43.125 186.350 ;
        RECT 41.800 186.170 42.765 186.180 ;
        RECT 41.460 186.000 41.630 186.090 ;
        RECT 42.090 186.010 42.765 186.170 ;
        RECT 39.500 185.810 40.240 185.840 ;
        RECT 39.500 185.510 40.415 185.810 ;
        RECT 40.090 185.335 40.415 185.510 ;
        RECT 39.120 184.780 39.375 185.310 ;
        RECT 39.545 184.600 39.850 185.060 ;
        RECT 40.095 184.980 40.415 185.335 ;
        RECT 40.585 185.550 41.125 185.920 ;
        RECT 41.460 185.830 41.865 186.000 ;
        RECT 40.585 185.150 40.825 185.550 ;
        RECT 41.305 185.380 41.525 185.660 ;
        RECT 40.995 185.210 41.525 185.380 ;
        RECT 40.995 184.980 41.165 185.210 ;
        RECT 41.695 185.050 41.865 185.830 ;
        RECT 42.035 185.220 42.385 185.840 ;
        RECT 42.555 185.220 42.765 186.010 ;
        RECT 42.955 186.040 44.455 186.210 ;
        RECT 42.955 185.350 43.125 186.040 ;
        RECT 44.815 185.870 44.985 186.650 ;
        RECT 45.790 186.520 45.960 186.650 ;
        RECT 43.295 185.700 44.985 185.870 ;
        RECT 45.155 186.090 45.620 186.480 ;
        RECT 45.790 186.350 46.185 186.520 ;
        RECT 43.295 185.520 43.465 185.700 ;
        RECT 40.095 184.810 41.165 184.980 ;
        RECT 41.335 184.600 41.525 185.040 ;
        RECT 41.695 184.770 42.645 185.050 ;
        RECT 42.955 184.960 43.215 185.350 ;
        RECT 43.635 185.280 44.425 185.530 ;
        RECT 42.865 184.790 43.215 184.960 ;
        RECT 43.425 184.600 43.755 185.060 ;
        RECT 44.630 184.990 44.800 185.700 ;
        RECT 45.155 185.500 45.325 186.090 ;
        RECT 44.970 185.280 45.325 185.500 ;
        RECT 45.495 185.280 45.845 185.900 ;
        RECT 46.015 184.990 46.185 186.350 ;
        RECT 46.550 186.180 46.875 186.965 ;
        RECT 46.355 185.130 46.815 186.180 ;
        RECT 44.630 184.820 45.485 184.990 ;
        RECT 45.690 184.820 46.185 184.990 ;
        RECT 46.355 184.600 46.685 184.960 ;
        RECT 47.045 184.860 47.215 186.980 ;
        RECT 47.385 186.650 47.715 187.150 ;
        RECT 47.885 186.480 48.140 186.980 ;
        RECT 47.390 186.310 48.140 186.480 ;
        RECT 47.390 185.320 47.620 186.310 ;
        RECT 47.790 185.490 48.140 186.140 ;
        RECT 48.355 186.010 48.585 187.150 ;
        RECT 48.755 186.000 49.085 186.980 ;
        RECT 49.255 186.010 49.465 187.150 ;
        RECT 48.335 185.590 48.665 185.840 ;
        RECT 47.390 185.150 48.140 185.320 ;
        RECT 47.385 184.600 47.715 184.980 ;
        RECT 47.885 184.860 48.140 185.150 ;
        RECT 48.355 184.600 48.585 185.420 ;
        RECT 48.835 185.400 49.085 186.000 ;
        RECT 49.700 185.960 49.955 186.840 ;
        RECT 50.125 186.010 50.430 187.150 ;
        RECT 50.770 186.770 51.100 187.150 ;
        RECT 51.280 186.600 51.450 186.890 ;
        RECT 51.620 186.690 51.870 187.150 ;
        RECT 50.650 186.430 51.450 186.600 ;
        RECT 52.040 186.640 52.910 186.980 ;
        RECT 48.755 184.770 49.085 185.400 ;
        RECT 49.255 184.600 49.465 185.420 ;
        RECT 49.700 185.310 49.910 185.960 ;
        RECT 50.650 185.840 50.820 186.430 ;
        RECT 52.040 186.260 52.210 186.640 ;
        RECT 53.145 186.520 53.315 186.980 ;
        RECT 53.485 186.690 53.855 187.150 ;
        RECT 54.150 186.550 54.320 186.890 ;
        RECT 54.490 186.720 54.820 187.150 ;
        RECT 55.055 186.550 55.225 186.890 ;
        RECT 50.990 186.090 52.210 186.260 ;
        RECT 52.380 186.180 52.840 186.470 ;
        RECT 53.145 186.350 53.705 186.520 ;
        RECT 54.150 186.380 55.225 186.550 ;
        RECT 55.395 186.650 56.075 186.980 ;
        RECT 56.290 186.650 56.540 186.980 ;
        RECT 56.710 186.690 56.960 187.150 ;
        RECT 53.535 186.210 53.705 186.350 ;
        RECT 52.380 186.170 53.345 186.180 ;
        RECT 52.040 186.000 52.210 186.090 ;
        RECT 52.670 186.010 53.345 186.170 ;
        RECT 50.080 185.810 50.820 185.840 ;
        RECT 50.080 185.510 50.995 185.810 ;
        RECT 50.670 185.335 50.995 185.510 ;
        RECT 49.700 184.780 49.955 185.310 ;
        RECT 50.125 184.600 50.430 185.060 ;
        RECT 50.675 184.980 50.995 185.335 ;
        RECT 51.165 185.550 51.705 185.920 ;
        RECT 52.040 185.830 52.445 186.000 ;
        RECT 51.165 185.150 51.405 185.550 ;
        RECT 51.885 185.380 52.105 185.660 ;
        RECT 51.575 185.210 52.105 185.380 ;
        RECT 51.575 184.980 51.745 185.210 ;
        RECT 52.275 185.050 52.445 185.830 ;
        RECT 52.615 185.220 52.965 185.840 ;
        RECT 53.135 185.220 53.345 186.010 ;
        RECT 53.535 186.040 55.035 186.210 ;
        RECT 53.535 185.350 53.705 186.040 ;
        RECT 55.395 185.870 55.565 186.650 ;
        RECT 56.370 186.520 56.540 186.650 ;
        RECT 53.875 185.700 55.565 185.870 ;
        RECT 55.735 186.090 56.200 186.480 ;
        RECT 56.370 186.350 56.765 186.520 ;
        RECT 53.875 185.520 54.045 185.700 ;
        RECT 50.675 184.810 51.745 184.980 ;
        RECT 51.915 184.600 52.105 185.040 ;
        RECT 52.275 184.770 53.225 185.050 ;
        RECT 53.535 184.960 53.795 185.350 ;
        RECT 54.215 185.280 55.005 185.530 ;
        RECT 53.445 184.790 53.795 184.960 ;
        RECT 54.005 184.600 54.335 185.060 ;
        RECT 55.210 184.990 55.380 185.700 ;
        RECT 55.735 185.500 55.905 186.090 ;
        RECT 55.550 185.280 55.905 185.500 ;
        RECT 56.075 185.280 56.425 185.900 ;
        RECT 56.595 184.990 56.765 186.350 ;
        RECT 57.130 186.180 57.455 186.965 ;
        RECT 56.935 185.130 57.395 186.180 ;
        RECT 55.210 184.820 56.065 184.990 ;
        RECT 56.270 184.820 56.765 184.990 ;
        RECT 56.935 184.600 57.265 184.960 ;
        RECT 57.625 184.860 57.795 186.980 ;
        RECT 57.965 186.650 58.295 187.150 ;
        RECT 58.465 186.480 58.720 186.980 ;
        RECT 57.970 186.310 58.720 186.480 ;
        RECT 57.970 185.320 58.200 186.310 ;
        RECT 58.370 185.490 58.720 186.140 ;
        RECT 58.895 186.060 60.565 187.150 ;
        RECT 58.895 185.540 59.645 186.060 ;
        RECT 59.815 185.370 60.565 185.890 ;
        RECT 57.970 185.150 58.720 185.320 ;
        RECT 57.965 184.600 58.295 184.980 ;
        RECT 58.465 184.860 58.720 185.150 ;
        RECT 58.895 184.600 60.565 185.370 ;
        RECT 60.735 185.340 60.995 186.965 ;
        RECT 62.745 186.700 63.075 187.150 ;
        RECT 61.175 186.310 63.785 186.520 ;
        RECT 61.175 185.510 61.395 186.310 ;
        RECT 61.635 185.510 61.935 186.130 ;
        RECT 62.105 185.510 62.435 186.130 ;
        RECT 62.605 185.510 62.925 186.130 ;
        RECT 63.095 185.510 63.445 186.130 ;
        RECT 63.615 185.340 63.785 186.310 ;
        RECT 63.955 185.985 64.245 187.150 ;
        RECT 64.415 186.060 66.085 187.150 ;
        RECT 66.260 186.715 71.605 187.150 ;
        RECT 64.415 185.540 65.165 186.060 ;
        RECT 65.335 185.370 66.085 185.890 ;
        RECT 67.850 185.465 68.200 186.715 ;
        RECT 71.835 186.010 72.045 187.150 ;
        RECT 72.215 186.000 72.545 186.980 ;
        RECT 72.715 186.010 72.945 187.150 ;
        RECT 73.530 186.170 73.785 186.840 ;
        RECT 73.965 186.350 74.250 187.150 ;
        RECT 74.430 186.430 74.760 186.940 ;
        RECT 60.735 185.170 62.575 185.340 ;
        RECT 61.005 184.600 61.335 184.995 ;
        RECT 61.505 184.815 61.705 185.170 ;
        RECT 61.875 184.600 62.205 185.000 ;
        RECT 62.375 184.825 62.575 185.170 ;
        RECT 62.745 184.600 63.075 185.340 ;
        RECT 63.310 185.170 63.785 185.340 ;
        RECT 63.310 184.920 63.480 185.170 ;
        RECT 63.955 184.600 64.245 185.325 ;
        RECT 64.415 184.600 66.085 185.370 ;
        RECT 69.680 185.145 70.020 185.975 ;
        RECT 66.260 184.600 71.605 185.145 ;
        RECT 71.835 184.600 72.045 185.420 ;
        RECT 72.215 185.400 72.465 186.000 ;
        RECT 72.635 185.590 72.965 185.840 ;
        RECT 72.215 184.770 72.545 185.400 ;
        RECT 72.715 184.600 72.945 185.420 ;
        RECT 73.530 185.310 73.710 186.170 ;
        RECT 74.430 185.840 74.680 186.430 ;
        RECT 75.030 186.280 75.200 186.890 ;
        RECT 75.370 186.460 75.700 187.150 ;
        RECT 75.930 186.600 76.170 186.890 ;
        RECT 76.370 186.770 76.790 187.150 ;
        RECT 76.970 186.680 77.600 186.930 ;
        RECT 78.070 186.770 78.400 187.150 ;
        RECT 76.970 186.600 77.140 186.680 ;
        RECT 78.570 186.600 78.740 186.890 ;
        RECT 78.920 186.770 79.300 187.150 ;
        RECT 79.540 186.765 80.370 186.935 ;
        RECT 75.930 186.430 77.140 186.600 ;
        RECT 73.880 185.510 74.680 185.840 ;
        RECT 73.530 185.110 73.785 185.310 ;
        RECT 73.445 184.940 73.785 185.110 ;
        RECT 73.530 184.780 73.785 184.940 ;
        RECT 73.965 184.600 74.250 185.060 ;
        RECT 74.430 184.860 74.680 185.510 ;
        RECT 74.880 186.260 75.200 186.280 ;
        RECT 74.880 186.090 76.800 186.260 ;
        RECT 74.880 185.195 75.070 186.090 ;
        RECT 76.970 185.920 77.140 186.430 ;
        RECT 77.310 186.170 77.830 186.480 ;
        RECT 75.240 185.750 77.140 185.920 ;
        RECT 75.240 185.690 75.570 185.750 ;
        RECT 75.720 185.520 76.050 185.580 ;
        RECT 75.390 185.250 76.050 185.520 ;
        RECT 74.880 184.865 75.200 185.195 ;
        RECT 75.380 184.600 76.040 185.080 ;
        RECT 76.240 184.990 76.410 185.750 ;
        RECT 77.310 185.580 77.490 185.990 ;
        RECT 76.580 185.410 76.910 185.530 ;
        RECT 77.660 185.410 77.830 186.170 ;
        RECT 76.580 185.240 77.830 185.410 ;
        RECT 78.000 186.350 79.370 186.600 ;
        RECT 78.000 185.580 78.190 186.350 ;
        RECT 79.120 186.090 79.370 186.350 ;
        RECT 78.360 185.920 78.610 186.080 ;
        RECT 79.540 185.920 79.710 186.765 ;
        RECT 80.605 186.480 80.775 186.980 ;
        RECT 80.945 186.650 81.275 187.150 ;
        RECT 79.880 186.090 80.380 186.470 ;
        RECT 80.605 186.310 81.300 186.480 ;
        RECT 78.360 185.750 79.710 185.920 ;
        RECT 79.290 185.710 79.710 185.750 ;
        RECT 78.000 185.240 78.420 185.580 ;
        RECT 78.710 185.250 79.120 185.580 ;
        RECT 76.240 184.820 77.090 184.990 ;
        RECT 77.650 184.600 77.970 185.060 ;
        RECT 78.170 184.810 78.420 185.240 ;
        RECT 78.710 184.600 79.120 185.040 ;
        RECT 79.290 184.980 79.460 185.710 ;
        RECT 79.630 185.160 79.980 185.530 ;
        RECT 80.160 185.220 80.380 186.090 ;
        RECT 80.550 185.520 80.960 186.140 ;
        RECT 81.130 185.340 81.300 186.310 ;
        RECT 80.605 185.150 81.300 185.340 ;
        RECT 79.290 184.780 80.305 184.980 ;
        RECT 80.605 184.820 80.775 185.150 ;
        RECT 80.945 184.600 81.275 184.980 ;
        RECT 81.490 184.860 81.715 186.980 ;
        RECT 81.885 186.650 82.215 187.150 ;
        RECT 82.385 186.480 82.555 186.980 ;
        RECT 82.820 186.715 88.165 187.150 ;
        RECT 81.890 186.310 82.555 186.480 ;
        RECT 81.890 185.320 82.120 186.310 ;
        RECT 82.290 185.490 82.640 186.140 ;
        RECT 84.410 185.465 84.760 186.715 ;
        RECT 88.375 186.010 88.605 187.150 ;
        RECT 88.775 186.000 89.105 186.980 ;
        RECT 89.275 186.010 89.485 187.150 ;
        RECT 81.890 185.150 82.555 185.320 ;
        RECT 81.885 184.600 82.215 184.980 ;
        RECT 82.385 184.860 82.555 185.150 ;
        RECT 86.240 185.145 86.580 185.975 ;
        RECT 88.355 185.590 88.685 185.840 ;
        RECT 82.820 184.600 88.165 185.145 ;
        RECT 88.375 184.600 88.605 185.420 ;
        RECT 88.855 185.400 89.105 186.000 ;
        RECT 89.715 185.985 90.005 187.150 ;
        RECT 90.180 186.480 90.435 186.980 ;
        RECT 90.605 186.650 90.935 187.150 ;
        RECT 90.180 186.310 90.930 186.480 ;
        RECT 90.180 185.490 90.530 186.140 ;
        RECT 88.775 184.770 89.105 185.400 ;
        RECT 89.275 184.600 89.485 185.420 ;
        RECT 89.715 184.600 90.005 185.325 ;
        RECT 90.700 185.320 90.930 186.310 ;
        RECT 90.180 185.150 90.930 185.320 ;
        RECT 90.180 184.860 90.435 185.150 ;
        RECT 90.605 184.600 90.935 184.980 ;
        RECT 91.105 184.860 91.275 186.980 ;
        RECT 91.445 186.180 91.770 186.965 ;
        RECT 91.940 186.690 92.190 187.150 ;
        RECT 92.360 186.650 92.610 186.980 ;
        RECT 92.825 186.650 93.505 186.980 ;
        RECT 92.360 186.520 92.530 186.650 ;
        RECT 92.135 186.350 92.530 186.520 ;
        RECT 91.505 185.130 91.965 186.180 ;
        RECT 92.135 184.990 92.305 186.350 ;
        RECT 92.700 186.090 93.165 186.480 ;
        RECT 92.475 185.280 92.825 185.900 ;
        RECT 92.995 185.500 93.165 186.090 ;
        RECT 93.335 185.870 93.505 186.650 ;
        RECT 93.675 186.550 93.845 186.890 ;
        RECT 94.080 186.720 94.410 187.150 ;
        RECT 94.580 186.550 94.750 186.890 ;
        RECT 95.045 186.690 95.415 187.150 ;
        RECT 93.675 186.380 94.750 186.550 ;
        RECT 95.585 186.520 95.755 186.980 ;
        RECT 95.990 186.640 96.860 186.980 ;
        RECT 97.030 186.690 97.280 187.150 ;
        RECT 95.195 186.350 95.755 186.520 ;
        RECT 95.195 186.210 95.365 186.350 ;
        RECT 93.865 186.040 95.365 186.210 ;
        RECT 96.060 186.180 96.520 186.470 ;
        RECT 93.335 185.700 95.025 185.870 ;
        RECT 92.995 185.280 93.350 185.500 ;
        RECT 93.520 184.990 93.690 185.700 ;
        RECT 93.895 185.280 94.685 185.530 ;
        RECT 94.855 185.520 95.025 185.700 ;
        RECT 95.195 185.350 95.365 186.040 ;
        RECT 91.635 184.600 91.965 184.960 ;
        RECT 92.135 184.820 92.630 184.990 ;
        RECT 92.835 184.820 93.690 184.990 ;
        RECT 94.565 184.600 94.895 185.060 ;
        RECT 95.105 184.960 95.365 185.350 ;
        RECT 95.555 186.170 96.520 186.180 ;
        RECT 96.690 186.260 96.860 186.640 ;
        RECT 97.450 186.600 97.620 186.890 ;
        RECT 97.800 186.770 98.130 187.150 ;
        RECT 97.450 186.430 98.250 186.600 ;
        RECT 95.555 186.010 96.230 186.170 ;
        RECT 96.690 186.090 97.910 186.260 ;
        RECT 95.555 185.220 95.765 186.010 ;
        RECT 96.690 186.000 96.860 186.090 ;
        RECT 95.935 185.220 96.285 185.840 ;
        RECT 96.455 185.830 96.860 186.000 ;
        RECT 96.455 185.050 96.625 185.830 ;
        RECT 96.795 185.380 97.015 185.660 ;
        RECT 97.195 185.550 97.735 185.920 ;
        RECT 98.080 185.840 98.250 186.430 ;
        RECT 98.470 186.010 98.775 187.150 ;
        RECT 98.945 185.960 99.200 186.840 ;
        RECT 98.080 185.810 98.820 185.840 ;
        RECT 96.795 185.210 97.325 185.380 ;
        RECT 95.105 184.790 95.455 184.960 ;
        RECT 95.675 184.770 96.625 185.050 ;
        RECT 96.795 184.600 96.985 185.040 ;
        RECT 97.155 184.980 97.325 185.210 ;
        RECT 97.495 185.150 97.735 185.550 ;
        RECT 97.905 185.510 98.820 185.810 ;
        RECT 97.905 185.335 98.230 185.510 ;
        RECT 97.905 184.980 98.225 185.335 ;
        RECT 98.990 185.310 99.200 185.960 ;
        RECT 99.375 186.060 101.045 187.150 ;
        RECT 101.305 186.220 101.475 186.980 ;
        RECT 101.655 186.390 101.985 187.150 ;
        RECT 99.375 185.540 100.125 186.060 ;
        RECT 101.305 186.050 101.970 186.220 ;
        RECT 102.155 186.075 102.425 186.980 ;
        RECT 101.800 185.905 101.970 186.050 ;
        RECT 100.295 185.370 101.045 185.890 ;
        RECT 101.235 185.500 101.565 185.870 ;
        RECT 101.800 185.575 102.085 185.905 ;
        RECT 97.155 184.810 98.225 184.980 ;
        RECT 98.470 184.600 98.775 185.060 ;
        RECT 98.945 184.780 99.200 185.310 ;
        RECT 99.375 184.600 101.045 185.370 ;
        RECT 101.800 185.320 101.970 185.575 ;
        RECT 101.305 185.150 101.970 185.320 ;
        RECT 102.255 185.275 102.425 186.075 ;
        RECT 102.595 186.390 103.110 186.800 ;
        RECT 103.345 186.390 103.515 187.150 ;
        RECT 103.685 186.810 105.715 186.980 ;
        RECT 102.595 185.580 102.935 186.390 ;
        RECT 103.685 186.145 103.855 186.810 ;
        RECT 104.250 186.470 105.375 186.640 ;
        RECT 103.105 185.955 103.855 186.145 ;
        RECT 104.025 186.130 105.035 186.300 ;
        RECT 102.595 185.410 103.825 185.580 ;
        RECT 101.305 184.770 101.475 185.150 ;
        RECT 101.655 184.600 101.985 184.980 ;
        RECT 102.165 184.770 102.425 185.275 ;
        RECT 102.870 184.805 103.115 185.410 ;
        RECT 103.335 184.600 103.845 185.135 ;
        RECT 104.025 184.770 104.215 186.130 ;
        RECT 104.385 185.450 104.660 185.930 ;
        RECT 104.385 185.280 104.665 185.450 ;
        RECT 104.865 185.330 105.035 186.130 ;
        RECT 105.205 185.340 105.375 186.470 ;
        RECT 105.545 185.840 105.715 186.810 ;
        RECT 105.885 186.010 106.055 187.150 ;
        RECT 106.225 186.010 106.560 186.980 ;
        RECT 105.545 185.510 105.740 185.840 ;
        RECT 105.965 185.510 106.220 185.840 ;
        RECT 105.965 185.340 106.135 185.510 ;
        RECT 106.390 185.340 106.560 186.010 ;
        RECT 104.385 184.770 104.660 185.280 ;
        RECT 105.205 185.170 106.135 185.340 ;
        RECT 105.205 185.135 105.380 185.170 ;
        RECT 104.850 184.770 105.380 185.135 ;
        RECT 105.805 184.600 106.135 185.000 ;
        RECT 106.305 184.770 106.560 185.340 ;
        RECT 106.735 186.010 107.120 186.980 ;
        RECT 107.290 186.690 107.615 187.150 ;
        RECT 108.135 186.520 108.415 186.980 ;
        RECT 107.290 186.300 108.415 186.520 ;
        RECT 106.735 185.340 107.015 186.010 ;
        RECT 107.290 185.840 107.740 186.300 ;
        RECT 108.605 186.130 109.005 186.980 ;
        RECT 109.405 186.690 109.675 187.150 ;
        RECT 109.845 186.520 110.130 186.980 ;
        RECT 107.185 185.510 107.740 185.840 ;
        RECT 107.910 185.570 109.005 186.130 ;
        RECT 107.290 185.400 107.740 185.510 ;
        RECT 106.735 184.770 107.120 185.340 ;
        RECT 107.290 185.230 108.415 185.400 ;
        RECT 107.290 184.600 107.615 185.060 ;
        RECT 108.135 184.770 108.415 185.230 ;
        RECT 108.605 184.770 109.005 185.570 ;
        RECT 109.175 186.300 110.130 186.520 ;
        RECT 109.175 185.400 109.385 186.300 ;
        RECT 109.555 185.570 110.245 186.130 ;
        RECT 110.875 186.060 114.385 187.150 ;
        RECT 114.555 186.060 115.765 187.150 ;
        RECT 110.875 185.540 112.565 186.060 ;
        RECT 109.175 185.230 110.130 185.400 ;
        RECT 112.735 185.370 114.385 185.890 ;
        RECT 114.555 185.520 115.075 186.060 ;
        RECT 109.405 184.600 109.675 185.060 ;
        RECT 109.845 184.770 110.130 185.230 ;
        RECT 110.875 184.600 114.385 185.370 ;
        RECT 115.245 185.350 115.765 185.890 ;
        RECT 114.555 184.600 115.765 185.350 ;
        RECT 10.510 184.430 115.850 184.600 ;
        RECT 10.595 183.680 11.805 184.430 ;
        RECT 10.595 183.140 11.115 183.680 ;
        RECT 12.435 183.660 14.105 184.430 ;
        RECT 14.280 183.885 19.625 184.430 ;
        RECT 19.800 183.885 25.145 184.430 ;
        RECT 11.285 182.970 11.805 183.510 ;
        RECT 10.595 181.880 11.805 182.970 ;
        RECT 12.435 182.970 13.185 183.490 ;
        RECT 13.355 183.140 14.105 183.660 ;
        RECT 12.435 181.880 14.105 182.970 ;
        RECT 15.870 182.315 16.220 183.565 ;
        RECT 17.700 183.055 18.040 183.885 ;
        RECT 21.390 182.315 21.740 183.565 ;
        RECT 23.220 183.055 23.560 183.885 ;
        RECT 25.315 183.705 25.605 184.430 ;
        RECT 25.835 183.610 26.045 184.430 ;
        RECT 26.215 183.630 26.545 184.260 ;
        RECT 14.280 181.880 19.625 182.315 ;
        RECT 19.800 181.880 25.145 182.315 ;
        RECT 25.315 181.880 25.605 183.045 ;
        RECT 26.215 183.030 26.465 183.630 ;
        RECT 26.715 183.610 26.945 184.430 ;
        RECT 27.155 183.680 28.365 184.430 ;
        RECT 28.625 183.880 28.795 184.260 ;
        RECT 28.975 184.050 29.305 184.430 ;
        RECT 28.625 183.710 29.290 183.880 ;
        RECT 29.485 183.755 29.745 184.260 ;
        RECT 26.635 183.190 26.965 183.440 ;
        RECT 25.835 181.880 26.045 183.020 ;
        RECT 26.215 182.050 26.545 183.030 ;
        RECT 26.715 181.880 26.945 183.020 ;
        RECT 27.155 182.970 27.675 183.510 ;
        RECT 27.845 183.140 28.365 183.680 ;
        RECT 28.555 183.160 28.885 183.530 ;
        RECT 29.120 183.455 29.290 183.710 ;
        RECT 29.120 183.125 29.405 183.455 ;
        RECT 29.120 182.980 29.290 183.125 ;
        RECT 27.155 181.880 28.365 182.970 ;
        RECT 28.625 182.810 29.290 182.980 ;
        RECT 29.575 182.955 29.745 183.755 ;
        RECT 28.625 182.050 28.795 182.810 ;
        RECT 28.975 181.880 29.305 182.640 ;
        RECT 29.475 182.050 29.745 182.955 ;
        RECT 29.915 183.755 30.175 184.260 ;
        RECT 30.355 184.050 30.685 184.430 ;
        RECT 30.865 183.880 31.035 184.260 ;
        RECT 29.915 182.955 30.085 183.755 ;
        RECT 30.370 183.710 31.035 183.880 ;
        RECT 30.370 183.455 30.540 183.710 ;
        RECT 31.295 183.660 32.965 184.430 ;
        RECT 33.225 183.880 33.395 184.260 ;
        RECT 33.575 184.050 33.905 184.430 ;
        RECT 33.225 183.710 33.890 183.880 ;
        RECT 34.085 183.755 34.345 184.260 ;
        RECT 30.255 183.125 30.540 183.455 ;
        RECT 30.775 183.160 31.105 183.530 ;
        RECT 30.370 182.980 30.540 183.125 ;
        RECT 29.915 182.050 30.185 182.955 ;
        RECT 30.370 182.810 31.035 182.980 ;
        RECT 30.355 181.880 30.685 182.640 ;
        RECT 30.865 182.050 31.035 182.810 ;
        RECT 31.295 182.970 32.045 183.490 ;
        RECT 32.215 183.140 32.965 183.660 ;
        RECT 33.155 183.160 33.485 183.530 ;
        RECT 33.720 183.455 33.890 183.710 ;
        RECT 33.720 183.125 34.005 183.455 ;
        RECT 33.720 182.980 33.890 183.125 ;
        RECT 31.295 181.880 32.965 182.970 ;
        RECT 33.225 182.810 33.890 182.980 ;
        RECT 34.175 182.955 34.345 183.755 ;
        RECT 34.630 183.800 34.915 184.260 ;
        RECT 35.085 183.970 35.355 184.430 ;
        RECT 34.630 183.630 35.585 183.800 ;
        RECT 33.225 182.050 33.395 182.810 ;
        RECT 33.575 181.880 33.905 182.640 ;
        RECT 34.075 182.050 34.345 182.955 ;
        RECT 34.515 182.900 35.205 183.460 ;
        RECT 35.375 182.730 35.585 183.630 ;
        RECT 34.630 182.510 35.585 182.730 ;
        RECT 35.755 183.460 36.155 184.260 ;
        RECT 36.345 183.800 36.625 184.260 ;
        RECT 37.145 183.970 37.470 184.430 ;
        RECT 36.345 183.630 37.470 183.800 ;
        RECT 37.640 183.690 38.025 184.260 ;
        RECT 37.020 183.520 37.470 183.630 ;
        RECT 35.755 182.900 36.850 183.460 ;
        RECT 37.020 183.190 37.575 183.520 ;
        RECT 34.630 182.050 34.915 182.510 ;
        RECT 35.085 181.880 35.355 182.340 ;
        RECT 35.755 182.050 36.155 182.900 ;
        RECT 37.020 182.730 37.470 183.190 ;
        RECT 37.745 183.020 38.025 183.690 ;
        RECT 38.470 183.620 38.715 184.225 ;
        RECT 38.935 183.895 39.445 184.430 ;
        RECT 36.345 182.510 37.470 182.730 ;
        RECT 36.345 182.050 36.625 182.510 ;
        RECT 37.145 181.880 37.470 182.340 ;
        RECT 37.640 182.050 38.025 183.020 ;
        RECT 38.195 183.450 39.425 183.620 ;
        RECT 38.195 182.640 38.535 183.450 ;
        RECT 38.705 182.885 39.455 183.075 ;
        RECT 38.195 182.230 38.710 182.640 ;
        RECT 38.945 181.880 39.115 182.640 ;
        RECT 39.285 182.220 39.455 182.885 ;
        RECT 39.625 182.900 39.815 184.260 ;
        RECT 39.985 184.090 40.260 184.260 ;
        RECT 39.985 183.920 40.265 184.090 ;
        RECT 39.985 183.100 40.260 183.920 ;
        RECT 40.450 183.895 40.980 184.260 ;
        RECT 41.405 184.030 41.735 184.430 ;
        RECT 40.805 183.860 40.980 183.895 ;
        RECT 40.465 182.900 40.635 183.700 ;
        RECT 39.625 182.730 40.635 182.900 ;
        RECT 40.805 183.690 41.735 183.860 ;
        RECT 41.905 183.690 42.160 184.260 ;
        RECT 40.805 182.560 40.975 183.690 ;
        RECT 41.565 183.520 41.735 183.690 ;
        RECT 39.850 182.390 40.975 182.560 ;
        RECT 41.145 183.190 41.340 183.520 ;
        RECT 41.565 183.190 41.820 183.520 ;
        RECT 41.145 182.220 41.315 183.190 ;
        RECT 41.990 183.020 42.160 183.690 ;
        RECT 42.610 183.620 42.855 184.225 ;
        RECT 43.075 183.895 43.585 184.430 ;
        RECT 39.285 182.050 41.315 182.220 ;
        RECT 41.485 181.880 41.655 183.020 ;
        RECT 41.825 182.050 42.160 183.020 ;
        RECT 42.335 183.450 43.565 183.620 ;
        RECT 42.335 182.640 42.675 183.450 ;
        RECT 42.845 182.885 43.595 183.075 ;
        RECT 42.335 182.230 42.850 182.640 ;
        RECT 43.085 181.880 43.255 182.640 ;
        RECT 43.425 182.220 43.595 182.885 ;
        RECT 43.765 182.900 43.955 184.260 ;
        RECT 44.125 183.410 44.400 184.260 ;
        RECT 44.590 183.895 45.120 184.260 ;
        RECT 45.545 184.030 45.875 184.430 ;
        RECT 44.945 183.860 45.120 183.895 ;
        RECT 44.125 183.240 44.405 183.410 ;
        RECT 44.125 183.100 44.400 183.240 ;
        RECT 44.605 182.900 44.775 183.700 ;
        RECT 43.765 182.730 44.775 182.900 ;
        RECT 44.945 183.690 45.875 183.860 ;
        RECT 46.045 183.690 46.300 184.260 ;
        RECT 44.945 182.560 45.115 183.690 ;
        RECT 45.705 183.520 45.875 183.690 ;
        RECT 43.990 182.390 45.115 182.560 ;
        RECT 45.285 183.190 45.480 183.520 ;
        RECT 45.705 183.190 45.960 183.520 ;
        RECT 45.285 182.220 45.455 183.190 ;
        RECT 46.130 183.020 46.300 183.690 ;
        RECT 47.210 183.620 47.455 184.225 ;
        RECT 47.675 183.895 48.185 184.430 ;
        RECT 43.425 182.050 45.455 182.220 ;
        RECT 45.625 181.880 45.795 183.020 ;
        RECT 45.965 182.050 46.300 183.020 ;
        RECT 46.935 183.450 48.165 183.620 ;
        RECT 46.935 182.640 47.275 183.450 ;
        RECT 47.445 182.885 48.195 183.075 ;
        RECT 46.935 182.230 47.450 182.640 ;
        RECT 47.685 181.880 47.855 182.640 ;
        RECT 48.025 182.220 48.195 182.885 ;
        RECT 48.365 182.900 48.555 184.260 ;
        RECT 48.725 183.410 49.000 184.260 ;
        RECT 49.190 183.895 49.720 184.260 ;
        RECT 50.145 184.030 50.475 184.430 ;
        RECT 49.545 183.860 49.720 183.895 ;
        RECT 48.725 183.240 49.005 183.410 ;
        RECT 48.725 183.100 49.000 183.240 ;
        RECT 49.205 182.900 49.375 183.700 ;
        RECT 48.365 182.730 49.375 182.900 ;
        RECT 49.545 183.690 50.475 183.860 ;
        RECT 50.645 183.690 50.900 184.260 ;
        RECT 51.075 183.705 51.365 184.430 ;
        RECT 51.625 183.880 51.795 184.260 ;
        RECT 51.975 184.050 52.305 184.430 ;
        RECT 51.625 183.710 52.290 183.880 ;
        RECT 52.485 183.755 52.745 184.260 ;
        RECT 49.545 182.560 49.715 183.690 ;
        RECT 50.305 183.520 50.475 183.690 ;
        RECT 48.590 182.390 49.715 182.560 ;
        RECT 49.885 183.190 50.080 183.520 ;
        RECT 50.305 183.190 50.560 183.520 ;
        RECT 49.885 182.220 50.055 183.190 ;
        RECT 50.730 183.020 50.900 183.690 ;
        RECT 51.555 183.160 51.885 183.530 ;
        RECT 52.120 183.455 52.290 183.710 ;
        RECT 52.120 183.125 52.405 183.455 ;
        RECT 48.025 182.050 50.055 182.220 ;
        RECT 50.225 181.880 50.395 183.020 ;
        RECT 50.565 182.050 50.900 183.020 ;
        RECT 51.075 181.880 51.365 183.045 ;
        RECT 52.120 182.980 52.290 183.125 ;
        RECT 51.625 182.810 52.290 182.980 ;
        RECT 52.575 182.955 52.745 183.755 ;
        RECT 53.835 183.660 57.345 184.430 ;
        RECT 57.785 184.035 58.115 184.430 ;
        RECT 58.285 183.860 58.485 184.215 ;
        RECT 58.655 184.030 58.985 184.430 ;
        RECT 59.155 183.860 59.355 184.205 ;
        RECT 51.625 182.050 51.795 182.810 ;
        RECT 51.975 181.880 52.305 182.640 ;
        RECT 52.475 182.050 52.745 182.955 ;
        RECT 53.835 182.970 55.525 183.490 ;
        RECT 55.695 183.140 57.345 183.660 ;
        RECT 57.515 183.690 59.355 183.860 ;
        RECT 59.525 183.690 59.855 184.430 ;
        RECT 60.090 183.860 60.260 184.110 ;
        RECT 60.090 183.690 60.565 183.860 ;
        RECT 60.930 183.690 61.180 184.430 ;
        RECT 53.835 181.880 57.345 182.970 ;
        RECT 57.515 182.065 57.775 183.690 ;
        RECT 57.955 182.720 58.175 183.520 ;
        RECT 58.415 182.900 58.715 183.520 ;
        RECT 58.885 182.900 59.215 183.520 ;
        RECT 59.385 182.900 59.705 183.520 ;
        RECT 59.875 182.900 60.225 183.520 ;
        RECT 60.395 182.720 60.565 183.690 ;
        RECT 61.350 183.610 61.705 184.135 ;
        RECT 61.875 183.620 62.080 184.430 ;
        RECT 62.250 183.790 62.580 184.260 ;
        RECT 62.750 183.960 62.920 184.430 ;
        RECT 63.090 183.790 63.420 184.260 ;
        RECT 63.590 183.960 64.315 184.430 ;
        RECT 64.485 183.790 64.815 184.260 ;
        RECT 64.985 183.960 65.155 184.430 ;
        RECT 65.325 183.790 65.655 184.260 ;
        RECT 61.535 183.440 61.705 183.610 ;
        RECT 62.250 183.610 65.655 183.790 ;
        RECT 65.825 183.610 66.085 184.430 ;
        RECT 62.250 183.440 62.455 183.610 ;
        RECT 57.955 182.510 60.565 182.720 ;
        RECT 60.735 183.230 61.365 183.440 ;
        RECT 61.535 183.270 61.850 183.440 ;
        RECT 60.735 182.560 60.985 183.230 ;
        RECT 61.535 182.480 61.705 183.270 ;
        RECT 62.135 183.060 62.455 183.440 ;
        RECT 62.635 183.230 63.355 183.440 ;
        RECT 63.535 183.230 64.750 183.440 ;
        RECT 64.930 183.230 66.070 183.440 ;
        RECT 62.135 182.890 62.540 183.060 ;
        RECT 59.525 181.880 59.855 182.330 ;
        RECT 60.930 181.880 61.180 182.380 ;
        RECT 61.350 182.065 61.705 182.480 ;
        RECT 61.875 182.220 62.120 182.720 ;
        RECT 62.290 182.390 62.540 182.890 ;
        RECT 62.710 182.890 63.895 183.060 ;
        RECT 62.710 182.220 62.960 182.890 ;
        RECT 61.875 182.050 62.960 182.220 ;
        RECT 63.130 182.220 63.340 182.720 ;
        RECT 63.510 182.390 63.895 182.890 ;
        RECT 64.065 182.890 66.085 183.060 ;
        RECT 64.065 182.390 64.395 182.890 ;
        RECT 64.565 182.220 64.775 182.720 ;
        RECT 63.130 182.050 64.775 182.220 ;
        RECT 64.945 182.050 65.195 182.890 ;
        RECT 65.365 181.880 65.575 182.720 ;
        RECT 65.745 182.050 66.085 182.890 ;
        RECT 66.255 182.050 66.515 184.260 ;
        RECT 66.685 184.050 67.015 184.430 ;
        RECT 67.225 183.520 67.420 184.095 ;
        RECT 67.690 183.520 67.875 184.100 ;
        RECT 66.685 182.600 66.855 183.520 ;
        RECT 67.165 183.190 67.420 183.520 ;
        RECT 67.645 183.190 67.875 183.520 ;
        RECT 68.125 184.090 69.605 184.260 ;
        RECT 68.125 183.190 68.295 184.090 ;
        RECT 68.465 183.590 69.015 183.920 ;
        RECT 69.205 183.760 69.605 184.090 ;
        RECT 69.785 184.050 70.115 184.430 ;
        RECT 70.425 183.930 70.685 184.260 ;
        RECT 67.225 182.880 67.420 183.190 ;
        RECT 67.690 182.880 67.875 183.190 ;
        RECT 68.465 182.600 68.635 183.590 ;
        RECT 69.205 183.280 69.375 183.760 ;
        RECT 69.955 183.570 70.165 183.750 ;
        RECT 69.545 183.400 70.165 183.570 ;
        RECT 66.685 182.430 68.635 182.600 ;
        RECT 68.805 183.110 69.375 183.280 ;
        RECT 70.515 183.230 70.685 183.930 ;
        RECT 70.855 183.660 72.525 184.430 ;
        RECT 68.805 182.600 68.975 183.110 ;
        RECT 69.555 183.060 70.685 183.230 ;
        RECT 69.555 182.940 69.725 183.060 ;
        RECT 69.145 182.770 69.725 182.940 ;
        RECT 68.805 182.430 69.545 182.600 ;
        RECT 69.995 182.560 70.345 182.890 ;
        RECT 66.685 181.880 67.015 182.260 ;
        RECT 67.440 182.050 67.610 182.430 ;
        RECT 67.870 181.880 68.200 182.260 ;
        RECT 68.395 182.050 68.565 182.430 ;
        RECT 68.775 181.880 69.105 182.260 ;
        RECT 69.355 182.050 69.545 182.430 ;
        RECT 70.515 182.380 70.685 183.060 ;
        RECT 69.785 181.880 70.115 182.260 ;
        RECT 70.425 182.050 70.685 182.380 ;
        RECT 70.855 182.970 71.605 183.490 ;
        RECT 71.775 183.140 72.525 183.660 ;
        RECT 72.970 183.620 73.215 184.225 ;
        RECT 73.435 183.895 73.945 184.430 ;
        RECT 72.695 183.450 73.925 183.620 ;
        RECT 70.855 181.880 72.525 182.970 ;
        RECT 72.695 182.640 73.035 183.450 ;
        RECT 73.205 182.885 73.955 183.075 ;
        RECT 72.695 182.230 73.210 182.640 ;
        RECT 73.445 181.880 73.615 182.640 ;
        RECT 73.785 182.220 73.955 182.885 ;
        RECT 74.125 182.900 74.315 184.260 ;
        RECT 74.485 183.410 74.760 184.260 ;
        RECT 74.950 183.895 75.480 184.260 ;
        RECT 75.905 184.030 76.235 184.430 ;
        RECT 75.305 183.860 75.480 183.895 ;
        RECT 74.485 183.240 74.765 183.410 ;
        RECT 74.485 183.100 74.760 183.240 ;
        RECT 74.965 182.900 75.135 183.700 ;
        RECT 74.125 182.730 75.135 182.900 ;
        RECT 75.305 183.690 76.235 183.860 ;
        RECT 76.405 183.690 76.660 184.260 ;
        RECT 76.835 183.705 77.125 184.430 ;
        RECT 77.385 183.780 77.555 184.260 ;
        RECT 77.735 183.950 77.975 184.430 ;
        RECT 78.225 183.780 78.395 184.260 ;
        RECT 78.565 183.950 78.895 184.430 ;
        RECT 79.065 183.780 79.235 184.260 ;
        RECT 75.305 182.560 75.475 183.690 ;
        RECT 76.065 183.520 76.235 183.690 ;
        RECT 74.350 182.390 75.475 182.560 ;
        RECT 75.645 183.190 75.840 183.520 ;
        RECT 76.065 183.190 76.320 183.520 ;
        RECT 75.645 182.220 75.815 183.190 ;
        RECT 76.490 183.020 76.660 183.690 ;
        RECT 77.385 183.610 78.020 183.780 ;
        RECT 78.225 183.610 79.235 183.780 ;
        RECT 79.405 183.630 79.735 184.430 ;
        RECT 80.145 183.880 80.315 184.260 ;
        RECT 80.495 184.050 80.825 184.430 ;
        RECT 80.145 183.710 80.810 183.880 ;
        RECT 81.005 183.755 81.265 184.260 ;
        RECT 81.495 183.950 81.775 184.430 ;
        RECT 81.945 183.780 82.205 184.170 ;
        RECT 82.380 183.950 82.635 184.430 ;
        RECT 82.805 183.780 83.100 184.170 ;
        RECT 83.280 183.950 83.555 184.430 ;
        RECT 83.725 183.930 84.025 184.260 ;
        RECT 77.850 183.440 78.020 183.610 ;
        RECT 77.300 183.200 77.680 183.440 ;
        RECT 77.850 183.270 78.350 183.440 ;
        RECT 73.785 182.050 75.815 182.220 ;
        RECT 75.985 181.880 76.155 183.020 ;
        RECT 76.325 182.050 76.660 183.020 ;
        RECT 76.835 181.880 77.125 183.045 ;
        RECT 77.850 183.030 78.020 183.270 ;
        RECT 78.740 183.070 79.235 183.610 ;
        RECT 80.075 183.160 80.405 183.530 ;
        RECT 80.640 183.455 80.810 183.710 ;
        RECT 77.305 182.860 78.020 183.030 ;
        RECT 78.225 182.900 79.235 183.070 ;
        RECT 80.640 183.125 80.925 183.455 ;
        RECT 77.305 182.050 77.635 182.860 ;
        RECT 77.805 181.880 78.045 182.680 ;
        RECT 78.225 182.050 78.395 182.900 ;
        RECT 78.565 181.880 78.895 182.680 ;
        RECT 79.065 182.050 79.235 182.900 ;
        RECT 79.405 181.880 79.735 183.030 ;
        RECT 80.640 182.980 80.810 183.125 ;
        RECT 80.145 182.810 80.810 182.980 ;
        RECT 81.095 182.955 81.265 183.755 ;
        RECT 80.145 182.050 80.315 182.810 ;
        RECT 80.495 181.880 80.825 182.640 ;
        RECT 80.995 182.050 81.265 182.955 ;
        RECT 81.450 183.610 83.100 183.780 ;
        RECT 81.450 183.100 81.855 183.610 ;
        RECT 82.025 183.270 83.165 183.440 ;
        RECT 81.450 182.930 82.205 183.100 ;
        RECT 81.490 181.880 81.775 182.750 ;
        RECT 81.945 182.680 82.205 182.930 ;
        RECT 82.995 183.020 83.165 183.270 ;
        RECT 83.335 183.190 83.685 183.760 ;
        RECT 83.855 183.020 84.025 183.930 ;
        RECT 82.995 182.850 84.025 183.020 ;
        RECT 81.945 182.510 83.065 182.680 ;
        RECT 81.945 182.050 82.205 182.510 ;
        RECT 82.380 181.880 82.635 182.340 ;
        RECT 82.805 182.050 83.065 182.510 ;
        RECT 83.235 181.880 83.545 182.680 ;
        RECT 83.715 182.050 84.025 182.850 ;
        RECT 84.200 183.720 84.455 184.250 ;
        RECT 84.625 183.970 84.930 184.430 ;
        RECT 85.175 184.050 86.245 184.220 ;
        RECT 84.200 183.070 84.410 183.720 ;
        RECT 85.175 183.695 85.495 184.050 ;
        RECT 85.170 183.520 85.495 183.695 ;
        RECT 84.580 183.220 85.495 183.520 ;
        RECT 85.665 183.480 85.905 183.880 ;
        RECT 86.075 183.820 86.245 184.050 ;
        RECT 86.415 183.990 86.605 184.430 ;
        RECT 86.775 183.980 87.725 184.260 ;
        RECT 87.945 184.070 88.295 184.240 ;
        RECT 86.075 183.650 86.605 183.820 ;
        RECT 84.580 183.190 85.320 183.220 ;
        RECT 84.200 182.190 84.455 183.070 ;
        RECT 84.625 181.880 84.930 183.020 ;
        RECT 85.150 182.600 85.320 183.190 ;
        RECT 85.665 183.110 86.205 183.480 ;
        RECT 86.385 183.370 86.605 183.650 ;
        RECT 86.775 183.200 86.945 183.980 ;
        RECT 86.540 183.030 86.945 183.200 ;
        RECT 87.115 183.190 87.465 183.810 ;
        RECT 86.540 182.940 86.710 183.030 ;
        RECT 87.635 183.020 87.845 183.810 ;
        RECT 85.490 182.770 86.710 182.940 ;
        RECT 87.170 182.860 87.845 183.020 ;
        RECT 85.150 182.430 85.950 182.600 ;
        RECT 85.270 181.880 85.600 182.260 ;
        RECT 85.780 182.140 85.950 182.430 ;
        RECT 86.540 182.390 86.710 182.770 ;
        RECT 86.880 182.850 87.845 182.860 ;
        RECT 88.035 183.680 88.295 184.070 ;
        RECT 88.505 183.970 88.835 184.430 ;
        RECT 89.710 184.040 90.565 184.210 ;
        RECT 90.770 184.040 91.265 184.210 ;
        RECT 91.435 184.070 91.765 184.430 ;
        RECT 88.035 182.990 88.205 183.680 ;
        RECT 88.375 183.330 88.545 183.510 ;
        RECT 88.715 183.500 89.505 183.750 ;
        RECT 89.710 183.330 89.880 184.040 ;
        RECT 90.050 183.530 90.405 183.750 ;
        RECT 88.375 183.160 90.065 183.330 ;
        RECT 86.880 182.560 87.340 182.850 ;
        RECT 88.035 182.820 89.535 182.990 ;
        RECT 88.035 182.680 88.205 182.820 ;
        RECT 87.645 182.510 88.205 182.680 ;
        RECT 86.120 181.880 86.370 182.340 ;
        RECT 86.540 182.050 87.410 182.390 ;
        RECT 87.645 182.050 87.815 182.510 ;
        RECT 88.650 182.480 89.725 182.650 ;
        RECT 87.985 181.880 88.355 182.340 ;
        RECT 88.650 182.140 88.820 182.480 ;
        RECT 88.990 181.880 89.320 182.310 ;
        RECT 89.555 182.140 89.725 182.480 ;
        RECT 89.895 182.380 90.065 183.160 ;
        RECT 90.235 182.940 90.405 183.530 ;
        RECT 90.575 183.130 90.925 183.750 ;
        RECT 90.235 182.550 90.700 182.940 ;
        RECT 91.095 182.680 91.265 184.040 ;
        RECT 91.435 182.850 91.895 183.900 ;
        RECT 90.870 182.510 91.265 182.680 ;
        RECT 90.870 182.380 91.040 182.510 ;
        RECT 89.895 182.050 90.575 182.380 ;
        RECT 90.790 182.050 91.040 182.380 ;
        RECT 91.210 181.880 91.460 182.340 ;
        RECT 91.630 182.065 91.955 182.850 ;
        RECT 92.125 182.050 92.295 184.170 ;
        RECT 92.465 184.050 92.795 184.430 ;
        RECT 92.965 183.880 93.220 184.170 ;
        RECT 92.470 183.710 93.220 183.880 ;
        RECT 92.470 182.720 92.700 183.710 ;
        RECT 93.670 183.620 93.915 184.225 ;
        RECT 94.135 183.895 94.645 184.430 ;
        RECT 92.870 182.890 93.220 183.540 ;
        RECT 93.395 183.450 94.625 183.620 ;
        RECT 92.470 182.550 93.220 182.720 ;
        RECT 92.465 181.880 92.795 182.380 ;
        RECT 92.965 182.050 93.220 182.550 ;
        RECT 93.395 182.640 93.735 183.450 ;
        RECT 93.905 182.885 94.655 183.075 ;
        RECT 93.395 182.230 93.910 182.640 ;
        RECT 94.145 181.880 94.315 182.640 ;
        RECT 94.485 182.220 94.655 182.885 ;
        RECT 94.825 182.900 95.015 184.260 ;
        RECT 95.185 183.750 95.460 184.260 ;
        RECT 95.650 183.895 96.180 184.260 ;
        RECT 96.605 184.030 96.935 184.430 ;
        RECT 96.005 183.860 96.180 183.895 ;
        RECT 95.185 183.580 95.465 183.750 ;
        RECT 95.185 183.100 95.460 183.580 ;
        RECT 95.665 182.900 95.835 183.700 ;
        RECT 94.825 182.730 95.835 182.900 ;
        RECT 96.005 183.690 96.935 183.860 ;
        RECT 97.105 183.690 97.360 184.260 ;
        RECT 96.005 182.560 96.175 183.690 ;
        RECT 96.765 183.520 96.935 183.690 ;
        RECT 95.050 182.390 96.175 182.560 ;
        RECT 96.345 183.190 96.540 183.520 ;
        RECT 96.765 183.190 97.020 183.520 ;
        RECT 96.345 182.220 96.515 183.190 ;
        RECT 97.190 183.020 97.360 183.690 ;
        RECT 98.730 183.620 98.975 184.225 ;
        RECT 99.195 183.895 99.705 184.430 ;
        RECT 94.485 182.050 96.515 182.220 ;
        RECT 96.685 181.880 96.855 183.020 ;
        RECT 97.025 182.050 97.360 183.020 ;
        RECT 98.455 183.450 99.685 183.620 ;
        RECT 98.455 182.640 98.795 183.450 ;
        RECT 98.965 182.885 99.715 183.075 ;
        RECT 98.455 182.230 98.970 182.640 ;
        RECT 99.205 181.880 99.375 182.640 ;
        RECT 99.545 182.220 99.715 182.885 ;
        RECT 99.885 182.900 100.075 184.260 ;
        RECT 100.245 184.090 100.520 184.260 ;
        RECT 100.245 183.920 100.525 184.090 ;
        RECT 100.245 183.100 100.520 183.920 ;
        RECT 100.710 183.895 101.240 184.260 ;
        RECT 101.665 184.030 101.995 184.430 ;
        RECT 101.065 183.860 101.240 183.895 ;
        RECT 100.725 182.900 100.895 183.700 ;
        RECT 99.885 182.730 100.895 182.900 ;
        RECT 101.065 183.690 101.995 183.860 ;
        RECT 102.165 183.690 102.420 184.260 ;
        RECT 102.595 183.705 102.885 184.430 ;
        RECT 101.065 182.560 101.235 183.690 ;
        RECT 101.825 183.520 101.995 183.690 ;
        RECT 100.110 182.390 101.235 182.560 ;
        RECT 101.405 183.190 101.600 183.520 ;
        RECT 101.825 183.190 102.080 183.520 ;
        RECT 101.405 182.220 101.575 183.190 ;
        RECT 102.250 183.020 102.420 183.690 ;
        RECT 103.115 183.610 103.325 184.430 ;
        RECT 103.495 183.630 103.825 184.260 ;
        RECT 99.545 182.050 101.575 182.220 ;
        RECT 101.745 181.880 101.915 183.020 ;
        RECT 102.085 182.050 102.420 183.020 ;
        RECT 102.595 181.880 102.885 183.045 ;
        RECT 103.495 183.030 103.745 183.630 ;
        RECT 103.995 183.610 104.225 184.430 ;
        RECT 105.360 183.720 105.615 184.250 ;
        RECT 105.785 183.970 106.090 184.430 ;
        RECT 106.335 184.050 107.405 184.220 ;
        RECT 103.915 183.190 104.245 183.440 ;
        RECT 105.360 183.070 105.570 183.720 ;
        RECT 106.335 183.695 106.655 184.050 ;
        RECT 106.330 183.520 106.655 183.695 ;
        RECT 105.740 183.220 106.655 183.520 ;
        RECT 106.825 183.480 107.065 183.880 ;
        RECT 107.235 183.820 107.405 184.050 ;
        RECT 107.575 183.990 107.765 184.430 ;
        RECT 107.935 183.980 108.885 184.260 ;
        RECT 109.105 184.070 109.455 184.240 ;
        RECT 107.235 183.650 107.765 183.820 ;
        RECT 105.740 183.190 106.480 183.220 ;
        RECT 103.115 181.880 103.325 183.020 ;
        RECT 103.495 182.050 103.825 183.030 ;
        RECT 103.995 181.880 104.225 183.020 ;
        RECT 105.360 182.190 105.615 183.070 ;
        RECT 105.785 181.880 106.090 183.020 ;
        RECT 106.310 182.600 106.480 183.190 ;
        RECT 106.825 183.110 107.365 183.480 ;
        RECT 107.545 183.370 107.765 183.650 ;
        RECT 107.935 183.200 108.105 183.980 ;
        RECT 107.700 183.030 108.105 183.200 ;
        RECT 108.275 183.190 108.625 183.810 ;
        RECT 107.700 182.940 107.870 183.030 ;
        RECT 108.795 183.020 109.005 183.810 ;
        RECT 106.650 182.770 107.870 182.940 ;
        RECT 108.330 182.860 109.005 183.020 ;
        RECT 106.310 182.430 107.110 182.600 ;
        RECT 106.430 181.880 106.760 182.260 ;
        RECT 106.940 182.140 107.110 182.430 ;
        RECT 107.700 182.390 107.870 182.770 ;
        RECT 108.040 182.850 109.005 182.860 ;
        RECT 109.195 183.680 109.455 184.070 ;
        RECT 109.665 183.970 109.995 184.430 ;
        RECT 110.870 184.040 111.725 184.210 ;
        RECT 111.930 184.040 112.425 184.210 ;
        RECT 112.595 184.070 112.925 184.430 ;
        RECT 109.195 182.990 109.365 183.680 ;
        RECT 109.535 183.330 109.705 183.510 ;
        RECT 109.875 183.500 110.665 183.750 ;
        RECT 110.870 183.330 111.040 184.040 ;
        RECT 111.210 183.530 111.565 183.750 ;
        RECT 109.535 183.160 111.225 183.330 ;
        RECT 108.040 182.560 108.500 182.850 ;
        RECT 109.195 182.820 110.695 182.990 ;
        RECT 109.195 182.680 109.365 182.820 ;
        RECT 108.805 182.510 109.365 182.680 ;
        RECT 107.280 181.880 107.530 182.340 ;
        RECT 107.700 182.050 108.570 182.390 ;
        RECT 108.805 182.050 108.975 182.510 ;
        RECT 109.810 182.480 110.885 182.650 ;
        RECT 109.145 181.880 109.515 182.340 ;
        RECT 109.810 182.140 109.980 182.480 ;
        RECT 110.150 181.880 110.480 182.310 ;
        RECT 110.715 182.140 110.885 182.480 ;
        RECT 111.055 182.380 111.225 183.160 ;
        RECT 111.395 182.940 111.565 183.530 ;
        RECT 111.735 183.130 112.085 183.750 ;
        RECT 111.395 182.550 111.860 182.940 ;
        RECT 112.255 182.680 112.425 184.040 ;
        RECT 112.595 182.850 113.055 183.900 ;
        RECT 112.030 182.510 112.425 182.680 ;
        RECT 112.030 182.380 112.200 182.510 ;
        RECT 111.055 182.050 111.735 182.380 ;
        RECT 111.950 182.050 112.200 182.380 ;
        RECT 112.370 181.880 112.620 182.340 ;
        RECT 112.790 182.065 113.115 182.850 ;
        RECT 113.285 182.050 113.455 184.170 ;
        RECT 113.625 184.050 113.955 184.430 ;
        RECT 114.125 183.880 114.380 184.170 ;
        RECT 113.630 183.710 114.380 183.880 ;
        RECT 113.630 182.720 113.860 183.710 ;
        RECT 114.555 183.680 115.765 184.430 ;
        RECT 114.030 182.890 114.380 183.540 ;
        RECT 114.555 182.970 115.075 183.510 ;
        RECT 115.245 183.140 115.765 183.680 ;
        RECT 113.630 182.550 114.380 182.720 ;
        RECT 113.625 181.880 113.955 182.380 ;
        RECT 114.125 182.050 114.380 182.550 ;
        RECT 114.555 181.880 115.765 182.970 ;
        RECT 10.510 181.710 115.850 181.880 ;
        RECT 10.595 180.620 11.805 181.710 ;
        RECT 10.595 179.910 11.115 180.450 ;
        RECT 11.285 180.080 11.805 180.620 ;
        RECT 12.435 180.545 12.725 181.710 ;
        RECT 12.895 180.620 14.105 181.710 ;
        RECT 14.280 181.275 19.625 181.710 ;
        RECT 12.895 180.080 13.415 180.620 ;
        RECT 13.585 179.910 14.105 180.450 ;
        RECT 15.870 180.025 16.220 181.275 ;
        RECT 19.910 181.080 20.195 181.540 ;
        RECT 20.365 181.250 20.635 181.710 ;
        RECT 19.910 180.860 20.865 181.080 ;
        RECT 10.595 179.160 11.805 179.910 ;
        RECT 12.435 179.160 12.725 179.885 ;
        RECT 12.895 179.160 14.105 179.910 ;
        RECT 17.700 179.705 18.040 180.535 ;
        RECT 19.795 180.130 20.485 180.690 ;
        RECT 20.655 179.960 20.865 180.860 ;
        RECT 19.910 179.790 20.865 179.960 ;
        RECT 21.035 180.690 21.435 181.540 ;
        RECT 21.625 181.080 21.905 181.540 ;
        RECT 22.425 181.250 22.750 181.710 ;
        RECT 21.625 180.860 22.750 181.080 ;
        RECT 21.035 180.130 22.130 180.690 ;
        RECT 22.300 180.400 22.750 180.860 ;
        RECT 22.920 180.570 23.305 181.540 ;
        RECT 23.590 181.080 23.875 181.540 ;
        RECT 24.045 181.250 24.315 181.710 ;
        RECT 23.590 180.860 24.545 181.080 ;
        RECT 14.280 179.160 19.625 179.705 ;
        RECT 19.910 179.330 20.195 179.790 ;
        RECT 20.365 179.160 20.635 179.620 ;
        RECT 21.035 179.330 21.435 180.130 ;
        RECT 22.300 180.070 22.855 180.400 ;
        RECT 22.300 179.960 22.750 180.070 ;
        RECT 21.625 179.790 22.750 179.960 ;
        RECT 23.025 179.900 23.305 180.570 ;
        RECT 23.475 180.130 24.165 180.690 ;
        RECT 24.335 179.960 24.545 180.860 ;
        RECT 21.625 179.330 21.905 179.790 ;
        RECT 22.425 179.160 22.750 179.620 ;
        RECT 22.920 179.330 23.305 179.900 ;
        RECT 23.590 179.790 24.545 179.960 ;
        RECT 24.715 180.690 25.115 181.540 ;
        RECT 25.305 181.080 25.585 181.540 ;
        RECT 26.105 181.250 26.430 181.710 ;
        RECT 25.305 180.860 26.430 181.080 ;
        RECT 24.715 180.130 25.810 180.690 ;
        RECT 25.980 180.400 26.430 180.860 ;
        RECT 26.600 180.570 26.985 181.540 ;
        RECT 23.590 179.330 23.875 179.790 ;
        RECT 24.045 179.160 24.315 179.620 ;
        RECT 24.715 179.330 25.115 180.130 ;
        RECT 25.980 180.070 26.535 180.400 ;
        RECT 25.980 179.960 26.430 180.070 ;
        RECT 25.305 179.790 26.430 179.960 ;
        RECT 26.705 179.900 26.985 180.570 ;
        RECT 27.155 180.950 27.670 181.360 ;
        RECT 27.905 180.950 28.075 181.710 ;
        RECT 28.245 181.370 30.275 181.540 ;
        RECT 27.155 180.140 27.495 180.950 ;
        RECT 28.245 180.705 28.415 181.370 ;
        RECT 28.810 181.030 29.935 181.200 ;
        RECT 27.665 180.515 28.415 180.705 ;
        RECT 28.585 180.690 29.595 180.860 ;
        RECT 27.155 179.970 28.385 180.140 ;
        RECT 25.305 179.330 25.585 179.790 ;
        RECT 26.105 179.160 26.430 179.620 ;
        RECT 26.600 179.330 26.985 179.900 ;
        RECT 27.430 179.365 27.675 179.970 ;
        RECT 27.895 179.160 28.405 179.695 ;
        RECT 28.585 179.330 28.775 180.690 ;
        RECT 28.945 179.670 29.220 180.490 ;
        RECT 29.425 179.890 29.595 180.690 ;
        RECT 29.765 179.900 29.935 181.030 ;
        RECT 30.105 180.400 30.275 181.370 ;
        RECT 30.445 180.570 30.615 181.710 ;
        RECT 30.785 180.570 31.120 181.540 ;
        RECT 31.385 180.780 31.555 181.540 ;
        RECT 31.735 180.950 32.065 181.710 ;
        RECT 31.385 180.610 32.050 180.780 ;
        RECT 32.235 180.635 32.505 181.540 ;
        RECT 30.105 180.070 30.300 180.400 ;
        RECT 30.525 180.070 30.780 180.400 ;
        RECT 30.525 179.900 30.695 180.070 ;
        RECT 30.950 179.900 31.120 180.570 ;
        RECT 31.880 180.465 32.050 180.610 ;
        RECT 31.315 180.060 31.645 180.430 ;
        RECT 31.880 180.135 32.165 180.465 ;
        RECT 29.765 179.730 30.695 179.900 ;
        RECT 29.765 179.695 29.940 179.730 ;
        RECT 28.945 179.500 29.225 179.670 ;
        RECT 28.945 179.330 29.220 179.500 ;
        RECT 29.410 179.330 29.940 179.695 ;
        RECT 30.365 179.160 30.695 179.560 ;
        RECT 30.865 179.330 31.120 179.900 ;
        RECT 31.880 179.880 32.050 180.135 ;
        RECT 31.385 179.710 32.050 179.880 ;
        RECT 32.335 179.835 32.505 180.635 ;
        RECT 32.675 180.620 34.345 181.710 ;
        RECT 34.720 180.740 35.050 181.540 ;
        RECT 35.220 180.910 35.550 181.710 ;
        RECT 35.850 180.740 36.180 181.540 ;
        RECT 36.825 180.910 37.075 181.710 ;
        RECT 32.675 180.100 33.425 180.620 ;
        RECT 34.720 180.570 37.155 180.740 ;
        RECT 37.345 180.570 37.515 181.710 ;
        RECT 37.685 180.570 38.025 181.540 ;
        RECT 33.595 179.930 34.345 180.450 ;
        RECT 34.515 180.150 34.865 180.400 ;
        RECT 35.050 179.940 35.220 180.570 ;
        RECT 35.390 180.150 35.720 180.350 ;
        RECT 35.890 180.150 36.220 180.350 ;
        RECT 36.390 180.150 36.810 180.350 ;
        RECT 36.985 180.320 37.155 180.570 ;
        RECT 36.985 180.150 37.680 180.320 ;
        RECT 31.385 179.330 31.555 179.710 ;
        RECT 31.735 179.160 32.065 179.540 ;
        RECT 32.245 179.330 32.505 179.835 ;
        RECT 32.675 179.160 34.345 179.930 ;
        RECT 34.720 179.330 35.220 179.940 ;
        RECT 35.850 179.810 37.075 179.980 ;
        RECT 37.850 179.960 38.025 180.570 ;
        RECT 38.195 180.545 38.485 181.710 ;
        RECT 38.655 180.620 39.865 181.710 ;
        RECT 38.655 180.080 39.175 180.620 ;
        RECT 40.095 180.570 40.305 181.710 ;
        RECT 40.475 180.560 40.805 181.540 ;
        RECT 40.975 180.570 41.205 181.710 ;
        RECT 41.530 181.080 41.815 181.540 ;
        RECT 41.985 181.250 42.255 181.710 ;
        RECT 41.530 180.860 42.485 181.080 ;
        RECT 35.850 179.330 36.180 179.810 ;
        RECT 36.350 179.160 36.575 179.620 ;
        RECT 36.745 179.330 37.075 179.810 ;
        RECT 37.265 179.160 37.515 179.960 ;
        RECT 37.685 179.330 38.025 179.960 ;
        RECT 39.345 179.910 39.865 180.450 ;
        RECT 38.195 179.160 38.485 179.885 ;
        RECT 38.655 179.160 39.865 179.910 ;
        RECT 40.095 179.160 40.305 179.980 ;
        RECT 40.475 179.960 40.725 180.560 ;
        RECT 40.895 180.150 41.225 180.400 ;
        RECT 41.415 180.130 42.105 180.690 ;
        RECT 40.475 179.330 40.805 179.960 ;
        RECT 40.975 179.160 41.205 179.980 ;
        RECT 42.275 179.960 42.485 180.860 ;
        RECT 41.530 179.790 42.485 179.960 ;
        RECT 42.655 180.690 43.055 181.540 ;
        RECT 43.245 181.080 43.525 181.540 ;
        RECT 44.045 181.250 44.370 181.710 ;
        RECT 43.245 180.860 44.370 181.080 ;
        RECT 42.655 180.130 43.750 180.690 ;
        RECT 43.920 180.400 44.370 180.860 ;
        RECT 44.540 180.570 44.925 181.540 ;
        RECT 41.530 179.330 41.815 179.790 ;
        RECT 41.985 179.160 42.255 179.620 ;
        RECT 42.655 179.330 43.055 180.130 ;
        RECT 43.920 180.070 44.475 180.400 ;
        RECT 43.920 179.960 44.370 180.070 ;
        RECT 43.245 179.790 44.370 179.960 ;
        RECT 44.645 179.900 44.925 180.570 ;
        RECT 43.245 179.330 43.525 179.790 ;
        RECT 44.045 179.160 44.370 179.620 ;
        RECT 44.540 179.330 44.925 179.900 ;
        RECT 45.560 180.520 45.815 181.400 ;
        RECT 45.985 180.570 46.290 181.710 ;
        RECT 46.630 181.330 46.960 181.710 ;
        RECT 47.140 181.160 47.310 181.450 ;
        RECT 47.480 181.250 47.730 181.710 ;
        RECT 46.510 180.990 47.310 181.160 ;
        RECT 47.900 181.200 48.770 181.540 ;
        RECT 45.560 179.870 45.770 180.520 ;
        RECT 46.510 180.400 46.680 180.990 ;
        RECT 47.900 180.820 48.070 181.200 ;
        RECT 49.005 181.080 49.175 181.540 ;
        RECT 49.345 181.250 49.715 181.710 ;
        RECT 50.010 181.110 50.180 181.450 ;
        RECT 50.350 181.280 50.680 181.710 ;
        RECT 50.915 181.110 51.085 181.450 ;
        RECT 46.850 180.650 48.070 180.820 ;
        RECT 48.240 180.740 48.700 181.030 ;
        RECT 49.005 180.910 49.565 181.080 ;
        RECT 50.010 180.940 51.085 181.110 ;
        RECT 51.255 181.210 51.935 181.540 ;
        RECT 52.150 181.210 52.400 181.540 ;
        RECT 52.570 181.250 52.820 181.710 ;
        RECT 49.395 180.770 49.565 180.910 ;
        RECT 48.240 180.730 49.205 180.740 ;
        RECT 47.900 180.560 48.070 180.650 ;
        RECT 48.530 180.570 49.205 180.730 ;
        RECT 45.940 180.370 46.680 180.400 ;
        RECT 45.940 180.070 46.855 180.370 ;
        RECT 46.530 179.895 46.855 180.070 ;
        RECT 45.560 179.340 45.815 179.870 ;
        RECT 45.985 179.160 46.290 179.620 ;
        RECT 46.535 179.540 46.855 179.895 ;
        RECT 47.025 180.110 47.565 180.480 ;
        RECT 47.900 180.390 48.305 180.560 ;
        RECT 47.025 179.710 47.265 180.110 ;
        RECT 47.745 179.940 47.965 180.220 ;
        RECT 47.435 179.770 47.965 179.940 ;
        RECT 47.435 179.540 47.605 179.770 ;
        RECT 48.135 179.610 48.305 180.390 ;
        RECT 48.475 179.780 48.825 180.400 ;
        RECT 48.995 179.780 49.205 180.570 ;
        RECT 49.395 180.600 50.895 180.770 ;
        RECT 49.395 179.910 49.565 180.600 ;
        RECT 51.255 180.430 51.425 181.210 ;
        RECT 52.230 181.080 52.400 181.210 ;
        RECT 49.735 180.260 51.425 180.430 ;
        RECT 51.595 180.650 52.060 181.040 ;
        RECT 52.230 180.910 52.625 181.080 ;
        RECT 49.735 180.080 49.905 180.260 ;
        RECT 46.535 179.370 47.605 179.540 ;
        RECT 47.775 179.160 47.965 179.600 ;
        RECT 48.135 179.330 49.085 179.610 ;
        RECT 49.395 179.520 49.655 179.910 ;
        RECT 50.075 179.840 50.865 180.090 ;
        RECT 49.305 179.350 49.655 179.520 ;
        RECT 49.865 179.160 50.195 179.620 ;
        RECT 51.070 179.550 51.240 180.260 ;
        RECT 51.595 180.060 51.765 180.650 ;
        RECT 51.410 179.840 51.765 180.060 ;
        RECT 51.935 179.840 52.285 180.460 ;
        RECT 52.455 179.550 52.625 180.910 ;
        RECT 52.990 180.740 53.315 181.525 ;
        RECT 52.795 179.690 53.255 180.740 ;
        RECT 51.070 179.380 51.925 179.550 ;
        RECT 52.130 179.380 52.625 179.550 ;
        RECT 52.795 179.160 53.125 179.520 ;
        RECT 53.485 179.420 53.655 181.540 ;
        RECT 53.825 181.210 54.155 181.710 ;
        RECT 54.325 181.040 54.580 181.540 ;
        RECT 53.830 180.870 54.580 181.040 ;
        RECT 53.830 179.880 54.060 180.870 ;
        RECT 54.230 180.050 54.580 180.700 ;
        RECT 55.675 180.620 59.185 181.710 ;
        RECT 55.675 180.100 57.365 180.620 ;
        RECT 59.395 180.570 59.625 181.710 ;
        RECT 59.795 180.560 60.125 181.540 ;
        RECT 60.295 180.570 60.505 181.710 ;
        RECT 61.445 181.260 61.775 181.710 ;
        RECT 60.735 180.870 63.345 181.080 ;
        RECT 57.535 179.930 59.185 180.450 ;
        RECT 59.375 180.150 59.705 180.400 ;
        RECT 53.830 179.710 54.580 179.880 ;
        RECT 53.825 179.160 54.155 179.540 ;
        RECT 54.325 179.420 54.580 179.710 ;
        RECT 55.675 179.160 59.185 179.930 ;
        RECT 59.395 179.160 59.625 179.980 ;
        RECT 59.875 179.960 60.125 180.560 ;
        RECT 59.795 179.330 60.125 179.960 ;
        RECT 60.295 179.160 60.505 179.980 ;
        RECT 60.735 179.900 60.905 180.870 ;
        RECT 61.075 180.070 61.425 180.690 ;
        RECT 61.595 180.070 61.915 180.690 ;
        RECT 62.085 180.070 62.415 180.690 ;
        RECT 62.585 180.070 62.885 180.690 ;
        RECT 63.125 180.070 63.345 180.870 ;
        RECT 63.525 179.900 63.785 181.525 ;
        RECT 63.955 180.545 64.245 181.710 ;
        RECT 64.415 180.620 65.625 181.710 ;
        RECT 65.795 180.620 69.305 181.710 ;
        RECT 69.475 180.740 69.785 181.540 ;
        RECT 69.955 180.910 70.265 181.710 ;
        RECT 70.435 181.080 70.695 181.540 ;
        RECT 70.865 181.250 71.120 181.710 ;
        RECT 71.295 181.080 71.555 181.540 ;
        RECT 70.435 180.910 71.555 181.080 ;
        RECT 64.415 180.080 64.935 180.620 ;
        RECT 65.105 179.910 65.625 180.450 ;
        RECT 65.795 180.100 67.485 180.620 ;
        RECT 69.475 180.570 70.505 180.740 ;
        RECT 67.655 179.930 69.305 180.450 ;
        RECT 60.735 179.730 61.210 179.900 ;
        RECT 61.040 179.480 61.210 179.730 ;
        RECT 61.445 179.160 61.775 179.900 ;
        RECT 61.945 179.730 63.785 179.900 ;
        RECT 61.945 179.385 62.145 179.730 ;
        RECT 62.315 179.160 62.645 179.560 ;
        RECT 62.815 179.375 63.015 179.730 ;
        RECT 63.185 179.160 63.515 179.555 ;
        RECT 63.955 179.160 64.245 179.885 ;
        RECT 64.415 179.160 65.625 179.910 ;
        RECT 65.795 179.160 69.305 179.930 ;
        RECT 69.475 179.660 69.645 180.570 ;
        RECT 69.815 179.830 70.165 180.400 ;
        RECT 70.335 180.320 70.505 180.570 ;
        RECT 71.295 180.660 71.555 180.910 ;
        RECT 71.725 180.840 72.010 181.710 ;
        RECT 71.295 180.490 72.050 180.660 ;
        RECT 70.335 180.150 71.475 180.320 ;
        RECT 71.645 179.980 72.050 180.490 ;
        RECT 72.695 180.620 74.365 181.710 ;
        RECT 72.695 180.100 73.445 180.620 ;
        RECT 74.540 180.520 74.795 181.400 ;
        RECT 74.965 180.570 75.270 181.710 ;
        RECT 75.610 181.330 75.940 181.710 ;
        RECT 76.120 181.160 76.290 181.450 ;
        RECT 76.460 181.250 76.710 181.710 ;
        RECT 75.490 180.990 76.290 181.160 ;
        RECT 76.880 181.200 77.750 181.540 ;
        RECT 70.400 179.810 72.050 179.980 ;
        RECT 73.615 179.930 74.365 180.450 ;
        RECT 69.475 179.330 69.775 179.660 ;
        RECT 69.945 179.160 70.220 179.640 ;
        RECT 70.400 179.420 70.695 179.810 ;
        RECT 70.865 179.160 71.120 179.640 ;
        RECT 71.295 179.420 71.555 179.810 ;
        RECT 71.725 179.160 72.005 179.640 ;
        RECT 72.695 179.160 74.365 179.930 ;
        RECT 74.540 179.870 74.750 180.520 ;
        RECT 75.490 180.400 75.660 180.990 ;
        RECT 76.880 180.820 77.050 181.200 ;
        RECT 77.985 181.080 78.155 181.540 ;
        RECT 78.325 181.250 78.695 181.710 ;
        RECT 78.990 181.110 79.160 181.450 ;
        RECT 79.330 181.280 79.660 181.710 ;
        RECT 79.895 181.110 80.065 181.450 ;
        RECT 75.830 180.650 77.050 180.820 ;
        RECT 77.220 180.740 77.680 181.030 ;
        RECT 77.985 180.910 78.545 181.080 ;
        RECT 78.990 180.940 80.065 181.110 ;
        RECT 80.235 181.210 80.915 181.540 ;
        RECT 81.130 181.210 81.380 181.540 ;
        RECT 81.550 181.250 81.800 181.710 ;
        RECT 78.375 180.770 78.545 180.910 ;
        RECT 77.220 180.730 78.185 180.740 ;
        RECT 76.880 180.560 77.050 180.650 ;
        RECT 77.510 180.570 78.185 180.730 ;
        RECT 74.920 180.370 75.660 180.400 ;
        RECT 74.920 180.070 75.835 180.370 ;
        RECT 75.510 179.895 75.835 180.070 ;
        RECT 74.540 179.340 74.795 179.870 ;
        RECT 74.965 179.160 75.270 179.620 ;
        RECT 75.515 179.540 75.835 179.895 ;
        RECT 76.005 180.110 76.545 180.480 ;
        RECT 76.880 180.390 77.285 180.560 ;
        RECT 76.005 179.710 76.245 180.110 ;
        RECT 76.725 179.940 76.945 180.220 ;
        RECT 76.415 179.770 76.945 179.940 ;
        RECT 76.415 179.540 76.585 179.770 ;
        RECT 77.115 179.610 77.285 180.390 ;
        RECT 77.455 179.780 77.805 180.400 ;
        RECT 77.975 179.780 78.185 180.570 ;
        RECT 78.375 180.600 79.875 180.770 ;
        RECT 78.375 179.910 78.545 180.600 ;
        RECT 80.235 180.430 80.405 181.210 ;
        RECT 81.210 181.080 81.380 181.210 ;
        RECT 78.715 180.260 80.405 180.430 ;
        RECT 80.575 180.650 81.040 181.040 ;
        RECT 81.210 180.910 81.605 181.080 ;
        RECT 78.715 180.080 78.885 180.260 ;
        RECT 75.515 179.370 76.585 179.540 ;
        RECT 76.755 179.160 76.945 179.600 ;
        RECT 77.115 179.330 78.065 179.610 ;
        RECT 78.375 179.520 78.635 179.910 ;
        RECT 79.055 179.840 79.845 180.090 ;
        RECT 78.285 179.350 78.635 179.520 ;
        RECT 78.845 179.160 79.175 179.620 ;
        RECT 80.050 179.550 80.220 180.260 ;
        RECT 80.575 180.060 80.745 180.650 ;
        RECT 80.390 179.840 80.745 180.060 ;
        RECT 80.915 179.840 81.265 180.460 ;
        RECT 81.435 179.550 81.605 180.910 ;
        RECT 81.970 180.740 82.295 181.525 ;
        RECT 81.775 179.690 82.235 180.740 ;
        RECT 80.050 179.380 80.905 179.550 ;
        RECT 81.110 179.380 81.605 179.550 ;
        RECT 81.775 179.160 82.105 179.520 ;
        RECT 82.465 179.420 82.635 181.540 ;
        RECT 82.805 181.210 83.135 181.710 ;
        RECT 83.305 181.040 83.560 181.540 ;
        RECT 82.810 180.870 83.560 181.040 ;
        RECT 82.810 179.880 83.040 180.870 ;
        RECT 83.210 180.050 83.560 180.700 ;
        RECT 83.735 180.635 84.005 181.540 ;
        RECT 84.175 180.950 84.505 181.710 ;
        RECT 84.685 180.780 84.855 181.540 ;
        RECT 82.810 179.710 83.560 179.880 ;
        RECT 82.805 179.160 83.135 179.540 ;
        RECT 83.305 179.420 83.560 179.710 ;
        RECT 83.735 179.835 83.905 180.635 ;
        RECT 84.190 180.610 84.855 180.780 ;
        RECT 84.190 180.465 84.360 180.610 ;
        RECT 84.075 180.135 84.360 180.465 ;
        RECT 86.035 180.570 86.420 181.540 ;
        RECT 86.590 181.250 86.915 181.710 ;
        RECT 87.435 181.080 87.715 181.540 ;
        RECT 86.590 180.860 87.715 181.080 ;
        RECT 84.190 179.880 84.360 180.135 ;
        RECT 84.595 180.060 84.925 180.430 ;
        RECT 86.035 179.900 86.315 180.570 ;
        RECT 86.590 180.400 87.040 180.860 ;
        RECT 87.905 180.690 88.305 181.540 ;
        RECT 88.705 181.250 88.975 181.710 ;
        RECT 89.145 181.080 89.430 181.540 ;
        RECT 86.485 180.070 87.040 180.400 ;
        RECT 87.210 180.130 88.305 180.690 ;
        RECT 86.590 179.960 87.040 180.070 ;
        RECT 83.735 179.330 83.995 179.835 ;
        RECT 84.190 179.710 84.855 179.880 ;
        RECT 84.175 179.160 84.505 179.540 ;
        RECT 84.685 179.330 84.855 179.710 ;
        RECT 86.035 179.330 86.420 179.900 ;
        RECT 86.590 179.790 87.715 179.960 ;
        RECT 86.590 179.160 86.915 179.620 ;
        RECT 87.435 179.330 87.715 179.790 ;
        RECT 87.905 179.330 88.305 180.130 ;
        RECT 88.475 180.860 89.430 181.080 ;
        RECT 88.475 179.960 88.685 180.860 ;
        RECT 88.855 180.130 89.545 180.690 ;
        RECT 89.715 180.545 90.005 181.710 ;
        RECT 90.235 180.570 90.445 181.710 ;
        RECT 90.615 180.560 90.945 181.540 ;
        RECT 91.115 180.570 91.345 181.710 ;
        RECT 91.555 180.635 91.825 181.540 ;
        RECT 91.995 180.950 92.325 181.710 ;
        RECT 92.505 180.780 92.675 181.540 ;
        RECT 88.475 179.790 89.430 179.960 ;
        RECT 88.705 179.160 88.975 179.620 ;
        RECT 89.145 179.330 89.430 179.790 ;
        RECT 89.715 179.160 90.005 179.885 ;
        RECT 90.235 179.160 90.445 179.980 ;
        RECT 90.615 179.960 90.865 180.560 ;
        RECT 91.035 180.150 91.365 180.400 ;
        RECT 90.615 179.330 90.945 179.960 ;
        RECT 91.115 179.160 91.345 179.980 ;
        RECT 91.555 179.835 91.725 180.635 ;
        RECT 92.010 180.610 92.675 180.780 ;
        RECT 92.010 180.465 92.180 180.610 ;
        RECT 91.895 180.135 92.180 180.465 ;
        RECT 92.935 180.570 93.320 181.540 ;
        RECT 93.490 181.250 93.815 181.710 ;
        RECT 94.335 181.080 94.615 181.540 ;
        RECT 93.490 180.860 94.615 181.080 ;
        RECT 92.010 179.880 92.180 180.135 ;
        RECT 92.415 180.060 92.745 180.430 ;
        RECT 92.935 179.900 93.215 180.570 ;
        RECT 93.490 180.400 93.940 180.860 ;
        RECT 94.805 180.690 95.205 181.540 ;
        RECT 95.605 181.250 95.875 181.710 ;
        RECT 96.045 181.080 96.330 181.540 ;
        RECT 93.385 180.070 93.940 180.400 ;
        RECT 94.110 180.130 95.205 180.690 ;
        RECT 93.490 179.960 93.940 180.070 ;
        RECT 91.555 179.330 91.815 179.835 ;
        RECT 92.010 179.710 92.675 179.880 ;
        RECT 91.995 179.160 92.325 179.540 ;
        RECT 92.505 179.330 92.675 179.710 ;
        RECT 92.935 179.330 93.320 179.900 ;
        RECT 93.490 179.790 94.615 179.960 ;
        RECT 93.490 179.160 93.815 179.620 ;
        RECT 94.335 179.330 94.615 179.790 ;
        RECT 94.805 179.330 95.205 180.130 ;
        RECT 95.375 180.860 96.330 181.080 ;
        RECT 95.375 179.960 95.585 180.860 ;
        RECT 95.755 180.130 96.445 180.690 ;
        RECT 97.075 180.620 98.745 181.710 ;
        RECT 97.075 180.100 97.825 180.620 ;
        RECT 98.920 180.520 99.175 181.400 ;
        RECT 99.345 180.570 99.650 181.710 ;
        RECT 99.990 181.330 100.320 181.710 ;
        RECT 100.500 181.160 100.670 181.450 ;
        RECT 100.840 181.250 101.090 181.710 ;
        RECT 99.870 180.990 100.670 181.160 ;
        RECT 101.260 181.200 102.130 181.540 ;
        RECT 95.375 179.790 96.330 179.960 ;
        RECT 97.995 179.930 98.745 180.450 ;
        RECT 95.605 179.160 95.875 179.620 ;
        RECT 96.045 179.330 96.330 179.790 ;
        RECT 97.075 179.160 98.745 179.930 ;
        RECT 98.920 179.870 99.130 180.520 ;
        RECT 99.870 180.400 100.040 180.990 ;
        RECT 101.260 180.820 101.430 181.200 ;
        RECT 102.365 181.080 102.535 181.540 ;
        RECT 102.705 181.250 103.075 181.710 ;
        RECT 103.370 181.110 103.540 181.450 ;
        RECT 103.710 181.280 104.040 181.710 ;
        RECT 104.275 181.110 104.445 181.450 ;
        RECT 100.210 180.650 101.430 180.820 ;
        RECT 101.600 180.740 102.060 181.030 ;
        RECT 102.365 180.910 102.925 181.080 ;
        RECT 103.370 180.940 104.445 181.110 ;
        RECT 104.615 181.210 105.295 181.540 ;
        RECT 105.510 181.210 105.760 181.540 ;
        RECT 105.930 181.250 106.180 181.710 ;
        RECT 102.755 180.770 102.925 180.910 ;
        RECT 101.600 180.730 102.565 180.740 ;
        RECT 101.260 180.560 101.430 180.650 ;
        RECT 101.890 180.570 102.565 180.730 ;
        RECT 99.300 180.370 100.040 180.400 ;
        RECT 99.300 180.070 100.215 180.370 ;
        RECT 99.890 179.895 100.215 180.070 ;
        RECT 98.920 179.340 99.175 179.870 ;
        RECT 99.345 179.160 99.650 179.620 ;
        RECT 99.895 179.540 100.215 179.895 ;
        RECT 100.385 180.110 100.925 180.480 ;
        RECT 101.260 180.390 101.665 180.560 ;
        RECT 100.385 179.710 100.625 180.110 ;
        RECT 101.105 179.940 101.325 180.220 ;
        RECT 100.795 179.770 101.325 179.940 ;
        RECT 100.795 179.540 100.965 179.770 ;
        RECT 101.495 179.610 101.665 180.390 ;
        RECT 101.835 179.780 102.185 180.400 ;
        RECT 102.355 179.780 102.565 180.570 ;
        RECT 102.755 180.600 104.255 180.770 ;
        RECT 102.755 179.910 102.925 180.600 ;
        RECT 104.615 180.430 104.785 181.210 ;
        RECT 105.590 181.080 105.760 181.210 ;
        RECT 103.095 180.260 104.785 180.430 ;
        RECT 104.955 180.650 105.420 181.040 ;
        RECT 105.590 180.910 105.985 181.080 ;
        RECT 103.095 180.080 103.265 180.260 ;
        RECT 99.895 179.370 100.965 179.540 ;
        RECT 101.135 179.160 101.325 179.600 ;
        RECT 101.495 179.330 102.445 179.610 ;
        RECT 102.755 179.520 103.015 179.910 ;
        RECT 103.435 179.840 104.225 180.090 ;
        RECT 102.665 179.350 103.015 179.520 ;
        RECT 103.225 179.160 103.555 179.620 ;
        RECT 104.430 179.550 104.600 180.260 ;
        RECT 104.955 180.060 105.125 180.650 ;
        RECT 104.770 179.840 105.125 180.060 ;
        RECT 105.295 179.840 105.645 180.460 ;
        RECT 105.815 179.550 105.985 180.910 ;
        RECT 106.350 180.740 106.675 181.525 ;
        RECT 106.155 179.690 106.615 180.740 ;
        RECT 104.430 179.380 105.285 179.550 ;
        RECT 105.490 179.380 105.985 179.550 ;
        RECT 106.155 179.160 106.485 179.520 ;
        RECT 106.845 179.420 107.015 181.540 ;
        RECT 107.185 181.210 107.515 181.710 ;
        RECT 107.685 181.040 107.940 181.540 ;
        RECT 107.190 180.870 107.940 181.040 ;
        RECT 107.190 179.880 107.420 180.870 ;
        RECT 107.590 180.050 107.940 180.700 ;
        RECT 108.155 180.570 108.385 181.710 ;
        RECT 108.555 180.560 108.885 181.540 ;
        RECT 109.055 180.570 109.265 181.710 ;
        RECT 110.505 180.780 110.675 181.540 ;
        RECT 110.855 180.950 111.185 181.710 ;
        RECT 110.505 180.610 111.170 180.780 ;
        RECT 111.355 180.635 111.625 181.540 ;
        RECT 108.135 180.150 108.465 180.400 ;
        RECT 107.190 179.710 107.940 179.880 ;
        RECT 107.185 179.160 107.515 179.540 ;
        RECT 107.685 179.420 107.940 179.710 ;
        RECT 108.155 179.160 108.385 179.980 ;
        RECT 108.635 179.960 108.885 180.560 ;
        RECT 111.000 180.465 111.170 180.610 ;
        RECT 110.435 180.060 110.765 180.430 ;
        RECT 111.000 180.135 111.285 180.465 ;
        RECT 108.555 179.330 108.885 179.960 ;
        RECT 109.055 179.160 109.265 179.980 ;
        RECT 111.000 179.880 111.170 180.135 ;
        RECT 110.505 179.710 111.170 179.880 ;
        RECT 111.455 179.835 111.625 180.635 ;
        RECT 111.795 180.620 114.385 181.710 ;
        RECT 114.555 180.620 115.765 181.710 ;
        RECT 111.795 180.100 113.005 180.620 ;
        RECT 113.175 179.930 114.385 180.450 ;
        RECT 114.555 180.080 115.075 180.620 ;
        RECT 110.505 179.330 110.675 179.710 ;
        RECT 110.855 179.160 111.185 179.540 ;
        RECT 111.365 179.330 111.625 179.835 ;
        RECT 111.795 179.160 114.385 179.930 ;
        RECT 115.245 179.910 115.765 180.450 ;
        RECT 114.555 179.160 115.765 179.910 ;
        RECT 10.510 178.990 115.850 179.160 ;
        RECT 10.595 178.240 11.805 178.990 ;
        RECT 10.595 177.700 11.115 178.240 ;
        RECT 11.975 178.220 15.485 178.990 ;
        RECT 11.285 177.530 11.805 178.070 ;
        RECT 10.595 176.440 11.805 177.530 ;
        RECT 11.975 177.530 13.665 178.050 ;
        RECT 13.835 177.700 15.485 178.220 ;
        RECT 15.770 178.360 16.055 178.820 ;
        RECT 16.225 178.530 16.495 178.990 ;
        RECT 15.770 178.190 16.725 178.360 ;
        RECT 11.975 176.440 15.485 177.530 ;
        RECT 15.655 177.460 16.345 178.020 ;
        RECT 16.515 177.290 16.725 178.190 ;
        RECT 15.770 177.070 16.725 177.290 ;
        RECT 16.895 178.020 17.295 178.820 ;
        RECT 17.485 178.360 17.765 178.820 ;
        RECT 18.285 178.530 18.610 178.990 ;
        RECT 17.485 178.190 18.610 178.360 ;
        RECT 18.780 178.250 19.165 178.820 ;
        RECT 18.160 178.080 18.610 178.190 ;
        RECT 16.895 177.460 17.990 178.020 ;
        RECT 18.160 177.750 18.715 178.080 ;
        RECT 15.770 176.610 16.055 177.070 ;
        RECT 16.225 176.440 16.495 176.900 ;
        RECT 16.895 176.610 17.295 177.460 ;
        RECT 18.160 177.290 18.610 177.750 ;
        RECT 18.885 177.580 19.165 178.250 ;
        RECT 19.855 178.170 20.065 178.990 ;
        RECT 20.235 178.190 20.565 178.820 ;
        RECT 20.235 177.590 20.485 178.190 ;
        RECT 20.735 178.170 20.965 178.990 ;
        RECT 21.450 178.180 21.695 178.785 ;
        RECT 21.915 178.455 22.425 178.990 ;
        RECT 21.175 178.010 22.405 178.180 ;
        RECT 20.655 177.750 20.985 178.000 ;
        RECT 17.485 177.070 18.610 177.290 ;
        RECT 17.485 176.610 17.765 177.070 ;
        RECT 18.285 176.440 18.610 176.900 ;
        RECT 18.780 176.610 19.165 177.580 ;
        RECT 19.855 176.440 20.065 177.580 ;
        RECT 20.235 176.610 20.565 177.590 ;
        RECT 20.735 176.440 20.965 177.580 ;
        RECT 21.175 177.200 21.515 178.010 ;
        RECT 21.685 177.445 22.435 177.635 ;
        RECT 21.175 176.790 21.690 177.200 ;
        RECT 21.925 176.440 22.095 177.200 ;
        RECT 22.265 176.780 22.435 177.445 ;
        RECT 22.605 177.460 22.795 178.820 ;
        RECT 22.965 178.310 23.240 178.820 ;
        RECT 23.430 178.455 23.960 178.820 ;
        RECT 24.385 178.590 24.715 178.990 ;
        RECT 23.785 178.420 23.960 178.455 ;
        RECT 22.965 178.140 23.245 178.310 ;
        RECT 22.965 177.660 23.240 178.140 ;
        RECT 23.445 177.460 23.615 178.260 ;
        RECT 22.605 177.290 23.615 177.460 ;
        RECT 23.785 178.250 24.715 178.420 ;
        RECT 24.885 178.250 25.140 178.820 ;
        RECT 25.315 178.265 25.605 178.990 ;
        RECT 23.785 177.120 23.955 178.250 ;
        RECT 24.545 178.080 24.715 178.250 ;
        RECT 22.830 176.950 23.955 177.120 ;
        RECT 24.125 177.750 24.320 178.080 ;
        RECT 24.545 177.750 24.800 178.080 ;
        RECT 24.125 176.780 24.295 177.750 ;
        RECT 24.970 177.580 25.140 178.250 ;
        RECT 26.900 178.210 27.400 178.820 ;
        RECT 26.695 177.750 27.045 178.000 ;
        RECT 22.265 176.610 24.295 176.780 ;
        RECT 24.465 176.440 24.635 177.580 ;
        RECT 24.805 176.610 25.140 177.580 ;
        RECT 25.315 176.440 25.605 177.605 ;
        RECT 27.230 177.580 27.400 178.210 ;
        RECT 28.030 178.340 28.360 178.820 ;
        RECT 28.530 178.530 28.755 178.990 ;
        RECT 28.925 178.340 29.255 178.820 ;
        RECT 28.030 178.170 29.255 178.340 ;
        RECT 29.445 178.190 29.695 178.990 ;
        RECT 29.865 178.190 30.205 178.820 ;
        RECT 27.570 177.800 27.900 178.000 ;
        RECT 28.070 177.800 28.400 178.000 ;
        RECT 28.570 177.800 28.990 178.000 ;
        RECT 29.165 177.830 29.860 178.000 ;
        RECT 29.165 177.580 29.335 177.830 ;
        RECT 30.030 177.580 30.205 178.190 ;
        RECT 26.900 177.410 29.335 177.580 ;
        RECT 26.900 176.610 27.230 177.410 ;
        RECT 27.400 176.440 27.730 177.240 ;
        RECT 28.030 176.610 28.360 177.410 ;
        RECT 29.005 176.440 29.255 177.240 ;
        RECT 29.525 176.440 29.695 177.580 ;
        RECT 29.865 176.610 30.205 177.580 ;
        RECT 30.380 178.250 30.635 178.820 ;
        RECT 30.805 178.590 31.135 178.990 ;
        RECT 31.560 178.455 32.090 178.820 ;
        RECT 32.280 178.650 32.555 178.820 ;
        RECT 32.275 178.480 32.555 178.650 ;
        RECT 31.560 178.420 31.735 178.455 ;
        RECT 30.805 178.250 31.735 178.420 ;
        RECT 30.380 177.580 30.550 178.250 ;
        RECT 30.805 178.080 30.975 178.250 ;
        RECT 30.720 177.750 30.975 178.080 ;
        RECT 31.200 177.750 31.395 178.080 ;
        RECT 30.380 176.610 30.715 177.580 ;
        RECT 30.885 176.440 31.055 177.580 ;
        RECT 31.225 176.780 31.395 177.750 ;
        RECT 31.565 177.120 31.735 178.250 ;
        RECT 31.905 177.460 32.075 178.260 ;
        RECT 32.280 177.660 32.555 178.480 ;
        RECT 32.725 177.460 32.915 178.820 ;
        RECT 33.095 178.455 33.605 178.990 ;
        RECT 33.825 178.180 34.070 178.785 ;
        RECT 34.515 178.240 35.725 178.990 ;
        RECT 33.115 178.010 34.345 178.180 ;
        RECT 31.905 177.290 32.915 177.460 ;
        RECT 33.085 177.445 33.835 177.635 ;
        RECT 31.565 176.950 32.690 177.120 ;
        RECT 33.085 176.780 33.255 177.445 ;
        RECT 34.005 177.200 34.345 178.010 ;
        RECT 31.225 176.610 33.255 176.780 ;
        RECT 33.425 176.440 33.595 177.200 ;
        RECT 33.830 176.790 34.345 177.200 ;
        RECT 34.515 177.530 35.035 178.070 ;
        RECT 35.205 177.700 35.725 178.240 ;
        RECT 36.100 178.210 36.600 178.820 ;
        RECT 35.895 177.750 36.245 178.000 ;
        RECT 36.430 177.580 36.600 178.210 ;
        RECT 37.230 178.340 37.560 178.820 ;
        RECT 37.730 178.530 37.955 178.990 ;
        RECT 38.125 178.340 38.455 178.820 ;
        RECT 37.230 178.170 38.455 178.340 ;
        RECT 38.645 178.190 38.895 178.990 ;
        RECT 39.065 178.190 39.405 178.820 ;
        RECT 39.780 178.210 40.280 178.820 ;
        RECT 36.770 177.800 37.100 178.000 ;
        RECT 37.270 177.800 37.600 178.000 ;
        RECT 37.770 177.800 38.190 178.000 ;
        RECT 38.365 177.830 39.060 178.000 ;
        RECT 38.365 177.580 38.535 177.830 ;
        RECT 39.230 177.580 39.405 178.190 ;
        RECT 39.575 177.750 39.925 178.000 ;
        RECT 40.110 177.580 40.280 178.210 ;
        RECT 40.910 178.340 41.240 178.820 ;
        RECT 41.410 178.530 41.635 178.990 ;
        RECT 41.805 178.340 42.135 178.820 ;
        RECT 40.910 178.170 42.135 178.340 ;
        RECT 42.325 178.190 42.575 178.990 ;
        RECT 42.745 178.190 43.085 178.820 ;
        RECT 43.370 178.360 43.655 178.820 ;
        RECT 43.825 178.530 44.095 178.990 ;
        RECT 43.370 178.190 44.325 178.360 ;
        RECT 40.450 177.800 40.780 178.000 ;
        RECT 40.950 177.800 41.280 178.000 ;
        RECT 41.450 177.800 41.870 178.000 ;
        RECT 42.045 177.830 42.740 178.000 ;
        RECT 42.045 177.580 42.215 177.830 ;
        RECT 42.910 177.580 43.085 178.190 ;
        RECT 34.515 176.440 35.725 177.530 ;
        RECT 36.100 177.410 38.535 177.580 ;
        RECT 36.100 176.610 36.430 177.410 ;
        RECT 36.600 176.440 36.930 177.240 ;
        RECT 37.230 176.610 37.560 177.410 ;
        RECT 38.205 176.440 38.455 177.240 ;
        RECT 38.725 176.440 38.895 177.580 ;
        RECT 39.065 176.610 39.405 177.580 ;
        RECT 39.780 177.410 42.215 177.580 ;
        RECT 39.780 176.610 40.110 177.410 ;
        RECT 40.280 176.440 40.610 177.240 ;
        RECT 40.910 176.610 41.240 177.410 ;
        RECT 41.885 176.440 42.135 177.240 ;
        RECT 42.405 176.440 42.575 177.580 ;
        RECT 42.745 176.610 43.085 177.580 ;
        RECT 43.255 177.460 43.945 178.020 ;
        RECT 44.115 177.290 44.325 178.190 ;
        RECT 43.370 177.070 44.325 177.290 ;
        RECT 44.495 178.020 44.895 178.820 ;
        RECT 45.085 178.360 45.365 178.820 ;
        RECT 45.885 178.530 46.210 178.990 ;
        RECT 45.085 178.190 46.210 178.360 ;
        RECT 46.380 178.250 46.765 178.820 ;
        RECT 45.760 178.080 46.210 178.190 ;
        RECT 44.495 177.460 45.590 178.020 ;
        RECT 45.760 177.750 46.315 178.080 ;
        RECT 43.370 176.610 43.655 177.070 ;
        RECT 43.825 176.440 44.095 176.900 ;
        RECT 44.495 176.610 44.895 177.460 ;
        RECT 45.760 177.290 46.210 177.750 ;
        RECT 46.485 177.580 46.765 178.250 ;
        RECT 47.210 178.180 47.455 178.785 ;
        RECT 47.675 178.455 48.185 178.990 ;
        RECT 45.085 177.070 46.210 177.290 ;
        RECT 45.085 176.610 45.365 177.070 ;
        RECT 45.885 176.440 46.210 176.900 ;
        RECT 46.380 176.610 46.765 177.580 ;
        RECT 46.935 178.010 48.165 178.180 ;
        RECT 46.935 177.200 47.275 178.010 ;
        RECT 47.445 177.445 48.195 177.635 ;
        RECT 46.935 176.790 47.450 177.200 ;
        RECT 47.685 176.440 47.855 177.200 ;
        RECT 48.025 176.780 48.195 177.445 ;
        RECT 48.365 177.460 48.555 178.820 ;
        RECT 48.725 177.970 49.000 178.820 ;
        RECT 49.190 178.455 49.720 178.820 ;
        RECT 50.145 178.590 50.475 178.990 ;
        RECT 49.545 178.420 49.720 178.455 ;
        RECT 48.725 177.800 49.005 177.970 ;
        RECT 48.725 177.660 49.000 177.800 ;
        RECT 49.205 177.460 49.375 178.260 ;
        RECT 48.365 177.290 49.375 177.460 ;
        RECT 49.545 178.250 50.475 178.420 ;
        RECT 50.645 178.250 50.900 178.820 ;
        RECT 51.075 178.265 51.365 178.990 ;
        RECT 49.545 177.120 49.715 178.250 ;
        RECT 50.305 178.080 50.475 178.250 ;
        RECT 48.590 176.950 49.715 177.120 ;
        RECT 49.885 177.750 50.080 178.080 ;
        RECT 50.305 177.750 50.560 178.080 ;
        RECT 49.885 176.780 50.055 177.750 ;
        RECT 50.730 177.580 50.900 178.250 ;
        RECT 51.535 178.250 51.920 178.820 ;
        RECT 52.090 178.530 52.415 178.990 ;
        RECT 52.935 178.360 53.215 178.820 ;
        RECT 48.025 176.610 50.055 176.780 ;
        RECT 50.225 176.440 50.395 177.580 ;
        RECT 50.565 176.610 50.900 177.580 ;
        RECT 51.075 176.440 51.365 177.605 ;
        RECT 51.535 177.580 51.815 178.250 ;
        RECT 52.090 178.190 53.215 178.360 ;
        RECT 52.090 178.080 52.540 178.190 ;
        RECT 51.985 177.750 52.540 178.080 ;
        RECT 53.405 178.020 53.805 178.820 ;
        RECT 54.205 178.530 54.475 178.990 ;
        RECT 54.645 178.360 54.930 178.820 ;
        RECT 55.275 178.510 55.555 178.990 ;
        RECT 51.535 176.610 51.920 177.580 ;
        RECT 52.090 177.290 52.540 177.750 ;
        RECT 52.710 177.460 53.805 178.020 ;
        RECT 52.090 177.070 53.215 177.290 ;
        RECT 52.090 176.440 52.415 176.900 ;
        RECT 52.935 176.610 53.215 177.070 ;
        RECT 53.405 176.610 53.805 177.460 ;
        RECT 53.975 178.190 54.930 178.360 ;
        RECT 55.725 178.340 55.985 178.730 ;
        RECT 56.160 178.510 56.415 178.990 ;
        RECT 56.585 178.340 56.880 178.730 ;
        RECT 57.060 178.510 57.335 178.990 ;
        RECT 57.505 178.490 57.805 178.820 ;
        RECT 53.975 177.290 54.185 178.190 ;
        RECT 55.230 178.170 56.880 178.340 ;
        RECT 54.355 177.460 55.045 178.020 ;
        RECT 55.230 177.660 55.635 178.170 ;
        RECT 55.805 177.830 56.945 178.000 ;
        RECT 55.230 177.490 55.985 177.660 ;
        RECT 53.975 177.070 54.930 177.290 ;
        RECT 54.205 176.440 54.475 176.900 ;
        RECT 54.645 176.610 54.930 177.070 ;
        RECT 55.270 176.440 55.555 177.310 ;
        RECT 55.725 177.240 55.985 177.490 ;
        RECT 56.775 177.580 56.945 177.830 ;
        RECT 57.115 177.750 57.465 178.320 ;
        RECT 57.635 177.580 57.805 178.490 ;
        RECT 58.065 178.340 58.235 178.820 ;
        RECT 58.415 178.510 58.655 178.990 ;
        RECT 58.905 178.340 59.075 178.820 ;
        RECT 59.245 178.510 59.575 178.990 ;
        RECT 59.745 178.340 59.915 178.820 ;
        RECT 58.065 178.170 58.700 178.340 ;
        RECT 58.905 178.170 59.915 178.340 ;
        RECT 60.085 178.190 60.415 178.990 ;
        RECT 60.825 178.440 60.995 178.820 ;
        RECT 61.210 178.610 61.540 178.990 ;
        RECT 60.825 178.270 61.540 178.440 ;
        RECT 58.530 178.000 58.700 178.170 ;
        RECT 57.980 177.760 58.360 178.000 ;
        RECT 58.530 177.830 59.030 178.000 ;
        RECT 58.530 177.590 58.700 177.830 ;
        RECT 59.420 177.630 59.915 178.170 ;
        RECT 60.735 177.720 61.090 178.090 ;
        RECT 61.370 178.080 61.540 178.270 ;
        RECT 61.710 178.245 61.965 178.820 ;
        RECT 61.370 177.750 61.625 178.080 ;
        RECT 56.775 177.410 57.805 177.580 ;
        RECT 55.725 177.070 56.845 177.240 ;
        RECT 55.725 176.610 55.985 177.070 ;
        RECT 56.160 176.440 56.415 176.900 ;
        RECT 56.585 176.610 56.845 177.070 ;
        RECT 57.015 176.440 57.325 177.240 ;
        RECT 57.495 176.610 57.805 177.410 ;
        RECT 57.985 177.420 58.700 177.590 ;
        RECT 58.905 177.460 59.915 177.630 ;
        RECT 57.985 176.610 58.315 177.420 ;
        RECT 58.485 176.440 58.725 177.240 ;
        RECT 58.905 176.610 59.075 177.460 ;
        RECT 59.245 176.440 59.575 177.240 ;
        RECT 59.745 176.610 59.915 177.460 ;
        RECT 60.085 176.440 60.415 177.590 ;
        RECT 61.370 177.540 61.540 177.750 ;
        RECT 60.825 177.370 61.540 177.540 ;
        RECT 61.795 177.515 61.965 178.245 ;
        RECT 62.140 178.150 62.400 178.990 ;
        RECT 62.665 178.440 62.835 178.820 ;
        RECT 63.050 178.610 63.380 178.990 ;
        RECT 62.665 178.270 63.380 178.440 ;
        RECT 62.575 177.720 62.930 178.090 ;
        RECT 63.210 178.080 63.380 178.270 ;
        RECT 63.550 178.245 63.805 178.820 ;
        RECT 63.210 177.750 63.465 178.080 ;
        RECT 60.825 176.610 60.995 177.370 ;
        RECT 61.210 176.440 61.540 177.200 ;
        RECT 61.710 176.610 61.965 177.515 ;
        RECT 62.140 176.440 62.400 177.590 ;
        RECT 63.210 177.540 63.380 177.750 ;
        RECT 62.665 177.370 63.380 177.540 ;
        RECT 63.635 177.515 63.805 178.245 ;
        RECT 63.980 178.150 64.240 178.990 ;
        RECT 64.425 178.460 64.755 178.820 ;
        RECT 64.925 178.630 65.255 178.990 ;
        RECT 65.455 178.460 65.785 178.820 ;
        RECT 64.425 178.250 65.785 178.460 ;
        RECT 66.295 178.230 67.005 178.820 ;
        RECT 67.265 178.440 67.435 178.820 ;
        RECT 67.650 178.610 67.980 178.990 ;
        RECT 67.265 178.270 67.980 178.440 ;
        RECT 64.415 177.750 64.725 178.080 ;
        RECT 64.935 177.750 65.310 178.080 ;
        RECT 65.630 177.750 66.125 178.080 ;
        RECT 62.665 176.610 62.835 177.370 ;
        RECT 63.050 176.440 63.380 177.200 ;
        RECT 63.550 176.610 63.805 177.515 ;
        RECT 63.980 176.440 64.240 177.590 ;
        RECT 64.425 176.440 64.755 177.500 ;
        RECT 64.935 176.780 65.105 177.750 ;
        RECT 65.275 177.260 65.605 177.480 ;
        RECT 65.800 177.460 66.125 177.750 ;
        RECT 66.300 177.460 66.630 178.000 ;
        RECT 66.800 177.260 67.005 178.230 ;
        RECT 67.175 177.720 67.530 178.090 ;
        RECT 67.810 178.080 67.980 178.270 ;
        RECT 68.150 178.245 68.405 178.820 ;
        RECT 67.810 177.750 68.065 178.080 ;
        RECT 67.810 177.540 67.980 177.750 ;
        RECT 65.275 177.030 67.005 177.260 ;
        RECT 65.275 176.630 65.605 177.030 ;
        RECT 65.775 176.440 66.105 176.800 ;
        RECT 66.305 176.610 67.005 177.030 ;
        RECT 67.265 177.370 67.980 177.540 ;
        RECT 68.235 177.515 68.405 178.245 ;
        RECT 68.580 178.150 68.840 178.990 ;
        RECT 69.130 178.360 69.415 178.820 ;
        RECT 69.585 178.530 69.855 178.990 ;
        RECT 69.130 178.190 70.085 178.360 ;
        RECT 67.265 176.610 67.435 177.370 ;
        RECT 67.650 176.440 67.980 177.200 ;
        RECT 68.150 176.610 68.405 177.515 ;
        RECT 68.580 176.440 68.840 177.590 ;
        RECT 69.015 177.460 69.705 178.020 ;
        RECT 69.875 177.290 70.085 178.190 ;
        RECT 69.130 177.070 70.085 177.290 ;
        RECT 70.255 178.020 70.655 178.820 ;
        RECT 70.845 178.360 71.125 178.820 ;
        RECT 71.645 178.530 71.970 178.990 ;
        RECT 70.845 178.190 71.970 178.360 ;
        RECT 72.140 178.250 72.525 178.820 ;
        RECT 71.520 178.080 71.970 178.190 ;
        RECT 70.255 177.460 71.350 178.020 ;
        RECT 71.520 177.750 72.075 178.080 ;
        RECT 69.130 176.610 69.415 177.070 ;
        RECT 69.585 176.440 69.855 176.900 ;
        RECT 70.255 176.610 70.655 177.460 ;
        RECT 71.520 177.290 71.970 177.750 ;
        RECT 72.245 177.580 72.525 178.250 ;
        RECT 72.970 178.180 73.215 178.785 ;
        RECT 73.435 178.455 73.945 178.990 ;
        RECT 70.845 177.070 71.970 177.290 ;
        RECT 70.845 176.610 71.125 177.070 ;
        RECT 71.645 176.440 71.970 176.900 ;
        RECT 72.140 176.610 72.525 177.580 ;
        RECT 72.695 178.010 73.925 178.180 ;
        RECT 72.695 177.200 73.035 178.010 ;
        RECT 73.205 177.445 73.955 177.635 ;
        RECT 72.695 176.790 73.210 177.200 ;
        RECT 73.445 176.440 73.615 177.200 ;
        RECT 73.785 176.780 73.955 177.445 ;
        RECT 74.125 177.460 74.315 178.820 ;
        RECT 74.485 177.970 74.760 178.820 ;
        RECT 74.950 178.455 75.480 178.820 ;
        RECT 75.905 178.590 76.235 178.990 ;
        RECT 75.305 178.420 75.480 178.455 ;
        RECT 74.485 177.800 74.765 177.970 ;
        RECT 74.485 177.660 74.760 177.800 ;
        RECT 74.965 177.460 75.135 178.260 ;
        RECT 74.125 177.290 75.135 177.460 ;
        RECT 75.305 178.250 76.235 178.420 ;
        RECT 76.405 178.250 76.660 178.820 ;
        RECT 76.835 178.265 77.125 178.990 ;
        RECT 77.410 178.360 77.695 178.820 ;
        RECT 77.865 178.530 78.135 178.990 ;
        RECT 75.305 177.120 75.475 178.250 ;
        RECT 76.065 178.080 76.235 178.250 ;
        RECT 74.350 176.950 75.475 177.120 ;
        RECT 75.645 177.750 75.840 178.080 ;
        RECT 76.065 177.750 76.320 178.080 ;
        RECT 75.645 176.780 75.815 177.750 ;
        RECT 76.490 177.580 76.660 178.250 ;
        RECT 77.410 178.190 78.365 178.360 ;
        RECT 73.785 176.610 75.815 176.780 ;
        RECT 75.985 176.440 76.155 177.580 ;
        RECT 76.325 176.610 76.660 177.580 ;
        RECT 76.835 176.440 77.125 177.605 ;
        RECT 77.295 177.460 77.985 178.020 ;
        RECT 78.155 177.290 78.365 178.190 ;
        RECT 77.410 177.070 78.365 177.290 ;
        RECT 78.535 178.020 78.935 178.820 ;
        RECT 79.125 178.360 79.405 178.820 ;
        RECT 79.925 178.530 80.250 178.990 ;
        RECT 79.125 178.190 80.250 178.360 ;
        RECT 80.420 178.250 80.805 178.820 ;
        RECT 79.800 178.080 80.250 178.190 ;
        RECT 78.535 177.460 79.630 178.020 ;
        RECT 79.800 177.750 80.355 178.080 ;
        RECT 77.410 176.610 77.695 177.070 ;
        RECT 77.865 176.440 78.135 176.900 ;
        RECT 78.535 176.610 78.935 177.460 ;
        RECT 79.800 177.290 80.250 177.750 ;
        RECT 80.525 177.580 80.805 178.250 ;
        RECT 81.035 178.170 81.245 178.990 ;
        RECT 81.415 178.190 81.745 178.820 ;
        RECT 81.415 177.590 81.665 178.190 ;
        RECT 81.915 178.170 82.145 178.990 ;
        RECT 83.390 178.360 83.675 178.820 ;
        RECT 83.845 178.530 84.115 178.990 ;
        RECT 83.390 178.190 84.345 178.360 ;
        RECT 81.835 177.750 82.165 178.000 ;
        RECT 79.125 177.070 80.250 177.290 ;
        RECT 79.125 176.610 79.405 177.070 ;
        RECT 79.925 176.440 80.250 176.900 ;
        RECT 80.420 176.610 80.805 177.580 ;
        RECT 81.035 176.440 81.245 177.580 ;
        RECT 81.415 176.610 81.745 177.590 ;
        RECT 81.915 176.440 82.145 177.580 ;
        RECT 83.275 177.460 83.965 178.020 ;
        RECT 84.135 177.290 84.345 178.190 ;
        RECT 83.390 177.070 84.345 177.290 ;
        RECT 84.515 178.020 84.915 178.820 ;
        RECT 85.105 178.360 85.385 178.820 ;
        RECT 85.905 178.530 86.230 178.990 ;
        RECT 85.105 178.190 86.230 178.360 ;
        RECT 86.400 178.250 86.785 178.820 ;
        RECT 85.780 178.080 86.230 178.190 ;
        RECT 84.515 177.460 85.610 178.020 ;
        RECT 85.780 177.750 86.335 178.080 ;
        RECT 83.390 176.610 83.675 177.070 ;
        RECT 83.845 176.440 84.115 176.900 ;
        RECT 84.515 176.610 84.915 177.460 ;
        RECT 85.780 177.290 86.230 177.750 ;
        RECT 86.505 177.580 86.785 178.250 ;
        RECT 85.105 177.070 86.230 177.290 ;
        RECT 85.105 176.610 85.385 177.070 ;
        RECT 85.905 176.440 86.230 176.900 ;
        RECT 86.400 176.610 86.785 177.580 ;
        RECT 86.960 178.250 87.215 178.820 ;
        RECT 87.385 178.590 87.715 178.990 ;
        RECT 88.140 178.455 88.670 178.820 ;
        RECT 88.860 178.650 89.135 178.820 ;
        RECT 88.855 178.480 89.135 178.650 ;
        RECT 88.140 178.420 88.315 178.455 ;
        RECT 87.385 178.250 88.315 178.420 ;
        RECT 86.960 177.580 87.130 178.250 ;
        RECT 87.385 178.080 87.555 178.250 ;
        RECT 87.300 177.750 87.555 178.080 ;
        RECT 87.780 177.750 87.975 178.080 ;
        RECT 86.960 176.610 87.295 177.580 ;
        RECT 87.465 176.440 87.635 177.580 ;
        RECT 87.805 176.780 87.975 177.750 ;
        RECT 88.145 177.120 88.315 178.250 ;
        RECT 88.485 177.460 88.655 178.260 ;
        RECT 88.860 177.660 89.135 178.480 ;
        RECT 89.305 177.460 89.495 178.820 ;
        RECT 89.675 178.455 90.185 178.990 ;
        RECT 90.405 178.180 90.650 178.785 ;
        RECT 91.210 178.360 91.495 178.820 ;
        RECT 91.665 178.530 91.935 178.990 ;
        RECT 91.210 178.190 92.165 178.360 ;
        RECT 89.695 178.010 90.925 178.180 ;
        RECT 88.485 177.290 89.495 177.460 ;
        RECT 89.665 177.445 90.415 177.635 ;
        RECT 88.145 176.950 89.270 177.120 ;
        RECT 89.665 176.780 89.835 177.445 ;
        RECT 90.585 177.200 90.925 178.010 ;
        RECT 91.095 177.460 91.785 178.020 ;
        RECT 91.955 177.290 92.165 178.190 ;
        RECT 87.805 176.610 89.835 176.780 ;
        RECT 90.005 176.440 90.175 177.200 ;
        RECT 90.410 176.790 90.925 177.200 ;
        RECT 91.210 177.070 92.165 177.290 ;
        RECT 92.335 178.020 92.735 178.820 ;
        RECT 92.925 178.360 93.205 178.820 ;
        RECT 93.725 178.530 94.050 178.990 ;
        RECT 92.925 178.190 94.050 178.360 ;
        RECT 94.220 178.250 94.605 178.820 ;
        RECT 93.600 178.080 94.050 178.190 ;
        RECT 92.335 177.460 93.430 178.020 ;
        RECT 93.600 177.750 94.155 178.080 ;
        RECT 91.210 176.610 91.495 177.070 ;
        RECT 91.665 176.440 91.935 176.900 ;
        RECT 92.335 176.610 92.735 177.460 ;
        RECT 93.600 177.290 94.050 177.750 ;
        RECT 94.325 177.580 94.605 178.250 ;
        RECT 92.925 177.070 94.050 177.290 ;
        RECT 92.925 176.610 93.205 177.070 ;
        RECT 93.725 176.440 94.050 176.900 ;
        RECT 94.220 176.610 94.605 177.580 ;
        RECT 94.775 178.190 95.115 178.820 ;
        RECT 95.285 178.190 95.535 178.990 ;
        RECT 95.725 178.340 96.055 178.820 ;
        RECT 96.225 178.530 96.450 178.990 ;
        RECT 96.620 178.340 96.950 178.820 ;
        RECT 94.775 177.580 94.950 178.190 ;
        RECT 95.725 178.170 96.950 178.340 ;
        RECT 97.580 178.210 98.080 178.820 ;
        RECT 95.120 177.830 95.815 178.000 ;
        RECT 95.645 177.580 95.815 177.830 ;
        RECT 95.990 177.800 96.410 178.000 ;
        RECT 96.580 177.800 96.910 178.000 ;
        RECT 97.080 177.800 97.410 178.000 ;
        RECT 97.580 177.580 97.750 178.210 ;
        RECT 98.455 178.190 98.795 178.820 ;
        RECT 98.965 178.190 99.215 178.990 ;
        RECT 99.405 178.340 99.735 178.820 ;
        RECT 99.905 178.530 100.130 178.990 ;
        RECT 100.300 178.340 100.630 178.820 ;
        RECT 97.935 177.750 98.285 178.000 ;
        RECT 98.455 177.580 98.630 178.190 ;
        RECT 99.405 178.170 100.630 178.340 ;
        RECT 101.260 178.210 101.760 178.820 ;
        RECT 102.595 178.265 102.885 178.990 ;
        RECT 98.800 177.830 99.495 178.000 ;
        RECT 99.325 177.580 99.495 177.830 ;
        RECT 99.670 177.800 100.090 178.000 ;
        RECT 100.260 177.800 100.590 178.000 ;
        RECT 100.760 177.800 101.090 178.000 ;
        RECT 101.260 177.580 101.430 178.210 ;
        RECT 104.250 178.180 104.495 178.785 ;
        RECT 104.715 178.455 105.225 178.990 ;
        RECT 103.975 178.010 105.205 178.180 ;
        RECT 101.615 177.750 101.965 178.000 ;
        RECT 94.775 176.610 95.115 177.580 ;
        RECT 95.285 176.440 95.455 177.580 ;
        RECT 95.645 177.410 98.080 177.580 ;
        RECT 95.725 176.440 95.975 177.240 ;
        RECT 96.620 176.610 96.950 177.410 ;
        RECT 97.250 176.440 97.580 177.240 ;
        RECT 97.750 176.610 98.080 177.410 ;
        RECT 98.455 176.610 98.795 177.580 ;
        RECT 98.965 176.440 99.135 177.580 ;
        RECT 99.325 177.410 101.760 177.580 ;
        RECT 99.405 176.440 99.655 177.240 ;
        RECT 100.300 176.610 100.630 177.410 ;
        RECT 100.930 176.440 101.260 177.240 ;
        RECT 101.430 176.610 101.760 177.410 ;
        RECT 102.595 176.440 102.885 177.605 ;
        RECT 103.975 177.200 104.315 178.010 ;
        RECT 104.485 177.445 105.235 177.635 ;
        RECT 103.975 176.790 104.490 177.200 ;
        RECT 104.725 176.440 104.895 177.200 ;
        RECT 105.065 176.780 105.235 177.445 ;
        RECT 105.405 177.460 105.595 178.820 ;
        RECT 105.765 178.650 106.040 178.820 ;
        RECT 105.765 178.480 106.045 178.650 ;
        RECT 105.765 177.660 106.040 178.480 ;
        RECT 106.230 178.455 106.760 178.820 ;
        RECT 107.185 178.590 107.515 178.990 ;
        RECT 106.585 178.420 106.760 178.455 ;
        RECT 106.245 177.460 106.415 178.260 ;
        RECT 105.405 177.290 106.415 177.460 ;
        RECT 106.585 178.250 107.515 178.420 ;
        RECT 107.685 178.250 107.940 178.820 ;
        RECT 106.585 177.120 106.755 178.250 ;
        RECT 107.345 178.080 107.515 178.250 ;
        RECT 105.630 176.950 106.755 177.120 ;
        RECT 106.925 177.750 107.120 178.080 ;
        RECT 107.345 177.750 107.600 178.080 ;
        RECT 106.925 176.780 107.095 177.750 ;
        RECT 107.770 177.580 107.940 178.250 ;
        RECT 108.230 178.360 108.515 178.820 ;
        RECT 108.685 178.530 108.955 178.990 ;
        RECT 108.230 178.190 109.185 178.360 ;
        RECT 105.065 176.610 107.095 176.780 ;
        RECT 107.265 176.440 107.435 177.580 ;
        RECT 107.605 176.610 107.940 177.580 ;
        RECT 108.115 177.460 108.805 178.020 ;
        RECT 108.975 177.290 109.185 178.190 ;
        RECT 108.230 177.070 109.185 177.290 ;
        RECT 109.355 178.020 109.755 178.820 ;
        RECT 109.945 178.360 110.225 178.820 ;
        RECT 110.745 178.530 111.070 178.990 ;
        RECT 109.945 178.190 111.070 178.360 ;
        RECT 111.240 178.250 111.625 178.820 ;
        RECT 110.620 178.080 111.070 178.190 ;
        RECT 109.355 177.460 110.450 178.020 ;
        RECT 110.620 177.750 111.175 178.080 ;
        RECT 108.230 176.610 108.515 177.070 ;
        RECT 108.685 176.440 108.955 176.900 ;
        RECT 109.355 176.610 109.755 177.460 ;
        RECT 110.620 177.290 111.070 177.750 ;
        RECT 111.345 177.580 111.625 178.250 ;
        RECT 111.795 178.220 114.385 178.990 ;
        RECT 114.555 178.240 115.765 178.990 ;
        RECT 109.945 177.070 111.070 177.290 ;
        RECT 109.945 176.610 110.225 177.070 ;
        RECT 110.745 176.440 111.070 176.900 ;
        RECT 111.240 176.610 111.625 177.580 ;
        RECT 111.795 177.530 113.005 178.050 ;
        RECT 113.175 177.700 114.385 178.220 ;
        RECT 114.555 177.530 115.075 178.070 ;
        RECT 115.245 177.700 115.765 178.240 ;
        RECT 111.795 176.440 114.385 177.530 ;
        RECT 114.555 176.440 115.765 177.530 ;
        RECT 10.510 176.270 115.850 176.440 ;
        RECT 10.595 175.180 11.805 176.270 ;
        RECT 10.595 174.470 11.115 175.010 ;
        RECT 11.285 174.640 11.805 175.180 ;
        RECT 12.435 175.105 12.725 176.270 ;
        RECT 13.355 175.180 15.025 176.270 ;
        RECT 13.355 174.660 14.105 175.180 ;
        RECT 15.200 175.080 15.455 175.960 ;
        RECT 15.625 175.130 15.930 176.270 ;
        RECT 16.270 175.890 16.600 176.270 ;
        RECT 16.780 175.720 16.950 176.010 ;
        RECT 17.120 175.810 17.370 176.270 ;
        RECT 16.150 175.550 16.950 175.720 ;
        RECT 17.540 175.760 18.410 176.100 ;
        RECT 14.275 174.490 15.025 175.010 ;
        RECT 10.595 173.720 11.805 174.470 ;
        RECT 12.435 173.720 12.725 174.445 ;
        RECT 13.355 173.720 15.025 174.490 ;
        RECT 15.200 174.430 15.410 175.080 ;
        RECT 16.150 174.960 16.320 175.550 ;
        RECT 17.540 175.380 17.710 175.760 ;
        RECT 18.645 175.640 18.815 176.100 ;
        RECT 18.985 175.810 19.355 176.270 ;
        RECT 19.650 175.670 19.820 176.010 ;
        RECT 19.990 175.840 20.320 176.270 ;
        RECT 20.555 175.670 20.725 176.010 ;
        RECT 16.490 175.210 17.710 175.380 ;
        RECT 17.880 175.300 18.340 175.590 ;
        RECT 18.645 175.470 19.205 175.640 ;
        RECT 19.650 175.500 20.725 175.670 ;
        RECT 20.895 175.770 21.575 176.100 ;
        RECT 21.790 175.770 22.040 176.100 ;
        RECT 22.210 175.810 22.460 176.270 ;
        RECT 19.035 175.330 19.205 175.470 ;
        RECT 17.880 175.290 18.845 175.300 ;
        RECT 17.540 175.120 17.710 175.210 ;
        RECT 18.170 175.130 18.845 175.290 ;
        RECT 15.580 174.930 16.320 174.960 ;
        RECT 15.580 174.630 16.495 174.930 ;
        RECT 16.170 174.455 16.495 174.630 ;
        RECT 15.200 173.900 15.455 174.430 ;
        RECT 15.625 173.720 15.930 174.180 ;
        RECT 16.175 174.100 16.495 174.455 ;
        RECT 16.665 174.670 17.205 175.040 ;
        RECT 17.540 174.950 17.945 175.120 ;
        RECT 16.665 174.270 16.905 174.670 ;
        RECT 17.385 174.500 17.605 174.780 ;
        RECT 17.075 174.330 17.605 174.500 ;
        RECT 17.075 174.100 17.245 174.330 ;
        RECT 17.775 174.170 17.945 174.950 ;
        RECT 18.115 174.340 18.465 174.960 ;
        RECT 18.635 174.340 18.845 175.130 ;
        RECT 19.035 175.160 20.535 175.330 ;
        RECT 19.035 174.470 19.205 175.160 ;
        RECT 20.895 174.990 21.065 175.770 ;
        RECT 21.870 175.640 22.040 175.770 ;
        RECT 19.375 174.820 21.065 174.990 ;
        RECT 21.235 175.210 21.700 175.600 ;
        RECT 21.870 175.470 22.265 175.640 ;
        RECT 19.375 174.640 19.545 174.820 ;
        RECT 16.175 173.930 17.245 174.100 ;
        RECT 17.415 173.720 17.605 174.160 ;
        RECT 17.775 173.890 18.725 174.170 ;
        RECT 19.035 174.080 19.295 174.470 ;
        RECT 19.715 174.400 20.505 174.650 ;
        RECT 18.945 173.910 19.295 174.080 ;
        RECT 19.505 173.720 19.835 174.180 ;
        RECT 20.710 174.110 20.880 174.820 ;
        RECT 21.235 174.620 21.405 175.210 ;
        RECT 21.050 174.400 21.405 174.620 ;
        RECT 21.575 174.400 21.925 175.020 ;
        RECT 22.095 174.110 22.265 175.470 ;
        RECT 22.630 175.300 22.955 176.085 ;
        RECT 22.435 174.250 22.895 175.300 ;
        RECT 20.710 173.940 21.565 174.110 ;
        RECT 21.770 173.940 22.265 174.110 ;
        RECT 22.435 173.720 22.765 174.080 ;
        RECT 23.125 173.980 23.295 176.100 ;
        RECT 23.465 175.770 23.795 176.270 ;
        RECT 23.965 175.600 24.220 176.100 ;
        RECT 23.470 175.430 24.220 175.600 ;
        RECT 23.470 174.440 23.700 175.430 ;
        RECT 23.870 174.610 24.220 175.260 ;
        RECT 24.400 175.080 24.655 175.960 ;
        RECT 24.825 175.130 25.130 176.270 ;
        RECT 25.470 175.890 25.800 176.270 ;
        RECT 25.980 175.720 26.150 176.010 ;
        RECT 26.320 175.810 26.570 176.270 ;
        RECT 25.350 175.550 26.150 175.720 ;
        RECT 26.740 175.760 27.610 176.100 ;
        RECT 23.470 174.270 24.220 174.440 ;
        RECT 23.465 173.720 23.795 174.100 ;
        RECT 23.965 173.980 24.220 174.270 ;
        RECT 24.400 174.430 24.610 175.080 ;
        RECT 25.350 174.960 25.520 175.550 ;
        RECT 26.740 175.380 26.910 175.760 ;
        RECT 27.845 175.640 28.015 176.100 ;
        RECT 28.185 175.810 28.555 176.270 ;
        RECT 28.850 175.670 29.020 176.010 ;
        RECT 29.190 175.840 29.520 176.270 ;
        RECT 29.755 175.670 29.925 176.010 ;
        RECT 25.690 175.210 26.910 175.380 ;
        RECT 27.080 175.300 27.540 175.590 ;
        RECT 27.845 175.470 28.405 175.640 ;
        RECT 28.850 175.500 29.925 175.670 ;
        RECT 30.095 175.770 30.775 176.100 ;
        RECT 30.990 175.770 31.240 176.100 ;
        RECT 31.410 175.810 31.660 176.270 ;
        RECT 28.235 175.330 28.405 175.470 ;
        RECT 27.080 175.290 28.045 175.300 ;
        RECT 26.740 175.120 26.910 175.210 ;
        RECT 27.370 175.130 28.045 175.290 ;
        RECT 24.780 174.930 25.520 174.960 ;
        RECT 24.780 174.630 25.695 174.930 ;
        RECT 25.370 174.455 25.695 174.630 ;
        RECT 24.400 173.900 24.655 174.430 ;
        RECT 24.825 173.720 25.130 174.180 ;
        RECT 25.375 174.100 25.695 174.455 ;
        RECT 25.865 174.670 26.405 175.040 ;
        RECT 26.740 174.950 27.145 175.120 ;
        RECT 25.865 174.270 26.105 174.670 ;
        RECT 26.585 174.500 26.805 174.780 ;
        RECT 26.275 174.330 26.805 174.500 ;
        RECT 26.275 174.100 26.445 174.330 ;
        RECT 26.975 174.170 27.145 174.950 ;
        RECT 27.315 174.340 27.665 174.960 ;
        RECT 27.835 174.340 28.045 175.130 ;
        RECT 28.235 175.160 29.735 175.330 ;
        RECT 28.235 174.470 28.405 175.160 ;
        RECT 30.095 174.990 30.265 175.770 ;
        RECT 31.070 175.640 31.240 175.770 ;
        RECT 28.575 174.820 30.265 174.990 ;
        RECT 30.435 175.210 30.900 175.600 ;
        RECT 31.070 175.470 31.465 175.640 ;
        RECT 28.575 174.640 28.745 174.820 ;
        RECT 25.375 173.930 26.445 174.100 ;
        RECT 26.615 173.720 26.805 174.160 ;
        RECT 26.975 173.890 27.925 174.170 ;
        RECT 28.235 174.080 28.495 174.470 ;
        RECT 28.915 174.400 29.705 174.650 ;
        RECT 28.145 173.910 28.495 174.080 ;
        RECT 28.705 173.720 29.035 174.180 ;
        RECT 29.910 174.110 30.080 174.820 ;
        RECT 30.435 174.620 30.605 175.210 ;
        RECT 30.250 174.400 30.605 174.620 ;
        RECT 30.775 174.400 31.125 175.020 ;
        RECT 31.295 174.110 31.465 175.470 ;
        RECT 31.830 175.300 32.155 176.085 ;
        RECT 31.635 174.250 32.095 175.300 ;
        RECT 29.910 173.940 30.765 174.110 ;
        RECT 30.970 173.940 31.465 174.110 ;
        RECT 31.635 173.720 31.965 174.080 ;
        RECT 32.325 173.980 32.495 176.100 ;
        RECT 32.665 175.770 32.995 176.270 ;
        RECT 33.165 175.600 33.420 176.100 ;
        RECT 32.670 175.430 33.420 175.600 ;
        RECT 32.670 174.440 32.900 175.430 ;
        RECT 34.720 175.300 35.050 176.100 ;
        RECT 35.220 175.470 35.550 176.270 ;
        RECT 35.850 175.300 36.180 176.100 ;
        RECT 36.825 175.470 37.075 176.270 ;
        RECT 33.070 174.610 33.420 175.260 ;
        RECT 34.720 175.130 37.155 175.300 ;
        RECT 37.345 175.130 37.515 176.270 ;
        RECT 37.685 175.130 38.025 176.100 ;
        RECT 34.515 174.710 34.865 174.960 ;
        RECT 35.050 174.500 35.220 175.130 ;
        RECT 35.390 174.710 35.720 174.910 ;
        RECT 35.890 174.710 36.220 174.910 ;
        RECT 36.390 174.710 36.810 174.910 ;
        RECT 36.985 174.880 37.155 175.130 ;
        RECT 36.985 174.710 37.680 174.880 ;
        RECT 32.670 174.270 33.420 174.440 ;
        RECT 32.665 173.720 32.995 174.100 ;
        RECT 33.165 173.980 33.420 174.270 ;
        RECT 34.720 173.890 35.220 174.500 ;
        RECT 35.850 174.370 37.075 174.540 ;
        RECT 37.850 174.520 38.025 175.130 ;
        RECT 38.195 175.105 38.485 176.270 ;
        RECT 39.320 175.300 39.650 176.100 ;
        RECT 39.820 175.470 40.150 176.270 ;
        RECT 40.450 175.300 40.780 176.100 ;
        RECT 41.425 175.470 41.675 176.270 ;
        RECT 39.320 175.130 41.755 175.300 ;
        RECT 41.945 175.130 42.115 176.270 ;
        RECT 42.285 175.130 42.625 176.100 ;
        RECT 39.115 174.710 39.465 174.960 ;
        RECT 35.850 173.890 36.180 174.370 ;
        RECT 36.350 173.720 36.575 174.180 ;
        RECT 36.745 173.890 37.075 174.370 ;
        RECT 37.265 173.720 37.515 174.520 ;
        RECT 37.685 173.890 38.025 174.520 ;
        RECT 39.650 174.500 39.820 175.130 ;
        RECT 39.990 174.710 40.320 174.910 ;
        RECT 40.490 174.710 40.820 174.910 ;
        RECT 40.990 174.710 41.410 174.910 ;
        RECT 41.585 174.880 41.755 175.130 ;
        RECT 41.585 174.710 42.280 174.880 ;
        RECT 38.195 173.720 38.485 174.445 ;
        RECT 39.320 173.890 39.820 174.500 ;
        RECT 40.450 174.370 41.675 174.540 ;
        RECT 42.450 174.520 42.625 175.130 ;
        RECT 40.450 173.890 40.780 174.370 ;
        RECT 40.950 173.720 41.175 174.180 ;
        RECT 41.345 173.890 41.675 174.370 ;
        RECT 41.865 173.720 42.115 174.520 ;
        RECT 42.285 173.890 42.625 174.520 ;
        RECT 42.795 175.130 43.135 176.100 ;
        RECT 43.305 175.130 43.475 176.270 ;
        RECT 43.745 175.470 43.995 176.270 ;
        RECT 44.640 175.300 44.970 176.100 ;
        RECT 45.270 175.470 45.600 176.270 ;
        RECT 45.770 175.300 46.100 176.100 ;
        RECT 46.590 175.640 46.875 176.100 ;
        RECT 47.045 175.810 47.315 176.270 ;
        RECT 46.590 175.420 47.545 175.640 ;
        RECT 43.665 175.130 46.100 175.300 ;
        RECT 42.795 174.520 42.970 175.130 ;
        RECT 43.665 174.880 43.835 175.130 ;
        RECT 43.140 174.710 43.835 174.880 ;
        RECT 44.010 174.710 44.430 174.910 ;
        RECT 44.600 174.710 44.930 174.910 ;
        RECT 45.100 174.710 45.430 174.910 ;
        RECT 42.795 173.890 43.135 174.520 ;
        RECT 43.305 173.720 43.555 174.520 ;
        RECT 43.745 174.370 44.970 174.540 ;
        RECT 43.745 173.890 44.075 174.370 ;
        RECT 44.245 173.720 44.470 174.180 ;
        RECT 44.640 173.890 44.970 174.370 ;
        RECT 45.600 174.500 45.770 175.130 ;
        RECT 45.955 174.710 46.305 174.960 ;
        RECT 46.475 174.690 47.165 175.250 ;
        RECT 47.335 174.520 47.545 175.420 ;
        RECT 45.600 173.890 46.100 174.500 ;
        RECT 46.590 174.350 47.545 174.520 ;
        RECT 47.715 175.250 48.115 176.100 ;
        RECT 48.305 175.640 48.585 176.100 ;
        RECT 49.105 175.810 49.430 176.270 ;
        RECT 48.305 175.420 49.430 175.640 ;
        RECT 47.715 174.690 48.810 175.250 ;
        RECT 48.980 174.960 49.430 175.420 ;
        RECT 49.600 175.130 49.985 176.100 ;
        RECT 46.590 173.890 46.875 174.350 ;
        RECT 47.045 173.720 47.315 174.180 ;
        RECT 47.715 173.890 48.115 174.690 ;
        RECT 48.980 174.630 49.535 174.960 ;
        RECT 48.980 174.520 49.430 174.630 ;
        RECT 48.305 174.350 49.430 174.520 ;
        RECT 49.705 174.460 49.985 175.130 ;
        RECT 51.075 175.510 51.590 175.920 ;
        RECT 51.825 175.510 51.995 176.270 ;
        RECT 52.165 175.930 54.195 176.100 ;
        RECT 51.075 174.700 51.415 175.510 ;
        RECT 52.165 175.265 52.335 175.930 ;
        RECT 52.730 175.590 53.855 175.760 ;
        RECT 51.585 175.075 52.335 175.265 ;
        RECT 52.505 175.250 53.515 175.420 ;
        RECT 51.075 174.530 52.305 174.700 ;
        RECT 48.305 173.890 48.585 174.350 ;
        RECT 49.105 173.720 49.430 174.180 ;
        RECT 49.600 173.890 49.985 174.460 ;
        RECT 51.350 173.925 51.595 174.530 ;
        RECT 51.815 173.720 52.325 174.255 ;
        RECT 52.505 173.890 52.695 175.250 ;
        RECT 52.865 174.570 53.140 175.050 ;
        RECT 52.865 174.400 53.145 174.570 ;
        RECT 53.345 174.450 53.515 175.250 ;
        RECT 53.685 174.460 53.855 175.590 ;
        RECT 54.025 174.960 54.195 175.930 ;
        RECT 54.365 175.130 54.535 176.270 ;
        RECT 54.705 175.130 55.040 176.100 ;
        RECT 55.275 175.130 55.485 176.270 ;
        RECT 54.025 174.630 54.220 174.960 ;
        RECT 54.445 174.630 54.700 174.960 ;
        RECT 54.445 174.460 54.615 174.630 ;
        RECT 54.870 174.460 55.040 175.130 ;
        RECT 55.655 175.120 55.985 176.100 ;
        RECT 56.155 175.130 56.385 176.270 ;
        RECT 56.685 175.340 56.855 176.100 ;
        RECT 57.035 175.510 57.365 176.270 ;
        RECT 56.685 175.170 57.350 175.340 ;
        RECT 57.535 175.195 57.805 176.100 ;
        RECT 52.865 173.890 53.140 174.400 ;
        RECT 53.685 174.290 54.615 174.460 ;
        RECT 53.685 174.255 53.860 174.290 ;
        RECT 53.330 173.890 53.860 174.255 ;
        RECT 54.285 173.720 54.615 174.120 ;
        RECT 54.785 173.890 55.040 174.460 ;
        RECT 55.275 173.720 55.485 174.540 ;
        RECT 55.655 174.520 55.905 175.120 ;
        RECT 57.180 175.025 57.350 175.170 ;
        RECT 56.075 174.710 56.405 174.960 ;
        RECT 56.615 174.620 56.945 174.990 ;
        RECT 57.180 174.695 57.465 175.025 ;
        RECT 55.655 173.890 55.985 174.520 ;
        RECT 56.155 173.720 56.385 174.540 ;
        RECT 57.180 174.440 57.350 174.695 ;
        RECT 56.685 174.270 57.350 174.440 ;
        RECT 57.635 174.395 57.805 175.195 ;
        RECT 58.435 175.180 60.105 176.270 ;
        RECT 58.435 174.660 59.185 175.180 ;
        RECT 60.280 175.120 60.540 176.270 ;
        RECT 60.715 175.195 60.970 176.100 ;
        RECT 61.140 175.510 61.470 176.270 ;
        RECT 61.685 175.340 61.855 176.100 ;
        RECT 59.355 174.490 60.105 175.010 ;
        RECT 56.685 173.890 56.855 174.270 ;
        RECT 57.035 173.720 57.365 174.100 ;
        RECT 57.545 173.890 57.805 174.395 ;
        RECT 58.435 173.720 60.105 174.490 ;
        RECT 60.280 173.720 60.540 174.560 ;
        RECT 60.715 174.465 60.885 175.195 ;
        RECT 61.140 175.170 61.855 175.340 ;
        RECT 61.140 174.960 61.310 175.170 ;
        RECT 62.120 175.120 62.380 176.270 ;
        RECT 62.555 175.195 62.810 176.100 ;
        RECT 62.980 175.510 63.310 176.270 ;
        RECT 63.525 175.340 63.695 176.100 ;
        RECT 61.055 174.630 61.310 174.960 ;
        RECT 60.715 173.890 60.970 174.465 ;
        RECT 61.140 174.440 61.310 174.630 ;
        RECT 61.590 174.620 61.945 174.990 ;
        RECT 61.140 174.270 61.855 174.440 ;
        RECT 61.140 173.720 61.470 174.100 ;
        RECT 61.685 173.890 61.855 174.270 ;
        RECT 62.120 173.720 62.380 174.560 ;
        RECT 62.555 174.465 62.725 175.195 ;
        RECT 62.980 175.170 63.695 175.340 ;
        RECT 62.980 174.960 63.150 175.170 ;
        RECT 63.955 175.105 64.245 176.270 ;
        RECT 64.415 175.180 66.085 176.270 ;
        RECT 62.895 174.630 63.150 174.960 ;
        RECT 62.555 173.890 62.810 174.465 ;
        RECT 62.980 174.440 63.150 174.630 ;
        RECT 63.430 174.620 63.785 174.990 ;
        RECT 64.415 174.660 65.165 175.180 ;
        RECT 66.255 175.130 66.595 176.100 ;
        RECT 66.765 175.130 66.935 176.270 ;
        RECT 67.205 175.470 67.455 176.270 ;
        RECT 68.100 175.300 68.430 176.100 ;
        RECT 68.730 175.470 69.060 176.270 ;
        RECT 69.230 175.300 69.560 176.100 ;
        RECT 67.125 175.130 69.560 175.300 ;
        RECT 69.935 175.130 70.275 176.100 ;
        RECT 70.445 175.130 70.615 176.270 ;
        RECT 70.885 175.470 71.135 176.270 ;
        RECT 71.780 175.300 72.110 176.100 ;
        RECT 72.410 175.470 72.740 176.270 ;
        RECT 72.910 175.300 73.240 176.100 ;
        RECT 70.805 175.130 73.240 175.300 ;
        RECT 73.615 175.130 73.955 176.100 ;
        RECT 74.125 175.130 74.295 176.270 ;
        RECT 74.565 175.470 74.815 176.270 ;
        RECT 75.460 175.300 75.790 176.100 ;
        RECT 76.090 175.470 76.420 176.270 ;
        RECT 76.590 175.300 76.920 176.100 ;
        RECT 78.225 175.460 78.520 176.270 ;
        RECT 74.485 175.130 76.920 175.300 ;
        RECT 65.335 174.490 66.085 175.010 ;
        RECT 62.980 174.270 63.695 174.440 ;
        RECT 62.980 173.720 63.310 174.100 ;
        RECT 63.525 173.890 63.695 174.270 ;
        RECT 63.955 173.720 64.245 174.445 ;
        RECT 64.415 173.720 66.085 174.490 ;
        RECT 66.255 174.520 66.430 175.130 ;
        RECT 67.125 174.880 67.295 175.130 ;
        RECT 66.600 174.710 67.295 174.880 ;
        RECT 67.470 174.710 67.890 174.910 ;
        RECT 68.060 174.710 68.390 174.910 ;
        RECT 68.560 174.710 68.890 174.910 ;
        RECT 66.255 173.890 66.595 174.520 ;
        RECT 66.765 173.720 67.015 174.520 ;
        RECT 67.205 174.370 68.430 174.540 ;
        RECT 67.205 173.890 67.535 174.370 ;
        RECT 67.705 173.720 67.930 174.180 ;
        RECT 68.100 173.890 68.430 174.370 ;
        RECT 69.060 174.500 69.230 175.130 ;
        RECT 69.415 174.710 69.765 174.960 ;
        RECT 69.935 174.520 70.110 175.130 ;
        RECT 70.805 174.880 70.975 175.130 ;
        RECT 70.280 174.710 70.975 174.880 ;
        RECT 71.150 174.710 71.570 174.910 ;
        RECT 71.740 174.710 72.070 174.910 ;
        RECT 72.240 174.710 72.570 174.910 ;
        RECT 69.060 173.890 69.560 174.500 ;
        RECT 69.935 173.890 70.275 174.520 ;
        RECT 70.445 173.720 70.695 174.520 ;
        RECT 70.885 174.370 72.110 174.540 ;
        RECT 70.885 173.890 71.215 174.370 ;
        RECT 71.385 173.720 71.610 174.180 ;
        RECT 71.780 173.890 72.110 174.370 ;
        RECT 72.740 174.500 72.910 175.130 ;
        RECT 73.095 174.710 73.445 174.960 ;
        RECT 73.615 174.520 73.790 175.130 ;
        RECT 74.485 174.880 74.655 175.130 ;
        RECT 73.960 174.710 74.655 174.880 ;
        RECT 74.830 174.710 75.250 174.910 ;
        RECT 75.420 174.710 75.750 174.910 ;
        RECT 75.920 174.710 76.250 174.910 ;
        RECT 72.740 173.890 73.240 174.500 ;
        RECT 73.615 173.890 73.955 174.520 ;
        RECT 74.125 173.720 74.375 174.520 ;
        RECT 74.565 174.370 75.790 174.540 ;
        RECT 74.565 173.890 74.895 174.370 ;
        RECT 75.065 173.720 75.290 174.180 ;
        RECT 75.460 173.890 75.790 174.370 ;
        RECT 76.420 174.500 76.590 175.130 ;
        RECT 78.700 174.960 78.945 176.100 ;
        RECT 79.120 175.460 79.380 176.270 ;
        RECT 79.980 176.265 86.255 176.270 ;
        RECT 79.560 174.960 79.810 176.095 ;
        RECT 79.980 175.470 80.240 176.265 ;
        RECT 80.410 175.370 80.670 176.095 ;
        RECT 80.840 175.540 81.100 176.265 ;
        RECT 81.270 175.370 81.530 176.095 ;
        RECT 81.700 175.540 81.960 176.265 ;
        RECT 82.130 175.370 82.390 176.095 ;
        RECT 82.560 175.540 82.820 176.265 ;
        RECT 82.990 175.370 83.250 176.095 ;
        RECT 83.420 175.540 83.665 176.265 ;
        RECT 83.835 175.370 84.095 176.095 ;
        RECT 84.280 175.540 84.525 176.265 ;
        RECT 84.695 175.370 84.955 176.095 ;
        RECT 85.140 175.540 85.385 176.265 ;
        RECT 85.555 175.370 85.815 176.095 ;
        RECT 86.000 175.540 86.255 176.265 ;
        RECT 80.410 175.355 85.815 175.370 ;
        RECT 86.425 175.355 86.715 176.095 ;
        RECT 86.885 175.525 87.155 176.270 ;
        RECT 80.410 175.130 87.155 175.355 ;
        RECT 88.425 175.340 88.595 176.100 ;
        RECT 88.775 175.510 89.105 176.270 ;
        RECT 88.425 175.170 89.090 175.340 ;
        RECT 89.275 175.195 89.545 176.100 ;
        RECT 76.775 174.710 77.125 174.960 ;
        RECT 76.420 173.890 76.920 174.500 ;
        RECT 78.215 174.400 78.530 174.960 ;
        RECT 78.700 174.710 85.820 174.960 ;
        RECT 78.215 173.720 78.520 174.230 ;
        RECT 78.700 173.900 78.950 174.710 ;
        RECT 79.120 173.720 79.380 174.245 ;
        RECT 79.560 173.900 79.810 174.710 ;
        RECT 85.990 174.540 87.155 175.130 ;
        RECT 88.920 175.025 89.090 175.170 ;
        RECT 88.355 174.620 88.685 174.990 ;
        RECT 88.920 174.695 89.205 175.025 ;
        RECT 80.410 174.370 87.155 174.540 ;
        RECT 88.920 174.440 89.090 174.695 ;
        RECT 79.980 173.720 80.240 174.280 ;
        RECT 80.410 173.915 80.670 174.370 ;
        RECT 80.840 173.720 81.100 174.200 ;
        RECT 81.270 173.915 81.530 174.370 ;
        RECT 81.700 173.720 81.960 174.200 ;
        RECT 82.130 173.915 82.390 174.370 ;
        RECT 82.560 173.720 82.805 174.200 ;
        RECT 82.975 173.915 83.250 174.370 ;
        RECT 83.420 173.720 83.665 174.200 ;
        RECT 83.835 173.915 84.095 174.370 ;
        RECT 84.275 173.720 84.525 174.200 ;
        RECT 84.695 173.915 84.955 174.370 ;
        RECT 85.135 173.720 85.385 174.200 ;
        RECT 85.555 173.915 85.815 174.370 ;
        RECT 85.995 173.720 86.255 174.200 ;
        RECT 86.425 173.915 86.685 174.370 ;
        RECT 88.425 174.270 89.090 174.440 ;
        RECT 89.375 174.395 89.545 175.195 ;
        RECT 89.715 175.105 90.005 176.270 ;
        RECT 90.175 175.130 90.515 176.100 ;
        RECT 90.685 175.130 90.855 176.270 ;
        RECT 91.125 175.470 91.375 176.270 ;
        RECT 92.020 175.300 92.350 176.100 ;
        RECT 92.650 175.470 92.980 176.270 ;
        RECT 93.150 175.300 93.480 176.100 ;
        RECT 91.045 175.130 93.480 175.300 ;
        RECT 94.980 175.300 95.310 176.100 ;
        RECT 95.480 175.470 95.810 176.270 ;
        RECT 96.110 175.300 96.440 176.100 ;
        RECT 97.085 175.470 97.335 176.270 ;
        RECT 94.980 175.130 97.415 175.300 ;
        RECT 97.605 175.130 97.775 176.270 ;
        RECT 97.945 175.130 98.285 176.100 ;
        RECT 90.175 174.520 90.350 175.130 ;
        RECT 91.045 174.880 91.215 175.130 ;
        RECT 90.520 174.710 91.215 174.880 ;
        RECT 91.390 174.710 91.810 174.910 ;
        RECT 91.980 174.710 92.310 174.910 ;
        RECT 92.480 174.710 92.810 174.910 ;
        RECT 86.855 173.720 87.155 174.200 ;
        RECT 88.425 173.890 88.595 174.270 ;
        RECT 88.775 173.720 89.105 174.100 ;
        RECT 89.285 173.890 89.545 174.395 ;
        RECT 89.715 173.720 90.005 174.445 ;
        RECT 90.175 173.890 90.515 174.520 ;
        RECT 90.685 173.720 90.935 174.520 ;
        RECT 91.125 174.370 92.350 174.540 ;
        RECT 91.125 173.890 91.455 174.370 ;
        RECT 91.625 173.720 91.850 174.180 ;
        RECT 92.020 173.890 92.350 174.370 ;
        RECT 92.980 174.500 93.150 175.130 ;
        RECT 93.335 174.710 93.685 174.960 ;
        RECT 94.775 174.710 95.125 174.960 ;
        RECT 95.310 174.500 95.480 175.130 ;
        RECT 95.650 174.710 95.980 174.910 ;
        RECT 96.150 174.710 96.480 174.910 ;
        RECT 96.650 174.710 97.070 174.910 ;
        RECT 97.245 174.880 97.415 175.130 ;
        RECT 97.245 174.710 97.940 174.880 ;
        RECT 98.110 174.570 98.285 175.130 ;
        RECT 98.455 175.180 101.045 176.270 ;
        RECT 101.330 175.640 101.615 176.100 ;
        RECT 101.785 175.810 102.055 176.270 ;
        RECT 101.330 175.420 102.285 175.640 ;
        RECT 98.455 174.660 99.665 175.180 ;
        RECT 92.980 173.890 93.480 174.500 ;
        RECT 94.980 173.890 95.480 174.500 ;
        RECT 96.110 174.370 97.335 174.540 ;
        RECT 98.055 174.520 98.285 174.570 ;
        RECT 96.110 173.890 96.440 174.370 ;
        RECT 96.610 173.720 96.835 174.180 ;
        RECT 97.005 173.890 97.335 174.370 ;
        RECT 97.525 173.720 97.775 174.520 ;
        RECT 97.945 173.890 98.285 174.520 ;
        RECT 99.835 174.490 101.045 175.010 ;
        RECT 101.215 174.690 101.905 175.250 ;
        RECT 102.075 174.520 102.285 175.420 ;
        RECT 98.455 173.720 101.045 174.490 ;
        RECT 101.330 174.350 102.285 174.520 ;
        RECT 102.455 175.250 102.855 176.100 ;
        RECT 103.045 175.640 103.325 176.100 ;
        RECT 103.845 175.810 104.170 176.270 ;
        RECT 103.045 175.420 104.170 175.640 ;
        RECT 102.455 174.690 103.550 175.250 ;
        RECT 103.720 174.960 104.170 175.420 ;
        RECT 104.340 175.130 104.725 176.100 ;
        RECT 101.330 173.890 101.615 174.350 ;
        RECT 101.785 173.720 102.055 174.180 ;
        RECT 102.455 173.890 102.855 174.690 ;
        RECT 103.720 174.630 104.275 174.960 ;
        RECT 103.720 174.520 104.170 174.630 ;
        RECT 103.045 174.350 104.170 174.520 ;
        RECT 104.445 174.460 104.725 175.130 ;
        RECT 103.045 173.890 103.325 174.350 ;
        RECT 103.845 173.720 104.170 174.180 ;
        RECT 104.340 173.890 104.725 174.460 ;
        RECT 104.895 175.130 105.235 176.100 ;
        RECT 105.405 175.130 105.575 176.270 ;
        RECT 105.845 175.470 106.095 176.270 ;
        RECT 106.740 175.300 107.070 176.100 ;
        RECT 107.370 175.470 107.700 176.270 ;
        RECT 107.870 175.300 108.200 176.100 ;
        RECT 105.765 175.130 108.200 175.300 ;
        RECT 108.780 175.300 109.110 176.100 ;
        RECT 109.280 175.470 109.610 176.270 ;
        RECT 109.910 175.300 110.240 176.100 ;
        RECT 110.885 175.470 111.135 176.270 ;
        RECT 108.780 175.130 111.215 175.300 ;
        RECT 111.405 175.130 111.575 176.270 ;
        RECT 111.745 175.130 112.085 176.100 ;
        RECT 104.895 174.520 105.070 175.130 ;
        RECT 105.765 174.880 105.935 175.130 ;
        RECT 105.240 174.710 105.935 174.880 ;
        RECT 106.105 174.740 106.530 174.910 ;
        RECT 106.110 174.710 106.530 174.740 ;
        RECT 106.700 174.710 107.030 174.910 ;
        RECT 107.200 174.710 107.530 174.910 ;
        RECT 104.895 173.890 105.235 174.520 ;
        RECT 105.405 173.720 105.655 174.520 ;
        RECT 105.845 174.370 107.070 174.540 ;
        RECT 105.845 173.890 106.175 174.370 ;
        RECT 106.345 173.720 106.570 174.180 ;
        RECT 106.740 173.890 107.070 174.370 ;
        RECT 107.700 174.500 107.870 175.130 ;
        RECT 108.055 174.710 108.405 174.960 ;
        RECT 108.575 174.710 108.925 174.960 ;
        RECT 109.110 174.500 109.280 175.130 ;
        RECT 109.450 174.710 109.780 174.910 ;
        RECT 109.950 174.710 110.280 174.910 ;
        RECT 110.450 174.710 110.870 174.910 ;
        RECT 111.045 174.880 111.215 175.130 ;
        RECT 111.045 174.710 111.740 174.880 ;
        RECT 107.700 173.890 108.200 174.500 ;
        RECT 108.780 173.890 109.280 174.500 ;
        RECT 109.910 174.370 111.135 174.540 ;
        RECT 111.910 174.520 112.085 175.130 ;
        RECT 109.910 173.890 110.240 174.370 ;
        RECT 110.410 173.720 110.635 174.180 ;
        RECT 110.805 173.890 111.135 174.370 ;
        RECT 111.325 173.720 111.575 174.520 ;
        RECT 111.745 173.890 112.085 174.520 ;
        RECT 112.255 175.195 112.525 176.100 ;
        RECT 112.695 175.510 113.025 176.270 ;
        RECT 113.205 175.340 113.375 176.100 ;
        RECT 112.255 174.395 112.425 175.195 ;
        RECT 112.710 175.170 113.375 175.340 ;
        RECT 114.555 175.180 115.765 176.270 ;
        RECT 112.710 175.025 112.880 175.170 ;
        RECT 112.595 174.695 112.880 175.025 ;
        RECT 112.710 174.440 112.880 174.695 ;
        RECT 113.115 174.620 113.445 174.990 ;
        RECT 114.555 174.640 115.075 175.180 ;
        RECT 115.245 174.470 115.765 175.010 ;
        RECT 112.255 173.890 112.515 174.395 ;
        RECT 112.710 174.270 113.375 174.440 ;
        RECT 112.695 173.720 113.025 174.100 ;
        RECT 113.205 173.890 113.375 174.270 ;
        RECT 114.555 173.720 115.765 174.470 ;
        RECT 10.510 173.550 115.850 173.720 ;
        RECT 10.595 172.800 11.805 173.550 ;
        RECT 10.595 172.260 11.115 172.800 ;
        RECT 11.975 172.780 14.565 173.550 ;
        RECT 14.740 173.005 20.085 173.550 ;
        RECT 11.285 172.090 11.805 172.630 ;
        RECT 10.595 171.000 11.805 172.090 ;
        RECT 11.975 172.090 13.185 172.610 ;
        RECT 13.355 172.260 14.565 172.780 ;
        RECT 11.975 171.000 14.565 172.090 ;
        RECT 16.330 171.435 16.680 172.685 ;
        RECT 18.160 172.175 18.500 173.005 ;
        RECT 20.315 172.730 20.525 173.550 ;
        RECT 20.695 172.750 21.025 173.380 ;
        RECT 20.695 172.150 20.945 172.750 ;
        RECT 21.195 172.730 21.425 173.550 ;
        RECT 21.635 172.810 22.020 173.380 ;
        RECT 22.190 173.090 22.515 173.550 ;
        RECT 23.035 172.920 23.315 173.380 ;
        RECT 21.115 172.310 21.445 172.560 ;
        RECT 14.740 171.000 20.085 171.435 ;
        RECT 20.315 171.000 20.525 172.140 ;
        RECT 20.695 171.170 21.025 172.150 ;
        RECT 21.635 172.140 21.915 172.810 ;
        RECT 22.190 172.750 23.315 172.920 ;
        RECT 22.190 172.640 22.640 172.750 ;
        RECT 22.085 172.310 22.640 172.640 ;
        RECT 23.505 172.580 23.905 173.380 ;
        RECT 24.305 173.090 24.575 173.550 ;
        RECT 24.745 172.920 25.030 173.380 ;
        RECT 21.195 171.000 21.425 172.140 ;
        RECT 21.635 171.170 22.020 172.140 ;
        RECT 22.190 171.850 22.640 172.310 ;
        RECT 22.810 172.020 23.905 172.580 ;
        RECT 22.190 171.630 23.315 171.850 ;
        RECT 22.190 171.000 22.515 171.460 ;
        RECT 23.035 171.170 23.315 171.630 ;
        RECT 23.505 171.170 23.905 172.020 ;
        RECT 24.075 172.750 25.030 172.920 ;
        RECT 25.315 172.825 25.605 173.550 ;
        RECT 25.775 172.800 26.985 173.550 ;
        RECT 24.075 171.850 24.285 172.750 ;
        RECT 24.455 172.020 25.145 172.580 ;
        RECT 24.075 171.630 25.030 171.850 ;
        RECT 24.305 171.000 24.575 171.460 ;
        RECT 24.745 171.170 25.030 171.630 ;
        RECT 25.315 171.000 25.605 172.165 ;
        RECT 25.775 172.090 26.295 172.630 ;
        RECT 26.465 172.260 26.985 172.800 ;
        RECT 27.155 172.875 27.415 173.380 ;
        RECT 27.595 173.170 27.925 173.550 ;
        RECT 28.105 173.000 28.275 173.380 ;
        RECT 25.775 171.000 26.985 172.090 ;
        RECT 27.155 172.075 27.325 172.875 ;
        RECT 27.610 172.830 28.275 173.000 ;
        RECT 27.610 172.575 27.780 172.830 ;
        RECT 29.200 172.770 29.700 173.380 ;
        RECT 27.495 172.245 27.780 172.575 ;
        RECT 28.015 172.280 28.345 172.650 ;
        RECT 28.995 172.310 29.345 172.560 ;
        RECT 27.610 172.100 27.780 172.245 ;
        RECT 29.530 172.140 29.700 172.770 ;
        RECT 30.330 172.900 30.660 173.380 ;
        RECT 30.830 173.090 31.055 173.550 ;
        RECT 31.225 172.900 31.555 173.380 ;
        RECT 30.330 172.730 31.555 172.900 ;
        RECT 31.745 172.750 31.995 173.550 ;
        RECT 32.165 172.750 32.505 173.380 ;
        RECT 29.870 172.360 30.200 172.560 ;
        RECT 30.370 172.360 30.700 172.560 ;
        RECT 30.870 172.360 31.290 172.560 ;
        RECT 31.465 172.390 32.160 172.560 ;
        RECT 31.465 172.140 31.635 172.390 ;
        RECT 32.330 172.140 32.505 172.750 ;
        RECT 27.155 171.170 27.425 172.075 ;
        RECT 27.610 171.930 28.275 172.100 ;
        RECT 27.595 171.000 27.925 171.760 ;
        RECT 28.105 171.170 28.275 171.930 ;
        RECT 29.200 171.970 31.635 172.140 ;
        RECT 29.200 171.170 29.530 171.970 ;
        RECT 29.700 171.000 30.030 171.800 ;
        RECT 30.330 171.170 30.660 171.970 ;
        RECT 31.305 171.000 31.555 171.800 ;
        RECT 31.825 171.000 31.995 172.140 ;
        RECT 32.165 171.170 32.505 172.140 ;
        RECT 32.675 172.750 33.015 173.380 ;
        RECT 33.185 172.750 33.435 173.550 ;
        RECT 33.625 172.900 33.955 173.380 ;
        RECT 34.125 173.090 34.350 173.550 ;
        RECT 34.520 172.900 34.850 173.380 ;
        RECT 32.675 172.140 32.850 172.750 ;
        RECT 33.625 172.730 34.850 172.900 ;
        RECT 35.480 172.770 35.980 173.380 ;
        RECT 36.355 172.800 37.565 173.550 ;
        RECT 33.020 172.390 33.715 172.560 ;
        RECT 33.545 172.140 33.715 172.390 ;
        RECT 33.890 172.360 34.310 172.560 ;
        RECT 34.480 172.360 34.810 172.560 ;
        RECT 34.980 172.360 35.310 172.560 ;
        RECT 35.480 172.140 35.650 172.770 ;
        RECT 35.835 172.310 36.185 172.560 ;
        RECT 32.675 171.170 33.015 172.140 ;
        RECT 33.185 171.000 33.355 172.140 ;
        RECT 33.545 171.970 35.980 172.140 ;
        RECT 33.625 171.000 33.875 171.800 ;
        RECT 34.520 171.170 34.850 171.970 ;
        RECT 35.150 171.000 35.480 171.800 ;
        RECT 35.650 171.170 35.980 171.970 ;
        RECT 36.355 172.090 36.875 172.630 ;
        RECT 37.045 172.260 37.565 172.800 ;
        RECT 37.735 172.750 38.075 173.380 ;
        RECT 38.245 172.750 38.495 173.550 ;
        RECT 38.685 172.900 39.015 173.380 ;
        RECT 39.185 173.090 39.410 173.550 ;
        RECT 39.580 172.900 39.910 173.380 ;
        RECT 37.735 172.140 37.910 172.750 ;
        RECT 38.685 172.730 39.910 172.900 ;
        RECT 40.540 172.770 41.040 173.380 ;
        RECT 41.505 173.070 41.805 173.550 ;
        RECT 41.975 172.900 42.235 173.355 ;
        RECT 42.405 173.070 42.665 173.550 ;
        RECT 42.845 172.900 43.105 173.355 ;
        RECT 43.275 173.070 43.525 173.550 ;
        RECT 43.705 172.900 43.965 173.355 ;
        RECT 44.135 173.070 44.385 173.550 ;
        RECT 44.565 172.900 44.825 173.355 ;
        RECT 44.995 173.070 45.240 173.550 ;
        RECT 45.410 172.900 45.685 173.355 ;
        RECT 45.855 173.070 46.100 173.550 ;
        RECT 46.270 172.900 46.530 173.355 ;
        RECT 46.700 173.070 46.960 173.550 ;
        RECT 47.130 172.900 47.390 173.355 ;
        RECT 47.560 173.070 47.820 173.550 ;
        RECT 47.990 172.900 48.250 173.355 ;
        RECT 48.420 172.990 48.680 173.550 ;
        RECT 38.080 172.390 38.775 172.560 ;
        RECT 38.605 172.140 38.775 172.390 ;
        RECT 38.950 172.360 39.370 172.560 ;
        RECT 39.540 172.360 39.870 172.560 ;
        RECT 40.040 172.360 40.370 172.560 ;
        RECT 40.540 172.140 40.710 172.770 ;
        RECT 41.505 172.730 48.250 172.900 ;
        RECT 40.895 172.310 41.245 172.560 ;
        RECT 41.505 172.140 42.670 172.730 ;
        RECT 48.850 172.560 49.100 173.370 ;
        RECT 49.280 173.025 49.540 173.550 ;
        RECT 49.710 172.560 49.960 173.370 ;
        RECT 50.140 173.040 50.445 173.550 ;
        RECT 42.840 172.310 49.960 172.560 ;
        RECT 50.130 172.310 50.445 172.870 ;
        RECT 51.075 172.825 51.365 173.550 ;
        RECT 51.540 172.840 51.795 173.370 ;
        RECT 51.965 173.090 52.270 173.550 ;
        RECT 52.515 173.170 53.585 173.340 ;
        RECT 36.355 171.000 37.565 172.090 ;
        RECT 37.735 171.170 38.075 172.140 ;
        RECT 38.245 171.000 38.415 172.140 ;
        RECT 38.605 171.970 41.040 172.140 ;
        RECT 38.685 171.000 38.935 171.800 ;
        RECT 39.580 171.170 39.910 171.970 ;
        RECT 40.210 171.000 40.540 171.800 ;
        RECT 40.710 171.170 41.040 171.970 ;
        RECT 41.505 171.915 48.250 172.140 ;
        RECT 41.505 171.000 41.775 171.745 ;
        RECT 41.945 171.175 42.235 171.915 ;
        RECT 42.845 171.900 48.250 171.915 ;
        RECT 42.405 171.005 42.660 171.730 ;
        RECT 42.845 171.175 43.105 171.900 ;
        RECT 43.275 171.005 43.520 171.730 ;
        RECT 43.705 171.175 43.965 171.900 ;
        RECT 44.135 171.005 44.380 171.730 ;
        RECT 44.565 171.175 44.825 171.900 ;
        RECT 44.995 171.005 45.240 171.730 ;
        RECT 45.410 171.175 45.670 171.900 ;
        RECT 45.840 171.005 46.100 171.730 ;
        RECT 46.270 171.175 46.530 171.900 ;
        RECT 46.700 171.005 46.960 171.730 ;
        RECT 47.130 171.175 47.390 171.900 ;
        RECT 47.560 171.005 47.820 171.730 ;
        RECT 47.990 171.175 48.250 171.900 ;
        RECT 48.420 171.005 48.680 171.800 ;
        RECT 48.850 171.175 49.100 172.310 ;
        RECT 42.405 171.000 48.680 171.005 ;
        RECT 49.280 171.000 49.540 171.810 ;
        RECT 49.715 171.170 49.960 172.310 ;
        RECT 51.540 172.190 51.750 172.840 ;
        RECT 52.515 172.815 52.835 173.170 ;
        RECT 52.510 172.640 52.835 172.815 ;
        RECT 51.920 172.340 52.835 172.640 ;
        RECT 53.005 172.600 53.245 173.000 ;
        RECT 53.415 172.940 53.585 173.170 ;
        RECT 53.755 173.110 53.945 173.550 ;
        RECT 54.115 173.100 55.065 173.380 ;
        RECT 55.285 173.190 55.635 173.360 ;
        RECT 53.415 172.770 53.945 172.940 ;
        RECT 51.920 172.310 52.660 172.340 ;
        RECT 50.140 171.000 50.435 171.810 ;
        RECT 51.075 171.000 51.365 172.165 ;
        RECT 51.540 171.310 51.795 172.190 ;
        RECT 51.965 171.000 52.270 172.140 ;
        RECT 52.490 171.720 52.660 172.310 ;
        RECT 53.005 172.230 53.545 172.600 ;
        RECT 53.725 172.490 53.945 172.770 ;
        RECT 54.115 172.320 54.285 173.100 ;
        RECT 53.880 172.150 54.285 172.320 ;
        RECT 54.455 172.310 54.805 172.930 ;
        RECT 53.880 172.060 54.050 172.150 ;
        RECT 54.975 172.140 55.185 172.930 ;
        RECT 52.830 171.890 54.050 172.060 ;
        RECT 54.510 171.980 55.185 172.140 ;
        RECT 52.490 171.550 53.290 171.720 ;
        RECT 52.610 171.000 52.940 171.380 ;
        RECT 53.120 171.260 53.290 171.550 ;
        RECT 53.880 171.510 54.050 171.890 ;
        RECT 54.220 171.970 55.185 171.980 ;
        RECT 55.375 172.800 55.635 173.190 ;
        RECT 55.845 173.090 56.175 173.550 ;
        RECT 57.050 173.160 57.905 173.330 ;
        RECT 58.110 173.160 58.605 173.330 ;
        RECT 58.775 173.190 59.105 173.550 ;
        RECT 55.375 172.110 55.545 172.800 ;
        RECT 55.715 172.450 55.885 172.630 ;
        RECT 56.055 172.620 56.845 172.870 ;
        RECT 57.050 172.450 57.220 173.160 ;
        RECT 57.390 172.650 57.745 172.870 ;
        RECT 55.715 172.280 57.405 172.450 ;
        RECT 54.220 171.680 54.680 171.970 ;
        RECT 55.375 171.940 56.875 172.110 ;
        RECT 55.375 171.800 55.545 171.940 ;
        RECT 54.985 171.630 55.545 171.800 ;
        RECT 53.460 171.000 53.710 171.460 ;
        RECT 53.880 171.170 54.750 171.510 ;
        RECT 54.985 171.170 55.155 171.630 ;
        RECT 55.990 171.600 57.065 171.770 ;
        RECT 55.325 171.000 55.695 171.460 ;
        RECT 55.990 171.260 56.160 171.600 ;
        RECT 56.330 171.000 56.660 171.430 ;
        RECT 56.895 171.260 57.065 171.600 ;
        RECT 57.235 171.500 57.405 172.280 ;
        RECT 57.575 172.060 57.745 172.650 ;
        RECT 57.915 172.250 58.265 172.870 ;
        RECT 57.575 171.670 58.040 172.060 ;
        RECT 58.435 171.800 58.605 173.160 ;
        RECT 58.775 171.970 59.235 173.020 ;
        RECT 58.210 171.630 58.605 171.800 ;
        RECT 58.210 171.500 58.380 171.630 ;
        RECT 57.235 171.170 57.915 171.500 ;
        RECT 58.130 171.170 58.380 171.500 ;
        RECT 58.550 171.000 58.800 171.460 ;
        RECT 58.970 171.185 59.295 171.970 ;
        RECT 59.465 171.170 59.635 173.290 ;
        RECT 59.805 173.170 60.135 173.550 ;
        RECT 60.305 173.000 60.560 173.290 ;
        RECT 59.810 172.830 60.560 173.000 ;
        RECT 59.810 171.840 60.040 172.830 ;
        RECT 61.655 172.780 65.165 173.550 ;
        RECT 65.340 173.005 70.685 173.550 ;
        RECT 60.210 172.010 60.560 172.660 ;
        RECT 61.655 172.090 63.345 172.610 ;
        RECT 63.515 172.260 65.165 172.780 ;
        RECT 59.810 171.670 60.560 171.840 ;
        RECT 59.805 171.000 60.135 171.500 ;
        RECT 60.305 171.170 60.560 171.670 ;
        RECT 61.655 171.000 65.165 172.090 ;
        RECT 66.930 171.435 67.280 172.685 ;
        RECT 68.760 172.175 69.100 173.005 ;
        RECT 70.855 172.750 71.195 173.380 ;
        RECT 71.365 172.750 71.615 173.550 ;
        RECT 71.805 172.900 72.135 173.380 ;
        RECT 72.305 173.090 72.530 173.550 ;
        RECT 72.700 172.900 73.030 173.380 ;
        RECT 70.855 172.140 71.030 172.750 ;
        RECT 71.805 172.730 73.030 172.900 ;
        RECT 73.660 172.770 74.160 173.380 ;
        RECT 74.995 172.780 76.665 173.550 ;
        RECT 76.835 172.825 77.125 173.550 ;
        RECT 77.755 172.780 81.265 173.550 ;
        RECT 71.200 172.390 71.895 172.560 ;
        RECT 71.725 172.140 71.895 172.390 ;
        RECT 72.070 172.360 72.490 172.560 ;
        RECT 72.660 172.360 72.990 172.560 ;
        RECT 73.160 172.360 73.490 172.560 ;
        RECT 73.660 172.140 73.830 172.770 ;
        RECT 74.015 172.310 74.365 172.560 ;
        RECT 65.340 171.000 70.685 171.435 ;
        RECT 70.855 171.170 71.195 172.140 ;
        RECT 71.365 171.000 71.535 172.140 ;
        RECT 71.725 171.970 74.160 172.140 ;
        RECT 71.805 171.000 72.055 171.800 ;
        RECT 72.700 171.170 73.030 171.970 ;
        RECT 73.330 171.000 73.660 171.800 ;
        RECT 73.830 171.170 74.160 171.970 ;
        RECT 74.995 172.090 75.745 172.610 ;
        RECT 75.915 172.260 76.665 172.780 ;
        RECT 74.995 171.000 76.665 172.090 ;
        RECT 76.835 171.000 77.125 172.165 ;
        RECT 77.755 172.090 79.445 172.610 ;
        RECT 79.615 172.260 81.265 172.780 ;
        RECT 81.475 172.730 81.705 173.550 ;
        RECT 81.875 172.750 82.205 173.380 ;
        RECT 81.455 172.310 81.785 172.560 ;
        RECT 81.955 172.150 82.205 172.750 ;
        RECT 82.375 172.730 82.585 173.550 ;
        RECT 82.820 173.000 83.075 173.290 ;
        RECT 83.245 173.170 83.575 173.550 ;
        RECT 82.820 172.830 83.570 173.000 ;
        RECT 77.755 171.000 81.265 172.090 ;
        RECT 81.475 171.000 81.705 172.140 ;
        RECT 81.875 171.170 82.205 172.150 ;
        RECT 82.375 171.000 82.585 172.140 ;
        RECT 82.820 172.010 83.170 172.660 ;
        RECT 83.340 171.840 83.570 172.830 ;
        RECT 82.820 171.670 83.570 171.840 ;
        RECT 82.820 171.170 83.075 171.670 ;
        RECT 83.245 171.000 83.575 171.500 ;
        RECT 83.745 171.170 83.915 173.290 ;
        RECT 84.275 173.190 84.605 173.550 ;
        RECT 84.775 173.160 85.270 173.330 ;
        RECT 85.475 173.160 86.330 173.330 ;
        RECT 84.145 171.970 84.605 173.020 ;
        RECT 84.085 171.185 84.410 171.970 ;
        RECT 84.775 171.800 84.945 173.160 ;
        RECT 85.115 172.250 85.465 172.870 ;
        RECT 85.635 172.650 85.990 172.870 ;
        RECT 85.635 172.060 85.805 172.650 ;
        RECT 86.160 172.450 86.330 173.160 ;
        RECT 87.205 173.090 87.535 173.550 ;
        RECT 87.745 173.190 88.095 173.360 ;
        RECT 86.535 172.620 87.325 172.870 ;
        RECT 87.745 172.800 88.005 173.190 ;
        RECT 88.315 173.100 89.265 173.380 ;
        RECT 89.435 173.110 89.625 173.550 ;
        RECT 89.795 173.170 90.865 173.340 ;
        RECT 87.495 172.450 87.665 172.630 ;
        RECT 84.775 171.630 85.170 171.800 ;
        RECT 85.340 171.670 85.805 172.060 ;
        RECT 85.975 172.280 87.665 172.450 ;
        RECT 85.000 171.500 85.170 171.630 ;
        RECT 85.975 171.500 86.145 172.280 ;
        RECT 87.835 172.110 88.005 172.800 ;
        RECT 86.505 171.940 88.005 172.110 ;
        RECT 88.195 172.140 88.405 172.930 ;
        RECT 88.575 172.310 88.925 172.930 ;
        RECT 89.095 172.320 89.265 173.100 ;
        RECT 89.795 172.940 89.965 173.170 ;
        RECT 89.435 172.770 89.965 172.940 ;
        RECT 89.435 172.490 89.655 172.770 ;
        RECT 90.135 172.600 90.375 173.000 ;
        RECT 89.095 172.150 89.500 172.320 ;
        RECT 89.835 172.230 90.375 172.600 ;
        RECT 90.545 172.815 90.865 173.170 ;
        RECT 91.110 173.090 91.415 173.550 ;
        RECT 91.585 172.840 91.840 173.370 ;
        RECT 90.545 172.640 90.870 172.815 ;
        RECT 90.545 172.340 91.460 172.640 ;
        RECT 90.720 172.310 91.460 172.340 ;
        RECT 88.195 171.980 88.870 172.140 ;
        RECT 89.330 172.060 89.500 172.150 ;
        RECT 88.195 171.970 89.160 171.980 ;
        RECT 87.835 171.800 88.005 171.940 ;
        RECT 84.580 171.000 84.830 171.460 ;
        RECT 85.000 171.170 85.250 171.500 ;
        RECT 85.465 171.170 86.145 171.500 ;
        RECT 86.315 171.600 87.390 171.770 ;
        RECT 87.835 171.630 88.395 171.800 ;
        RECT 88.700 171.680 89.160 171.970 ;
        RECT 89.330 171.890 90.550 172.060 ;
        RECT 86.315 171.260 86.485 171.600 ;
        RECT 86.720 171.000 87.050 171.430 ;
        RECT 87.220 171.260 87.390 171.600 ;
        RECT 87.685 171.000 88.055 171.460 ;
        RECT 88.225 171.170 88.395 171.630 ;
        RECT 89.330 171.510 89.500 171.890 ;
        RECT 90.720 171.720 90.890 172.310 ;
        RECT 91.630 172.190 91.840 172.840 ;
        RECT 88.630 171.170 89.500 171.510 ;
        RECT 90.090 171.550 90.890 171.720 ;
        RECT 89.670 171.000 89.920 171.460 ;
        RECT 90.090 171.260 90.260 171.550 ;
        RECT 90.440 171.000 90.770 171.380 ;
        RECT 91.110 171.000 91.415 172.140 ;
        RECT 91.585 171.310 91.840 172.190 ;
        RECT 92.015 172.810 92.400 173.380 ;
        RECT 92.570 173.090 92.895 173.550 ;
        RECT 93.415 172.920 93.695 173.380 ;
        RECT 92.015 172.140 92.295 172.810 ;
        RECT 92.570 172.750 93.695 172.920 ;
        RECT 92.570 172.640 93.020 172.750 ;
        RECT 92.465 172.310 93.020 172.640 ;
        RECT 93.885 172.580 94.285 173.380 ;
        RECT 94.685 173.090 94.955 173.550 ;
        RECT 95.125 172.920 95.410 173.380 ;
        RECT 92.015 171.170 92.400 172.140 ;
        RECT 92.570 171.850 93.020 172.310 ;
        RECT 93.190 172.020 94.285 172.580 ;
        RECT 92.570 171.630 93.695 171.850 ;
        RECT 92.570 171.000 92.895 171.460 ;
        RECT 93.415 171.170 93.695 171.630 ;
        RECT 93.885 171.170 94.285 172.020 ;
        RECT 94.455 172.750 95.410 172.920 ;
        RECT 95.695 172.780 98.285 173.550 ;
        RECT 94.455 171.850 94.665 172.750 ;
        RECT 94.835 172.020 95.525 172.580 ;
        RECT 95.695 172.090 96.905 172.610 ;
        RECT 97.075 172.260 98.285 172.780 ;
        RECT 98.730 172.740 98.975 173.345 ;
        RECT 99.195 173.015 99.705 173.550 ;
        RECT 98.455 172.570 99.685 172.740 ;
        RECT 94.455 171.630 95.410 171.850 ;
        RECT 94.685 171.000 94.955 171.460 ;
        RECT 95.125 171.170 95.410 171.630 ;
        RECT 95.695 171.000 98.285 172.090 ;
        RECT 98.455 171.760 98.795 172.570 ;
        RECT 98.965 172.005 99.715 172.195 ;
        RECT 98.455 171.350 98.970 171.760 ;
        RECT 99.205 171.000 99.375 171.760 ;
        RECT 99.545 171.340 99.715 172.005 ;
        RECT 99.885 172.020 100.075 173.380 ;
        RECT 100.245 172.530 100.520 173.380 ;
        RECT 100.710 173.015 101.240 173.380 ;
        RECT 101.665 173.150 101.995 173.550 ;
        RECT 101.065 172.980 101.240 173.015 ;
        RECT 100.245 172.360 100.525 172.530 ;
        RECT 100.245 172.220 100.520 172.360 ;
        RECT 100.725 172.020 100.895 172.820 ;
        RECT 99.885 171.850 100.895 172.020 ;
        RECT 101.065 172.810 101.995 172.980 ;
        RECT 102.165 172.810 102.420 173.380 ;
        RECT 102.595 172.825 102.885 173.550 ;
        RECT 101.065 171.680 101.235 172.810 ;
        RECT 101.825 172.640 101.995 172.810 ;
        RECT 100.110 171.510 101.235 171.680 ;
        RECT 101.405 172.310 101.600 172.640 ;
        RECT 101.825 172.310 102.080 172.640 ;
        RECT 101.405 171.340 101.575 172.310 ;
        RECT 102.250 172.140 102.420 172.810 ;
        RECT 103.095 172.730 103.325 173.550 ;
        RECT 103.495 172.750 103.825 173.380 ;
        RECT 103.075 172.310 103.405 172.560 ;
        RECT 99.545 171.170 101.575 171.340 ;
        RECT 101.745 171.000 101.915 172.140 ;
        RECT 102.085 171.170 102.420 172.140 ;
        RECT 102.595 171.000 102.885 172.165 ;
        RECT 103.575 172.150 103.825 172.750 ;
        RECT 103.995 172.730 104.205 173.550 ;
        RECT 104.440 172.840 104.695 173.370 ;
        RECT 104.865 173.090 105.170 173.550 ;
        RECT 105.415 173.170 106.485 173.340 ;
        RECT 103.095 171.000 103.325 172.140 ;
        RECT 103.495 171.170 103.825 172.150 ;
        RECT 104.440 172.190 104.650 172.840 ;
        RECT 105.415 172.815 105.735 173.170 ;
        RECT 105.410 172.640 105.735 172.815 ;
        RECT 104.820 172.340 105.735 172.640 ;
        RECT 105.905 172.600 106.145 173.000 ;
        RECT 106.315 172.940 106.485 173.170 ;
        RECT 106.655 173.110 106.845 173.550 ;
        RECT 107.015 173.100 107.965 173.380 ;
        RECT 108.185 173.190 108.535 173.360 ;
        RECT 106.315 172.770 106.845 172.940 ;
        RECT 104.820 172.310 105.560 172.340 ;
        RECT 103.995 171.000 104.205 172.140 ;
        RECT 104.440 171.310 104.695 172.190 ;
        RECT 104.865 171.000 105.170 172.140 ;
        RECT 105.390 171.720 105.560 172.310 ;
        RECT 105.905 172.230 106.445 172.600 ;
        RECT 106.625 172.490 106.845 172.770 ;
        RECT 107.015 172.320 107.185 173.100 ;
        RECT 106.780 172.150 107.185 172.320 ;
        RECT 107.355 172.310 107.705 172.930 ;
        RECT 106.780 172.060 106.950 172.150 ;
        RECT 107.875 172.140 108.085 172.930 ;
        RECT 105.730 171.890 106.950 172.060 ;
        RECT 107.410 171.980 108.085 172.140 ;
        RECT 105.390 171.550 106.190 171.720 ;
        RECT 105.510 171.000 105.840 171.380 ;
        RECT 106.020 171.260 106.190 171.550 ;
        RECT 106.780 171.510 106.950 171.890 ;
        RECT 107.120 171.970 108.085 171.980 ;
        RECT 108.275 172.800 108.535 173.190 ;
        RECT 108.745 173.090 109.075 173.550 ;
        RECT 109.950 173.160 110.805 173.330 ;
        RECT 111.010 173.160 111.505 173.330 ;
        RECT 111.675 173.190 112.005 173.550 ;
        RECT 108.275 172.110 108.445 172.800 ;
        RECT 108.615 172.450 108.785 172.630 ;
        RECT 108.955 172.620 109.745 172.870 ;
        RECT 109.950 172.450 110.120 173.160 ;
        RECT 110.290 172.650 110.645 172.870 ;
        RECT 108.615 172.280 110.305 172.450 ;
        RECT 107.120 171.680 107.580 171.970 ;
        RECT 108.275 171.940 109.775 172.110 ;
        RECT 108.275 171.800 108.445 171.940 ;
        RECT 107.885 171.630 108.445 171.800 ;
        RECT 106.360 171.000 106.610 171.460 ;
        RECT 106.780 171.170 107.650 171.510 ;
        RECT 107.885 171.170 108.055 171.630 ;
        RECT 108.890 171.600 109.965 171.770 ;
        RECT 108.225 171.000 108.595 171.460 ;
        RECT 108.890 171.260 109.060 171.600 ;
        RECT 109.230 171.000 109.560 171.430 ;
        RECT 109.795 171.260 109.965 171.600 ;
        RECT 110.135 171.500 110.305 172.280 ;
        RECT 110.475 172.060 110.645 172.650 ;
        RECT 110.815 172.250 111.165 172.870 ;
        RECT 110.475 171.670 110.940 172.060 ;
        RECT 111.335 171.800 111.505 173.160 ;
        RECT 111.675 171.970 112.135 173.020 ;
        RECT 111.110 171.630 111.505 171.800 ;
        RECT 111.110 171.500 111.280 171.630 ;
        RECT 110.135 171.170 110.815 171.500 ;
        RECT 111.030 171.170 111.280 171.500 ;
        RECT 111.450 171.000 111.700 171.460 ;
        RECT 111.870 171.185 112.195 171.970 ;
        RECT 112.365 171.170 112.535 173.290 ;
        RECT 112.705 173.170 113.035 173.550 ;
        RECT 113.205 173.000 113.460 173.290 ;
        RECT 112.710 172.830 113.460 173.000 ;
        RECT 112.710 171.840 112.940 172.830 ;
        RECT 114.555 172.800 115.765 173.550 ;
        RECT 113.110 172.010 113.460 172.660 ;
        RECT 114.555 172.090 115.075 172.630 ;
        RECT 115.245 172.260 115.765 172.800 ;
        RECT 112.710 171.670 113.460 171.840 ;
        RECT 112.705 171.000 113.035 171.500 ;
        RECT 113.205 171.170 113.460 171.670 ;
        RECT 114.555 171.000 115.765 172.090 ;
        RECT 10.510 170.830 115.850 171.000 ;
        RECT 10.595 169.740 11.805 170.830 ;
        RECT 10.595 169.030 11.115 169.570 ;
        RECT 11.285 169.200 11.805 169.740 ;
        RECT 12.435 169.665 12.725 170.830 ;
        RECT 13.355 169.740 15.945 170.830 ;
        RECT 16.120 170.395 21.465 170.830 ;
        RECT 13.355 169.220 14.565 169.740 ;
        RECT 14.735 169.050 15.945 169.570 ;
        RECT 17.710 169.145 18.060 170.395 ;
        RECT 21.725 170.085 21.995 170.830 ;
        RECT 22.625 170.825 28.900 170.830 ;
        RECT 22.165 169.915 22.455 170.655 ;
        RECT 22.625 170.100 22.880 170.825 ;
        RECT 23.065 169.930 23.325 170.655 ;
        RECT 23.495 170.100 23.740 170.825 ;
        RECT 23.925 169.930 24.185 170.655 ;
        RECT 24.355 170.100 24.600 170.825 ;
        RECT 24.785 169.930 25.045 170.655 ;
        RECT 25.215 170.100 25.460 170.825 ;
        RECT 25.630 169.930 25.890 170.655 ;
        RECT 26.060 170.100 26.320 170.825 ;
        RECT 26.490 169.930 26.750 170.655 ;
        RECT 26.920 170.100 27.180 170.825 ;
        RECT 27.350 169.930 27.610 170.655 ;
        RECT 27.780 170.100 28.040 170.825 ;
        RECT 28.210 169.930 28.470 170.655 ;
        RECT 28.640 170.030 28.900 170.825 ;
        RECT 23.065 169.915 28.470 169.930 ;
        RECT 21.725 169.690 28.470 169.915 ;
        RECT 10.595 168.280 11.805 169.030 ;
        RECT 12.435 168.280 12.725 169.005 ;
        RECT 13.355 168.280 15.945 169.050 ;
        RECT 19.540 168.825 19.880 169.655 ;
        RECT 21.725 169.100 22.890 169.690 ;
        RECT 29.070 169.520 29.320 170.655 ;
        RECT 29.500 170.020 29.760 170.830 ;
        RECT 29.935 169.520 30.180 170.660 ;
        RECT 30.360 170.020 30.655 170.830 ;
        RECT 31.815 169.690 32.025 170.830 ;
        RECT 32.195 169.680 32.525 170.660 ;
        RECT 32.695 169.690 32.925 170.830 ;
        RECT 33.595 169.740 36.185 170.830 ;
        RECT 23.060 169.270 30.180 169.520 ;
        RECT 21.725 168.930 28.470 169.100 ;
        RECT 16.120 168.280 21.465 168.825 ;
        RECT 21.725 168.280 22.025 168.760 ;
        RECT 22.195 168.475 22.455 168.930 ;
        RECT 22.625 168.280 22.885 168.760 ;
        RECT 23.065 168.475 23.325 168.930 ;
        RECT 23.495 168.280 23.745 168.760 ;
        RECT 23.925 168.475 24.185 168.930 ;
        RECT 24.355 168.280 24.605 168.760 ;
        RECT 24.785 168.475 25.045 168.930 ;
        RECT 25.215 168.280 25.460 168.760 ;
        RECT 25.630 168.475 25.905 168.930 ;
        RECT 26.075 168.280 26.320 168.760 ;
        RECT 26.490 168.475 26.750 168.930 ;
        RECT 26.920 168.280 27.180 168.760 ;
        RECT 27.350 168.475 27.610 168.930 ;
        RECT 27.780 168.280 28.040 168.760 ;
        RECT 28.210 168.475 28.470 168.930 ;
        RECT 28.640 168.280 28.900 168.840 ;
        RECT 29.070 168.460 29.320 169.270 ;
        RECT 29.500 168.280 29.760 168.805 ;
        RECT 29.930 168.460 30.180 169.270 ;
        RECT 30.350 168.960 30.665 169.520 ;
        RECT 30.360 168.280 30.665 168.790 ;
        RECT 31.815 168.280 32.025 169.100 ;
        RECT 32.195 169.080 32.445 169.680 ;
        RECT 32.615 169.270 32.945 169.520 ;
        RECT 33.595 169.220 34.805 169.740 ;
        RECT 36.395 169.690 36.625 170.830 ;
        RECT 36.795 169.680 37.125 170.660 ;
        RECT 37.295 169.690 37.505 170.830 ;
        RECT 32.195 168.450 32.525 169.080 ;
        RECT 32.695 168.280 32.925 169.100 ;
        RECT 34.975 169.050 36.185 169.570 ;
        RECT 36.375 169.270 36.705 169.520 ;
        RECT 33.595 168.280 36.185 169.050 ;
        RECT 36.395 168.280 36.625 169.100 ;
        RECT 36.875 169.080 37.125 169.680 ;
        RECT 38.195 169.665 38.485 170.830 ;
        RECT 39.115 169.740 41.705 170.830 ;
        RECT 39.115 169.220 40.325 169.740 ;
        RECT 41.875 169.690 42.260 170.660 ;
        RECT 42.430 170.370 42.755 170.830 ;
        RECT 43.275 170.200 43.555 170.660 ;
        RECT 42.430 169.980 43.555 170.200 ;
        RECT 36.795 168.450 37.125 169.080 ;
        RECT 37.295 168.280 37.505 169.100 ;
        RECT 40.495 169.050 41.705 169.570 ;
        RECT 38.195 168.280 38.485 169.005 ;
        RECT 39.115 168.280 41.705 169.050 ;
        RECT 41.875 169.020 42.155 169.690 ;
        RECT 42.430 169.520 42.880 169.980 ;
        RECT 43.745 169.810 44.145 170.660 ;
        RECT 44.545 170.370 44.815 170.830 ;
        RECT 44.985 170.200 45.270 170.660 ;
        RECT 42.325 169.190 42.880 169.520 ;
        RECT 43.050 169.250 44.145 169.810 ;
        RECT 42.430 169.080 42.880 169.190 ;
        RECT 41.875 168.450 42.260 169.020 ;
        RECT 42.430 168.910 43.555 169.080 ;
        RECT 42.430 168.280 42.755 168.740 ;
        RECT 43.275 168.450 43.555 168.910 ;
        RECT 43.745 168.450 44.145 169.250 ;
        RECT 44.315 169.980 45.270 170.200 ;
        RECT 45.615 169.995 45.870 170.830 ;
        RECT 44.315 169.080 44.525 169.980 ;
        RECT 46.040 169.825 46.300 170.630 ;
        RECT 46.470 169.995 46.730 170.830 ;
        RECT 46.900 169.825 47.155 170.630 ;
        RECT 44.695 169.250 45.385 169.810 ;
        RECT 45.555 169.655 47.155 169.825 ;
        RECT 45.555 169.090 45.835 169.655 ;
        RECT 47.400 169.640 47.655 170.520 ;
        RECT 47.825 169.690 48.130 170.830 ;
        RECT 48.470 170.450 48.800 170.830 ;
        RECT 48.980 170.280 49.150 170.570 ;
        RECT 49.320 170.370 49.570 170.830 ;
        RECT 48.350 170.110 49.150 170.280 ;
        RECT 49.740 170.320 50.610 170.660 ;
        RECT 46.005 169.260 47.225 169.485 ;
        RECT 44.315 168.910 45.270 169.080 ;
        RECT 45.555 168.920 46.285 169.090 ;
        RECT 44.545 168.280 44.815 168.740 ;
        RECT 44.985 168.450 45.270 168.910 ;
        RECT 45.560 168.280 45.890 168.750 ;
        RECT 46.060 168.475 46.285 168.920 ;
        RECT 47.400 168.990 47.610 169.640 ;
        RECT 48.350 169.520 48.520 170.110 ;
        RECT 49.740 169.940 49.910 170.320 ;
        RECT 50.845 170.200 51.015 170.660 ;
        RECT 51.185 170.370 51.555 170.830 ;
        RECT 51.850 170.230 52.020 170.570 ;
        RECT 52.190 170.400 52.520 170.830 ;
        RECT 52.755 170.230 52.925 170.570 ;
        RECT 48.690 169.770 49.910 169.940 ;
        RECT 50.080 169.860 50.540 170.150 ;
        RECT 50.845 170.030 51.405 170.200 ;
        RECT 51.850 170.060 52.925 170.230 ;
        RECT 53.095 170.330 53.775 170.660 ;
        RECT 53.990 170.330 54.240 170.660 ;
        RECT 54.410 170.370 54.660 170.830 ;
        RECT 51.235 169.890 51.405 170.030 ;
        RECT 50.080 169.850 51.045 169.860 ;
        RECT 49.740 169.680 49.910 169.770 ;
        RECT 50.370 169.690 51.045 169.850 ;
        RECT 47.780 169.490 48.520 169.520 ;
        RECT 47.780 169.190 48.695 169.490 ;
        RECT 48.370 169.015 48.695 169.190 ;
        RECT 46.455 168.280 46.750 168.805 ;
        RECT 47.400 168.460 47.655 168.990 ;
        RECT 47.825 168.280 48.130 168.740 ;
        RECT 48.375 168.660 48.695 169.015 ;
        RECT 48.865 169.230 49.405 169.600 ;
        RECT 49.740 169.510 50.145 169.680 ;
        RECT 48.865 168.830 49.105 169.230 ;
        RECT 49.585 169.060 49.805 169.340 ;
        RECT 49.275 168.890 49.805 169.060 ;
        RECT 49.275 168.660 49.445 168.890 ;
        RECT 49.975 168.730 50.145 169.510 ;
        RECT 50.315 168.900 50.665 169.520 ;
        RECT 50.835 168.900 51.045 169.690 ;
        RECT 51.235 169.720 52.735 169.890 ;
        RECT 51.235 169.030 51.405 169.720 ;
        RECT 53.095 169.550 53.265 170.330 ;
        RECT 54.070 170.200 54.240 170.330 ;
        RECT 51.575 169.380 53.265 169.550 ;
        RECT 53.435 169.770 53.900 170.160 ;
        RECT 54.070 170.030 54.465 170.200 ;
        RECT 51.575 169.200 51.745 169.380 ;
        RECT 48.375 168.490 49.445 168.660 ;
        RECT 49.615 168.280 49.805 168.720 ;
        RECT 49.975 168.450 50.925 168.730 ;
        RECT 51.235 168.640 51.495 169.030 ;
        RECT 51.915 168.960 52.705 169.210 ;
        RECT 51.145 168.470 51.495 168.640 ;
        RECT 51.705 168.280 52.035 168.740 ;
        RECT 52.910 168.670 53.080 169.380 ;
        RECT 53.435 169.180 53.605 169.770 ;
        RECT 53.250 168.960 53.605 169.180 ;
        RECT 53.775 168.960 54.125 169.580 ;
        RECT 54.295 168.670 54.465 170.030 ;
        RECT 54.830 169.860 55.155 170.645 ;
        RECT 54.635 168.810 55.095 169.860 ;
        RECT 52.910 168.500 53.765 168.670 ;
        RECT 53.970 168.500 54.465 168.670 ;
        RECT 54.635 168.280 54.965 168.640 ;
        RECT 55.325 168.540 55.495 170.660 ;
        RECT 55.665 170.330 55.995 170.830 ;
        RECT 56.165 170.160 56.420 170.660 ;
        RECT 55.670 169.990 56.420 170.160 ;
        RECT 55.670 169.000 55.900 169.990 ;
        RECT 56.070 169.170 56.420 169.820 ;
        RECT 56.595 169.740 60.105 170.830 ;
        RECT 56.595 169.220 58.285 169.740 ;
        RECT 60.280 169.680 60.540 170.830 ;
        RECT 60.715 169.755 60.970 170.660 ;
        RECT 61.140 170.070 61.470 170.830 ;
        RECT 61.685 169.900 61.855 170.660 ;
        RECT 58.455 169.050 60.105 169.570 ;
        RECT 55.670 168.830 56.420 169.000 ;
        RECT 55.665 168.280 55.995 168.660 ;
        RECT 56.165 168.540 56.420 168.830 ;
        RECT 56.595 168.280 60.105 169.050 ;
        RECT 60.280 168.280 60.540 169.120 ;
        RECT 60.715 169.025 60.885 169.755 ;
        RECT 61.140 169.730 61.855 169.900 ;
        RECT 61.140 169.520 61.310 169.730 ;
        RECT 62.120 169.680 62.380 170.830 ;
        RECT 62.555 169.755 62.810 170.660 ;
        RECT 62.980 170.070 63.310 170.830 ;
        RECT 63.525 169.900 63.695 170.660 ;
        RECT 61.055 169.190 61.310 169.520 ;
        RECT 60.715 168.450 60.970 169.025 ;
        RECT 61.140 169.000 61.310 169.190 ;
        RECT 61.590 169.180 61.945 169.550 ;
        RECT 61.140 168.830 61.855 169.000 ;
        RECT 61.140 168.280 61.470 168.660 ;
        RECT 61.685 168.450 61.855 168.830 ;
        RECT 62.120 168.280 62.380 169.120 ;
        RECT 62.555 169.025 62.725 169.755 ;
        RECT 62.980 169.730 63.695 169.900 ;
        RECT 62.980 169.520 63.150 169.730 ;
        RECT 63.955 169.665 64.245 170.830 ;
        RECT 65.340 170.395 70.685 170.830 ;
        RECT 62.895 169.190 63.150 169.520 ;
        RECT 62.555 168.450 62.810 169.025 ;
        RECT 62.980 169.000 63.150 169.190 ;
        RECT 63.430 169.180 63.785 169.550 ;
        RECT 66.930 169.145 67.280 170.395 ;
        RECT 71.230 169.850 71.485 170.520 ;
        RECT 71.665 170.030 71.950 170.830 ;
        RECT 72.130 170.110 72.460 170.620 ;
        RECT 71.230 169.810 71.410 169.850 ;
        RECT 62.980 168.830 63.695 169.000 ;
        RECT 62.980 168.280 63.310 168.660 ;
        RECT 63.525 168.450 63.695 168.830 ;
        RECT 63.955 168.280 64.245 169.005 ;
        RECT 68.760 168.825 69.100 169.655 ;
        RECT 71.145 169.640 71.410 169.810 ;
        RECT 71.230 168.990 71.410 169.640 ;
        RECT 72.130 169.520 72.380 170.110 ;
        RECT 72.730 169.960 72.900 170.570 ;
        RECT 73.070 170.140 73.400 170.830 ;
        RECT 73.630 170.280 73.870 170.570 ;
        RECT 74.070 170.450 74.490 170.830 ;
        RECT 74.670 170.360 75.300 170.610 ;
        RECT 75.770 170.450 76.100 170.830 ;
        RECT 74.670 170.280 74.840 170.360 ;
        RECT 76.270 170.280 76.440 170.570 ;
        RECT 76.620 170.450 77.000 170.830 ;
        RECT 77.240 170.445 78.070 170.615 ;
        RECT 73.630 170.110 74.840 170.280 ;
        RECT 71.580 169.190 72.380 169.520 ;
        RECT 65.340 168.280 70.685 168.825 ;
        RECT 71.230 168.460 71.485 168.990 ;
        RECT 71.665 168.280 71.950 168.740 ;
        RECT 72.130 168.540 72.380 169.190 ;
        RECT 72.580 169.940 72.900 169.960 ;
        RECT 72.580 169.770 74.500 169.940 ;
        RECT 72.580 168.875 72.770 169.770 ;
        RECT 74.670 169.600 74.840 170.110 ;
        RECT 75.010 169.850 75.530 170.160 ;
        RECT 72.940 169.430 74.840 169.600 ;
        RECT 72.940 169.370 73.270 169.430 ;
        RECT 73.420 169.200 73.750 169.260 ;
        RECT 73.090 168.930 73.750 169.200 ;
        RECT 72.580 168.545 72.900 168.875 ;
        RECT 73.080 168.280 73.740 168.760 ;
        RECT 73.940 168.670 74.110 169.430 ;
        RECT 75.010 169.260 75.190 169.670 ;
        RECT 74.280 169.090 74.610 169.210 ;
        RECT 75.360 169.090 75.530 169.850 ;
        RECT 74.280 168.920 75.530 169.090 ;
        RECT 75.700 170.030 77.070 170.280 ;
        RECT 75.700 169.260 75.890 170.030 ;
        RECT 76.820 169.770 77.070 170.030 ;
        RECT 76.060 169.600 76.310 169.760 ;
        RECT 77.240 169.600 77.410 170.445 ;
        RECT 78.305 170.160 78.475 170.660 ;
        RECT 78.645 170.330 78.975 170.830 ;
        RECT 77.580 169.770 78.080 170.150 ;
        RECT 78.305 169.990 79.000 170.160 ;
        RECT 76.060 169.430 77.410 169.600 ;
        RECT 76.990 169.390 77.410 169.430 ;
        RECT 75.700 168.920 76.120 169.260 ;
        RECT 76.410 168.930 76.820 169.260 ;
        RECT 73.940 168.500 74.790 168.670 ;
        RECT 75.350 168.280 75.670 168.740 ;
        RECT 75.870 168.490 76.120 168.920 ;
        RECT 76.410 168.280 76.820 168.720 ;
        RECT 76.990 168.660 77.160 169.390 ;
        RECT 77.330 168.840 77.680 169.210 ;
        RECT 77.860 168.900 78.080 169.770 ;
        RECT 78.250 169.200 78.660 169.820 ;
        RECT 78.830 169.020 79.000 169.990 ;
        RECT 78.305 168.830 79.000 169.020 ;
        RECT 76.990 168.460 78.005 168.660 ;
        RECT 78.305 168.500 78.475 168.830 ;
        RECT 78.645 168.280 78.975 168.660 ;
        RECT 79.190 168.540 79.415 170.660 ;
        RECT 79.585 170.330 79.915 170.830 ;
        RECT 80.085 170.160 80.255 170.660 ;
        RECT 79.590 169.990 80.255 170.160 ;
        RECT 79.590 169.000 79.820 169.990 ;
        RECT 79.990 169.170 80.340 169.820 ;
        RECT 80.515 169.740 83.105 170.830 ;
        RECT 83.275 170.070 83.790 170.480 ;
        RECT 84.025 170.070 84.195 170.830 ;
        RECT 84.365 170.490 86.395 170.660 ;
        RECT 80.515 169.220 81.725 169.740 ;
        RECT 81.895 169.050 83.105 169.570 ;
        RECT 83.275 169.260 83.615 170.070 ;
        RECT 84.365 169.825 84.535 170.490 ;
        RECT 84.930 170.150 86.055 170.320 ;
        RECT 83.785 169.635 84.535 169.825 ;
        RECT 84.705 169.810 85.715 169.980 ;
        RECT 83.275 169.090 84.505 169.260 ;
        RECT 79.590 168.830 80.255 169.000 ;
        RECT 79.585 168.280 79.915 168.660 ;
        RECT 80.085 168.540 80.255 168.830 ;
        RECT 80.515 168.280 83.105 169.050 ;
        RECT 83.550 168.485 83.795 169.090 ;
        RECT 84.015 168.280 84.525 168.815 ;
        RECT 84.705 168.450 84.895 169.810 ;
        RECT 85.065 169.470 85.340 169.610 ;
        RECT 85.065 169.300 85.345 169.470 ;
        RECT 85.065 168.450 85.340 169.300 ;
        RECT 85.545 169.010 85.715 169.810 ;
        RECT 85.885 169.020 86.055 170.150 ;
        RECT 86.225 169.520 86.395 170.490 ;
        RECT 86.565 169.690 86.735 170.830 ;
        RECT 86.905 169.690 87.240 170.660 ;
        RECT 86.225 169.190 86.420 169.520 ;
        RECT 86.645 169.190 86.900 169.520 ;
        RECT 86.645 169.020 86.815 169.190 ;
        RECT 87.070 169.020 87.240 169.690 ;
        RECT 85.885 168.850 86.815 169.020 ;
        RECT 85.885 168.815 86.060 168.850 ;
        RECT 85.530 168.450 86.060 168.815 ;
        RECT 86.485 168.280 86.815 168.680 ;
        RECT 86.985 168.450 87.240 169.020 ;
        RECT 87.875 169.755 88.145 170.660 ;
        RECT 88.315 170.070 88.645 170.830 ;
        RECT 88.825 169.900 88.995 170.660 ;
        RECT 87.875 168.955 88.045 169.755 ;
        RECT 88.330 169.730 88.995 169.900 ;
        RECT 88.330 169.585 88.500 169.730 ;
        RECT 89.715 169.665 90.005 170.830 ;
        RECT 90.175 169.740 92.765 170.830 ;
        RECT 88.215 169.255 88.500 169.585 ;
        RECT 88.330 169.000 88.500 169.255 ;
        RECT 88.735 169.180 89.065 169.550 ;
        RECT 90.175 169.220 91.385 169.740 ;
        RECT 92.975 169.690 93.205 170.830 ;
        RECT 93.375 169.680 93.705 170.660 ;
        RECT 93.875 169.690 94.085 170.830 ;
        RECT 94.430 170.200 94.715 170.660 ;
        RECT 94.885 170.370 95.155 170.830 ;
        RECT 94.430 169.980 95.385 170.200 ;
        RECT 91.555 169.050 92.765 169.570 ;
        RECT 92.955 169.270 93.285 169.520 ;
        RECT 87.875 168.450 88.135 168.955 ;
        RECT 88.330 168.830 88.995 169.000 ;
        RECT 88.315 168.280 88.645 168.660 ;
        RECT 88.825 168.450 88.995 168.830 ;
        RECT 89.715 168.280 90.005 169.005 ;
        RECT 90.175 168.280 92.765 169.050 ;
        RECT 92.975 168.280 93.205 169.100 ;
        RECT 93.455 169.080 93.705 169.680 ;
        RECT 94.315 169.250 95.005 169.810 ;
        RECT 93.375 168.450 93.705 169.080 ;
        RECT 93.875 168.280 94.085 169.100 ;
        RECT 95.175 169.080 95.385 169.980 ;
        RECT 94.430 168.910 95.385 169.080 ;
        RECT 95.555 169.810 95.955 170.660 ;
        RECT 96.145 170.200 96.425 170.660 ;
        RECT 96.945 170.370 97.270 170.830 ;
        RECT 96.145 169.980 97.270 170.200 ;
        RECT 95.555 169.250 96.650 169.810 ;
        RECT 96.820 169.520 97.270 169.980 ;
        RECT 97.440 169.690 97.825 170.660 ;
        RECT 98.005 170.020 98.300 170.830 ;
        RECT 94.430 168.450 94.715 168.910 ;
        RECT 94.885 168.280 95.155 168.740 ;
        RECT 95.555 168.450 95.955 169.250 ;
        RECT 96.820 169.190 97.375 169.520 ;
        RECT 96.820 169.080 97.270 169.190 ;
        RECT 96.145 168.910 97.270 169.080 ;
        RECT 97.545 169.020 97.825 169.690 ;
        RECT 98.480 169.520 98.725 170.660 ;
        RECT 98.900 170.020 99.160 170.830 ;
        RECT 99.760 170.825 106.035 170.830 ;
        RECT 99.340 169.520 99.590 170.655 ;
        RECT 99.760 170.030 100.020 170.825 ;
        RECT 100.190 169.930 100.450 170.655 ;
        RECT 100.620 170.100 100.880 170.825 ;
        RECT 101.050 169.930 101.310 170.655 ;
        RECT 101.480 170.100 101.740 170.825 ;
        RECT 101.910 169.930 102.170 170.655 ;
        RECT 102.340 170.100 102.600 170.825 ;
        RECT 102.770 169.930 103.030 170.655 ;
        RECT 103.200 170.100 103.445 170.825 ;
        RECT 103.615 169.930 103.875 170.655 ;
        RECT 104.060 170.100 104.305 170.825 ;
        RECT 104.475 169.930 104.735 170.655 ;
        RECT 104.920 170.100 105.165 170.825 ;
        RECT 105.335 169.930 105.595 170.655 ;
        RECT 105.780 170.100 106.035 170.825 ;
        RECT 100.190 169.915 105.595 169.930 ;
        RECT 106.205 169.915 106.495 170.655 ;
        RECT 106.665 170.085 106.935 170.830 ;
        RECT 100.190 169.690 106.935 169.915 ;
        RECT 96.145 168.450 96.425 168.910 ;
        RECT 96.945 168.280 97.270 168.740 ;
        RECT 97.440 168.450 97.825 169.020 ;
        RECT 97.995 168.960 98.310 169.520 ;
        RECT 98.480 169.270 105.600 169.520 ;
        RECT 97.995 168.280 98.300 168.790 ;
        RECT 98.480 168.460 98.730 169.270 ;
        RECT 98.900 168.280 99.160 168.805 ;
        RECT 99.340 168.460 99.590 169.270 ;
        RECT 105.770 169.100 106.935 169.690 ;
        RECT 107.325 169.660 107.655 170.830 ;
        RECT 107.855 169.490 108.185 170.660 ;
        RECT 108.385 169.660 108.715 170.830 ;
        RECT 108.915 169.490 109.275 170.660 ;
        RECT 109.445 169.690 109.775 170.830 ;
        RECT 109.960 170.405 110.295 170.830 ;
        RECT 110.465 170.225 110.650 170.630 ;
        RECT 109.985 170.050 110.650 170.225 ;
        RECT 110.855 170.050 111.185 170.830 ;
        RECT 107.855 169.210 109.275 169.490 ;
        RECT 100.190 168.930 106.935 169.100 ;
        RECT 99.760 168.280 100.020 168.840 ;
        RECT 100.190 168.475 100.450 168.930 ;
        RECT 100.620 168.280 100.880 168.760 ;
        RECT 101.050 168.475 101.310 168.930 ;
        RECT 101.480 168.280 101.740 168.760 ;
        RECT 101.910 168.475 102.170 168.930 ;
        RECT 102.340 168.280 102.585 168.760 ;
        RECT 102.755 168.475 103.030 168.930 ;
        RECT 103.200 168.280 103.445 168.760 ;
        RECT 103.615 168.475 103.875 168.930 ;
        RECT 104.055 168.280 104.305 168.760 ;
        RECT 104.475 168.475 104.735 168.930 ;
        RECT 104.915 168.280 105.165 168.760 ;
        RECT 105.335 168.475 105.595 168.930 ;
        RECT 105.775 168.280 106.035 168.760 ;
        RECT 106.205 168.475 106.465 168.930 ;
        RECT 106.635 168.280 106.935 168.760 ;
        RECT 107.865 168.280 108.195 168.970 ;
        RECT 108.915 168.875 109.275 169.210 ;
        RECT 109.445 168.940 109.785 169.520 ;
        RECT 109.985 169.020 110.325 170.050 ;
        RECT 111.355 169.860 111.625 170.630 ;
        RECT 110.495 169.690 111.625 169.860 ;
        RECT 110.495 169.190 110.745 169.690 ;
        RECT 108.655 168.450 109.275 168.875 ;
        RECT 109.985 168.850 110.670 169.020 ;
        RECT 110.925 168.940 111.285 169.520 ;
        RECT 109.445 168.280 109.775 168.770 ;
        RECT 109.960 168.280 110.295 168.680 ;
        RECT 110.465 168.450 110.670 168.850 ;
        RECT 111.455 168.780 111.625 169.690 ;
        RECT 111.795 169.740 114.385 170.830 ;
        RECT 114.555 169.740 115.765 170.830 ;
        RECT 111.795 169.220 113.005 169.740 ;
        RECT 113.175 169.050 114.385 169.570 ;
        RECT 114.555 169.200 115.075 169.740 ;
        RECT 110.880 168.280 111.155 168.760 ;
        RECT 111.365 168.450 111.625 168.780 ;
        RECT 111.795 168.280 114.385 169.050 ;
        RECT 115.245 169.030 115.765 169.570 ;
        RECT 114.555 168.280 115.765 169.030 ;
        RECT 10.510 168.110 115.850 168.280 ;
        RECT 10.595 167.360 11.805 168.110 ;
        RECT 10.595 166.820 11.115 167.360 ;
        RECT 12.435 167.340 14.105 168.110 ;
        RECT 14.280 167.565 19.625 168.110 ;
        RECT 11.285 166.650 11.805 167.190 ;
        RECT 10.595 165.560 11.805 166.650 ;
        RECT 12.435 166.650 13.185 167.170 ;
        RECT 13.355 166.820 14.105 167.340 ;
        RECT 12.435 165.560 14.105 166.650 ;
        RECT 15.870 165.995 16.220 167.245 ;
        RECT 17.700 166.735 18.040 167.565 ;
        RECT 19.855 167.290 20.065 168.110 ;
        RECT 20.235 167.310 20.565 167.940 ;
        RECT 20.235 166.710 20.485 167.310 ;
        RECT 20.735 167.290 20.965 168.110 ;
        RECT 21.265 167.560 21.435 167.940 ;
        RECT 21.615 167.730 21.945 168.110 ;
        RECT 21.265 167.390 21.930 167.560 ;
        RECT 22.125 167.435 22.385 167.940 ;
        RECT 20.655 166.870 20.985 167.120 ;
        RECT 21.195 166.840 21.525 167.210 ;
        RECT 21.760 167.135 21.930 167.390 ;
        RECT 21.760 166.805 22.045 167.135 ;
        RECT 14.280 165.560 19.625 165.995 ;
        RECT 19.855 165.560 20.065 166.700 ;
        RECT 20.235 165.730 20.565 166.710 ;
        RECT 20.735 165.560 20.965 166.700 ;
        RECT 21.760 166.660 21.930 166.805 ;
        RECT 21.265 166.490 21.930 166.660 ;
        RECT 22.215 166.635 22.385 167.435 ;
        RECT 22.595 167.290 22.825 168.110 ;
        RECT 22.995 167.310 23.325 167.940 ;
        RECT 22.575 166.870 22.905 167.120 ;
        RECT 23.075 166.710 23.325 167.310 ;
        RECT 23.495 167.290 23.705 168.110 ;
        RECT 24.025 167.560 24.195 167.940 ;
        RECT 24.375 167.730 24.705 168.110 ;
        RECT 24.025 167.390 24.690 167.560 ;
        RECT 24.885 167.435 25.145 167.940 ;
        RECT 23.955 166.840 24.285 167.210 ;
        RECT 24.520 167.135 24.690 167.390 ;
        RECT 21.265 165.730 21.435 166.490 ;
        RECT 21.615 165.560 21.945 166.320 ;
        RECT 22.115 165.730 22.385 166.635 ;
        RECT 22.595 165.560 22.825 166.700 ;
        RECT 22.995 165.730 23.325 166.710 ;
        RECT 24.520 166.805 24.805 167.135 ;
        RECT 23.495 165.560 23.705 166.700 ;
        RECT 24.520 166.660 24.690 166.805 ;
        RECT 24.025 166.490 24.690 166.660 ;
        RECT 24.975 166.635 25.145 167.435 ;
        RECT 25.315 167.385 25.605 168.110 ;
        RECT 26.810 167.480 27.095 167.940 ;
        RECT 27.265 167.650 27.535 168.110 ;
        RECT 26.810 167.310 27.765 167.480 ;
        RECT 24.025 165.730 24.195 166.490 ;
        RECT 24.375 165.560 24.705 166.320 ;
        RECT 24.875 165.730 25.145 166.635 ;
        RECT 25.315 165.560 25.605 166.725 ;
        RECT 26.695 166.580 27.385 167.140 ;
        RECT 27.555 166.410 27.765 167.310 ;
        RECT 26.810 166.190 27.765 166.410 ;
        RECT 27.935 167.140 28.335 167.940 ;
        RECT 28.525 167.480 28.805 167.940 ;
        RECT 29.325 167.650 29.650 168.110 ;
        RECT 28.525 167.310 29.650 167.480 ;
        RECT 29.820 167.370 30.205 167.940 ;
        RECT 29.200 167.200 29.650 167.310 ;
        RECT 27.935 166.580 29.030 167.140 ;
        RECT 29.200 166.870 29.755 167.200 ;
        RECT 26.810 165.730 27.095 166.190 ;
        RECT 27.265 165.560 27.535 166.020 ;
        RECT 27.935 165.730 28.335 166.580 ;
        RECT 29.200 166.410 29.650 166.870 ;
        RECT 29.925 166.700 30.205 167.370 ;
        RECT 30.490 167.480 30.775 167.940 ;
        RECT 30.945 167.650 31.215 168.110 ;
        RECT 30.490 167.310 31.445 167.480 ;
        RECT 28.525 166.190 29.650 166.410 ;
        RECT 28.525 165.730 28.805 166.190 ;
        RECT 29.325 165.560 29.650 166.020 ;
        RECT 29.820 165.730 30.205 166.700 ;
        RECT 30.375 166.580 31.065 167.140 ;
        RECT 31.235 166.410 31.445 167.310 ;
        RECT 30.490 166.190 31.445 166.410 ;
        RECT 31.615 167.140 32.015 167.940 ;
        RECT 32.205 167.480 32.485 167.940 ;
        RECT 33.005 167.650 33.330 168.110 ;
        RECT 32.205 167.310 33.330 167.480 ;
        RECT 33.500 167.370 33.885 167.940 ;
        RECT 32.880 167.200 33.330 167.310 ;
        RECT 31.615 166.580 32.710 167.140 ;
        RECT 32.880 166.870 33.435 167.200 ;
        RECT 30.490 165.730 30.775 166.190 ;
        RECT 30.945 165.560 31.215 166.020 ;
        RECT 31.615 165.730 32.015 166.580 ;
        RECT 32.880 166.410 33.330 166.870 ;
        RECT 33.605 166.700 33.885 167.370 ;
        RECT 34.170 167.480 34.455 167.940 ;
        RECT 34.625 167.650 34.895 168.110 ;
        RECT 34.170 167.310 35.125 167.480 ;
        RECT 32.205 166.190 33.330 166.410 ;
        RECT 32.205 165.730 32.485 166.190 ;
        RECT 33.005 165.560 33.330 166.020 ;
        RECT 33.500 165.730 33.885 166.700 ;
        RECT 34.055 166.580 34.745 167.140 ;
        RECT 34.915 166.410 35.125 167.310 ;
        RECT 34.170 166.190 35.125 166.410 ;
        RECT 35.295 167.140 35.695 167.940 ;
        RECT 35.885 167.480 36.165 167.940 ;
        RECT 36.685 167.650 37.010 168.110 ;
        RECT 35.885 167.310 37.010 167.480 ;
        RECT 37.180 167.370 37.565 167.940 ;
        RECT 36.560 167.200 37.010 167.310 ;
        RECT 35.295 166.580 36.390 167.140 ;
        RECT 36.560 166.870 37.115 167.200 ;
        RECT 34.170 165.730 34.455 166.190 ;
        RECT 34.625 165.560 34.895 166.020 ;
        RECT 35.295 165.730 35.695 166.580 ;
        RECT 36.560 166.410 37.010 166.870 ;
        RECT 37.285 166.700 37.565 167.370 ;
        RECT 35.885 166.190 37.010 166.410 ;
        RECT 35.885 165.730 36.165 166.190 ;
        RECT 36.685 165.560 37.010 166.020 ;
        RECT 37.180 165.730 37.565 166.700 ;
        RECT 37.740 167.400 37.995 167.930 ;
        RECT 38.165 167.650 38.470 168.110 ;
        RECT 38.715 167.730 39.785 167.900 ;
        RECT 37.740 166.750 37.950 167.400 ;
        RECT 38.715 167.375 39.035 167.730 ;
        RECT 38.710 167.200 39.035 167.375 ;
        RECT 38.120 166.900 39.035 167.200 ;
        RECT 39.205 167.160 39.445 167.560 ;
        RECT 39.615 167.500 39.785 167.730 ;
        RECT 39.955 167.670 40.145 168.110 ;
        RECT 40.315 167.660 41.265 167.940 ;
        RECT 41.485 167.750 41.835 167.920 ;
        RECT 39.615 167.330 40.145 167.500 ;
        RECT 38.120 166.870 38.860 166.900 ;
        RECT 37.740 165.870 37.995 166.750 ;
        RECT 38.165 165.560 38.470 166.700 ;
        RECT 38.690 166.280 38.860 166.870 ;
        RECT 39.205 166.790 39.745 167.160 ;
        RECT 39.925 167.050 40.145 167.330 ;
        RECT 40.315 166.880 40.485 167.660 ;
        RECT 40.080 166.710 40.485 166.880 ;
        RECT 40.655 166.870 41.005 167.490 ;
        RECT 40.080 166.620 40.250 166.710 ;
        RECT 41.175 166.700 41.385 167.490 ;
        RECT 39.030 166.450 40.250 166.620 ;
        RECT 40.710 166.540 41.385 166.700 ;
        RECT 38.690 166.110 39.490 166.280 ;
        RECT 38.810 165.560 39.140 165.940 ;
        RECT 39.320 165.820 39.490 166.110 ;
        RECT 40.080 166.070 40.250 166.450 ;
        RECT 40.420 166.530 41.385 166.540 ;
        RECT 41.575 167.360 41.835 167.750 ;
        RECT 42.045 167.650 42.375 168.110 ;
        RECT 43.250 167.720 44.105 167.890 ;
        RECT 44.310 167.720 44.805 167.890 ;
        RECT 44.975 167.750 45.305 168.110 ;
        RECT 41.575 166.670 41.745 167.360 ;
        RECT 41.915 167.010 42.085 167.190 ;
        RECT 42.255 167.180 43.045 167.430 ;
        RECT 43.250 167.010 43.420 167.720 ;
        RECT 43.590 167.210 43.945 167.430 ;
        RECT 41.915 166.840 43.605 167.010 ;
        RECT 40.420 166.240 40.880 166.530 ;
        RECT 41.575 166.500 43.075 166.670 ;
        RECT 41.575 166.360 41.745 166.500 ;
        RECT 41.185 166.190 41.745 166.360 ;
        RECT 39.660 165.560 39.910 166.020 ;
        RECT 40.080 165.730 40.950 166.070 ;
        RECT 41.185 165.730 41.355 166.190 ;
        RECT 42.190 166.160 43.265 166.330 ;
        RECT 41.525 165.560 41.895 166.020 ;
        RECT 42.190 165.820 42.360 166.160 ;
        RECT 42.530 165.560 42.860 165.990 ;
        RECT 43.095 165.820 43.265 166.160 ;
        RECT 43.435 166.060 43.605 166.840 ;
        RECT 43.775 166.620 43.945 167.210 ;
        RECT 44.115 166.810 44.465 167.430 ;
        RECT 43.775 166.230 44.240 166.620 ;
        RECT 44.635 166.360 44.805 167.720 ;
        RECT 44.975 166.530 45.435 167.580 ;
        RECT 44.410 166.190 44.805 166.360 ;
        RECT 44.410 166.060 44.580 166.190 ;
        RECT 43.435 165.730 44.115 166.060 ;
        RECT 44.330 165.730 44.580 166.060 ;
        RECT 44.750 165.560 45.000 166.020 ;
        RECT 45.170 165.745 45.495 166.530 ;
        RECT 45.665 165.730 45.835 167.850 ;
        RECT 46.005 167.730 46.335 168.110 ;
        RECT 46.505 167.560 46.760 167.850 ;
        RECT 46.010 167.390 46.760 167.560 ;
        RECT 46.010 166.400 46.240 167.390 ;
        RECT 46.935 167.340 49.525 168.110 ;
        RECT 46.410 166.570 46.760 167.220 ;
        RECT 46.935 166.650 48.145 167.170 ;
        RECT 48.315 166.820 49.525 167.340 ;
        RECT 49.735 167.290 49.965 168.110 ;
        RECT 50.135 167.310 50.465 167.940 ;
        RECT 49.715 166.870 50.045 167.120 ;
        RECT 50.215 166.710 50.465 167.310 ;
        RECT 50.635 167.290 50.845 168.110 ;
        RECT 51.075 167.385 51.365 168.110 ;
        RECT 51.535 167.340 53.205 168.110 ;
        RECT 46.010 166.230 46.760 166.400 ;
        RECT 46.005 165.560 46.335 166.060 ;
        RECT 46.505 165.730 46.760 166.230 ;
        RECT 46.935 165.560 49.525 166.650 ;
        RECT 49.735 165.560 49.965 166.700 ;
        RECT 50.135 165.730 50.465 166.710 ;
        RECT 50.635 165.560 50.845 166.700 ;
        RECT 51.075 165.560 51.365 166.725 ;
        RECT 51.535 166.650 52.285 167.170 ;
        RECT 52.455 166.820 53.205 167.340 ;
        RECT 53.525 167.310 53.855 168.110 ;
        RECT 54.025 167.460 54.195 167.940 ;
        RECT 54.365 167.630 54.695 168.110 ;
        RECT 54.865 167.460 55.035 167.940 ;
        RECT 55.285 167.630 55.525 168.110 ;
        RECT 55.705 167.460 55.875 167.940 ;
        RECT 54.025 167.290 55.035 167.460 ;
        RECT 55.240 167.290 55.875 167.460 ;
        RECT 57.055 167.340 60.565 168.110 ;
        RECT 54.025 167.090 54.520 167.290 ;
        RECT 55.240 167.120 55.410 167.290 ;
        RECT 54.025 166.920 54.525 167.090 ;
        RECT 54.910 166.950 55.410 167.120 ;
        RECT 54.025 166.750 54.520 166.920 ;
        RECT 51.535 165.560 53.205 166.650 ;
        RECT 53.525 165.560 53.855 166.710 ;
        RECT 54.025 166.580 55.035 166.750 ;
        RECT 54.025 165.730 54.195 166.580 ;
        RECT 54.365 165.560 54.695 166.360 ;
        RECT 54.865 165.730 55.035 166.580 ;
        RECT 55.240 166.710 55.410 166.950 ;
        RECT 55.580 166.880 55.960 167.120 ;
        RECT 55.240 166.540 55.955 166.710 ;
        RECT 55.215 165.560 55.455 166.360 ;
        RECT 55.625 165.730 55.955 166.540 ;
        RECT 57.055 166.650 58.745 167.170 ;
        RECT 58.915 166.820 60.565 167.340 ;
        RECT 60.735 167.610 61.035 167.940 ;
        RECT 61.205 167.630 61.480 168.110 ;
        RECT 60.735 166.700 60.905 167.610 ;
        RECT 61.660 167.460 61.955 167.850 ;
        RECT 62.125 167.630 62.380 168.110 ;
        RECT 62.555 167.460 62.815 167.850 ;
        RECT 62.985 167.630 63.265 168.110 ;
        RECT 63.505 167.580 63.835 167.940 ;
        RECT 64.005 167.750 64.335 168.110 ;
        RECT 64.535 167.580 64.865 167.940 ;
        RECT 61.075 166.870 61.425 167.440 ;
        RECT 61.660 167.290 63.310 167.460 ;
        RECT 63.505 167.370 64.865 167.580 ;
        RECT 65.375 167.350 66.085 167.940 ;
        RECT 61.595 166.950 62.735 167.120 ;
        RECT 61.595 166.700 61.765 166.950 ;
        RECT 62.905 166.780 63.310 167.290 ;
        RECT 65.855 167.260 66.085 167.350 ;
        RECT 66.530 167.300 66.775 167.905 ;
        RECT 66.995 167.575 67.505 168.110 ;
        RECT 63.495 166.870 63.805 167.200 ;
        RECT 64.015 166.870 64.390 167.200 ;
        RECT 64.710 166.870 65.205 167.200 ;
        RECT 57.055 165.560 60.565 166.650 ;
        RECT 60.735 166.530 61.765 166.700 ;
        RECT 62.555 166.610 63.310 166.780 ;
        RECT 60.735 165.730 61.045 166.530 ;
        RECT 62.555 166.360 62.815 166.610 ;
        RECT 61.215 165.560 61.525 166.360 ;
        RECT 61.695 166.190 62.815 166.360 ;
        RECT 61.695 165.730 61.955 166.190 ;
        RECT 62.125 165.560 62.380 166.020 ;
        RECT 62.555 165.730 62.815 166.190 ;
        RECT 62.985 165.560 63.270 166.430 ;
        RECT 63.505 165.560 63.835 166.620 ;
        RECT 64.015 165.945 64.185 166.870 ;
        RECT 64.355 166.380 64.685 166.600 ;
        RECT 64.880 166.580 65.205 166.870 ;
        RECT 65.380 166.580 65.710 167.120 ;
        RECT 65.880 166.380 66.085 167.260 ;
        RECT 64.355 166.150 66.085 166.380 ;
        RECT 64.355 165.750 64.685 166.150 ;
        RECT 64.855 165.560 65.185 165.920 ;
        RECT 65.385 165.730 66.085 166.150 ;
        RECT 66.255 167.130 67.485 167.300 ;
        RECT 66.255 166.320 66.595 167.130 ;
        RECT 66.765 166.565 67.515 166.755 ;
        RECT 66.255 165.910 66.770 166.320 ;
        RECT 67.005 165.560 67.175 166.320 ;
        RECT 67.345 165.900 67.515 166.565 ;
        RECT 67.685 166.580 67.875 167.940 ;
        RECT 68.045 167.090 68.320 167.940 ;
        RECT 68.510 167.575 69.040 167.940 ;
        RECT 69.465 167.710 69.795 168.110 ;
        RECT 68.865 167.540 69.040 167.575 ;
        RECT 68.045 166.920 68.325 167.090 ;
        RECT 68.045 166.780 68.320 166.920 ;
        RECT 68.525 166.580 68.695 167.380 ;
        RECT 67.685 166.410 68.695 166.580 ;
        RECT 68.865 167.370 69.795 167.540 ;
        RECT 69.965 167.370 70.220 167.940 ;
        RECT 68.865 166.240 69.035 167.370 ;
        RECT 69.625 167.200 69.795 167.370 ;
        RECT 67.910 166.070 69.035 166.240 ;
        RECT 69.205 166.870 69.400 167.200 ;
        RECT 69.625 166.870 69.880 167.200 ;
        RECT 69.205 165.900 69.375 166.870 ;
        RECT 70.050 166.700 70.220 167.370 ;
        RECT 70.670 167.300 70.915 167.905 ;
        RECT 71.135 167.575 71.645 168.110 ;
        RECT 67.345 165.730 69.375 165.900 ;
        RECT 69.545 165.560 69.715 166.700 ;
        RECT 69.885 165.730 70.220 166.700 ;
        RECT 70.395 167.130 71.625 167.300 ;
        RECT 70.395 166.320 70.735 167.130 ;
        RECT 70.905 166.565 71.655 166.755 ;
        RECT 70.395 165.910 70.910 166.320 ;
        RECT 71.145 165.560 71.315 166.320 ;
        RECT 71.485 165.900 71.655 166.565 ;
        RECT 71.825 166.580 72.015 167.940 ;
        RECT 72.185 167.090 72.460 167.940 ;
        RECT 72.650 167.575 73.180 167.940 ;
        RECT 73.605 167.710 73.935 168.110 ;
        RECT 73.005 167.540 73.180 167.575 ;
        RECT 72.185 166.920 72.465 167.090 ;
        RECT 72.185 166.780 72.460 166.920 ;
        RECT 72.665 166.580 72.835 167.380 ;
        RECT 71.825 166.410 72.835 166.580 ;
        RECT 73.005 167.370 73.935 167.540 ;
        RECT 74.105 167.370 74.360 167.940 ;
        RECT 73.005 166.240 73.175 167.370 ;
        RECT 73.765 167.200 73.935 167.370 ;
        RECT 72.050 166.070 73.175 166.240 ;
        RECT 73.345 166.870 73.540 167.200 ;
        RECT 73.765 166.870 74.020 167.200 ;
        RECT 73.345 165.900 73.515 166.870 ;
        RECT 74.190 166.700 74.360 167.370 ;
        RECT 75.055 167.290 75.265 168.110 ;
        RECT 75.435 167.310 75.765 167.940 ;
        RECT 75.435 166.710 75.685 167.310 ;
        RECT 75.935 167.290 76.165 168.110 ;
        RECT 76.835 167.385 77.125 168.110 ;
        RECT 77.385 167.560 77.555 167.940 ;
        RECT 77.735 167.730 78.065 168.110 ;
        RECT 77.385 167.390 78.050 167.560 ;
        RECT 78.245 167.435 78.505 167.940 ;
        RECT 75.855 166.870 76.185 167.120 ;
        RECT 77.315 166.840 77.645 167.210 ;
        RECT 77.880 167.135 78.050 167.390 ;
        RECT 77.880 166.805 78.165 167.135 ;
        RECT 71.485 165.730 73.515 165.900 ;
        RECT 73.685 165.560 73.855 166.700 ;
        RECT 74.025 165.730 74.360 166.700 ;
        RECT 75.055 165.560 75.265 166.700 ;
        RECT 75.435 165.730 75.765 166.710 ;
        RECT 75.935 165.560 76.165 166.700 ;
        RECT 76.835 165.560 77.125 166.725 ;
        RECT 77.880 166.660 78.050 166.805 ;
        RECT 77.385 166.490 78.050 166.660 ;
        RECT 78.335 166.635 78.505 167.435 ;
        RECT 79.135 167.340 81.725 168.110 ;
        RECT 81.900 167.565 87.245 168.110 ;
        RECT 77.385 165.730 77.555 166.490 ;
        RECT 77.735 165.560 78.065 166.320 ;
        RECT 78.235 165.730 78.505 166.635 ;
        RECT 79.135 166.650 80.345 167.170 ;
        RECT 80.515 166.820 81.725 167.340 ;
        RECT 79.135 165.560 81.725 166.650 ;
        RECT 83.490 165.995 83.840 167.245 ;
        RECT 85.320 166.735 85.660 167.565 ;
        RECT 87.455 167.290 87.685 168.110 ;
        RECT 87.855 167.310 88.185 167.940 ;
        RECT 87.435 166.870 87.765 167.120 ;
        RECT 87.935 166.710 88.185 167.310 ;
        RECT 88.355 167.290 88.565 168.110 ;
        RECT 88.910 167.480 89.195 167.940 ;
        RECT 89.365 167.650 89.635 168.110 ;
        RECT 88.910 167.310 89.865 167.480 ;
        RECT 81.900 165.560 87.245 165.995 ;
        RECT 87.455 165.560 87.685 166.700 ;
        RECT 87.855 165.730 88.185 166.710 ;
        RECT 88.355 165.560 88.565 166.700 ;
        RECT 88.795 166.580 89.485 167.140 ;
        RECT 89.655 166.410 89.865 167.310 ;
        RECT 88.910 166.190 89.865 166.410 ;
        RECT 90.035 167.140 90.435 167.940 ;
        RECT 90.625 167.480 90.905 167.940 ;
        RECT 91.425 167.650 91.750 168.110 ;
        RECT 90.625 167.310 91.750 167.480 ;
        RECT 91.920 167.370 92.305 167.940 ;
        RECT 91.300 167.200 91.750 167.310 ;
        RECT 90.035 166.580 91.130 167.140 ;
        RECT 91.300 166.870 91.855 167.200 ;
        RECT 88.910 165.730 89.195 166.190 ;
        RECT 89.365 165.560 89.635 166.020 ;
        RECT 90.035 165.730 90.435 166.580 ;
        RECT 91.300 166.410 91.750 166.870 ;
        RECT 92.025 166.700 92.305 167.370 ;
        RECT 90.625 166.190 91.750 166.410 ;
        RECT 90.625 165.730 90.905 166.190 ;
        RECT 91.425 165.560 91.750 166.020 ;
        RECT 91.920 165.730 92.305 166.700 ;
        RECT 92.480 167.400 92.735 167.930 ;
        RECT 92.905 167.650 93.210 168.110 ;
        RECT 93.455 167.730 94.525 167.900 ;
        RECT 92.480 166.750 92.690 167.400 ;
        RECT 93.455 167.375 93.775 167.730 ;
        RECT 93.450 167.200 93.775 167.375 ;
        RECT 92.860 166.900 93.775 167.200 ;
        RECT 93.945 167.160 94.185 167.560 ;
        RECT 94.355 167.500 94.525 167.730 ;
        RECT 94.695 167.670 94.885 168.110 ;
        RECT 95.055 167.660 96.005 167.940 ;
        RECT 96.225 167.750 96.575 167.920 ;
        RECT 94.355 167.330 94.885 167.500 ;
        RECT 92.860 166.870 93.600 166.900 ;
        RECT 92.480 165.870 92.735 166.750 ;
        RECT 92.905 165.560 93.210 166.700 ;
        RECT 93.430 166.280 93.600 166.870 ;
        RECT 93.945 166.790 94.485 167.160 ;
        RECT 94.665 167.050 94.885 167.330 ;
        RECT 95.055 166.880 95.225 167.660 ;
        RECT 94.820 166.710 95.225 166.880 ;
        RECT 95.395 166.870 95.745 167.490 ;
        RECT 94.820 166.620 94.990 166.710 ;
        RECT 95.915 166.700 96.125 167.490 ;
        RECT 93.770 166.450 94.990 166.620 ;
        RECT 95.450 166.540 96.125 166.700 ;
        RECT 93.430 166.110 94.230 166.280 ;
        RECT 93.550 165.560 93.880 165.940 ;
        RECT 94.060 165.820 94.230 166.110 ;
        RECT 94.820 166.070 94.990 166.450 ;
        RECT 95.160 166.530 96.125 166.540 ;
        RECT 96.315 167.360 96.575 167.750 ;
        RECT 96.785 167.650 97.115 168.110 ;
        RECT 97.990 167.720 98.845 167.890 ;
        RECT 99.050 167.720 99.545 167.890 ;
        RECT 99.715 167.750 100.045 168.110 ;
        RECT 96.315 166.670 96.485 167.360 ;
        RECT 96.655 167.010 96.825 167.190 ;
        RECT 96.995 167.180 97.785 167.430 ;
        RECT 97.990 167.010 98.160 167.720 ;
        RECT 98.330 167.210 98.685 167.430 ;
        RECT 96.655 166.840 98.345 167.010 ;
        RECT 95.160 166.240 95.620 166.530 ;
        RECT 96.315 166.500 97.815 166.670 ;
        RECT 96.315 166.360 96.485 166.500 ;
        RECT 95.925 166.190 96.485 166.360 ;
        RECT 94.400 165.560 94.650 166.020 ;
        RECT 94.820 165.730 95.690 166.070 ;
        RECT 95.925 165.730 96.095 166.190 ;
        RECT 96.930 166.160 98.005 166.330 ;
        RECT 96.265 165.560 96.635 166.020 ;
        RECT 96.930 165.820 97.100 166.160 ;
        RECT 97.270 165.560 97.600 165.990 ;
        RECT 97.835 165.820 98.005 166.160 ;
        RECT 98.175 166.060 98.345 166.840 ;
        RECT 98.515 166.620 98.685 167.210 ;
        RECT 98.855 166.810 99.205 167.430 ;
        RECT 98.515 166.230 98.980 166.620 ;
        RECT 99.375 166.360 99.545 167.720 ;
        RECT 99.715 166.530 100.175 167.580 ;
        RECT 99.150 166.190 99.545 166.360 ;
        RECT 99.150 166.060 99.320 166.190 ;
        RECT 98.175 165.730 98.855 166.060 ;
        RECT 99.070 165.730 99.320 166.060 ;
        RECT 99.490 165.560 99.740 166.020 ;
        RECT 99.910 165.745 100.235 166.530 ;
        RECT 100.405 165.730 100.575 167.850 ;
        RECT 100.745 167.730 101.075 168.110 ;
        RECT 101.245 167.560 101.500 167.850 ;
        RECT 100.750 167.390 101.500 167.560 ;
        RECT 100.750 166.400 100.980 167.390 ;
        RECT 102.595 167.385 102.885 168.110 ;
        RECT 103.555 167.290 103.785 168.110 ;
        RECT 103.955 167.310 104.285 167.940 ;
        RECT 101.150 166.570 101.500 167.220 ;
        RECT 103.535 166.870 103.865 167.120 ;
        RECT 100.750 166.230 101.500 166.400 ;
        RECT 100.745 165.560 101.075 166.060 ;
        RECT 101.245 165.730 101.500 166.230 ;
        RECT 102.595 165.560 102.885 166.725 ;
        RECT 104.035 166.710 104.285 167.310 ;
        RECT 104.455 167.290 104.665 168.110 ;
        RECT 104.900 167.400 105.155 167.930 ;
        RECT 105.325 167.650 105.630 168.110 ;
        RECT 105.875 167.730 106.945 167.900 ;
        RECT 103.555 165.560 103.785 166.700 ;
        RECT 103.955 165.730 104.285 166.710 ;
        RECT 104.900 166.750 105.110 167.400 ;
        RECT 105.875 167.375 106.195 167.730 ;
        RECT 105.870 167.200 106.195 167.375 ;
        RECT 105.280 166.900 106.195 167.200 ;
        RECT 106.365 167.160 106.605 167.560 ;
        RECT 106.775 167.500 106.945 167.730 ;
        RECT 107.115 167.670 107.305 168.110 ;
        RECT 107.475 167.660 108.425 167.940 ;
        RECT 108.645 167.750 108.995 167.920 ;
        RECT 106.775 167.330 107.305 167.500 ;
        RECT 105.280 166.870 106.020 166.900 ;
        RECT 104.455 165.560 104.665 166.700 ;
        RECT 104.900 165.870 105.155 166.750 ;
        RECT 105.325 165.560 105.630 166.700 ;
        RECT 105.850 166.280 106.020 166.870 ;
        RECT 106.365 166.790 106.905 167.160 ;
        RECT 107.085 167.050 107.305 167.330 ;
        RECT 107.475 166.880 107.645 167.660 ;
        RECT 107.240 166.710 107.645 166.880 ;
        RECT 107.815 166.870 108.165 167.490 ;
        RECT 107.240 166.620 107.410 166.710 ;
        RECT 108.335 166.700 108.545 167.490 ;
        RECT 106.190 166.450 107.410 166.620 ;
        RECT 107.870 166.540 108.545 166.700 ;
        RECT 105.850 166.110 106.650 166.280 ;
        RECT 105.970 165.560 106.300 165.940 ;
        RECT 106.480 165.820 106.650 166.110 ;
        RECT 107.240 166.070 107.410 166.450 ;
        RECT 107.580 166.530 108.545 166.540 ;
        RECT 108.735 167.360 108.995 167.750 ;
        RECT 109.205 167.650 109.535 168.110 ;
        RECT 110.410 167.720 111.265 167.890 ;
        RECT 111.470 167.720 111.965 167.890 ;
        RECT 112.135 167.750 112.465 168.110 ;
        RECT 108.735 166.670 108.905 167.360 ;
        RECT 109.075 167.010 109.245 167.190 ;
        RECT 109.415 167.180 110.205 167.430 ;
        RECT 110.410 167.010 110.580 167.720 ;
        RECT 110.750 167.210 111.105 167.430 ;
        RECT 109.075 166.840 110.765 167.010 ;
        RECT 107.580 166.240 108.040 166.530 ;
        RECT 108.735 166.500 110.235 166.670 ;
        RECT 108.735 166.360 108.905 166.500 ;
        RECT 108.345 166.190 108.905 166.360 ;
        RECT 106.820 165.560 107.070 166.020 ;
        RECT 107.240 165.730 108.110 166.070 ;
        RECT 108.345 165.730 108.515 166.190 ;
        RECT 109.350 166.160 110.425 166.330 ;
        RECT 108.685 165.560 109.055 166.020 ;
        RECT 109.350 165.820 109.520 166.160 ;
        RECT 109.690 165.560 110.020 165.990 ;
        RECT 110.255 165.820 110.425 166.160 ;
        RECT 110.595 166.060 110.765 166.840 ;
        RECT 110.935 166.620 111.105 167.210 ;
        RECT 111.275 166.810 111.625 167.430 ;
        RECT 110.935 166.230 111.400 166.620 ;
        RECT 111.795 166.360 111.965 167.720 ;
        RECT 112.135 166.530 112.595 167.580 ;
        RECT 111.570 166.190 111.965 166.360 ;
        RECT 111.570 166.060 111.740 166.190 ;
        RECT 110.595 165.730 111.275 166.060 ;
        RECT 111.490 165.730 111.740 166.060 ;
        RECT 111.910 165.560 112.160 166.020 ;
        RECT 112.330 165.745 112.655 166.530 ;
        RECT 112.825 165.730 112.995 167.850 ;
        RECT 113.165 167.730 113.495 168.110 ;
        RECT 113.665 167.560 113.920 167.850 ;
        RECT 113.170 167.390 113.920 167.560 ;
        RECT 113.170 166.400 113.400 167.390 ;
        RECT 114.555 167.360 115.765 168.110 ;
        RECT 113.570 166.570 113.920 167.220 ;
        RECT 114.555 166.650 115.075 167.190 ;
        RECT 115.245 166.820 115.765 167.360 ;
        RECT 113.170 166.230 113.920 166.400 ;
        RECT 113.165 165.560 113.495 166.060 ;
        RECT 113.665 165.730 113.920 166.230 ;
        RECT 114.555 165.560 115.765 166.650 ;
        RECT 10.510 165.390 115.850 165.560 ;
        RECT 10.595 164.300 11.805 165.390 ;
        RECT 10.595 163.590 11.115 164.130 ;
        RECT 11.285 163.760 11.805 164.300 ;
        RECT 12.435 164.225 12.725 165.390 ;
        RECT 12.895 164.300 16.405 165.390 ;
        RECT 12.895 163.780 14.585 164.300 ;
        RECT 16.580 164.200 16.835 165.080 ;
        RECT 17.005 164.250 17.310 165.390 ;
        RECT 17.650 165.010 17.980 165.390 ;
        RECT 18.160 164.840 18.330 165.130 ;
        RECT 18.500 164.930 18.750 165.390 ;
        RECT 17.530 164.670 18.330 164.840 ;
        RECT 18.920 164.880 19.790 165.220 ;
        RECT 14.755 163.610 16.405 164.130 ;
        RECT 10.595 162.840 11.805 163.590 ;
        RECT 12.435 162.840 12.725 163.565 ;
        RECT 12.895 162.840 16.405 163.610 ;
        RECT 16.580 163.550 16.790 164.200 ;
        RECT 17.530 164.080 17.700 164.670 ;
        RECT 18.920 164.500 19.090 164.880 ;
        RECT 20.025 164.760 20.195 165.220 ;
        RECT 20.365 164.930 20.735 165.390 ;
        RECT 21.030 164.790 21.200 165.130 ;
        RECT 21.370 164.960 21.700 165.390 ;
        RECT 21.935 164.790 22.105 165.130 ;
        RECT 17.870 164.330 19.090 164.500 ;
        RECT 19.260 164.420 19.720 164.710 ;
        RECT 20.025 164.590 20.585 164.760 ;
        RECT 21.030 164.620 22.105 164.790 ;
        RECT 22.275 164.890 22.955 165.220 ;
        RECT 23.170 164.890 23.420 165.220 ;
        RECT 23.590 164.930 23.840 165.390 ;
        RECT 20.415 164.450 20.585 164.590 ;
        RECT 19.260 164.410 20.225 164.420 ;
        RECT 18.920 164.240 19.090 164.330 ;
        RECT 19.550 164.250 20.225 164.410 ;
        RECT 16.960 164.050 17.700 164.080 ;
        RECT 16.960 163.750 17.875 164.050 ;
        RECT 17.550 163.575 17.875 163.750 ;
        RECT 16.580 163.020 16.835 163.550 ;
        RECT 17.005 162.840 17.310 163.300 ;
        RECT 17.555 163.220 17.875 163.575 ;
        RECT 18.045 163.790 18.585 164.160 ;
        RECT 18.920 164.070 19.325 164.240 ;
        RECT 18.045 163.390 18.285 163.790 ;
        RECT 18.765 163.620 18.985 163.900 ;
        RECT 18.455 163.450 18.985 163.620 ;
        RECT 18.455 163.220 18.625 163.450 ;
        RECT 19.155 163.290 19.325 164.070 ;
        RECT 19.495 163.460 19.845 164.080 ;
        RECT 20.015 163.460 20.225 164.250 ;
        RECT 20.415 164.280 21.915 164.450 ;
        RECT 20.415 163.590 20.585 164.280 ;
        RECT 22.275 164.110 22.445 164.890 ;
        RECT 23.250 164.760 23.420 164.890 ;
        RECT 20.755 163.940 22.445 164.110 ;
        RECT 22.615 164.330 23.080 164.720 ;
        RECT 23.250 164.590 23.645 164.760 ;
        RECT 20.755 163.760 20.925 163.940 ;
        RECT 17.555 163.050 18.625 163.220 ;
        RECT 18.795 162.840 18.985 163.280 ;
        RECT 19.155 163.010 20.105 163.290 ;
        RECT 20.415 163.200 20.675 163.590 ;
        RECT 21.095 163.520 21.885 163.770 ;
        RECT 20.325 163.030 20.675 163.200 ;
        RECT 20.885 162.840 21.215 163.300 ;
        RECT 22.090 163.230 22.260 163.940 ;
        RECT 22.615 163.740 22.785 164.330 ;
        RECT 22.430 163.520 22.785 163.740 ;
        RECT 22.955 163.520 23.305 164.140 ;
        RECT 23.475 163.230 23.645 164.590 ;
        RECT 24.010 164.420 24.335 165.205 ;
        RECT 23.815 163.370 24.275 164.420 ;
        RECT 22.090 163.060 22.945 163.230 ;
        RECT 23.150 163.060 23.645 163.230 ;
        RECT 23.815 162.840 24.145 163.200 ;
        RECT 24.505 163.100 24.675 165.220 ;
        RECT 24.845 164.890 25.175 165.390 ;
        RECT 25.345 164.720 25.600 165.220 ;
        RECT 24.850 164.550 25.600 164.720 ;
        RECT 24.850 163.560 25.080 164.550 ;
        RECT 25.250 163.730 25.600 164.380 ;
        RECT 26.365 164.220 26.695 165.390 ;
        RECT 26.895 164.050 27.225 165.220 ;
        RECT 27.425 164.220 27.755 165.390 ;
        RECT 27.955 164.050 28.315 165.220 ;
        RECT 28.485 164.250 28.815 165.390 ;
        RECT 29.000 164.200 29.255 165.080 ;
        RECT 29.425 164.250 29.730 165.390 ;
        RECT 30.070 165.010 30.400 165.390 ;
        RECT 30.580 164.840 30.750 165.130 ;
        RECT 30.920 164.930 31.170 165.390 ;
        RECT 29.950 164.670 30.750 164.840 ;
        RECT 31.340 164.880 32.210 165.220 ;
        RECT 26.895 163.770 28.315 164.050 ;
        RECT 24.850 163.390 25.600 163.560 ;
        RECT 24.845 162.840 25.175 163.220 ;
        RECT 25.345 163.100 25.600 163.390 ;
        RECT 26.905 162.840 27.235 163.530 ;
        RECT 27.955 163.435 28.315 163.770 ;
        RECT 28.485 163.500 28.825 164.080 ;
        RECT 29.000 163.550 29.210 164.200 ;
        RECT 29.950 164.080 30.120 164.670 ;
        RECT 31.340 164.500 31.510 164.880 ;
        RECT 32.445 164.760 32.615 165.220 ;
        RECT 32.785 164.930 33.155 165.390 ;
        RECT 33.450 164.790 33.620 165.130 ;
        RECT 33.790 164.960 34.120 165.390 ;
        RECT 34.355 164.790 34.525 165.130 ;
        RECT 30.290 164.330 31.510 164.500 ;
        RECT 31.680 164.420 32.140 164.710 ;
        RECT 32.445 164.590 33.005 164.760 ;
        RECT 33.450 164.620 34.525 164.790 ;
        RECT 34.695 164.890 35.375 165.220 ;
        RECT 35.590 164.890 35.840 165.220 ;
        RECT 36.010 164.930 36.260 165.390 ;
        RECT 32.835 164.450 33.005 164.590 ;
        RECT 31.680 164.410 32.645 164.420 ;
        RECT 31.340 164.240 31.510 164.330 ;
        RECT 31.970 164.250 32.645 164.410 ;
        RECT 29.380 164.050 30.120 164.080 ;
        RECT 29.380 163.750 30.295 164.050 ;
        RECT 29.970 163.575 30.295 163.750 ;
        RECT 27.695 163.010 28.315 163.435 ;
        RECT 28.485 162.840 28.815 163.330 ;
        RECT 29.000 163.020 29.255 163.550 ;
        RECT 29.425 162.840 29.730 163.300 ;
        RECT 29.975 163.220 30.295 163.575 ;
        RECT 30.465 163.790 31.005 164.160 ;
        RECT 31.340 164.070 31.745 164.240 ;
        RECT 30.465 163.390 30.705 163.790 ;
        RECT 31.185 163.620 31.405 163.900 ;
        RECT 30.875 163.450 31.405 163.620 ;
        RECT 30.875 163.220 31.045 163.450 ;
        RECT 31.575 163.290 31.745 164.070 ;
        RECT 31.915 163.460 32.265 164.080 ;
        RECT 32.435 163.460 32.645 164.250 ;
        RECT 32.835 164.280 34.335 164.450 ;
        RECT 32.835 163.590 33.005 164.280 ;
        RECT 34.695 164.110 34.865 164.890 ;
        RECT 35.670 164.760 35.840 164.890 ;
        RECT 33.175 163.940 34.865 164.110 ;
        RECT 35.035 164.330 35.500 164.720 ;
        RECT 35.670 164.590 36.065 164.760 ;
        RECT 33.175 163.760 33.345 163.940 ;
        RECT 29.975 163.050 31.045 163.220 ;
        RECT 31.215 162.840 31.405 163.280 ;
        RECT 31.575 163.010 32.525 163.290 ;
        RECT 32.835 163.200 33.095 163.590 ;
        RECT 33.515 163.520 34.305 163.770 ;
        RECT 32.745 163.030 33.095 163.200 ;
        RECT 33.305 162.840 33.635 163.300 ;
        RECT 34.510 163.230 34.680 163.940 ;
        RECT 35.035 163.740 35.205 164.330 ;
        RECT 34.850 163.520 35.205 163.740 ;
        RECT 35.375 163.520 35.725 164.140 ;
        RECT 35.895 163.230 36.065 164.590 ;
        RECT 36.430 164.420 36.755 165.205 ;
        RECT 36.235 163.370 36.695 164.420 ;
        RECT 34.510 163.060 35.365 163.230 ;
        RECT 35.570 163.060 36.065 163.230 ;
        RECT 36.235 162.840 36.565 163.200 ;
        RECT 36.925 163.100 37.095 165.220 ;
        RECT 37.265 164.890 37.595 165.390 ;
        RECT 37.765 164.720 38.020 165.220 ;
        RECT 37.270 164.550 38.020 164.720 ;
        RECT 37.270 163.560 37.500 164.550 ;
        RECT 37.670 163.730 38.020 164.380 ;
        RECT 38.195 164.225 38.485 165.390 ;
        RECT 38.655 164.315 38.925 165.220 ;
        RECT 39.095 164.630 39.425 165.390 ;
        RECT 39.605 164.460 39.775 165.220 ;
        RECT 37.270 163.390 38.020 163.560 ;
        RECT 37.265 162.840 37.595 163.220 ;
        RECT 37.765 163.100 38.020 163.390 ;
        RECT 38.195 162.840 38.485 163.565 ;
        RECT 38.655 163.515 38.825 164.315 ;
        RECT 39.110 164.290 39.775 164.460 ;
        RECT 40.035 164.300 41.705 165.390 ;
        RECT 41.875 164.630 42.390 165.040 ;
        RECT 42.625 164.630 42.795 165.390 ;
        RECT 42.965 165.050 44.995 165.220 ;
        RECT 39.110 164.145 39.280 164.290 ;
        RECT 38.995 163.815 39.280 164.145 ;
        RECT 39.110 163.560 39.280 163.815 ;
        RECT 39.515 163.740 39.845 164.110 ;
        RECT 40.035 163.780 40.785 164.300 ;
        RECT 40.955 163.610 41.705 164.130 ;
        RECT 41.875 163.820 42.215 164.630 ;
        RECT 42.965 164.385 43.135 165.050 ;
        RECT 43.530 164.710 44.655 164.880 ;
        RECT 42.385 164.195 43.135 164.385 ;
        RECT 43.305 164.370 44.315 164.540 ;
        RECT 41.875 163.650 43.105 163.820 ;
        RECT 38.655 163.010 38.915 163.515 ;
        RECT 39.110 163.390 39.775 163.560 ;
        RECT 39.095 162.840 39.425 163.220 ;
        RECT 39.605 163.010 39.775 163.390 ;
        RECT 40.035 162.840 41.705 163.610 ;
        RECT 42.150 163.045 42.395 163.650 ;
        RECT 42.615 162.840 43.125 163.375 ;
        RECT 43.305 163.010 43.495 164.370 ;
        RECT 43.665 164.030 43.940 164.170 ;
        RECT 43.665 163.860 43.945 164.030 ;
        RECT 43.665 163.010 43.940 163.860 ;
        RECT 44.145 163.570 44.315 164.370 ;
        RECT 44.485 163.580 44.655 164.710 ;
        RECT 44.825 164.080 44.995 165.050 ;
        RECT 45.165 164.250 45.335 165.390 ;
        RECT 45.505 164.250 45.840 165.220 ;
        RECT 44.825 163.750 45.020 164.080 ;
        RECT 45.245 163.750 45.500 164.080 ;
        RECT 45.245 163.580 45.415 163.750 ;
        RECT 45.670 163.580 45.840 164.250 ;
        RECT 46.015 164.630 46.530 165.040 ;
        RECT 46.765 164.630 46.935 165.390 ;
        RECT 47.105 165.050 49.135 165.220 ;
        RECT 46.015 163.820 46.355 164.630 ;
        RECT 47.105 164.385 47.275 165.050 ;
        RECT 47.670 164.710 48.795 164.880 ;
        RECT 46.525 164.195 47.275 164.385 ;
        RECT 47.445 164.370 48.455 164.540 ;
        RECT 46.015 163.650 47.245 163.820 ;
        RECT 44.485 163.410 45.415 163.580 ;
        RECT 44.485 163.375 44.660 163.410 ;
        RECT 44.130 163.010 44.660 163.375 ;
        RECT 45.085 162.840 45.415 163.240 ;
        RECT 45.585 163.010 45.840 163.580 ;
        RECT 46.290 163.045 46.535 163.650 ;
        RECT 46.755 162.840 47.265 163.375 ;
        RECT 47.445 163.010 47.635 164.370 ;
        RECT 47.805 164.030 48.080 164.170 ;
        RECT 47.805 163.860 48.085 164.030 ;
        RECT 47.805 163.010 48.080 163.860 ;
        RECT 48.285 163.570 48.455 164.370 ;
        RECT 48.625 163.580 48.795 164.710 ;
        RECT 48.965 164.080 49.135 165.050 ;
        RECT 49.305 164.250 49.475 165.390 ;
        RECT 49.645 164.250 49.980 165.220 ;
        RECT 48.965 163.750 49.160 164.080 ;
        RECT 49.385 163.750 49.640 164.080 ;
        RECT 49.385 163.580 49.555 163.750 ;
        RECT 49.810 163.580 49.980 164.250 ;
        RECT 50.155 164.300 51.825 165.390 ;
        RECT 52.085 164.460 52.255 165.220 ;
        RECT 52.435 164.630 52.765 165.390 ;
        RECT 50.155 163.780 50.905 164.300 ;
        RECT 52.085 164.290 52.750 164.460 ;
        RECT 52.935 164.315 53.205 165.220 ;
        RECT 54.350 164.520 54.635 165.390 ;
        RECT 54.805 164.760 55.065 165.220 ;
        RECT 55.240 164.930 55.495 165.390 ;
        RECT 55.665 164.760 55.925 165.220 ;
        RECT 54.805 164.590 55.925 164.760 ;
        RECT 56.095 164.590 56.405 165.390 ;
        RECT 54.805 164.340 55.065 164.590 ;
        RECT 56.575 164.420 56.885 165.220 ;
        RECT 52.580 164.145 52.750 164.290 ;
        RECT 51.075 163.610 51.825 164.130 ;
        RECT 52.015 163.740 52.345 164.110 ;
        RECT 52.580 163.815 52.865 164.145 ;
        RECT 48.625 163.410 49.555 163.580 ;
        RECT 48.625 163.375 48.800 163.410 ;
        RECT 48.270 163.010 48.800 163.375 ;
        RECT 49.225 162.840 49.555 163.240 ;
        RECT 49.725 163.010 49.980 163.580 ;
        RECT 50.155 162.840 51.825 163.610 ;
        RECT 52.580 163.560 52.750 163.815 ;
        RECT 52.085 163.390 52.750 163.560 ;
        RECT 53.035 163.515 53.205 164.315 ;
        RECT 52.085 163.010 52.255 163.390 ;
        RECT 52.435 162.840 52.765 163.220 ;
        RECT 52.945 163.010 53.205 163.515 ;
        RECT 54.310 164.170 55.065 164.340 ;
        RECT 55.855 164.250 56.885 164.420 ;
        RECT 54.310 163.660 54.715 164.170 ;
        RECT 55.855 164.000 56.025 164.250 ;
        RECT 54.885 163.830 56.025 164.000 ;
        RECT 54.310 163.490 55.960 163.660 ;
        RECT 56.195 163.510 56.545 164.080 ;
        RECT 54.355 162.840 54.635 163.320 ;
        RECT 54.805 163.100 55.065 163.490 ;
        RECT 55.240 162.840 55.495 163.320 ;
        RECT 55.665 163.100 55.960 163.490 ;
        RECT 56.715 163.340 56.885 164.250 ;
        RECT 57.205 164.240 57.535 165.390 ;
        RECT 57.705 164.370 57.875 165.220 ;
        RECT 58.045 164.590 58.375 165.390 ;
        RECT 58.545 164.370 58.715 165.220 ;
        RECT 58.895 164.590 59.135 165.390 ;
        RECT 59.305 164.410 59.635 165.220 ;
        RECT 59.870 164.520 60.155 165.390 ;
        RECT 60.325 164.760 60.585 165.220 ;
        RECT 60.760 164.930 61.015 165.390 ;
        RECT 61.185 164.760 61.445 165.220 ;
        RECT 60.325 164.590 61.445 164.760 ;
        RECT 61.615 164.590 61.925 165.390 ;
        RECT 57.705 164.200 58.715 164.370 ;
        RECT 58.920 164.240 59.635 164.410 ;
        RECT 60.325 164.340 60.585 164.590 ;
        RECT 62.095 164.420 62.405 165.220 ;
        RECT 57.705 163.660 58.200 164.200 ;
        RECT 58.920 164.000 59.090 164.240 ;
        RECT 59.830 164.170 60.585 164.340 ;
        RECT 61.375 164.250 62.405 164.420 ;
        RECT 58.590 163.830 59.090 164.000 ;
        RECT 59.260 163.830 59.640 164.070 ;
        RECT 58.920 163.660 59.090 163.830 ;
        RECT 59.830 163.660 60.235 164.170 ;
        RECT 61.375 164.000 61.545 164.250 ;
        RECT 60.405 163.830 61.545 164.000 ;
        RECT 56.140 162.840 56.415 163.320 ;
        RECT 56.585 163.010 56.885 163.340 ;
        RECT 57.205 162.840 57.535 163.640 ;
        RECT 57.705 163.490 58.715 163.660 ;
        RECT 58.920 163.490 59.555 163.660 ;
        RECT 59.830 163.490 61.480 163.660 ;
        RECT 61.715 163.510 62.065 164.080 ;
        RECT 57.705 163.010 57.875 163.490 ;
        RECT 58.045 162.840 58.375 163.320 ;
        RECT 58.545 163.010 58.715 163.490 ;
        RECT 58.965 162.840 59.205 163.320 ;
        RECT 59.385 163.010 59.555 163.490 ;
        RECT 59.875 162.840 60.155 163.320 ;
        RECT 60.325 163.100 60.585 163.490 ;
        RECT 60.760 162.840 61.015 163.320 ;
        RECT 61.185 163.100 61.480 163.490 ;
        RECT 62.235 163.340 62.405 164.250 ;
        RECT 62.575 164.300 63.785 165.390 ;
        RECT 62.575 163.760 63.095 164.300 ;
        RECT 63.955 164.225 64.245 165.390 ;
        RECT 64.415 164.300 67.925 165.390 ;
        RECT 68.470 164.410 68.725 165.080 ;
        RECT 68.905 164.590 69.190 165.390 ;
        RECT 69.370 164.670 69.700 165.180 ;
        RECT 68.470 164.370 68.650 164.410 ;
        RECT 63.265 163.590 63.785 164.130 ;
        RECT 64.415 163.780 66.105 164.300 ;
        RECT 68.385 164.200 68.650 164.370 ;
        RECT 66.275 163.610 67.925 164.130 ;
        RECT 61.660 162.840 61.935 163.320 ;
        RECT 62.105 163.010 62.405 163.340 ;
        RECT 62.575 162.840 63.785 163.590 ;
        RECT 63.955 162.840 64.245 163.565 ;
        RECT 64.415 162.840 67.925 163.610 ;
        RECT 68.470 163.550 68.650 164.200 ;
        RECT 69.370 164.080 69.620 164.670 ;
        RECT 69.970 164.520 70.140 165.130 ;
        RECT 70.310 164.700 70.640 165.390 ;
        RECT 70.870 164.840 71.110 165.130 ;
        RECT 71.310 165.010 71.730 165.390 ;
        RECT 71.910 164.920 72.540 165.170 ;
        RECT 73.010 165.010 73.340 165.390 ;
        RECT 71.910 164.840 72.080 164.920 ;
        RECT 73.510 164.840 73.680 165.130 ;
        RECT 73.860 165.010 74.240 165.390 ;
        RECT 74.480 165.005 75.310 165.175 ;
        RECT 70.870 164.670 72.080 164.840 ;
        RECT 68.820 163.750 69.620 164.080 ;
        RECT 68.470 163.020 68.725 163.550 ;
        RECT 68.905 162.840 69.190 163.300 ;
        RECT 69.370 163.100 69.620 163.750 ;
        RECT 69.820 164.500 70.140 164.520 ;
        RECT 69.820 164.330 71.740 164.500 ;
        RECT 69.820 163.435 70.010 164.330 ;
        RECT 71.910 164.160 72.080 164.670 ;
        RECT 72.250 164.410 72.770 164.720 ;
        RECT 70.180 163.990 72.080 164.160 ;
        RECT 70.180 163.930 70.510 163.990 ;
        RECT 70.660 163.760 70.990 163.820 ;
        RECT 70.330 163.490 70.990 163.760 ;
        RECT 69.820 163.105 70.140 163.435 ;
        RECT 70.320 162.840 70.980 163.320 ;
        RECT 71.180 163.230 71.350 163.990 ;
        RECT 72.250 163.820 72.430 164.230 ;
        RECT 71.520 163.650 71.850 163.770 ;
        RECT 72.600 163.650 72.770 164.410 ;
        RECT 71.520 163.480 72.770 163.650 ;
        RECT 72.940 164.590 74.310 164.840 ;
        RECT 72.940 163.820 73.130 164.590 ;
        RECT 74.060 164.330 74.310 164.590 ;
        RECT 73.300 164.160 73.550 164.320 ;
        RECT 74.480 164.160 74.650 165.005 ;
        RECT 75.545 164.720 75.715 165.220 ;
        RECT 75.885 164.890 76.215 165.390 ;
        RECT 74.820 164.330 75.320 164.710 ;
        RECT 75.545 164.550 76.240 164.720 ;
        RECT 73.300 163.990 74.650 164.160 ;
        RECT 74.230 163.950 74.650 163.990 ;
        RECT 72.940 163.480 73.360 163.820 ;
        RECT 73.650 163.490 74.060 163.820 ;
        RECT 71.180 163.060 72.030 163.230 ;
        RECT 72.590 162.840 72.910 163.300 ;
        RECT 73.110 163.050 73.360 163.480 ;
        RECT 73.650 162.840 74.060 163.280 ;
        RECT 74.230 163.220 74.400 163.950 ;
        RECT 74.570 163.400 74.920 163.770 ;
        RECT 75.100 163.460 75.320 164.330 ;
        RECT 75.490 163.760 75.900 164.380 ;
        RECT 76.070 163.580 76.240 164.550 ;
        RECT 75.545 163.390 76.240 163.580 ;
        RECT 74.230 163.020 75.245 163.220 ;
        RECT 75.545 163.060 75.715 163.390 ;
        RECT 75.885 162.840 76.215 163.220 ;
        RECT 76.430 163.100 76.655 165.220 ;
        RECT 76.825 164.890 77.155 165.390 ;
        RECT 77.325 164.720 77.495 165.220 ;
        RECT 76.830 164.550 77.495 164.720 ;
        RECT 76.830 163.560 77.060 164.550 ;
        RECT 77.230 163.730 77.580 164.380 ;
        RECT 77.755 164.315 78.025 165.220 ;
        RECT 78.195 164.630 78.525 165.390 ;
        RECT 78.705 164.460 78.875 165.220 ;
        RECT 79.140 164.955 84.485 165.390 ;
        RECT 76.830 163.390 77.495 163.560 ;
        RECT 76.825 162.840 77.155 163.220 ;
        RECT 77.325 163.100 77.495 163.390 ;
        RECT 77.755 163.515 77.925 164.315 ;
        RECT 78.210 164.290 78.875 164.460 ;
        RECT 78.210 164.145 78.380 164.290 ;
        RECT 78.095 163.815 78.380 164.145 ;
        RECT 78.210 163.560 78.380 163.815 ;
        RECT 78.615 163.740 78.945 164.110 ;
        RECT 80.730 163.705 81.080 164.955 ;
        RECT 84.655 164.630 85.170 165.040 ;
        RECT 85.405 164.630 85.575 165.390 ;
        RECT 85.745 165.050 87.775 165.220 ;
        RECT 77.755 163.010 78.015 163.515 ;
        RECT 78.210 163.390 78.875 163.560 ;
        RECT 78.195 162.840 78.525 163.220 ;
        RECT 78.705 163.010 78.875 163.390 ;
        RECT 82.560 163.385 82.900 164.215 ;
        RECT 84.655 163.820 84.995 164.630 ;
        RECT 85.745 164.385 85.915 165.050 ;
        RECT 86.310 164.710 87.435 164.880 ;
        RECT 85.165 164.195 85.915 164.385 ;
        RECT 86.085 164.370 87.095 164.540 ;
        RECT 84.655 163.650 85.885 163.820 ;
        RECT 79.140 162.840 84.485 163.385 ;
        RECT 84.930 163.045 85.175 163.650 ;
        RECT 85.395 162.840 85.905 163.375 ;
        RECT 86.085 163.010 86.275 164.370 ;
        RECT 86.445 163.690 86.720 164.170 ;
        RECT 86.445 163.520 86.725 163.690 ;
        RECT 86.925 163.570 87.095 164.370 ;
        RECT 87.265 163.580 87.435 164.710 ;
        RECT 87.605 164.080 87.775 165.050 ;
        RECT 87.945 164.250 88.115 165.390 ;
        RECT 88.285 164.250 88.620 165.220 ;
        RECT 87.605 163.750 87.800 164.080 ;
        RECT 88.025 163.750 88.280 164.080 ;
        RECT 88.025 163.580 88.195 163.750 ;
        RECT 88.450 163.580 88.620 164.250 ;
        RECT 89.715 164.225 90.005 165.390 ;
        RECT 91.095 164.630 91.610 165.040 ;
        RECT 91.845 164.630 92.015 165.390 ;
        RECT 92.185 165.050 94.215 165.220 ;
        RECT 91.095 163.820 91.435 164.630 ;
        RECT 92.185 164.385 92.355 165.050 ;
        RECT 92.750 164.710 93.875 164.880 ;
        RECT 91.605 164.195 92.355 164.385 ;
        RECT 92.525 164.370 93.535 164.540 ;
        RECT 91.095 163.650 92.325 163.820 ;
        RECT 86.445 163.010 86.720 163.520 ;
        RECT 87.265 163.410 88.195 163.580 ;
        RECT 87.265 163.375 87.440 163.410 ;
        RECT 86.910 163.010 87.440 163.375 ;
        RECT 87.865 162.840 88.195 163.240 ;
        RECT 88.365 163.010 88.620 163.580 ;
        RECT 89.715 162.840 90.005 163.565 ;
        RECT 91.370 163.045 91.615 163.650 ;
        RECT 91.835 162.840 92.345 163.375 ;
        RECT 92.525 163.010 92.715 164.370 ;
        RECT 92.885 164.030 93.160 164.170 ;
        RECT 92.885 163.860 93.165 164.030 ;
        RECT 92.885 163.010 93.160 163.860 ;
        RECT 93.365 163.570 93.535 164.370 ;
        RECT 93.705 163.580 93.875 164.710 ;
        RECT 94.045 164.080 94.215 165.050 ;
        RECT 94.385 164.250 94.555 165.390 ;
        RECT 94.725 164.250 95.060 165.220 ;
        RECT 95.325 164.460 95.495 165.220 ;
        RECT 95.675 164.630 96.005 165.390 ;
        RECT 95.325 164.290 95.990 164.460 ;
        RECT 96.175 164.315 96.445 165.220 ;
        RECT 94.045 163.750 94.240 164.080 ;
        RECT 94.465 163.750 94.720 164.080 ;
        RECT 94.465 163.580 94.635 163.750 ;
        RECT 94.890 163.580 95.060 164.250 ;
        RECT 95.820 164.145 95.990 164.290 ;
        RECT 95.255 163.740 95.585 164.110 ;
        RECT 95.820 163.815 96.105 164.145 ;
        RECT 93.705 163.410 94.635 163.580 ;
        RECT 93.705 163.375 93.880 163.410 ;
        RECT 93.350 163.010 93.880 163.375 ;
        RECT 94.305 162.840 94.635 163.240 ;
        RECT 94.805 163.010 95.060 163.580 ;
        RECT 95.820 163.560 95.990 163.815 ;
        RECT 95.325 163.390 95.990 163.560 ;
        RECT 96.275 163.515 96.445 164.315 ;
        RECT 95.325 163.010 95.495 163.390 ;
        RECT 95.675 162.840 96.005 163.220 ;
        RECT 96.185 163.010 96.445 163.515 ;
        RECT 96.620 164.250 96.955 165.220 ;
        RECT 97.125 164.250 97.295 165.390 ;
        RECT 97.465 165.050 99.495 165.220 ;
        RECT 96.620 163.580 96.790 164.250 ;
        RECT 97.465 164.080 97.635 165.050 ;
        RECT 96.960 163.750 97.215 164.080 ;
        RECT 97.440 163.750 97.635 164.080 ;
        RECT 97.805 164.710 98.930 164.880 ;
        RECT 97.045 163.580 97.215 163.750 ;
        RECT 97.805 163.580 97.975 164.710 ;
        RECT 96.620 163.010 96.875 163.580 ;
        RECT 97.045 163.410 97.975 163.580 ;
        RECT 98.145 164.370 99.155 164.540 ;
        RECT 98.145 163.570 98.315 164.370 ;
        RECT 97.800 163.375 97.975 163.410 ;
        RECT 97.045 162.840 97.375 163.240 ;
        RECT 97.800 163.010 98.330 163.375 ;
        RECT 98.520 163.350 98.795 164.170 ;
        RECT 98.515 163.180 98.795 163.350 ;
        RECT 98.520 163.010 98.795 163.180 ;
        RECT 98.965 163.010 99.155 164.370 ;
        RECT 99.325 164.385 99.495 165.050 ;
        RECT 99.665 164.630 99.835 165.390 ;
        RECT 100.070 164.630 100.585 165.040 ;
        RECT 99.325 164.195 100.075 164.385 ;
        RECT 100.245 163.820 100.585 164.630 ;
        RECT 101.715 164.250 101.945 165.390 ;
        RECT 102.115 164.240 102.445 165.220 ;
        RECT 102.615 164.250 102.825 165.390 ;
        RECT 101.695 163.830 102.025 164.080 ;
        RECT 99.355 163.650 100.585 163.820 ;
        RECT 99.335 162.840 99.845 163.375 ;
        RECT 100.065 163.045 100.310 163.650 ;
        RECT 101.715 162.840 101.945 163.660 ;
        RECT 102.195 163.640 102.445 164.240 ;
        RECT 103.060 164.200 103.315 165.080 ;
        RECT 103.485 164.250 103.790 165.390 ;
        RECT 104.130 165.010 104.460 165.390 ;
        RECT 104.640 164.840 104.810 165.130 ;
        RECT 104.980 164.930 105.230 165.390 ;
        RECT 104.010 164.670 104.810 164.840 ;
        RECT 105.400 164.880 106.270 165.220 ;
        RECT 102.115 163.010 102.445 163.640 ;
        RECT 102.615 162.840 102.825 163.660 ;
        RECT 103.060 163.550 103.270 164.200 ;
        RECT 104.010 164.080 104.180 164.670 ;
        RECT 105.400 164.500 105.570 164.880 ;
        RECT 106.505 164.760 106.675 165.220 ;
        RECT 106.845 164.930 107.215 165.390 ;
        RECT 107.510 164.790 107.680 165.130 ;
        RECT 107.850 164.960 108.180 165.390 ;
        RECT 108.415 164.790 108.585 165.130 ;
        RECT 104.350 164.330 105.570 164.500 ;
        RECT 105.740 164.420 106.200 164.710 ;
        RECT 106.505 164.590 107.065 164.760 ;
        RECT 107.510 164.620 108.585 164.790 ;
        RECT 108.755 164.890 109.435 165.220 ;
        RECT 109.650 164.890 109.900 165.220 ;
        RECT 110.070 164.930 110.320 165.390 ;
        RECT 106.895 164.450 107.065 164.590 ;
        RECT 105.740 164.410 106.705 164.420 ;
        RECT 105.400 164.240 105.570 164.330 ;
        RECT 106.030 164.250 106.705 164.410 ;
        RECT 103.440 164.050 104.180 164.080 ;
        RECT 103.440 163.750 104.355 164.050 ;
        RECT 104.030 163.575 104.355 163.750 ;
        RECT 103.060 163.020 103.315 163.550 ;
        RECT 103.485 162.840 103.790 163.300 ;
        RECT 104.035 163.220 104.355 163.575 ;
        RECT 104.525 163.790 105.065 164.160 ;
        RECT 105.400 164.070 105.805 164.240 ;
        RECT 104.525 163.390 104.765 163.790 ;
        RECT 105.245 163.620 105.465 163.900 ;
        RECT 104.935 163.450 105.465 163.620 ;
        RECT 104.935 163.220 105.105 163.450 ;
        RECT 105.635 163.290 105.805 164.070 ;
        RECT 105.975 163.460 106.325 164.080 ;
        RECT 106.495 163.460 106.705 164.250 ;
        RECT 106.895 164.280 108.395 164.450 ;
        RECT 106.895 163.590 107.065 164.280 ;
        RECT 108.755 164.110 108.925 164.890 ;
        RECT 109.730 164.760 109.900 164.890 ;
        RECT 107.235 163.940 108.925 164.110 ;
        RECT 109.095 164.330 109.560 164.720 ;
        RECT 109.730 164.590 110.125 164.760 ;
        RECT 107.235 163.760 107.405 163.940 ;
        RECT 104.035 163.050 105.105 163.220 ;
        RECT 105.275 162.840 105.465 163.280 ;
        RECT 105.635 163.010 106.585 163.290 ;
        RECT 106.895 163.200 107.155 163.590 ;
        RECT 107.575 163.520 108.365 163.770 ;
        RECT 106.805 163.030 107.155 163.200 ;
        RECT 107.365 162.840 107.695 163.300 ;
        RECT 108.570 163.230 108.740 163.940 ;
        RECT 109.095 163.740 109.265 164.330 ;
        RECT 108.910 163.520 109.265 163.740 ;
        RECT 109.435 163.520 109.785 164.140 ;
        RECT 109.955 163.230 110.125 164.590 ;
        RECT 110.490 164.420 110.815 165.205 ;
        RECT 110.295 163.370 110.755 164.420 ;
        RECT 108.570 163.060 109.425 163.230 ;
        RECT 109.630 163.060 110.125 163.230 ;
        RECT 110.295 162.840 110.625 163.200 ;
        RECT 110.985 163.100 111.155 165.220 ;
        RECT 111.325 164.890 111.655 165.390 ;
        RECT 111.825 164.720 112.080 165.220 ;
        RECT 111.330 164.550 112.080 164.720 ;
        RECT 111.330 163.560 111.560 164.550 ;
        RECT 111.730 163.730 112.080 164.380 ;
        RECT 112.255 164.315 112.525 165.220 ;
        RECT 112.695 164.630 113.025 165.390 ;
        RECT 113.205 164.460 113.375 165.220 ;
        RECT 111.330 163.390 112.080 163.560 ;
        RECT 111.325 162.840 111.655 163.220 ;
        RECT 111.825 163.100 112.080 163.390 ;
        RECT 112.255 163.515 112.425 164.315 ;
        RECT 112.710 164.290 113.375 164.460 ;
        RECT 114.555 164.300 115.765 165.390 ;
        RECT 112.710 164.145 112.880 164.290 ;
        RECT 112.595 163.815 112.880 164.145 ;
        RECT 112.710 163.560 112.880 163.815 ;
        RECT 113.115 163.740 113.445 164.110 ;
        RECT 114.555 163.760 115.075 164.300 ;
        RECT 115.245 163.590 115.765 164.130 ;
        RECT 112.255 163.010 112.515 163.515 ;
        RECT 112.710 163.390 113.375 163.560 ;
        RECT 112.695 162.840 113.025 163.220 ;
        RECT 113.205 163.010 113.375 163.390 ;
        RECT 114.555 162.840 115.765 163.590 ;
        RECT 10.510 162.670 115.850 162.840 ;
        RECT 10.595 161.920 11.805 162.670 ;
        RECT 10.595 161.380 11.115 161.920 ;
        RECT 12.435 161.900 15.025 162.670 ;
        RECT 11.285 161.210 11.805 161.750 ;
        RECT 10.595 160.120 11.805 161.210 ;
        RECT 12.435 161.210 13.645 161.730 ;
        RECT 13.815 161.380 15.025 161.900 ;
        RECT 15.235 161.850 15.465 162.670 ;
        RECT 15.635 161.870 15.965 162.500 ;
        RECT 15.215 161.430 15.545 161.680 ;
        RECT 15.715 161.270 15.965 161.870 ;
        RECT 16.135 161.850 16.345 162.670 ;
        RECT 16.850 161.860 17.095 162.465 ;
        RECT 17.315 162.135 17.825 162.670 ;
        RECT 12.435 160.120 15.025 161.210 ;
        RECT 15.235 160.120 15.465 161.260 ;
        RECT 15.635 160.290 15.965 161.270 ;
        RECT 16.575 161.690 17.805 161.860 ;
        RECT 16.135 160.120 16.345 161.260 ;
        RECT 16.575 160.880 16.915 161.690 ;
        RECT 17.085 161.125 17.835 161.315 ;
        RECT 16.575 160.470 17.090 160.880 ;
        RECT 17.325 160.120 17.495 160.880 ;
        RECT 17.665 160.460 17.835 161.125 ;
        RECT 18.005 161.140 18.195 162.500 ;
        RECT 18.365 161.650 18.640 162.500 ;
        RECT 18.830 162.135 19.360 162.500 ;
        RECT 19.785 162.270 20.115 162.670 ;
        RECT 19.185 162.100 19.360 162.135 ;
        RECT 18.365 161.480 18.645 161.650 ;
        RECT 18.365 161.340 18.640 161.480 ;
        RECT 18.845 161.140 19.015 161.940 ;
        RECT 18.005 160.970 19.015 161.140 ;
        RECT 19.185 161.930 20.115 162.100 ;
        RECT 20.285 161.930 20.540 162.500 ;
        RECT 19.185 160.800 19.355 161.930 ;
        RECT 19.945 161.760 20.115 161.930 ;
        RECT 18.230 160.630 19.355 160.800 ;
        RECT 19.525 161.430 19.720 161.760 ;
        RECT 19.945 161.430 20.200 161.760 ;
        RECT 19.525 160.460 19.695 161.430 ;
        RECT 20.370 161.260 20.540 161.930 ;
        RECT 17.665 160.290 19.695 160.460 ;
        RECT 19.865 160.120 20.035 161.260 ;
        RECT 20.205 160.290 20.540 161.260 ;
        RECT 20.720 161.930 20.975 162.500 ;
        RECT 21.145 162.270 21.475 162.670 ;
        RECT 21.900 162.135 22.430 162.500 ;
        RECT 21.900 162.100 22.075 162.135 ;
        RECT 21.145 161.930 22.075 162.100 ;
        RECT 20.720 161.260 20.890 161.930 ;
        RECT 21.145 161.760 21.315 161.930 ;
        RECT 21.060 161.430 21.315 161.760 ;
        RECT 21.540 161.430 21.735 161.760 ;
        RECT 20.720 160.290 21.055 161.260 ;
        RECT 21.225 160.120 21.395 161.260 ;
        RECT 21.565 160.460 21.735 161.430 ;
        RECT 21.905 160.800 22.075 161.930 ;
        RECT 22.245 161.140 22.415 161.940 ;
        RECT 22.620 161.650 22.895 162.500 ;
        RECT 22.615 161.480 22.895 161.650 ;
        RECT 22.620 161.340 22.895 161.480 ;
        RECT 23.065 161.140 23.255 162.500 ;
        RECT 23.435 162.135 23.945 162.670 ;
        RECT 24.165 161.860 24.410 162.465 ;
        RECT 25.315 161.945 25.605 162.670 ;
        RECT 25.780 162.120 26.035 162.410 ;
        RECT 26.205 162.290 26.535 162.670 ;
        RECT 25.780 161.950 26.530 162.120 ;
        RECT 23.455 161.690 24.685 161.860 ;
        RECT 22.245 160.970 23.255 161.140 ;
        RECT 23.425 161.125 24.175 161.315 ;
        RECT 21.905 160.630 23.030 160.800 ;
        RECT 23.425 160.460 23.595 161.125 ;
        RECT 24.345 160.880 24.685 161.690 ;
        RECT 21.565 160.290 23.595 160.460 ;
        RECT 23.765 160.120 23.935 160.880 ;
        RECT 24.170 160.470 24.685 160.880 ;
        RECT 25.315 160.120 25.605 161.285 ;
        RECT 25.780 161.130 26.130 161.780 ;
        RECT 26.300 160.960 26.530 161.950 ;
        RECT 25.780 160.790 26.530 160.960 ;
        RECT 25.780 160.290 26.035 160.790 ;
        RECT 26.205 160.120 26.535 160.620 ;
        RECT 26.705 160.290 26.875 162.410 ;
        RECT 27.235 162.310 27.565 162.670 ;
        RECT 27.735 162.280 28.230 162.450 ;
        RECT 28.435 162.280 29.290 162.450 ;
        RECT 27.105 161.090 27.565 162.140 ;
        RECT 27.045 160.305 27.370 161.090 ;
        RECT 27.735 160.920 27.905 162.280 ;
        RECT 28.075 161.370 28.425 161.990 ;
        RECT 28.595 161.770 28.950 161.990 ;
        RECT 28.595 161.180 28.765 161.770 ;
        RECT 29.120 161.570 29.290 162.280 ;
        RECT 30.165 162.210 30.495 162.670 ;
        RECT 30.705 162.310 31.055 162.480 ;
        RECT 29.495 161.740 30.285 161.990 ;
        RECT 30.705 161.920 30.965 162.310 ;
        RECT 31.275 162.220 32.225 162.500 ;
        RECT 32.395 162.230 32.585 162.670 ;
        RECT 32.755 162.290 33.825 162.460 ;
        RECT 30.455 161.570 30.625 161.750 ;
        RECT 27.735 160.750 28.130 160.920 ;
        RECT 28.300 160.790 28.765 161.180 ;
        RECT 28.935 161.400 30.625 161.570 ;
        RECT 27.960 160.620 28.130 160.750 ;
        RECT 28.935 160.620 29.105 161.400 ;
        RECT 30.795 161.230 30.965 161.920 ;
        RECT 29.465 161.060 30.965 161.230 ;
        RECT 31.155 161.260 31.365 162.050 ;
        RECT 31.535 161.430 31.885 162.050 ;
        RECT 32.055 161.440 32.225 162.220 ;
        RECT 32.755 162.060 32.925 162.290 ;
        RECT 32.395 161.890 32.925 162.060 ;
        RECT 32.395 161.610 32.615 161.890 ;
        RECT 33.095 161.720 33.335 162.120 ;
        RECT 32.055 161.270 32.460 161.440 ;
        RECT 32.795 161.350 33.335 161.720 ;
        RECT 33.505 161.935 33.825 162.290 ;
        RECT 34.070 162.210 34.375 162.670 ;
        RECT 34.545 161.960 34.800 162.490 ;
        RECT 33.505 161.760 33.830 161.935 ;
        RECT 33.505 161.460 34.420 161.760 ;
        RECT 33.680 161.430 34.420 161.460 ;
        RECT 31.155 161.100 31.830 161.260 ;
        RECT 32.290 161.180 32.460 161.270 ;
        RECT 31.155 161.090 32.120 161.100 ;
        RECT 30.795 160.920 30.965 161.060 ;
        RECT 27.540 160.120 27.790 160.580 ;
        RECT 27.960 160.290 28.210 160.620 ;
        RECT 28.425 160.290 29.105 160.620 ;
        RECT 29.275 160.720 30.350 160.890 ;
        RECT 30.795 160.750 31.355 160.920 ;
        RECT 31.660 160.800 32.120 161.090 ;
        RECT 32.290 161.010 33.510 161.180 ;
        RECT 29.275 160.380 29.445 160.720 ;
        RECT 29.680 160.120 30.010 160.550 ;
        RECT 30.180 160.380 30.350 160.720 ;
        RECT 30.645 160.120 31.015 160.580 ;
        RECT 31.185 160.290 31.355 160.750 ;
        RECT 32.290 160.630 32.460 161.010 ;
        RECT 33.680 160.840 33.850 161.430 ;
        RECT 34.590 161.310 34.800 161.960 ;
        RECT 31.590 160.290 32.460 160.630 ;
        RECT 33.050 160.670 33.850 160.840 ;
        RECT 32.630 160.120 32.880 160.580 ;
        RECT 33.050 160.380 33.220 160.670 ;
        RECT 33.400 160.120 33.730 160.500 ;
        RECT 34.070 160.120 34.375 161.260 ;
        RECT 34.545 160.430 34.800 161.310 ;
        RECT 35.440 161.930 35.695 162.500 ;
        RECT 35.865 162.270 36.195 162.670 ;
        RECT 36.620 162.135 37.150 162.500 ;
        RECT 36.620 162.100 36.795 162.135 ;
        RECT 35.865 161.930 36.795 162.100 ;
        RECT 37.340 161.990 37.615 162.500 ;
        RECT 35.440 161.260 35.610 161.930 ;
        RECT 35.865 161.760 36.035 161.930 ;
        RECT 35.780 161.430 36.035 161.760 ;
        RECT 36.260 161.430 36.455 161.760 ;
        RECT 35.440 160.290 35.775 161.260 ;
        RECT 35.945 160.120 36.115 161.260 ;
        RECT 36.285 160.460 36.455 161.430 ;
        RECT 36.625 160.800 36.795 161.930 ;
        RECT 36.965 161.140 37.135 161.940 ;
        RECT 37.335 161.820 37.615 161.990 ;
        RECT 37.340 161.340 37.615 161.820 ;
        RECT 37.785 161.140 37.975 162.500 ;
        RECT 38.155 162.135 38.665 162.670 ;
        RECT 38.885 161.860 39.130 162.465 ;
        RECT 39.575 161.920 40.785 162.670 ;
        RECT 38.175 161.690 39.405 161.860 ;
        RECT 36.965 160.970 37.975 161.140 ;
        RECT 38.145 161.125 38.895 161.315 ;
        RECT 36.625 160.630 37.750 160.800 ;
        RECT 38.145 160.460 38.315 161.125 ;
        RECT 39.065 160.880 39.405 161.690 ;
        RECT 36.285 160.290 38.315 160.460 ;
        RECT 38.485 160.120 38.655 160.880 ;
        RECT 38.890 160.470 39.405 160.880 ;
        RECT 39.575 161.210 40.095 161.750 ;
        RECT 40.265 161.380 40.785 161.920 ;
        RECT 41.160 161.890 41.660 162.500 ;
        RECT 40.955 161.430 41.305 161.680 ;
        RECT 41.490 161.260 41.660 161.890 ;
        RECT 42.290 162.020 42.620 162.500 ;
        RECT 42.790 162.210 43.015 162.670 ;
        RECT 43.185 162.020 43.515 162.500 ;
        RECT 42.290 161.850 43.515 162.020 ;
        RECT 43.705 161.870 43.955 162.670 ;
        RECT 44.125 161.870 44.465 162.500 ;
        RECT 41.830 161.480 42.160 161.680 ;
        RECT 42.330 161.480 42.660 161.680 ;
        RECT 42.830 161.480 43.250 161.680 ;
        RECT 43.425 161.510 44.120 161.680 ;
        RECT 43.425 161.260 43.595 161.510 ;
        RECT 44.290 161.260 44.465 161.870 ;
        RECT 39.575 160.120 40.785 161.210 ;
        RECT 41.160 161.090 43.595 161.260 ;
        RECT 41.160 160.290 41.490 161.090 ;
        RECT 41.660 160.120 41.990 160.920 ;
        RECT 42.290 160.290 42.620 161.090 ;
        RECT 43.265 160.120 43.515 160.920 ;
        RECT 43.785 160.120 43.955 161.260 ;
        RECT 44.125 160.290 44.465 161.260 ;
        RECT 45.095 161.995 45.355 162.500 ;
        RECT 45.535 162.290 45.865 162.670 ;
        RECT 46.045 162.120 46.215 162.500 ;
        RECT 45.095 161.195 45.265 161.995 ;
        RECT 45.550 161.950 46.215 162.120 ;
        RECT 45.550 161.695 45.720 161.950 ;
        RECT 46.935 161.900 49.525 162.670 ;
        RECT 45.435 161.365 45.720 161.695 ;
        RECT 45.955 161.400 46.285 161.770 ;
        RECT 45.550 161.220 45.720 161.365 ;
        RECT 45.095 160.290 45.365 161.195 ;
        RECT 45.550 161.050 46.215 161.220 ;
        RECT 45.535 160.120 45.865 160.880 ;
        RECT 46.045 160.290 46.215 161.050 ;
        RECT 46.935 161.210 48.145 161.730 ;
        RECT 48.315 161.380 49.525 161.900 ;
        RECT 49.735 161.850 49.965 162.670 ;
        RECT 50.135 161.870 50.465 162.500 ;
        RECT 49.715 161.430 50.045 161.680 ;
        RECT 50.215 161.270 50.465 161.870 ;
        RECT 50.635 161.850 50.845 162.670 ;
        RECT 51.075 161.945 51.365 162.670 ;
        RECT 52.000 162.125 57.345 162.670 ;
        RECT 46.935 160.120 49.525 161.210 ;
        RECT 49.735 160.120 49.965 161.260 ;
        RECT 50.135 160.290 50.465 161.270 ;
        RECT 50.635 160.120 50.845 161.260 ;
        RECT 51.075 160.120 51.365 161.285 ;
        RECT 53.590 160.555 53.940 161.805 ;
        RECT 55.420 161.295 55.760 162.125 ;
        RECT 57.520 161.830 57.780 162.670 ;
        RECT 57.955 161.925 58.210 162.500 ;
        RECT 58.380 162.290 58.710 162.670 ;
        RECT 58.925 162.120 59.095 162.500 ;
        RECT 58.380 161.950 59.095 162.120 ;
        RECT 52.000 160.120 57.345 160.555 ;
        RECT 57.520 160.120 57.780 161.270 ;
        RECT 57.955 161.195 58.125 161.925 ;
        RECT 58.380 161.760 58.550 161.950 ;
        RECT 59.360 161.830 59.620 162.670 ;
        RECT 59.795 161.925 60.050 162.500 ;
        RECT 60.220 162.290 60.550 162.670 ;
        RECT 60.765 162.120 60.935 162.500 ;
        RECT 60.220 161.950 60.935 162.120 ;
        RECT 61.285 162.120 61.455 162.500 ;
        RECT 61.670 162.290 62.000 162.670 ;
        RECT 61.285 161.950 62.000 162.120 ;
        RECT 58.295 161.430 58.550 161.760 ;
        RECT 58.380 161.220 58.550 161.430 ;
        RECT 58.830 161.400 59.185 161.770 ;
        RECT 57.955 160.290 58.210 161.195 ;
        RECT 58.380 161.050 59.095 161.220 ;
        RECT 58.380 160.120 58.710 160.880 ;
        RECT 58.925 160.290 59.095 161.050 ;
        RECT 59.360 160.120 59.620 161.270 ;
        RECT 59.795 161.195 59.965 161.925 ;
        RECT 60.220 161.760 60.390 161.950 ;
        RECT 60.135 161.430 60.390 161.760 ;
        RECT 60.220 161.220 60.390 161.430 ;
        RECT 60.670 161.400 61.025 161.770 ;
        RECT 61.195 161.400 61.550 161.770 ;
        RECT 61.830 161.760 62.000 161.950 ;
        RECT 62.170 161.925 62.425 162.500 ;
        RECT 61.830 161.430 62.085 161.760 ;
        RECT 61.830 161.220 62.000 161.430 ;
        RECT 59.795 160.290 60.050 161.195 ;
        RECT 60.220 161.050 60.935 161.220 ;
        RECT 60.220 160.120 60.550 160.880 ;
        RECT 60.765 160.290 60.935 161.050 ;
        RECT 61.285 161.050 62.000 161.220 ;
        RECT 62.255 161.195 62.425 161.925 ;
        RECT 62.600 161.830 62.860 162.670 ;
        RECT 63.125 162.120 63.295 162.500 ;
        RECT 63.510 162.290 63.840 162.670 ;
        RECT 63.125 161.950 63.840 162.120 ;
        RECT 63.035 161.400 63.390 161.770 ;
        RECT 63.670 161.760 63.840 161.950 ;
        RECT 64.010 161.925 64.265 162.500 ;
        RECT 63.670 161.430 63.925 161.760 ;
        RECT 61.285 160.290 61.455 161.050 ;
        RECT 61.670 160.120 62.000 160.880 ;
        RECT 62.170 160.290 62.425 161.195 ;
        RECT 62.600 160.120 62.860 161.270 ;
        RECT 63.670 161.220 63.840 161.430 ;
        RECT 63.125 161.050 63.840 161.220 ;
        RECT 64.095 161.195 64.265 161.925 ;
        RECT 64.440 161.830 64.700 162.670 ;
        RECT 65.800 162.125 71.145 162.670 ;
        RECT 63.125 160.290 63.295 161.050 ;
        RECT 63.510 160.120 63.840 160.880 ;
        RECT 64.010 160.290 64.265 161.195 ;
        RECT 64.440 160.120 64.700 161.270 ;
        RECT 67.390 160.555 67.740 161.805 ;
        RECT 69.220 161.295 69.560 162.125 ;
        RECT 71.375 161.850 71.585 162.670 ;
        RECT 71.755 161.870 72.085 162.500 ;
        RECT 71.755 161.270 72.005 161.870 ;
        RECT 72.255 161.850 72.485 162.670 ;
        RECT 72.970 161.860 73.215 162.465 ;
        RECT 73.435 162.135 73.945 162.670 ;
        RECT 72.695 161.690 73.925 161.860 ;
        RECT 72.175 161.430 72.505 161.680 ;
        RECT 65.800 160.120 71.145 160.555 ;
        RECT 71.375 160.120 71.585 161.260 ;
        RECT 71.755 160.290 72.085 161.270 ;
        RECT 72.255 160.120 72.485 161.260 ;
        RECT 72.695 160.880 73.035 161.690 ;
        RECT 73.205 161.125 73.955 161.315 ;
        RECT 72.695 160.470 73.210 160.880 ;
        RECT 73.445 160.120 73.615 160.880 ;
        RECT 73.785 160.460 73.955 161.125 ;
        RECT 74.125 161.140 74.315 162.500 ;
        RECT 74.485 161.650 74.760 162.500 ;
        RECT 74.950 162.135 75.480 162.500 ;
        RECT 75.905 162.270 76.235 162.670 ;
        RECT 75.305 162.100 75.480 162.135 ;
        RECT 74.485 161.480 74.765 161.650 ;
        RECT 74.485 161.340 74.760 161.480 ;
        RECT 74.965 161.140 75.135 161.940 ;
        RECT 74.125 160.970 75.135 161.140 ;
        RECT 75.305 161.930 76.235 162.100 ;
        RECT 76.405 161.930 76.660 162.500 ;
        RECT 76.835 161.945 77.125 162.670 ;
        RECT 75.305 160.800 75.475 161.930 ;
        RECT 76.065 161.760 76.235 161.930 ;
        RECT 74.350 160.630 75.475 160.800 ;
        RECT 75.645 161.430 75.840 161.760 ;
        RECT 76.065 161.430 76.320 161.760 ;
        RECT 75.645 160.460 75.815 161.430 ;
        RECT 76.490 161.260 76.660 161.930 ;
        RECT 77.355 161.850 77.565 162.670 ;
        RECT 77.735 161.870 78.065 162.500 ;
        RECT 73.785 160.290 75.815 160.460 ;
        RECT 75.985 160.120 76.155 161.260 ;
        RECT 76.325 160.290 76.660 161.260 ;
        RECT 76.835 160.120 77.125 161.285 ;
        RECT 77.735 161.270 77.985 161.870 ;
        RECT 78.235 161.850 78.465 162.670 ;
        RECT 79.225 162.120 79.395 162.500 ;
        RECT 79.575 162.290 79.905 162.670 ;
        RECT 79.225 161.950 79.890 162.120 ;
        RECT 80.085 161.995 80.345 162.500 ;
        RECT 78.155 161.430 78.485 161.680 ;
        RECT 79.155 161.400 79.485 161.770 ;
        RECT 79.720 161.695 79.890 161.950 ;
        RECT 79.720 161.365 80.005 161.695 ;
        RECT 77.355 160.120 77.565 161.260 ;
        RECT 77.735 160.290 78.065 161.270 ;
        RECT 78.235 160.120 78.465 161.260 ;
        RECT 79.720 161.220 79.890 161.365 ;
        RECT 79.225 161.050 79.890 161.220 ;
        RECT 80.175 161.195 80.345 161.995 ;
        RECT 80.890 161.990 81.145 162.490 ;
        RECT 81.325 162.210 81.610 162.670 ;
        RECT 80.805 161.960 81.145 161.990 ;
        RECT 80.805 161.820 81.070 161.960 ;
        RECT 79.225 160.290 79.395 161.050 ;
        RECT 79.575 160.120 79.905 160.880 ;
        RECT 80.075 160.290 80.345 161.195 ;
        RECT 80.890 161.100 81.070 161.820 ;
        RECT 81.790 161.760 82.040 162.410 ;
        RECT 81.240 161.430 82.040 161.760 ;
        RECT 80.890 160.430 81.145 161.100 ;
        RECT 81.325 160.120 81.610 160.920 ;
        RECT 81.790 160.840 82.040 161.430 ;
        RECT 82.240 162.075 82.560 162.405 ;
        RECT 82.740 162.190 83.400 162.670 ;
        RECT 83.600 162.280 84.450 162.450 ;
        RECT 82.240 161.180 82.430 162.075 ;
        RECT 82.750 161.750 83.410 162.020 ;
        RECT 83.080 161.690 83.410 161.750 ;
        RECT 82.600 161.520 82.930 161.580 ;
        RECT 83.600 161.520 83.770 162.280 ;
        RECT 85.010 162.210 85.330 162.670 ;
        RECT 85.530 162.030 85.780 162.460 ;
        RECT 86.070 162.230 86.480 162.670 ;
        RECT 86.650 162.290 87.665 162.490 ;
        RECT 83.940 161.860 85.190 162.030 ;
        RECT 83.940 161.740 84.270 161.860 ;
        RECT 82.600 161.350 84.500 161.520 ;
        RECT 82.240 161.010 84.160 161.180 ;
        RECT 82.240 160.990 82.560 161.010 ;
        RECT 81.790 160.330 82.120 160.840 ;
        RECT 82.390 160.380 82.560 160.990 ;
        RECT 84.330 160.840 84.500 161.350 ;
        RECT 84.670 161.280 84.850 161.690 ;
        RECT 85.020 161.100 85.190 161.860 ;
        RECT 82.730 160.120 83.060 160.810 ;
        RECT 83.290 160.670 84.500 160.840 ;
        RECT 84.670 160.790 85.190 161.100 ;
        RECT 85.360 161.690 85.780 162.030 ;
        RECT 86.070 161.690 86.480 162.020 ;
        RECT 85.360 160.920 85.550 161.690 ;
        RECT 86.650 161.560 86.820 162.290 ;
        RECT 87.965 162.120 88.135 162.450 ;
        RECT 88.305 162.290 88.635 162.670 ;
        RECT 86.990 161.740 87.340 162.110 ;
        RECT 86.650 161.520 87.070 161.560 ;
        RECT 85.720 161.350 87.070 161.520 ;
        RECT 85.720 161.190 85.970 161.350 ;
        RECT 86.480 160.920 86.730 161.180 ;
        RECT 85.360 160.670 86.730 160.920 ;
        RECT 83.290 160.380 83.530 160.670 ;
        RECT 84.330 160.590 84.500 160.670 ;
        RECT 83.730 160.120 84.150 160.500 ;
        RECT 84.330 160.340 84.960 160.590 ;
        RECT 85.430 160.120 85.760 160.500 ;
        RECT 85.930 160.380 86.100 160.670 ;
        RECT 86.900 160.505 87.070 161.350 ;
        RECT 87.520 161.180 87.740 162.050 ;
        RECT 87.965 161.930 88.660 162.120 ;
        RECT 87.240 160.800 87.740 161.180 ;
        RECT 87.910 161.130 88.320 161.750 ;
        RECT 88.490 160.960 88.660 161.930 ;
        RECT 87.965 160.790 88.660 160.960 ;
        RECT 86.280 160.120 86.660 160.500 ;
        RECT 86.900 160.335 87.730 160.505 ;
        RECT 87.965 160.290 88.135 160.790 ;
        RECT 88.305 160.120 88.635 160.620 ;
        RECT 88.850 160.290 89.075 162.410 ;
        RECT 89.245 162.290 89.575 162.670 ;
        RECT 89.745 162.120 89.915 162.410 ;
        RECT 89.250 161.950 89.915 162.120 ;
        RECT 90.550 161.960 90.805 162.490 ;
        RECT 90.985 162.210 91.270 162.670 ;
        RECT 89.250 160.960 89.480 161.950 ;
        RECT 89.650 161.130 90.000 161.780 ;
        RECT 90.550 161.100 90.730 161.960 ;
        RECT 91.450 161.760 91.700 162.410 ;
        RECT 90.900 161.430 91.700 161.760 ;
        RECT 89.250 160.790 89.915 160.960 ;
        RECT 89.245 160.120 89.575 160.620 ;
        RECT 89.745 160.290 89.915 160.790 ;
        RECT 90.550 160.630 90.805 161.100 ;
        RECT 90.465 160.460 90.805 160.630 ;
        RECT 90.550 160.430 90.805 160.460 ;
        RECT 90.985 160.120 91.270 160.920 ;
        RECT 91.450 160.840 91.700 161.430 ;
        RECT 91.900 162.075 92.220 162.405 ;
        RECT 92.400 162.190 93.060 162.670 ;
        RECT 93.260 162.280 94.110 162.450 ;
        RECT 91.900 161.180 92.090 162.075 ;
        RECT 92.410 161.750 93.070 162.020 ;
        RECT 92.740 161.690 93.070 161.750 ;
        RECT 92.260 161.520 92.590 161.580 ;
        RECT 93.260 161.520 93.430 162.280 ;
        RECT 94.670 162.210 94.990 162.670 ;
        RECT 95.190 162.030 95.440 162.460 ;
        RECT 95.730 162.230 96.140 162.670 ;
        RECT 96.310 162.290 97.325 162.490 ;
        RECT 93.600 161.860 94.850 162.030 ;
        RECT 93.600 161.740 93.930 161.860 ;
        RECT 92.260 161.350 94.160 161.520 ;
        RECT 91.900 161.010 93.820 161.180 ;
        RECT 91.900 160.990 92.220 161.010 ;
        RECT 91.450 160.330 91.780 160.840 ;
        RECT 92.050 160.380 92.220 160.990 ;
        RECT 93.990 160.840 94.160 161.350 ;
        RECT 94.330 161.280 94.510 161.690 ;
        RECT 94.680 161.100 94.850 161.860 ;
        RECT 92.390 160.120 92.720 160.810 ;
        RECT 92.950 160.670 94.160 160.840 ;
        RECT 94.330 160.790 94.850 161.100 ;
        RECT 95.020 161.690 95.440 162.030 ;
        RECT 95.730 161.690 96.140 162.020 ;
        RECT 95.020 160.920 95.210 161.690 ;
        RECT 96.310 161.560 96.480 162.290 ;
        RECT 97.625 162.120 97.795 162.450 ;
        RECT 97.965 162.290 98.295 162.670 ;
        RECT 96.650 161.740 97.000 162.110 ;
        RECT 96.310 161.520 96.730 161.560 ;
        RECT 95.380 161.350 96.730 161.520 ;
        RECT 95.380 161.190 95.630 161.350 ;
        RECT 96.140 160.920 96.390 161.180 ;
        RECT 95.020 160.670 96.390 160.920 ;
        RECT 92.950 160.380 93.190 160.670 ;
        RECT 93.990 160.590 94.160 160.670 ;
        RECT 93.390 160.120 93.810 160.500 ;
        RECT 93.990 160.340 94.620 160.590 ;
        RECT 95.090 160.120 95.420 160.500 ;
        RECT 95.590 160.380 95.760 160.670 ;
        RECT 96.560 160.505 96.730 161.350 ;
        RECT 97.180 161.180 97.400 162.050 ;
        RECT 97.625 161.930 98.320 162.120 ;
        RECT 96.900 160.800 97.400 161.180 ;
        RECT 97.570 161.130 97.980 161.750 ;
        RECT 98.150 160.960 98.320 161.930 ;
        RECT 97.625 160.790 98.320 160.960 ;
        RECT 95.940 160.120 96.320 160.500 ;
        RECT 96.560 160.335 97.390 160.505 ;
        RECT 97.625 160.290 97.795 160.790 ;
        RECT 97.965 160.120 98.295 160.620 ;
        RECT 98.510 160.290 98.735 162.410 ;
        RECT 98.905 162.290 99.235 162.670 ;
        RECT 99.405 162.120 99.575 162.410 ;
        RECT 98.910 161.950 99.575 162.120 ;
        RECT 98.910 160.960 99.140 161.950 ;
        RECT 99.985 161.870 100.315 162.670 ;
        RECT 100.485 162.020 100.655 162.500 ;
        RECT 100.825 162.190 101.155 162.670 ;
        RECT 101.325 162.020 101.495 162.500 ;
        RECT 101.745 162.190 101.985 162.670 ;
        RECT 102.165 162.020 102.335 162.500 ;
        RECT 100.485 161.850 101.495 162.020 ;
        RECT 101.700 161.850 102.335 162.020 ;
        RECT 102.595 161.945 102.885 162.670 ;
        RECT 103.330 161.860 103.575 162.465 ;
        RECT 103.795 162.135 104.305 162.670 ;
        RECT 99.310 161.130 99.660 161.780 ;
        RECT 100.485 161.310 100.980 161.850 ;
        RECT 101.700 161.680 101.870 161.850 ;
        RECT 103.055 161.690 104.285 161.860 ;
        RECT 101.370 161.510 101.870 161.680 ;
        RECT 98.910 160.790 99.575 160.960 ;
        RECT 98.905 160.120 99.235 160.620 ;
        RECT 99.405 160.290 99.575 160.790 ;
        RECT 99.985 160.120 100.315 161.270 ;
        RECT 100.485 161.140 101.495 161.310 ;
        RECT 100.485 160.290 100.655 161.140 ;
        RECT 100.825 160.120 101.155 160.920 ;
        RECT 101.325 160.290 101.495 161.140 ;
        RECT 101.700 161.270 101.870 161.510 ;
        RECT 102.040 161.440 102.420 161.680 ;
        RECT 101.700 161.100 102.415 161.270 ;
        RECT 101.675 160.120 101.915 160.920 ;
        RECT 102.085 160.290 102.415 161.100 ;
        RECT 102.595 160.120 102.885 161.285 ;
        RECT 103.055 160.880 103.395 161.690 ;
        RECT 103.565 161.125 104.315 161.315 ;
        RECT 103.055 160.470 103.570 160.880 ;
        RECT 103.805 160.120 103.975 160.880 ;
        RECT 104.145 160.460 104.315 161.125 ;
        RECT 104.485 161.140 104.675 162.500 ;
        RECT 104.845 161.990 105.120 162.500 ;
        RECT 105.310 162.135 105.840 162.500 ;
        RECT 106.265 162.270 106.595 162.670 ;
        RECT 105.665 162.100 105.840 162.135 ;
        RECT 104.845 161.820 105.125 161.990 ;
        RECT 104.845 161.340 105.120 161.820 ;
        RECT 105.325 161.140 105.495 161.940 ;
        RECT 104.485 160.970 105.495 161.140 ;
        RECT 105.665 161.930 106.595 162.100 ;
        RECT 106.765 161.930 107.020 162.500 ;
        RECT 105.665 160.800 105.835 161.930 ;
        RECT 106.425 161.760 106.595 161.930 ;
        RECT 104.710 160.630 105.835 160.800 ;
        RECT 106.005 161.430 106.200 161.760 ;
        RECT 106.425 161.430 106.680 161.760 ;
        RECT 106.005 160.460 106.175 161.430 ;
        RECT 106.850 161.260 107.020 161.930 ;
        RECT 104.145 160.290 106.175 160.460 ;
        RECT 106.345 160.120 106.515 161.260 ;
        RECT 106.685 160.290 107.020 161.260 ;
        RECT 107.195 161.930 107.580 162.500 ;
        RECT 107.750 162.210 108.075 162.670 ;
        RECT 108.595 162.040 108.875 162.500 ;
        RECT 107.195 161.260 107.475 161.930 ;
        RECT 107.750 161.870 108.875 162.040 ;
        RECT 107.750 161.760 108.200 161.870 ;
        RECT 107.645 161.430 108.200 161.760 ;
        RECT 109.065 161.700 109.465 162.500 ;
        RECT 109.865 162.210 110.135 162.670 ;
        RECT 110.305 162.040 110.590 162.500 ;
        RECT 107.195 160.290 107.580 161.260 ;
        RECT 107.750 160.970 108.200 161.430 ;
        RECT 108.370 161.140 109.465 161.700 ;
        RECT 107.750 160.750 108.875 160.970 ;
        RECT 107.750 160.120 108.075 160.580 ;
        RECT 108.595 160.290 108.875 160.750 ;
        RECT 109.065 160.290 109.465 161.140 ;
        RECT 109.635 161.870 110.590 162.040 ;
        RECT 110.990 162.040 111.275 162.500 ;
        RECT 111.445 162.210 111.715 162.670 ;
        RECT 110.990 161.870 111.945 162.040 ;
        RECT 109.635 160.970 109.845 161.870 ;
        RECT 110.015 161.140 110.705 161.700 ;
        RECT 110.875 161.140 111.565 161.700 ;
        RECT 111.735 160.970 111.945 161.870 ;
        RECT 109.635 160.750 110.590 160.970 ;
        RECT 109.865 160.120 110.135 160.580 ;
        RECT 110.305 160.290 110.590 160.750 ;
        RECT 110.990 160.750 111.945 160.970 ;
        RECT 112.115 161.700 112.515 162.500 ;
        RECT 112.705 162.040 112.985 162.500 ;
        RECT 113.505 162.210 113.830 162.670 ;
        RECT 112.705 161.870 113.830 162.040 ;
        RECT 114.000 161.930 114.385 162.500 ;
        RECT 113.380 161.760 113.830 161.870 ;
        RECT 112.115 161.140 113.210 161.700 ;
        RECT 113.380 161.430 113.935 161.760 ;
        RECT 110.990 160.290 111.275 160.750 ;
        RECT 111.445 160.120 111.715 160.580 ;
        RECT 112.115 160.290 112.515 161.140 ;
        RECT 113.380 160.970 113.830 161.430 ;
        RECT 114.105 161.260 114.385 161.930 ;
        RECT 114.555 161.920 115.765 162.670 ;
        RECT 112.705 160.750 113.830 160.970 ;
        RECT 112.705 160.290 112.985 160.750 ;
        RECT 113.505 160.120 113.830 160.580 ;
        RECT 114.000 160.290 114.385 161.260 ;
        RECT 114.555 161.210 115.075 161.750 ;
        RECT 115.245 161.380 115.765 161.920 ;
        RECT 114.555 160.120 115.765 161.210 ;
        RECT 10.510 159.950 115.850 160.120 ;
        RECT 10.595 158.860 11.805 159.950 ;
        RECT 10.595 158.150 11.115 158.690 ;
        RECT 11.285 158.320 11.805 158.860 ;
        RECT 12.435 158.785 12.725 159.950 ;
        RECT 13.270 159.610 13.525 159.640 ;
        RECT 13.185 159.440 13.525 159.610 ;
        RECT 13.270 158.970 13.525 159.440 ;
        RECT 13.705 159.150 13.990 159.950 ;
        RECT 14.170 159.230 14.500 159.740 ;
        RECT 10.595 157.400 11.805 158.150 ;
        RECT 12.435 157.400 12.725 158.125 ;
        RECT 13.270 158.110 13.450 158.970 ;
        RECT 14.170 158.640 14.420 159.230 ;
        RECT 14.770 159.080 14.940 159.690 ;
        RECT 15.110 159.260 15.440 159.950 ;
        RECT 15.670 159.400 15.910 159.690 ;
        RECT 16.110 159.570 16.530 159.950 ;
        RECT 16.710 159.480 17.340 159.730 ;
        RECT 17.810 159.570 18.140 159.950 ;
        RECT 16.710 159.400 16.880 159.480 ;
        RECT 18.310 159.400 18.480 159.690 ;
        RECT 18.660 159.570 19.040 159.950 ;
        RECT 19.280 159.565 20.110 159.735 ;
        RECT 15.670 159.230 16.880 159.400 ;
        RECT 13.620 158.310 14.420 158.640 ;
        RECT 13.270 157.580 13.525 158.110 ;
        RECT 13.705 157.400 13.990 157.860 ;
        RECT 14.170 157.660 14.420 158.310 ;
        RECT 14.620 159.060 14.940 159.080 ;
        RECT 14.620 158.890 16.540 159.060 ;
        RECT 14.620 157.995 14.810 158.890 ;
        RECT 16.710 158.720 16.880 159.230 ;
        RECT 17.050 158.970 17.570 159.280 ;
        RECT 14.980 158.550 16.880 158.720 ;
        RECT 14.980 158.490 15.310 158.550 ;
        RECT 15.460 158.320 15.790 158.380 ;
        RECT 15.130 158.050 15.790 158.320 ;
        RECT 14.620 157.665 14.940 157.995 ;
        RECT 15.120 157.400 15.780 157.880 ;
        RECT 15.980 157.790 16.150 158.550 ;
        RECT 17.050 158.380 17.230 158.790 ;
        RECT 16.320 158.210 16.650 158.330 ;
        RECT 17.400 158.210 17.570 158.970 ;
        RECT 16.320 158.040 17.570 158.210 ;
        RECT 17.740 159.150 19.110 159.400 ;
        RECT 17.740 158.380 17.930 159.150 ;
        RECT 18.860 158.890 19.110 159.150 ;
        RECT 18.100 158.720 18.350 158.880 ;
        RECT 19.280 158.720 19.450 159.565 ;
        RECT 20.345 159.280 20.515 159.780 ;
        RECT 20.685 159.450 21.015 159.950 ;
        RECT 19.620 158.890 20.120 159.270 ;
        RECT 20.345 159.110 21.040 159.280 ;
        RECT 18.100 158.550 19.450 158.720 ;
        RECT 19.030 158.510 19.450 158.550 ;
        RECT 17.740 158.040 18.160 158.380 ;
        RECT 18.450 158.050 18.860 158.380 ;
        RECT 15.980 157.620 16.830 157.790 ;
        RECT 17.390 157.400 17.710 157.860 ;
        RECT 17.910 157.610 18.160 158.040 ;
        RECT 18.450 157.400 18.860 157.840 ;
        RECT 19.030 157.780 19.200 158.510 ;
        RECT 19.370 157.960 19.720 158.330 ;
        RECT 19.900 158.020 20.120 158.890 ;
        RECT 20.290 158.320 20.700 158.940 ;
        RECT 20.870 158.140 21.040 159.110 ;
        RECT 20.345 157.950 21.040 158.140 ;
        RECT 19.030 157.580 20.045 157.780 ;
        RECT 20.345 157.620 20.515 157.950 ;
        RECT 20.685 157.400 21.015 157.780 ;
        RECT 21.230 157.660 21.455 159.780 ;
        RECT 21.625 159.450 21.955 159.950 ;
        RECT 22.125 159.280 22.295 159.780 ;
        RECT 21.630 159.110 22.295 159.280 ;
        RECT 21.630 158.120 21.860 159.110 ;
        RECT 22.030 158.290 22.380 158.940 ;
        RECT 22.555 158.875 22.825 159.780 ;
        RECT 22.995 159.190 23.325 159.950 ;
        RECT 23.505 159.020 23.675 159.780 ;
        RECT 21.630 157.950 22.295 158.120 ;
        RECT 21.625 157.400 21.955 157.780 ;
        RECT 22.125 157.660 22.295 157.950 ;
        RECT 22.555 158.075 22.725 158.875 ;
        RECT 23.010 158.850 23.675 159.020 ;
        RECT 23.935 158.860 25.145 159.950 ;
        RECT 25.430 159.320 25.715 159.780 ;
        RECT 25.885 159.490 26.155 159.950 ;
        RECT 25.430 159.100 26.385 159.320 ;
        RECT 23.010 158.705 23.180 158.850 ;
        RECT 22.895 158.375 23.180 158.705 ;
        RECT 23.010 158.120 23.180 158.375 ;
        RECT 23.415 158.300 23.745 158.670 ;
        RECT 23.935 158.320 24.455 158.860 ;
        RECT 24.625 158.150 25.145 158.690 ;
        RECT 25.315 158.370 26.005 158.930 ;
        RECT 26.175 158.200 26.385 159.100 ;
        RECT 22.555 157.570 22.815 158.075 ;
        RECT 23.010 157.950 23.675 158.120 ;
        RECT 22.995 157.400 23.325 157.780 ;
        RECT 23.505 157.570 23.675 157.950 ;
        RECT 23.935 157.400 25.145 158.150 ;
        RECT 25.430 158.030 26.385 158.200 ;
        RECT 26.555 158.930 26.955 159.780 ;
        RECT 27.145 159.320 27.425 159.780 ;
        RECT 27.945 159.490 28.270 159.950 ;
        RECT 27.145 159.100 28.270 159.320 ;
        RECT 26.555 158.370 27.650 158.930 ;
        RECT 27.820 158.640 28.270 159.100 ;
        RECT 28.440 158.810 28.825 159.780 ;
        RECT 25.430 157.570 25.715 158.030 ;
        RECT 25.885 157.400 26.155 157.860 ;
        RECT 26.555 157.570 26.955 158.370 ;
        RECT 27.820 158.310 28.375 158.640 ;
        RECT 27.820 158.200 28.270 158.310 ;
        RECT 27.145 158.030 28.270 158.200 ;
        RECT 28.545 158.140 28.825 158.810 ;
        RECT 27.145 157.570 27.425 158.030 ;
        RECT 27.945 157.400 28.270 157.860 ;
        RECT 28.440 157.570 28.825 158.140 ;
        RECT 29.000 158.810 29.335 159.780 ;
        RECT 29.505 158.810 29.675 159.950 ;
        RECT 29.845 159.610 31.875 159.780 ;
        RECT 29.000 158.140 29.170 158.810 ;
        RECT 29.845 158.640 30.015 159.610 ;
        RECT 29.340 158.310 29.595 158.640 ;
        RECT 29.820 158.310 30.015 158.640 ;
        RECT 30.185 159.270 31.310 159.440 ;
        RECT 29.425 158.140 29.595 158.310 ;
        RECT 30.185 158.140 30.355 159.270 ;
        RECT 29.000 157.570 29.255 158.140 ;
        RECT 29.425 157.970 30.355 158.140 ;
        RECT 30.525 158.930 31.535 159.100 ;
        RECT 30.525 158.130 30.695 158.930 ;
        RECT 30.900 158.590 31.175 158.730 ;
        RECT 30.895 158.420 31.175 158.590 ;
        RECT 30.180 157.935 30.355 157.970 ;
        RECT 29.425 157.400 29.755 157.800 ;
        RECT 30.180 157.570 30.710 157.935 ;
        RECT 30.900 157.570 31.175 158.420 ;
        RECT 31.345 157.570 31.535 158.930 ;
        RECT 31.705 158.945 31.875 159.610 ;
        RECT 32.045 159.190 32.215 159.950 ;
        RECT 32.450 159.190 32.965 159.600 ;
        RECT 31.705 158.755 32.455 158.945 ;
        RECT 32.625 158.380 32.965 159.190 ;
        RECT 31.735 158.210 32.965 158.380 ;
        RECT 33.135 158.860 34.345 159.950 ;
        RECT 33.135 158.320 33.655 158.860 ;
        RECT 34.515 158.810 34.855 159.780 ;
        RECT 35.025 158.810 35.195 159.950 ;
        RECT 35.465 159.150 35.715 159.950 ;
        RECT 36.360 158.980 36.690 159.780 ;
        RECT 36.990 159.150 37.320 159.950 ;
        RECT 37.490 158.980 37.820 159.780 ;
        RECT 35.385 158.810 37.820 158.980 ;
        RECT 31.715 157.400 32.225 157.935 ;
        RECT 32.445 157.605 32.690 158.210 ;
        RECT 33.825 158.150 34.345 158.690 ;
        RECT 33.135 157.400 34.345 158.150 ;
        RECT 34.515 158.200 34.690 158.810 ;
        RECT 35.385 158.560 35.555 158.810 ;
        RECT 34.860 158.390 35.555 158.560 ;
        RECT 35.730 158.390 36.150 158.590 ;
        RECT 36.320 158.390 36.650 158.590 ;
        RECT 36.820 158.390 37.150 158.590 ;
        RECT 34.515 157.570 34.855 158.200 ;
        RECT 35.025 157.400 35.275 158.200 ;
        RECT 35.465 158.050 36.690 158.220 ;
        RECT 35.465 157.570 35.795 158.050 ;
        RECT 35.965 157.400 36.190 157.860 ;
        RECT 36.360 157.570 36.690 158.050 ;
        RECT 37.320 158.180 37.490 158.810 ;
        RECT 38.195 158.785 38.485 159.950 ;
        RECT 38.655 158.860 39.865 159.950 ;
        RECT 40.240 158.980 40.570 159.780 ;
        RECT 40.740 159.150 41.070 159.950 ;
        RECT 41.370 158.980 41.700 159.780 ;
        RECT 42.345 159.150 42.595 159.950 ;
        RECT 37.675 158.390 38.025 158.640 ;
        RECT 38.655 158.320 39.175 158.860 ;
        RECT 40.240 158.810 42.675 158.980 ;
        RECT 42.865 158.810 43.035 159.950 ;
        RECT 43.205 158.810 43.545 159.780 ;
        RECT 37.320 157.570 37.820 158.180 ;
        RECT 39.345 158.150 39.865 158.690 ;
        RECT 40.035 158.390 40.385 158.640 ;
        RECT 40.570 158.180 40.740 158.810 ;
        RECT 40.910 158.390 41.240 158.590 ;
        RECT 41.410 158.390 41.740 158.590 ;
        RECT 41.910 158.390 42.330 158.590 ;
        RECT 42.505 158.560 42.675 158.810 ;
        RECT 42.505 158.390 43.200 158.560 ;
        RECT 38.195 157.400 38.485 158.125 ;
        RECT 38.655 157.400 39.865 158.150 ;
        RECT 40.240 157.570 40.740 158.180 ;
        RECT 41.370 158.050 42.595 158.220 ;
        RECT 43.370 158.200 43.545 158.810 ;
        RECT 41.370 157.570 41.700 158.050 ;
        RECT 41.870 157.400 42.095 157.860 ;
        RECT 42.265 157.570 42.595 158.050 ;
        RECT 42.785 157.400 43.035 158.200 ;
        RECT 43.205 157.570 43.545 158.200 ;
        RECT 43.715 158.810 44.055 159.780 ;
        RECT 44.225 158.810 44.395 159.950 ;
        RECT 44.665 159.150 44.915 159.950 ;
        RECT 45.560 158.980 45.890 159.780 ;
        RECT 46.190 159.150 46.520 159.950 ;
        RECT 46.690 158.980 47.020 159.780 ;
        RECT 44.585 158.810 47.020 158.980 ;
        RECT 47.770 158.970 48.025 159.640 ;
        RECT 48.205 159.150 48.490 159.950 ;
        RECT 48.670 159.230 49.000 159.740 ;
        RECT 43.715 158.760 43.945 158.810 ;
        RECT 43.715 158.200 43.890 158.760 ;
        RECT 44.585 158.560 44.755 158.810 ;
        RECT 44.060 158.390 44.755 158.560 ;
        RECT 44.930 158.390 45.350 158.590 ;
        RECT 45.520 158.390 45.850 158.590 ;
        RECT 46.020 158.390 46.350 158.590 ;
        RECT 43.715 157.570 44.055 158.200 ;
        RECT 44.225 157.400 44.475 158.200 ;
        RECT 44.665 158.050 45.890 158.220 ;
        RECT 44.665 157.570 44.995 158.050 ;
        RECT 45.165 157.400 45.390 157.860 ;
        RECT 45.560 157.570 45.890 158.050 ;
        RECT 46.520 158.180 46.690 158.810 ;
        RECT 46.875 158.390 47.225 158.640 ;
        RECT 46.520 157.570 47.020 158.180 ;
        RECT 47.770 158.110 47.950 158.970 ;
        RECT 48.670 158.640 48.920 159.230 ;
        RECT 49.270 159.080 49.440 159.690 ;
        RECT 49.610 159.260 49.940 159.950 ;
        RECT 50.170 159.400 50.410 159.690 ;
        RECT 50.610 159.570 51.030 159.950 ;
        RECT 51.210 159.480 51.840 159.730 ;
        RECT 52.310 159.570 52.640 159.950 ;
        RECT 51.210 159.400 51.380 159.480 ;
        RECT 52.810 159.400 52.980 159.690 ;
        RECT 53.160 159.570 53.540 159.950 ;
        RECT 53.780 159.565 54.610 159.735 ;
        RECT 50.170 159.230 51.380 159.400 ;
        RECT 48.120 158.310 48.920 158.640 ;
        RECT 47.770 157.910 48.025 158.110 ;
        RECT 47.685 157.740 48.025 157.910 ;
        RECT 47.770 157.580 48.025 157.740 ;
        RECT 48.205 157.400 48.490 157.860 ;
        RECT 48.670 157.660 48.920 158.310 ;
        RECT 49.120 159.060 49.440 159.080 ;
        RECT 49.120 158.890 51.040 159.060 ;
        RECT 49.120 157.995 49.310 158.890 ;
        RECT 51.210 158.720 51.380 159.230 ;
        RECT 51.550 158.970 52.070 159.280 ;
        RECT 49.480 158.550 51.380 158.720 ;
        RECT 49.480 158.490 49.810 158.550 ;
        RECT 49.960 158.320 50.290 158.380 ;
        RECT 49.630 158.050 50.290 158.320 ;
        RECT 49.120 157.665 49.440 157.995 ;
        RECT 49.620 157.400 50.280 157.880 ;
        RECT 50.480 157.790 50.650 158.550 ;
        RECT 51.550 158.380 51.730 158.790 ;
        RECT 50.820 158.210 51.150 158.330 ;
        RECT 51.900 158.210 52.070 158.970 ;
        RECT 50.820 158.040 52.070 158.210 ;
        RECT 52.240 159.150 53.610 159.400 ;
        RECT 52.240 158.380 52.430 159.150 ;
        RECT 53.360 158.890 53.610 159.150 ;
        RECT 52.600 158.720 52.850 158.880 ;
        RECT 53.780 158.720 53.950 159.565 ;
        RECT 54.845 159.280 55.015 159.780 ;
        RECT 55.185 159.450 55.515 159.950 ;
        RECT 54.120 158.890 54.620 159.270 ;
        RECT 54.845 159.110 55.540 159.280 ;
        RECT 52.600 158.550 53.950 158.720 ;
        RECT 53.530 158.510 53.950 158.550 ;
        RECT 52.240 158.040 52.660 158.380 ;
        RECT 52.950 158.050 53.360 158.380 ;
        RECT 50.480 157.620 51.330 157.790 ;
        RECT 51.890 157.400 52.210 157.860 ;
        RECT 52.410 157.610 52.660 158.040 ;
        RECT 52.950 157.400 53.360 157.840 ;
        RECT 53.530 157.780 53.700 158.510 ;
        RECT 53.870 157.960 54.220 158.330 ;
        RECT 54.400 158.020 54.620 158.890 ;
        RECT 54.790 158.320 55.200 158.940 ;
        RECT 55.370 158.140 55.540 159.110 ;
        RECT 54.845 157.950 55.540 158.140 ;
        RECT 53.530 157.580 54.545 157.780 ;
        RECT 54.845 157.620 55.015 157.950 ;
        RECT 55.185 157.400 55.515 157.780 ;
        RECT 55.730 157.660 55.955 159.780 ;
        RECT 56.125 159.450 56.455 159.950 ;
        RECT 56.625 159.280 56.795 159.780 ;
        RECT 56.130 159.110 56.795 159.280 ;
        RECT 56.130 158.120 56.360 159.110 ;
        RECT 56.530 158.290 56.880 158.940 ;
        RECT 57.205 158.800 57.535 159.950 ;
        RECT 57.705 158.930 57.875 159.780 ;
        RECT 58.045 159.150 58.375 159.950 ;
        RECT 58.545 158.930 58.715 159.780 ;
        RECT 58.895 159.150 59.135 159.950 ;
        RECT 59.305 158.970 59.635 159.780 ;
        RECT 57.705 158.760 58.715 158.930 ;
        RECT 58.920 158.800 59.635 158.970 ;
        RECT 60.275 158.860 61.945 159.950 ;
        RECT 57.705 158.220 58.200 158.760 ;
        RECT 58.920 158.560 59.090 158.800 ;
        RECT 58.590 158.390 59.090 158.560 ;
        RECT 59.260 158.390 59.640 158.630 ;
        RECT 58.920 158.220 59.090 158.390 ;
        RECT 60.275 158.340 61.025 158.860 ;
        RECT 62.120 158.800 62.380 159.950 ;
        RECT 62.555 158.875 62.810 159.780 ;
        RECT 62.980 159.190 63.310 159.950 ;
        RECT 63.525 159.020 63.695 159.780 ;
        RECT 56.130 157.950 56.795 158.120 ;
        RECT 56.125 157.400 56.455 157.780 ;
        RECT 56.625 157.660 56.795 157.950 ;
        RECT 57.205 157.400 57.535 158.200 ;
        RECT 57.705 158.050 58.715 158.220 ;
        RECT 58.920 158.050 59.555 158.220 ;
        RECT 61.195 158.170 61.945 158.690 ;
        RECT 57.705 157.570 57.875 158.050 ;
        RECT 58.045 157.400 58.375 157.880 ;
        RECT 58.545 157.570 58.715 158.050 ;
        RECT 58.965 157.400 59.205 157.880 ;
        RECT 59.385 157.570 59.555 158.050 ;
        RECT 60.275 157.400 61.945 158.170 ;
        RECT 62.120 157.400 62.380 158.240 ;
        RECT 62.555 158.145 62.725 158.875 ;
        RECT 62.980 158.850 63.695 159.020 ;
        RECT 62.980 158.640 63.150 158.850 ;
        RECT 63.955 158.785 64.245 159.950 ;
        RECT 64.875 158.860 67.465 159.950 ;
        RECT 62.895 158.310 63.150 158.640 ;
        RECT 62.555 157.570 62.810 158.145 ;
        RECT 62.980 158.120 63.150 158.310 ;
        RECT 63.430 158.300 63.785 158.670 ;
        RECT 64.875 158.340 66.085 158.860 ;
        RECT 67.635 158.810 67.975 159.780 ;
        RECT 68.145 158.810 68.315 159.950 ;
        RECT 68.585 159.150 68.835 159.950 ;
        RECT 69.480 158.980 69.810 159.780 ;
        RECT 70.110 159.150 70.440 159.950 ;
        RECT 70.610 158.980 70.940 159.780 ;
        RECT 68.505 158.810 70.940 158.980 ;
        RECT 71.775 158.860 73.445 159.950 ;
        RECT 73.990 158.970 74.245 159.640 ;
        RECT 74.425 159.150 74.710 159.950 ;
        RECT 74.890 159.230 75.220 159.740 ;
        RECT 66.255 158.170 67.465 158.690 ;
        RECT 62.980 157.950 63.695 158.120 ;
        RECT 62.980 157.400 63.310 157.780 ;
        RECT 63.525 157.570 63.695 157.950 ;
        RECT 63.955 157.400 64.245 158.125 ;
        RECT 64.875 157.400 67.465 158.170 ;
        RECT 67.635 158.200 67.810 158.810 ;
        RECT 68.505 158.560 68.675 158.810 ;
        RECT 67.980 158.390 68.675 158.560 ;
        RECT 68.850 158.390 69.270 158.590 ;
        RECT 69.440 158.390 69.770 158.590 ;
        RECT 69.940 158.390 70.270 158.590 ;
        RECT 67.635 157.570 67.975 158.200 ;
        RECT 68.145 157.400 68.395 158.200 ;
        RECT 68.585 158.050 69.810 158.220 ;
        RECT 68.585 157.570 68.915 158.050 ;
        RECT 69.085 157.400 69.310 157.860 ;
        RECT 69.480 157.570 69.810 158.050 ;
        RECT 70.440 158.180 70.610 158.810 ;
        RECT 70.795 158.390 71.145 158.640 ;
        RECT 71.775 158.340 72.525 158.860 ;
        RECT 70.440 157.570 70.940 158.180 ;
        RECT 72.695 158.170 73.445 158.690 ;
        RECT 71.775 157.400 73.445 158.170 ;
        RECT 73.990 158.110 74.170 158.970 ;
        RECT 74.890 158.640 75.140 159.230 ;
        RECT 75.490 159.080 75.660 159.690 ;
        RECT 75.830 159.260 76.160 159.950 ;
        RECT 76.390 159.400 76.630 159.690 ;
        RECT 76.830 159.570 77.250 159.950 ;
        RECT 77.430 159.480 78.060 159.730 ;
        RECT 78.530 159.570 78.860 159.950 ;
        RECT 77.430 159.400 77.600 159.480 ;
        RECT 79.030 159.400 79.200 159.690 ;
        RECT 79.380 159.570 79.760 159.950 ;
        RECT 80.000 159.565 80.830 159.735 ;
        RECT 76.390 159.230 77.600 159.400 ;
        RECT 74.340 158.310 75.140 158.640 ;
        RECT 73.990 157.910 74.245 158.110 ;
        RECT 73.905 157.740 74.245 157.910 ;
        RECT 73.990 157.580 74.245 157.740 ;
        RECT 74.425 157.400 74.710 157.860 ;
        RECT 74.890 157.660 75.140 158.310 ;
        RECT 75.340 159.060 75.660 159.080 ;
        RECT 75.340 158.890 77.260 159.060 ;
        RECT 75.340 157.995 75.530 158.890 ;
        RECT 77.430 158.720 77.600 159.230 ;
        RECT 77.770 158.970 78.290 159.280 ;
        RECT 75.700 158.550 77.600 158.720 ;
        RECT 75.700 158.490 76.030 158.550 ;
        RECT 76.180 158.320 76.510 158.380 ;
        RECT 75.850 158.050 76.510 158.320 ;
        RECT 75.340 157.665 75.660 157.995 ;
        RECT 75.840 157.400 76.500 157.880 ;
        RECT 76.700 157.790 76.870 158.550 ;
        RECT 77.770 158.380 77.950 158.790 ;
        RECT 77.040 158.210 77.370 158.330 ;
        RECT 78.120 158.210 78.290 158.970 ;
        RECT 77.040 158.040 78.290 158.210 ;
        RECT 78.460 159.150 79.830 159.400 ;
        RECT 78.460 158.380 78.650 159.150 ;
        RECT 79.580 158.890 79.830 159.150 ;
        RECT 78.820 158.720 79.070 158.880 ;
        RECT 80.000 158.720 80.170 159.565 ;
        RECT 81.065 159.280 81.235 159.780 ;
        RECT 81.405 159.450 81.735 159.950 ;
        RECT 80.340 158.890 80.840 159.270 ;
        RECT 81.065 159.110 81.760 159.280 ;
        RECT 78.820 158.550 80.170 158.720 ;
        RECT 79.750 158.510 80.170 158.550 ;
        RECT 78.460 158.040 78.880 158.380 ;
        RECT 79.170 158.050 79.580 158.380 ;
        RECT 76.700 157.620 77.550 157.790 ;
        RECT 78.110 157.400 78.430 157.860 ;
        RECT 78.630 157.610 78.880 158.040 ;
        RECT 79.170 157.400 79.580 157.840 ;
        RECT 79.750 157.780 79.920 158.510 ;
        RECT 80.090 157.960 80.440 158.330 ;
        RECT 80.620 158.020 80.840 158.890 ;
        RECT 81.010 158.320 81.420 158.940 ;
        RECT 81.590 158.140 81.760 159.110 ;
        RECT 81.065 157.950 81.760 158.140 ;
        RECT 79.750 157.580 80.765 157.780 ;
        RECT 81.065 157.620 81.235 157.950 ;
        RECT 81.405 157.400 81.735 157.780 ;
        RECT 81.950 157.660 82.175 159.780 ;
        RECT 82.345 159.450 82.675 159.950 ;
        RECT 82.845 159.280 83.015 159.780 ;
        RECT 82.350 159.110 83.015 159.280 ;
        RECT 82.350 158.120 82.580 159.110 ;
        RECT 82.750 158.290 83.100 158.940 ;
        RECT 84.255 158.810 84.465 159.950 ;
        RECT 84.635 158.800 84.965 159.780 ;
        RECT 85.135 158.810 85.365 159.950 ;
        RECT 86.240 158.980 86.570 159.780 ;
        RECT 86.740 159.150 87.070 159.950 ;
        RECT 87.370 158.980 87.700 159.780 ;
        RECT 88.345 159.150 88.595 159.950 ;
        RECT 86.240 158.810 88.675 158.980 ;
        RECT 88.865 158.810 89.035 159.950 ;
        RECT 89.205 158.810 89.545 159.780 ;
        RECT 82.350 157.950 83.015 158.120 ;
        RECT 82.345 157.400 82.675 157.780 ;
        RECT 82.845 157.660 83.015 157.950 ;
        RECT 84.255 157.400 84.465 158.220 ;
        RECT 84.635 158.200 84.885 158.800 ;
        RECT 85.055 158.390 85.385 158.640 ;
        RECT 86.035 158.390 86.385 158.640 ;
        RECT 84.635 157.570 84.965 158.200 ;
        RECT 85.135 157.400 85.365 158.220 ;
        RECT 86.570 158.180 86.740 158.810 ;
        RECT 86.910 158.390 87.240 158.590 ;
        RECT 87.410 158.390 87.740 158.590 ;
        RECT 87.910 158.390 88.330 158.590 ;
        RECT 88.505 158.560 88.675 158.810 ;
        RECT 88.505 158.390 89.200 158.560 ;
        RECT 86.240 157.570 86.740 158.180 ;
        RECT 87.370 158.050 88.595 158.220 ;
        RECT 89.370 158.200 89.545 158.810 ;
        RECT 89.715 158.785 90.005 159.950 ;
        RECT 90.175 158.875 90.445 159.780 ;
        RECT 90.615 159.190 90.945 159.950 ;
        RECT 91.125 159.020 91.295 159.780 ;
        RECT 87.370 157.570 87.700 158.050 ;
        RECT 87.870 157.400 88.095 157.860 ;
        RECT 88.265 157.570 88.595 158.050 ;
        RECT 88.785 157.400 89.035 158.200 ;
        RECT 89.205 157.570 89.545 158.200 ;
        RECT 89.715 157.400 90.005 158.125 ;
        RECT 90.175 158.075 90.345 158.875 ;
        RECT 90.630 158.850 91.295 159.020 ;
        RECT 90.630 158.705 90.800 158.850 ;
        RECT 90.515 158.375 90.800 158.705 ;
        RECT 92.475 158.810 92.860 159.780 ;
        RECT 93.030 159.490 93.355 159.950 ;
        RECT 93.875 159.320 94.155 159.780 ;
        RECT 93.030 159.100 94.155 159.320 ;
        RECT 90.630 158.120 90.800 158.375 ;
        RECT 91.035 158.300 91.365 158.670 ;
        RECT 92.475 158.140 92.755 158.810 ;
        RECT 93.030 158.640 93.480 159.100 ;
        RECT 94.345 158.930 94.745 159.780 ;
        RECT 95.145 159.490 95.415 159.950 ;
        RECT 95.585 159.320 95.870 159.780 ;
        RECT 92.925 158.310 93.480 158.640 ;
        RECT 93.650 158.370 94.745 158.930 ;
        RECT 93.030 158.200 93.480 158.310 ;
        RECT 90.175 157.570 90.435 158.075 ;
        RECT 90.630 157.950 91.295 158.120 ;
        RECT 90.615 157.400 90.945 157.780 ;
        RECT 91.125 157.570 91.295 157.950 ;
        RECT 92.475 157.570 92.860 158.140 ;
        RECT 93.030 158.030 94.155 158.200 ;
        RECT 93.030 157.400 93.355 157.860 ;
        RECT 93.875 157.570 94.155 158.030 ;
        RECT 94.345 157.570 94.745 158.370 ;
        RECT 94.915 159.100 95.870 159.320 ;
        RECT 94.915 158.200 95.125 159.100 ;
        RECT 96.245 159.020 96.415 159.780 ;
        RECT 96.595 159.190 96.925 159.950 ;
        RECT 95.295 158.370 95.985 158.930 ;
        RECT 96.245 158.850 96.910 159.020 ;
        RECT 97.095 158.875 97.365 159.780 ;
        RECT 96.740 158.705 96.910 158.850 ;
        RECT 96.175 158.300 96.505 158.670 ;
        RECT 96.740 158.375 97.025 158.705 ;
        RECT 94.915 158.030 95.870 158.200 ;
        RECT 96.740 158.120 96.910 158.375 ;
        RECT 95.145 157.400 95.415 157.860 ;
        RECT 95.585 157.570 95.870 158.030 ;
        RECT 96.245 157.950 96.910 158.120 ;
        RECT 97.195 158.075 97.365 158.875 ;
        RECT 97.740 158.980 98.070 159.780 ;
        RECT 98.240 159.150 98.570 159.950 ;
        RECT 98.870 158.980 99.200 159.780 ;
        RECT 99.845 159.150 100.095 159.950 ;
        RECT 97.740 158.810 100.175 158.980 ;
        RECT 100.365 158.810 100.535 159.950 ;
        RECT 100.705 158.810 101.045 159.780 ;
        RECT 97.535 158.390 97.885 158.640 ;
        RECT 98.070 158.180 98.240 158.810 ;
        RECT 98.410 158.390 98.740 158.590 ;
        RECT 98.910 158.390 99.240 158.590 ;
        RECT 99.410 158.390 99.830 158.590 ;
        RECT 100.005 158.560 100.175 158.810 ;
        RECT 100.005 158.390 100.700 158.560 ;
        RECT 96.245 157.570 96.415 157.950 ;
        RECT 96.595 157.400 96.925 157.780 ;
        RECT 97.105 157.570 97.365 158.075 ;
        RECT 97.740 157.570 98.240 158.180 ;
        RECT 98.870 158.050 100.095 158.220 ;
        RECT 100.870 158.200 101.045 158.810 ;
        RECT 101.675 158.860 103.345 159.950 ;
        RECT 103.515 159.190 104.030 159.600 ;
        RECT 104.265 159.190 104.435 159.950 ;
        RECT 104.605 159.610 106.635 159.780 ;
        RECT 101.675 158.340 102.425 158.860 ;
        RECT 98.870 157.570 99.200 158.050 ;
        RECT 99.370 157.400 99.595 157.860 ;
        RECT 99.765 157.570 100.095 158.050 ;
        RECT 100.285 157.400 100.535 158.200 ;
        RECT 100.705 157.570 101.045 158.200 ;
        RECT 102.595 158.170 103.345 158.690 ;
        RECT 103.515 158.380 103.855 159.190 ;
        RECT 104.605 158.945 104.775 159.610 ;
        RECT 105.170 159.270 106.295 159.440 ;
        RECT 104.025 158.755 104.775 158.945 ;
        RECT 104.945 158.930 105.955 159.100 ;
        RECT 103.515 158.210 104.745 158.380 ;
        RECT 101.675 157.400 103.345 158.170 ;
        RECT 103.790 157.605 104.035 158.210 ;
        RECT 104.255 157.400 104.765 157.935 ;
        RECT 104.945 157.570 105.135 158.930 ;
        RECT 105.305 158.590 105.580 158.730 ;
        RECT 105.305 158.420 105.585 158.590 ;
        RECT 105.305 157.570 105.580 158.420 ;
        RECT 105.785 158.130 105.955 158.930 ;
        RECT 106.125 158.140 106.295 159.270 ;
        RECT 106.465 158.640 106.635 159.610 ;
        RECT 106.805 158.810 106.975 159.950 ;
        RECT 107.145 158.810 107.480 159.780 ;
        RECT 106.465 158.310 106.660 158.640 ;
        RECT 106.885 158.310 107.140 158.640 ;
        RECT 106.885 158.140 107.055 158.310 ;
        RECT 107.310 158.140 107.480 158.810 ;
        RECT 108.115 158.860 109.785 159.950 ;
        RECT 110.045 159.020 110.215 159.780 ;
        RECT 110.395 159.190 110.725 159.950 ;
        RECT 108.115 158.340 108.865 158.860 ;
        RECT 110.045 158.850 110.710 159.020 ;
        RECT 110.895 158.875 111.165 159.780 ;
        RECT 110.540 158.705 110.710 158.850 ;
        RECT 109.035 158.170 109.785 158.690 ;
        RECT 109.975 158.300 110.305 158.670 ;
        RECT 110.540 158.375 110.825 158.705 ;
        RECT 106.125 157.970 107.055 158.140 ;
        RECT 106.125 157.935 106.300 157.970 ;
        RECT 105.770 157.570 106.300 157.935 ;
        RECT 106.725 157.400 107.055 157.800 ;
        RECT 107.225 157.570 107.480 158.140 ;
        RECT 108.115 157.400 109.785 158.170 ;
        RECT 110.540 158.120 110.710 158.375 ;
        RECT 110.045 157.950 110.710 158.120 ;
        RECT 110.995 158.075 111.165 158.875 ;
        RECT 111.795 158.860 114.385 159.950 ;
        RECT 114.555 158.860 115.765 159.950 ;
        RECT 111.795 158.340 113.005 158.860 ;
        RECT 113.175 158.170 114.385 158.690 ;
        RECT 114.555 158.320 115.075 158.860 ;
        RECT 110.045 157.570 110.215 157.950 ;
        RECT 110.395 157.400 110.725 157.780 ;
        RECT 110.905 157.570 111.165 158.075 ;
        RECT 111.795 157.400 114.385 158.170 ;
        RECT 115.245 158.150 115.765 158.690 ;
        RECT 114.555 157.400 115.765 158.150 ;
        RECT 10.510 157.230 115.850 157.400 ;
        RECT 10.595 156.480 11.805 157.230 ;
        RECT 10.595 155.940 11.115 156.480 ;
        RECT 12.435 156.460 15.025 157.230 ;
        RECT 11.285 155.770 11.805 156.310 ;
        RECT 10.595 154.680 11.805 155.770 ;
        RECT 12.435 155.770 13.645 156.290 ;
        RECT 13.815 155.940 15.025 156.460 ;
        RECT 15.235 156.410 15.465 157.230 ;
        RECT 15.635 156.430 15.965 157.060 ;
        RECT 15.215 155.990 15.545 156.240 ;
        RECT 15.715 155.830 15.965 156.430 ;
        RECT 16.135 156.410 16.345 157.230 ;
        RECT 16.850 156.420 17.095 157.025 ;
        RECT 17.315 156.695 17.825 157.230 ;
        RECT 12.435 154.680 15.025 155.770 ;
        RECT 15.235 154.680 15.465 155.820 ;
        RECT 15.635 154.850 15.965 155.830 ;
        RECT 16.575 156.250 17.805 156.420 ;
        RECT 16.135 154.680 16.345 155.820 ;
        RECT 16.575 155.440 16.915 156.250 ;
        RECT 17.085 155.685 17.835 155.875 ;
        RECT 16.575 155.030 17.090 155.440 ;
        RECT 17.325 154.680 17.495 155.440 ;
        RECT 17.665 155.020 17.835 155.685 ;
        RECT 18.005 155.700 18.195 157.060 ;
        RECT 18.365 156.210 18.640 157.060 ;
        RECT 18.830 156.695 19.360 157.060 ;
        RECT 19.785 156.830 20.115 157.230 ;
        RECT 19.185 156.660 19.360 156.695 ;
        RECT 18.365 156.040 18.645 156.210 ;
        RECT 18.365 155.900 18.640 156.040 ;
        RECT 18.845 155.700 19.015 156.500 ;
        RECT 18.005 155.530 19.015 155.700 ;
        RECT 19.185 156.490 20.115 156.660 ;
        RECT 20.285 156.490 20.540 157.060 ;
        RECT 19.185 155.360 19.355 156.490 ;
        RECT 19.945 156.320 20.115 156.490 ;
        RECT 18.230 155.190 19.355 155.360 ;
        RECT 19.525 155.990 19.720 156.320 ;
        RECT 19.945 155.990 20.200 156.320 ;
        RECT 19.525 155.020 19.695 155.990 ;
        RECT 20.370 155.820 20.540 156.490 ;
        RECT 17.665 154.850 19.695 155.020 ;
        RECT 19.865 154.680 20.035 155.820 ;
        RECT 20.205 154.850 20.540 155.820 ;
        RECT 21.635 156.490 22.020 157.060 ;
        RECT 22.190 156.770 22.515 157.230 ;
        RECT 23.035 156.600 23.315 157.060 ;
        RECT 21.635 155.820 21.915 156.490 ;
        RECT 22.190 156.430 23.315 156.600 ;
        RECT 22.190 156.320 22.640 156.430 ;
        RECT 22.085 155.990 22.640 156.320 ;
        RECT 23.505 156.260 23.905 157.060 ;
        RECT 24.305 156.770 24.575 157.230 ;
        RECT 24.745 156.600 25.030 157.060 ;
        RECT 21.635 154.850 22.020 155.820 ;
        RECT 22.190 155.530 22.640 155.990 ;
        RECT 22.810 155.700 23.905 156.260 ;
        RECT 22.190 155.310 23.315 155.530 ;
        RECT 22.190 154.680 22.515 155.140 ;
        RECT 23.035 154.850 23.315 155.310 ;
        RECT 23.505 154.850 23.905 155.700 ;
        RECT 24.075 156.430 25.030 156.600 ;
        RECT 25.315 156.505 25.605 157.230 ;
        RECT 25.890 156.600 26.175 157.060 ;
        RECT 26.345 156.770 26.615 157.230 ;
        RECT 25.890 156.430 26.845 156.600 ;
        RECT 24.075 155.530 24.285 156.430 ;
        RECT 24.455 155.700 25.145 156.260 ;
        RECT 24.075 155.310 25.030 155.530 ;
        RECT 24.305 154.680 24.575 155.140 ;
        RECT 24.745 154.850 25.030 155.310 ;
        RECT 25.315 154.680 25.605 155.845 ;
        RECT 25.775 155.700 26.465 156.260 ;
        RECT 26.635 155.530 26.845 156.430 ;
        RECT 25.890 155.310 26.845 155.530 ;
        RECT 27.015 156.260 27.415 157.060 ;
        RECT 27.605 156.600 27.885 157.060 ;
        RECT 28.405 156.770 28.730 157.230 ;
        RECT 27.605 156.430 28.730 156.600 ;
        RECT 28.900 156.490 29.285 157.060 ;
        RECT 28.280 156.320 28.730 156.430 ;
        RECT 27.015 155.700 28.110 156.260 ;
        RECT 28.280 155.990 28.835 156.320 ;
        RECT 25.890 154.850 26.175 155.310 ;
        RECT 26.345 154.680 26.615 155.140 ;
        RECT 27.015 154.850 27.415 155.700 ;
        RECT 28.280 155.530 28.730 155.990 ;
        RECT 29.005 155.820 29.285 156.490 ;
        RECT 27.605 155.310 28.730 155.530 ;
        RECT 27.605 154.850 27.885 155.310 ;
        RECT 28.405 154.680 28.730 155.140 ;
        RECT 28.900 154.850 29.285 155.820 ;
        RECT 29.455 156.430 29.795 157.060 ;
        RECT 29.965 156.430 30.215 157.230 ;
        RECT 30.405 156.580 30.735 157.060 ;
        RECT 30.905 156.770 31.130 157.230 ;
        RECT 31.300 156.580 31.630 157.060 ;
        RECT 29.455 155.820 29.630 156.430 ;
        RECT 30.405 156.410 31.630 156.580 ;
        RECT 32.260 156.450 32.760 157.060 ;
        RECT 33.800 156.450 34.300 157.060 ;
        RECT 29.800 156.070 30.495 156.240 ;
        RECT 30.325 155.820 30.495 156.070 ;
        RECT 30.670 156.040 31.090 156.240 ;
        RECT 31.260 156.040 31.590 156.240 ;
        RECT 31.760 156.040 32.090 156.240 ;
        RECT 32.260 155.820 32.430 156.450 ;
        RECT 32.615 155.990 32.965 156.240 ;
        RECT 33.595 155.990 33.945 156.240 ;
        RECT 34.130 155.820 34.300 156.450 ;
        RECT 34.930 156.580 35.260 157.060 ;
        RECT 35.430 156.770 35.655 157.230 ;
        RECT 35.825 156.580 36.155 157.060 ;
        RECT 34.930 156.410 36.155 156.580 ;
        RECT 36.345 156.430 36.595 157.230 ;
        RECT 36.765 156.430 37.105 157.060 ;
        RECT 37.480 156.450 37.980 157.060 ;
        RECT 34.470 156.040 34.800 156.240 ;
        RECT 34.970 156.040 35.300 156.240 ;
        RECT 35.470 156.040 35.890 156.240 ;
        RECT 36.065 156.070 36.760 156.240 ;
        RECT 36.065 155.820 36.235 156.070 ;
        RECT 36.930 155.820 37.105 156.430 ;
        RECT 37.275 155.990 37.625 156.240 ;
        RECT 37.810 155.820 37.980 156.450 ;
        RECT 38.610 156.580 38.940 157.060 ;
        RECT 39.110 156.770 39.335 157.230 ;
        RECT 39.505 156.580 39.835 157.060 ;
        RECT 38.610 156.410 39.835 156.580 ;
        RECT 40.025 156.430 40.275 157.230 ;
        RECT 40.445 156.430 40.785 157.060 ;
        RECT 41.415 156.460 44.005 157.230 ;
        RECT 44.180 156.685 49.525 157.230 ;
        RECT 38.150 156.040 38.480 156.240 ;
        RECT 38.650 156.040 38.980 156.240 ;
        RECT 39.150 156.040 39.570 156.240 ;
        RECT 39.745 156.070 40.440 156.240 ;
        RECT 39.745 155.820 39.915 156.070 ;
        RECT 40.610 155.820 40.785 156.430 ;
        RECT 29.455 154.850 29.795 155.820 ;
        RECT 29.965 154.680 30.135 155.820 ;
        RECT 30.325 155.650 32.760 155.820 ;
        RECT 30.405 154.680 30.655 155.480 ;
        RECT 31.300 154.850 31.630 155.650 ;
        RECT 31.930 154.680 32.260 155.480 ;
        RECT 32.430 154.850 32.760 155.650 ;
        RECT 33.800 155.650 36.235 155.820 ;
        RECT 33.800 154.850 34.130 155.650 ;
        RECT 34.300 154.680 34.630 155.480 ;
        RECT 34.930 154.850 35.260 155.650 ;
        RECT 35.905 154.680 36.155 155.480 ;
        RECT 36.425 154.680 36.595 155.820 ;
        RECT 36.765 154.850 37.105 155.820 ;
        RECT 37.480 155.650 39.915 155.820 ;
        RECT 37.480 154.850 37.810 155.650 ;
        RECT 37.980 154.680 38.310 155.480 ;
        RECT 38.610 154.850 38.940 155.650 ;
        RECT 39.585 154.680 39.835 155.480 ;
        RECT 40.105 154.680 40.275 155.820 ;
        RECT 40.445 154.850 40.785 155.820 ;
        RECT 41.415 155.770 42.625 156.290 ;
        RECT 42.795 155.940 44.005 156.460 ;
        RECT 41.415 154.680 44.005 155.770 ;
        RECT 45.770 155.115 46.120 156.365 ;
        RECT 47.600 155.855 47.940 156.685 ;
        RECT 49.785 156.680 49.955 157.060 ;
        RECT 50.135 156.850 50.465 157.230 ;
        RECT 49.785 156.510 50.450 156.680 ;
        RECT 50.645 156.555 50.905 157.060 ;
        RECT 49.715 155.960 50.045 156.330 ;
        RECT 50.280 156.255 50.450 156.510 ;
        RECT 50.280 155.925 50.565 156.255 ;
        RECT 50.280 155.780 50.450 155.925 ;
        RECT 49.785 155.610 50.450 155.780 ;
        RECT 50.735 155.755 50.905 156.555 ;
        RECT 51.075 156.505 51.365 157.230 ;
        RECT 51.910 156.520 52.165 157.050 ;
        RECT 52.345 156.770 52.630 157.230 ;
        RECT 44.180 154.680 49.525 155.115 ;
        RECT 49.785 154.850 49.955 155.610 ;
        RECT 50.135 154.680 50.465 155.440 ;
        RECT 50.635 154.850 50.905 155.755 ;
        RECT 51.075 154.680 51.365 155.845 ;
        RECT 51.910 155.660 52.090 156.520 ;
        RECT 52.810 156.320 53.060 156.970 ;
        RECT 52.260 155.990 53.060 156.320 ;
        RECT 51.910 155.190 52.165 155.660 ;
        RECT 51.825 155.020 52.165 155.190 ;
        RECT 51.910 154.990 52.165 155.020 ;
        RECT 52.345 154.680 52.630 155.480 ;
        RECT 52.810 155.400 53.060 155.990 ;
        RECT 53.260 156.635 53.580 156.965 ;
        RECT 53.760 156.750 54.420 157.230 ;
        RECT 54.620 156.840 55.470 157.010 ;
        RECT 53.260 155.740 53.450 156.635 ;
        RECT 53.770 156.310 54.430 156.580 ;
        RECT 54.100 156.250 54.430 156.310 ;
        RECT 53.620 156.080 53.950 156.140 ;
        RECT 54.620 156.080 54.790 156.840 ;
        RECT 56.030 156.770 56.350 157.230 ;
        RECT 56.550 156.590 56.800 157.020 ;
        RECT 57.090 156.790 57.500 157.230 ;
        RECT 57.670 156.850 58.685 157.050 ;
        RECT 54.960 156.420 56.210 156.590 ;
        RECT 54.960 156.300 55.290 156.420 ;
        RECT 53.620 155.910 55.520 156.080 ;
        RECT 53.260 155.570 55.180 155.740 ;
        RECT 53.260 155.550 53.580 155.570 ;
        RECT 52.810 154.890 53.140 155.400 ;
        RECT 53.410 154.940 53.580 155.550 ;
        RECT 55.350 155.400 55.520 155.910 ;
        RECT 55.690 155.840 55.870 156.250 ;
        RECT 56.040 155.660 56.210 156.420 ;
        RECT 53.750 154.680 54.080 155.370 ;
        RECT 54.310 155.230 55.520 155.400 ;
        RECT 55.690 155.350 56.210 155.660 ;
        RECT 56.380 156.250 56.800 156.590 ;
        RECT 57.090 156.250 57.500 156.580 ;
        RECT 56.380 155.480 56.570 156.250 ;
        RECT 57.670 156.120 57.840 156.850 ;
        RECT 58.985 156.680 59.155 157.010 ;
        RECT 59.325 156.850 59.655 157.230 ;
        RECT 58.010 156.300 58.360 156.670 ;
        RECT 57.670 156.080 58.090 156.120 ;
        RECT 56.740 155.910 58.090 156.080 ;
        RECT 56.740 155.750 56.990 155.910 ;
        RECT 57.500 155.480 57.750 155.740 ;
        RECT 56.380 155.230 57.750 155.480 ;
        RECT 54.310 154.940 54.550 155.230 ;
        RECT 55.350 155.150 55.520 155.230 ;
        RECT 54.750 154.680 55.170 155.060 ;
        RECT 55.350 154.900 55.980 155.150 ;
        RECT 56.450 154.680 56.780 155.060 ;
        RECT 56.950 154.940 57.120 155.230 ;
        RECT 57.920 155.065 58.090 155.910 ;
        RECT 58.540 155.740 58.760 156.610 ;
        RECT 58.985 156.490 59.680 156.680 ;
        RECT 58.260 155.360 58.760 155.740 ;
        RECT 58.930 155.690 59.340 156.310 ;
        RECT 59.510 155.520 59.680 156.490 ;
        RECT 58.985 155.350 59.680 155.520 ;
        RECT 57.300 154.680 57.680 155.060 ;
        RECT 57.920 154.895 58.750 155.065 ;
        RECT 58.985 154.850 59.155 155.350 ;
        RECT 59.325 154.680 59.655 155.180 ;
        RECT 59.870 154.850 60.095 156.970 ;
        RECT 60.265 156.850 60.595 157.230 ;
        RECT 60.765 156.680 60.935 156.970 ;
        RECT 60.270 156.510 60.935 156.680 ;
        RECT 60.270 155.520 60.500 156.510 ;
        RECT 61.200 156.390 61.460 157.230 ;
        RECT 61.635 156.485 61.890 157.060 ;
        RECT 62.060 156.850 62.390 157.230 ;
        RECT 62.605 156.680 62.775 157.060 ;
        RECT 62.060 156.510 62.775 156.680 ;
        RECT 63.125 156.680 63.295 157.060 ;
        RECT 63.510 156.850 63.840 157.230 ;
        RECT 63.125 156.510 63.840 156.680 ;
        RECT 60.670 155.690 61.020 156.340 ;
        RECT 60.270 155.350 60.935 155.520 ;
        RECT 60.265 154.680 60.595 155.180 ;
        RECT 60.765 154.850 60.935 155.350 ;
        RECT 61.200 154.680 61.460 155.830 ;
        RECT 61.635 155.755 61.805 156.485 ;
        RECT 62.060 156.320 62.230 156.510 ;
        RECT 61.975 155.990 62.230 156.320 ;
        RECT 62.060 155.780 62.230 155.990 ;
        RECT 62.510 155.960 62.865 156.330 ;
        RECT 63.035 155.960 63.390 156.330 ;
        RECT 63.670 156.320 63.840 156.510 ;
        RECT 64.010 156.485 64.265 157.060 ;
        RECT 63.670 155.990 63.925 156.320 ;
        RECT 63.670 155.780 63.840 155.990 ;
        RECT 61.635 154.850 61.890 155.755 ;
        RECT 62.060 155.610 62.775 155.780 ;
        RECT 62.060 154.680 62.390 155.440 ;
        RECT 62.605 154.850 62.775 155.610 ;
        RECT 63.125 155.610 63.840 155.780 ;
        RECT 64.095 155.755 64.265 156.485 ;
        RECT 64.440 156.390 64.700 157.230 ;
        RECT 65.080 156.450 65.580 157.060 ;
        RECT 64.875 155.990 65.225 156.240 ;
        RECT 63.125 154.850 63.295 155.610 ;
        RECT 63.510 154.680 63.840 155.440 ;
        RECT 64.010 154.850 64.265 155.755 ;
        RECT 64.440 154.680 64.700 155.830 ;
        RECT 65.410 155.820 65.580 156.450 ;
        RECT 66.210 156.580 66.540 157.060 ;
        RECT 66.710 156.770 66.935 157.230 ;
        RECT 67.105 156.580 67.435 157.060 ;
        RECT 66.210 156.410 67.435 156.580 ;
        RECT 67.625 156.430 67.875 157.230 ;
        RECT 68.045 156.430 68.385 157.060 ;
        RECT 65.750 156.040 66.080 156.240 ;
        RECT 66.250 156.040 66.580 156.240 ;
        RECT 66.750 156.040 67.170 156.240 ;
        RECT 67.345 156.070 68.040 156.240 ;
        RECT 67.345 155.820 67.515 156.070 ;
        RECT 68.210 155.820 68.385 156.430 ;
        RECT 65.080 155.650 67.515 155.820 ;
        RECT 65.080 154.850 65.410 155.650 ;
        RECT 65.580 154.680 65.910 155.480 ;
        RECT 66.210 154.850 66.540 155.650 ;
        RECT 67.185 154.680 67.435 155.480 ;
        RECT 67.705 154.680 67.875 155.820 ;
        RECT 68.045 154.850 68.385 155.820 ;
        RECT 68.555 156.430 68.895 157.060 ;
        RECT 69.065 156.430 69.315 157.230 ;
        RECT 69.505 156.580 69.835 157.060 ;
        RECT 70.005 156.770 70.230 157.230 ;
        RECT 70.400 156.580 70.730 157.060 ;
        RECT 68.555 155.820 68.730 156.430 ;
        RECT 69.505 156.410 70.730 156.580 ;
        RECT 71.360 156.450 71.860 157.060 ;
        RECT 73.155 156.460 76.665 157.230 ;
        RECT 76.835 156.505 77.125 157.230 ;
        RECT 78.215 156.460 81.725 157.230 ;
        RECT 81.900 156.685 87.245 157.230 ;
        RECT 68.900 156.070 69.595 156.240 ;
        RECT 69.425 155.820 69.595 156.070 ;
        RECT 69.770 156.040 70.190 156.240 ;
        RECT 70.360 156.040 70.690 156.240 ;
        RECT 70.860 156.040 71.190 156.240 ;
        RECT 71.360 155.820 71.530 156.450 ;
        RECT 71.715 155.990 72.065 156.240 ;
        RECT 68.555 154.850 68.895 155.820 ;
        RECT 69.065 154.680 69.235 155.820 ;
        RECT 69.425 155.650 71.860 155.820 ;
        RECT 69.505 154.680 69.755 155.480 ;
        RECT 70.400 154.850 70.730 155.650 ;
        RECT 71.030 154.680 71.360 155.480 ;
        RECT 71.530 154.850 71.860 155.650 ;
        RECT 73.155 155.770 74.845 156.290 ;
        RECT 75.015 155.940 76.665 156.460 ;
        RECT 73.155 154.680 76.665 155.770 ;
        RECT 76.835 154.680 77.125 155.845 ;
        RECT 78.215 155.770 79.905 156.290 ;
        RECT 80.075 155.940 81.725 156.460 ;
        RECT 78.215 154.680 81.725 155.770 ;
        RECT 83.490 155.115 83.840 156.365 ;
        RECT 85.320 155.855 85.660 156.685 ;
        RECT 87.415 156.430 87.755 157.060 ;
        RECT 87.925 156.430 88.175 157.230 ;
        RECT 88.365 156.580 88.695 157.060 ;
        RECT 88.865 156.770 89.090 157.230 ;
        RECT 89.260 156.580 89.590 157.060 ;
        RECT 87.415 155.820 87.590 156.430 ;
        RECT 88.365 156.410 89.590 156.580 ;
        RECT 90.220 156.450 90.720 157.060 ;
        RECT 91.095 156.460 93.685 157.230 ;
        RECT 87.760 156.070 88.455 156.240 ;
        RECT 88.285 155.820 88.455 156.070 ;
        RECT 88.630 156.040 89.050 156.240 ;
        RECT 89.220 156.040 89.550 156.240 ;
        RECT 89.720 156.040 90.050 156.240 ;
        RECT 90.220 155.820 90.390 156.450 ;
        RECT 90.575 155.990 90.925 156.240 ;
        RECT 81.900 154.680 87.245 155.115 ;
        RECT 87.415 154.850 87.755 155.820 ;
        RECT 87.925 154.680 88.095 155.820 ;
        RECT 88.285 155.650 90.720 155.820 ;
        RECT 88.365 154.680 88.615 155.480 ;
        RECT 89.260 154.850 89.590 155.650 ;
        RECT 89.890 154.680 90.220 155.480 ;
        RECT 90.390 154.850 90.720 155.650 ;
        RECT 91.095 155.770 92.305 156.290 ;
        RECT 92.475 155.940 93.685 156.460 ;
        RECT 93.855 156.430 94.195 157.060 ;
        RECT 94.365 156.430 94.615 157.230 ;
        RECT 94.805 156.580 95.135 157.060 ;
        RECT 95.305 156.770 95.530 157.230 ;
        RECT 95.700 156.580 96.030 157.060 ;
        RECT 93.855 155.820 94.030 156.430 ;
        RECT 94.805 156.410 96.030 156.580 ;
        RECT 96.660 156.450 97.160 157.060 ;
        RECT 97.535 156.480 98.745 157.230 ;
        RECT 94.200 156.070 94.895 156.240 ;
        RECT 94.725 155.820 94.895 156.070 ;
        RECT 95.070 156.040 95.490 156.240 ;
        RECT 95.660 156.040 95.990 156.240 ;
        RECT 96.160 156.040 96.490 156.240 ;
        RECT 96.660 155.820 96.830 156.450 ;
        RECT 97.015 155.990 97.365 156.240 ;
        RECT 91.095 154.680 93.685 155.770 ;
        RECT 93.855 154.850 94.195 155.820 ;
        RECT 94.365 154.680 94.535 155.820 ;
        RECT 94.725 155.650 97.160 155.820 ;
        RECT 94.805 154.680 95.055 155.480 ;
        RECT 95.700 154.850 96.030 155.650 ;
        RECT 96.330 154.680 96.660 155.480 ;
        RECT 96.830 154.850 97.160 155.650 ;
        RECT 97.535 155.770 98.055 156.310 ;
        RECT 98.225 155.940 98.745 156.480 ;
        RECT 98.915 156.430 99.255 157.060 ;
        RECT 99.425 156.430 99.675 157.230 ;
        RECT 99.865 156.580 100.195 157.060 ;
        RECT 100.365 156.770 100.590 157.230 ;
        RECT 100.760 156.580 101.090 157.060 ;
        RECT 98.915 155.820 99.090 156.430 ;
        RECT 99.865 156.410 101.090 156.580 ;
        RECT 101.720 156.450 102.220 157.060 ;
        RECT 102.595 156.505 102.885 157.230 ;
        RECT 103.055 156.460 104.725 157.230 ;
        RECT 99.260 156.070 99.955 156.240 ;
        RECT 99.785 155.820 99.955 156.070 ;
        RECT 100.130 156.040 100.550 156.240 ;
        RECT 100.720 156.040 101.050 156.240 ;
        RECT 101.220 156.040 101.550 156.240 ;
        RECT 101.720 155.820 101.890 156.450 ;
        RECT 102.075 155.990 102.425 156.240 ;
        RECT 97.535 154.680 98.745 155.770 ;
        RECT 98.915 154.850 99.255 155.820 ;
        RECT 99.425 154.680 99.595 155.820 ;
        RECT 99.785 155.650 102.220 155.820 ;
        RECT 99.865 154.680 100.115 155.480 ;
        RECT 100.760 154.850 101.090 155.650 ;
        RECT 101.390 154.680 101.720 155.480 ;
        RECT 101.890 154.850 102.220 155.650 ;
        RECT 102.595 154.680 102.885 155.845 ;
        RECT 103.055 155.770 103.805 156.290 ;
        RECT 103.975 155.940 104.725 156.460 ;
        RECT 105.010 156.600 105.295 157.060 ;
        RECT 105.465 156.770 105.735 157.230 ;
        RECT 105.010 156.430 105.965 156.600 ;
        RECT 103.055 154.680 104.725 155.770 ;
        RECT 104.895 155.700 105.585 156.260 ;
        RECT 105.755 155.530 105.965 156.430 ;
        RECT 105.010 155.310 105.965 155.530 ;
        RECT 106.135 156.260 106.535 157.060 ;
        RECT 106.725 156.600 107.005 157.060 ;
        RECT 107.525 156.770 107.850 157.230 ;
        RECT 106.725 156.430 107.850 156.600 ;
        RECT 108.020 156.490 108.405 157.060 ;
        RECT 107.400 156.320 107.850 156.430 ;
        RECT 106.135 155.700 107.230 156.260 ;
        RECT 107.400 155.990 107.955 156.320 ;
        RECT 105.010 154.850 105.295 155.310 ;
        RECT 105.465 154.680 105.735 155.140 ;
        RECT 106.135 154.850 106.535 155.700 ;
        RECT 107.400 155.530 107.850 155.990 ;
        RECT 108.125 155.820 108.405 156.490 ;
        RECT 108.665 156.580 108.835 157.060 ;
        RECT 109.015 156.750 109.255 157.230 ;
        RECT 109.505 156.580 109.675 157.060 ;
        RECT 109.845 156.750 110.175 157.230 ;
        RECT 110.345 156.580 110.515 157.060 ;
        RECT 108.665 156.410 109.300 156.580 ;
        RECT 109.505 156.410 110.515 156.580 ;
        RECT 110.685 156.430 111.015 157.230 ;
        RECT 111.795 156.460 114.385 157.230 ;
        RECT 114.555 156.480 115.765 157.230 ;
        RECT 109.130 156.240 109.300 156.410 ;
        RECT 108.580 156.000 108.960 156.240 ;
        RECT 109.130 156.070 109.630 156.240 ;
        RECT 109.130 155.830 109.300 156.070 ;
        RECT 110.020 155.870 110.515 156.410 ;
        RECT 106.725 155.310 107.850 155.530 ;
        RECT 106.725 154.850 107.005 155.310 ;
        RECT 107.525 154.680 107.850 155.140 ;
        RECT 108.020 154.850 108.405 155.820 ;
        RECT 108.585 155.660 109.300 155.830 ;
        RECT 109.505 155.700 110.515 155.870 ;
        RECT 108.585 154.850 108.915 155.660 ;
        RECT 109.085 154.680 109.325 155.480 ;
        RECT 109.505 154.850 109.675 155.700 ;
        RECT 109.845 154.680 110.175 155.480 ;
        RECT 110.345 154.850 110.515 155.700 ;
        RECT 110.685 154.680 111.015 155.830 ;
        RECT 111.795 155.770 113.005 156.290 ;
        RECT 113.175 155.940 114.385 156.460 ;
        RECT 114.555 155.770 115.075 156.310 ;
        RECT 115.245 155.940 115.765 156.480 ;
        RECT 111.795 154.680 114.385 155.770 ;
        RECT 114.555 154.680 115.765 155.770 ;
        RECT 10.510 154.510 115.850 154.680 ;
        RECT 10.595 153.420 11.805 154.510 ;
        RECT 10.595 152.710 11.115 153.250 ;
        RECT 11.285 152.880 11.805 153.420 ;
        RECT 12.435 153.345 12.725 154.510 ;
        RECT 13.270 154.170 13.525 154.200 ;
        RECT 13.185 154.000 13.525 154.170 ;
        RECT 13.270 153.530 13.525 154.000 ;
        RECT 13.705 153.710 13.990 154.510 ;
        RECT 14.170 153.790 14.500 154.300 ;
        RECT 10.595 151.960 11.805 152.710 ;
        RECT 12.435 151.960 12.725 152.685 ;
        RECT 13.270 152.670 13.450 153.530 ;
        RECT 14.170 153.200 14.420 153.790 ;
        RECT 14.770 153.640 14.940 154.250 ;
        RECT 15.110 153.820 15.440 154.510 ;
        RECT 15.670 153.960 15.910 154.250 ;
        RECT 16.110 154.130 16.530 154.510 ;
        RECT 16.710 154.040 17.340 154.290 ;
        RECT 17.810 154.130 18.140 154.510 ;
        RECT 16.710 153.960 16.880 154.040 ;
        RECT 18.310 153.960 18.480 154.250 ;
        RECT 18.660 154.130 19.040 154.510 ;
        RECT 19.280 154.125 20.110 154.295 ;
        RECT 15.670 153.790 16.880 153.960 ;
        RECT 13.620 152.870 14.420 153.200 ;
        RECT 13.270 152.140 13.525 152.670 ;
        RECT 13.705 151.960 13.990 152.420 ;
        RECT 14.170 152.220 14.420 152.870 ;
        RECT 14.620 153.620 14.940 153.640 ;
        RECT 14.620 153.450 16.540 153.620 ;
        RECT 14.620 152.555 14.810 153.450 ;
        RECT 16.710 153.280 16.880 153.790 ;
        RECT 17.050 153.530 17.570 153.840 ;
        RECT 14.980 153.110 16.880 153.280 ;
        RECT 14.980 153.050 15.310 153.110 ;
        RECT 15.460 152.880 15.790 152.940 ;
        RECT 15.130 152.610 15.790 152.880 ;
        RECT 14.620 152.225 14.940 152.555 ;
        RECT 15.120 151.960 15.780 152.440 ;
        RECT 15.980 152.350 16.150 153.110 ;
        RECT 17.050 152.940 17.230 153.350 ;
        RECT 16.320 152.770 16.650 152.890 ;
        RECT 17.400 152.770 17.570 153.530 ;
        RECT 16.320 152.600 17.570 152.770 ;
        RECT 17.740 153.710 19.110 153.960 ;
        RECT 17.740 152.940 17.930 153.710 ;
        RECT 18.860 153.450 19.110 153.710 ;
        RECT 18.100 153.280 18.350 153.440 ;
        RECT 19.280 153.280 19.450 154.125 ;
        RECT 20.345 153.840 20.515 154.340 ;
        RECT 20.685 154.010 21.015 154.510 ;
        RECT 19.620 153.450 20.120 153.830 ;
        RECT 20.345 153.670 21.040 153.840 ;
        RECT 18.100 153.110 19.450 153.280 ;
        RECT 19.030 153.070 19.450 153.110 ;
        RECT 17.740 152.600 18.160 152.940 ;
        RECT 18.450 152.610 18.860 152.940 ;
        RECT 15.980 152.180 16.830 152.350 ;
        RECT 17.390 151.960 17.710 152.420 ;
        RECT 17.910 152.170 18.160 152.600 ;
        RECT 18.450 151.960 18.860 152.400 ;
        RECT 19.030 152.340 19.200 153.070 ;
        RECT 19.370 152.520 19.720 152.890 ;
        RECT 19.900 152.580 20.120 153.450 ;
        RECT 20.290 152.880 20.700 153.500 ;
        RECT 20.870 152.700 21.040 153.670 ;
        RECT 20.345 152.510 21.040 152.700 ;
        RECT 19.030 152.140 20.045 152.340 ;
        RECT 20.345 152.180 20.515 152.510 ;
        RECT 20.685 151.960 21.015 152.340 ;
        RECT 21.230 152.220 21.455 154.340 ;
        RECT 21.625 154.010 21.955 154.510 ;
        RECT 22.125 153.840 22.295 154.340 ;
        RECT 21.630 153.670 22.295 153.840 ;
        RECT 21.630 152.680 21.860 153.670 ;
        RECT 22.030 152.850 22.380 153.500 ;
        RECT 22.555 153.435 22.825 154.340 ;
        RECT 22.995 153.750 23.325 154.510 ;
        RECT 23.505 153.580 23.675 154.340 ;
        RECT 21.630 152.510 22.295 152.680 ;
        RECT 21.625 151.960 21.955 152.340 ;
        RECT 22.125 152.220 22.295 152.510 ;
        RECT 22.555 152.635 22.725 153.435 ;
        RECT 23.010 153.410 23.675 153.580 ;
        RECT 24.395 153.420 27.905 154.510 ;
        RECT 23.010 153.265 23.180 153.410 ;
        RECT 22.895 152.935 23.180 153.265 ;
        RECT 23.010 152.680 23.180 152.935 ;
        RECT 23.415 152.860 23.745 153.230 ;
        RECT 24.395 152.900 26.085 153.420 ;
        RECT 28.080 153.370 28.415 154.340 ;
        RECT 28.585 153.370 28.755 154.510 ;
        RECT 28.925 154.170 30.955 154.340 ;
        RECT 26.255 152.730 27.905 153.250 ;
        RECT 22.555 152.130 22.815 152.635 ;
        RECT 23.010 152.510 23.675 152.680 ;
        RECT 22.995 151.960 23.325 152.340 ;
        RECT 23.505 152.130 23.675 152.510 ;
        RECT 24.395 151.960 27.905 152.730 ;
        RECT 28.080 152.700 28.250 153.370 ;
        RECT 28.925 153.200 29.095 154.170 ;
        RECT 28.420 152.870 28.675 153.200 ;
        RECT 28.900 152.870 29.095 153.200 ;
        RECT 29.265 153.830 30.390 154.000 ;
        RECT 28.505 152.700 28.675 152.870 ;
        RECT 29.265 152.700 29.435 153.830 ;
        RECT 28.080 152.130 28.335 152.700 ;
        RECT 28.505 152.530 29.435 152.700 ;
        RECT 29.605 153.490 30.615 153.660 ;
        RECT 29.605 152.690 29.775 153.490 ;
        RECT 29.980 153.150 30.255 153.290 ;
        RECT 29.975 152.980 30.255 153.150 ;
        RECT 29.260 152.495 29.435 152.530 ;
        RECT 28.505 151.960 28.835 152.360 ;
        RECT 29.260 152.130 29.790 152.495 ;
        RECT 29.980 152.130 30.255 152.980 ;
        RECT 30.425 152.130 30.615 153.490 ;
        RECT 30.785 153.505 30.955 154.170 ;
        RECT 31.125 153.750 31.295 154.510 ;
        RECT 31.530 153.750 32.045 154.160 ;
        RECT 32.680 154.075 38.025 154.510 ;
        RECT 30.785 153.315 31.535 153.505 ;
        RECT 31.705 152.940 32.045 153.750 ;
        RECT 30.815 152.770 32.045 152.940 ;
        RECT 34.270 152.825 34.620 154.075 ;
        RECT 38.195 153.345 38.485 154.510 ;
        RECT 39.575 153.420 43.085 154.510 ;
        RECT 43.260 154.075 48.605 154.510 ;
        RECT 30.795 151.960 31.305 152.495 ;
        RECT 31.525 152.165 31.770 152.770 ;
        RECT 36.100 152.505 36.440 153.335 ;
        RECT 39.575 152.900 41.265 153.420 ;
        RECT 41.435 152.730 43.085 153.250 ;
        RECT 44.850 152.825 45.200 154.075 ;
        RECT 48.780 153.370 49.115 154.340 ;
        RECT 49.285 153.370 49.455 154.510 ;
        RECT 49.625 154.170 51.655 154.340 ;
        RECT 32.680 151.960 38.025 152.505 ;
        RECT 38.195 151.960 38.485 152.685 ;
        RECT 39.575 151.960 43.085 152.730 ;
        RECT 46.680 152.505 47.020 153.335 ;
        RECT 48.780 152.700 48.950 153.370 ;
        RECT 49.625 153.200 49.795 154.170 ;
        RECT 49.120 152.870 49.375 153.200 ;
        RECT 49.600 152.870 49.795 153.200 ;
        RECT 49.965 153.830 51.090 154.000 ;
        RECT 49.205 152.700 49.375 152.870 ;
        RECT 49.965 152.700 50.135 153.830 ;
        RECT 43.260 151.960 48.605 152.505 ;
        RECT 48.780 152.130 49.035 152.700 ;
        RECT 49.205 152.530 50.135 152.700 ;
        RECT 50.305 153.490 51.315 153.660 ;
        RECT 50.305 152.690 50.475 153.490 ;
        RECT 49.960 152.495 50.135 152.530 ;
        RECT 49.205 151.960 49.535 152.360 ;
        RECT 49.960 152.130 50.490 152.495 ;
        RECT 50.680 152.470 50.955 153.290 ;
        RECT 50.675 152.300 50.955 152.470 ;
        RECT 50.680 152.130 50.955 152.300 ;
        RECT 51.125 152.130 51.315 153.490 ;
        RECT 51.485 153.505 51.655 154.170 ;
        RECT 51.825 153.750 51.995 154.510 ;
        RECT 52.230 153.750 52.745 154.160 ;
        RECT 51.485 153.315 52.235 153.505 ;
        RECT 52.405 152.940 52.745 153.750 ;
        RECT 51.515 152.770 52.745 152.940 ;
        RECT 52.920 153.370 53.255 154.340 ;
        RECT 53.425 153.370 53.595 154.510 ;
        RECT 53.765 154.170 55.795 154.340 ;
        RECT 51.495 151.960 52.005 152.495 ;
        RECT 52.225 152.165 52.470 152.770 ;
        RECT 52.920 152.700 53.090 153.370 ;
        RECT 53.765 153.200 53.935 154.170 ;
        RECT 53.260 152.870 53.515 153.200 ;
        RECT 53.740 152.870 53.935 153.200 ;
        RECT 54.105 153.830 55.230 154.000 ;
        RECT 53.345 152.700 53.515 152.870 ;
        RECT 54.105 152.700 54.275 153.830 ;
        RECT 52.920 152.130 53.175 152.700 ;
        RECT 53.345 152.530 54.275 152.700 ;
        RECT 54.445 153.490 55.455 153.660 ;
        RECT 54.445 152.690 54.615 153.490 ;
        RECT 54.100 152.495 54.275 152.530 ;
        RECT 53.345 151.960 53.675 152.360 ;
        RECT 54.100 152.130 54.630 152.495 ;
        RECT 54.820 152.470 55.095 153.290 ;
        RECT 54.815 152.300 55.095 152.470 ;
        RECT 54.820 152.130 55.095 152.300 ;
        RECT 55.265 152.130 55.455 153.490 ;
        RECT 55.625 153.505 55.795 154.170 ;
        RECT 55.965 153.750 56.135 154.510 ;
        RECT 56.370 153.750 56.885 154.160 ;
        RECT 55.625 153.315 56.375 153.505 ;
        RECT 56.545 152.940 56.885 153.750 ;
        RECT 58.065 153.580 58.235 154.340 ;
        RECT 58.415 153.750 58.745 154.510 ;
        RECT 58.065 153.410 58.730 153.580 ;
        RECT 58.915 153.435 59.185 154.340 ;
        RECT 58.560 153.265 58.730 153.410 ;
        RECT 55.655 152.770 56.885 152.940 ;
        RECT 57.995 152.860 58.325 153.230 ;
        RECT 58.560 152.935 58.845 153.265 ;
        RECT 55.635 151.960 56.145 152.495 ;
        RECT 56.365 152.165 56.610 152.770 ;
        RECT 58.560 152.680 58.730 152.935 ;
        RECT 58.065 152.510 58.730 152.680 ;
        RECT 59.015 152.635 59.185 153.435 ;
        RECT 59.360 153.360 59.620 154.510 ;
        RECT 59.795 153.435 60.050 154.340 ;
        RECT 60.220 153.750 60.550 154.510 ;
        RECT 60.765 153.580 60.935 154.340 ;
        RECT 58.065 152.130 58.235 152.510 ;
        RECT 58.415 151.960 58.745 152.340 ;
        RECT 58.925 152.130 59.185 152.635 ;
        RECT 59.360 151.960 59.620 152.800 ;
        RECT 59.795 152.705 59.965 153.435 ;
        RECT 60.220 153.410 60.935 153.580 ;
        RECT 60.220 153.200 60.390 153.410 ;
        RECT 61.200 153.360 61.460 154.510 ;
        RECT 61.635 153.435 61.890 154.340 ;
        RECT 62.060 153.750 62.390 154.510 ;
        RECT 62.605 153.580 62.775 154.340 ;
        RECT 60.135 152.870 60.390 153.200 ;
        RECT 59.795 152.130 60.050 152.705 ;
        RECT 60.220 152.680 60.390 152.870 ;
        RECT 60.670 152.860 61.025 153.230 ;
        RECT 60.220 152.510 60.935 152.680 ;
        RECT 60.220 151.960 60.550 152.340 ;
        RECT 60.765 152.130 60.935 152.510 ;
        RECT 61.200 151.960 61.460 152.800 ;
        RECT 61.635 152.705 61.805 153.435 ;
        RECT 62.060 153.410 62.775 153.580 ;
        RECT 62.060 153.200 62.230 153.410 ;
        RECT 63.955 153.345 64.245 154.510 ;
        RECT 64.420 153.360 64.680 154.510 ;
        RECT 64.855 153.435 65.110 154.340 ;
        RECT 65.280 153.750 65.610 154.510 ;
        RECT 65.825 153.580 65.995 154.340 ;
        RECT 61.975 152.870 62.230 153.200 ;
        RECT 61.635 152.130 61.890 152.705 ;
        RECT 62.060 152.680 62.230 152.870 ;
        RECT 62.510 152.860 62.865 153.230 ;
        RECT 62.060 152.510 62.775 152.680 ;
        RECT 62.060 151.960 62.390 152.340 ;
        RECT 62.605 152.130 62.775 152.510 ;
        RECT 63.955 151.960 64.245 152.685 ;
        RECT 64.420 151.960 64.680 152.800 ;
        RECT 64.855 152.705 65.025 153.435 ;
        RECT 65.280 153.410 65.995 153.580 ;
        RECT 66.265 153.450 66.595 154.510 ;
        RECT 65.280 153.200 65.450 153.410 ;
        RECT 65.195 152.870 65.450 153.200 ;
        RECT 64.855 152.130 65.110 152.705 ;
        RECT 65.280 152.680 65.450 152.870 ;
        RECT 65.730 152.860 66.085 153.230 ;
        RECT 66.775 153.200 66.945 154.125 ;
        RECT 67.115 153.920 67.445 154.320 ;
        RECT 67.615 154.150 67.945 154.510 ;
        RECT 68.145 153.920 68.845 154.340 ;
        RECT 67.115 153.690 68.845 153.920 ;
        RECT 67.115 153.470 67.445 153.690 ;
        RECT 67.640 153.200 67.965 153.490 ;
        RECT 66.255 152.870 66.565 153.200 ;
        RECT 66.775 152.870 67.150 153.200 ;
        RECT 67.470 152.870 67.965 153.200 ;
        RECT 68.140 152.950 68.470 153.490 ;
        RECT 68.640 152.720 68.845 153.690 ;
        RECT 65.280 152.510 65.995 152.680 ;
        RECT 65.280 151.960 65.610 152.340 ;
        RECT 65.825 152.130 65.995 152.510 ;
        RECT 66.265 152.490 67.625 152.700 ;
        RECT 66.265 152.130 66.595 152.490 ;
        RECT 66.765 151.960 67.095 152.320 ;
        RECT 67.295 152.130 67.625 152.490 ;
        RECT 68.135 152.130 68.845 152.720 ;
        RECT 69.015 153.370 69.355 154.340 ;
        RECT 69.525 153.370 69.695 154.510 ;
        RECT 69.965 153.710 70.215 154.510 ;
        RECT 70.860 153.540 71.190 154.340 ;
        RECT 71.490 153.710 71.820 154.510 ;
        RECT 71.990 153.540 72.320 154.340 ;
        RECT 69.885 153.370 72.320 153.540 ;
        RECT 73.155 153.420 75.745 154.510 ;
        RECT 75.920 154.075 81.265 154.510 ;
        RECT 69.015 152.810 69.190 153.370 ;
        RECT 69.885 153.120 70.055 153.370 ;
        RECT 69.360 152.950 70.055 153.120 ;
        RECT 70.230 152.950 70.650 153.150 ;
        RECT 70.820 152.950 71.150 153.150 ;
        RECT 71.320 152.950 71.650 153.150 ;
        RECT 69.015 152.760 69.245 152.810 ;
        RECT 69.015 152.130 69.355 152.760 ;
        RECT 69.525 151.960 69.775 152.760 ;
        RECT 69.965 152.610 71.190 152.780 ;
        RECT 69.965 152.130 70.295 152.610 ;
        RECT 70.465 151.960 70.690 152.420 ;
        RECT 70.860 152.130 71.190 152.610 ;
        RECT 71.820 152.740 71.990 153.370 ;
        RECT 72.175 152.950 72.525 153.200 ;
        RECT 73.155 152.900 74.365 153.420 ;
        RECT 71.820 152.130 72.320 152.740 ;
        RECT 74.535 152.730 75.745 153.250 ;
        RECT 77.510 152.825 77.860 154.075 ;
        RECT 81.495 153.370 81.705 154.510 ;
        RECT 81.875 153.360 82.205 154.340 ;
        RECT 82.375 153.370 82.605 154.510 ;
        RECT 82.905 153.580 83.075 154.340 ;
        RECT 83.255 153.750 83.585 154.510 ;
        RECT 82.905 153.410 83.570 153.580 ;
        RECT 83.755 153.435 84.025 154.340 ;
        RECT 73.155 151.960 75.745 152.730 ;
        RECT 79.340 152.505 79.680 153.335 ;
        RECT 75.920 151.960 81.265 152.505 ;
        RECT 81.495 151.960 81.705 152.780 ;
        RECT 81.875 152.760 82.125 153.360 ;
        RECT 83.400 153.265 83.570 153.410 ;
        RECT 82.295 152.950 82.625 153.200 ;
        RECT 82.835 152.860 83.165 153.230 ;
        RECT 83.400 152.935 83.685 153.265 ;
        RECT 81.875 152.130 82.205 152.760 ;
        RECT 82.375 151.960 82.605 152.780 ;
        RECT 83.400 152.680 83.570 152.935 ;
        RECT 82.905 152.510 83.570 152.680 ;
        RECT 83.855 152.635 84.025 153.435 ;
        RECT 84.655 153.420 88.165 154.510 ;
        RECT 84.655 152.900 86.345 153.420 ;
        RECT 88.375 153.370 88.605 154.510 ;
        RECT 88.775 153.360 89.105 154.340 ;
        RECT 89.275 153.370 89.485 154.510 ;
        RECT 86.515 152.730 88.165 153.250 ;
        RECT 88.355 152.950 88.685 153.200 ;
        RECT 82.905 152.130 83.075 152.510 ;
        RECT 83.255 151.960 83.585 152.340 ;
        RECT 83.765 152.130 84.025 152.635 ;
        RECT 84.655 151.960 88.165 152.730 ;
        RECT 88.375 151.960 88.605 152.780 ;
        RECT 88.855 152.760 89.105 153.360 ;
        RECT 89.715 153.345 90.005 154.510 ;
        RECT 90.180 154.075 95.525 154.510 ;
        RECT 91.770 152.825 92.120 154.075 ;
        RECT 95.695 153.370 96.035 154.340 ;
        RECT 96.205 153.370 96.375 154.510 ;
        RECT 96.645 153.710 96.895 154.510 ;
        RECT 97.540 153.540 97.870 154.340 ;
        RECT 98.170 153.710 98.500 154.510 ;
        RECT 98.670 153.540 99.000 154.340 ;
        RECT 99.950 153.880 100.235 154.340 ;
        RECT 100.405 154.050 100.675 154.510 ;
        RECT 99.950 153.660 100.905 153.880 ;
        RECT 96.565 153.370 99.000 153.540 ;
        RECT 88.775 152.130 89.105 152.760 ;
        RECT 89.275 151.960 89.485 152.780 ;
        RECT 89.715 151.960 90.005 152.685 ;
        RECT 93.600 152.505 93.940 153.335 ;
        RECT 95.695 152.760 95.870 153.370 ;
        RECT 96.565 153.120 96.735 153.370 ;
        RECT 96.040 152.950 96.735 153.120 ;
        RECT 96.910 152.950 97.330 153.150 ;
        RECT 97.500 152.950 97.830 153.150 ;
        RECT 98.000 152.950 98.330 153.150 ;
        RECT 90.180 151.960 95.525 152.505 ;
        RECT 95.695 152.130 96.035 152.760 ;
        RECT 96.205 151.960 96.455 152.760 ;
        RECT 96.645 152.610 97.870 152.780 ;
        RECT 96.645 152.130 96.975 152.610 ;
        RECT 97.145 151.960 97.370 152.420 ;
        RECT 97.540 152.130 97.870 152.610 ;
        RECT 98.500 152.740 98.670 153.370 ;
        RECT 98.855 152.950 99.205 153.200 ;
        RECT 99.835 152.930 100.525 153.490 ;
        RECT 100.695 152.760 100.905 153.660 ;
        RECT 98.500 152.130 99.000 152.740 ;
        RECT 99.950 152.590 100.905 152.760 ;
        RECT 101.075 153.490 101.475 154.340 ;
        RECT 101.665 153.880 101.945 154.340 ;
        RECT 102.465 154.050 102.790 154.510 ;
        RECT 101.665 153.660 102.790 153.880 ;
        RECT 101.075 152.930 102.170 153.490 ;
        RECT 102.340 153.200 102.790 153.660 ;
        RECT 102.960 153.370 103.345 154.340 ;
        RECT 99.950 152.130 100.235 152.590 ;
        RECT 100.405 151.960 100.675 152.420 ;
        RECT 101.075 152.130 101.475 152.930 ;
        RECT 102.340 152.870 102.895 153.200 ;
        RECT 102.340 152.760 102.790 152.870 ;
        RECT 101.665 152.590 102.790 152.760 ;
        RECT 103.065 152.700 103.345 153.370 ;
        RECT 103.515 153.750 104.030 154.160 ;
        RECT 104.265 153.750 104.435 154.510 ;
        RECT 104.605 154.170 106.635 154.340 ;
        RECT 103.515 152.940 103.855 153.750 ;
        RECT 104.605 153.505 104.775 154.170 ;
        RECT 105.170 153.830 106.295 154.000 ;
        RECT 104.025 153.315 104.775 153.505 ;
        RECT 104.945 153.490 105.955 153.660 ;
        RECT 103.515 152.770 104.745 152.940 ;
        RECT 101.665 152.130 101.945 152.590 ;
        RECT 102.465 151.960 102.790 152.420 ;
        RECT 102.960 152.130 103.345 152.700 ;
        RECT 103.790 152.165 104.035 152.770 ;
        RECT 104.255 151.960 104.765 152.495 ;
        RECT 104.945 152.130 105.135 153.490 ;
        RECT 105.305 152.470 105.580 153.290 ;
        RECT 105.785 152.690 105.955 153.490 ;
        RECT 106.125 152.700 106.295 153.830 ;
        RECT 106.465 153.200 106.635 154.170 ;
        RECT 106.805 153.370 106.975 154.510 ;
        RECT 107.145 153.370 107.480 154.340 ;
        RECT 106.465 152.870 106.660 153.200 ;
        RECT 106.885 152.870 107.140 153.200 ;
        RECT 106.885 152.700 107.055 152.870 ;
        RECT 107.310 152.700 107.480 153.370 ;
        RECT 107.655 153.420 109.325 154.510 ;
        RECT 109.585 153.580 109.755 154.340 ;
        RECT 109.935 153.750 110.265 154.510 ;
        RECT 107.655 152.900 108.405 153.420 ;
        RECT 109.585 153.410 110.250 153.580 ;
        RECT 110.435 153.435 110.705 154.340 ;
        RECT 110.080 153.265 110.250 153.410 ;
        RECT 108.575 152.730 109.325 153.250 ;
        RECT 109.515 152.860 109.845 153.230 ;
        RECT 110.080 152.935 110.365 153.265 ;
        RECT 106.125 152.530 107.055 152.700 ;
        RECT 106.125 152.495 106.300 152.530 ;
        RECT 105.305 152.300 105.585 152.470 ;
        RECT 105.305 152.130 105.580 152.300 ;
        RECT 105.770 152.130 106.300 152.495 ;
        RECT 106.725 151.960 107.055 152.360 ;
        RECT 107.225 152.130 107.480 152.700 ;
        RECT 107.655 151.960 109.325 152.730 ;
        RECT 110.080 152.680 110.250 152.935 ;
        RECT 109.585 152.510 110.250 152.680 ;
        RECT 110.535 152.635 110.705 153.435 ;
        RECT 110.875 153.420 114.385 154.510 ;
        RECT 114.555 153.420 115.765 154.510 ;
        RECT 110.875 152.900 112.565 153.420 ;
        RECT 112.735 152.730 114.385 153.250 ;
        RECT 114.555 152.880 115.075 153.420 ;
        RECT 109.585 152.130 109.755 152.510 ;
        RECT 109.935 151.960 110.265 152.340 ;
        RECT 110.445 152.130 110.705 152.635 ;
        RECT 110.875 151.960 114.385 152.730 ;
        RECT 115.245 152.710 115.765 153.250 ;
        RECT 114.555 151.960 115.765 152.710 ;
        RECT 10.510 151.790 115.850 151.960 ;
        RECT 10.595 151.040 11.805 151.790 ;
        RECT 11.975 151.040 13.185 151.790 ;
        RECT 10.595 150.500 11.115 151.040 ;
        RECT 11.285 150.330 11.805 150.870 ;
        RECT 10.595 149.240 11.805 150.330 ;
        RECT 11.975 150.330 12.495 150.870 ;
        RECT 12.665 150.500 13.185 151.040 ;
        RECT 13.355 151.020 16.865 151.790 ;
        RECT 13.355 150.330 15.045 150.850 ;
        RECT 15.215 150.500 16.865 151.020 ;
        RECT 17.310 150.980 17.555 151.585 ;
        RECT 17.775 151.255 18.285 151.790 ;
        RECT 17.035 150.810 18.265 150.980 ;
        RECT 11.975 149.240 13.185 150.330 ;
        RECT 13.355 149.240 16.865 150.330 ;
        RECT 17.035 150.000 17.375 150.810 ;
        RECT 17.545 150.245 18.295 150.435 ;
        RECT 17.035 149.590 17.550 150.000 ;
        RECT 17.785 149.240 17.955 150.000 ;
        RECT 18.125 149.580 18.295 150.245 ;
        RECT 18.465 150.260 18.655 151.620 ;
        RECT 18.825 151.110 19.100 151.620 ;
        RECT 19.290 151.255 19.820 151.620 ;
        RECT 20.245 151.390 20.575 151.790 ;
        RECT 19.645 151.220 19.820 151.255 ;
        RECT 18.825 150.940 19.105 151.110 ;
        RECT 18.825 150.460 19.100 150.940 ;
        RECT 19.305 150.260 19.475 151.060 ;
        RECT 18.465 150.090 19.475 150.260 ;
        RECT 19.645 151.050 20.575 151.220 ;
        RECT 20.745 151.050 21.000 151.620 ;
        RECT 19.645 149.920 19.815 151.050 ;
        RECT 20.405 150.880 20.575 151.050 ;
        RECT 18.690 149.750 19.815 149.920 ;
        RECT 19.985 150.550 20.180 150.880 ;
        RECT 20.405 150.550 20.660 150.880 ;
        RECT 19.985 149.580 20.155 150.550 ;
        RECT 20.830 150.380 21.000 151.050 ;
        RECT 21.175 151.020 23.765 151.790 ;
        RECT 18.125 149.410 20.155 149.580 ;
        RECT 20.325 149.240 20.495 150.380 ;
        RECT 20.665 149.410 21.000 150.380 ;
        RECT 21.175 150.330 22.385 150.850 ;
        RECT 22.555 150.500 23.765 151.020 ;
        RECT 23.975 150.970 24.205 151.790 ;
        RECT 24.375 150.990 24.705 151.620 ;
        RECT 23.955 150.550 24.285 150.800 ;
        RECT 24.455 150.390 24.705 150.990 ;
        RECT 24.875 150.970 25.085 151.790 ;
        RECT 25.315 151.065 25.605 151.790 ;
        RECT 26.150 151.080 26.405 151.610 ;
        RECT 26.585 151.330 26.870 151.790 ;
        RECT 26.150 150.770 26.330 151.080 ;
        RECT 27.050 150.880 27.300 151.530 ;
        RECT 26.065 150.600 26.330 150.770 ;
        RECT 21.175 149.240 23.765 150.330 ;
        RECT 23.975 149.240 24.205 150.380 ;
        RECT 24.375 149.410 24.705 150.390 ;
        RECT 24.875 149.240 25.085 150.380 ;
        RECT 25.315 149.240 25.605 150.405 ;
        RECT 26.150 150.220 26.330 150.600 ;
        RECT 26.500 150.550 27.300 150.880 ;
        RECT 26.150 149.550 26.405 150.220 ;
        RECT 26.585 149.240 26.870 150.040 ;
        RECT 27.050 149.960 27.300 150.550 ;
        RECT 27.500 151.195 27.820 151.525 ;
        RECT 28.000 151.310 28.660 151.790 ;
        RECT 28.860 151.400 29.710 151.570 ;
        RECT 27.500 150.300 27.690 151.195 ;
        RECT 28.010 150.870 28.670 151.140 ;
        RECT 28.340 150.810 28.670 150.870 ;
        RECT 27.860 150.640 28.190 150.700 ;
        RECT 28.860 150.640 29.030 151.400 ;
        RECT 30.270 151.330 30.590 151.790 ;
        RECT 30.790 151.150 31.040 151.580 ;
        RECT 31.330 151.350 31.740 151.790 ;
        RECT 31.910 151.410 32.925 151.610 ;
        RECT 29.200 150.980 30.450 151.150 ;
        RECT 29.200 150.860 29.530 150.980 ;
        RECT 27.860 150.470 29.760 150.640 ;
        RECT 27.500 150.130 29.420 150.300 ;
        RECT 27.500 150.110 27.820 150.130 ;
        RECT 27.050 149.450 27.380 149.960 ;
        RECT 27.650 149.500 27.820 150.110 ;
        RECT 29.590 149.960 29.760 150.470 ;
        RECT 29.930 150.400 30.110 150.810 ;
        RECT 30.280 150.220 30.450 150.980 ;
        RECT 27.990 149.240 28.320 149.930 ;
        RECT 28.550 149.790 29.760 149.960 ;
        RECT 29.930 149.910 30.450 150.220 ;
        RECT 30.620 150.810 31.040 151.150 ;
        RECT 31.330 150.810 31.740 151.140 ;
        RECT 30.620 150.040 30.810 150.810 ;
        RECT 31.910 150.680 32.080 151.410 ;
        RECT 33.225 151.240 33.395 151.570 ;
        RECT 33.565 151.410 33.895 151.790 ;
        RECT 32.250 150.860 32.600 151.230 ;
        RECT 31.910 150.640 32.330 150.680 ;
        RECT 30.980 150.470 32.330 150.640 ;
        RECT 30.980 150.310 31.230 150.470 ;
        RECT 31.740 150.040 31.990 150.300 ;
        RECT 30.620 149.790 31.990 150.040 ;
        RECT 28.550 149.500 28.790 149.790 ;
        RECT 29.590 149.710 29.760 149.790 ;
        RECT 28.990 149.240 29.410 149.620 ;
        RECT 29.590 149.460 30.220 149.710 ;
        RECT 30.690 149.240 31.020 149.620 ;
        RECT 31.190 149.500 31.360 149.790 ;
        RECT 32.160 149.625 32.330 150.470 ;
        RECT 32.780 150.300 33.000 151.170 ;
        RECT 33.225 151.050 33.920 151.240 ;
        RECT 32.500 149.920 33.000 150.300 ;
        RECT 33.170 150.250 33.580 150.870 ;
        RECT 33.750 150.080 33.920 151.050 ;
        RECT 33.225 149.910 33.920 150.080 ;
        RECT 31.540 149.240 31.920 149.620 ;
        RECT 32.160 149.455 32.990 149.625 ;
        RECT 33.225 149.410 33.395 149.910 ;
        RECT 33.565 149.240 33.895 149.740 ;
        RECT 34.110 149.410 34.335 151.530 ;
        RECT 34.505 151.410 34.835 151.790 ;
        RECT 35.005 151.240 35.175 151.530 ;
        RECT 34.510 151.070 35.175 151.240 ;
        RECT 34.510 150.080 34.740 151.070 ;
        RECT 35.435 150.990 35.775 151.620 ;
        RECT 35.945 150.990 36.195 151.790 ;
        RECT 36.385 151.140 36.715 151.620 ;
        RECT 36.885 151.330 37.110 151.790 ;
        RECT 37.280 151.140 37.610 151.620 ;
        RECT 34.910 150.250 35.260 150.900 ;
        RECT 35.435 150.380 35.610 150.990 ;
        RECT 36.385 150.970 37.610 151.140 ;
        RECT 38.240 151.010 38.740 151.620 ;
        RECT 39.115 151.040 40.325 151.790 ;
        RECT 40.505 151.290 40.835 151.790 ;
        RECT 41.035 151.220 41.205 151.570 ;
        RECT 41.405 151.390 41.735 151.790 ;
        RECT 41.905 151.220 42.075 151.570 ;
        RECT 42.245 151.390 42.625 151.790 ;
        RECT 35.780 150.630 36.475 150.800 ;
        RECT 36.305 150.380 36.475 150.630 ;
        RECT 36.650 150.600 37.070 150.800 ;
        RECT 37.240 150.600 37.570 150.800 ;
        RECT 37.740 150.600 38.070 150.800 ;
        RECT 38.240 150.380 38.410 151.010 ;
        RECT 38.595 150.550 38.945 150.800 ;
        RECT 34.510 149.910 35.175 150.080 ;
        RECT 34.505 149.240 34.835 149.740 ;
        RECT 35.005 149.410 35.175 149.910 ;
        RECT 35.435 149.410 35.775 150.380 ;
        RECT 35.945 149.240 36.115 150.380 ;
        RECT 36.305 150.210 38.740 150.380 ;
        RECT 36.385 149.240 36.635 150.040 ;
        RECT 37.280 149.410 37.610 150.210 ;
        RECT 37.910 149.240 38.240 150.040 ;
        RECT 38.410 149.410 38.740 150.210 ;
        RECT 39.115 150.330 39.635 150.870 ;
        RECT 39.805 150.500 40.325 151.040 ;
        RECT 40.500 150.550 40.850 151.120 ;
        RECT 41.035 151.050 42.645 151.220 ;
        RECT 42.815 151.115 43.085 151.460 ;
        RECT 42.475 150.880 42.645 151.050 ;
        RECT 41.020 150.430 41.730 150.880 ;
        RECT 41.900 150.550 42.305 150.880 ;
        RECT 42.475 150.550 42.745 150.880 ;
        RECT 39.115 149.240 40.325 150.330 ;
        RECT 40.500 150.090 40.820 150.380 ;
        RECT 41.015 150.260 41.730 150.430 ;
        RECT 42.475 150.380 42.645 150.550 ;
        RECT 42.915 150.380 43.085 151.115 ;
        RECT 41.920 150.210 42.645 150.380 ;
        RECT 41.920 150.090 42.090 150.210 ;
        RECT 40.500 149.920 42.090 150.090 ;
        RECT 40.500 149.460 42.155 149.750 ;
        RECT 42.325 149.240 42.605 150.040 ;
        RECT 42.815 149.410 43.085 150.380 ;
        RECT 43.255 151.115 43.525 151.460 ;
        RECT 43.715 151.390 44.095 151.790 ;
        RECT 44.265 151.220 44.435 151.570 ;
        RECT 44.605 151.390 44.935 151.790 ;
        RECT 45.135 151.220 45.305 151.570 ;
        RECT 45.505 151.290 45.835 151.790 ;
        RECT 43.255 150.380 43.425 151.115 ;
        RECT 43.695 151.050 45.305 151.220 ;
        RECT 43.695 150.880 43.865 151.050 ;
        RECT 43.595 150.550 43.865 150.880 ;
        RECT 44.035 150.550 44.440 150.880 ;
        RECT 43.695 150.380 43.865 150.550 ;
        RECT 43.255 149.410 43.525 150.380 ;
        RECT 43.695 150.210 44.420 150.380 ;
        RECT 44.610 150.260 45.320 150.880 ;
        RECT 45.490 150.550 45.840 151.120 ;
        RECT 46.475 150.990 46.815 151.620 ;
        RECT 46.985 150.990 47.235 151.790 ;
        RECT 47.425 151.140 47.755 151.620 ;
        RECT 47.925 151.330 48.150 151.790 ;
        RECT 48.320 151.140 48.650 151.620 ;
        RECT 46.475 150.940 46.705 150.990 ;
        RECT 47.425 150.970 48.650 151.140 ;
        RECT 49.280 151.010 49.780 151.620 ;
        RECT 51.075 151.065 51.365 151.790 ;
        RECT 46.475 150.380 46.650 150.940 ;
        RECT 46.820 150.630 47.515 150.800 ;
        RECT 47.345 150.380 47.515 150.630 ;
        RECT 47.690 150.600 48.110 150.800 ;
        RECT 48.280 150.600 48.610 150.800 ;
        RECT 48.780 150.600 49.110 150.800 ;
        RECT 49.280 150.380 49.450 151.010 ;
        RECT 52.035 150.970 52.265 151.790 ;
        RECT 52.435 150.990 52.765 151.620 ;
        RECT 49.635 150.550 49.985 150.800 ;
        RECT 52.015 150.550 52.345 150.800 ;
        RECT 44.250 150.090 44.420 150.210 ;
        RECT 45.520 150.090 45.840 150.380 ;
        RECT 43.735 149.240 44.015 150.040 ;
        RECT 44.250 149.920 45.840 150.090 ;
        RECT 44.185 149.460 45.840 149.750 ;
        RECT 46.475 149.410 46.815 150.380 ;
        RECT 46.985 149.240 47.155 150.380 ;
        RECT 47.345 150.210 49.780 150.380 ;
        RECT 47.425 149.240 47.675 150.040 ;
        RECT 48.320 149.410 48.650 150.210 ;
        RECT 48.950 149.240 49.280 150.040 ;
        RECT 49.450 149.410 49.780 150.210 ;
        RECT 51.075 149.240 51.365 150.405 ;
        RECT 52.515 150.390 52.765 150.990 ;
        RECT 52.935 150.970 53.145 151.790 ;
        RECT 53.465 151.240 53.635 151.620 ;
        RECT 53.815 151.410 54.145 151.790 ;
        RECT 53.465 151.070 54.130 151.240 ;
        RECT 54.325 151.115 54.585 151.620 ;
        RECT 54.845 151.310 55.145 151.790 ;
        RECT 55.315 151.140 55.575 151.595 ;
        RECT 55.745 151.310 56.005 151.790 ;
        RECT 56.185 151.140 56.445 151.595 ;
        RECT 56.615 151.310 56.865 151.790 ;
        RECT 57.045 151.140 57.305 151.595 ;
        RECT 57.475 151.310 57.725 151.790 ;
        RECT 57.905 151.140 58.165 151.595 ;
        RECT 58.335 151.310 58.580 151.790 ;
        RECT 58.750 151.140 59.025 151.595 ;
        RECT 59.195 151.310 59.440 151.790 ;
        RECT 59.610 151.140 59.870 151.595 ;
        RECT 60.040 151.310 60.300 151.790 ;
        RECT 60.470 151.140 60.730 151.595 ;
        RECT 60.900 151.310 61.160 151.790 ;
        RECT 61.330 151.140 61.590 151.595 ;
        RECT 61.760 151.230 62.020 151.790 ;
        RECT 53.395 150.520 53.725 150.890 ;
        RECT 53.960 150.815 54.130 151.070 ;
        RECT 52.035 149.240 52.265 150.380 ;
        RECT 52.435 149.410 52.765 150.390 ;
        RECT 53.960 150.485 54.245 150.815 ;
        RECT 52.935 149.240 53.145 150.380 ;
        RECT 53.960 150.340 54.130 150.485 ;
        RECT 53.465 150.170 54.130 150.340 ;
        RECT 54.415 150.315 54.585 151.115 ;
        RECT 53.465 149.410 53.635 150.170 ;
        RECT 53.815 149.240 54.145 150.000 ;
        RECT 54.315 149.410 54.585 150.315 ;
        RECT 54.845 150.970 61.590 151.140 ;
        RECT 54.845 150.380 56.010 150.970 ;
        RECT 62.190 150.800 62.440 151.610 ;
        RECT 62.620 151.265 62.880 151.790 ;
        RECT 63.050 150.800 63.300 151.610 ;
        RECT 63.480 151.280 63.785 151.790 ;
        RECT 64.015 151.310 64.295 151.790 ;
        RECT 64.465 151.140 64.725 151.530 ;
        RECT 64.900 151.310 65.155 151.790 ;
        RECT 65.325 151.140 65.620 151.530 ;
        RECT 65.800 151.310 66.075 151.790 ;
        RECT 66.245 151.290 66.545 151.620 ;
        RECT 56.180 150.550 63.300 150.800 ;
        RECT 63.470 150.550 63.785 151.110 ;
        RECT 63.970 150.970 65.620 151.140 ;
        RECT 54.845 150.155 61.590 150.380 ;
        RECT 54.845 149.240 55.115 149.985 ;
        RECT 55.285 149.415 55.575 150.155 ;
        RECT 56.185 150.140 61.590 150.155 ;
        RECT 55.745 149.245 56.000 149.970 ;
        RECT 56.185 149.415 56.445 150.140 ;
        RECT 56.615 149.245 56.860 149.970 ;
        RECT 57.045 149.415 57.305 150.140 ;
        RECT 57.475 149.245 57.720 149.970 ;
        RECT 57.905 149.415 58.165 150.140 ;
        RECT 58.335 149.245 58.580 149.970 ;
        RECT 58.750 149.415 59.010 150.140 ;
        RECT 59.180 149.245 59.440 149.970 ;
        RECT 59.610 149.415 59.870 150.140 ;
        RECT 60.040 149.245 60.300 149.970 ;
        RECT 60.470 149.415 60.730 150.140 ;
        RECT 60.900 149.245 61.160 149.970 ;
        RECT 61.330 149.415 61.590 150.140 ;
        RECT 61.760 149.245 62.020 150.040 ;
        RECT 62.190 149.415 62.440 150.550 ;
        RECT 55.745 149.240 62.020 149.245 ;
        RECT 62.620 149.240 62.880 150.050 ;
        RECT 63.055 149.410 63.300 150.550 ;
        RECT 63.970 150.460 64.375 150.970 ;
        RECT 64.545 150.630 65.685 150.800 ;
        RECT 63.970 150.290 64.725 150.460 ;
        RECT 63.480 149.240 63.775 150.050 ;
        RECT 64.010 149.240 64.295 150.110 ;
        RECT 64.465 150.040 64.725 150.290 ;
        RECT 65.515 150.380 65.685 150.630 ;
        RECT 65.855 150.550 66.205 151.120 ;
        RECT 66.375 150.380 66.545 151.290 ;
        RECT 66.715 151.040 67.925 151.790 ;
        RECT 65.515 150.210 66.545 150.380 ;
        RECT 64.465 149.870 65.585 150.040 ;
        RECT 64.465 149.410 64.725 149.870 ;
        RECT 64.900 149.240 65.155 149.700 ;
        RECT 65.325 149.410 65.585 149.870 ;
        RECT 65.755 149.240 66.065 150.040 ;
        RECT 66.235 149.410 66.545 150.210 ;
        RECT 66.715 150.330 67.235 150.870 ;
        RECT 67.405 150.500 67.925 151.040 ;
        RECT 68.095 151.115 68.365 151.460 ;
        RECT 68.555 151.390 68.935 151.790 ;
        RECT 69.105 151.220 69.275 151.570 ;
        RECT 69.445 151.390 69.775 151.790 ;
        RECT 69.975 151.220 70.145 151.570 ;
        RECT 70.345 151.290 70.675 151.790 ;
        RECT 70.855 151.290 71.155 151.620 ;
        RECT 71.325 151.310 71.600 151.790 ;
        RECT 68.095 150.380 68.265 151.115 ;
        RECT 68.535 151.050 70.145 151.220 ;
        RECT 68.535 150.880 68.705 151.050 ;
        RECT 68.435 150.550 68.705 150.880 ;
        RECT 68.875 150.550 69.280 150.880 ;
        RECT 68.535 150.380 68.705 150.550 ;
        RECT 69.450 150.430 70.160 150.880 ;
        RECT 70.330 150.550 70.680 151.120 ;
        RECT 66.715 149.240 67.925 150.330 ;
        RECT 68.095 149.410 68.365 150.380 ;
        RECT 68.535 150.210 69.260 150.380 ;
        RECT 69.450 150.260 70.165 150.430 ;
        RECT 70.855 150.380 71.025 151.290 ;
        RECT 71.780 151.140 72.075 151.530 ;
        RECT 72.245 151.310 72.500 151.790 ;
        RECT 72.675 151.140 72.935 151.530 ;
        RECT 73.105 151.310 73.385 151.790 ;
        RECT 71.195 150.550 71.545 151.120 ;
        RECT 71.780 150.970 73.430 151.140 ;
        RECT 74.075 151.020 76.665 151.790 ;
        RECT 76.835 151.065 77.125 151.790 ;
        RECT 77.670 151.080 77.925 151.610 ;
        RECT 78.105 151.330 78.390 151.790 ;
        RECT 71.715 150.630 72.855 150.800 ;
        RECT 71.715 150.380 71.885 150.630 ;
        RECT 73.025 150.460 73.430 150.970 ;
        RECT 69.090 150.090 69.260 150.210 ;
        RECT 70.360 150.090 70.680 150.380 ;
        RECT 68.575 149.240 68.855 150.040 ;
        RECT 69.090 149.920 70.680 150.090 ;
        RECT 70.855 150.210 71.885 150.380 ;
        RECT 72.675 150.290 73.430 150.460 ;
        RECT 74.075 150.330 75.285 150.850 ;
        RECT 75.455 150.500 76.665 151.020 ;
        RECT 69.025 149.460 70.680 149.750 ;
        RECT 70.855 149.410 71.165 150.210 ;
        RECT 72.675 150.040 72.935 150.290 ;
        RECT 71.335 149.240 71.645 150.040 ;
        RECT 71.815 149.870 72.935 150.040 ;
        RECT 71.815 149.410 72.075 149.870 ;
        RECT 72.245 149.240 72.500 149.700 ;
        RECT 72.675 149.410 72.935 149.870 ;
        RECT 73.105 149.240 73.390 150.110 ;
        RECT 74.075 149.240 76.665 150.330 ;
        RECT 76.835 149.240 77.125 150.405 ;
        RECT 77.670 150.220 77.850 151.080 ;
        RECT 78.570 150.880 78.820 151.530 ;
        RECT 78.020 150.550 78.820 150.880 ;
        RECT 77.670 149.750 77.925 150.220 ;
        RECT 77.585 149.580 77.925 149.750 ;
        RECT 77.670 149.550 77.925 149.580 ;
        RECT 78.105 149.240 78.390 150.040 ;
        RECT 78.570 149.960 78.820 150.550 ;
        RECT 79.020 151.195 79.340 151.525 ;
        RECT 79.520 151.310 80.180 151.790 ;
        RECT 80.380 151.400 81.230 151.570 ;
        RECT 79.020 150.300 79.210 151.195 ;
        RECT 79.530 150.870 80.190 151.140 ;
        RECT 79.860 150.810 80.190 150.870 ;
        RECT 79.380 150.640 79.710 150.700 ;
        RECT 80.380 150.640 80.550 151.400 ;
        RECT 81.790 151.330 82.110 151.790 ;
        RECT 82.310 151.150 82.560 151.580 ;
        RECT 82.850 151.350 83.260 151.790 ;
        RECT 83.430 151.410 84.445 151.610 ;
        RECT 80.720 150.980 81.970 151.150 ;
        RECT 80.720 150.860 81.050 150.980 ;
        RECT 79.380 150.470 81.280 150.640 ;
        RECT 79.020 150.130 80.940 150.300 ;
        RECT 79.020 150.110 79.340 150.130 ;
        RECT 78.570 149.450 78.900 149.960 ;
        RECT 79.170 149.500 79.340 150.110 ;
        RECT 81.110 149.960 81.280 150.470 ;
        RECT 81.450 150.400 81.630 150.810 ;
        RECT 81.800 150.220 81.970 150.980 ;
        RECT 79.510 149.240 79.840 149.930 ;
        RECT 80.070 149.790 81.280 149.960 ;
        RECT 81.450 149.910 81.970 150.220 ;
        RECT 82.140 150.810 82.560 151.150 ;
        RECT 82.850 150.810 83.260 151.140 ;
        RECT 82.140 150.040 82.330 150.810 ;
        RECT 83.430 150.680 83.600 151.410 ;
        RECT 84.745 151.240 84.915 151.570 ;
        RECT 85.085 151.410 85.415 151.790 ;
        RECT 83.770 150.860 84.120 151.230 ;
        RECT 83.430 150.640 83.850 150.680 ;
        RECT 82.500 150.470 83.850 150.640 ;
        RECT 82.500 150.310 82.750 150.470 ;
        RECT 83.260 150.040 83.510 150.300 ;
        RECT 82.140 149.790 83.510 150.040 ;
        RECT 80.070 149.500 80.310 149.790 ;
        RECT 81.110 149.710 81.280 149.790 ;
        RECT 80.510 149.240 80.930 149.620 ;
        RECT 81.110 149.460 81.740 149.710 ;
        RECT 82.210 149.240 82.540 149.620 ;
        RECT 82.710 149.500 82.880 149.790 ;
        RECT 83.680 149.625 83.850 150.470 ;
        RECT 84.300 150.300 84.520 151.170 ;
        RECT 84.745 151.050 85.440 151.240 ;
        RECT 84.020 149.920 84.520 150.300 ;
        RECT 84.690 150.250 85.100 150.870 ;
        RECT 85.270 150.080 85.440 151.050 ;
        RECT 84.745 149.910 85.440 150.080 ;
        RECT 83.060 149.240 83.440 149.620 ;
        RECT 83.680 149.455 84.510 149.625 ;
        RECT 84.745 149.410 84.915 149.910 ;
        RECT 85.085 149.240 85.415 149.740 ;
        RECT 85.630 149.410 85.855 151.530 ;
        RECT 86.025 151.410 86.355 151.790 ;
        RECT 86.525 151.240 86.695 151.530 ;
        RECT 86.030 151.070 86.695 151.240 ;
        RECT 86.960 151.080 87.215 151.610 ;
        RECT 87.385 151.330 87.690 151.790 ;
        RECT 87.935 151.410 89.005 151.580 ;
        RECT 86.030 150.080 86.260 151.070 ;
        RECT 86.430 150.250 86.780 150.900 ;
        RECT 86.960 150.430 87.170 151.080 ;
        RECT 87.935 151.055 88.255 151.410 ;
        RECT 87.930 150.880 88.255 151.055 ;
        RECT 87.340 150.580 88.255 150.880 ;
        RECT 88.425 150.840 88.665 151.240 ;
        RECT 88.835 151.180 89.005 151.410 ;
        RECT 89.175 151.350 89.365 151.790 ;
        RECT 89.535 151.340 90.485 151.620 ;
        RECT 90.705 151.430 91.055 151.600 ;
        RECT 88.835 151.010 89.365 151.180 ;
        RECT 87.340 150.550 88.080 150.580 ;
        RECT 86.030 149.910 86.695 150.080 ;
        RECT 86.025 149.240 86.355 149.740 ;
        RECT 86.525 149.410 86.695 149.910 ;
        RECT 86.960 149.550 87.215 150.430 ;
        RECT 87.385 149.240 87.690 150.380 ;
        RECT 87.910 149.960 88.080 150.550 ;
        RECT 88.425 150.470 88.965 150.840 ;
        RECT 89.145 150.730 89.365 151.010 ;
        RECT 89.535 150.560 89.705 151.340 ;
        RECT 89.300 150.390 89.705 150.560 ;
        RECT 89.875 150.550 90.225 151.170 ;
        RECT 89.300 150.300 89.470 150.390 ;
        RECT 90.395 150.380 90.605 151.170 ;
        RECT 88.250 150.130 89.470 150.300 ;
        RECT 89.930 150.220 90.605 150.380 ;
        RECT 87.910 149.790 88.710 149.960 ;
        RECT 88.030 149.240 88.360 149.620 ;
        RECT 88.540 149.500 88.710 149.790 ;
        RECT 89.300 149.750 89.470 150.130 ;
        RECT 89.640 150.210 90.605 150.220 ;
        RECT 90.795 151.040 91.055 151.430 ;
        RECT 91.265 151.330 91.595 151.790 ;
        RECT 92.470 151.400 93.325 151.570 ;
        RECT 93.530 151.400 94.025 151.570 ;
        RECT 94.195 151.430 94.525 151.790 ;
        RECT 90.795 150.350 90.965 151.040 ;
        RECT 91.135 150.690 91.305 150.870 ;
        RECT 91.475 150.860 92.265 151.110 ;
        RECT 92.470 150.690 92.640 151.400 ;
        RECT 92.810 150.890 93.165 151.110 ;
        RECT 91.135 150.520 92.825 150.690 ;
        RECT 89.640 149.920 90.100 150.210 ;
        RECT 90.795 150.180 92.295 150.350 ;
        RECT 90.795 150.040 90.965 150.180 ;
        RECT 90.405 149.870 90.965 150.040 ;
        RECT 88.880 149.240 89.130 149.700 ;
        RECT 89.300 149.410 90.170 149.750 ;
        RECT 90.405 149.410 90.575 149.870 ;
        RECT 91.410 149.840 92.485 150.010 ;
        RECT 90.745 149.240 91.115 149.700 ;
        RECT 91.410 149.500 91.580 149.840 ;
        RECT 91.750 149.240 92.080 149.670 ;
        RECT 92.315 149.500 92.485 149.840 ;
        RECT 92.655 149.740 92.825 150.520 ;
        RECT 92.995 150.300 93.165 150.890 ;
        RECT 93.335 150.490 93.685 151.110 ;
        RECT 92.995 149.910 93.460 150.300 ;
        RECT 93.855 150.040 94.025 151.400 ;
        RECT 94.195 150.210 94.655 151.260 ;
        RECT 93.630 149.870 94.025 150.040 ;
        RECT 93.630 149.740 93.800 149.870 ;
        RECT 92.655 149.410 93.335 149.740 ;
        RECT 93.550 149.410 93.800 149.740 ;
        RECT 93.970 149.240 94.220 149.700 ;
        RECT 94.390 149.425 94.715 150.210 ;
        RECT 94.885 149.410 95.055 151.530 ;
        RECT 95.225 151.410 95.555 151.790 ;
        RECT 95.725 151.240 95.980 151.530 ;
        RECT 95.230 151.070 95.980 151.240 ;
        RECT 96.155 151.115 96.425 151.460 ;
        RECT 96.615 151.390 96.995 151.790 ;
        RECT 97.165 151.220 97.335 151.570 ;
        RECT 97.505 151.390 97.835 151.790 ;
        RECT 98.035 151.220 98.205 151.570 ;
        RECT 98.405 151.290 98.735 151.790 ;
        RECT 95.230 150.080 95.460 151.070 ;
        RECT 95.630 150.250 95.980 150.900 ;
        RECT 96.155 150.380 96.325 151.115 ;
        RECT 96.595 151.050 98.205 151.220 ;
        RECT 96.595 150.880 96.765 151.050 ;
        RECT 96.495 150.550 96.765 150.880 ;
        RECT 96.935 150.550 97.340 150.880 ;
        RECT 96.595 150.380 96.765 150.550 ;
        RECT 97.510 150.430 98.220 150.880 ;
        RECT 98.390 150.550 98.740 151.120 ;
        RECT 98.915 150.990 99.255 151.620 ;
        RECT 99.425 150.990 99.675 151.790 ;
        RECT 99.865 151.140 100.195 151.620 ;
        RECT 100.365 151.330 100.590 151.790 ;
        RECT 100.760 151.140 101.090 151.620 ;
        RECT 98.915 150.940 99.145 150.990 ;
        RECT 99.865 150.970 101.090 151.140 ;
        RECT 101.720 151.010 102.220 151.620 ;
        RECT 102.595 151.065 102.885 151.790 ;
        RECT 95.230 149.910 95.980 150.080 ;
        RECT 95.225 149.240 95.555 149.740 ;
        RECT 95.725 149.410 95.980 149.910 ;
        RECT 96.155 149.410 96.425 150.380 ;
        RECT 96.595 150.210 97.320 150.380 ;
        RECT 97.510 150.260 98.225 150.430 ;
        RECT 98.915 150.380 99.090 150.940 ;
        RECT 99.260 150.630 99.955 150.800 ;
        RECT 100.130 150.770 100.550 150.800 ;
        RECT 99.785 150.380 99.955 150.630 ;
        RECT 100.125 150.600 100.550 150.770 ;
        RECT 100.720 150.600 101.050 150.800 ;
        RECT 101.220 150.600 101.550 150.800 ;
        RECT 101.720 150.380 101.890 151.010 ;
        RECT 103.555 150.970 103.785 151.790 ;
        RECT 103.955 150.990 104.285 151.620 ;
        RECT 102.075 150.550 102.425 150.800 ;
        RECT 103.535 150.550 103.865 150.800 ;
        RECT 97.150 150.090 97.320 150.210 ;
        RECT 98.420 150.090 98.740 150.380 ;
        RECT 96.635 149.240 96.915 150.040 ;
        RECT 97.150 149.920 98.740 150.090 ;
        RECT 97.085 149.460 98.740 149.750 ;
        RECT 98.915 149.410 99.255 150.380 ;
        RECT 99.425 149.240 99.595 150.380 ;
        RECT 99.785 150.210 102.220 150.380 ;
        RECT 99.865 149.240 100.115 150.040 ;
        RECT 100.760 149.410 101.090 150.210 ;
        RECT 101.390 149.240 101.720 150.040 ;
        RECT 101.890 149.410 102.220 150.210 ;
        RECT 102.595 149.240 102.885 150.405 ;
        RECT 104.035 150.390 104.285 150.990 ;
        RECT 104.455 150.970 104.665 151.790 ;
        RECT 104.900 151.080 105.155 151.610 ;
        RECT 105.325 151.330 105.630 151.790 ;
        RECT 105.875 151.410 106.945 151.580 ;
        RECT 103.555 149.240 103.785 150.380 ;
        RECT 103.955 149.410 104.285 150.390 ;
        RECT 104.900 150.430 105.110 151.080 ;
        RECT 105.875 151.055 106.195 151.410 ;
        RECT 105.870 150.880 106.195 151.055 ;
        RECT 105.280 150.580 106.195 150.880 ;
        RECT 106.365 150.840 106.605 151.240 ;
        RECT 106.775 151.180 106.945 151.410 ;
        RECT 107.115 151.350 107.305 151.790 ;
        RECT 107.475 151.340 108.425 151.620 ;
        RECT 108.645 151.430 108.995 151.600 ;
        RECT 106.775 151.010 107.305 151.180 ;
        RECT 105.280 150.550 106.020 150.580 ;
        RECT 104.455 149.240 104.665 150.380 ;
        RECT 104.900 149.550 105.155 150.430 ;
        RECT 105.325 149.240 105.630 150.380 ;
        RECT 105.850 149.960 106.020 150.550 ;
        RECT 106.365 150.470 106.905 150.840 ;
        RECT 107.085 150.730 107.305 151.010 ;
        RECT 107.475 150.560 107.645 151.340 ;
        RECT 107.240 150.390 107.645 150.560 ;
        RECT 107.815 150.550 108.165 151.170 ;
        RECT 107.240 150.300 107.410 150.390 ;
        RECT 108.335 150.380 108.545 151.170 ;
        RECT 106.190 150.130 107.410 150.300 ;
        RECT 107.870 150.220 108.545 150.380 ;
        RECT 105.850 149.790 106.650 149.960 ;
        RECT 105.970 149.240 106.300 149.620 ;
        RECT 106.480 149.500 106.650 149.790 ;
        RECT 107.240 149.750 107.410 150.130 ;
        RECT 107.580 150.210 108.545 150.220 ;
        RECT 108.735 151.040 108.995 151.430 ;
        RECT 109.205 151.330 109.535 151.790 ;
        RECT 110.410 151.400 111.265 151.570 ;
        RECT 111.470 151.400 111.965 151.570 ;
        RECT 112.135 151.430 112.465 151.790 ;
        RECT 108.735 150.350 108.905 151.040 ;
        RECT 109.075 150.690 109.245 150.870 ;
        RECT 109.415 150.860 110.205 151.110 ;
        RECT 110.410 150.690 110.580 151.400 ;
        RECT 110.750 150.890 111.105 151.110 ;
        RECT 109.075 150.520 110.765 150.690 ;
        RECT 107.580 149.920 108.040 150.210 ;
        RECT 108.735 150.180 110.235 150.350 ;
        RECT 108.735 150.040 108.905 150.180 ;
        RECT 108.345 149.870 108.905 150.040 ;
        RECT 106.820 149.240 107.070 149.700 ;
        RECT 107.240 149.410 108.110 149.750 ;
        RECT 108.345 149.410 108.515 149.870 ;
        RECT 109.350 149.840 110.425 150.010 ;
        RECT 108.685 149.240 109.055 149.700 ;
        RECT 109.350 149.500 109.520 149.840 ;
        RECT 109.690 149.240 110.020 149.670 ;
        RECT 110.255 149.500 110.425 149.840 ;
        RECT 110.595 149.740 110.765 150.520 ;
        RECT 110.935 150.300 111.105 150.890 ;
        RECT 111.275 150.490 111.625 151.110 ;
        RECT 110.935 149.910 111.400 150.300 ;
        RECT 111.795 150.040 111.965 151.400 ;
        RECT 112.135 150.210 112.595 151.260 ;
        RECT 111.570 149.870 111.965 150.040 ;
        RECT 111.570 149.740 111.740 149.870 ;
        RECT 110.595 149.410 111.275 149.740 ;
        RECT 111.490 149.410 111.740 149.740 ;
        RECT 111.910 149.240 112.160 149.700 ;
        RECT 112.330 149.425 112.655 150.210 ;
        RECT 112.825 149.410 112.995 151.530 ;
        RECT 113.165 151.410 113.495 151.790 ;
        RECT 113.665 151.240 113.920 151.530 ;
        RECT 113.170 151.070 113.920 151.240 ;
        RECT 113.170 150.080 113.400 151.070 ;
        RECT 114.555 151.040 115.765 151.790 ;
        RECT 113.570 150.250 113.920 150.900 ;
        RECT 114.555 150.330 115.075 150.870 ;
        RECT 115.245 150.500 115.765 151.040 ;
        RECT 113.170 149.910 113.920 150.080 ;
        RECT 113.165 149.240 113.495 149.740 ;
        RECT 113.665 149.410 113.920 149.910 ;
        RECT 114.555 149.240 115.765 150.330 ;
        RECT 10.510 149.070 115.850 149.240 ;
        RECT 10.595 147.980 11.805 149.070 ;
        RECT 10.595 147.270 11.115 147.810 ;
        RECT 11.285 147.440 11.805 147.980 ;
        RECT 12.435 147.905 12.725 149.070 ;
        RECT 13.270 148.090 13.525 148.760 ;
        RECT 13.705 148.270 13.990 149.070 ;
        RECT 14.170 148.350 14.500 148.860 ;
        RECT 13.270 148.050 13.450 148.090 ;
        RECT 13.185 147.880 13.450 148.050 ;
        RECT 10.595 146.520 11.805 147.270 ;
        RECT 12.435 146.520 12.725 147.245 ;
        RECT 13.270 147.230 13.450 147.880 ;
        RECT 14.170 147.760 14.420 148.350 ;
        RECT 14.770 148.200 14.940 148.810 ;
        RECT 15.110 148.380 15.440 149.070 ;
        RECT 15.670 148.520 15.910 148.810 ;
        RECT 16.110 148.690 16.530 149.070 ;
        RECT 16.710 148.600 17.340 148.850 ;
        RECT 17.810 148.690 18.140 149.070 ;
        RECT 16.710 148.520 16.880 148.600 ;
        RECT 18.310 148.520 18.480 148.810 ;
        RECT 18.660 148.690 19.040 149.070 ;
        RECT 19.280 148.685 20.110 148.855 ;
        RECT 15.670 148.350 16.880 148.520 ;
        RECT 13.620 147.430 14.420 147.760 ;
        RECT 13.270 146.700 13.525 147.230 ;
        RECT 13.705 146.520 13.990 146.980 ;
        RECT 14.170 146.780 14.420 147.430 ;
        RECT 14.620 148.180 14.940 148.200 ;
        RECT 14.620 148.010 16.540 148.180 ;
        RECT 14.620 147.115 14.810 148.010 ;
        RECT 16.710 147.840 16.880 148.350 ;
        RECT 17.050 148.090 17.570 148.400 ;
        RECT 14.980 147.670 16.880 147.840 ;
        RECT 14.980 147.610 15.310 147.670 ;
        RECT 15.460 147.440 15.790 147.500 ;
        RECT 15.130 147.170 15.790 147.440 ;
        RECT 14.620 146.785 14.940 147.115 ;
        RECT 15.120 146.520 15.780 147.000 ;
        RECT 15.980 146.910 16.150 147.670 ;
        RECT 17.050 147.500 17.230 147.910 ;
        RECT 16.320 147.330 16.650 147.450 ;
        RECT 17.400 147.330 17.570 148.090 ;
        RECT 16.320 147.160 17.570 147.330 ;
        RECT 17.740 148.270 19.110 148.520 ;
        RECT 17.740 147.500 17.930 148.270 ;
        RECT 18.860 148.010 19.110 148.270 ;
        RECT 18.100 147.840 18.350 148.000 ;
        RECT 19.280 147.840 19.450 148.685 ;
        RECT 20.345 148.400 20.515 148.900 ;
        RECT 20.685 148.570 21.015 149.070 ;
        RECT 19.620 148.010 20.120 148.390 ;
        RECT 20.345 148.230 21.040 148.400 ;
        RECT 18.100 147.670 19.450 147.840 ;
        RECT 19.030 147.630 19.450 147.670 ;
        RECT 17.740 147.160 18.160 147.500 ;
        RECT 18.450 147.170 18.860 147.500 ;
        RECT 15.980 146.740 16.830 146.910 ;
        RECT 17.390 146.520 17.710 146.980 ;
        RECT 17.910 146.730 18.160 147.160 ;
        RECT 18.450 146.520 18.860 146.960 ;
        RECT 19.030 146.900 19.200 147.630 ;
        RECT 19.370 147.080 19.720 147.450 ;
        RECT 19.900 147.140 20.120 148.010 ;
        RECT 20.290 147.440 20.700 148.060 ;
        RECT 20.870 147.260 21.040 148.230 ;
        RECT 20.345 147.070 21.040 147.260 ;
        RECT 19.030 146.700 20.045 146.900 ;
        RECT 20.345 146.740 20.515 147.070 ;
        RECT 20.685 146.520 21.015 146.900 ;
        RECT 21.230 146.780 21.455 148.900 ;
        RECT 21.625 148.570 21.955 149.070 ;
        RECT 22.125 148.400 22.295 148.900 ;
        RECT 21.630 148.230 22.295 148.400 ;
        RECT 21.630 147.240 21.860 148.230 ;
        RECT 22.030 147.410 22.380 148.060 ;
        RECT 22.555 147.980 23.765 149.070 ;
        RECT 22.555 147.440 23.075 147.980 ;
        RECT 23.940 147.930 24.275 148.900 ;
        RECT 24.445 147.930 24.615 149.070 ;
        RECT 24.785 148.730 26.815 148.900 ;
        RECT 23.245 147.270 23.765 147.810 ;
        RECT 21.630 147.070 22.295 147.240 ;
        RECT 21.625 146.520 21.955 146.900 ;
        RECT 22.125 146.780 22.295 147.070 ;
        RECT 22.555 146.520 23.765 147.270 ;
        RECT 23.940 147.260 24.110 147.930 ;
        RECT 24.785 147.760 24.955 148.730 ;
        RECT 24.280 147.430 24.535 147.760 ;
        RECT 24.760 147.430 24.955 147.760 ;
        RECT 25.125 148.390 26.250 148.560 ;
        RECT 24.365 147.260 24.535 147.430 ;
        RECT 25.125 147.260 25.295 148.390 ;
        RECT 23.940 146.690 24.195 147.260 ;
        RECT 24.365 147.090 25.295 147.260 ;
        RECT 25.465 148.050 26.475 148.220 ;
        RECT 25.465 147.250 25.635 148.050 ;
        RECT 25.840 147.710 26.115 147.850 ;
        RECT 25.835 147.540 26.115 147.710 ;
        RECT 25.120 147.055 25.295 147.090 ;
        RECT 24.365 146.520 24.695 146.920 ;
        RECT 25.120 146.690 25.650 147.055 ;
        RECT 25.840 146.690 26.115 147.540 ;
        RECT 26.285 146.690 26.475 148.050 ;
        RECT 26.645 148.065 26.815 148.730 ;
        RECT 26.985 148.310 27.155 149.070 ;
        RECT 27.390 148.310 27.905 148.720 ;
        RECT 26.645 147.875 27.395 148.065 ;
        RECT 27.565 147.500 27.905 148.310 ;
        RECT 29.085 148.140 29.255 148.900 ;
        RECT 29.435 148.310 29.765 149.070 ;
        RECT 29.085 147.970 29.750 148.140 ;
        RECT 29.935 147.995 30.205 148.900 ;
        RECT 29.580 147.825 29.750 147.970 ;
        RECT 26.675 147.330 27.905 147.500 ;
        RECT 29.015 147.420 29.345 147.790 ;
        RECT 29.580 147.495 29.865 147.825 ;
        RECT 26.655 146.520 27.165 147.055 ;
        RECT 27.385 146.725 27.630 147.330 ;
        RECT 29.580 147.240 29.750 147.495 ;
        RECT 29.085 147.070 29.750 147.240 ;
        RECT 30.035 147.195 30.205 147.995 ;
        RECT 30.580 148.100 30.910 148.900 ;
        RECT 31.080 148.270 31.410 149.070 ;
        RECT 31.710 148.100 32.040 148.900 ;
        RECT 32.685 148.270 32.935 149.070 ;
        RECT 30.580 147.930 33.015 148.100 ;
        RECT 33.205 147.930 33.375 149.070 ;
        RECT 33.545 147.930 33.885 148.900 ;
        RECT 30.375 147.510 30.725 147.760 ;
        RECT 30.910 147.300 31.080 147.930 ;
        RECT 31.250 147.510 31.580 147.710 ;
        RECT 31.750 147.510 32.080 147.710 ;
        RECT 32.250 147.510 32.670 147.710 ;
        RECT 32.845 147.680 33.015 147.930 ;
        RECT 32.845 147.510 33.540 147.680 ;
        RECT 29.085 146.690 29.255 147.070 ;
        RECT 29.435 146.520 29.765 146.900 ;
        RECT 29.945 146.690 30.205 147.195 ;
        RECT 30.580 146.690 31.080 147.300 ;
        RECT 31.710 147.170 32.935 147.340 ;
        RECT 33.710 147.320 33.885 147.930 ;
        RECT 34.055 147.980 36.645 149.070 ;
        RECT 34.055 147.460 35.265 147.980 ;
        RECT 36.855 147.930 37.085 149.070 ;
        RECT 37.255 147.920 37.585 148.900 ;
        RECT 37.755 147.930 37.965 149.070 ;
        RECT 31.710 146.690 32.040 147.170 ;
        RECT 32.210 146.520 32.435 146.980 ;
        RECT 32.605 146.690 32.935 147.170 ;
        RECT 33.125 146.520 33.375 147.320 ;
        RECT 33.545 146.690 33.885 147.320 ;
        RECT 35.435 147.290 36.645 147.810 ;
        RECT 36.835 147.510 37.165 147.760 ;
        RECT 34.055 146.520 36.645 147.290 ;
        RECT 36.855 146.520 37.085 147.340 ;
        RECT 37.335 147.320 37.585 147.920 ;
        RECT 38.195 147.905 38.485 149.070 ;
        RECT 38.655 147.980 41.245 149.070 ;
        RECT 41.420 148.560 43.075 148.850 ;
        RECT 41.420 148.220 43.010 148.390 ;
        RECT 43.245 148.270 43.525 149.070 ;
        RECT 38.655 147.460 39.865 147.980 ;
        RECT 41.420 147.930 41.740 148.220 ;
        RECT 42.840 148.100 43.010 148.220 ;
        RECT 41.935 147.880 42.650 148.050 ;
        RECT 42.840 147.930 43.565 148.100 ;
        RECT 43.735 147.930 44.005 148.900 ;
        RECT 37.255 146.690 37.585 147.320 ;
        RECT 37.755 146.520 37.965 147.340 ;
        RECT 40.035 147.290 41.245 147.810 ;
        RECT 38.195 146.520 38.485 147.245 ;
        RECT 38.655 146.520 41.245 147.290 ;
        RECT 41.420 147.190 41.770 147.760 ;
        RECT 41.940 147.430 42.650 147.880 ;
        RECT 43.395 147.760 43.565 147.930 ;
        RECT 42.820 147.430 43.225 147.760 ;
        RECT 43.395 147.430 43.665 147.760 ;
        RECT 43.395 147.260 43.565 147.430 ;
        RECT 41.955 147.090 43.565 147.260 ;
        RECT 43.835 147.195 44.005 147.930 ;
        RECT 41.425 146.520 41.755 147.020 ;
        RECT 41.955 146.740 42.125 147.090 ;
        RECT 42.325 146.520 42.655 146.920 ;
        RECT 42.825 146.740 42.995 147.090 ;
        RECT 43.165 146.520 43.545 146.920 ;
        RECT 43.735 146.850 44.005 147.195 ;
        RECT 44.175 147.930 44.515 148.900 ;
        RECT 44.685 147.930 44.855 149.070 ;
        RECT 45.125 148.270 45.375 149.070 ;
        RECT 46.020 148.100 46.350 148.900 ;
        RECT 46.650 148.270 46.980 149.070 ;
        RECT 47.150 148.100 47.480 148.900 ;
        RECT 45.045 147.930 47.480 148.100 ;
        RECT 48.775 147.930 49.115 148.900 ;
        RECT 49.285 147.930 49.455 149.070 ;
        RECT 49.725 148.270 49.975 149.070 ;
        RECT 50.620 148.100 50.950 148.900 ;
        RECT 51.250 148.270 51.580 149.070 ;
        RECT 51.750 148.100 52.080 148.900 ;
        RECT 49.645 147.930 52.080 148.100 ;
        RECT 53.750 148.090 54.005 148.760 ;
        RECT 54.185 148.270 54.470 149.070 ;
        RECT 54.650 148.350 54.980 148.860 ;
        RECT 53.750 148.050 53.930 148.090 ;
        RECT 44.175 147.320 44.350 147.930 ;
        RECT 45.045 147.680 45.215 147.930 ;
        RECT 44.520 147.510 45.215 147.680 ;
        RECT 45.390 147.510 45.810 147.710 ;
        RECT 45.980 147.510 46.310 147.710 ;
        RECT 46.480 147.510 46.810 147.710 ;
        RECT 44.175 146.690 44.515 147.320 ;
        RECT 44.685 146.520 44.935 147.320 ;
        RECT 45.125 147.170 46.350 147.340 ;
        RECT 45.125 146.690 45.455 147.170 ;
        RECT 45.625 146.520 45.850 146.980 ;
        RECT 46.020 146.690 46.350 147.170 ;
        RECT 46.980 147.300 47.150 147.930 ;
        RECT 47.335 147.510 47.685 147.760 ;
        RECT 48.775 147.370 48.950 147.930 ;
        RECT 49.645 147.680 49.815 147.930 ;
        RECT 49.120 147.510 49.815 147.680 ;
        RECT 49.990 147.510 50.410 147.710 ;
        RECT 50.580 147.510 50.910 147.710 ;
        RECT 51.080 147.510 51.410 147.710 ;
        RECT 48.775 147.320 49.005 147.370 ;
        RECT 46.980 146.690 47.480 147.300 ;
        RECT 48.775 146.690 49.115 147.320 ;
        RECT 49.285 146.520 49.535 147.320 ;
        RECT 49.725 147.170 50.950 147.340 ;
        RECT 49.725 146.690 50.055 147.170 ;
        RECT 50.225 146.520 50.450 146.980 ;
        RECT 50.620 146.690 50.950 147.170 ;
        RECT 51.580 147.300 51.750 147.930 ;
        RECT 53.665 147.880 53.930 148.050 ;
        RECT 51.935 147.510 52.285 147.760 ;
        RECT 51.580 146.690 52.080 147.300 ;
        RECT 53.750 147.230 53.930 147.880 ;
        RECT 54.650 147.760 54.900 148.350 ;
        RECT 55.250 148.200 55.420 148.810 ;
        RECT 55.590 148.380 55.920 149.070 ;
        RECT 56.150 148.520 56.390 148.810 ;
        RECT 56.590 148.690 57.010 149.070 ;
        RECT 57.190 148.600 57.820 148.850 ;
        RECT 58.290 148.690 58.620 149.070 ;
        RECT 57.190 148.520 57.360 148.600 ;
        RECT 58.790 148.520 58.960 148.810 ;
        RECT 59.140 148.690 59.520 149.070 ;
        RECT 59.760 148.685 60.590 148.855 ;
        RECT 56.150 148.350 57.360 148.520 ;
        RECT 54.100 147.430 54.900 147.760 ;
        RECT 53.750 146.700 54.005 147.230 ;
        RECT 54.185 146.520 54.470 146.980 ;
        RECT 54.650 146.780 54.900 147.430 ;
        RECT 55.100 148.180 55.420 148.200 ;
        RECT 55.100 148.010 57.020 148.180 ;
        RECT 55.100 147.115 55.290 148.010 ;
        RECT 57.190 147.840 57.360 148.350 ;
        RECT 57.530 148.090 58.050 148.400 ;
        RECT 55.460 147.670 57.360 147.840 ;
        RECT 55.460 147.610 55.790 147.670 ;
        RECT 55.940 147.440 56.270 147.500 ;
        RECT 55.610 147.170 56.270 147.440 ;
        RECT 55.100 146.785 55.420 147.115 ;
        RECT 55.600 146.520 56.260 147.000 ;
        RECT 56.460 146.910 56.630 147.670 ;
        RECT 57.530 147.500 57.710 147.910 ;
        RECT 56.800 147.330 57.130 147.450 ;
        RECT 57.880 147.330 58.050 148.090 ;
        RECT 56.800 147.160 58.050 147.330 ;
        RECT 58.220 148.270 59.590 148.520 ;
        RECT 58.220 147.500 58.410 148.270 ;
        RECT 59.340 148.010 59.590 148.270 ;
        RECT 58.580 147.840 58.830 148.000 ;
        RECT 59.760 147.840 59.930 148.685 ;
        RECT 60.825 148.400 60.995 148.900 ;
        RECT 61.165 148.570 61.495 149.070 ;
        RECT 60.100 148.010 60.600 148.390 ;
        RECT 60.825 148.230 61.520 148.400 ;
        RECT 58.580 147.670 59.930 147.840 ;
        RECT 59.510 147.630 59.930 147.670 ;
        RECT 58.220 147.160 58.640 147.500 ;
        RECT 58.930 147.170 59.340 147.500 ;
        RECT 56.460 146.740 57.310 146.910 ;
        RECT 57.870 146.520 58.190 146.980 ;
        RECT 58.390 146.730 58.640 147.160 ;
        RECT 58.930 146.520 59.340 146.960 ;
        RECT 59.510 146.900 59.680 147.630 ;
        RECT 59.850 147.080 60.200 147.450 ;
        RECT 60.380 147.140 60.600 148.010 ;
        RECT 60.770 147.440 61.180 148.060 ;
        RECT 61.350 147.260 61.520 148.230 ;
        RECT 60.825 147.070 61.520 147.260 ;
        RECT 59.510 146.700 60.525 146.900 ;
        RECT 60.825 146.740 60.995 147.070 ;
        RECT 61.165 146.520 61.495 146.900 ;
        RECT 61.710 146.780 61.935 148.900 ;
        RECT 62.105 148.570 62.435 149.070 ;
        RECT 62.605 148.400 62.775 148.900 ;
        RECT 62.110 148.230 62.775 148.400 ;
        RECT 62.110 147.240 62.340 148.230 ;
        RECT 62.510 147.410 62.860 148.060 ;
        RECT 63.955 147.905 64.245 149.070 ;
        RECT 64.415 147.930 64.685 148.900 ;
        RECT 64.895 148.270 65.175 149.070 ;
        RECT 65.345 148.560 67.000 148.850 ;
        RECT 65.410 148.220 67.000 148.390 ;
        RECT 65.410 148.100 65.580 148.220 ;
        RECT 64.855 147.930 65.580 148.100 ;
        RECT 62.110 147.070 62.775 147.240 ;
        RECT 62.105 146.520 62.435 146.900 ;
        RECT 62.605 146.780 62.775 147.070 ;
        RECT 63.955 146.520 64.245 147.245 ;
        RECT 64.415 147.195 64.585 147.930 ;
        RECT 64.855 147.760 65.025 147.930 ;
        RECT 64.755 147.430 65.025 147.760 ;
        RECT 65.195 147.430 65.600 147.760 ;
        RECT 65.770 147.430 66.480 148.050 ;
        RECT 66.680 147.930 67.000 148.220 ;
        RECT 67.380 148.100 67.710 148.900 ;
        RECT 67.880 148.270 68.210 149.070 ;
        RECT 68.510 148.100 68.840 148.900 ;
        RECT 69.485 148.270 69.735 149.070 ;
        RECT 67.380 147.930 69.815 148.100 ;
        RECT 70.005 147.930 70.175 149.070 ;
        RECT 70.345 147.930 70.685 148.900 ;
        RECT 64.855 147.260 65.025 147.430 ;
        RECT 64.415 146.850 64.685 147.195 ;
        RECT 64.855 147.090 66.465 147.260 ;
        RECT 66.650 147.190 67.000 147.760 ;
        RECT 67.175 147.510 67.525 147.760 ;
        RECT 67.710 147.300 67.880 147.930 ;
        RECT 68.050 147.510 68.380 147.710 ;
        RECT 68.550 147.510 68.880 147.710 ;
        RECT 69.050 147.510 69.470 147.710 ;
        RECT 69.645 147.680 69.815 147.930 ;
        RECT 69.645 147.510 70.340 147.680 ;
        RECT 64.875 146.520 65.255 146.920 ;
        RECT 65.425 146.740 65.595 147.090 ;
        RECT 65.765 146.520 66.095 146.920 ;
        RECT 66.295 146.740 66.465 147.090 ;
        RECT 66.665 146.520 66.995 147.020 ;
        RECT 67.380 146.690 67.880 147.300 ;
        RECT 68.510 147.170 69.735 147.340 ;
        RECT 70.510 147.320 70.685 147.930 ;
        RECT 68.510 146.690 68.840 147.170 ;
        RECT 69.010 146.520 69.235 146.980 ;
        RECT 69.405 146.690 69.735 147.170 ;
        RECT 69.925 146.520 70.175 147.320 ;
        RECT 70.345 146.690 70.685 147.320 ;
        RECT 70.855 147.930 71.195 148.900 ;
        RECT 71.365 147.930 71.535 149.070 ;
        RECT 71.805 148.270 72.055 149.070 ;
        RECT 72.700 148.100 73.030 148.900 ;
        RECT 73.330 148.270 73.660 149.070 ;
        RECT 73.830 148.100 74.160 148.900 ;
        RECT 71.725 147.930 74.160 148.100 ;
        RECT 74.625 148.140 74.795 148.900 ;
        RECT 74.975 148.310 75.305 149.070 ;
        RECT 74.625 147.970 75.290 148.140 ;
        RECT 75.475 147.995 75.745 148.900 ;
        RECT 76.005 148.400 76.175 148.900 ;
        RECT 76.345 148.570 76.675 149.070 ;
        RECT 76.005 148.230 76.670 148.400 ;
        RECT 70.855 147.370 71.030 147.930 ;
        RECT 71.725 147.680 71.895 147.930 ;
        RECT 71.200 147.510 71.895 147.680 ;
        RECT 72.070 147.510 72.490 147.710 ;
        RECT 72.660 147.510 72.990 147.710 ;
        RECT 73.160 147.510 73.490 147.710 ;
        RECT 70.855 147.320 71.085 147.370 ;
        RECT 70.855 146.690 71.195 147.320 ;
        RECT 71.365 146.520 71.615 147.320 ;
        RECT 71.805 147.170 73.030 147.340 ;
        RECT 71.805 146.690 72.135 147.170 ;
        RECT 72.305 146.520 72.530 146.980 ;
        RECT 72.700 146.690 73.030 147.170 ;
        RECT 73.660 147.300 73.830 147.930 ;
        RECT 75.120 147.825 75.290 147.970 ;
        RECT 74.015 147.510 74.365 147.760 ;
        RECT 74.555 147.420 74.885 147.790 ;
        RECT 75.120 147.495 75.405 147.825 ;
        RECT 73.660 146.690 74.160 147.300 ;
        RECT 75.120 147.240 75.290 147.495 ;
        RECT 74.625 147.070 75.290 147.240 ;
        RECT 75.575 147.195 75.745 147.995 ;
        RECT 75.920 147.410 76.270 148.060 ;
        RECT 76.440 147.240 76.670 148.230 ;
        RECT 74.625 146.690 74.795 147.070 ;
        RECT 74.975 146.520 75.305 146.900 ;
        RECT 75.485 146.690 75.745 147.195 ;
        RECT 76.005 147.070 76.670 147.240 ;
        RECT 76.005 146.780 76.175 147.070 ;
        RECT 76.345 146.520 76.675 146.900 ;
        RECT 76.845 146.780 77.070 148.900 ;
        RECT 77.285 148.570 77.615 149.070 ;
        RECT 77.785 148.400 77.955 148.900 ;
        RECT 78.190 148.685 79.020 148.855 ;
        RECT 79.260 148.690 79.640 149.070 ;
        RECT 77.260 148.230 77.955 148.400 ;
        RECT 77.260 147.260 77.430 148.230 ;
        RECT 77.600 147.440 78.010 148.060 ;
        RECT 78.180 148.010 78.680 148.390 ;
        RECT 77.260 147.070 77.955 147.260 ;
        RECT 78.180 147.140 78.400 148.010 ;
        RECT 78.850 147.840 79.020 148.685 ;
        RECT 79.820 148.520 79.990 148.810 ;
        RECT 80.160 148.690 80.490 149.070 ;
        RECT 80.960 148.600 81.590 148.850 ;
        RECT 81.770 148.690 82.190 149.070 ;
        RECT 81.420 148.520 81.590 148.600 ;
        RECT 82.390 148.520 82.630 148.810 ;
        RECT 79.190 148.270 80.560 148.520 ;
        RECT 79.190 148.010 79.440 148.270 ;
        RECT 79.950 147.840 80.200 148.000 ;
        RECT 78.850 147.670 80.200 147.840 ;
        RECT 78.850 147.630 79.270 147.670 ;
        RECT 78.580 147.080 78.930 147.450 ;
        RECT 77.285 146.520 77.615 146.900 ;
        RECT 77.785 146.740 77.955 147.070 ;
        RECT 79.100 146.900 79.270 147.630 ;
        RECT 80.370 147.500 80.560 148.270 ;
        RECT 79.440 147.170 79.850 147.500 ;
        RECT 80.140 147.160 80.560 147.500 ;
        RECT 80.730 148.090 81.250 148.400 ;
        RECT 81.420 148.350 82.630 148.520 ;
        RECT 82.860 148.380 83.190 149.070 ;
        RECT 80.730 147.330 80.900 148.090 ;
        RECT 81.070 147.500 81.250 147.910 ;
        RECT 81.420 147.840 81.590 148.350 ;
        RECT 83.360 148.200 83.530 148.810 ;
        RECT 83.800 148.350 84.130 148.860 ;
        RECT 83.360 148.180 83.680 148.200 ;
        RECT 81.760 148.010 83.680 148.180 ;
        RECT 81.420 147.670 83.320 147.840 ;
        RECT 81.650 147.330 81.980 147.450 ;
        RECT 80.730 147.160 81.980 147.330 ;
        RECT 78.255 146.700 79.270 146.900 ;
        RECT 79.440 146.520 79.850 146.960 ;
        RECT 80.140 146.730 80.390 147.160 ;
        RECT 80.590 146.520 80.910 146.980 ;
        RECT 82.150 146.910 82.320 147.670 ;
        RECT 82.990 147.610 83.320 147.670 ;
        RECT 82.510 147.440 82.840 147.500 ;
        RECT 82.510 147.170 83.170 147.440 ;
        RECT 83.490 147.115 83.680 148.010 ;
        RECT 81.470 146.740 82.320 146.910 ;
        RECT 82.520 146.520 83.180 147.000 ;
        RECT 83.360 146.785 83.680 147.115 ;
        RECT 83.880 147.760 84.130 148.350 ;
        RECT 84.310 148.270 84.595 149.070 ;
        RECT 84.775 148.090 85.030 148.760 ;
        RECT 83.880 147.430 84.680 147.760 ;
        RECT 83.880 146.780 84.130 147.430 ;
        RECT 84.850 147.230 85.030 148.090 ;
        RECT 85.575 148.310 86.090 148.720 ;
        RECT 86.325 148.310 86.495 149.070 ;
        RECT 86.665 148.730 88.695 148.900 ;
        RECT 85.575 147.500 85.915 148.310 ;
        RECT 86.665 148.065 86.835 148.730 ;
        RECT 87.230 148.390 88.355 148.560 ;
        RECT 86.085 147.875 86.835 148.065 ;
        RECT 87.005 148.050 88.015 148.220 ;
        RECT 85.575 147.330 86.805 147.500 ;
        RECT 84.775 147.030 85.030 147.230 ;
        RECT 84.310 146.520 84.595 146.980 ;
        RECT 84.775 146.860 85.115 147.030 ;
        RECT 84.775 146.700 85.030 146.860 ;
        RECT 85.850 146.725 86.095 147.330 ;
        RECT 86.315 146.520 86.825 147.055 ;
        RECT 87.005 146.690 87.195 148.050 ;
        RECT 87.365 147.710 87.640 147.850 ;
        RECT 87.365 147.540 87.645 147.710 ;
        RECT 87.365 146.690 87.640 147.540 ;
        RECT 87.845 147.250 88.015 148.050 ;
        RECT 88.185 147.260 88.355 148.390 ;
        RECT 88.525 147.760 88.695 148.730 ;
        RECT 88.865 147.930 89.035 149.070 ;
        RECT 89.205 147.930 89.540 148.900 ;
        RECT 88.525 147.430 88.720 147.760 ;
        RECT 88.945 147.430 89.200 147.760 ;
        RECT 88.945 147.260 89.115 147.430 ;
        RECT 89.370 147.260 89.540 147.930 ;
        RECT 89.715 147.905 90.005 149.070 ;
        RECT 90.175 147.980 91.845 149.070 ;
        RECT 92.105 148.140 92.275 148.900 ;
        RECT 92.455 148.310 92.785 149.070 ;
        RECT 90.175 147.460 90.925 147.980 ;
        RECT 92.105 147.970 92.770 148.140 ;
        RECT 92.955 147.995 93.225 148.900 ;
        RECT 92.600 147.825 92.770 147.970 ;
        RECT 91.095 147.290 91.845 147.810 ;
        RECT 92.035 147.420 92.365 147.790 ;
        RECT 92.600 147.495 92.885 147.825 ;
        RECT 88.185 147.090 89.115 147.260 ;
        RECT 88.185 147.055 88.360 147.090 ;
        RECT 87.830 146.690 88.360 147.055 ;
        RECT 88.785 146.520 89.115 146.920 ;
        RECT 89.285 146.690 89.540 147.260 ;
        RECT 89.715 146.520 90.005 147.245 ;
        RECT 90.175 146.520 91.845 147.290 ;
        RECT 92.600 147.240 92.770 147.495 ;
        RECT 92.105 147.070 92.770 147.240 ;
        RECT 93.055 147.195 93.225 147.995 ;
        RECT 92.105 146.690 92.275 147.070 ;
        RECT 92.455 146.520 92.785 146.900 ;
        RECT 92.965 146.690 93.225 147.195 ;
        RECT 94.315 147.930 94.585 148.900 ;
        RECT 94.795 148.270 95.075 149.070 ;
        RECT 95.245 148.560 96.900 148.850 ;
        RECT 95.310 148.220 96.900 148.390 ;
        RECT 95.310 148.100 95.480 148.220 ;
        RECT 94.755 147.930 95.480 148.100 ;
        RECT 94.315 147.195 94.485 147.930 ;
        RECT 94.755 147.760 94.925 147.930 ;
        RECT 95.670 147.880 96.385 148.050 ;
        RECT 96.580 147.930 96.900 148.220 ;
        RECT 97.075 147.930 97.415 148.900 ;
        RECT 97.585 147.930 97.755 149.070 ;
        RECT 98.025 148.270 98.275 149.070 ;
        RECT 98.920 148.100 99.250 148.900 ;
        RECT 99.550 148.270 99.880 149.070 ;
        RECT 100.050 148.100 100.380 148.900 ;
        RECT 97.945 147.930 100.380 148.100 ;
        RECT 100.755 148.310 101.270 148.720 ;
        RECT 101.505 148.310 101.675 149.070 ;
        RECT 101.845 148.730 103.875 148.900 ;
        RECT 94.655 147.430 94.925 147.760 ;
        RECT 95.095 147.430 95.500 147.760 ;
        RECT 95.670 147.430 96.380 147.880 ;
        RECT 94.755 147.260 94.925 147.430 ;
        RECT 94.315 146.850 94.585 147.195 ;
        RECT 94.755 147.090 96.365 147.260 ;
        RECT 96.550 147.190 96.900 147.760 ;
        RECT 97.075 147.370 97.250 147.930 ;
        RECT 97.945 147.680 98.115 147.930 ;
        RECT 97.420 147.510 98.115 147.680 ;
        RECT 98.290 147.510 98.710 147.710 ;
        RECT 98.880 147.510 99.210 147.710 ;
        RECT 99.380 147.510 99.710 147.710 ;
        RECT 97.075 147.320 97.305 147.370 ;
        RECT 94.775 146.520 95.155 146.920 ;
        RECT 95.325 146.740 95.495 147.090 ;
        RECT 95.665 146.520 95.995 146.920 ;
        RECT 96.195 146.740 96.365 147.090 ;
        RECT 96.565 146.520 96.895 147.020 ;
        RECT 97.075 146.690 97.415 147.320 ;
        RECT 97.585 146.520 97.835 147.320 ;
        RECT 98.025 147.170 99.250 147.340 ;
        RECT 98.025 146.690 98.355 147.170 ;
        RECT 98.525 146.520 98.750 146.980 ;
        RECT 98.920 146.690 99.250 147.170 ;
        RECT 99.880 147.300 100.050 147.930 ;
        RECT 100.235 147.510 100.585 147.760 ;
        RECT 100.755 147.500 101.095 148.310 ;
        RECT 101.845 148.065 102.015 148.730 ;
        RECT 102.410 148.390 103.535 148.560 ;
        RECT 101.265 147.875 102.015 148.065 ;
        RECT 102.185 148.050 103.195 148.220 ;
        RECT 100.755 147.330 101.985 147.500 ;
        RECT 99.880 146.690 100.380 147.300 ;
        RECT 101.030 146.725 101.275 147.330 ;
        RECT 101.495 146.520 102.005 147.055 ;
        RECT 102.185 146.690 102.375 148.050 ;
        RECT 102.545 147.370 102.820 147.850 ;
        RECT 102.545 147.200 102.825 147.370 ;
        RECT 103.025 147.250 103.195 148.050 ;
        RECT 103.365 147.260 103.535 148.390 ;
        RECT 103.705 147.760 103.875 148.730 ;
        RECT 104.045 147.930 104.215 149.070 ;
        RECT 104.385 147.930 104.720 148.900 ;
        RECT 103.705 147.430 103.900 147.760 ;
        RECT 104.125 147.430 104.380 147.760 ;
        RECT 104.125 147.260 104.295 147.430 ;
        RECT 104.550 147.260 104.720 147.930 ;
        RECT 105.270 148.090 105.525 148.760 ;
        RECT 105.705 148.270 105.990 149.070 ;
        RECT 106.170 148.350 106.500 148.860 ;
        RECT 105.270 147.370 105.450 148.090 ;
        RECT 106.170 147.760 106.420 148.350 ;
        RECT 106.770 148.200 106.940 148.810 ;
        RECT 107.110 148.380 107.440 149.070 ;
        RECT 107.670 148.520 107.910 148.810 ;
        RECT 108.110 148.690 108.530 149.070 ;
        RECT 108.710 148.600 109.340 148.850 ;
        RECT 109.810 148.690 110.140 149.070 ;
        RECT 108.710 148.520 108.880 148.600 ;
        RECT 110.310 148.520 110.480 148.810 ;
        RECT 110.660 148.690 111.040 149.070 ;
        RECT 111.280 148.685 112.110 148.855 ;
        RECT 107.670 148.350 108.880 148.520 ;
        RECT 105.620 147.430 106.420 147.760 ;
        RECT 102.545 146.690 102.820 147.200 ;
        RECT 103.365 147.090 104.295 147.260 ;
        RECT 103.365 147.055 103.540 147.090 ;
        RECT 103.010 146.690 103.540 147.055 ;
        RECT 103.965 146.520 104.295 146.920 ;
        RECT 104.465 146.690 104.720 147.260 ;
        RECT 105.185 147.230 105.450 147.370 ;
        RECT 105.185 147.200 105.525 147.230 ;
        RECT 105.270 146.700 105.525 147.200 ;
        RECT 105.705 146.520 105.990 146.980 ;
        RECT 106.170 146.780 106.420 147.430 ;
        RECT 106.620 148.180 106.940 148.200 ;
        RECT 106.620 148.010 108.540 148.180 ;
        RECT 106.620 147.115 106.810 148.010 ;
        RECT 108.710 147.840 108.880 148.350 ;
        RECT 109.050 148.090 109.570 148.400 ;
        RECT 106.980 147.670 108.880 147.840 ;
        RECT 106.980 147.610 107.310 147.670 ;
        RECT 107.460 147.440 107.790 147.500 ;
        RECT 107.130 147.170 107.790 147.440 ;
        RECT 106.620 146.785 106.940 147.115 ;
        RECT 107.120 146.520 107.780 147.000 ;
        RECT 107.980 146.910 108.150 147.670 ;
        RECT 109.050 147.500 109.230 147.910 ;
        RECT 108.320 147.330 108.650 147.450 ;
        RECT 109.400 147.330 109.570 148.090 ;
        RECT 108.320 147.160 109.570 147.330 ;
        RECT 109.740 148.270 111.110 148.520 ;
        RECT 109.740 147.500 109.930 148.270 ;
        RECT 110.860 148.010 111.110 148.270 ;
        RECT 110.100 147.840 110.350 148.000 ;
        RECT 111.280 147.840 111.450 148.685 ;
        RECT 112.345 148.400 112.515 148.900 ;
        RECT 112.685 148.570 113.015 149.070 ;
        RECT 111.620 148.010 112.120 148.390 ;
        RECT 112.345 148.230 113.040 148.400 ;
        RECT 110.100 147.670 111.450 147.840 ;
        RECT 111.030 147.630 111.450 147.670 ;
        RECT 109.740 147.160 110.160 147.500 ;
        RECT 110.450 147.170 110.860 147.500 ;
        RECT 107.980 146.740 108.830 146.910 ;
        RECT 109.390 146.520 109.710 146.980 ;
        RECT 109.910 146.730 110.160 147.160 ;
        RECT 110.450 146.520 110.860 146.960 ;
        RECT 111.030 146.900 111.200 147.630 ;
        RECT 111.370 147.080 111.720 147.450 ;
        RECT 111.900 147.140 112.120 148.010 ;
        RECT 112.290 147.440 112.700 148.060 ;
        RECT 112.870 147.260 113.040 148.230 ;
        RECT 112.345 147.070 113.040 147.260 ;
        RECT 111.030 146.700 112.045 146.900 ;
        RECT 112.345 146.740 112.515 147.070 ;
        RECT 112.685 146.520 113.015 146.900 ;
        RECT 113.230 146.780 113.455 148.900 ;
        RECT 113.625 148.570 113.955 149.070 ;
        RECT 114.125 148.400 114.295 148.900 ;
        RECT 113.630 148.230 114.295 148.400 ;
        RECT 113.630 147.240 113.860 148.230 ;
        RECT 114.030 147.410 114.380 148.060 ;
        RECT 114.555 147.980 115.765 149.070 ;
        RECT 114.555 147.440 115.075 147.980 ;
        RECT 115.245 147.270 115.765 147.810 ;
        RECT 113.630 147.070 114.295 147.240 ;
        RECT 113.625 146.520 113.955 146.900 ;
        RECT 114.125 146.780 114.295 147.070 ;
        RECT 114.555 146.520 115.765 147.270 ;
        RECT 10.510 146.350 115.850 146.520 ;
        RECT 10.595 145.600 11.805 146.350 ;
        RECT 10.595 145.060 11.115 145.600 ;
        RECT 12.435 145.580 14.105 146.350 ;
        RECT 11.285 144.890 11.805 145.430 ;
        RECT 10.595 143.800 11.805 144.890 ;
        RECT 12.435 144.890 13.185 145.410 ;
        RECT 13.355 145.060 14.105 145.580 ;
        RECT 14.335 145.530 14.545 146.350 ;
        RECT 14.715 145.550 15.045 146.180 ;
        RECT 14.715 144.950 14.965 145.550 ;
        RECT 15.215 145.530 15.445 146.350 ;
        RECT 16.030 145.640 16.285 146.170 ;
        RECT 16.465 145.890 16.750 146.350 ;
        RECT 15.135 145.110 15.465 145.360 ;
        RECT 16.030 144.990 16.210 145.640 ;
        RECT 16.930 145.440 17.180 146.090 ;
        RECT 16.380 145.110 17.180 145.440 ;
        RECT 12.435 143.800 14.105 144.890 ;
        RECT 14.335 143.800 14.545 144.940 ;
        RECT 14.715 143.970 15.045 144.950 ;
        RECT 15.215 143.800 15.445 144.940 ;
        RECT 15.945 144.820 16.210 144.990 ;
        RECT 16.030 144.780 16.210 144.820 ;
        RECT 16.030 144.110 16.285 144.780 ;
        RECT 16.465 143.800 16.750 144.600 ;
        RECT 16.930 144.520 17.180 145.110 ;
        RECT 17.380 145.755 17.700 146.085 ;
        RECT 17.880 145.870 18.540 146.350 ;
        RECT 18.740 145.960 19.590 146.130 ;
        RECT 17.380 144.860 17.570 145.755 ;
        RECT 17.890 145.430 18.550 145.700 ;
        RECT 18.220 145.370 18.550 145.430 ;
        RECT 17.740 145.200 18.070 145.260 ;
        RECT 18.740 145.200 18.910 145.960 ;
        RECT 20.150 145.890 20.470 146.350 ;
        RECT 20.670 145.710 20.920 146.140 ;
        RECT 21.210 145.910 21.620 146.350 ;
        RECT 21.790 145.970 22.805 146.170 ;
        RECT 19.080 145.540 20.330 145.710 ;
        RECT 19.080 145.420 19.410 145.540 ;
        RECT 17.740 145.030 19.640 145.200 ;
        RECT 17.380 144.690 19.300 144.860 ;
        RECT 17.380 144.670 17.700 144.690 ;
        RECT 16.930 144.010 17.260 144.520 ;
        RECT 17.530 144.060 17.700 144.670 ;
        RECT 19.470 144.520 19.640 145.030 ;
        RECT 19.810 144.960 19.990 145.370 ;
        RECT 20.160 144.780 20.330 145.540 ;
        RECT 17.870 143.800 18.200 144.490 ;
        RECT 18.430 144.350 19.640 144.520 ;
        RECT 19.810 144.470 20.330 144.780 ;
        RECT 20.500 145.370 20.920 145.710 ;
        RECT 21.210 145.370 21.620 145.700 ;
        RECT 20.500 144.600 20.690 145.370 ;
        RECT 21.790 145.240 21.960 145.970 ;
        RECT 23.105 145.800 23.275 146.130 ;
        RECT 23.445 145.970 23.775 146.350 ;
        RECT 22.130 145.420 22.480 145.790 ;
        RECT 21.790 145.200 22.210 145.240 ;
        RECT 20.860 145.030 22.210 145.200 ;
        RECT 20.860 144.870 21.110 145.030 ;
        RECT 21.620 144.600 21.870 144.860 ;
        RECT 20.500 144.350 21.870 144.600 ;
        RECT 18.430 144.060 18.670 144.350 ;
        RECT 19.470 144.270 19.640 144.350 ;
        RECT 18.870 143.800 19.290 144.180 ;
        RECT 19.470 144.020 20.100 144.270 ;
        RECT 20.570 143.800 20.900 144.180 ;
        RECT 21.070 144.060 21.240 144.350 ;
        RECT 22.040 144.185 22.210 145.030 ;
        RECT 22.660 144.860 22.880 145.730 ;
        RECT 23.105 145.610 23.800 145.800 ;
        RECT 22.380 144.480 22.880 144.860 ;
        RECT 23.050 144.810 23.460 145.430 ;
        RECT 23.630 144.640 23.800 145.610 ;
        RECT 23.105 144.470 23.800 144.640 ;
        RECT 21.420 143.800 21.800 144.180 ;
        RECT 22.040 144.015 22.870 144.185 ;
        RECT 23.105 143.970 23.275 144.470 ;
        RECT 23.445 143.800 23.775 144.300 ;
        RECT 23.990 143.970 24.215 146.090 ;
        RECT 24.385 145.970 24.715 146.350 ;
        RECT 24.885 145.800 25.055 146.090 ;
        RECT 24.390 145.630 25.055 145.800 ;
        RECT 24.390 144.640 24.620 145.630 ;
        RECT 25.315 145.625 25.605 146.350 ;
        RECT 25.775 145.675 26.035 146.180 ;
        RECT 26.215 145.970 26.545 146.350 ;
        RECT 26.725 145.800 26.895 146.180 ;
        RECT 24.790 144.810 25.140 145.460 ;
        RECT 24.390 144.470 25.055 144.640 ;
        RECT 24.385 143.800 24.715 144.300 ;
        RECT 24.885 143.970 25.055 144.470 ;
        RECT 25.315 143.800 25.605 144.965 ;
        RECT 25.775 144.875 25.945 145.675 ;
        RECT 26.230 145.630 26.895 145.800 ;
        RECT 26.230 145.375 26.400 145.630 ;
        RECT 27.155 145.580 29.745 146.350 ;
        RECT 26.115 145.045 26.400 145.375 ;
        RECT 26.635 145.080 26.965 145.450 ;
        RECT 26.230 144.900 26.400 145.045 ;
        RECT 25.775 143.970 26.045 144.875 ;
        RECT 26.230 144.730 26.895 144.900 ;
        RECT 26.215 143.800 26.545 144.560 ;
        RECT 26.725 143.970 26.895 144.730 ;
        RECT 27.155 144.890 28.365 145.410 ;
        RECT 28.535 145.060 29.745 145.580 ;
        RECT 29.915 145.550 30.255 146.180 ;
        RECT 30.425 145.550 30.675 146.350 ;
        RECT 30.865 145.700 31.195 146.180 ;
        RECT 31.365 145.890 31.590 146.350 ;
        RECT 31.760 145.700 32.090 146.180 ;
        RECT 29.915 144.940 30.090 145.550 ;
        RECT 30.865 145.530 32.090 145.700 ;
        RECT 32.720 145.570 33.220 146.180 ;
        RECT 34.145 145.800 34.315 146.090 ;
        RECT 34.485 145.970 34.815 146.350 ;
        RECT 34.145 145.630 34.810 145.800 ;
        RECT 30.260 145.190 30.955 145.360 ;
        RECT 31.130 145.330 31.550 145.360 ;
        RECT 30.785 144.940 30.955 145.190 ;
        RECT 31.125 145.160 31.550 145.330 ;
        RECT 31.720 145.160 32.050 145.360 ;
        RECT 32.220 145.160 32.550 145.360 ;
        RECT 32.720 144.940 32.890 145.570 ;
        RECT 33.075 145.110 33.425 145.360 ;
        RECT 27.155 143.800 29.745 144.890 ;
        RECT 29.915 143.970 30.255 144.940 ;
        RECT 30.425 143.800 30.595 144.940 ;
        RECT 30.785 144.770 33.220 144.940 ;
        RECT 34.060 144.810 34.410 145.460 ;
        RECT 30.865 143.800 31.115 144.600 ;
        RECT 31.760 143.970 32.090 144.770 ;
        RECT 32.390 143.800 32.720 144.600 ;
        RECT 32.890 143.970 33.220 144.770 ;
        RECT 34.580 144.640 34.810 145.630 ;
        RECT 34.145 144.470 34.810 144.640 ;
        RECT 34.145 143.970 34.315 144.470 ;
        RECT 34.485 143.800 34.815 144.300 ;
        RECT 34.985 143.970 35.210 146.090 ;
        RECT 35.425 145.970 35.755 146.350 ;
        RECT 35.925 145.800 36.095 146.130 ;
        RECT 36.395 145.970 37.410 146.170 ;
        RECT 35.400 145.610 36.095 145.800 ;
        RECT 35.400 144.640 35.570 145.610 ;
        RECT 35.740 144.810 36.150 145.430 ;
        RECT 36.320 144.860 36.540 145.730 ;
        RECT 36.720 145.420 37.070 145.790 ;
        RECT 37.240 145.240 37.410 145.970 ;
        RECT 37.580 145.910 37.990 146.350 ;
        RECT 38.280 145.710 38.530 146.140 ;
        RECT 38.730 145.890 39.050 146.350 ;
        RECT 39.610 145.960 40.460 146.130 ;
        RECT 37.580 145.370 37.990 145.700 ;
        RECT 38.280 145.370 38.700 145.710 ;
        RECT 36.990 145.200 37.410 145.240 ;
        RECT 36.990 145.030 38.340 145.200 ;
        RECT 35.400 144.470 36.095 144.640 ;
        RECT 36.320 144.480 36.820 144.860 ;
        RECT 35.425 143.800 35.755 144.300 ;
        RECT 35.925 143.970 36.095 144.470 ;
        RECT 36.990 144.185 37.160 145.030 ;
        RECT 38.090 144.870 38.340 145.030 ;
        RECT 37.330 144.600 37.580 144.860 ;
        RECT 38.510 144.600 38.700 145.370 ;
        RECT 37.330 144.350 38.700 144.600 ;
        RECT 38.870 145.540 40.120 145.710 ;
        RECT 38.870 144.780 39.040 145.540 ;
        RECT 39.790 145.420 40.120 145.540 ;
        RECT 39.210 144.960 39.390 145.370 ;
        RECT 40.290 145.200 40.460 145.960 ;
        RECT 40.660 145.870 41.320 146.350 ;
        RECT 41.500 145.755 41.820 146.085 ;
        RECT 40.650 145.430 41.310 145.700 ;
        RECT 40.650 145.370 40.980 145.430 ;
        RECT 41.130 145.200 41.460 145.260 ;
        RECT 39.560 145.030 41.460 145.200 ;
        RECT 38.870 144.470 39.390 144.780 ;
        RECT 39.560 144.520 39.730 145.030 ;
        RECT 41.630 144.860 41.820 145.755 ;
        RECT 39.900 144.690 41.820 144.860 ;
        RECT 41.500 144.670 41.820 144.690 ;
        RECT 42.020 145.440 42.270 146.090 ;
        RECT 42.450 145.890 42.735 146.350 ;
        RECT 42.915 145.640 43.170 146.170 ;
        RECT 42.020 145.110 42.820 145.440 ;
        RECT 39.560 144.350 40.770 144.520 ;
        RECT 36.330 144.015 37.160 144.185 ;
        RECT 37.400 143.800 37.780 144.180 ;
        RECT 37.960 144.060 38.130 144.350 ;
        RECT 39.560 144.270 39.730 144.350 ;
        RECT 38.300 143.800 38.630 144.180 ;
        RECT 39.100 144.020 39.730 144.270 ;
        RECT 39.910 143.800 40.330 144.180 ;
        RECT 40.530 144.060 40.770 144.350 ;
        RECT 41.000 143.800 41.330 144.490 ;
        RECT 41.500 144.060 41.670 144.670 ;
        RECT 42.020 144.520 42.270 145.110 ;
        RECT 42.990 144.990 43.170 145.640 ;
        RECT 44.180 145.610 44.435 146.180 ;
        RECT 44.605 145.950 44.935 146.350 ;
        RECT 45.360 145.815 45.890 146.180 ;
        RECT 46.080 146.010 46.355 146.180 ;
        RECT 46.075 145.840 46.355 146.010 ;
        RECT 45.360 145.780 45.535 145.815 ;
        RECT 44.605 145.610 45.535 145.780 ;
        RECT 42.990 144.820 43.255 144.990 ;
        RECT 44.180 144.940 44.350 145.610 ;
        RECT 44.605 145.440 44.775 145.610 ;
        RECT 44.520 145.110 44.775 145.440 ;
        RECT 45.000 145.110 45.195 145.440 ;
        RECT 42.990 144.780 43.170 144.820 ;
        RECT 41.940 144.010 42.270 144.520 ;
        RECT 42.450 143.800 42.735 144.600 ;
        RECT 42.915 144.110 43.170 144.780 ;
        RECT 44.180 143.970 44.515 144.940 ;
        RECT 44.685 143.800 44.855 144.940 ;
        RECT 45.025 144.140 45.195 145.110 ;
        RECT 45.365 144.480 45.535 145.610 ;
        RECT 45.705 144.820 45.875 145.620 ;
        RECT 46.080 145.020 46.355 145.840 ;
        RECT 46.525 144.820 46.715 146.180 ;
        RECT 46.895 145.815 47.405 146.350 ;
        RECT 47.625 145.540 47.870 146.145 ;
        RECT 48.315 145.580 50.905 146.350 ;
        RECT 51.075 145.625 51.365 146.350 ;
        RECT 51.535 145.580 53.205 146.350 ;
        RECT 46.915 145.370 48.145 145.540 ;
        RECT 45.705 144.650 46.715 144.820 ;
        RECT 46.885 144.805 47.635 144.995 ;
        RECT 45.365 144.310 46.490 144.480 ;
        RECT 46.885 144.140 47.055 144.805 ;
        RECT 47.805 144.560 48.145 145.370 ;
        RECT 45.025 143.970 47.055 144.140 ;
        RECT 47.225 143.800 47.395 144.560 ;
        RECT 47.630 144.150 48.145 144.560 ;
        RECT 48.315 144.890 49.525 145.410 ;
        RECT 49.695 145.060 50.905 145.580 ;
        RECT 48.315 143.800 50.905 144.890 ;
        RECT 51.075 143.800 51.365 144.965 ;
        RECT 51.535 144.890 52.285 145.410 ;
        RECT 52.455 145.060 53.205 145.580 ;
        RECT 53.415 145.530 53.645 146.350 ;
        RECT 53.815 145.550 54.145 146.180 ;
        RECT 53.395 145.110 53.725 145.360 ;
        RECT 53.895 144.950 54.145 145.550 ;
        RECT 54.315 145.530 54.525 146.350 ;
        RECT 55.030 145.540 55.275 146.145 ;
        RECT 55.495 145.815 56.005 146.350 ;
        RECT 51.535 143.800 53.205 144.890 ;
        RECT 53.415 143.800 53.645 144.940 ;
        RECT 53.815 143.970 54.145 144.950 ;
        RECT 54.755 145.370 55.985 145.540 ;
        RECT 54.315 143.800 54.525 144.940 ;
        RECT 54.755 144.560 55.095 145.370 ;
        RECT 55.265 144.805 56.015 144.995 ;
        RECT 54.755 144.150 55.270 144.560 ;
        RECT 55.505 143.800 55.675 144.560 ;
        RECT 55.845 144.140 56.015 144.805 ;
        RECT 56.185 144.820 56.375 146.180 ;
        RECT 56.545 145.330 56.820 146.180 ;
        RECT 57.010 145.815 57.540 146.180 ;
        RECT 57.965 145.950 58.295 146.350 ;
        RECT 57.365 145.780 57.540 145.815 ;
        RECT 56.545 145.160 56.825 145.330 ;
        RECT 56.545 145.020 56.820 145.160 ;
        RECT 57.025 144.820 57.195 145.620 ;
        RECT 56.185 144.650 57.195 144.820 ;
        RECT 57.365 145.610 58.295 145.780 ;
        RECT 58.465 145.610 58.720 146.180 ;
        RECT 57.365 144.480 57.535 145.610 ;
        RECT 58.125 145.440 58.295 145.610 ;
        RECT 56.410 144.310 57.535 144.480 ;
        RECT 57.705 145.110 57.900 145.440 ;
        RECT 58.125 145.110 58.380 145.440 ;
        RECT 57.705 144.140 57.875 145.110 ;
        RECT 58.550 144.940 58.720 145.610 ;
        RECT 58.895 145.600 60.105 146.350 ;
        RECT 60.280 145.805 65.625 146.350 ;
        RECT 55.845 143.970 57.875 144.140 ;
        RECT 58.045 143.800 58.215 144.940 ;
        RECT 58.385 143.970 58.720 144.940 ;
        RECT 58.895 144.890 59.415 145.430 ;
        RECT 59.585 145.060 60.105 145.600 ;
        RECT 58.895 143.800 60.105 144.890 ;
        RECT 61.870 144.235 62.220 145.485 ;
        RECT 63.700 144.975 64.040 145.805 ;
        RECT 65.885 145.800 66.055 146.180 ;
        RECT 66.270 145.970 66.600 146.350 ;
        RECT 65.885 145.630 66.600 145.800 ;
        RECT 65.795 145.080 66.150 145.450 ;
        RECT 66.430 145.440 66.600 145.630 ;
        RECT 66.770 145.605 67.025 146.180 ;
        RECT 66.430 145.110 66.685 145.440 ;
        RECT 66.430 144.900 66.600 145.110 ;
        RECT 65.885 144.730 66.600 144.900 ;
        RECT 66.855 144.875 67.025 145.605 ;
        RECT 67.200 145.510 67.460 146.350 ;
        RECT 67.635 145.600 68.845 146.350 ;
        RECT 60.280 143.800 65.625 144.235 ;
        RECT 65.885 143.970 66.055 144.730 ;
        RECT 66.270 143.800 66.600 144.560 ;
        RECT 66.770 143.970 67.025 144.875 ;
        RECT 67.200 143.800 67.460 144.950 ;
        RECT 67.635 144.890 68.155 145.430 ;
        RECT 68.325 145.060 68.845 145.600 ;
        RECT 69.015 145.580 72.525 146.350 ;
        RECT 69.015 144.890 70.705 145.410 ;
        RECT 70.875 145.060 72.525 145.580 ;
        RECT 72.970 145.540 73.215 146.145 ;
        RECT 73.435 145.815 73.945 146.350 ;
        RECT 72.695 145.370 73.925 145.540 ;
        RECT 67.635 143.800 68.845 144.890 ;
        RECT 69.015 143.800 72.525 144.890 ;
        RECT 72.695 144.560 73.035 145.370 ;
        RECT 73.205 144.805 73.955 144.995 ;
        RECT 72.695 144.150 73.210 144.560 ;
        RECT 73.445 143.800 73.615 144.560 ;
        RECT 73.785 144.140 73.955 144.805 ;
        RECT 74.125 144.820 74.315 146.180 ;
        RECT 74.485 145.330 74.760 146.180 ;
        RECT 74.950 145.815 75.480 146.180 ;
        RECT 75.905 145.950 76.235 146.350 ;
        RECT 75.305 145.780 75.480 145.815 ;
        RECT 74.485 145.160 74.765 145.330 ;
        RECT 74.485 145.020 74.760 145.160 ;
        RECT 74.965 144.820 75.135 145.620 ;
        RECT 74.125 144.650 75.135 144.820 ;
        RECT 75.305 145.610 76.235 145.780 ;
        RECT 76.405 145.610 76.660 146.180 ;
        RECT 76.835 145.625 77.125 146.350 ;
        RECT 75.305 144.480 75.475 145.610 ;
        RECT 76.065 145.440 76.235 145.610 ;
        RECT 74.350 144.310 75.475 144.480 ;
        RECT 75.645 145.110 75.840 145.440 ;
        RECT 76.065 145.110 76.320 145.440 ;
        RECT 75.645 144.140 75.815 145.110 ;
        RECT 76.490 144.940 76.660 145.610 ;
        RECT 78.030 145.540 78.275 146.145 ;
        RECT 78.495 145.815 79.005 146.350 ;
        RECT 77.755 145.370 78.985 145.540 ;
        RECT 73.785 143.970 75.815 144.140 ;
        RECT 75.985 143.800 76.155 144.940 ;
        RECT 76.325 143.970 76.660 144.940 ;
        RECT 76.835 143.800 77.125 144.965 ;
        RECT 77.755 144.560 78.095 145.370 ;
        RECT 78.265 144.805 79.015 144.995 ;
        RECT 77.755 144.150 78.270 144.560 ;
        RECT 78.505 143.800 78.675 144.560 ;
        RECT 78.845 144.140 79.015 144.805 ;
        RECT 79.185 144.820 79.375 146.180 ;
        RECT 79.545 146.010 79.820 146.180 ;
        RECT 79.545 145.840 79.825 146.010 ;
        RECT 79.545 145.020 79.820 145.840 ;
        RECT 80.010 145.815 80.540 146.180 ;
        RECT 80.965 145.950 81.295 146.350 ;
        RECT 80.365 145.780 80.540 145.815 ;
        RECT 80.025 144.820 80.195 145.620 ;
        RECT 79.185 144.650 80.195 144.820 ;
        RECT 80.365 145.610 81.295 145.780 ;
        RECT 81.465 145.610 81.720 146.180 ;
        RECT 80.365 144.480 80.535 145.610 ;
        RECT 81.125 145.440 81.295 145.610 ;
        RECT 79.410 144.310 80.535 144.480 ;
        RECT 80.705 145.110 80.900 145.440 ;
        RECT 81.125 145.110 81.380 145.440 ;
        RECT 80.705 144.140 80.875 145.110 ;
        RECT 81.550 144.940 81.720 145.610 ;
        RECT 81.955 145.530 82.165 146.350 ;
        RECT 82.335 145.550 82.665 146.180 ;
        RECT 82.335 144.950 82.585 145.550 ;
        RECT 82.835 145.530 83.065 146.350 ;
        RECT 83.850 145.720 84.135 146.180 ;
        RECT 84.305 145.890 84.575 146.350 ;
        RECT 83.850 145.550 84.805 145.720 ;
        RECT 82.755 145.110 83.085 145.360 ;
        RECT 78.845 143.970 80.875 144.140 ;
        RECT 81.045 143.800 81.215 144.940 ;
        RECT 81.385 143.970 81.720 144.940 ;
        RECT 81.955 143.800 82.165 144.940 ;
        RECT 82.335 143.970 82.665 144.950 ;
        RECT 82.835 143.800 83.065 144.940 ;
        RECT 83.735 144.820 84.425 145.380 ;
        RECT 84.595 144.650 84.805 145.550 ;
        RECT 83.850 144.430 84.805 144.650 ;
        RECT 84.975 145.380 85.375 146.180 ;
        RECT 85.565 145.720 85.845 146.180 ;
        RECT 86.365 145.890 86.690 146.350 ;
        RECT 85.565 145.550 86.690 145.720 ;
        RECT 86.860 145.610 87.245 146.180 ;
        RECT 86.240 145.440 86.690 145.550 ;
        RECT 84.975 144.820 86.070 145.380 ;
        RECT 86.240 145.110 86.795 145.440 ;
        RECT 83.850 143.970 84.135 144.430 ;
        RECT 84.305 143.800 84.575 144.260 ;
        RECT 84.975 143.970 85.375 144.820 ;
        RECT 86.240 144.650 86.690 145.110 ;
        RECT 86.965 144.940 87.245 145.610 ;
        RECT 87.875 145.580 90.465 146.350 ;
        RECT 90.640 145.805 95.985 146.350 ;
        RECT 85.565 144.430 86.690 144.650 ;
        RECT 85.565 143.970 85.845 144.430 ;
        RECT 86.365 143.800 86.690 144.260 ;
        RECT 86.860 143.970 87.245 144.940 ;
        RECT 87.875 144.890 89.085 145.410 ;
        RECT 89.255 145.060 90.465 145.580 ;
        RECT 87.875 143.800 90.465 144.890 ;
        RECT 92.230 144.235 92.580 145.485 ;
        RECT 94.060 144.975 94.400 145.805 ;
        RECT 96.155 145.675 96.425 146.020 ;
        RECT 96.615 145.950 96.995 146.350 ;
        RECT 97.165 145.780 97.335 146.130 ;
        RECT 97.505 145.950 97.835 146.350 ;
        RECT 98.035 145.780 98.205 146.130 ;
        RECT 98.405 145.850 98.735 146.350 ;
        RECT 96.155 144.940 96.325 145.675 ;
        RECT 96.595 145.610 98.205 145.780 ;
        RECT 96.595 145.440 96.765 145.610 ;
        RECT 96.495 145.110 96.765 145.440 ;
        RECT 96.935 145.110 97.340 145.440 ;
        RECT 96.595 144.940 96.765 145.110 ;
        RECT 97.510 144.990 98.220 145.440 ;
        RECT 98.390 145.110 98.740 145.680 ;
        RECT 98.915 145.550 99.255 146.180 ;
        RECT 99.425 145.550 99.675 146.350 ;
        RECT 99.865 145.700 100.195 146.180 ;
        RECT 100.365 145.890 100.590 146.350 ;
        RECT 100.760 145.700 101.090 146.180 ;
        RECT 98.915 145.500 99.145 145.550 ;
        RECT 99.865 145.530 101.090 145.700 ;
        RECT 101.720 145.570 102.220 146.180 ;
        RECT 102.595 145.625 102.885 146.350 ;
        RECT 103.055 145.600 104.265 146.350 ;
        RECT 90.640 143.800 95.985 144.235 ;
        RECT 96.155 143.970 96.425 144.940 ;
        RECT 96.595 144.770 97.320 144.940 ;
        RECT 97.510 144.820 98.225 144.990 ;
        RECT 98.915 144.940 99.090 145.500 ;
        RECT 99.260 145.190 99.955 145.360 ;
        RECT 99.785 144.940 99.955 145.190 ;
        RECT 100.130 145.160 100.550 145.360 ;
        RECT 100.720 145.160 101.050 145.360 ;
        RECT 101.220 145.160 101.550 145.360 ;
        RECT 101.720 144.940 101.890 145.570 ;
        RECT 102.075 145.110 102.425 145.360 ;
        RECT 97.150 144.650 97.320 144.770 ;
        RECT 98.420 144.650 98.740 144.940 ;
        RECT 96.635 143.800 96.915 144.600 ;
        RECT 97.150 144.480 98.740 144.650 ;
        RECT 97.085 144.020 98.740 144.310 ;
        RECT 98.915 143.970 99.255 144.940 ;
        RECT 99.425 143.800 99.595 144.940 ;
        RECT 99.785 144.770 102.220 144.940 ;
        RECT 99.865 143.800 100.115 144.600 ;
        RECT 100.760 143.970 101.090 144.770 ;
        RECT 101.390 143.800 101.720 144.600 ;
        RECT 101.890 143.970 102.220 144.770 ;
        RECT 102.595 143.800 102.885 144.965 ;
        RECT 103.055 144.890 103.575 145.430 ;
        RECT 103.745 145.060 104.265 145.600 ;
        RECT 104.435 145.580 107.945 146.350 ;
        RECT 104.435 144.890 106.125 145.410 ;
        RECT 106.295 145.060 107.945 145.580 ;
        RECT 108.155 145.530 108.385 146.350 ;
        RECT 108.555 145.550 108.885 146.180 ;
        RECT 108.135 145.110 108.465 145.360 ;
        RECT 108.635 144.950 108.885 145.550 ;
        RECT 109.055 145.530 109.265 146.350 ;
        RECT 110.045 145.800 110.215 146.180 ;
        RECT 110.395 145.970 110.725 146.350 ;
        RECT 110.045 145.630 110.710 145.800 ;
        RECT 110.905 145.675 111.165 146.180 ;
        RECT 109.975 145.080 110.305 145.450 ;
        RECT 110.540 145.375 110.710 145.630 ;
        RECT 103.055 143.800 104.265 144.890 ;
        RECT 104.435 143.800 107.945 144.890 ;
        RECT 108.155 143.800 108.385 144.940 ;
        RECT 108.555 143.970 108.885 144.950 ;
        RECT 110.540 145.045 110.825 145.375 ;
        RECT 109.055 143.800 109.265 144.940 ;
        RECT 110.540 144.900 110.710 145.045 ;
        RECT 110.045 144.730 110.710 144.900 ;
        RECT 110.995 144.875 111.165 145.675 ;
        RECT 111.795 145.580 114.385 146.350 ;
        RECT 114.555 145.600 115.765 146.350 ;
        RECT 110.045 143.970 110.215 144.730 ;
        RECT 110.395 143.800 110.725 144.560 ;
        RECT 110.895 143.970 111.165 144.875 ;
        RECT 111.795 144.890 113.005 145.410 ;
        RECT 113.175 145.060 114.385 145.580 ;
        RECT 114.555 144.890 115.075 145.430 ;
        RECT 115.245 145.060 115.765 145.600 ;
        RECT 111.795 143.800 114.385 144.890 ;
        RECT 114.555 143.800 115.765 144.890 ;
        RECT 10.510 143.630 115.850 143.800 ;
        RECT 10.595 142.540 11.805 143.630 ;
        RECT 10.595 141.830 11.115 142.370 ;
        RECT 11.285 142.000 11.805 142.540 ;
        RECT 12.435 142.465 12.725 143.630 ;
        RECT 13.820 143.195 19.165 143.630 ;
        RECT 15.410 141.945 15.760 143.195 ;
        RECT 19.425 142.700 19.595 143.460 ;
        RECT 19.775 142.870 20.105 143.630 ;
        RECT 19.425 142.530 20.090 142.700 ;
        RECT 20.275 142.555 20.545 143.460 ;
        RECT 10.595 141.080 11.805 141.830 ;
        RECT 12.435 141.080 12.725 141.805 ;
        RECT 17.240 141.625 17.580 142.455 ;
        RECT 19.920 142.385 20.090 142.530 ;
        RECT 19.355 141.980 19.685 142.350 ;
        RECT 19.920 142.055 20.205 142.385 ;
        RECT 19.920 141.800 20.090 142.055 ;
        RECT 19.425 141.630 20.090 141.800 ;
        RECT 20.375 141.755 20.545 142.555 ;
        RECT 20.775 142.490 20.985 143.630 ;
        RECT 21.155 142.480 21.485 143.460 ;
        RECT 21.655 142.490 21.885 143.630 ;
        RECT 22.095 142.540 23.305 143.630 ;
        RECT 23.475 142.540 26.985 143.630 ;
        RECT 27.160 143.195 32.505 143.630 ;
        RECT 32.680 143.195 38.025 143.630 ;
        RECT 13.820 141.080 19.165 141.625 ;
        RECT 19.425 141.250 19.595 141.630 ;
        RECT 19.775 141.080 20.105 141.460 ;
        RECT 20.285 141.250 20.545 141.755 ;
        RECT 20.775 141.080 20.985 141.900 ;
        RECT 21.155 141.880 21.405 142.480 ;
        RECT 21.575 142.070 21.905 142.320 ;
        RECT 22.095 142.000 22.615 142.540 ;
        RECT 21.155 141.250 21.485 141.880 ;
        RECT 21.655 141.080 21.885 141.900 ;
        RECT 22.785 141.830 23.305 142.370 ;
        RECT 23.475 142.020 25.165 142.540 ;
        RECT 25.335 141.850 26.985 142.370 ;
        RECT 28.750 141.945 29.100 143.195 ;
        RECT 22.095 141.080 23.305 141.830 ;
        RECT 23.475 141.080 26.985 141.850 ;
        RECT 30.580 141.625 30.920 142.455 ;
        RECT 34.270 141.945 34.620 143.195 ;
        RECT 38.195 142.465 38.485 143.630 ;
        RECT 39.115 142.540 41.705 143.630 ;
        RECT 41.875 142.555 42.145 143.460 ;
        RECT 42.315 142.870 42.645 143.630 ;
        RECT 42.825 142.700 42.995 143.460 ;
        RECT 36.100 141.625 36.440 142.455 ;
        RECT 39.115 142.020 40.325 142.540 ;
        RECT 40.495 141.850 41.705 142.370 ;
        RECT 27.160 141.080 32.505 141.625 ;
        RECT 32.680 141.080 38.025 141.625 ;
        RECT 38.195 141.080 38.485 141.805 ;
        RECT 39.115 141.080 41.705 141.850 ;
        RECT 41.875 141.755 42.045 142.555 ;
        RECT 42.330 142.530 42.995 142.700 ;
        RECT 42.330 142.385 42.500 142.530 ;
        RECT 42.215 142.055 42.500 142.385 ;
        RECT 43.255 142.490 43.595 143.460 ;
        RECT 43.765 142.490 43.935 143.630 ;
        RECT 44.205 142.830 44.455 143.630 ;
        RECT 45.100 142.660 45.430 143.460 ;
        RECT 45.730 142.830 46.060 143.630 ;
        RECT 46.230 142.660 46.560 143.460 ;
        RECT 44.125 142.490 46.560 142.660 ;
        RECT 46.935 142.540 48.145 143.630 ;
        RECT 42.330 141.800 42.500 142.055 ;
        RECT 42.735 141.980 43.065 142.350 ;
        RECT 43.255 141.880 43.430 142.490 ;
        RECT 44.125 142.240 44.295 142.490 ;
        RECT 43.600 142.070 44.295 142.240 ;
        RECT 44.470 142.070 44.890 142.270 ;
        RECT 45.060 142.070 45.390 142.270 ;
        RECT 45.560 142.070 45.890 142.270 ;
        RECT 41.875 141.250 42.135 141.755 ;
        RECT 42.330 141.630 42.995 141.800 ;
        RECT 42.315 141.080 42.645 141.460 ;
        RECT 42.825 141.250 42.995 141.630 ;
        RECT 43.255 141.250 43.595 141.880 ;
        RECT 43.765 141.080 44.015 141.880 ;
        RECT 44.205 141.730 45.430 141.900 ;
        RECT 44.205 141.250 44.535 141.730 ;
        RECT 44.705 141.080 44.930 141.540 ;
        RECT 45.100 141.250 45.430 141.730 ;
        RECT 46.060 141.860 46.230 142.490 ;
        RECT 46.415 142.070 46.765 142.320 ;
        RECT 46.935 142.000 47.455 142.540 ;
        RECT 48.315 142.490 48.655 143.460 ;
        RECT 48.825 142.490 48.995 143.630 ;
        RECT 49.265 142.830 49.515 143.630 ;
        RECT 50.160 142.660 50.490 143.460 ;
        RECT 50.790 142.830 51.120 143.630 ;
        RECT 51.290 142.660 51.620 143.460 ;
        RECT 49.185 142.490 51.620 142.660 ;
        RECT 51.995 142.540 53.205 143.630 ;
        RECT 46.060 141.250 46.560 141.860 ;
        RECT 47.625 141.830 48.145 142.370 ;
        RECT 46.935 141.080 48.145 141.830 ;
        RECT 48.315 141.880 48.490 142.490 ;
        RECT 49.185 142.240 49.355 142.490 ;
        RECT 48.660 142.070 49.355 142.240 ;
        RECT 49.530 142.070 49.950 142.270 ;
        RECT 50.120 142.070 50.450 142.270 ;
        RECT 50.620 142.070 50.950 142.270 ;
        RECT 48.315 141.250 48.655 141.880 ;
        RECT 48.825 141.080 49.075 141.880 ;
        RECT 49.265 141.730 50.490 141.900 ;
        RECT 49.265 141.250 49.595 141.730 ;
        RECT 49.765 141.080 49.990 141.540 ;
        RECT 50.160 141.250 50.490 141.730 ;
        RECT 51.120 141.860 51.290 142.490 ;
        RECT 51.475 142.070 51.825 142.320 ;
        RECT 51.995 142.000 52.515 142.540 ;
        RECT 53.415 142.490 53.645 143.630 ;
        RECT 53.815 142.480 54.145 143.460 ;
        RECT 54.315 142.490 54.525 143.630 ;
        RECT 51.120 141.250 51.620 141.860 ;
        RECT 52.685 141.830 53.205 142.370 ;
        RECT 53.395 142.070 53.725 142.320 ;
        RECT 51.995 141.080 53.205 141.830 ;
        RECT 53.415 141.080 53.645 141.900 ;
        RECT 53.895 141.880 54.145 142.480 ;
        RECT 54.760 142.440 55.015 143.320 ;
        RECT 55.185 142.490 55.490 143.630 ;
        RECT 55.830 143.250 56.160 143.630 ;
        RECT 56.340 143.080 56.510 143.370 ;
        RECT 56.680 143.170 56.930 143.630 ;
        RECT 55.710 142.910 56.510 143.080 ;
        RECT 57.100 143.120 57.970 143.460 ;
        RECT 53.815 141.250 54.145 141.880 ;
        RECT 54.315 141.080 54.525 141.900 ;
        RECT 54.760 141.790 54.970 142.440 ;
        RECT 55.710 142.320 55.880 142.910 ;
        RECT 57.100 142.740 57.270 143.120 ;
        RECT 58.205 143.000 58.375 143.460 ;
        RECT 58.545 143.170 58.915 143.630 ;
        RECT 59.210 143.030 59.380 143.370 ;
        RECT 59.550 143.200 59.880 143.630 ;
        RECT 60.115 143.030 60.285 143.370 ;
        RECT 56.050 142.570 57.270 142.740 ;
        RECT 57.440 142.660 57.900 142.950 ;
        RECT 58.205 142.830 58.765 143.000 ;
        RECT 59.210 142.860 60.285 143.030 ;
        RECT 60.455 143.130 61.135 143.460 ;
        RECT 61.350 143.130 61.600 143.460 ;
        RECT 61.770 143.170 62.020 143.630 ;
        RECT 58.595 142.690 58.765 142.830 ;
        RECT 57.440 142.650 58.405 142.660 ;
        RECT 57.100 142.480 57.270 142.570 ;
        RECT 57.730 142.490 58.405 142.650 ;
        RECT 55.140 142.290 55.880 142.320 ;
        RECT 55.140 141.990 56.055 142.290 ;
        RECT 55.730 141.815 56.055 141.990 ;
        RECT 54.760 141.260 55.015 141.790 ;
        RECT 55.185 141.080 55.490 141.540 ;
        RECT 55.735 141.460 56.055 141.815 ;
        RECT 56.225 142.030 56.765 142.400 ;
        RECT 57.100 142.310 57.505 142.480 ;
        RECT 56.225 141.630 56.465 142.030 ;
        RECT 56.945 141.860 57.165 142.140 ;
        RECT 56.635 141.690 57.165 141.860 ;
        RECT 56.635 141.460 56.805 141.690 ;
        RECT 57.335 141.530 57.505 142.310 ;
        RECT 57.675 141.700 58.025 142.320 ;
        RECT 58.195 141.700 58.405 142.490 ;
        RECT 58.595 142.520 60.095 142.690 ;
        RECT 58.595 141.830 58.765 142.520 ;
        RECT 60.455 142.350 60.625 143.130 ;
        RECT 61.430 143.000 61.600 143.130 ;
        RECT 58.935 142.180 60.625 142.350 ;
        RECT 60.795 142.570 61.260 142.960 ;
        RECT 61.430 142.830 61.825 143.000 ;
        RECT 58.935 142.000 59.105 142.180 ;
        RECT 55.735 141.290 56.805 141.460 ;
        RECT 56.975 141.080 57.165 141.520 ;
        RECT 57.335 141.250 58.285 141.530 ;
        RECT 58.595 141.440 58.855 141.830 ;
        RECT 59.275 141.760 60.065 142.010 ;
        RECT 58.505 141.270 58.855 141.440 ;
        RECT 59.065 141.080 59.395 141.540 ;
        RECT 60.270 141.470 60.440 142.180 ;
        RECT 60.795 141.980 60.965 142.570 ;
        RECT 60.610 141.760 60.965 141.980 ;
        RECT 61.135 141.760 61.485 142.380 ;
        RECT 61.655 141.470 61.825 142.830 ;
        RECT 62.190 142.660 62.515 143.445 ;
        RECT 61.995 141.610 62.455 142.660 ;
        RECT 60.270 141.300 61.125 141.470 ;
        RECT 61.330 141.300 61.825 141.470 ;
        RECT 61.995 141.080 62.325 141.440 ;
        RECT 62.685 141.340 62.855 143.460 ;
        RECT 63.025 143.130 63.355 143.630 ;
        RECT 63.525 142.960 63.780 143.460 ;
        RECT 63.030 142.790 63.780 142.960 ;
        RECT 63.030 141.800 63.260 142.790 ;
        RECT 63.430 141.970 63.780 142.620 ;
        RECT 63.955 142.465 64.245 143.630 ;
        RECT 64.415 142.540 67.005 143.630 ;
        RECT 64.415 142.020 65.625 142.540 ;
        RECT 67.175 142.490 67.445 143.460 ;
        RECT 67.655 142.830 67.935 143.630 ;
        RECT 68.105 143.120 69.760 143.410 ;
        RECT 68.170 142.780 69.760 142.950 ;
        RECT 68.170 142.660 68.340 142.780 ;
        RECT 67.615 142.490 68.340 142.660 ;
        RECT 65.795 141.850 67.005 142.370 ;
        RECT 63.030 141.630 63.780 141.800 ;
        RECT 63.025 141.080 63.355 141.460 ;
        RECT 63.525 141.340 63.780 141.630 ;
        RECT 63.955 141.080 64.245 141.805 ;
        RECT 64.415 141.080 67.005 141.850 ;
        RECT 67.175 141.755 67.345 142.490 ;
        RECT 67.615 142.320 67.785 142.490 ;
        RECT 68.530 142.440 69.245 142.610 ;
        RECT 69.440 142.490 69.760 142.780 ;
        RECT 69.935 142.490 70.275 143.460 ;
        RECT 70.445 142.490 70.615 143.630 ;
        RECT 70.885 142.830 71.135 143.630 ;
        RECT 71.780 142.660 72.110 143.460 ;
        RECT 72.410 142.830 72.740 143.630 ;
        RECT 72.910 142.660 73.240 143.460 ;
        RECT 70.805 142.490 73.240 142.660 ;
        RECT 73.990 142.650 74.245 143.320 ;
        RECT 74.425 142.830 74.710 143.630 ;
        RECT 74.890 142.910 75.220 143.420 ;
        RECT 67.515 141.990 67.785 142.320 ;
        RECT 67.955 141.990 68.360 142.320 ;
        RECT 68.530 141.990 69.240 142.440 ;
        RECT 67.615 141.820 67.785 141.990 ;
        RECT 67.175 141.410 67.445 141.755 ;
        RECT 67.615 141.650 69.225 141.820 ;
        RECT 69.410 141.750 69.760 142.320 ;
        RECT 69.935 141.930 70.110 142.490 ;
        RECT 70.805 142.240 70.975 142.490 ;
        RECT 70.280 142.070 70.975 142.240 ;
        RECT 71.150 142.070 71.570 142.270 ;
        RECT 71.740 142.070 72.070 142.270 ;
        RECT 72.240 142.070 72.570 142.270 ;
        RECT 69.935 141.880 70.165 141.930 ;
        RECT 67.635 141.080 68.015 141.480 ;
        RECT 68.185 141.300 68.355 141.650 ;
        RECT 68.525 141.080 68.855 141.480 ;
        RECT 69.055 141.300 69.225 141.650 ;
        RECT 69.425 141.080 69.755 141.580 ;
        RECT 69.935 141.250 70.275 141.880 ;
        RECT 70.445 141.080 70.695 141.880 ;
        RECT 70.885 141.730 72.110 141.900 ;
        RECT 70.885 141.250 71.215 141.730 ;
        RECT 71.385 141.080 71.610 141.540 ;
        RECT 71.780 141.250 72.110 141.730 ;
        RECT 72.740 141.860 72.910 142.490 ;
        RECT 73.095 142.070 73.445 142.320 ;
        RECT 73.990 141.930 74.170 142.650 ;
        RECT 74.890 142.320 75.140 142.910 ;
        RECT 75.490 142.760 75.660 143.370 ;
        RECT 75.830 142.940 76.160 143.630 ;
        RECT 76.390 143.080 76.630 143.370 ;
        RECT 76.830 143.250 77.250 143.630 ;
        RECT 77.430 143.160 78.060 143.410 ;
        RECT 78.530 143.250 78.860 143.630 ;
        RECT 77.430 143.080 77.600 143.160 ;
        RECT 79.030 143.080 79.200 143.370 ;
        RECT 79.380 143.250 79.760 143.630 ;
        RECT 80.000 143.245 80.830 143.415 ;
        RECT 76.390 142.910 77.600 143.080 ;
        RECT 74.340 141.990 75.140 142.320 ;
        RECT 72.740 141.250 73.240 141.860 ;
        RECT 73.905 141.790 74.170 141.930 ;
        RECT 73.905 141.760 74.245 141.790 ;
        RECT 73.990 141.260 74.245 141.760 ;
        RECT 74.425 141.080 74.710 141.540 ;
        RECT 74.890 141.340 75.140 141.990 ;
        RECT 75.340 142.740 75.660 142.760 ;
        RECT 75.340 142.570 77.260 142.740 ;
        RECT 75.340 141.675 75.530 142.570 ;
        RECT 77.430 142.400 77.600 142.910 ;
        RECT 77.770 142.650 78.290 142.960 ;
        RECT 75.700 142.230 77.600 142.400 ;
        RECT 75.700 142.170 76.030 142.230 ;
        RECT 76.180 142.000 76.510 142.060 ;
        RECT 75.850 141.730 76.510 142.000 ;
        RECT 75.340 141.345 75.660 141.675 ;
        RECT 75.840 141.080 76.500 141.560 ;
        RECT 76.700 141.470 76.870 142.230 ;
        RECT 77.770 142.060 77.950 142.470 ;
        RECT 77.040 141.890 77.370 142.010 ;
        RECT 78.120 141.890 78.290 142.650 ;
        RECT 77.040 141.720 78.290 141.890 ;
        RECT 78.460 142.830 79.830 143.080 ;
        RECT 78.460 142.060 78.650 142.830 ;
        RECT 79.580 142.570 79.830 142.830 ;
        RECT 78.820 142.400 79.070 142.560 ;
        RECT 80.000 142.400 80.170 143.245 ;
        RECT 81.065 142.960 81.235 143.460 ;
        RECT 81.405 143.130 81.735 143.630 ;
        RECT 80.340 142.570 80.840 142.950 ;
        RECT 81.065 142.790 81.760 142.960 ;
        RECT 78.820 142.230 80.170 142.400 ;
        RECT 79.750 142.190 80.170 142.230 ;
        RECT 78.460 141.720 78.880 142.060 ;
        RECT 79.170 141.730 79.580 142.060 ;
        RECT 76.700 141.300 77.550 141.470 ;
        RECT 78.110 141.080 78.430 141.540 ;
        RECT 78.630 141.290 78.880 141.720 ;
        RECT 79.170 141.080 79.580 141.520 ;
        RECT 79.750 141.460 79.920 142.190 ;
        RECT 80.090 141.640 80.440 142.010 ;
        RECT 80.620 141.700 80.840 142.570 ;
        RECT 81.010 142.000 81.420 142.620 ;
        RECT 81.590 141.820 81.760 142.790 ;
        RECT 81.065 141.630 81.760 141.820 ;
        RECT 79.750 141.260 80.765 141.460 ;
        RECT 81.065 141.300 81.235 141.630 ;
        RECT 81.405 141.080 81.735 141.460 ;
        RECT 81.950 141.340 82.175 143.460 ;
        RECT 82.345 143.130 82.675 143.630 ;
        RECT 82.845 142.960 83.015 143.460 ;
        RECT 84.200 143.195 89.545 143.630 ;
        RECT 82.350 142.790 83.015 142.960 ;
        RECT 82.350 141.800 82.580 142.790 ;
        RECT 82.750 141.970 83.100 142.620 ;
        RECT 85.790 141.945 86.140 143.195 ;
        RECT 89.715 142.465 90.005 143.630 ;
        RECT 90.175 142.540 93.685 143.630 ;
        RECT 93.860 143.195 99.205 143.630 ;
        RECT 99.380 143.195 104.725 143.630 ;
        RECT 82.350 141.630 83.015 141.800 ;
        RECT 82.345 141.080 82.675 141.460 ;
        RECT 82.845 141.340 83.015 141.630 ;
        RECT 87.620 141.625 87.960 142.455 ;
        RECT 90.175 142.020 91.865 142.540 ;
        RECT 92.035 141.850 93.685 142.370 ;
        RECT 95.450 141.945 95.800 143.195 ;
        RECT 84.200 141.080 89.545 141.625 ;
        RECT 89.715 141.080 90.005 141.805 ;
        RECT 90.175 141.080 93.685 141.850 ;
        RECT 97.280 141.625 97.620 142.455 ;
        RECT 100.970 141.945 101.320 143.195 ;
        RECT 104.895 142.870 105.410 143.280 ;
        RECT 105.645 142.870 105.815 143.630 ;
        RECT 105.985 143.290 108.015 143.460 ;
        RECT 102.800 141.625 103.140 142.455 ;
        RECT 104.895 142.060 105.235 142.870 ;
        RECT 105.985 142.625 106.155 143.290 ;
        RECT 106.550 142.950 107.675 143.120 ;
        RECT 105.405 142.435 106.155 142.625 ;
        RECT 106.325 142.610 107.335 142.780 ;
        RECT 104.895 141.890 106.125 142.060 ;
        RECT 93.860 141.080 99.205 141.625 ;
        RECT 99.380 141.080 104.725 141.625 ;
        RECT 105.170 141.285 105.415 141.890 ;
        RECT 105.635 141.080 106.145 141.615 ;
        RECT 106.325 141.250 106.515 142.610 ;
        RECT 106.685 142.270 106.960 142.410 ;
        RECT 106.685 142.100 106.965 142.270 ;
        RECT 106.685 141.250 106.960 142.100 ;
        RECT 107.165 141.810 107.335 142.610 ;
        RECT 107.505 141.820 107.675 142.950 ;
        RECT 107.845 142.320 108.015 143.290 ;
        RECT 108.185 142.490 108.355 143.630 ;
        RECT 108.525 142.490 108.860 143.460 ;
        RECT 109.075 142.490 109.305 143.630 ;
        RECT 107.845 141.990 108.040 142.320 ;
        RECT 108.265 141.990 108.520 142.320 ;
        RECT 108.265 141.820 108.435 141.990 ;
        RECT 108.690 141.820 108.860 142.490 ;
        RECT 109.475 142.480 109.805 143.460 ;
        RECT 109.975 142.490 110.185 143.630 ;
        RECT 110.875 142.540 114.385 143.630 ;
        RECT 114.555 142.540 115.765 143.630 ;
        RECT 109.055 142.070 109.385 142.320 ;
        RECT 107.505 141.650 108.435 141.820 ;
        RECT 107.505 141.615 107.680 141.650 ;
        RECT 107.150 141.250 107.680 141.615 ;
        RECT 108.105 141.080 108.435 141.480 ;
        RECT 108.605 141.250 108.860 141.820 ;
        RECT 109.075 141.080 109.305 141.900 ;
        RECT 109.555 141.880 109.805 142.480 ;
        RECT 110.875 142.020 112.565 142.540 ;
        RECT 109.475 141.250 109.805 141.880 ;
        RECT 109.975 141.080 110.185 141.900 ;
        RECT 112.735 141.850 114.385 142.370 ;
        RECT 114.555 142.000 115.075 142.540 ;
        RECT 110.875 141.080 114.385 141.850 ;
        RECT 115.245 141.830 115.765 142.370 ;
        RECT 114.555 141.080 115.765 141.830 ;
        RECT 10.510 140.910 115.850 141.080 ;
        RECT 10.595 140.160 11.805 140.910 ;
        RECT 10.595 139.620 11.115 140.160 ;
        RECT 12.435 140.140 15.945 140.910 ;
        RECT 11.285 139.450 11.805 139.990 ;
        RECT 10.595 138.360 11.805 139.450 ;
        RECT 12.435 139.450 14.125 139.970 ;
        RECT 14.295 139.620 15.945 140.140 ;
        RECT 16.155 140.090 16.385 140.910 ;
        RECT 16.555 140.110 16.885 140.740 ;
        RECT 16.135 139.670 16.465 139.920 ;
        RECT 16.635 139.510 16.885 140.110 ;
        RECT 17.055 140.090 17.265 140.910 ;
        RECT 17.955 140.140 19.625 140.910 ;
        RECT 19.800 140.365 25.145 140.910 ;
        RECT 12.435 138.360 15.945 139.450 ;
        RECT 16.155 138.360 16.385 139.500 ;
        RECT 16.555 138.530 16.885 139.510 ;
        RECT 17.055 138.360 17.265 139.500 ;
        RECT 17.955 139.450 18.705 139.970 ;
        RECT 18.875 139.620 19.625 140.140 ;
        RECT 17.955 138.360 19.625 139.450 ;
        RECT 21.390 138.795 21.740 140.045 ;
        RECT 23.220 139.535 23.560 140.365 ;
        RECT 25.315 140.185 25.605 140.910 ;
        RECT 26.235 140.140 28.825 140.910 ;
        RECT 19.800 138.360 25.145 138.795 ;
        RECT 25.315 138.360 25.605 139.525 ;
        RECT 26.235 139.450 27.445 139.970 ;
        RECT 27.615 139.620 28.825 140.140 ;
        RECT 28.995 140.235 29.265 140.580 ;
        RECT 29.455 140.510 29.835 140.910 ;
        RECT 30.005 140.340 30.175 140.690 ;
        RECT 30.345 140.510 30.675 140.910 ;
        RECT 30.875 140.340 31.045 140.690 ;
        RECT 31.245 140.410 31.575 140.910 ;
        RECT 28.995 139.500 29.165 140.235 ;
        RECT 29.435 140.170 31.045 140.340 ;
        RECT 29.435 140.000 29.605 140.170 ;
        RECT 29.335 139.670 29.605 140.000 ;
        RECT 29.775 139.670 30.180 140.000 ;
        RECT 29.435 139.500 29.605 139.670 ;
        RECT 26.235 138.360 28.825 139.450 ;
        RECT 28.995 138.530 29.265 139.500 ;
        RECT 29.435 139.330 30.160 139.500 ;
        RECT 30.350 139.380 31.060 140.000 ;
        RECT 31.230 139.670 31.580 140.240 ;
        RECT 32.215 140.140 34.805 140.910 ;
        RECT 29.990 139.210 30.160 139.330 ;
        RECT 31.260 139.210 31.580 139.500 ;
        RECT 29.475 138.360 29.755 139.160 ;
        RECT 29.990 139.040 31.580 139.210 ;
        RECT 32.215 139.450 33.425 139.970 ;
        RECT 33.595 139.620 34.805 140.140 ;
        RECT 34.975 140.235 35.245 140.580 ;
        RECT 35.435 140.510 35.815 140.910 ;
        RECT 35.985 140.340 36.155 140.690 ;
        RECT 36.325 140.510 36.655 140.910 ;
        RECT 36.855 140.340 37.025 140.690 ;
        RECT 37.225 140.410 37.555 140.910 ;
        RECT 37.745 140.410 38.075 140.910 ;
        RECT 34.975 139.500 35.145 140.235 ;
        RECT 35.415 140.170 37.025 140.340 ;
        RECT 38.275 140.340 38.445 140.690 ;
        RECT 38.645 140.510 38.975 140.910 ;
        RECT 39.145 140.340 39.315 140.690 ;
        RECT 39.485 140.510 39.865 140.910 ;
        RECT 35.415 140.000 35.585 140.170 ;
        RECT 35.315 139.670 35.585 140.000 ;
        RECT 35.755 139.670 36.160 140.000 ;
        RECT 35.415 139.500 35.585 139.670 ;
        RECT 36.330 139.550 37.040 140.000 ;
        RECT 37.210 139.670 37.560 140.240 ;
        RECT 37.740 139.670 38.090 140.240 ;
        RECT 38.275 140.170 39.885 140.340 ;
        RECT 40.055 140.235 40.325 140.580 ;
        RECT 40.505 140.410 40.835 140.910 ;
        RECT 41.035 140.340 41.205 140.690 ;
        RECT 41.405 140.510 41.735 140.910 ;
        RECT 41.905 140.340 42.075 140.690 ;
        RECT 42.245 140.510 42.625 140.910 ;
        RECT 39.715 140.000 39.885 140.170 ;
        RECT 29.925 138.580 31.580 138.870 ;
        RECT 32.215 138.360 34.805 139.450 ;
        RECT 34.975 138.530 35.245 139.500 ;
        RECT 35.415 139.330 36.140 139.500 ;
        RECT 36.330 139.380 37.045 139.550 ;
        RECT 35.970 139.210 36.140 139.330 ;
        RECT 37.240 139.210 37.560 139.500 ;
        RECT 35.455 138.360 35.735 139.160 ;
        RECT 35.970 139.040 37.560 139.210 ;
        RECT 37.740 139.210 38.060 139.500 ;
        RECT 38.260 139.380 38.970 140.000 ;
        RECT 39.140 139.670 39.545 140.000 ;
        RECT 39.715 139.670 39.985 140.000 ;
        RECT 39.715 139.500 39.885 139.670 ;
        RECT 40.155 139.500 40.325 140.235 ;
        RECT 40.500 139.670 40.850 140.240 ;
        RECT 41.035 140.170 42.645 140.340 ;
        RECT 42.815 140.235 43.085 140.580 ;
        RECT 42.475 140.000 42.645 140.170 ;
        RECT 39.160 139.330 39.885 139.500 ;
        RECT 39.160 139.210 39.330 139.330 ;
        RECT 37.740 139.040 39.330 139.210 ;
        RECT 35.905 138.580 37.560 138.870 ;
        RECT 37.740 138.580 39.395 138.870 ;
        RECT 39.565 138.360 39.845 139.160 ;
        RECT 40.055 138.530 40.325 139.500 ;
        RECT 40.500 139.210 40.820 139.500 ;
        RECT 41.020 139.380 41.730 140.000 ;
        RECT 41.900 139.670 42.305 140.000 ;
        RECT 42.475 139.670 42.745 140.000 ;
        RECT 42.475 139.500 42.645 139.670 ;
        RECT 42.915 139.500 43.085 140.235 ;
        RECT 41.920 139.330 42.645 139.500 ;
        RECT 41.920 139.210 42.090 139.330 ;
        RECT 40.500 139.040 42.090 139.210 ;
        RECT 40.500 138.580 42.155 138.870 ;
        RECT 42.325 138.360 42.605 139.160 ;
        RECT 42.815 138.530 43.085 139.500 ;
        RECT 43.255 140.110 43.595 140.740 ;
        RECT 43.765 140.110 44.015 140.910 ;
        RECT 44.205 140.260 44.535 140.740 ;
        RECT 44.705 140.450 44.930 140.910 ;
        RECT 45.100 140.260 45.430 140.740 ;
        RECT 43.255 139.550 43.430 140.110 ;
        RECT 44.205 140.090 45.430 140.260 ;
        RECT 46.060 140.130 46.560 140.740 ;
        RECT 47.395 140.140 50.905 140.910 ;
        RECT 51.075 140.185 51.365 140.910 ;
        RECT 51.535 140.140 53.205 140.910 ;
        RECT 43.600 139.750 44.295 139.920 ;
        RECT 43.255 139.500 43.485 139.550 ;
        RECT 44.125 139.500 44.295 139.750 ;
        RECT 44.470 139.720 44.890 139.920 ;
        RECT 45.060 139.720 45.390 139.920 ;
        RECT 45.560 139.720 45.890 139.920 ;
        RECT 46.060 139.500 46.230 140.130 ;
        RECT 46.415 139.670 46.765 139.920 ;
        RECT 43.255 138.530 43.595 139.500 ;
        RECT 43.765 138.360 43.935 139.500 ;
        RECT 44.125 139.330 46.560 139.500 ;
        RECT 44.205 138.360 44.455 139.160 ;
        RECT 45.100 138.530 45.430 139.330 ;
        RECT 45.730 138.360 46.060 139.160 ;
        RECT 46.230 138.530 46.560 139.330 ;
        RECT 47.395 139.450 49.085 139.970 ;
        RECT 49.255 139.620 50.905 140.140 ;
        RECT 47.395 138.360 50.905 139.450 ;
        RECT 51.075 138.360 51.365 139.525 ;
        RECT 51.535 139.450 52.285 139.970 ;
        RECT 52.455 139.620 53.205 140.140 ;
        RECT 53.490 140.280 53.775 140.740 ;
        RECT 53.945 140.450 54.215 140.910 ;
        RECT 53.490 140.110 54.445 140.280 ;
        RECT 51.535 138.360 53.205 139.450 ;
        RECT 53.375 139.380 54.065 139.940 ;
        RECT 54.235 139.210 54.445 140.110 ;
        RECT 53.490 138.990 54.445 139.210 ;
        RECT 54.615 139.940 55.015 140.740 ;
        RECT 55.205 140.280 55.485 140.740 ;
        RECT 56.005 140.450 56.330 140.910 ;
        RECT 55.205 140.110 56.330 140.280 ;
        RECT 56.500 140.170 56.885 140.740 ;
        RECT 55.880 140.000 56.330 140.110 ;
        RECT 54.615 139.380 55.710 139.940 ;
        RECT 55.880 139.670 56.435 140.000 ;
        RECT 53.490 138.530 53.775 138.990 ;
        RECT 53.945 138.360 54.215 138.820 ;
        RECT 54.615 138.530 55.015 139.380 ;
        RECT 55.880 139.210 56.330 139.670 ;
        RECT 56.605 139.500 56.885 140.170 ;
        RECT 57.790 140.100 58.035 140.705 ;
        RECT 58.255 140.375 58.765 140.910 ;
        RECT 55.205 138.990 56.330 139.210 ;
        RECT 55.205 138.530 55.485 138.990 ;
        RECT 56.005 138.360 56.330 138.820 ;
        RECT 56.500 138.530 56.885 139.500 ;
        RECT 57.515 139.930 58.745 140.100 ;
        RECT 57.515 139.120 57.855 139.930 ;
        RECT 58.025 139.365 58.775 139.555 ;
        RECT 57.515 138.710 58.030 139.120 ;
        RECT 58.265 138.360 58.435 139.120 ;
        RECT 58.605 138.700 58.775 139.365 ;
        RECT 58.945 139.380 59.135 140.740 ;
        RECT 59.305 139.890 59.580 140.740 ;
        RECT 59.770 140.375 60.300 140.740 ;
        RECT 60.725 140.510 61.055 140.910 ;
        RECT 60.125 140.340 60.300 140.375 ;
        RECT 59.305 139.720 59.585 139.890 ;
        RECT 59.305 139.580 59.580 139.720 ;
        RECT 59.785 139.380 59.955 140.180 ;
        RECT 58.945 139.210 59.955 139.380 ;
        RECT 60.125 140.170 61.055 140.340 ;
        RECT 61.225 140.170 61.480 140.740 ;
        RECT 61.745 140.360 61.915 140.740 ;
        RECT 62.095 140.530 62.425 140.910 ;
        RECT 61.745 140.190 62.410 140.360 ;
        RECT 62.605 140.235 62.865 140.740 ;
        RECT 60.125 139.040 60.295 140.170 ;
        RECT 60.885 140.000 61.055 140.170 ;
        RECT 59.170 138.870 60.295 139.040 ;
        RECT 60.465 139.670 60.660 140.000 ;
        RECT 60.885 139.670 61.140 140.000 ;
        RECT 60.465 138.700 60.635 139.670 ;
        RECT 61.310 139.500 61.480 140.170 ;
        RECT 61.675 139.640 62.005 140.010 ;
        RECT 62.240 139.935 62.410 140.190 ;
        RECT 58.605 138.530 60.635 138.700 ;
        RECT 60.805 138.360 60.975 139.500 ;
        RECT 61.145 138.530 61.480 139.500 ;
        RECT 62.240 139.605 62.525 139.935 ;
        RECT 62.240 139.460 62.410 139.605 ;
        RECT 61.745 139.290 62.410 139.460 ;
        RECT 62.695 139.435 62.865 140.235 ;
        RECT 63.495 140.140 66.085 140.910 ;
        RECT 61.745 138.530 61.915 139.290 ;
        RECT 62.095 138.360 62.425 139.120 ;
        RECT 62.595 138.530 62.865 139.435 ;
        RECT 63.495 139.450 64.705 139.970 ;
        RECT 64.875 139.620 66.085 140.140 ;
        RECT 66.255 140.235 66.525 140.580 ;
        RECT 66.715 140.510 67.095 140.910 ;
        RECT 67.265 140.340 67.435 140.690 ;
        RECT 67.605 140.510 67.935 140.910 ;
        RECT 68.135 140.340 68.305 140.690 ;
        RECT 68.505 140.410 68.835 140.910 ;
        RECT 66.255 139.500 66.425 140.235 ;
        RECT 66.695 140.170 68.305 140.340 ;
        RECT 66.695 140.000 66.865 140.170 ;
        RECT 66.595 139.670 66.865 140.000 ;
        RECT 67.035 139.670 67.440 140.000 ;
        RECT 66.695 139.500 66.865 139.670 ;
        RECT 67.610 139.550 68.320 140.000 ;
        RECT 68.490 139.670 68.840 140.240 ;
        RECT 69.015 140.110 69.355 140.740 ;
        RECT 69.525 140.110 69.775 140.910 ;
        RECT 69.965 140.260 70.295 140.740 ;
        RECT 70.465 140.450 70.690 140.910 ;
        RECT 70.860 140.260 71.190 140.740 ;
        RECT 69.015 140.060 69.245 140.110 ;
        RECT 69.965 140.090 71.190 140.260 ;
        RECT 71.820 140.130 72.320 140.740 ;
        RECT 63.495 138.360 66.085 139.450 ;
        RECT 66.255 138.530 66.525 139.500 ;
        RECT 66.695 139.330 67.420 139.500 ;
        RECT 67.610 139.380 68.325 139.550 ;
        RECT 69.015 139.500 69.190 140.060 ;
        RECT 69.360 139.750 70.055 139.920 ;
        RECT 69.885 139.500 70.055 139.750 ;
        RECT 70.230 139.720 70.650 139.920 ;
        RECT 70.820 139.720 71.150 139.920 ;
        RECT 71.320 139.720 71.650 139.920 ;
        RECT 71.820 139.500 71.990 140.130 ;
        RECT 72.970 140.100 73.215 140.705 ;
        RECT 73.435 140.375 73.945 140.910 ;
        RECT 72.695 139.930 73.925 140.100 ;
        RECT 72.175 139.670 72.525 139.920 ;
        RECT 67.250 139.210 67.420 139.330 ;
        RECT 68.520 139.210 68.840 139.500 ;
        RECT 66.735 138.360 67.015 139.160 ;
        RECT 67.250 139.040 68.840 139.210 ;
        RECT 67.185 138.580 68.840 138.870 ;
        RECT 69.015 138.530 69.355 139.500 ;
        RECT 69.525 138.360 69.695 139.500 ;
        RECT 69.885 139.330 72.320 139.500 ;
        RECT 69.965 138.360 70.215 139.160 ;
        RECT 70.860 138.530 71.190 139.330 ;
        RECT 71.490 138.360 71.820 139.160 ;
        RECT 71.990 138.530 72.320 139.330 ;
        RECT 72.695 139.120 73.035 139.930 ;
        RECT 73.205 139.365 73.955 139.555 ;
        RECT 72.695 138.710 73.210 139.120 ;
        RECT 73.445 138.360 73.615 139.120 ;
        RECT 73.785 138.700 73.955 139.365 ;
        RECT 74.125 139.380 74.315 140.740 ;
        RECT 74.485 139.890 74.760 140.740 ;
        RECT 74.950 140.375 75.480 140.740 ;
        RECT 75.905 140.510 76.235 140.910 ;
        RECT 75.305 140.340 75.480 140.375 ;
        RECT 74.485 139.720 74.765 139.890 ;
        RECT 74.485 139.580 74.760 139.720 ;
        RECT 74.965 139.380 75.135 140.180 ;
        RECT 74.125 139.210 75.135 139.380 ;
        RECT 75.305 140.170 76.235 140.340 ;
        RECT 76.405 140.170 76.660 140.740 ;
        RECT 76.835 140.185 77.125 140.910 ;
        RECT 77.845 140.360 78.015 140.740 ;
        RECT 78.195 140.530 78.525 140.910 ;
        RECT 77.845 140.190 78.510 140.360 ;
        RECT 78.705 140.235 78.965 140.740 ;
        RECT 75.305 139.040 75.475 140.170 ;
        RECT 76.065 140.000 76.235 140.170 ;
        RECT 74.350 138.870 75.475 139.040 ;
        RECT 75.645 139.670 75.840 140.000 ;
        RECT 76.065 139.670 76.320 140.000 ;
        RECT 75.645 138.700 75.815 139.670 ;
        RECT 76.490 139.500 76.660 140.170 ;
        RECT 77.775 139.640 78.105 140.010 ;
        RECT 78.340 139.935 78.510 140.190 ;
        RECT 78.340 139.605 78.625 139.935 ;
        RECT 73.785 138.530 75.815 138.700 ;
        RECT 75.985 138.360 76.155 139.500 ;
        RECT 76.325 138.530 76.660 139.500 ;
        RECT 76.835 138.360 77.125 139.525 ;
        RECT 78.340 139.460 78.510 139.605 ;
        RECT 77.845 139.290 78.510 139.460 ;
        RECT 78.795 139.435 78.965 140.235 ;
        RECT 79.195 140.090 79.405 140.910 ;
        RECT 79.575 140.110 79.905 140.740 ;
        RECT 79.575 139.510 79.825 140.110 ;
        RECT 80.075 140.090 80.305 140.910 ;
        RECT 80.515 140.140 83.105 140.910 ;
        RECT 79.995 139.670 80.325 139.920 ;
        RECT 77.845 138.530 78.015 139.290 ;
        RECT 78.195 138.360 78.525 139.120 ;
        RECT 78.695 138.530 78.965 139.435 ;
        RECT 79.195 138.360 79.405 139.500 ;
        RECT 79.575 138.530 79.905 139.510 ;
        RECT 80.075 138.360 80.305 139.500 ;
        RECT 80.515 139.450 81.725 139.970 ;
        RECT 81.895 139.620 83.105 140.140 ;
        RECT 83.550 140.100 83.795 140.705 ;
        RECT 84.015 140.375 84.525 140.910 ;
        RECT 83.275 139.930 84.505 140.100 ;
        RECT 80.515 138.360 83.105 139.450 ;
        RECT 83.275 139.120 83.615 139.930 ;
        RECT 83.785 139.365 84.535 139.555 ;
        RECT 83.275 138.710 83.790 139.120 ;
        RECT 84.025 138.360 84.195 139.120 ;
        RECT 84.365 138.700 84.535 139.365 ;
        RECT 84.705 139.380 84.895 140.740 ;
        RECT 85.065 140.230 85.340 140.740 ;
        RECT 85.530 140.375 86.060 140.740 ;
        RECT 86.485 140.510 86.815 140.910 ;
        RECT 85.885 140.340 86.060 140.375 ;
        RECT 85.065 140.060 85.345 140.230 ;
        RECT 85.065 139.580 85.340 140.060 ;
        RECT 85.545 139.380 85.715 140.180 ;
        RECT 84.705 139.210 85.715 139.380 ;
        RECT 85.885 140.170 86.815 140.340 ;
        RECT 86.985 140.170 87.240 140.740 ;
        RECT 85.885 139.040 86.055 140.170 ;
        RECT 86.645 140.000 86.815 140.170 ;
        RECT 84.930 138.870 86.055 139.040 ;
        RECT 86.225 139.670 86.420 140.000 ;
        RECT 86.645 139.670 86.900 140.000 ;
        RECT 86.225 138.700 86.395 139.670 ;
        RECT 87.070 139.500 87.240 140.170 ;
        RECT 87.415 140.140 89.085 140.910 ;
        RECT 84.365 138.530 86.395 138.700 ;
        RECT 86.565 138.360 86.735 139.500 ;
        RECT 86.905 138.530 87.240 139.500 ;
        RECT 87.415 139.450 88.165 139.970 ;
        RECT 88.335 139.620 89.085 140.140 ;
        RECT 89.255 140.110 89.595 140.740 ;
        RECT 89.765 140.110 90.015 140.910 ;
        RECT 90.205 140.260 90.535 140.740 ;
        RECT 90.705 140.450 90.930 140.910 ;
        RECT 91.100 140.260 91.430 140.740 ;
        RECT 89.255 139.550 89.430 140.110 ;
        RECT 90.205 140.090 91.430 140.260 ;
        RECT 92.060 140.130 92.560 140.740 ;
        RECT 89.600 139.750 90.295 139.920 ;
        RECT 90.470 139.890 90.890 139.920 ;
        RECT 89.255 139.500 89.485 139.550 ;
        RECT 90.125 139.500 90.295 139.750 ;
        RECT 90.465 139.720 90.890 139.890 ;
        RECT 91.060 139.720 91.390 139.920 ;
        RECT 91.560 139.720 91.890 139.920 ;
        RECT 92.060 139.500 92.230 140.130 ;
        RECT 93.210 140.100 93.455 140.705 ;
        RECT 93.675 140.375 94.185 140.910 ;
        RECT 92.935 139.930 94.165 140.100 ;
        RECT 92.415 139.670 92.765 139.920 ;
        RECT 87.415 138.360 89.085 139.450 ;
        RECT 89.255 138.530 89.595 139.500 ;
        RECT 89.765 138.360 89.935 139.500 ;
        RECT 90.125 139.330 92.560 139.500 ;
        RECT 90.205 138.360 90.455 139.160 ;
        RECT 91.100 138.530 91.430 139.330 ;
        RECT 91.730 138.360 92.060 139.160 ;
        RECT 92.230 138.530 92.560 139.330 ;
        RECT 92.935 139.120 93.275 139.930 ;
        RECT 93.445 139.365 94.195 139.555 ;
        RECT 92.935 138.710 93.450 139.120 ;
        RECT 93.685 138.360 93.855 139.120 ;
        RECT 94.025 138.700 94.195 139.365 ;
        RECT 94.365 139.380 94.555 140.740 ;
        RECT 94.725 139.890 95.000 140.740 ;
        RECT 95.190 140.375 95.720 140.740 ;
        RECT 96.145 140.510 96.475 140.910 ;
        RECT 95.545 140.340 95.720 140.375 ;
        RECT 94.725 139.720 95.005 139.890 ;
        RECT 94.725 139.580 95.000 139.720 ;
        RECT 95.205 139.380 95.375 140.180 ;
        RECT 94.365 139.210 95.375 139.380 ;
        RECT 95.545 140.170 96.475 140.340 ;
        RECT 96.645 140.170 96.900 140.740 ;
        RECT 95.545 139.040 95.715 140.170 ;
        RECT 96.305 140.000 96.475 140.170 ;
        RECT 94.590 138.870 95.715 139.040 ;
        RECT 95.885 139.670 96.080 140.000 ;
        RECT 96.305 139.670 96.560 140.000 ;
        RECT 95.885 138.700 96.055 139.670 ;
        RECT 96.730 139.500 96.900 140.170 ;
        RECT 97.075 140.140 98.745 140.910 ;
        RECT 94.025 138.530 96.055 138.700 ;
        RECT 96.225 138.360 96.395 139.500 ;
        RECT 96.565 138.530 96.900 139.500 ;
        RECT 97.075 139.450 97.825 139.970 ;
        RECT 97.995 139.620 98.745 140.140 ;
        RECT 99.120 140.130 99.620 140.740 ;
        RECT 98.915 139.670 99.265 139.920 ;
        RECT 99.450 139.500 99.620 140.130 ;
        RECT 100.250 140.260 100.580 140.740 ;
        RECT 100.750 140.450 100.975 140.910 ;
        RECT 101.145 140.260 101.475 140.740 ;
        RECT 100.250 140.090 101.475 140.260 ;
        RECT 101.665 140.110 101.915 140.910 ;
        RECT 102.085 140.110 102.425 140.740 ;
        RECT 102.595 140.185 102.885 140.910 ;
        RECT 99.790 139.720 100.120 139.920 ;
        RECT 100.290 139.720 100.620 139.920 ;
        RECT 100.790 139.720 101.210 139.920 ;
        RECT 101.385 139.750 102.080 139.920 ;
        RECT 101.385 139.500 101.555 139.750 ;
        RECT 102.250 139.500 102.425 140.110 ;
        RECT 103.555 140.090 103.785 140.910 ;
        RECT 103.955 140.110 104.285 140.740 ;
        RECT 103.535 139.670 103.865 139.920 ;
        RECT 97.075 138.360 98.745 139.450 ;
        RECT 99.120 139.330 101.555 139.500 ;
        RECT 99.120 138.530 99.450 139.330 ;
        RECT 99.620 138.360 99.950 139.160 ;
        RECT 100.250 138.530 100.580 139.330 ;
        RECT 101.225 138.360 101.475 139.160 ;
        RECT 101.745 138.360 101.915 139.500 ;
        RECT 102.085 138.530 102.425 139.500 ;
        RECT 102.595 138.360 102.885 139.525 ;
        RECT 104.035 139.510 104.285 140.110 ;
        RECT 104.455 140.090 104.665 140.910 ;
        RECT 105.270 140.200 105.525 140.730 ;
        RECT 105.705 140.450 105.990 140.910 ;
        RECT 105.270 139.550 105.450 140.200 ;
        RECT 106.170 140.000 106.420 140.650 ;
        RECT 105.620 139.670 106.420 140.000 ;
        RECT 103.555 138.360 103.785 139.500 ;
        RECT 103.955 138.530 104.285 139.510 ;
        RECT 104.455 138.360 104.665 139.500 ;
        RECT 105.185 139.380 105.450 139.550 ;
        RECT 105.270 139.340 105.450 139.380 ;
        RECT 105.270 138.670 105.525 139.340 ;
        RECT 105.705 138.360 105.990 139.160 ;
        RECT 106.170 139.080 106.420 139.670 ;
        RECT 106.620 140.315 106.940 140.645 ;
        RECT 107.120 140.430 107.780 140.910 ;
        RECT 107.980 140.520 108.830 140.690 ;
        RECT 106.620 139.420 106.810 140.315 ;
        RECT 107.130 139.990 107.790 140.260 ;
        RECT 107.460 139.930 107.790 139.990 ;
        RECT 106.980 139.760 107.310 139.820 ;
        RECT 107.980 139.760 108.150 140.520 ;
        RECT 109.390 140.450 109.710 140.910 ;
        RECT 109.910 140.270 110.160 140.700 ;
        RECT 110.450 140.470 110.860 140.910 ;
        RECT 111.030 140.530 112.045 140.730 ;
        RECT 108.320 140.100 109.570 140.270 ;
        RECT 108.320 139.980 108.650 140.100 ;
        RECT 106.980 139.590 108.880 139.760 ;
        RECT 106.620 139.250 108.540 139.420 ;
        RECT 106.620 139.230 106.940 139.250 ;
        RECT 106.170 138.570 106.500 139.080 ;
        RECT 106.770 138.620 106.940 139.230 ;
        RECT 108.710 139.080 108.880 139.590 ;
        RECT 109.050 139.520 109.230 139.930 ;
        RECT 109.400 139.340 109.570 140.100 ;
        RECT 107.110 138.360 107.440 139.050 ;
        RECT 107.670 138.910 108.880 139.080 ;
        RECT 109.050 139.030 109.570 139.340 ;
        RECT 109.740 139.930 110.160 140.270 ;
        RECT 110.450 139.930 110.860 140.260 ;
        RECT 109.740 139.160 109.930 139.930 ;
        RECT 111.030 139.800 111.200 140.530 ;
        RECT 112.345 140.360 112.515 140.690 ;
        RECT 112.685 140.530 113.015 140.910 ;
        RECT 111.370 139.980 111.720 140.350 ;
        RECT 111.030 139.760 111.450 139.800 ;
        RECT 110.100 139.590 111.450 139.760 ;
        RECT 110.100 139.430 110.350 139.590 ;
        RECT 110.860 139.160 111.110 139.420 ;
        RECT 109.740 138.910 111.110 139.160 ;
        RECT 107.670 138.620 107.910 138.910 ;
        RECT 108.710 138.830 108.880 138.910 ;
        RECT 108.110 138.360 108.530 138.740 ;
        RECT 108.710 138.580 109.340 138.830 ;
        RECT 109.810 138.360 110.140 138.740 ;
        RECT 110.310 138.620 110.480 138.910 ;
        RECT 111.280 138.745 111.450 139.590 ;
        RECT 111.900 139.420 112.120 140.290 ;
        RECT 112.345 140.170 113.040 140.360 ;
        RECT 111.620 139.040 112.120 139.420 ;
        RECT 112.290 139.370 112.700 139.990 ;
        RECT 112.870 139.200 113.040 140.170 ;
        RECT 112.345 139.030 113.040 139.200 ;
        RECT 110.660 138.360 111.040 138.740 ;
        RECT 111.280 138.575 112.110 138.745 ;
        RECT 112.345 138.530 112.515 139.030 ;
        RECT 112.685 138.360 113.015 138.860 ;
        RECT 113.230 138.530 113.455 140.650 ;
        RECT 113.625 140.530 113.955 140.910 ;
        RECT 114.125 140.360 114.295 140.650 ;
        RECT 113.630 140.190 114.295 140.360 ;
        RECT 113.630 139.200 113.860 140.190 ;
        RECT 114.555 140.160 115.765 140.910 ;
        RECT 114.030 139.370 114.380 140.020 ;
        RECT 114.555 139.450 115.075 139.990 ;
        RECT 115.245 139.620 115.765 140.160 ;
        RECT 113.630 139.030 114.295 139.200 ;
        RECT 113.625 138.360 113.955 138.860 ;
        RECT 114.125 138.530 114.295 139.030 ;
        RECT 114.555 138.360 115.765 139.450 ;
        RECT 10.510 138.190 115.850 138.360 ;
        RECT 10.595 137.100 11.805 138.190 ;
        RECT 10.595 136.390 11.115 136.930 ;
        RECT 11.285 136.560 11.805 137.100 ;
        RECT 12.435 137.025 12.725 138.190 ;
        RECT 12.985 137.520 13.155 138.020 ;
        RECT 13.325 137.690 13.655 138.190 ;
        RECT 12.985 137.350 13.650 137.520 ;
        RECT 12.900 136.530 13.250 137.180 ;
        RECT 10.595 135.640 11.805 136.390 ;
        RECT 12.435 135.640 12.725 136.365 ;
        RECT 13.420 136.360 13.650 137.350 ;
        RECT 12.985 136.190 13.650 136.360 ;
        RECT 12.985 135.900 13.155 136.190 ;
        RECT 13.325 135.640 13.655 136.020 ;
        RECT 13.825 135.900 14.050 138.020 ;
        RECT 14.265 137.690 14.595 138.190 ;
        RECT 14.765 137.520 14.935 138.020 ;
        RECT 15.170 137.805 16.000 137.975 ;
        RECT 16.240 137.810 16.620 138.190 ;
        RECT 14.240 137.350 14.935 137.520 ;
        RECT 14.240 136.380 14.410 137.350 ;
        RECT 14.580 136.560 14.990 137.180 ;
        RECT 15.160 137.130 15.660 137.510 ;
        RECT 14.240 136.190 14.935 136.380 ;
        RECT 15.160 136.260 15.380 137.130 ;
        RECT 15.830 136.960 16.000 137.805 ;
        RECT 16.800 137.640 16.970 137.930 ;
        RECT 17.140 137.810 17.470 138.190 ;
        RECT 17.940 137.720 18.570 137.970 ;
        RECT 18.750 137.810 19.170 138.190 ;
        RECT 18.400 137.640 18.570 137.720 ;
        RECT 19.370 137.640 19.610 137.930 ;
        RECT 16.170 137.390 17.540 137.640 ;
        RECT 16.170 137.130 16.420 137.390 ;
        RECT 16.930 136.960 17.180 137.120 ;
        RECT 15.830 136.790 17.180 136.960 ;
        RECT 15.830 136.750 16.250 136.790 ;
        RECT 15.560 136.200 15.910 136.570 ;
        RECT 14.265 135.640 14.595 136.020 ;
        RECT 14.765 135.860 14.935 136.190 ;
        RECT 16.080 136.020 16.250 136.750 ;
        RECT 17.350 136.620 17.540 137.390 ;
        RECT 16.420 136.290 16.830 136.620 ;
        RECT 17.120 136.280 17.540 136.620 ;
        RECT 17.710 137.210 18.230 137.520 ;
        RECT 18.400 137.470 19.610 137.640 ;
        RECT 19.840 137.500 20.170 138.190 ;
        RECT 17.710 136.450 17.880 137.210 ;
        RECT 18.050 136.620 18.230 137.030 ;
        RECT 18.400 136.960 18.570 137.470 ;
        RECT 20.340 137.320 20.510 137.930 ;
        RECT 20.780 137.470 21.110 137.980 ;
        RECT 20.340 137.300 20.660 137.320 ;
        RECT 18.740 137.130 20.660 137.300 ;
        RECT 18.400 136.790 20.300 136.960 ;
        RECT 18.630 136.450 18.960 136.570 ;
        RECT 17.710 136.280 18.960 136.450 ;
        RECT 15.235 135.820 16.250 136.020 ;
        RECT 16.420 135.640 16.830 136.080 ;
        RECT 17.120 135.850 17.370 136.280 ;
        RECT 17.570 135.640 17.890 136.100 ;
        RECT 19.130 136.030 19.300 136.790 ;
        RECT 19.970 136.730 20.300 136.790 ;
        RECT 19.490 136.560 19.820 136.620 ;
        RECT 19.490 136.290 20.150 136.560 ;
        RECT 20.470 136.235 20.660 137.130 ;
        RECT 18.450 135.860 19.300 136.030 ;
        RECT 19.500 135.640 20.160 136.120 ;
        RECT 20.340 135.905 20.660 136.235 ;
        RECT 20.860 136.880 21.110 137.470 ;
        RECT 21.290 137.390 21.575 138.190 ;
        RECT 21.755 137.210 22.010 137.880 ;
        RECT 20.860 136.550 21.660 136.880 ;
        RECT 20.860 135.900 21.110 136.550 ;
        RECT 21.830 136.350 22.010 137.210 ;
        RECT 22.555 137.100 25.145 138.190 ;
        RECT 25.315 137.115 25.585 138.020 ;
        RECT 25.755 137.430 26.085 138.190 ;
        RECT 26.265 137.260 26.435 138.020 ;
        RECT 27.815 137.520 28.095 138.190 ;
        RECT 22.555 136.580 23.765 137.100 ;
        RECT 23.935 136.410 25.145 136.930 ;
        RECT 21.755 136.150 22.010 136.350 ;
        RECT 21.290 135.640 21.575 136.100 ;
        RECT 21.755 135.980 22.095 136.150 ;
        RECT 21.755 135.820 22.010 135.980 ;
        RECT 22.555 135.640 25.145 136.410 ;
        RECT 25.315 136.315 25.485 137.115 ;
        RECT 25.770 137.090 26.435 137.260 ;
        RECT 28.265 137.300 28.565 137.850 ;
        RECT 28.765 137.470 29.095 138.190 ;
        RECT 29.285 137.470 29.745 138.020 ;
        RECT 25.770 136.945 25.940 137.090 ;
        RECT 25.655 136.615 25.940 136.945 ;
        RECT 25.770 136.360 25.940 136.615 ;
        RECT 26.175 136.540 26.505 136.910 ;
        RECT 27.630 136.880 27.895 137.240 ;
        RECT 28.265 137.130 29.205 137.300 ;
        RECT 29.035 136.880 29.205 137.130 ;
        RECT 27.630 136.630 28.305 136.880 ;
        RECT 28.525 136.630 28.865 136.880 ;
        RECT 29.035 136.550 29.325 136.880 ;
        RECT 29.035 136.460 29.205 136.550 ;
        RECT 25.315 135.810 25.575 136.315 ;
        RECT 25.770 136.190 26.435 136.360 ;
        RECT 25.755 135.640 26.085 136.020 ;
        RECT 26.265 135.810 26.435 136.190 ;
        RECT 27.815 136.270 29.205 136.460 ;
        RECT 27.815 135.910 28.145 136.270 ;
        RECT 29.495 136.100 29.745 137.470 ;
        RECT 28.765 135.640 29.015 136.100 ;
        RECT 29.185 135.810 29.745 136.100 ;
        RECT 29.915 137.050 30.185 138.020 ;
        RECT 30.395 137.390 30.675 138.190 ;
        RECT 30.845 137.680 32.500 137.970 ;
        RECT 30.910 137.340 32.500 137.510 ;
        RECT 30.910 137.220 31.080 137.340 ;
        RECT 30.355 137.050 31.080 137.220 ;
        RECT 29.915 136.315 30.085 137.050 ;
        RECT 30.355 136.880 30.525 137.050 ;
        RECT 30.255 136.550 30.525 136.880 ;
        RECT 30.695 136.550 31.100 136.880 ;
        RECT 31.270 136.550 31.980 137.170 ;
        RECT 32.180 137.050 32.500 137.340 ;
        RECT 33.135 137.050 33.405 138.020 ;
        RECT 33.615 137.390 33.895 138.190 ;
        RECT 34.065 137.680 35.720 137.970 ;
        RECT 34.130 137.340 35.720 137.510 ;
        RECT 34.130 137.220 34.300 137.340 ;
        RECT 33.575 137.050 34.300 137.220 ;
        RECT 30.355 136.380 30.525 136.550 ;
        RECT 29.915 135.970 30.185 136.315 ;
        RECT 30.355 136.210 31.965 136.380 ;
        RECT 32.150 136.310 32.500 136.880 ;
        RECT 33.135 136.315 33.305 137.050 ;
        RECT 33.575 136.880 33.745 137.050 ;
        RECT 34.490 137.000 35.205 137.170 ;
        RECT 35.400 137.050 35.720 137.340 ;
        RECT 36.355 137.100 38.025 138.190 ;
        RECT 33.475 136.550 33.745 136.880 ;
        RECT 33.915 136.550 34.320 136.880 ;
        RECT 34.490 136.550 35.200 137.000 ;
        RECT 33.575 136.380 33.745 136.550 ;
        RECT 30.375 135.640 30.755 136.040 ;
        RECT 30.925 135.860 31.095 136.210 ;
        RECT 31.265 135.640 31.595 136.040 ;
        RECT 31.795 135.860 31.965 136.210 ;
        RECT 32.165 135.640 32.495 136.140 ;
        RECT 33.135 135.970 33.405 136.315 ;
        RECT 33.575 136.210 35.185 136.380 ;
        RECT 35.370 136.310 35.720 136.880 ;
        RECT 36.355 136.580 37.105 137.100 ;
        RECT 38.195 137.025 38.485 138.190 ;
        RECT 38.660 137.755 44.005 138.190 ;
        RECT 37.275 136.410 38.025 136.930 ;
        RECT 40.250 136.505 40.600 137.755 ;
        RECT 44.175 137.115 44.445 138.020 ;
        RECT 44.615 137.430 44.945 138.190 ;
        RECT 45.125 137.260 45.295 138.020 ;
        RECT 33.595 135.640 33.975 136.040 ;
        RECT 34.145 135.860 34.315 136.210 ;
        RECT 34.485 135.640 34.815 136.040 ;
        RECT 35.015 135.860 35.185 136.210 ;
        RECT 35.385 135.640 35.715 136.140 ;
        RECT 36.355 135.640 38.025 136.410 ;
        RECT 38.195 135.640 38.485 136.365 ;
        RECT 42.080 136.185 42.420 137.015 ;
        RECT 44.175 136.315 44.345 137.115 ;
        RECT 44.630 137.090 45.295 137.260 ;
        RECT 44.630 136.945 44.800 137.090 ;
        RECT 44.515 136.615 44.800 136.945 ;
        RECT 45.560 137.050 45.895 138.020 ;
        RECT 46.065 137.050 46.235 138.190 ;
        RECT 46.405 137.850 48.435 138.020 ;
        RECT 44.630 136.360 44.800 136.615 ;
        RECT 45.035 136.540 45.365 136.910 ;
        RECT 45.560 136.380 45.730 137.050 ;
        RECT 46.405 136.880 46.575 137.850 ;
        RECT 45.900 136.550 46.155 136.880 ;
        RECT 46.380 136.550 46.575 136.880 ;
        RECT 46.745 137.510 47.870 137.680 ;
        RECT 45.985 136.380 46.155 136.550 ;
        RECT 46.745 136.380 46.915 137.510 ;
        RECT 38.660 135.640 44.005 136.185 ;
        RECT 44.175 135.810 44.435 136.315 ;
        RECT 44.630 136.190 45.295 136.360 ;
        RECT 44.615 135.640 44.945 136.020 ;
        RECT 45.125 135.810 45.295 136.190 ;
        RECT 45.560 135.810 45.815 136.380 ;
        RECT 45.985 136.210 46.915 136.380 ;
        RECT 47.085 137.170 48.095 137.340 ;
        RECT 47.085 136.370 47.255 137.170 ;
        RECT 47.460 136.830 47.735 136.970 ;
        RECT 47.455 136.660 47.735 136.830 ;
        RECT 46.740 136.175 46.915 136.210 ;
        RECT 45.985 135.640 46.315 136.040 ;
        RECT 46.740 135.810 47.270 136.175 ;
        RECT 47.460 135.810 47.735 136.660 ;
        RECT 47.905 135.810 48.095 137.170 ;
        RECT 48.265 137.185 48.435 137.850 ;
        RECT 48.605 137.430 48.775 138.190 ;
        RECT 49.010 137.430 49.525 137.840 ;
        RECT 48.265 136.995 49.015 137.185 ;
        RECT 49.185 136.620 49.525 137.430 ;
        RECT 48.295 136.450 49.525 136.620 ;
        RECT 49.695 137.050 50.035 138.020 ;
        RECT 50.205 137.050 50.375 138.190 ;
        RECT 50.645 137.390 50.895 138.190 ;
        RECT 51.540 137.220 51.870 138.020 ;
        RECT 52.170 137.390 52.500 138.190 ;
        RECT 52.670 137.220 53.000 138.020 ;
        RECT 50.565 137.050 53.000 137.220 ;
        RECT 53.375 137.050 53.715 138.020 ;
        RECT 53.885 137.050 54.055 138.190 ;
        RECT 54.325 137.390 54.575 138.190 ;
        RECT 55.220 137.220 55.550 138.020 ;
        RECT 55.850 137.390 56.180 138.190 ;
        RECT 56.350 137.220 56.680 138.020 ;
        RECT 54.245 137.050 56.680 137.220 ;
        RECT 57.055 137.100 58.725 138.190 ;
        RECT 48.275 135.640 48.785 136.175 ;
        RECT 49.005 135.845 49.250 136.450 ;
        RECT 49.695 136.440 49.870 137.050 ;
        RECT 50.565 136.800 50.735 137.050 ;
        RECT 50.040 136.630 50.735 136.800 ;
        RECT 50.910 136.630 51.330 136.830 ;
        RECT 51.500 136.630 51.830 136.830 ;
        RECT 52.000 136.630 52.330 136.830 ;
        RECT 49.695 135.810 50.035 136.440 ;
        RECT 50.205 135.640 50.455 136.440 ;
        RECT 50.645 136.290 51.870 136.460 ;
        RECT 50.645 135.810 50.975 136.290 ;
        RECT 51.145 135.640 51.370 136.100 ;
        RECT 51.540 135.810 51.870 136.290 ;
        RECT 52.500 136.420 52.670 137.050 ;
        RECT 52.855 136.630 53.205 136.880 ;
        RECT 53.375 136.440 53.550 137.050 ;
        RECT 54.245 136.800 54.415 137.050 ;
        RECT 53.720 136.630 54.415 136.800 ;
        RECT 54.590 136.630 55.010 136.830 ;
        RECT 55.180 136.630 55.510 136.830 ;
        RECT 55.680 136.630 56.010 136.830 ;
        RECT 52.500 135.810 53.000 136.420 ;
        RECT 53.375 135.810 53.715 136.440 ;
        RECT 53.885 135.640 54.135 136.440 ;
        RECT 54.325 136.290 55.550 136.460 ;
        RECT 54.325 135.810 54.655 136.290 ;
        RECT 54.825 135.640 55.050 136.100 ;
        RECT 55.220 135.810 55.550 136.290 ;
        RECT 56.180 136.420 56.350 137.050 ;
        RECT 56.535 136.630 56.885 136.880 ;
        RECT 57.055 136.580 57.805 137.100 ;
        RECT 58.935 137.050 59.165 138.190 ;
        RECT 59.335 137.040 59.665 138.020 ;
        RECT 59.835 137.050 60.045 138.190 ;
        RECT 60.280 137.800 60.615 138.020 ;
        RECT 61.620 137.810 61.975 138.190 ;
        RECT 60.280 137.180 60.535 137.800 ;
        RECT 60.785 137.640 61.015 137.680 ;
        RECT 62.145 137.640 62.395 138.020 ;
        RECT 60.785 137.440 62.395 137.640 ;
        RECT 60.785 137.350 60.970 137.440 ;
        RECT 61.560 137.430 62.395 137.440 ;
        RECT 62.645 137.410 62.895 138.190 ;
        RECT 63.065 137.340 63.325 138.020 ;
        RECT 61.125 137.240 61.455 137.270 ;
        RECT 61.125 137.180 62.925 137.240 ;
        RECT 60.280 137.070 62.985 137.180 ;
        RECT 56.180 135.810 56.680 136.420 ;
        RECT 57.975 136.410 58.725 136.930 ;
        RECT 58.915 136.630 59.245 136.880 ;
        RECT 57.055 135.640 58.725 136.410 ;
        RECT 58.935 135.640 59.165 136.460 ;
        RECT 59.415 136.440 59.665 137.040 ;
        RECT 60.280 137.010 61.455 137.070 ;
        RECT 62.785 137.035 62.985 137.070 ;
        RECT 60.275 136.630 60.765 136.830 ;
        RECT 60.955 136.630 61.430 136.840 ;
        RECT 59.335 135.810 59.665 136.440 ;
        RECT 59.835 135.640 60.045 136.460 ;
        RECT 60.280 135.640 60.735 136.405 ;
        RECT 61.210 136.230 61.430 136.630 ;
        RECT 61.675 136.630 62.005 136.840 ;
        RECT 61.675 136.230 61.885 136.630 ;
        RECT 62.175 136.595 62.585 136.900 ;
        RECT 62.815 136.460 62.985 137.035 ;
        RECT 62.715 136.340 62.985 136.460 ;
        RECT 62.140 136.295 62.985 136.340 ;
        RECT 62.140 136.170 62.895 136.295 ;
        RECT 62.140 136.020 62.310 136.170 ;
        RECT 63.155 136.150 63.325 137.340 ;
        RECT 63.955 137.025 64.245 138.190 ;
        RECT 64.875 137.100 67.465 138.190 ;
        RECT 67.640 137.755 72.985 138.190 ;
        RECT 73.160 137.755 78.505 138.190 ;
        RECT 79.050 137.850 79.305 137.880 ;
        RECT 64.875 136.580 66.085 137.100 ;
        RECT 66.255 136.410 67.465 136.930 ;
        RECT 69.230 136.505 69.580 137.755 ;
        RECT 63.095 136.140 63.325 136.150 ;
        RECT 61.010 135.810 62.310 136.020 ;
        RECT 62.565 135.640 62.895 136.000 ;
        RECT 63.065 135.810 63.325 136.140 ;
        RECT 63.955 135.640 64.245 136.365 ;
        RECT 64.875 135.640 67.465 136.410 ;
        RECT 71.060 136.185 71.400 137.015 ;
        RECT 74.750 136.505 75.100 137.755 ;
        RECT 78.965 137.680 79.305 137.850 ;
        RECT 79.050 137.210 79.305 137.680 ;
        RECT 79.485 137.390 79.770 138.190 ;
        RECT 79.950 137.470 80.280 137.980 ;
        RECT 76.580 136.185 76.920 137.015 ;
        RECT 79.050 136.350 79.230 137.210 ;
        RECT 79.950 136.880 80.200 137.470 ;
        RECT 80.550 137.320 80.720 137.930 ;
        RECT 80.890 137.500 81.220 138.190 ;
        RECT 81.450 137.640 81.690 137.930 ;
        RECT 81.890 137.810 82.310 138.190 ;
        RECT 82.490 137.720 83.120 137.970 ;
        RECT 83.590 137.810 83.920 138.190 ;
        RECT 82.490 137.640 82.660 137.720 ;
        RECT 84.090 137.640 84.260 137.930 ;
        RECT 84.440 137.810 84.820 138.190 ;
        RECT 85.060 137.805 85.890 137.975 ;
        RECT 81.450 137.470 82.660 137.640 ;
        RECT 79.400 136.550 80.200 136.880 ;
        RECT 67.640 135.640 72.985 136.185 ;
        RECT 73.160 135.640 78.505 136.185 ;
        RECT 79.050 135.820 79.305 136.350 ;
        RECT 79.485 135.640 79.770 136.100 ;
        RECT 79.950 135.900 80.200 136.550 ;
        RECT 80.400 137.300 80.720 137.320 ;
        RECT 80.400 137.130 82.320 137.300 ;
        RECT 80.400 136.235 80.590 137.130 ;
        RECT 82.490 136.960 82.660 137.470 ;
        RECT 82.830 137.210 83.350 137.520 ;
        RECT 80.760 136.790 82.660 136.960 ;
        RECT 80.760 136.730 81.090 136.790 ;
        RECT 81.240 136.560 81.570 136.620 ;
        RECT 80.910 136.290 81.570 136.560 ;
        RECT 80.400 135.905 80.720 136.235 ;
        RECT 80.900 135.640 81.560 136.120 ;
        RECT 81.760 136.030 81.930 136.790 ;
        RECT 82.830 136.620 83.010 137.030 ;
        RECT 82.100 136.450 82.430 136.570 ;
        RECT 83.180 136.450 83.350 137.210 ;
        RECT 82.100 136.280 83.350 136.450 ;
        RECT 83.520 137.390 84.890 137.640 ;
        RECT 83.520 136.620 83.710 137.390 ;
        RECT 84.640 137.130 84.890 137.390 ;
        RECT 83.880 136.960 84.130 137.120 ;
        RECT 85.060 136.960 85.230 137.805 ;
        RECT 86.125 137.520 86.295 138.020 ;
        RECT 86.465 137.690 86.795 138.190 ;
        RECT 85.400 137.130 85.900 137.510 ;
        RECT 86.125 137.350 86.820 137.520 ;
        RECT 83.880 136.790 85.230 136.960 ;
        RECT 84.810 136.750 85.230 136.790 ;
        RECT 83.520 136.280 83.940 136.620 ;
        RECT 84.230 136.290 84.640 136.620 ;
        RECT 81.760 135.860 82.610 136.030 ;
        RECT 83.170 135.640 83.490 136.100 ;
        RECT 83.690 135.850 83.940 136.280 ;
        RECT 84.230 135.640 84.640 136.080 ;
        RECT 84.810 136.020 84.980 136.750 ;
        RECT 85.150 136.200 85.500 136.570 ;
        RECT 85.680 136.260 85.900 137.130 ;
        RECT 86.070 136.560 86.480 137.180 ;
        RECT 86.650 136.380 86.820 137.350 ;
        RECT 86.125 136.190 86.820 136.380 ;
        RECT 84.810 135.820 85.825 136.020 ;
        RECT 86.125 135.860 86.295 136.190 ;
        RECT 86.465 135.640 86.795 136.020 ;
        RECT 87.010 135.900 87.235 138.020 ;
        RECT 87.405 137.690 87.735 138.190 ;
        RECT 87.905 137.520 88.075 138.020 ;
        RECT 87.410 137.350 88.075 137.520 ;
        RECT 87.410 136.360 87.640 137.350 ;
        RECT 87.810 136.530 88.160 137.180 ;
        RECT 88.335 137.115 88.605 138.020 ;
        RECT 88.775 137.430 89.105 138.190 ;
        RECT 89.285 137.260 89.455 138.020 ;
        RECT 87.410 136.190 88.075 136.360 ;
        RECT 87.405 135.640 87.735 136.020 ;
        RECT 87.905 135.900 88.075 136.190 ;
        RECT 88.335 136.315 88.505 137.115 ;
        RECT 88.790 137.090 89.455 137.260 ;
        RECT 88.790 136.945 88.960 137.090 ;
        RECT 89.715 137.025 90.005 138.190 ;
        RECT 90.550 137.850 90.805 137.880 ;
        RECT 90.465 137.680 90.805 137.850 ;
        RECT 90.550 137.210 90.805 137.680 ;
        RECT 90.985 137.390 91.270 138.190 ;
        RECT 91.450 137.470 91.780 137.980 ;
        RECT 88.675 136.615 88.960 136.945 ;
        RECT 88.790 136.360 88.960 136.615 ;
        RECT 89.195 136.540 89.525 136.910 ;
        RECT 88.335 135.810 88.595 136.315 ;
        RECT 88.790 136.190 89.455 136.360 ;
        RECT 88.775 135.640 89.105 136.020 ;
        RECT 89.285 135.810 89.455 136.190 ;
        RECT 89.715 135.640 90.005 136.365 ;
        RECT 90.550 136.350 90.730 137.210 ;
        RECT 91.450 136.880 91.700 137.470 ;
        RECT 92.050 137.320 92.220 137.930 ;
        RECT 92.390 137.500 92.720 138.190 ;
        RECT 92.950 137.640 93.190 137.930 ;
        RECT 93.390 137.810 93.810 138.190 ;
        RECT 93.990 137.720 94.620 137.970 ;
        RECT 95.090 137.810 95.420 138.190 ;
        RECT 93.990 137.640 94.160 137.720 ;
        RECT 95.590 137.640 95.760 137.930 ;
        RECT 95.940 137.810 96.320 138.190 ;
        RECT 96.560 137.805 97.390 137.975 ;
        RECT 92.950 137.470 94.160 137.640 ;
        RECT 90.900 136.550 91.700 136.880 ;
        RECT 90.550 135.820 90.805 136.350 ;
        RECT 90.985 135.640 91.270 136.100 ;
        RECT 91.450 135.900 91.700 136.550 ;
        RECT 91.900 137.300 92.220 137.320 ;
        RECT 91.900 137.130 93.820 137.300 ;
        RECT 91.900 136.235 92.090 137.130 ;
        RECT 93.990 136.960 94.160 137.470 ;
        RECT 94.330 137.210 94.850 137.520 ;
        RECT 92.260 136.790 94.160 136.960 ;
        RECT 92.260 136.730 92.590 136.790 ;
        RECT 92.740 136.560 93.070 136.620 ;
        RECT 92.410 136.290 93.070 136.560 ;
        RECT 91.900 135.905 92.220 136.235 ;
        RECT 92.400 135.640 93.060 136.120 ;
        RECT 93.260 136.030 93.430 136.790 ;
        RECT 94.330 136.620 94.510 137.030 ;
        RECT 93.600 136.450 93.930 136.570 ;
        RECT 94.680 136.450 94.850 137.210 ;
        RECT 93.600 136.280 94.850 136.450 ;
        RECT 95.020 137.390 96.390 137.640 ;
        RECT 95.020 136.620 95.210 137.390 ;
        RECT 96.140 137.130 96.390 137.390 ;
        RECT 95.380 136.960 95.630 137.120 ;
        RECT 96.560 136.960 96.730 137.805 ;
        RECT 97.625 137.520 97.795 138.020 ;
        RECT 97.965 137.690 98.295 138.190 ;
        RECT 96.900 137.130 97.400 137.510 ;
        RECT 97.625 137.350 98.320 137.520 ;
        RECT 95.380 136.790 96.730 136.960 ;
        RECT 96.310 136.750 96.730 136.790 ;
        RECT 95.020 136.280 95.440 136.620 ;
        RECT 95.730 136.290 96.140 136.620 ;
        RECT 93.260 135.860 94.110 136.030 ;
        RECT 94.670 135.640 94.990 136.100 ;
        RECT 95.190 135.850 95.440 136.280 ;
        RECT 95.730 135.640 96.140 136.080 ;
        RECT 96.310 136.020 96.480 136.750 ;
        RECT 96.650 136.200 97.000 136.570 ;
        RECT 97.180 136.260 97.400 137.130 ;
        RECT 97.570 136.560 97.980 137.180 ;
        RECT 98.150 136.380 98.320 137.350 ;
        RECT 97.625 136.190 98.320 136.380 ;
        RECT 96.310 135.820 97.325 136.020 ;
        RECT 97.625 135.860 97.795 136.190 ;
        RECT 97.965 135.640 98.295 136.020 ;
        RECT 98.510 135.900 98.735 138.020 ;
        RECT 98.905 137.690 99.235 138.190 ;
        RECT 99.405 137.520 99.575 138.020 ;
        RECT 98.910 137.350 99.575 137.520 ;
        RECT 98.910 136.360 99.140 137.350 ;
        RECT 99.310 136.530 99.660 137.180 ;
        RECT 99.835 137.115 100.105 138.020 ;
        RECT 100.275 137.430 100.605 138.190 ;
        RECT 100.785 137.260 100.955 138.020 ;
        RECT 102.510 137.850 102.765 137.880 ;
        RECT 102.425 137.680 102.765 137.850 ;
        RECT 98.910 136.190 99.575 136.360 ;
        RECT 98.905 135.640 99.235 136.020 ;
        RECT 99.405 135.900 99.575 136.190 ;
        RECT 99.835 136.315 100.005 137.115 ;
        RECT 100.290 137.090 100.955 137.260 ;
        RECT 102.510 137.210 102.765 137.680 ;
        RECT 102.945 137.390 103.230 138.190 ;
        RECT 103.410 137.470 103.740 137.980 ;
        RECT 100.290 136.945 100.460 137.090 ;
        RECT 100.175 136.615 100.460 136.945 ;
        RECT 100.290 136.360 100.460 136.615 ;
        RECT 100.695 136.540 101.025 136.910 ;
        RECT 99.835 135.810 100.095 136.315 ;
        RECT 100.290 136.190 100.955 136.360 ;
        RECT 100.275 135.640 100.605 136.020 ;
        RECT 100.785 135.810 100.955 136.190 ;
        RECT 102.510 136.350 102.690 137.210 ;
        RECT 103.410 136.880 103.660 137.470 ;
        RECT 104.010 137.320 104.180 137.930 ;
        RECT 104.350 137.500 104.680 138.190 ;
        RECT 104.910 137.640 105.150 137.930 ;
        RECT 105.350 137.810 105.770 138.190 ;
        RECT 105.950 137.720 106.580 137.970 ;
        RECT 107.050 137.810 107.380 138.190 ;
        RECT 105.950 137.640 106.120 137.720 ;
        RECT 107.550 137.640 107.720 137.930 ;
        RECT 107.900 137.810 108.280 138.190 ;
        RECT 108.520 137.805 109.350 137.975 ;
        RECT 104.910 137.470 106.120 137.640 ;
        RECT 102.860 136.550 103.660 136.880 ;
        RECT 102.510 135.820 102.765 136.350 ;
        RECT 102.945 135.640 103.230 136.100 ;
        RECT 103.410 135.900 103.660 136.550 ;
        RECT 103.860 137.300 104.180 137.320 ;
        RECT 103.860 137.130 105.780 137.300 ;
        RECT 103.860 136.235 104.050 137.130 ;
        RECT 105.950 136.960 106.120 137.470 ;
        RECT 106.290 137.210 106.810 137.520 ;
        RECT 104.220 136.790 106.120 136.960 ;
        RECT 104.220 136.730 104.550 136.790 ;
        RECT 104.700 136.560 105.030 136.620 ;
        RECT 104.370 136.290 105.030 136.560 ;
        RECT 103.860 135.905 104.180 136.235 ;
        RECT 104.360 135.640 105.020 136.120 ;
        RECT 105.220 136.030 105.390 136.790 ;
        RECT 106.290 136.620 106.470 137.030 ;
        RECT 105.560 136.450 105.890 136.570 ;
        RECT 106.640 136.450 106.810 137.210 ;
        RECT 105.560 136.280 106.810 136.450 ;
        RECT 106.980 137.390 108.350 137.640 ;
        RECT 106.980 136.620 107.170 137.390 ;
        RECT 108.100 137.130 108.350 137.390 ;
        RECT 107.340 136.960 107.590 137.120 ;
        RECT 108.520 136.960 108.690 137.805 ;
        RECT 109.585 137.520 109.755 138.020 ;
        RECT 109.925 137.690 110.255 138.190 ;
        RECT 108.860 137.130 109.360 137.510 ;
        RECT 109.585 137.350 110.280 137.520 ;
        RECT 107.340 136.790 108.690 136.960 ;
        RECT 108.270 136.750 108.690 136.790 ;
        RECT 106.980 136.280 107.400 136.620 ;
        RECT 107.690 136.290 108.100 136.620 ;
        RECT 105.220 135.860 106.070 136.030 ;
        RECT 106.630 135.640 106.950 136.100 ;
        RECT 107.150 135.850 107.400 136.280 ;
        RECT 107.690 135.640 108.100 136.080 ;
        RECT 108.270 136.020 108.440 136.750 ;
        RECT 108.610 136.200 108.960 136.570 ;
        RECT 109.140 136.260 109.360 137.130 ;
        RECT 109.530 136.560 109.940 137.180 ;
        RECT 110.110 136.380 110.280 137.350 ;
        RECT 109.585 136.190 110.280 136.380 ;
        RECT 108.270 135.820 109.285 136.020 ;
        RECT 109.585 135.860 109.755 136.190 ;
        RECT 109.925 135.640 110.255 136.020 ;
        RECT 110.470 135.900 110.695 138.020 ;
        RECT 110.865 137.690 111.195 138.190 ;
        RECT 111.365 137.520 111.535 138.020 ;
        RECT 110.870 137.350 111.535 137.520 ;
        RECT 110.870 136.360 111.100 137.350 ;
        RECT 111.885 137.260 112.055 138.020 ;
        RECT 112.235 137.430 112.565 138.190 ;
        RECT 111.270 136.530 111.620 137.180 ;
        RECT 111.885 137.090 112.550 137.260 ;
        RECT 112.735 137.115 113.005 138.020 ;
        RECT 112.380 136.945 112.550 137.090 ;
        RECT 111.815 136.540 112.145 136.910 ;
        RECT 112.380 136.615 112.665 136.945 ;
        RECT 112.380 136.360 112.550 136.615 ;
        RECT 110.870 136.190 111.535 136.360 ;
        RECT 110.865 135.640 111.195 136.020 ;
        RECT 111.365 135.900 111.535 136.190 ;
        RECT 111.885 136.190 112.550 136.360 ;
        RECT 112.835 136.315 113.005 137.115 ;
        RECT 113.175 137.100 114.385 138.190 ;
        RECT 114.555 137.100 115.765 138.190 ;
        RECT 113.175 136.560 113.695 137.100 ;
        RECT 113.865 136.390 114.385 136.930 ;
        RECT 114.555 136.560 115.075 137.100 ;
        RECT 115.245 136.390 115.765 136.930 ;
        RECT 111.885 135.810 112.055 136.190 ;
        RECT 112.235 135.640 112.565 136.020 ;
        RECT 112.745 135.810 113.005 136.315 ;
        RECT 113.175 135.640 114.385 136.390 ;
        RECT 114.555 135.640 115.765 136.390 ;
        RECT 10.510 135.470 115.850 135.640 ;
        RECT 10.595 134.720 11.805 135.470 ;
        RECT 12.985 134.920 13.155 135.300 ;
        RECT 13.335 135.090 13.665 135.470 ;
        RECT 12.985 134.750 13.650 134.920 ;
        RECT 13.845 134.795 14.105 135.300 ;
        RECT 10.595 134.180 11.115 134.720 ;
        RECT 11.285 134.010 11.805 134.550 ;
        RECT 12.915 134.200 13.245 134.570 ;
        RECT 13.480 134.495 13.650 134.750 ;
        RECT 13.480 134.165 13.765 134.495 ;
        RECT 13.480 134.020 13.650 134.165 ;
        RECT 10.595 132.920 11.805 134.010 ;
        RECT 12.985 133.850 13.650 134.020 ;
        RECT 13.935 133.995 14.105 134.795 ;
        RECT 14.315 134.650 14.545 135.470 ;
        RECT 14.715 134.670 15.045 135.300 ;
        RECT 14.295 134.230 14.625 134.480 ;
        RECT 14.795 134.070 15.045 134.670 ;
        RECT 15.215 134.650 15.425 135.470 ;
        RECT 16.030 134.760 16.285 135.290 ;
        RECT 16.465 135.010 16.750 135.470 ;
        RECT 12.985 133.090 13.155 133.850 ;
        RECT 13.335 132.920 13.665 133.680 ;
        RECT 13.835 133.090 14.105 133.995 ;
        RECT 14.315 132.920 14.545 134.060 ;
        RECT 14.715 133.090 15.045 134.070 ;
        RECT 15.215 132.920 15.425 134.060 ;
        RECT 16.030 133.900 16.210 134.760 ;
        RECT 16.930 134.560 17.180 135.210 ;
        RECT 16.380 134.230 17.180 134.560 ;
        RECT 16.030 133.430 16.285 133.900 ;
        RECT 15.945 133.260 16.285 133.430 ;
        RECT 16.030 133.230 16.285 133.260 ;
        RECT 16.465 132.920 16.750 133.720 ;
        RECT 16.930 133.640 17.180 134.230 ;
        RECT 17.380 134.875 17.700 135.205 ;
        RECT 17.880 134.990 18.540 135.470 ;
        RECT 18.740 135.080 19.590 135.250 ;
        RECT 17.380 133.980 17.570 134.875 ;
        RECT 17.890 134.550 18.550 134.820 ;
        RECT 18.220 134.490 18.550 134.550 ;
        RECT 17.740 134.320 18.070 134.380 ;
        RECT 18.740 134.320 18.910 135.080 ;
        RECT 20.150 135.010 20.470 135.470 ;
        RECT 20.670 134.830 20.920 135.260 ;
        RECT 21.210 135.030 21.620 135.470 ;
        RECT 21.790 135.090 22.805 135.290 ;
        RECT 19.080 134.660 20.330 134.830 ;
        RECT 19.080 134.540 19.410 134.660 ;
        RECT 17.740 134.150 19.640 134.320 ;
        RECT 17.380 133.810 19.300 133.980 ;
        RECT 17.380 133.790 17.700 133.810 ;
        RECT 16.930 133.130 17.260 133.640 ;
        RECT 17.530 133.180 17.700 133.790 ;
        RECT 19.470 133.640 19.640 134.150 ;
        RECT 19.810 134.080 19.990 134.490 ;
        RECT 20.160 133.900 20.330 134.660 ;
        RECT 17.870 132.920 18.200 133.610 ;
        RECT 18.430 133.470 19.640 133.640 ;
        RECT 19.810 133.590 20.330 133.900 ;
        RECT 20.500 134.490 20.920 134.830 ;
        RECT 21.210 134.490 21.620 134.820 ;
        RECT 20.500 133.720 20.690 134.490 ;
        RECT 21.790 134.360 21.960 135.090 ;
        RECT 23.105 134.920 23.275 135.250 ;
        RECT 23.445 135.090 23.775 135.470 ;
        RECT 22.130 134.540 22.480 134.910 ;
        RECT 21.790 134.320 22.210 134.360 ;
        RECT 20.860 134.150 22.210 134.320 ;
        RECT 20.860 133.990 21.110 134.150 ;
        RECT 21.620 133.720 21.870 133.980 ;
        RECT 20.500 133.470 21.870 133.720 ;
        RECT 18.430 133.180 18.670 133.470 ;
        RECT 19.470 133.390 19.640 133.470 ;
        RECT 18.870 132.920 19.290 133.300 ;
        RECT 19.470 133.140 20.100 133.390 ;
        RECT 20.570 132.920 20.900 133.300 ;
        RECT 21.070 133.180 21.240 133.470 ;
        RECT 22.040 133.305 22.210 134.150 ;
        RECT 22.660 133.980 22.880 134.850 ;
        RECT 23.105 134.730 23.800 134.920 ;
        RECT 22.380 133.600 22.880 133.980 ;
        RECT 23.050 133.930 23.460 134.550 ;
        RECT 23.630 133.760 23.800 134.730 ;
        RECT 23.105 133.590 23.800 133.760 ;
        RECT 21.420 132.920 21.800 133.300 ;
        RECT 22.040 133.135 22.870 133.305 ;
        RECT 23.105 133.090 23.275 133.590 ;
        RECT 23.445 132.920 23.775 133.420 ;
        RECT 23.990 133.090 24.215 135.210 ;
        RECT 24.385 135.090 24.715 135.470 ;
        RECT 24.885 134.920 25.055 135.210 ;
        RECT 24.390 134.750 25.055 134.920 ;
        RECT 24.390 133.760 24.620 134.750 ;
        RECT 25.315 134.745 25.605 135.470 ;
        RECT 25.780 134.730 26.035 135.300 ;
        RECT 26.205 135.070 26.535 135.470 ;
        RECT 26.960 134.935 27.490 135.300 ;
        RECT 26.960 134.900 27.135 134.935 ;
        RECT 26.205 134.730 27.135 134.900 ;
        RECT 24.790 133.930 25.140 134.580 ;
        RECT 24.390 133.590 25.055 133.760 ;
        RECT 24.385 132.920 24.715 133.420 ;
        RECT 24.885 133.090 25.055 133.590 ;
        RECT 25.315 132.920 25.605 134.085 ;
        RECT 25.780 134.060 25.950 134.730 ;
        RECT 26.205 134.560 26.375 134.730 ;
        RECT 26.120 134.230 26.375 134.560 ;
        RECT 26.600 134.230 26.795 134.560 ;
        RECT 25.780 133.090 26.115 134.060 ;
        RECT 26.285 132.920 26.455 134.060 ;
        RECT 26.625 133.260 26.795 134.230 ;
        RECT 26.965 133.600 27.135 134.730 ;
        RECT 27.305 133.940 27.475 134.740 ;
        RECT 27.680 134.450 27.955 135.300 ;
        RECT 27.675 134.280 27.955 134.450 ;
        RECT 27.680 134.140 27.955 134.280 ;
        RECT 28.125 133.940 28.315 135.300 ;
        RECT 28.495 134.935 29.005 135.470 ;
        RECT 29.225 134.660 29.470 135.265 ;
        RECT 29.915 134.700 31.585 135.470 ;
        RECT 28.515 134.490 29.745 134.660 ;
        RECT 27.305 133.770 28.315 133.940 ;
        RECT 28.485 133.925 29.235 134.115 ;
        RECT 26.965 133.430 28.090 133.600 ;
        RECT 28.485 133.260 28.655 133.925 ;
        RECT 29.405 133.680 29.745 134.490 ;
        RECT 26.625 133.090 28.655 133.260 ;
        RECT 28.825 132.920 28.995 133.680 ;
        RECT 29.230 133.270 29.745 133.680 ;
        RECT 29.915 134.010 30.665 134.530 ;
        RECT 30.835 134.180 31.585 134.700 ;
        RECT 31.755 134.795 32.025 135.140 ;
        RECT 32.215 135.070 32.595 135.470 ;
        RECT 32.765 134.900 32.935 135.250 ;
        RECT 33.105 135.070 33.435 135.470 ;
        RECT 33.635 134.900 33.805 135.250 ;
        RECT 34.005 134.970 34.335 135.470 ;
        RECT 31.755 134.060 31.925 134.795 ;
        RECT 32.195 134.730 33.805 134.900 ;
        RECT 34.715 134.840 35.045 135.200 ;
        RECT 35.665 135.010 35.915 135.470 ;
        RECT 36.085 135.010 36.645 135.300 ;
        RECT 32.195 134.560 32.365 134.730 ;
        RECT 32.095 134.230 32.365 134.560 ;
        RECT 32.535 134.230 32.940 134.560 ;
        RECT 32.195 134.060 32.365 134.230 ;
        RECT 29.915 132.920 31.585 134.010 ;
        RECT 31.755 133.090 32.025 134.060 ;
        RECT 32.195 133.890 32.920 134.060 ;
        RECT 33.110 133.940 33.820 134.560 ;
        RECT 33.990 134.230 34.340 134.800 ;
        RECT 34.715 134.650 36.105 134.840 ;
        RECT 35.935 134.560 36.105 134.650 ;
        RECT 34.530 134.230 35.205 134.480 ;
        RECT 35.425 134.230 35.765 134.480 ;
        RECT 35.935 134.230 36.225 134.560 ;
        RECT 32.750 133.770 32.920 133.890 ;
        RECT 34.020 133.770 34.340 134.060 ;
        RECT 34.530 133.870 34.795 134.230 ;
        RECT 35.935 133.980 36.105 134.230 ;
        RECT 32.235 132.920 32.515 133.720 ;
        RECT 32.750 133.600 34.340 133.770 ;
        RECT 35.165 133.810 36.105 133.980 ;
        RECT 32.685 133.140 34.340 133.430 ;
        RECT 34.715 132.920 34.995 133.590 ;
        RECT 35.165 133.260 35.465 133.810 ;
        RECT 36.395 133.640 36.645 135.010 ;
        RECT 36.815 134.700 40.325 135.470 ;
        RECT 35.665 132.920 35.995 133.640 ;
        RECT 36.185 133.090 36.645 133.640 ;
        RECT 36.815 134.010 38.505 134.530 ;
        RECT 38.675 134.180 40.325 134.700 ;
        RECT 40.695 134.840 41.025 135.200 ;
        RECT 41.645 135.010 41.895 135.470 ;
        RECT 42.065 135.010 42.625 135.300 ;
        RECT 40.695 134.650 42.085 134.840 ;
        RECT 41.915 134.560 42.085 134.650 ;
        RECT 40.510 134.230 41.185 134.480 ;
        RECT 41.405 134.230 41.745 134.480 ;
        RECT 41.915 134.230 42.205 134.560 ;
        RECT 36.815 132.920 40.325 134.010 ;
        RECT 40.510 133.870 40.775 134.230 ;
        RECT 41.915 133.980 42.085 134.230 ;
        RECT 41.145 133.810 42.085 133.980 ;
        RECT 40.695 132.920 40.975 133.590 ;
        RECT 41.145 133.260 41.445 133.810 ;
        RECT 42.375 133.640 42.625 135.010 ;
        RECT 41.645 132.920 41.975 133.640 ;
        RECT 42.165 133.090 42.625 133.640 ;
        RECT 43.715 134.670 44.055 135.300 ;
        RECT 44.225 134.670 44.475 135.470 ;
        RECT 44.665 134.820 44.995 135.300 ;
        RECT 45.165 135.010 45.390 135.470 ;
        RECT 45.560 134.820 45.890 135.300 ;
        RECT 43.715 134.620 43.945 134.670 ;
        RECT 44.665 134.650 45.890 134.820 ;
        RECT 46.520 134.690 47.020 135.300 ;
        RECT 43.715 134.060 43.890 134.620 ;
        RECT 44.060 134.310 44.755 134.480 ;
        RECT 44.585 134.060 44.755 134.310 ;
        RECT 44.930 134.280 45.350 134.480 ;
        RECT 45.520 134.280 45.850 134.480 ;
        RECT 46.020 134.280 46.350 134.480 ;
        RECT 46.520 134.060 46.690 134.690 ;
        RECT 47.395 134.670 47.735 135.300 ;
        RECT 47.905 134.670 48.155 135.470 ;
        RECT 48.345 134.820 48.675 135.300 ;
        RECT 48.845 135.010 49.070 135.470 ;
        RECT 49.240 134.820 49.570 135.300 ;
        RECT 46.875 134.230 47.225 134.480 ;
        RECT 47.395 134.060 47.570 134.670 ;
        RECT 48.345 134.650 49.570 134.820 ;
        RECT 50.200 134.690 50.700 135.300 ;
        RECT 51.075 134.745 51.365 135.470 ;
        RECT 51.535 134.700 53.205 135.470 ;
        RECT 47.740 134.310 48.435 134.480 ;
        RECT 48.265 134.060 48.435 134.310 ;
        RECT 48.610 134.280 49.030 134.480 ;
        RECT 49.200 134.280 49.530 134.480 ;
        RECT 49.700 134.280 50.030 134.480 ;
        RECT 50.200 134.060 50.370 134.690 ;
        RECT 50.555 134.230 50.905 134.480 ;
        RECT 43.715 133.090 44.055 134.060 ;
        RECT 44.225 132.920 44.395 134.060 ;
        RECT 44.585 133.890 47.020 134.060 ;
        RECT 44.665 132.920 44.915 133.720 ;
        RECT 45.560 133.090 45.890 133.890 ;
        RECT 46.190 132.920 46.520 133.720 ;
        RECT 46.690 133.090 47.020 133.890 ;
        RECT 47.395 133.090 47.735 134.060 ;
        RECT 47.905 132.920 48.075 134.060 ;
        RECT 48.265 133.890 50.700 134.060 ;
        RECT 48.345 132.920 48.595 133.720 ;
        RECT 49.240 133.090 49.570 133.890 ;
        RECT 49.870 132.920 50.200 133.720 ;
        RECT 50.370 133.090 50.700 133.890 ;
        RECT 51.075 132.920 51.365 134.085 ;
        RECT 51.535 134.010 52.285 134.530 ;
        RECT 52.455 134.180 53.205 134.700 ;
        RECT 53.490 134.840 53.775 135.300 ;
        RECT 53.945 135.010 54.215 135.470 ;
        RECT 53.490 134.670 54.445 134.840 ;
        RECT 51.535 132.920 53.205 134.010 ;
        RECT 53.375 133.940 54.065 134.500 ;
        RECT 54.235 133.770 54.445 134.670 ;
        RECT 53.490 133.550 54.445 133.770 ;
        RECT 54.615 134.500 55.015 135.300 ;
        RECT 55.205 134.840 55.485 135.300 ;
        RECT 56.005 135.010 56.330 135.470 ;
        RECT 55.205 134.670 56.330 134.840 ;
        RECT 56.500 134.730 56.885 135.300 ;
        RECT 57.430 134.790 57.685 135.290 ;
        RECT 57.865 135.010 58.150 135.470 ;
        RECT 55.880 134.560 56.330 134.670 ;
        RECT 54.615 133.940 55.710 134.500 ;
        RECT 55.880 134.230 56.435 134.560 ;
        RECT 53.490 133.090 53.775 133.550 ;
        RECT 53.945 132.920 54.215 133.380 ;
        RECT 54.615 133.090 55.015 133.940 ;
        RECT 55.880 133.770 56.330 134.230 ;
        RECT 56.605 134.060 56.885 134.730 ;
        RECT 57.345 134.760 57.685 134.790 ;
        RECT 57.345 134.620 57.610 134.760 ;
        RECT 55.205 133.550 56.330 133.770 ;
        RECT 55.205 133.090 55.485 133.550 ;
        RECT 56.005 132.920 56.330 133.380 ;
        RECT 56.500 133.090 56.885 134.060 ;
        RECT 57.430 133.900 57.610 134.620 ;
        RECT 58.330 134.560 58.580 135.210 ;
        RECT 57.780 134.230 58.580 134.560 ;
        RECT 57.430 133.230 57.685 133.900 ;
        RECT 57.865 132.920 58.150 133.720 ;
        RECT 58.330 133.640 58.580 134.230 ;
        RECT 58.780 134.875 59.100 135.205 ;
        RECT 59.280 134.990 59.940 135.470 ;
        RECT 60.140 135.080 60.990 135.250 ;
        RECT 58.780 133.980 58.970 134.875 ;
        RECT 59.290 134.550 59.950 134.820 ;
        RECT 59.620 134.490 59.950 134.550 ;
        RECT 59.140 134.320 59.470 134.380 ;
        RECT 60.140 134.320 60.310 135.080 ;
        RECT 61.550 135.010 61.870 135.470 ;
        RECT 62.070 134.830 62.320 135.260 ;
        RECT 62.610 135.030 63.020 135.470 ;
        RECT 63.190 135.090 64.205 135.290 ;
        RECT 60.480 134.660 61.730 134.830 ;
        RECT 60.480 134.540 60.810 134.660 ;
        RECT 59.140 134.150 61.040 134.320 ;
        RECT 58.780 133.810 60.700 133.980 ;
        RECT 58.780 133.790 59.100 133.810 ;
        RECT 58.330 133.130 58.660 133.640 ;
        RECT 58.930 133.180 59.100 133.790 ;
        RECT 60.870 133.640 61.040 134.150 ;
        RECT 61.210 134.080 61.390 134.490 ;
        RECT 61.560 133.900 61.730 134.660 ;
        RECT 59.270 132.920 59.600 133.610 ;
        RECT 59.830 133.470 61.040 133.640 ;
        RECT 61.210 133.590 61.730 133.900 ;
        RECT 61.900 134.490 62.320 134.830 ;
        RECT 62.610 134.490 63.020 134.820 ;
        RECT 61.900 133.720 62.090 134.490 ;
        RECT 63.190 134.360 63.360 135.090 ;
        RECT 64.505 134.920 64.675 135.250 ;
        RECT 64.845 135.090 65.175 135.470 ;
        RECT 63.530 134.540 63.880 134.910 ;
        RECT 63.190 134.320 63.610 134.360 ;
        RECT 62.260 134.150 63.610 134.320 ;
        RECT 62.260 133.990 62.510 134.150 ;
        RECT 63.020 133.720 63.270 133.980 ;
        RECT 61.900 133.470 63.270 133.720 ;
        RECT 59.830 133.180 60.070 133.470 ;
        RECT 60.870 133.390 61.040 133.470 ;
        RECT 60.270 132.920 60.690 133.300 ;
        RECT 60.870 133.140 61.500 133.390 ;
        RECT 61.970 132.920 62.300 133.300 ;
        RECT 62.470 133.180 62.640 133.470 ;
        RECT 63.440 133.305 63.610 134.150 ;
        RECT 64.060 133.980 64.280 134.850 ;
        RECT 64.505 134.730 65.200 134.920 ;
        RECT 63.780 133.600 64.280 133.980 ;
        RECT 64.450 133.930 64.860 134.550 ;
        RECT 65.030 133.760 65.200 134.730 ;
        RECT 64.505 133.590 65.200 133.760 ;
        RECT 62.820 132.920 63.200 133.300 ;
        RECT 63.440 133.135 64.270 133.305 ;
        RECT 64.505 133.090 64.675 133.590 ;
        RECT 64.845 132.920 65.175 133.420 ;
        RECT 65.390 133.090 65.615 135.210 ;
        RECT 65.785 135.090 66.115 135.470 ;
        RECT 66.285 134.920 66.455 135.210 ;
        RECT 65.790 134.750 66.455 134.920 ;
        RECT 65.790 133.760 66.020 134.750 ;
        RECT 66.715 134.720 67.925 135.470 ;
        RECT 66.190 133.930 66.540 134.580 ;
        RECT 66.715 134.010 67.235 134.550 ;
        RECT 67.405 134.180 67.925 134.720 ;
        RECT 68.295 134.840 68.625 135.200 ;
        RECT 69.245 135.010 69.495 135.470 ;
        RECT 69.665 135.010 70.225 135.300 ;
        RECT 68.295 134.650 69.685 134.840 ;
        RECT 69.515 134.560 69.685 134.650 ;
        RECT 68.110 134.230 68.785 134.480 ;
        RECT 69.005 134.230 69.345 134.480 ;
        RECT 69.515 134.230 69.805 134.560 ;
        RECT 65.790 133.590 66.455 133.760 ;
        RECT 65.785 132.920 66.115 133.420 ;
        RECT 66.285 133.090 66.455 133.590 ;
        RECT 66.715 132.920 67.925 134.010 ;
        RECT 68.110 133.870 68.375 134.230 ;
        RECT 69.515 133.980 69.685 134.230 ;
        RECT 68.745 133.810 69.685 133.980 ;
        RECT 68.295 132.920 68.575 133.590 ;
        RECT 68.745 133.260 69.045 133.810 ;
        RECT 69.975 133.640 70.225 135.010 ;
        RECT 69.245 132.920 69.575 133.640 ;
        RECT 69.765 133.090 70.225 133.640 ;
        RECT 70.395 135.010 70.955 135.300 ;
        RECT 71.125 135.010 71.375 135.470 ;
        RECT 70.395 133.640 70.645 135.010 ;
        RECT 71.995 134.840 72.325 135.200 ;
        RECT 70.935 134.650 72.325 134.840 ;
        RECT 73.155 134.700 76.665 135.470 ;
        RECT 76.835 134.745 77.125 135.470 ;
        RECT 77.295 134.720 78.505 135.470 ;
        RECT 70.935 134.560 71.105 134.650 ;
        RECT 70.815 134.230 71.105 134.560 ;
        RECT 71.275 134.230 71.615 134.480 ;
        RECT 71.835 134.230 72.510 134.480 ;
        RECT 70.935 133.980 71.105 134.230 ;
        RECT 70.935 133.810 71.875 133.980 ;
        RECT 72.245 133.870 72.510 134.230 ;
        RECT 73.155 134.010 74.845 134.530 ;
        RECT 75.015 134.180 76.665 134.700 ;
        RECT 70.395 133.090 70.855 133.640 ;
        RECT 71.045 132.920 71.375 133.640 ;
        RECT 71.575 133.260 71.875 133.810 ;
        RECT 72.045 132.920 72.325 133.590 ;
        RECT 73.155 132.920 76.665 134.010 ;
        RECT 76.835 132.920 77.125 134.085 ;
        RECT 77.295 134.010 77.815 134.550 ;
        RECT 77.985 134.180 78.505 134.720 ;
        RECT 78.675 134.700 82.185 135.470 ;
        RECT 78.675 134.010 80.365 134.530 ;
        RECT 80.535 134.180 82.185 134.700 ;
        RECT 82.415 134.650 82.625 135.470 ;
        RECT 82.795 134.670 83.125 135.300 ;
        RECT 82.795 134.070 83.045 134.670 ;
        RECT 83.295 134.650 83.525 135.470 ;
        RECT 83.735 134.700 87.245 135.470 ;
        RECT 87.425 134.970 87.755 135.470 ;
        RECT 87.955 134.900 88.125 135.250 ;
        RECT 88.325 135.070 88.655 135.470 ;
        RECT 88.825 134.900 88.995 135.250 ;
        RECT 89.165 135.070 89.545 135.470 ;
        RECT 83.215 134.230 83.545 134.480 ;
        RECT 77.295 132.920 78.505 134.010 ;
        RECT 78.675 132.920 82.185 134.010 ;
        RECT 82.415 132.920 82.625 134.060 ;
        RECT 82.795 133.090 83.125 134.070 ;
        RECT 83.295 132.920 83.525 134.060 ;
        RECT 83.735 134.010 85.425 134.530 ;
        RECT 85.595 134.180 87.245 134.700 ;
        RECT 87.420 134.230 87.770 134.800 ;
        RECT 87.955 134.730 89.565 134.900 ;
        RECT 89.735 134.795 90.005 135.140 ;
        RECT 89.395 134.560 89.565 134.730 ;
        RECT 83.735 132.920 87.245 134.010 ;
        RECT 87.420 133.770 87.740 134.060 ;
        RECT 87.940 133.940 88.650 134.560 ;
        RECT 88.820 134.230 89.225 134.560 ;
        RECT 89.395 134.230 89.665 134.560 ;
        RECT 89.395 134.060 89.565 134.230 ;
        RECT 89.835 134.060 90.005 134.795 ;
        RECT 91.135 134.650 91.365 135.470 ;
        RECT 91.535 134.670 91.865 135.300 ;
        RECT 91.115 134.230 91.445 134.480 ;
        RECT 91.615 134.070 91.865 134.670 ;
        RECT 92.035 134.650 92.245 135.470 ;
        RECT 92.945 134.970 93.275 135.470 ;
        RECT 93.475 134.900 93.645 135.250 ;
        RECT 93.845 135.070 94.175 135.470 ;
        RECT 94.345 134.900 94.515 135.250 ;
        RECT 94.685 135.070 95.065 135.470 ;
        RECT 92.940 134.230 93.290 134.800 ;
        RECT 93.475 134.730 95.085 134.900 ;
        RECT 95.255 134.795 95.525 135.140 ;
        RECT 94.915 134.560 95.085 134.730 ;
        RECT 88.840 133.890 89.565 134.060 ;
        RECT 88.840 133.770 89.010 133.890 ;
        RECT 87.420 133.600 89.010 133.770 ;
        RECT 87.420 133.140 89.075 133.430 ;
        RECT 89.245 132.920 89.525 133.720 ;
        RECT 89.735 133.090 90.005 134.060 ;
        RECT 91.135 132.920 91.365 134.060 ;
        RECT 91.535 133.090 91.865 134.070 ;
        RECT 92.035 132.920 92.245 134.060 ;
        RECT 92.940 133.770 93.260 134.060 ;
        RECT 93.460 133.940 94.170 134.560 ;
        RECT 94.340 134.230 94.745 134.560 ;
        RECT 94.915 134.230 95.185 134.560 ;
        RECT 94.915 134.060 95.085 134.230 ;
        RECT 95.355 134.060 95.525 134.795 ;
        RECT 94.360 133.890 95.085 134.060 ;
        RECT 94.360 133.770 94.530 133.890 ;
        RECT 92.940 133.600 94.530 133.770 ;
        RECT 92.940 133.140 94.595 133.430 ;
        RECT 94.765 132.920 95.045 133.720 ;
        RECT 95.255 133.090 95.525 134.060 ;
        RECT 95.695 134.670 96.035 135.300 ;
        RECT 96.205 134.670 96.455 135.470 ;
        RECT 96.645 134.820 96.975 135.300 ;
        RECT 97.145 135.010 97.370 135.470 ;
        RECT 97.540 134.820 97.870 135.300 ;
        RECT 95.695 134.620 95.925 134.670 ;
        RECT 96.645 134.650 97.870 134.820 ;
        RECT 98.500 134.690 99.000 135.300 ;
        RECT 99.375 134.795 99.645 135.140 ;
        RECT 99.835 135.070 100.215 135.470 ;
        RECT 100.385 134.900 100.555 135.250 ;
        RECT 100.725 135.070 101.055 135.470 ;
        RECT 101.255 134.900 101.425 135.250 ;
        RECT 101.625 134.970 101.955 135.470 ;
        RECT 95.695 134.060 95.870 134.620 ;
        RECT 96.040 134.310 96.735 134.480 ;
        RECT 96.565 134.060 96.735 134.310 ;
        RECT 96.910 134.280 97.330 134.480 ;
        RECT 97.500 134.280 97.830 134.480 ;
        RECT 98.000 134.280 98.330 134.480 ;
        RECT 98.500 134.060 98.670 134.690 ;
        RECT 98.855 134.230 99.205 134.480 ;
        RECT 99.375 134.060 99.545 134.795 ;
        RECT 99.815 134.730 101.425 134.900 ;
        RECT 99.815 134.560 99.985 134.730 ;
        RECT 99.715 134.230 99.985 134.560 ;
        RECT 100.155 134.230 100.560 134.560 ;
        RECT 99.815 134.060 99.985 134.230 ;
        RECT 100.730 134.110 101.440 134.560 ;
        RECT 101.610 134.230 101.960 134.800 ;
        RECT 102.595 134.745 102.885 135.470 ;
        RECT 103.330 134.660 103.575 135.265 ;
        RECT 103.795 134.935 104.305 135.470 ;
        RECT 103.055 134.490 104.285 134.660 ;
        RECT 95.695 133.090 96.035 134.060 ;
        RECT 96.205 132.920 96.375 134.060 ;
        RECT 96.565 133.890 99.000 134.060 ;
        RECT 96.645 132.920 96.895 133.720 ;
        RECT 97.540 133.090 97.870 133.890 ;
        RECT 98.170 132.920 98.500 133.720 ;
        RECT 98.670 133.090 99.000 133.890 ;
        RECT 99.375 133.090 99.645 134.060 ;
        RECT 99.815 133.890 100.540 134.060 ;
        RECT 100.730 133.940 101.445 134.110 ;
        RECT 100.370 133.770 100.540 133.890 ;
        RECT 101.640 133.770 101.960 134.060 ;
        RECT 99.855 132.920 100.135 133.720 ;
        RECT 100.370 133.600 101.960 133.770 ;
        RECT 100.305 133.140 101.960 133.430 ;
        RECT 102.595 132.920 102.885 134.085 ;
        RECT 103.055 133.680 103.395 134.490 ;
        RECT 103.565 133.925 104.315 134.115 ;
        RECT 103.055 133.270 103.570 133.680 ;
        RECT 103.805 132.920 103.975 133.680 ;
        RECT 104.145 133.260 104.315 133.925 ;
        RECT 104.485 133.940 104.675 135.300 ;
        RECT 104.845 135.130 105.120 135.300 ;
        RECT 104.845 134.960 105.125 135.130 ;
        RECT 104.845 134.140 105.120 134.960 ;
        RECT 105.310 134.935 105.840 135.300 ;
        RECT 106.265 135.070 106.595 135.470 ;
        RECT 105.665 134.900 105.840 134.935 ;
        RECT 105.325 133.940 105.495 134.740 ;
        RECT 104.485 133.770 105.495 133.940 ;
        RECT 105.665 134.730 106.595 134.900 ;
        RECT 106.765 134.730 107.020 135.300 ;
        RECT 107.745 134.920 107.915 135.300 ;
        RECT 108.095 135.090 108.425 135.470 ;
        RECT 107.745 134.750 108.410 134.920 ;
        RECT 108.605 134.795 108.865 135.300 ;
        RECT 109.040 134.925 114.385 135.470 ;
        RECT 105.665 133.600 105.835 134.730 ;
        RECT 106.425 134.560 106.595 134.730 ;
        RECT 104.710 133.430 105.835 133.600 ;
        RECT 106.005 134.230 106.200 134.560 ;
        RECT 106.425 134.230 106.680 134.560 ;
        RECT 106.005 133.260 106.175 134.230 ;
        RECT 106.850 134.060 107.020 134.730 ;
        RECT 107.675 134.200 108.005 134.570 ;
        RECT 108.240 134.495 108.410 134.750 ;
        RECT 104.145 133.090 106.175 133.260 ;
        RECT 106.345 132.920 106.515 134.060 ;
        RECT 106.685 133.090 107.020 134.060 ;
        RECT 108.240 134.165 108.525 134.495 ;
        RECT 108.240 134.020 108.410 134.165 ;
        RECT 107.745 133.850 108.410 134.020 ;
        RECT 108.695 133.995 108.865 134.795 ;
        RECT 107.745 133.090 107.915 133.850 ;
        RECT 108.095 132.920 108.425 133.680 ;
        RECT 108.595 133.090 108.865 133.995 ;
        RECT 110.630 133.355 110.980 134.605 ;
        RECT 112.460 134.095 112.800 134.925 ;
        RECT 114.555 134.720 115.765 135.470 ;
        RECT 114.555 134.010 115.075 134.550 ;
        RECT 115.245 134.180 115.765 134.720 ;
        RECT 109.040 132.920 114.385 133.355 ;
        RECT 114.555 132.920 115.765 134.010 ;
        RECT 10.510 132.750 115.850 132.920 ;
        RECT 10.595 131.660 11.805 132.750 ;
        RECT 10.595 130.950 11.115 131.490 ;
        RECT 11.285 131.120 11.805 131.660 ;
        RECT 12.435 131.585 12.725 132.750 ;
        RECT 12.895 131.990 13.410 132.400 ;
        RECT 13.645 131.990 13.815 132.750 ;
        RECT 13.985 132.410 16.015 132.580 ;
        RECT 12.895 131.180 13.235 131.990 ;
        RECT 13.985 131.745 14.155 132.410 ;
        RECT 14.550 132.070 15.675 132.240 ;
        RECT 13.405 131.555 14.155 131.745 ;
        RECT 14.325 131.730 15.335 131.900 ;
        RECT 12.895 131.010 14.125 131.180 ;
        RECT 10.595 130.200 11.805 130.950 ;
        RECT 12.435 130.200 12.725 130.925 ;
        RECT 13.170 130.405 13.415 131.010 ;
        RECT 13.635 130.200 14.145 130.735 ;
        RECT 14.325 130.370 14.515 131.730 ;
        RECT 14.685 131.050 14.960 131.530 ;
        RECT 14.685 130.880 14.965 131.050 ;
        RECT 15.165 130.930 15.335 131.730 ;
        RECT 15.505 130.940 15.675 132.070 ;
        RECT 15.845 131.440 16.015 132.410 ;
        RECT 16.185 131.610 16.355 132.750 ;
        RECT 16.525 131.610 16.860 132.580 ;
        RECT 15.845 131.110 16.040 131.440 ;
        RECT 16.265 131.110 16.520 131.440 ;
        RECT 16.265 130.940 16.435 131.110 ;
        RECT 16.690 130.940 16.860 131.610 ;
        RECT 14.685 130.370 14.960 130.880 ;
        RECT 15.505 130.770 16.435 130.940 ;
        RECT 15.505 130.735 15.680 130.770 ;
        RECT 15.150 130.370 15.680 130.735 ;
        RECT 16.105 130.200 16.435 130.600 ;
        RECT 16.605 130.370 16.860 130.940 ;
        RECT 17.040 131.610 17.375 132.580 ;
        RECT 17.545 131.610 17.715 132.750 ;
        RECT 17.885 132.410 19.915 132.580 ;
        RECT 17.040 130.940 17.210 131.610 ;
        RECT 17.885 131.440 18.055 132.410 ;
        RECT 17.380 131.110 17.635 131.440 ;
        RECT 17.860 131.110 18.055 131.440 ;
        RECT 18.225 132.070 19.350 132.240 ;
        RECT 17.465 130.940 17.635 131.110 ;
        RECT 18.225 130.940 18.395 132.070 ;
        RECT 17.040 130.370 17.295 130.940 ;
        RECT 17.465 130.770 18.395 130.940 ;
        RECT 18.565 131.730 19.575 131.900 ;
        RECT 18.565 130.930 18.735 131.730 ;
        RECT 18.220 130.735 18.395 130.770 ;
        RECT 17.465 130.200 17.795 130.600 ;
        RECT 18.220 130.370 18.750 130.735 ;
        RECT 18.940 130.710 19.215 131.530 ;
        RECT 18.935 130.540 19.215 130.710 ;
        RECT 18.940 130.370 19.215 130.540 ;
        RECT 19.385 130.370 19.575 131.730 ;
        RECT 19.745 131.745 19.915 132.410 ;
        RECT 20.085 131.990 20.255 132.750 ;
        RECT 20.490 131.990 21.005 132.400 ;
        RECT 21.180 132.315 26.525 132.750 ;
        RECT 19.745 131.555 20.495 131.745 ;
        RECT 20.665 131.180 21.005 131.990 ;
        RECT 19.775 131.010 21.005 131.180 ;
        RECT 22.770 131.065 23.120 132.315 ;
        RECT 26.895 132.080 27.175 132.750 ;
        RECT 27.345 131.860 27.645 132.410 ;
        RECT 27.845 132.030 28.175 132.750 ;
        RECT 28.365 132.030 28.825 132.580 ;
        RECT 19.755 130.200 20.265 130.735 ;
        RECT 20.485 130.405 20.730 131.010 ;
        RECT 24.600 130.745 24.940 131.575 ;
        RECT 26.710 131.440 26.975 131.800 ;
        RECT 27.345 131.690 28.285 131.860 ;
        RECT 28.115 131.440 28.285 131.690 ;
        RECT 26.710 131.190 27.385 131.440 ;
        RECT 27.605 131.190 27.945 131.440 ;
        RECT 28.115 131.110 28.405 131.440 ;
        RECT 28.115 131.020 28.285 131.110 ;
        RECT 26.895 130.830 28.285 131.020 ;
        RECT 21.180 130.200 26.525 130.745 ;
        RECT 26.895 130.470 27.225 130.830 ;
        RECT 28.575 130.660 28.825 132.030 ;
        RECT 27.845 130.200 28.095 130.660 ;
        RECT 28.265 130.370 28.825 130.660 ;
        RECT 29.000 131.610 29.335 132.580 ;
        RECT 29.505 131.610 29.675 132.750 ;
        RECT 29.845 132.410 31.875 132.580 ;
        RECT 29.000 130.940 29.170 131.610 ;
        RECT 29.845 131.440 30.015 132.410 ;
        RECT 29.340 131.110 29.595 131.440 ;
        RECT 29.820 131.110 30.015 131.440 ;
        RECT 30.185 132.070 31.310 132.240 ;
        RECT 29.425 130.940 29.595 131.110 ;
        RECT 30.185 130.940 30.355 132.070 ;
        RECT 29.000 130.370 29.255 130.940 ;
        RECT 29.425 130.770 30.355 130.940 ;
        RECT 30.525 131.730 31.535 131.900 ;
        RECT 30.525 130.930 30.695 131.730 ;
        RECT 30.180 130.735 30.355 130.770 ;
        RECT 29.425 130.200 29.755 130.600 ;
        RECT 30.180 130.370 30.710 130.735 ;
        RECT 30.900 130.710 31.175 131.530 ;
        RECT 30.895 130.540 31.175 130.710 ;
        RECT 30.900 130.370 31.175 130.540 ;
        RECT 31.345 130.370 31.535 131.730 ;
        RECT 31.705 131.745 31.875 132.410 ;
        RECT 32.045 131.990 32.215 132.750 ;
        RECT 32.450 131.990 32.965 132.400 ;
        RECT 31.705 131.555 32.455 131.745 ;
        RECT 32.625 131.180 32.965 131.990 ;
        RECT 31.735 131.010 32.965 131.180 ;
        RECT 33.135 131.660 34.345 132.750 ;
        RECT 34.515 131.660 38.025 132.750 ;
        RECT 33.135 131.120 33.655 131.660 ;
        RECT 31.715 130.200 32.225 130.735 ;
        RECT 32.445 130.405 32.690 131.010 ;
        RECT 33.825 130.950 34.345 131.490 ;
        RECT 34.515 131.140 36.205 131.660 ;
        RECT 38.195 131.585 38.485 132.750 ;
        RECT 39.115 131.660 40.785 132.750 ;
        RECT 41.155 132.080 41.435 132.750 ;
        RECT 41.605 131.860 41.905 132.410 ;
        RECT 42.105 132.030 42.435 132.750 ;
        RECT 42.625 132.030 43.085 132.580 ;
        RECT 36.375 130.970 38.025 131.490 ;
        RECT 39.115 131.140 39.865 131.660 ;
        RECT 40.035 130.970 40.785 131.490 ;
        RECT 40.970 131.440 41.235 131.800 ;
        RECT 41.605 131.690 42.545 131.860 ;
        RECT 42.375 131.440 42.545 131.690 ;
        RECT 40.970 131.190 41.645 131.440 ;
        RECT 41.865 131.190 42.205 131.440 ;
        RECT 42.375 131.110 42.665 131.440 ;
        RECT 42.375 131.020 42.545 131.110 ;
        RECT 33.135 130.200 34.345 130.950 ;
        RECT 34.515 130.200 38.025 130.970 ;
        RECT 38.195 130.200 38.485 130.925 ;
        RECT 39.115 130.200 40.785 130.970 ;
        RECT 41.155 130.830 42.545 131.020 ;
        RECT 41.155 130.470 41.485 130.830 ;
        RECT 42.835 130.660 43.085 132.030 ;
        RECT 43.345 132.080 43.515 132.580 ;
        RECT 43.685 132.250 44.015 132.750 ;
        RECT 43.345 131.910 44.010 132.080 ;
        RECT 43.260 131.090 43.610 131.740 ;
        RECT 43.780 130.920 44.010 131.910 ;
        RECT 42.105 130.200 42.355 130.660 ;
        RECT 42.525 130.370 43.085 130.660 ;
        RECT 43.345 130.750 44.010 130.920 ;
        RECT 43.345 130.460 43.515 130.750 ;
        RECT 43.685 130.200 44.015 130.580 ;
        RECT 44.185 130.460 44.410 132.580 ;
        RECT 44.625 132.250 44.955 132.750 ;
        RECT 45.125 132.080 45.295 132.580 ;
        RECT 45.530 132.365 46.360 132.535 ;
        RECT 46.600 132.370 46.980 132.750 ;
        RECT 44.600 131.910 45.295 132.080 ;
        RECT 44.600 130.940 44.770 131.910 ;
        RECT 44.940 131.120 45.350 131.740 ;
        RECT 45.520 131.690 46.020 132.070 ;
        RECT 44.600 130.750 45.295 130.940 ;
        RECT 45.520 130.820 45.740 131.690 ;
        RECT 46.190 131.520 46.360 132.365 ;
        RECT 47.160 132.200 47.330 132.490 ;
        RECT 47.500 132.370 47.830 132.750 ;
        RECT 48.300 132.280 48.930 132.530 ;
        RECT 49.110 132.370 49.530 132.750 ;
        RECT 48.760 132.200 48.930 132.280 ;
        RECT 49.730 132.200 49.970 132.490 ;
        RECT 46.530 131.950 47.900 132.200 ;
        RECT 46.530 131.690 46.780 131.950 ;
        RECT 47.290 131.520 47.540 131.680 ;
        RECT 46.190 131.350 47.540 131.520 ;
        RECT 46.190 131.310 46.610 131.350 ;
        RECT 45.920 130.760 46.270 131.130 ;
        RECT 44.625 130.200 44.955 130.580 ;
        RECT 45.125 130.420 45.295 130.750 ;
        RECT 46.440 130.580 46.610 131.310 ;
        RECT 47.710 131.180 47.900 131.950 ;
        RECT 46.780 130.850 47.190 131.180 ;
        RECT 47.480 130.840 47.900 131.180 ;
        RECT 48.070 131.770 48.590 132.080 ;
        RECT 48.760 132.030 49.970 132.200 ;
        RECT 50.200 132.060 50.530 132.750 ;
        RECT 48.070 131.010 48.240 131.770 ;
        RECT 48.410 131.180 48.590 131.590 ;
        RECT 48.760 131.520 48.930 132.030 ;
        RECT 50.700 131.880 50.870 132.490 ;
        RECT 51.140 132.030 51.470 132.540 ;
        RECT 50.700 131.860 51.020 131.880 ;
        RECT 49.100 131.690 51.020 131.860 ;
        RECT 48.760 131.350 50.660 131.520 ;
        RECT 48.990 131.010 49.320 131.130 ;
        RECT 48.070 130.840 49.320 131.010 ;
        RECT 45.595 130.380 46.610 130.580 ;
        RECT 46.780 130.200 47.190 130.640 ;
        RECT 47.480 130.410 47.730 130.840 ;
        RECT 47.930 130.200 48.250 130.660 ;
        RECT 49.490 130.590 49.660 131.350 ;
        RECT 50.330 131.290 50.660 131.350 ;
        RECT 49.850 131.120 50.180 131.180 ;
        RECT 49.850 130.850 50.510 131.120 ;
        RECT 50.830 130.795 51.020 131.690 ;
        RECT 48.810 130.420 49.660 130.590 ;
        RECT 49.860 130.200 50.520 130.680 ;
        RECT 50.700 130.465 51.020 130.795 ;
        RECT 51.220 131.440 51.470 132.030 ;
        RECT 51.650 131.950 51.935 132.750 ;
        RECT 52.115 132.410 52.370 132.440 ;
        RECT 52.115 132.240 52.455 132.410 ;
        RECT 52.115 131.770 52.370 132.240 ;
        RECT 51.220 131.110 52.020 131.440 ;
        RECT 51.220 130.460 51.470 131.110 ;
        RECT 52.190 130.910 52.370 131.770 ;
        RECT 52.915 131.660 54.125 132.750 ;
        RECT 54.300 132.315 59.645 132.750 ;
        RECT 59.820 132.325 60.155 132.750 ;
        RECT 52.915 131.120 53.435 131.660 ;
        RECT 53.605 130.950 54.125 131.490 ;
        RECT 55.890 131.065 56.240 132.315 ;
        RECT 60.325 132.145 60.510 132.550 ;
        RECT 59.845 131.970 60.510 132.145 ;
        RECT 60.715 131.970 61.045 132.750 ;
        RECT 51.650 130.200 51.935 130.660 ;
        RECT 52.115 130.380 52.370 130.910 ;
        RECT 52.915 130.200 54.125 130.950 ;
        RECT 57.720 130.745 58.060 131.575 ;
        RECT 59.845 130.940 60.185 131.970 ;
        RECT 61.215 131.780 61.485 132.550 ;
        RECT 61.855 132.080 62.135 132.750 ;
        RECT 62.305 131.860 62.605 132.410 ;
        RECT 62.805 132.030 63.135 132.750 ;
        RECT 63.325 132.030 63.785 132.580 ;
        RECT 60.355 131.610 61.485 131.780 ;
        RECT 60.355 131.110 60.605 131.610 ;
        RECT 59.845 130.770 60.530 130.940 ;
        RECT 60.785 130.860 61.145 131.440 ;
        RECT 54.300 130.200 59.645 130.745 ;
        RECT 59.820 130.200 60.155 130.600 ;
        RECT 60.325 130.370 60.530 130.770 ;
        RECT 61.315 130.700 61.485 131.610 ;
        RECT 61.670 131.440 61.935 131.800 ;
        RECT 62.305 131.690 63.245 131.860 ;
        RECT 63.075 131.440 63.245 131.690 ;
        RECT 61.670 131.190 62.345 131.440 ;
        RECT 62.565 131.190 62.905 131.440 ;
        RECT 63.075 131.110 63.365 131.440 ;
        RECT 63.075 131.020 63.245 131.110 ;
        RECT 60.740 130.200 61.015 130.680 ;
        RECT 61.225 130.370 61.485 130.700 ;
        RECT 61.855 130.830 63.245 131.020 ;
        RECT 61.855 130.470 62.185 130.830 ;
        RECT 63.535 130.660 63.785 132.030 ;
        RECT 63.955 131.585 64.245 132.750 ;
        RECT 64.415 131.780 64.685 132.550 ;
        RECT 64.855 131.970 65.185 132.750 ;
        RECT 65.390 132.145 65.575 132.550 ;
        RECT 65.745 132.325 66.080 132.750 ;
        RECT 65.390 131.970 66.055 132.145 ;
        RECT 64.415 131.610 65.545 131.780 ;
        RECT 62.805 130.200 63.055 130.660 ;
        RECT 63.225 130.370 63.785 130.660 ;
        RECT 63.955 130.200 64.245 130.925 ;
        RECT 64.415 130.700 64.585 131.610 ;
        RECT 64.755 130.860 65.115 131.440 ;
        RECT 65.295 131.110 65.545 131.610 ;
        RECT 65.715 130.940 66.055 131.970 ;
        RECT 65.370 130.770 66.055 130.940 ;
        RECT 66.255 132.030 66.715 132.580 ;
        RECT 66.905 132.030 67.235 132.750 ;
        RECT 64.415 130.370 64.675 130.700 ;
        RECT 64.885 130.200 65.160 130.680 ;
        RECT 65.370 130.370 65.575 130.770 ;
        RECT 66.255 130.660 66.505 132.030 ;
        RECT 67.435 131.860 67.735 132.410 ;
        RECT 67.905 132.080 68.185 132.750 ;
        RECT 66.795 131.690 67.735 131.860 ;
        RECT 68.555 132.030 69.015 132.580 ;
        RECT 69.205 132.030 69.535 132.750 ;
        RECT 66.795 131.440 66.965 131.690 ;
        RECT 68.105 131.440 68.370 131.800 ;
        RECT 66.675 131.110 66.965 131.440 ;
        RECT 67.135 131.190 67.475 131.440 ;
        RECT 67.695 131.190 68.370 131.440 ;
        RECT 66.795 131.020 66.965 131.110 ;
        RECT 66.795 130.830 68.185 131.020 ;
        RECT 65.745 130.200 66.080 130.600 ;
        RECT 66.255 130.370 66.815 130.660 ;
        RECT 66.985 130.200 67.235 130.660 ;
        RECT 67.855 130.470 68.185 130.830 ;
        RECT 68.555 130.660 68.805 132.030 ;
        RECT 69.735 131.860 70.035 132.410 ;
        RECT 70.205 132.080 70.485 132.750 ;
        RECT 69.095 131.690 70.035 131.860 ;
        RECT 71.775 131.990 72.290 132.400 ;
        RECT 72.525 131.990 72.695 132.750 ;
        RECT 72.865 132.410 74.895 132.580 ;
        RECT 69.095 131.440 69.265 131.690 ;
        RECT 70.405 131.440 70.670 131.800 ;
        RECT 68.975 131.110 69.265 131.440 ;
        RECT 69.435 131.190 69.775 131.440 ;
        RECT 69.995 131.190 70.670 131.440 ;
        RECT 69.095 131.020 69.265 131.110 ;
        RECT 71.775 131.180 72.115 131.990 ;
        RECT 72.865 131.745 73.035 132.410 ;
        RECT 73.430 132.070 74.555 132.240 ;
        RECT 72.285 131.555 73.035 131.745 ;
        RECT 73.205 131.730 74.215 131.900 ;
        RECT 69.095 130.830 70.485 131.020 ;
        RECT 71.775 131.010 73.005 131.180 ;
        RECT 68.555 130.370 69.115 130.660 ;
        RECT 69.285 130.200 69.535 130.660 ;
        RECT 70.155 130.470 70.485 130.830 ;
        RECT 72.050 130.405 72.295 131.010 ;
        RECT 72.515 130.200 73.025 130.735 ;
        RECT 73.205 130.370 73.395 131.730 ;
        RECT 73.565 131.050 73.840 131.530 ;
        RECT 73.565 130.880 73.845 131.050 ;
        RECT 74.045 130.930 74.215 131.730 ;
        RECT 74.385 130.940 74.555 132.070 ;
        RECT 74.725 131.440 74.895 132.410 ;
        RECT 75.065 131.610 75.235 132.750 ;
        RECT 75.405 131.610 75.740 132.580 ;
        RECT 74.725 131.110 74.920 131.440 ;
        RECT 75.145 131.110 75.400 131.440 ;
        RECT 75.145 130.940 75.315 131.110 ;
        RECT 75.570 130.940 75.740 131.610 ;
        RECT 75.915 131.660 78.505 132.750 ;
        RECT 78.680 132.315 84.025 132.750 ;
        RECT 84.200 132.315 89.545 132.750 ;
        RECT 75.915 131.140 77.125 131.660 ;
        RECT 77.295 130.970 78.505 131.490 ;
        RECT 80.270 131.065 80.620 132.315 ;
        RECT 73.565 130.370 73.840 130.880 ;
        RECT 74.385 130.770 75.315 130.940 ;
        RECT 74.385 130.735 74.560 130.770 ;
        RECT 74.030 130.370 74.560 130.735 ;
        RECT 74.985 130.200 75.315 130.600 ;
        RECT 75.485 130.370 75.740 130.940 ;
        RECT 75.915 130.200 78.505 130.970 ;
        RECT 82.100 130.745 82.440 131.575 ;
        RECT 85.790 131.065 86.140 132.315 ;
        RECT 89.715 131.585 90.005 132.750 ;
        RECT 90.175 131.660 91.385 132.750 ;
        RECT 91.560 132.315 96.905 132.750 ;
        RECT 87.620 130.745 87.960 131.575 ;
        RECT 90.175 131.120 90.695 131.660 ;
        RECT 90.865 130.950 91.385 131.490 ;
        RECT 93.150 131.065 93.500 132.315 ;
        RECT 97.275 132.080 97.555 132.750 ;
        RECT 97.725 131.860 98.025 132.410 ;
        RECT 98.225 132.030 98.555 132.750 ;
        RECT 98.745 132.030 99.205 132.580 ;
        RECT 78.680 130.200 84.025 130.745 ;
        RECT 84.200 130.200 89.545 130.745 ;
        RECT 89.715 130.200 90.005 130.925 ;
        RECT 90.175 130.200 91.385 130.950 ;
        RECT 94.980 130.745 95.320 131.575 ;
        RECT 97.090 131.440 97.355 131.800 ;
        RECT 97.725 131.690 98.665 131.860 ;
        RECT 98.495 131.440 98.665 131.690 ;
        RECT 97.090 131.190 97.765 131.440 ;
        RECT 97.985 131.190 98.325 131.440 ;
        RECT 98.495 131.110 98.785 131.440 ;
        RECT 98.495 131.020 98.665 131.110 ;
        RECT 97.275 130.830 98.665 131.020 ;
        RECT 91.560 130.200 96.905 130.745 ;
        RECT 97.275 130.470 97.605 130.830 ;
        RECT 98.955 130.660 99.205 132.030 ;
        RECT 98.225 130.200 98.475 130.660 ;
        RECT 98.645 130.370 99.205 130.660 ;
        RECT 99.375 132.030 99.835 132.580 ;
        RECT 100.025 132.030 100.355 132.750 ;
        RECT 99.375 130.660 99.625 132.030 ;
        RECT 100.555 131.860 100.855 132.410 ;
        RECT 101.025 132.080 101.305 132.750 ;
        RECT 99.915 131.690 100.855 131.860 ;
        RECT 99.915 131.440 100.085 131.690 ;
        RECT 101.225 131.440 101.490 131.800 ;
        RECT 99.795 131.110 100.085 131.440 ;
        RECT 100.255 131.190 100.595 131.440 ;
        RECT 100.815 131.190 101.490 131.440 ;
        RECT 101.675 131.660 103.345 132.750 ;
        RECT 103.520 132.315 108.865 132.750 ;
        RECT 109.040 132.315 114.385 132.750 ;
        RECT 101.675 131.140 102.425 131.660 ;
        RECT 99.915 131.020 100.085 131.110 ;
        RECT 99.915 130.830 101.305 131.020 ;
        RECT 102.595 130.970 103.345 131.490 ;
        RECT 105.110 131.065 105.460 132.315 ;
        RECT 99.375 130.370 99.935 130.660 ;
        RECT 100.105 130.200 100.355 130.660 ;
        RECT 100.975 130.470 101.305 130.830 ;
        RECT 101.675 130.200 103.345 130.970 ;
        RECT 106.940 130.745 107.280 131.575 ;
        RECT 110.630 131.065 110.980 132.315 ;
        RECT 114.555 131.660 115.765 132.750 ;
        RECT 112.460 130.745 112.800 131.575 ;
        RECT 114.555 131.120 115.075 131.660 ;
        RECT 115.245 130.950 115.765 131.490 ;
        RECT 103.520 130.200 108.865 130.745 ;
        RECT 109.040 130.200 114.385 130.745 ;
        RECT 114.555 130.200 115.765 130.950 ;
        RECT 10.510 130.030 115.850 130.200 ;
        RECT 10.595 129.280 11.805 130.030 ;
        RECT 12.985 129.480 13.155 129.770 ;
        RECT 13.325 129.650 13.655 130.030 ;
        RECT 12.985 129.310 13.650 129.480 ;
        RECT 10.595 128.740 11.115 129.280 ;
        RECT 11.285 128.570 11.805 129.110 ;
        RECT 10.595 127.480 11.805 128.570 ;
        RECT 12.900 128.490 13.250 129.140 ;
        RECT 13.420 128.320 13.650 129.310 ;
        RECT 12.985 128.150 13.650 128.320 ;
        RECT 12.985 127.650 13.155 128.150 ;
        RECT 13.325 127.480 13.655 127.980 ;
        RECT 13.825 127.650 14.050 129.770 ;
        RECT 14.265 129.650 14.595 130.030 ;
        RECT 14.765 129.480 14.935 129.810 ;
        RECT 15.235 129.650 16.250 129.850 ;
        RECT 14.240 129.290 14.935 129.480 ;
        RECT 14.240 128.320 14.410 129.290 ;
        RECT 14.580 128.490 14.990 129.110 ;
        RECT 15.160 128.540 15.380 129.410 ;
        RECT 15.560 129.100 15.910 129.470 ;
        RECT 16.080 128.920 16.250 129.650 ;
        RECT 16.420 129.590 16.830 130.030 ;
        RECT 17.120 129.390 17.370 129.820 ;
        RECT 17.570 129.570 17.890 130.030 ;
        RECT 18.450 129.640 19.300 129.810 ;
        RECT 16.420 129.050 16.830 129.380 ;
        RECT 17.120 129.050 17.540 129.390 ;
        RECT 15.830 128.880 16.250 128.920 ;
        RECT 15.830 128.710 17.180 128.880 ;
        RECT 14.240 128.150 14.935 128.320 ;
        RECT 15.160 128.160 15.660 128.540 ;
        RECT 14.265 127.480 14.595 127.980 ;
        RECT 14.765 127.650 14.935 128.150 ;
        RECT 15.830 127.865 16.000 128.710 ;
        RECT 16.930 128.550 17.180 128.710 ;
        RECT 16.170 128.280 16.420 128.540 ;
        RECT 17.350 128.280 17.540 129.050 ;
        RECT 16.170 128.030 17.540 128.280 ;
        RECT 17.710 129.220 18.960 129.390 ;
        RECT 17.710 128.460 17.880 129.220 ;
        RECT 18.630 129.100 18.960 129.220 ;
        RECT 18.050 128.640 18.230 129.050 ;
        RECT 19.130 128.880 19.300 129.640 ;
        RECT 19.500 129.550 20.160 130.030 ;
        RECT 20.340 129.435 20.660 129.765 ;
        RECT 19.490 129.110 20.150 129.380 ;
        RECT 19.490 129.050 19.820 129.110 ;
        RECT 19.970 128.880 20.300 128.940 ;
        RECT 18.400 128.710 20.300 128.880 ;
        RECT 17.710 128.150 18.230 128.460 ;
        RECT 18.400 128.200 18.570 128.710 ;
        RECT 20.470 128.540 20.660 129.435 ;
        RECT 18.740 128.370 20.660 128.540 ;
        RECT 20.340 128.350 20.660 128.370 ;
        RECT 20.860 129.120 21.110 129.770 ;
        RECT 21.290 129.570 21.575 130.030 ;
        RECT 21.755 129.690 22.010 129.850 ;
        RECT 21.755 129.520 22.095 129.690 ;
        RECT 21.755 129.320 22.010 129.520 ;
        RECT 20.860 128.790 21.660 129.120 ;
        RECT 18.400 128.030 19.610 128.200 ;
        RECT 15.170 127.695 16.000 127.865 ;
        RECT 16.240 127.480 16.620 127.860 ;
        RECT 16.800 127.740 16.970 128.030 ;
        RECT 18.400 127.950 18.570 128.030 ;
        RECT 17.140 127.480 17.470 127.860 ;
        RECT 17.940 127.700 18.570 127.950 ;
        RECT 18.750 127.480 19.170 127.860 ;
        RECT 19.370 127.740 19.610 128.030 ;
        RECT 19.840 127.480 20.170 128.170 ;
        RECT 20.340 127.740 20.510 128.350 ;
        RECT 20.860 128.200 21.110 128.790 ;
        RECT 21.830 128.460 22.010 129.320 ;
        RECT 22.555 129.260 25.145 130.030 ;
        RECT 25.315 129.305 25.605 130.030 ;
        RECT 25.865 129.480 26.035 129.770 ;
        RECT 26.205 129.650 26.535 130.030 ;
        RECT 25.865 129.310 26.530 129.480 ;
        RECT 20.780 127.690 21.110 128.200 ;
        RECT 21.290 127.480 21.575 128.280 ;
        RECT 21.755 127.790 22.010 128.460 ;
        RECT 22.555 128.570 23.765 129.090 ;
        RECT 23.935 128.740 25.145 129.260 ;
        RECT 22.555 127.480 25.145 128.570 ;
        RECT 25.315 127.480 25.605 128.645 ;
        RECT 25.780 128.490 26.130 129.140 ;
        RECT 26.300 128.320 26.530 129.310 ;
        RECT 25.865 128.150 26.530 128.320 ;
        RECT 25.865 127.650 26.035 128.150 ;
        RECT 26.205 127.480 26.535 127.980 ;
        RECT 26.705 127.650 26.930 129.770 ;
        RECT 27.145 129.650 27.475 130.030 ;
        RECT 27.645 129.480 27.815 129.810 ;
        RECT 28.115 129.650 29.130 129.850 ;
        RECT 27.120 129.290 27.815 129.480 ;
        RECT 27.120 128.320 27.290 129.290 ;
        RECT 27.460 128.490 27.870 129.110 ;
        RECT 28.040 128.540 28.260 129.410 ;
        RECT 28.440 129.100 28.790 129.470 ;
        RECT 28.960 128.920 29.130 129.650 ;
        RECT 29.300 129.590 29.710 130.030 ;
        RECT 30.000 129.390 30.250 129.820 ;
        RECT 30.450 129.570 30.770 130.030 ;
        RECT 31.330 129.640 32.180 129.810 ;
        RECT 29.300 129.050 29.710 129.380 ;
        RECT 30.000 129.050 30.420 129.390 ;
        RECT 28.710 128.880 29.130 128.920 ;
        RECT 28.710 128.710 30.060 128.880 ;
        RECT 27.120 128.150 27.815 128.320 ;
        RECT 28.040 128.160 28.540 128.540 ;
        RECT 27.145 127.480 27.475 127.980 ;
        RECT 27.645 127.650 27.815 128.150 ;
        RECT 28.710 127.865 28.880 128.710 ;
        RECT 29.810 128.550 30.060 128.710 ;
        RECT 29.050 128.280 29.300 128.540 ;
        RECT 30.230 128.280 30.420 129.050 ;
        RECT 29.050 128.030 30.420 128.280 ;
        RECT 30.590 129.220 31.840 129.390 ;
        RECT 30.590 128.460 30.760 129.220 ;
        RECT 31.510 129.100 31.840 129.220 ;
        RECT 30.930 128.640 31.110 129.050 ;
        RECT 32.010 128.880 32.180 129.640 ;
        RECT 32.380 129.550 33.040 130.030 ;
        RECT 33.220 129.435 33.540 129.765 ;
        RECT 32.370 129.110 33.030 129.380 ;
        RECT 32.370 129.050 32.700 129.110 ;
        RECT 32.850 128.880 33.180 128.940 ;
        RECT 31.280 128.710 33.180 128.880 ;
        RECT 30.590 128.150 31.110 128.460 ;
        RECT 31.280 128.200 31.450 128.710 ;
        RECT 33.350 128.540 33.540 129.435 ;
        RECT 31.620 128.370 33.540 128.540 ;
        RECT 33.220 128.350 33.540 128.370 ;
        RECT 33.740 129.120 33.990 129.770 ;
        RECT 34.170 129.570 34.455 130.030 ;
        RECT 34.635 129.690 34.890 129.850 ;
        RECT 34.635 129.520 34.975 129.690 ;
        RECT 34.635 129.320 34.890 129.520 ;
        RECT 33.740 128.790 34.540 129.120 ;
        RECT 31.280 128.030 32.490 128.200 ;
        RECT 28.050 127.695 28.880 127.865 ;
        RECT 29.120 127.480 29.500 127.860 ;
        RECT 29.680 127.740 29.850 128.030 ;
        RECT 31.280 127.950 31.450 128.030 ;
        RECT 30.020 127.480 30.350 127.860 ;
        RECT 30.820 127.700 31.450 127.950 ;
        RECT 31.630 127.480 32.050 127.860 ;
        RECT 32.250 127.740 32.490 128.030 ;
        RECT 32.720 127.480 33.050 128.170 ;
        RECT 33.220 127.740 33.390 128.350 ;
        RECT 33.740 128.200 33.990 128.790 ;
        RECT 34.710 128.460 34.890 129.320 ;
        RECT 36.095 129.400 36.425 129.760 ;
        RECT 37.045 129.570 37.295 130.030 ;
        RECT 37.465 129.570 38.025 129.860 ;
        RECT 36.095 129.210 37.485 129.400 ;
        RECT 37.315 129.120 37.485 129.210 ;
        RECT 33.660 127.690 33.990 128.200 ;
        RECT 34.170 127.480 34.455 128.280 ;
        RECT 34.635 127.790 34.890 128.460 ;
        RECT 35.910 128.790 36.585 129.040 ;
        RECT 36.805 128.790 37.145 129.040 ;
        RECT 37.315 128.790 37.605 129.120 ;
        RECT 35.910 128.430 36.175 128.790 ;
        RECT 37.315 128.540 37.485 128.790 ;
        RECT 36.545 128.370 37.485 128.540 ;
        RECT 36.095 127.480 36.375 128.150 ;
        RECT 36.545 127.820 36.845 128.370 ;
        RECT 37.775 128.200 38.025 129.570 ;
        RECT 37.045 127.480 37.375 128.200 ;
        RECT 37.565 127.650 38.025 128.200 ;
        RECT 38.195 129.570 38.755 129.860 ;
        RECT 38.925 129.570 39.175 130.030 ;
        RECT 38.195 128.200 38.445 129.570 ;
        RECT 39.795 129.400 40.125 129.760 ;
        RECT 38.735 129.210 40.125 129.400 ;
        RECT 40.695 129.400 41.025 129.760 ;
        RECT 41.645 129.570 41.895 130.030 ;
        RECT 42.065 129.570 42.625 129.860 ;
        RECT 40.695 129.210 42.085 129.400 ;
        RECT 38.735 129.120 38.905 129.210 ;
        RECT 38.615 128.790 38.905 129.120 ;
        RECT 41.915 129.120 42.085 129.210 ;
        RECT 39.075 128.790 39.415 129.040 ;
        RECT 39.635 128.790 40.310 129.040 ;
        RECT 38.735 128.540 38.905 128.790 ;
        RECT 38.735 128.370 39.675 128.540 ;
        RECT 40.045 128.430 40.310 128.790 ;
        RECT 40.510 128.790 41.185 129.040 ;
        RECT 41.405 128.790 41.745 129.040 ;
        RECT 41.915 128.790 42.205 129.120 ;
        RECT 40.510 128.430 40.775 128.790 ;
        RECT 41.915 128.540 42.085 128.790 ;
        RECT 38.195 127.650 38.655 128.200 ;
        RECT 38.845 127.480 39.175 128.200 ;
        RECT 39.375 127.820 39.675 128.370 ;
        RECT 41.145 128.370 42.085 128.540 ;
        RECT 39.845 127.480 40.125 128.150 ;
        RECT 40.695 127.480 40.975 128.150 ;
        RECT 41.145 127.820 41.445 128.370 ;
        RECT 42.375 128.200 42.625 129.570 ;
        RECT 42.855 129.550 43.135 130.030 ;
        RECT 43.305 129.380 43.565 129.770 ;
        RECT 43.740 129.550 43.995 130.030 ;
        RECT 44.165 129.380 44.460 129.770 ;
        RECT 44.640 129.550 44.915 130.030 ;
        RECT 45.085 129.530 45.385 129.860 ;
        RECT 42.810 129.210 44.460 129.380 ;
        RECT 42.810 128.700 43.215 129.210 ;
        RECT 43.385 128.870 44.525 129.040 ;
        RECT 42.810 128.530 43.565 128.700 ;
        RECT 41.645 127.480 41.975 128.200 ;
        RECT 42.165 127.650 42.625 128.200 ;
        RECT 42.850 127.480 43.135 128.350 ;
        RECT 43.305 128.280 43.565 128.530 ;
        RECT 44.355 128.620 44.525 128.870 ;
        RECT 44.695 128.790 45.045 129.360 ;
        RECT 45.215 128.620 45.385 129.530 ;
        RECT 45.615 129.210 45.825 130.030 ;
        RECT 45.995 129.230 46.325 129.860 ;
        RECT 45.995 128.630 46.245 129.230 ;
        RECT 46.495 129.210 46.725 130.030 ;
        RECT 47.210 129.220 47.455 129.825 ;
        RECT 47.675 129.495 48.185 130.030 ;
        RECT 46.935 129.050 48.165 129.220 ;
        RECT 46.415 128.790 46.745 129.040 ;
        RECT 44.355 128.450 45.385 128.620 ;
        RECT 43.305 128.110 44.425 128.280 ;
        RECT 43.305 127.650 43.565 128.110 ;
        RECT 43.740 127.480 43.995 127.940 ;
        RECT 44.165 127.650 44.425 128.110 ;
        RECT 44.595 127.480 44.905 128.280 ;
        RECT 45.075 127.650 45.385 128.450 ;
        RECT 45.615 127.480 45.825 128.620 ;
        RECT 45.995 127.650 46.325 128.630 ;
        RECT 46.495 127.480 46.725 128.620 ;
        RECT 46.935 128.240 47.275 129.050 ;
        RECT 47.445 128.485 48.195 128.675 ;
        RECT 46.935 127.830 47.450 128.240 ;
        RECT 47.685 127.480 47.855 128.240 ;
        RECT 48.025 127.820 48.195 128.485 ;
        RECT 48.365 128.500 48.555 129.860 ;
        RECT 48.725 129.690 49.000 129.860 ;
        RECT 48.725 129.520 49.005 129.690 ;
        RECT 48.725 128.700 49.000 129.520 ;
        RECT 49.190 129.495 49.720 129.860 ;
        RECT 50.145 129.630 50.475 130.030 ;
        RECT 49.545 129.460 49.720 129.495 ;
        RECT 49.205 128.500 49.375 129.300 ;
        RECT 48.365 128.330 49.375 128.500 ;
        RECT 49.545 129.290 50.475 129.460 ;
        RECT 50.645 129.290 50.900 129.860 ;
        RECT 51.075 129.305 51.365 130.030 ;
        RECT 49.545 128.160 49.715 129.290 ;
        RECT 50.305 129.120 50.475 129.290 ;
        RECT 48.590 127.990 49.715 128.160 ;
        RECT 49.885 128.790 50.080 129.120 ;
        RECT 50.305 128.790 50.560 129.120 ;
        RECT 49.885 127.820 50.055 128.790 ;
        RECT 50.730 128.620 50.900 129.290 ;
        RECT 51.995 129.260 53.665 130.030 ;
        RECT 48.025 127.650 50.055 127.820 ;
        RECT 50.225 127.480 50.395 128.620 ;
        RECT 50.565 127.650 50.900 128.620 ;
        RECT 51.075 127.480 51.365 128.645 ;
        RECT 51.995 128.570 52.745 129.090 ;
        RECT 52.915 128.740 53.665 129.260 ;
        RECT 53.875 129.210 54.105 130.030 ;
        RECT 54.275 129.230 54.605 129.860 ;
        RECT 53.855 128.790 54.185 129.040 ;
        RECT 54.355 128.630 54.605 129.230 ;
        RECT 54.775 129.210 54.985 130.030 ;
        RECT 55.765 129.480 55.935 129.860 ;
        RECT 56.115 129.650 56.445 130.030 ;
        RECT 55.765 129.310 56.430 129.480 ;
        RECT 56.625 129.355 56.885 129.860 ;
        RECT 55.695 128.760 56.025 129.130 ;
        RECT 56.260 129.055 56.430 129.310 ;
        RECT 51.995 127.480 53.665 128.570 ;
        RECT 53.875 127.480 54.105 128.620 ;
        RECT 54.275 127.650 54.605 128.630 ;
        RECT 56.260 128.725 56.545 129.055 ;
        RECT 54.775 127.480 54.985 128.620 ;
        RECT 56.260 128.580 56.430 128.725 ;
        RECT 55.765 128.410 56.430 128.580 ;
        RECT 56.715 128.555 56.885 129.355 ;
        RECT 57.055 129.260 58.725 130.030 ;
        RECT 58.900 129.485 64.245 130.030 ;
        RECT 64.415 129.530 64.715 129.860 ;
        RECT 64.885 129.550 65.160 130.030 ;
        RECT 55.765 127.650 55.935 128.410 ;
        RECT 56.115 127.480 56.445 128.240 ;
        RECT 56.615 127.650 56.885 128.555 ;
        RECT 57.055 128.570 57.805 129.090 ;
        RECT 57.975 128.740 58.725 129.260 ;
        RECT 57.055 127.480 58.725 128.570 ;
        RECT 60.490 127.915 60.840 129.165 ;
        RECT 62.320 128.655 62.660 129.485 ;
        RECT 64.415 128.620 64.585 129.530 ;
        RECT 65.340 129.380 65.635 129.770 ;
        RECT 65.805 129.550 66.060 130.030 ;
        RECT 66.235 129.380 66.495 129.770 ;
        RECT 66.665 129.550 66.945 130.030 ;
        RECT 64.755 128.790 65.105 129.360 ;
        RECT 65.340 129.210 66.990 129.380 ;
        RECT 65.275 128.870 66.415 129.040 ;
        RECT 65.275 128.620 65.445 128.870 ;
        RECT 66.585 128.700 66.990 129.210 ;
        RECT 64.415 128.450 65.445 128.620 ;
        RECT 66.235 128.530 66.990 128.700 ;
        RECT 67.550 129.320 67.805 129.850 ;
        RECT 67.985 129.570 68.270 130.030 ;
        RECT 67.550 128.670 67.730 129.320 ;
        RECT 68.450 129.120 68.700 129.770 ;
        RECT 67.900 128.790 68.700 129.120 ;
        RECT 58.900 127.480 64.245 127.915 ;
        RECT 64.415 127.650 64.725 128.450 ;
        RECT 66.235 128.280 66.495 128.530 ;
        RECT 67.465 128.500 67.730 128.670 ;
        RECT 67.550 128.460 67.730 128.500 ;
        RECT 64.895 127.480 65.205 128.280 ;
        RECT 65.375 128.110 66.495 128.280 ;
        RECT 65.375 127.650 65.635 128.110 ;
        RECT 65.805 127.480 66.060 127.940 ;
        RECT 66.235 127.650 66.495 128.110 ;
        RECT 66.665 127.480 66.950 128.350 ;
        RECT 67.550 127.790 67.805 128.460 ;
        RECT 67.985 127.480 68.270 128.280 ;
        RECT 68.450 128.200 68.700 128.790 ;
        RECT 68.900 129.435 69.220 129.765 ;
        RECT 69.400 129.550 70.060 130.030 ;
        RECT 70.260 129.640 71.110 129.810 ;
        RECT 68.900 128.540 69.090 129.435 ;
        RECT 69.410 129.110 70.070 129.380 ;
        RECT 69.740 129.050 70.070 129.110 ;
        RECT 69.260 128.880 69.590 128.940 ;
        RECT 70.260 128.880 70.430 129.640 ;
        RECT 71.670 129.570 71.990 130.030 ;
        RECT 72.190 129.390 72.440 129.820 ;
        RECT 72.730 129.590 73.140 130.030 ;
        RECT 73.310 129.650 74.325 129.850 ;
        RECT 70.600 129.220 71.850 129.390 ;
        RECT 70.600 129.100 70.930 129.220 ;
        RECT 69.260 128.710 71.160 128.880 ;
        RECT 68.900 128.370 70.820 128.540 ;
        RECT 68.900 128.350 69.220 128.370 ;
        RECT 68.450 127.690 68.780 128.200 ;
        RECT 69.050 127.740 69.220 128.350 ;
        RECT 70.990 128.200 71.160 128.710 ;
        RECT 71.330 128.640 71.510 129.050 ;
        RECT 71.680 128.460 71.850 129.220 ;
        RECT 69.390 127.480 69.720 128.170 ;
        RECT 69.950 128.030 71.160 128.200 ;
        RECT 71.330 128.150 71.850 128.460 ;
        RECT 72.020 129.050 72.440 129.390 ;
        RECT 72.730 129.050 73.140 129.380 ;
        RECT 72.020 128.280 72.210 129.050 ;
        RECT 73.310 128.920 73.480 129.650 ;
        RECT 74.625 129.480 74.795 129.810 ;
        RECT 74.965 129.650 75.295 130.030 ;
        RECT 73.650 129.100 74.000 129.470 ;
        RECT 73.310 128.880 73.730 128.920 ;
        RECT 72.380 128.710 73.730 128.880 ;
        RECT 72.380 128.550 72.630 128.710 ;
        RECT 73.140 128.280 73.390 128.540 ;
        RECT 72.020 128.030 73.390 128.280 ;
        RECT 69.950 127.740 70.190 128.030 ;
        RECT 70.990 127.950 71.160 128.030 ;
        RECT 70.390 127.480 70.810 127.860 ;
        RECT 70.990 127.700 71.620 127.950 ;
        RECT 72.090 127.480 72.420 127.860 ;
        RECT 72.590 127.740 72.760 128.030 ;
        RECT 73.560 127.865 73.730 128.710 ;
        RECT 74.180 128.540 74.400 129.410 ;
        RECT 74.625 129.290 75.320 129.480 ;
        RECT 73.900 128.160 74.400 128.540 ;
        RECT 74.570 128.490 74.980 129.110 ;
        RECT 75.150 128.320 75.320 129.290 ;
        RECT 74.625 128.150 75.320 128.320 ;
        RECT 72.940 127.480 73.320 127.860 ;
        RECT 73.560 127.695 74.390 127.865 ;
        RECT 74.625 127.650 74.795 128.150 ;
        RECT 74.965 127.480 75.295 127.980 ;
        RECT 75.510 127.650 75.735 129.770 ;
        RECT 75.905 129.650 76.235 130.030 ;
        RECT 76.405 129.480 76.575 129.770 ;
        RECT 75.910 129.310 76.575 129.480 ;
        RECT 75.910 128.320 76.140 129.310 ;
        RECT 76.835 129.305 77.125 130.030 ;
        RECT 77.295 129.355 77.555 129.860 ;
        RECT 77.735 129.650 78.065 130.030 ;
        RECT 78.245 129.480 78.415 129.860 ;
        RECT 76.310 128.490 76.660 129.140 ;
        RECT 75.910 128.150 76.575 128.320 ;
        RECT 75.905 127.480 76.235 127.980 ;
        RECT 76.405 127.650 76.575 128.150 ;
        RECT 76.835 127.480 77.125 128.645 ;
        RECT 77.295 128.555 77.465 129.355 ;
        RECT 77.750 129.310 78.415 129.480 ;
        RECT 77.750 129.055 77.920 129.310 ;
        RECT 79.135 129.260 80.805 130.030 ;
        RECT 77.635 128.725 77.920 129.055 ;
        RECT 78.155 128.760 78.485 129.130 ;
        RECT 77.750 128.580 77.920 128.725 ;
        RECT 77.295 127.650 77.565 128.555 ;
        RECT 77.750 128.410 78.415 128.580 ;
        RECT 77.735 127.480 78.065 128.240 ;
        RECT 78.245 127.650 78.415 128.410 ;
        RECT 79.135 128.570 79.885 129.090 ;
        RECT 80.055 128.740 80.805 129.260 ;
        RECT 81.250 129.220 81.495 129.825 ;
        RECT 81.715 129.495 82.225 130.030 ;
        RECT 80.975 129.050 82.205 129.220 ;
        RECT 79.135 127.480 80.805 128.570 ;
        RECT 80.975 128.240 81.315 129.050 ;
        RECT 81.485 128.485 82.235 128.675 ;
        RECT 80.975 127.830 81.490 128.240 ;
        RECT 81.725 127.480 81.895 128.240 ;
        RECT 82.065 127.820 82.235 128.485 ;
        RECT 82.405 128.500 82.595 129.860 ;
        RECT 82.765 129.350 83.040 129.860 ;
        RECT 83.230 129.495 83.760 129.860 ;
        RECT 84.185 129.630 84.515 130.030 ;
        RECT 83.585 129.460 83.760 129.495 ;
        RECT 82.765 129.180 83.045 129.350 ;
        RECT 82.765 128.700 83.040 129.180 ;
        RECT 83.245 128.500 83.415 129.300 ;
        RECT 82.405 128.330 83.415 128.500 ;
        RECT 83.585 129.290 84.515 129.460 ;
        RECT 84.685 129.290 84.940 129.860 ;
        RECT 83.585 128.160 83.755 129.290 ;
        RECT 84.345 129.120 84.515 129.290 ;
        RECT 82.630 127.990 83.755 128.160 ;
        RECT 83.925 128.790 84.120 129.120 ;
        RECT 84.345 128.790 84.600 129.120 ;
        RECT 83.925 127.820 84.095 128.790 ;
        RECT 84.770 128.620 84.940 129.290 ;
        RECT 82.065 127.650 84.095 127.820 ;
        RECT 84.265 127.480 84.435 128.620 ;
        RECT 84.605 127.650 84.940 128.620 ;
        RECT 85.575 129.355 85.835 129.860 ;
        RECT 86.015 129.650 86.345 130.030 ;
        RECT 86.525 129.480 86.695 129.860 ;
        RECT 85.575 128.555 85.745 129.355 ;
        RECT 86.030 129.310 86.695 129.480 ;
        RECT 87.155 129.400 87.485 129.760 ;
        RECT 88.105 129.570 88.355 130.030 ;
        RECT 88.525 129.570 89.085 129.860 ;
        RECT 86.030 129.055 86.200 129.310 ;
        RECT 87.155 129.210 88.545 129.400 ;
        RECT 85.915 128.725 86.200 129.055 ;
        RECT 86.435 128.760 86.765 129.130 ;
        RECT 88.375 129.120 88.545 129.210 ;
        RECT 86.970 128.790 87.645 129.040 ;
        RECT 87.865 128.790 88.205 129.040 ;
        RECT 88.375 128.790 88.665 129.120 ;
        RECT 86.030 128.580 86.200 128.725 ;
        RECT 85.575 127.650 85.845 128.555 ;
        RECT 86.030 128.410 86.695 128.580 ;
        RECT 86.970 128.430 87.235 128.790 ;
        RECT 88.375 128.540 88.545 128.790 ;
        RECT 86.015 127.480 86.345 128.240 ;
        RECT 86.525 127.650 86.695 128.410 ;
        RECT 87.605 128.370 88.545 128.540 ;
        RECT 87.155 127.480 87.435 128.150 ;
        RECT 87.605 127.820 87.905 128.370 ;
        RECT 88.835 128.200 89.085 129.570 ;
        RECT 89.715 129.260 93.225 130.030 ;
        RECT 88.105 127.480 88.435 128.200 ;
        RECT 88.625 127.650 89.085 128.200 ;
        RECT 89.715 128.570 91.405 129.090 ;
        RECT 91.575 128.740 93.225 129.260 ;
        RECT 93.395 129.570 93.955 129.860 ;
        RECT 94.125 129.570 94.375 130.030 ;
        RECT 89.715 127.480 93.225 128.570 ;
        RECT 93.395 128.200 93.645 129.570 ;
        RECT 94.995 129.400 95.325 129.760 ;
        RECT 93.935 129.210 95.325 129.400 ;
        RECT 96.155 129.570 96.715 129.860 ;
        RECT 96.885 129.570 97.135 130.030 ;
        RECT 93.935 129.120 94.105 129.210 ;
        RECT 93.815 128.790 94.105 129.120 ;
        RECT 94.275 128.790 94.615 129.040 ;
        RECT 94.835 128.790 95.510 129.040 ;
        RECT 93.935 128.540 94.105 128.790 ;
        RECT 93.935 128.370 94.875 128.540 ;
        RECT 95.245 128.430 95.510 128.790 ;
        RECT 93.395 127.650 93.855 128.200 ;
        RECT 94.045 127.480 94.375 128.200 ;
        RECT 94.575 127.820 94.875 128.370 ;
        RECT 96.155 128.200 96.405 129.570 ;
        RECT 97.755 129.400 98.085 129.760 ;
        RECT 96.695 129.210 98.085 129.400 ;
        RECT 98.730 129.220 98.975 129.825 ;
        RECT 99.195 129.495 99.705 130.030 ;
        RECT 96.695 129.120 96.865 129.210 ;
        RECT 96.575 128.790 96.865 129.120 ;
        RECT 98.455 129.050 99.685 129.220 ;
        RECT 97.035 128.790 97.375 129.040 ;
        RECT 97.595 128.790 98.270 129.040 ;
        RECT 96.695 128.540 96.865 128.790 ;
        RECT 96.695 128.370 97.635 128.540 ;
        RECT 98.005 128.430 98.270 128.790 ;
        RECT 95.045 127.480 95.325 128.150 ;
        RECT 96.155 127.650 96.615 128.200 ;
        RECT 96.805 127.480 97.135 128.200 ;
        RECT 97.335 127.820 97.635 128.370 ;
        RECT 98.455 128.240 98.795 129.050 ;
        RECT 98.965 128.485 99.715 128.675 ;
        RECT 97.805 127.480 98.085 128.150 ;
        RECT 98.455 127.830 98.970 128.240 ;
        RECT 99.205 127.480 99.375 128.240 ;
        RECT 99.545 127.820 99.715 128.485 ;
        RECT 99.885 128.500 100.075 129.860 ;
        RECT 100.245 129.010 100.520 129.860 ;
        RECT 100.710 129.495 101.240 129.860 ;
        RECT 101.665 129.630 101.995 130.030 ;
        RECT 101.065 129.460 101.240 129.495 ;
        RECT 100.245 128.840 100.525 129.010 ;
        RECT 100.245 128.700 100.520 128.840 ;
        RECT 100.725 128.500 100.895 129.300 ;
        RECT 99.885 128.330 100.895 128.500 ;
        RECT 101.065 129.290 101.995 129.460 ;
        RECT 102.165 129.290 102.420 129.860 ;
        RECT 102.595 129.305 102.885 130.030 ;
        RECT 103.055 129.570 103.615 129.860 ;
        RECT 103.785 129.570 104.035 130.030 ;
        RECT 101.065 128.160 101.235 129.290 ;
        RECT 101.825 129.120 101.995 129.290 ;
        RECT 100.110 127.990 101.235 128.160 ;
        RECT 101.405 128.790 101.600 129.120 ;
        RECT 101.825 128.790 102.080 129.120 ;
        RECT 101.405 127.820 101.575 128.790 ;
        RECT 102.250 128.620 102.420 129.290 ;
        RECT 99.545 127.650 101.575 127.820 ;
        RECT 101.745 127.480 101.915 128.620 ;
        RECT 102.085 127.650 102.420 128.620 ;
        RECT 102.595 127.480 102.885 128.645 ;
        RECT 103.055 128.200 103.305 129.570 ;
        RECT 104.655 129.400 104.985 129.760 ;
        RECT 103.595 129.210 104.985 129.400 ;
        RECT 105.355 129.280 106.565 130.030 ;
        RECT 103.595 129.120 103.765 129.210 ;
        RECT 103.475 128.790 103.765 129.120 ;
        RECT 103.935 128.790 104.275 129.040 ;
        RECT 104.495 128.790 105.170 129.040 ;
        RECT 103.595 128.540 103.765 128.790 ;
        RECT 103.595 128.370 104.535 128.540 ;
        RECT 104.905 128.430 105.170 128.790 ;
        RECT 105.355 128.570 105.875 129.110 ;
        RECT 106.045 128.740 106.565 129.280 ;
        RECT 106.775 129.210 107.005 130.030 ;
        RECT 107.175 129.230 107.505 129.860 ;
        RECT 106.755 128.790 107.085 129.040 ;
        RECT 107.255 128.630 107.505 129.230 ;
        RECT 107.675 129.210 107.885 130.030 ;
        RECT 108.665 129.480 108.835 129.860 ;
        RECT 109.015 129.650 109.345 130.030 ;
        RECT 108.665 129.310 109.330 129.480 ;
        RECT 109.525 129.355 109.785 129.860 ;
        RECT 108.595 128.760 108.925 129.130 ;
        RECT 109.160 129.055 109.330 129.310 ;
        RECT 103.055 127.650 103.515 128.200 ;
        RECT 103.705 127.480 104.035 128.200 ;
        RECT 104.235 127.820 104.535 128.370 ;
        RECT 104.705 127.480 104.985 128.150 ;
        RECT 105.355 127.480 106.565 128.570 ;
        RECT 106.775 127.480 107.005 128.620 ;
        RECT 107.175 127.650 107.505 128.630 ;
        RECT 109.160 128.725 109.445 129.055 ;
        RECT 107.675 127.480 107.885 128.620 ;
        RECT 109.160 128.580 109.330 128.725 ;
        RECT 108.665 128.410 109.330 128.580 ;
        RECT 109.615 128.555 109.785 129.355 ;
        RECT 110.875 129.260 114.385 130.030 ;
        RECT 114.555 129.280 115.765 130.030 ;
        RECT 108.665 127.650 108.835 128.410 ;
        RECT 109.015 127.480 109.345 128.240 ;
        RECT 109.515 127.650 109.785 128.555 ;
        RECT 110.875 128.570 112.565 129.090 ;
        RECT 112.735 128.740 114.385 129.260 ;
        RECT 114.555 128.570 115.075 129.110 ;
        RECT 115.245 128.740 115.765 129.280 ;
        RECT 110.875 127.480 114.385 128.570 ;
        RECT 114.555 127.480 115.765 128.570 ;
        RECT 10.510 127.310 115.850 127.480 ;
        RECT 10.595 126.220 11.805 127.310 ;
        RECT 10.595 125.510 11.115 126.050 ;
        RECT 11.285 125.680 11.805 126.220 ;
        RECT 12.435 126.145 12.725 127.310 ;
        RECT 12.895 126.220 14.565 127.310 ;
        RECT 12.895 125.700 13.645 126.220 ;
        RECT 14.775 126.170 15.005 127.310 ;
        RECT 15.175 126.160 15.505 127.140 ;
        RECT 15.675 126.170 15.885 127.310 ;
        RECT 16.115 126.235 16.385 127.140 ;
        RECT 16.555 126.550 16.885 127.310 ;
        RECT 17.065 126.380 17.235 127.140 ;
        RECT 13.815 125.530 14.565 126.050 ;
        RECT 14.755 125.750 15.085 126.000 ;
        RECT 10.595 124.760 11.805 125.510 ;
        RECT 12.435 124.760 12.725 125.485 ;
        RECT 12.895 124.760 14.565 125.530 ;
        RECT 14.775 124.760 15.005 125.580 ;
        RECT 15.255 125.560 15.505 126.160 ;
        RECT 15.175 124.930 15.505 125.560 ;
        RECT 15.675 124.760 15.885 125.580 ;
        RECT 16.115 125.435 16.285 126.235 ;
        RECT 16.570 126.210 17.235 126.380 ;
        RECT 16.570 126.065 16.740 126.210 ;
        RECT 16.455 125.735 16.740 126.065 ;
        RECT 17.500 126.170 17.835 127.140 ;
        RECT 18.005 126.170 18.175 127.310 ;
        RECT 18.345 126.970 20.375 127.140 ;
        RECT 16.570 125.480 16.740 125.735 ;
        RECT 16.975 125.660 17.305 126.030 ;
        RECT 17.500 125.500 17.670 126.170 ;
        RECT 18.345 126.000 18.515 126.970 ;
        RECT 17.840 125.670 18.095 126.000 ;
        RECT 18.320 125.670 18.515 126.000 ;
        RECT 18.685 126.630 19.810 126.800 ;
        RECT 17.925 125.500 18.095 125.670 ;
        RECT 18.685 125.500 18.855 126.630 ;
        RECT 16.115 124.930 16.375 125.435 ;
        RECT 16.570 125.310 17.235 125.480 ;
        RECT 16.555 124.760 16.885 125.140 ;
        RECT 17.065 124.930 17.235 125.310 ;
        RECT 17.500 124.930 17.755 125.500 ;
        RECT 17.925 125.330 18.855 125.500 ;
        RECT 19.025 126.290 20.035 126.460 ;
        RECT 19.025 125.490 19.195 126.290 ;
        RECT 19.400 125.610 19.675 126.090 ;
        RECT 19.395 125.440 19.675 125.610 ;
        RECT 18.680 125.295 18.855 125.330 ;
        RECT 17.925 124.760 18.255 125.160 ;
        RECT 18.680 124.930 19.210 125.295 ;
        RECT 19.400 124.930 19.675 125.440 ;
        RECT 19.845 124.930 20.035 126.290 ;
        RECT 20.205 126.305 20.375 126.970 ;
        RECT 20.545 126.550 20.715 127.310 ;
        RECT 20.950 126.550 21.465 126.960 ;
        RECT 20.205 126.115 20.955 126.305 ;
        RECT 21.125 125.740 21.465 126.550 ;
        RECT 20.235 125.570 21.465 125.740 ;
        RECT 21.635 126.235 21.905 127.140 ;
        RECT 22.075 126.550 22.405 127.310 ;
        RECT 22.585 126.380 22.755 127.140 ;
        RECT 20.215 124.760 20.725 125.295 ;
        RECT 20.945 124.965 21.190 125.570 ;
        RECT 21.635 125.435 21.805 126.235 ;
        RECT 22.090 126.210 22.755 126.380 ;
        RECT 23.015 126.220 26.525 127.310 ;
        RECT 22.090 126.065 22.260 126.210 ;
        RECT 21.975 125.735 22.260 126.065 ;
        RECT 22.090 125.480 22.260 125.735 ;
        RECT 22.495 125.660 22.825 126.030 ;
        RECT 23.015 125.700 24.705 126.220 ;
        RECT 26.735 126.170 26.965 127.310 ;
        RECT 27.135 126.160 27.465 127.140 ;
        RECT 27.635 126.170 27.845 127.310 ;
        RECT 28.115 126.170 28.345 127.310 ;
        RECT 28.515 126.160 28.845 127.140 ;
        RECT 29.015 126.170 29.225 127.310 ;
        RECT 29.455 126.235 29.725 127.140 ;
        RECT 29.895 126.550 30.225 127.310 ;
        RECT 30.405 126.380 30.575 127.140 ;
        RECT 31.035 126.640 31.315 127.310 ;
        RECT 24.875 125.530 26.525 126.050 ;
        RECT 26.715 125.750 27.045 126.000 ;
        RECT 21.635 124.930 21.895 125.435 ;
        RECT 22.090 125.310 22.755 125.480 ;
        RECT 22.075 124.760 22.405 125.140 ;
        RECT 22.585 124.930 22.755 125.310 ;
        RECT 23.015 124.760 26.525 125.530 ;
        RECT 26.735 124.760 26.965 125.580 ;
        RECT 27.215 125.560 27.465 126.160 ;
        RECT 28.095 125.750 28.425 126.000 ;
        RECT 27.135 124.930 27.465 125.560 ;
        RECT 27.635 124.760 27.845 125.580 ;
        RECT 28.115 124.760 28.345 125.580 ;
        RECT 28.595 125.560 28.845 126.160 ;
        RECT 28.515 124.930 28.845 125.560 ;
        RECT 29.015 124.760 29.225 125.580 ;
        RECT 29.455 125.435 29.625 126.235 ;
        RECT 29.910 126.210 30.575 126.380 ;
        RECT 31.485 126.420 31.785 126.970 ;
        RECT 31.985 126.590 32.315 127.310 ;
        RECT 32.505 126.590 32.965 127.140 ;
        RECT 29.910 126.065 30.080 126.210 ;
        RECT 29.795 125.735 30.080 126.065 ;
        RECT 29.910 125.480 30.080 125.735 ;
        RECT 30.315 125.660 30.645 126.030 ;
        RECT 30.850 126.000 31.115 126.360 ;
        RECT 31.485 126.250 32.425 126.420 ;
        RECT 32.255 126.000 32.425 126.250 ;
        RECT 30.850 125.750 31.525 126.000 ;
        RECT 31.745 125.750 32.085 126.000 ;
        RECT 32.255 125.670 32.545 126.000 ;
        RECT 32.255 125.580 32.425 125.670 ;
        RECT 29.455 124.930 29.715 125.435 ;
        RECT 29.910 125.310 30.575 125.480 ;
        RECT 29.895 124.760 30.225 125.140 ;
        RECT 30.405 124.930 30.575 125.310 ;
        RECT 31.035 125.390 32.425 125.580 ;
        RECT 31.035 125.030 31.365 125.390 ;
        RECT 32.715 125.220 32.965 126.590 ;
        RECT 33.135 126.550 33.650 126.960 ;
        RECT 33.885 126.550 34.055 127.310 ;
        RECT 34.225 126.970 36.255 127.140 ;
        RECT 33.135 125.740 33.475 126.550 ;
        RECT 34.225 126.305 34.395 126.970 ;
        RECT 34.790 126.630 35.915 126.800 ;
        RECT 33.645 126.115 34.395 126.305 ;
        RECT 34.565 126.290 35.575 126.460 ;
        RECT 33.135 125.570 34.365 125.740 ;
        RECT 31.985 124.760 32.235 125.220 ;
        RECT 32.405 124.930 32.965 125.220 ;
        RECT 33.410 124.965 33.655 125.570 ;
        RECT 33.875 124.760 34.385 125.295 ;
        RECT 34.565 124.930 34.755 126.290 ;
        RECT 34.925 125.950 35.200 126.090 ;
        RECT 34.925 125.780 35.205 125.950 ;
        RECT 34.925 124.930 35.200 125.780 ;
        RECT 35.405 125.490 35.575 126.290 ;
        RECT 35.745 125.500 35.915 126.630 ;
        RECT 36.085 126.000 36.255 126.970 ;
        RECT 36.425 126.170 36.595 127.310 ;
        RECT 36.765 126.170 37.100 127.140 ;
        RECT 36.085 125.670 36.280 126.000 ;
        RECT 36.505 125.670 36.760 126.000 ;
        RECT 36.505 125.500 36.675 125.670 ;
        RECT 36.930 125.500 37.100 126.170 ;
        RECT 38.195 126.145 38.485 127.310 ;
        RECT 38.655 126.220 40.325 127.310 ;
        RECT 40.695 126.640 40.975 127.310 ;
        RECT 41.145 126.420 41.445 126.970 ;
        RECT 41.645 126.590 41.975 127.310 ;
        RECT 42.165 126.590 42.625 127.140 ;
        RECT 38.655 125.700 39.405 126.220 ;
        RECT 39.575 125.530 40.325 126.050 ;
        RECT 40.510 126.000 40.775 126.360 ;
        RECT 41.145 126.250 42.085 126.420 ;
        RECT 41.915 126.000 42.085 126.250 ;
        RECT 40.510 125.750 41.185 126.000 ;
        RECT 41.405 125.750 41.745 126.000 ;
        RECT 41.915 125.670 42.205 126.000 ;
        RECT 41.915 125.580 42.085 125.670 ;
        RECT 35.745 125.330 36.675 125.500 ;
        RECT 35.745 125.295 35.920 125.330 ;
        RECT 35.390 124.930 35.920 125.295 ;
        RECT 36.345 124.760 36.675 125.160 ;
        RECT 36.845 124.930 37.100 125.500 ;
        RECT 38.195 124.760 38.485 125.485 ;
        RECT 38.655 124.760 40.325 125.530 ;
        RECT 40.695 125.390 42.085 125.580 ;
        RECT 40.695 125.030 41.025 125.390 ;
        RECT 42.375 125.220 42.625 126.590 ;
        RECT 43.755 126.170 43.985 127.310 ;
        RECT 44.155 126.160 44.485 127.140 ;
        RECT 44.655 126.170 44.865 127.310 ;
        RECT 45.100 126.875 50.445 127.310 ;
        RECT 50.990 126.970 51.245 127.000 ;
        RECT 43.735 125.750 44.065 126.000 ;
        RECT 41.645 124.760 41.895 125.220 ;
        RECT 42.065 124.930 42.625 125.220 ;
        RECT 43.755 124.760 43.985 125.580 ;
        RECT 44.235 125.560 44.485 126.160 ;
        RECT 46.690 125.625 47.040 126.875 ;
        RECT 50.905 126.800 51.245 126.970 ;
        RECT 50.990 126.330 51.245 126.800 ;
        RECT 51.425 126.510 51.710 127.310 ;
        RECT 51.890 126.590 52.220 127.100 ;
        RECT 44.155 124.930 44.485 125.560 ;
        RECT 44.655 124.760 44.865 125.580 ;
        RECT 48.520 125.305 48.860 126.135 ;
        RECT 50.990 125.470 51.170 126.330 ;
        RECT 51.890 126.000 52.140 126.590 ;
        RECT 52.490 126.440 52.660 127.050 ;
        RECT 52.830 126.620 53.160 127.310 ;
        RECT 53.390 126.760 53.630 127.050 ;
        RECT 53.830 126.930 54.250 127.310 ;
        RECT 54.430 126.840 55.060 127.090 ;
        RECT 55.530 126.930 55.860 127.310 ;
        RECT 54.430 126.760 54.600 126.840 ;
        RECT 56.030 126.760 56.200 127.050 ;
        RECT 56.380 126.930 56.760 127.310 ;
        RECT 57.000 126.925 57.830 127.095 ;
        RECT 53.390 126.590 54.600 126.760 ;
        RECT 51.340 125.670 52.140 126.000 ;
        RECT 45.100 124.760 50.445 125.305 ;
        RECT 50.990 124.940 51.245 125.470 ;
        RECT 51.425 124.760 51.710 125.220 ;
        RECT 51.890 125.020 52.140 125.670 ;
        RECT 52.340 126.420 52.660 126.440 ;
        RECT 52.340 126.250 54.260 126.420 ;
        RECT 52.340 125.355 52.530 126.250 ;
        RECT 54.430 126.080 54.600 126.590 ;
        RECT 54.770 126.330 55.290 126.640 ;
        RECT 52.700 125.910 54.600 126.080 ;
        RECT 52.700 125.850 53.030 125.910 ;
        RECT 53.180 125.680 53.510 125.740 ;
        RECT 52.850 125.410 53.510 125.680 ;
        RECT 52.340 125.025 52.660 125.355 ;
        RECT 52.840 124.760 53.500 125.240 ;
        RECT 53.700 125.150 53.870 125.910 ;
        RECT 54.770 125.740 54.950 126.150 ;
        RECT 54.040 125.570 54.370 125.690 ;
        RECT 55.120 125.570 55.290 126.330 ;
        RECT 54.040 125.400 55.290 125.570 ;
        RECT 55.460 126.510 56.830 126.760 ;
        RECT 55.460 125.740 55.650 126.510 ;
        RECT 56.580 126.250 56.830 126.510 ;
        RECT 55.820 126.080 56.070 126.240 ;
        RECT 57.000 126.080 57.170 126.925 ;
        RECT 58.065 126.640 58.235 127.140 ;
        RECT 58.405 126.810 58.735 127.310 ;
        RECT 57.340 126.250 57.840 126.630 ;
        RECT 58.065 126.470 58.760 126.640 ;
        RECT 55.820 125.910 57.170 126.080 ;
        RECT 56.750 125.870 57.170 125.910 ;
        RECT 55.460 125.400 55.880 125.740 ;
        RECT 56.170 125.410 56.580 125.740 ;
        RECT 53.700 124.980 54.550 125.150 ;
        RECT 55.110 124.760 55.430 125.220 ;
        RECT 55.630 124.970 55.880 125.400 ;
        RECT 56.170 124.760 56.580 125.200 ;
        RECT 56.750 125.140 56.920 125.870 ;
        RECT 57.090 125.320 57.440 125.690 ;
        RECT 57.620 125.380 57.840 126.250 ;
        RECT 58.010 125.680 58.420 126.300 ;
        RECT 58.590 125.500 58.760 126.470 ;
        RECT 58.065 125.310 58.760 125.500 ;
        RECT 56.750 124.940 57.765 125.140 ;
        RECT 58.065 124.980 58.235 125.310 ;
        RECT 58.405 124.760 58.735 125.140 ;
        RECT 58.950 125.020 59.175 127.140 ;
        RECT 59.345 126.810 59.675 127.310 ;
        RECT 59.845 126.640 60.015 127.140 ;
        RECT 59.350 126.470 60.015 126.640 ;
        RECT 59.350 125.480 59.580 126.470 ;
        RECT 59.750 125.650 60.100 126.300 ;
        RECT 60.275 126.220 63.785 127.310 ;
        RECT 60.275 125.700 61.965 126.220 ;
        RECT 63.955 126.145 64.245 127.310 ;
        RECT 64.875 126.220 68.385 127.310 ;
        RECT 68.555 126.550 69.070 126.960 ;
        RECT 69.305 126.550 69.475 127.310 ;
        RECT 69.645 126.970 71.675 127.140 ;
        RECT 62.135 125.530 63.785 126.050 ;
        RECT 64.875 125.700 66.565 126.220 ;
        RECT 66.735 125.530 68.385 126.050 ;
        RECT 68.555 125.740 68.895 126.550 ;
        RECT 69.645 126.305 69.815 126.970 ;
        RECT 70.210 126.630 71.335 126.800 ;
        RECT 69.065 126.115 69.815 126.305 ;
        RECT 69.985 126.290 70.995 126.460 ;
        RECT 68.555 125.570 69.785 125.740 ;
        RECT 59.350 125.310 60.015 125.480 ;
        RECT 59.345 124.760 59.675 125.140 ;
        RECT 59.845 125.020 60.015 125.310 ;
        RECT 60.275 124.760 63.785 125.530 ;
        RECT 63.955 124.760 64.245 125.485 ;
        RECT 64.875 124.760 68.385 125.530 ;
        RECT 68.830 124.965 69.075 125.570 ;
        RECT 69.295 124.760 69.805 125.295 ;
        RECT 69.985 124.930 70.175 126.290 ;
        RECT 70.345 125.270 70.620 126.090 ;
        RECT 70.825 125.490 70.995 126.290 ;
        RECT 71.165 125.500 71.335 126.630 ;
        RECT 71.505 126.000 71.675 126.970 ;
        RECT 71.845 126.170 72.015 127.310 ;
        RECT 72.185 126.170 72.520 127.140 ;
        RECT 71.505 125.670 71.700 126.000 ;
        RECT 71.925 125.670 72.180 126.000 ;
        RECT 71.925 125.500 72.095 125.670 ;
        RECT 72.350 125.500 72.520 126.170 ;
        RECT 72.695 126.220 74.365 127.310 ;
        RECT 72.695 125.700 73.445 126.220 ;
        RECT 74.595 126.170 74.805 127.310 ;
        RECT 74.975 126.160 75.305 127.140 ;
        RECT 75.475 126.170 75.705 127.310 ;
        RECT 76.375 126.220 78.045 127.310 ;
        RECT 78.275 126.475 78.530 127.310 ;
        RECT 78.700 126.305 78.960 127.110 ;
        RECT 79.130 126.475 79.390 127.310 ;
        RECT 79.560 126.305 79.815 127.110 ;
        RECT 80.145 126.640 80.315 127.140 ;
        RECT 80.485 126.810 80.815 127.310 ;
        RECT 80.145 126.470 80.810 126.640 ;
        RECT 73.615 125.530 74.365 126.050 ;
        RECT 71.165 125.330 72.095 125.500 ;
        RECT 71.165 125.295 71.340 125.330 ;
        RECT 70.345 125.100 70.625 125.270 ;
        RECT 70.345 124.930 70.620 125.100 ;
        RECT 70.810 124.930 71.340 125.295 ;
        RECT 71.765 124.760 72.095 125.160 ;
        RECT 72.265 124.930 72.520 125.500 ;
        RECT 72.695 124.760 74.365 125.530 ;
        RECT 74.595 124.760 74.805 125.580 ;
        RECT 74.975 125.560 75.225 126.160 ;
        RECT 75.395 125.750 75.725 126.000 ;
        RECT 76.375 125.700 77.125 126.220 ;
        RECT 78.215 126.135 79.815 126.305 ;
        RECT 74.975 124.930 75.305 125.560 ;
        RECT 75.475 124.760 75.705 125.580 ;
        RECT 77.295 125.530 78.045 126.050 ;
        RECT 76.375 124.760 78.045 125.530 ;
        RECT 78.215 125.570 78.495 126.135 ;
        RECT 78.665 125.740 79.885 125.965 ;
        RECT 80.060 125.650 80.410 126.300 ;
        RECT 78.215 125.400 78.945 125.570 ;
        RECT 80.580 125.480 80.810 126.470 ;
        RECT 78.220 124.760 78.550 125.230 ;
        RECT 78.720 124.955 78.945 125.400 ;
        RECT 80.145 125.310 80.810 125.480 ;
        RECT 79.115 124.760 79.410 125.285 ;
        RECT 80.145 125.020 80.315 125.310 ;
        RECT 80.485 124.760 80.815 125.140 ;
        RECT 80.985 125.020 81.210 127.140 ;
        RECT 81.425 126.810 81.755 127.310 ;
        RECT 81.925 126.640 82.095 127.140 ;
        RECT 82.330 126.925 83.160 127.095 ;
        RECT 83.400 126.930 83.780 127.310 ;
        RECT 81.400 126.470 82.095 126.640 ;
        RECT 81.400 125.500 81.570 126.470 ;
        RECT 81.740 125.680 82.150 126.300 ;
        RECT 82.320 126.250 82.820 126.630 ;
        RECT 81.400 125.310 82.095 125.500 ;
        RECT 82.320 125.380 82.540 126.250 ;
        RECT 82.990 126.080 83.160 126.925 ;
        RECT 83.960 126.760 84.130 127.050 ;
        RECT 84.300 126.930 84.630 127.310 ;
        RECT 85.100 126.840 85.730 127.090 ;
        RECT 85.910 126.930 86.330 127.310 ;
        RECT 85.560 126.760 85.730 126.840 ;
        RECT 86.530 126.760 86.770 127.050 ;
        RECT 83.330 126.510 84.700 126.760 ;
        RECT 83.330 126.250 83.580 126.510 ;
        RECT 84.090 126.080 84.340 126.240 ;
        RECT 82.990 125.910 84.340 126.080 ;
        RECT 82.990 125.870 83.410 125.910 ;
        RECT 82.720 125.320 83.070 125.690 ;
        RECT 81.425 124.760 81.755 125.140 ;
        RECT 81.925 124.980 82.095 125.310 ;
        RECT 83.240 125.140 83.410 125.870 ;
        RECT 84.510 125.740 84.700 126.510 ;
        RECT 83.580 125.410 83.990 125.740 ;
        RECT 84.280 125.400 84.700 125.740 ;
        RECT 84.870 126.330 85.390 126.640 ;
        RECT 85.560 126.590 86.770 126.760 ;
        RECT 87.000 126.620 87.330 127.310 ;
        RECT 84.870 125.570 85.040 126.330 ;
        RECT 85.210 125.740 85.390 126.150 ;
        RECT 85.560 126.080 85.730 126.590 ;
        RECT 87.500 126.440 87.670 127.050 ;
        RECT 87.940 126.590 88.270 127.100 ;
        RECT 87.500 126.420 87.820 126.440 ;
        RECT 85.900 126.250 87.820 126.420 ;
        RECT 85.560 125.910 87.460 126.080 ;
        RECT 85.790 125.570 86.120 125.690 ;
        RECT 84.870 125.400 86.120 125.570 ;
        RECT 82.395 124.940 83.410 125.140 ;
        RECT 83.580 124.760 83.990 125.200 ;
        RECT 84.280 124.970 84.530 125.400 ;
        RECT 84.730 124.760 85.050 125.220 ;
        RECT 86.290 125.150 86.460 125.910 ;
        RECT 87.130 125.850 87.460 125.910 ;
        RECT 86.650 125.680 86.980 125.740 ;
        RECT 86.650 125.410 87.310 125.680 ;
        RECT 87.630 125.355 87.820 126.250 ;
        RECT 85.610 124.980 86.460 125.150 ;
        RECT 86.660 124.760 87.320 125.240 ;
        RECT 87.500 125.025 87.820 125.355 ;
        RECT 88.020 126.000 88.270 126.590 ;
        RECT 88.450 126.510 88.735 127.310 ;
        RECT 88.915 126.970 89.170 127.000 ;
        RECT 88.915 126.800 89.255 126.970 ;
        RECT 88.915 126.330 89.170 126.800 ;
        RECT 88.020 125.670 88.820 126.000 ;
        RECT 88.020 125.020 88.270 125.670 ;
        RECT 88.990 125.470 89.170 126.330 ;
        RECT 89.715 126.145 90.005 127.310 ;
        RECT 90.635 126.220 92.305 127.310 ;
        RECT 90.635 125.700 91.385 126.220 ;
        RECT 92.515 126.170 92.745 127.310 ;
        RECT 92.915 126.160 93.245 127.140 ;
        RECT 93.415 126.170 93.625 127.310 ;
        RECT 93.855 126.550 94.370 126.960 ;
        RECT 94.605 126.550 94.775 127.310 ;
        RECT 94.945 126.970 96.975 127.140 ;
        RECT 91.555 125.530 92.305 126.050 ;
        RECT 92.495 125.750 92.825 126.000 ;
        RECT 88.450 124.760 88.735 125.220 ;
        RECT 88.915 124.940 89.170 125.470 ;
        RECT 89.715 124.760 90.005 125.485 ;
        RECT 90.635 124.760 92.305 125.530 ;
        RECT 92.515 124.760 92.745 125.580 ;
        RECT 92.995 125.560 93.245 126.160 ;
        RECT 93.855 125.740 94.195 126.550 ;
        RECT 94.945 126.305 95.115 126.970 ;
        RECT 95.510 126.630 96.635 126.800 ;
        RECT 94.365 126.115 95.115 126.305 ;
        RECT 95.285 126.290 96.295 126.460 ;
        RECT 92.915 124.930 93.245 125.560 ;
        RECT 93.415 124.760 93.625 125.580 ;
        RECT 93.855 125.570 95.085 125.740 ;
        RECT 94.130 124.965 94.375 125.570 ;
        RECT 94.595 124.760 95.105 125.295 ;
        RECT 95.285 124.930 95.475 126.290 ;
        RECT 95.645 125.610 95.920 126.090 ;
        RECT 95.645 125.440 95.925 125.610 ;
        RECT 96.125 125.490 96.295 126.290 ;
        RECT 96.465 125.500 96.635 126.630 ;
        RECT 96.805 126.000 96.975 126.970 ;
        RECT 97.145 126.170 97.315 127.310 ;
        RECT 97.485 126.170 97.820 127.140 ;
        RECT 96.805 125.670 97.000 126.000 ;
        RECT 97.225 125.670 97.480 126.000 ;
        RECT 97.225 125.500 97.395 125.670 ;
        RECT 97.650 125.500 97.820 126.170 ;
        RECT 97.995 126.220 99.665 127.310 ;
        RECT 99.835 126.550 100.350 126.960 ;
        RECT 100.585 126.550 100.755 127.310 ;
        RECT 100.925 126.970 102.955 127.140 ;
        RECT 97.995 125.700 98.745 126.220 ;
        RECT 98.915 125.530 99.665 126.050 ;
        RECT 99.835 125.740 100.175 126.550 ;
        RECT 100.925 126.305 101.095 126.970 ;
        RECT 101.490 126.630 102.615 126.800 ;
        RECT 100.345 126.115 101.095 126.305 ;
        RECT 101.265 126.290 102.275 126.460 ;
        RECT 99.835 125.570 101.065 125.740 ;
        RECT 95.645 124.930 95.920 125.440 ;
        RECT 96.465 125.330 97.395 125.500 ;
        RECT 96.465 125.295 96.640 125.330 ;
        RECT 96.110 124.930 96.640 125.295 ;
        RECT 97.065 124.760 97.395 125.160 ;
        RECT 97.565 124.930 97.820 125.500 ;
        RECT 97.995 124.760 99.665 125.530 ;
        RECT 100.110 124.965 100.355 125.570 ;
        RECT 100.575 124.760 101.085 125.295 ;
        RECT 101.265 124.930 101.455 126.290 ;
        RECT 101.625 125.950 101.900 126.090 ;
        RECT 101.625 125.780 101.905 125.950 ;
        RECT 101.625 124.930 101.900 125.780 ;
        RECT 102.105 125.490 102.275 126.290 ;
        RECT 102.445 125.500 102.615 126.630 ;
        RECT 102.785 126.000 102.955 126.970 ;
        RECT 103.125 126.170 103.295 127.310 ;
        RECT 103.465 126.170 103.800 127.140 ;
        RECT 102.785 125.670 102.980 126.000 ;
        RECT 103.205 125.670 103.460 126.000 ;
        RECT 103.205 125.500 103.375 125.670 ;
        RECT 103.630 125.500 103.800 126.170 ;
        RECT 104.350 126.330 104.605 127.000 ;
        RECT 104.785 126.510 105.070 127.310 ;
        RECT 105.250 126.590 105.580 127.100 ;
        RECT 104.350 125.950 104.530 126.330 ;
        RECT 105.250 126.000 105.500 126.590 ;
        RECT 105.850 126.440 106.020 127.050 ;
        RECT 106.190 126.620 106.520 127.310 ;
        RECT 106.750 126.760 106.990 127.050 ;
        RECT 107.190 126.930 107.610 127.310 ;
        RECT 107.790 126.840 108.420 127.090 ;
        RECT 108.890 126.930 109.220 127.310 ;
        RECT 107.790 126.760 107.960 126.840 ;
        RECT 109.390 126.760 109.560 127.050 ;
        RECT 109.740 126.930 110.120 127.310 ;
        RECT 110.360 126.925 111.190 127.095 ;
        RECT 106.750 126.590 107.960 126.760 ;
        RECT 104.265 125.780 104.530 125.950 ;
        RECT 102.445 125.330 103.375 125.500 ;
        RECT 102.445 125.295 102.620 125.330 ;
        RECT 102.090 124.930 102.620 125.295 ;
        RECT 103.045 124.760 103.375 125.160 ;
        RECT 103.545 124.930 103.800 125.500 ;
        RECT 104.350 125.470 104.530 125.780 ;
        RECT 104.700 125.670 105.500 126.000 ;
        RECT 104.350 124.940 104.605 125.470 ;
        RECT 104.785 124.760 105.070 125.220 ;
        RECT 105.250 125.020 105.500 125.670 ;
        RECT 105.700 126.420 106.020 126.440 ;
        RECT 105.700 126.250 107.620 126.420 ;
        RECT 105.700 125.355 105.890 126.250 ;
        RECT 107.790 126.080 107.960 126.590 ;
        RECT 108.130 126.330 108.650 126.640 ;
        RECT 106.060 125.910 107.960 126.080 ;
        RECT 106.060 125.850 106.390 125.910 ;
        RECT 106.540 125.680 106.870 125.740 ;
        RECT 106.210 125.410 106.870 125.680 ;
        RECT 105.700 125.025 106.020 125.355 ;
        RECT 106.200 124.760 106.860 125.240 ;
        RECT 107.060 125.150 107.230 125.910 ;
        RECT 108.130 125.740 108.310 126.150 ;
        RECT 107.400 125.570 107.730 125.690 ;
        RECT 108.480 125.570 108.650 126.330 ;
        RECT 107.400 125.400 108.650 125.570 ;
        RECT 108.820 126.510 110.190 126.760 ;
        RECT 108.820 125.740 109.010 126.510 ;
        RECT 109.940 126.250 110.190 126.510 ;
        RECT 109.180 126.080 109.430 126.240 ;
        RECT 110.360 126.080 110.530 126.925 ;
        RECT 111.425 126.640 111.595 127.140 ;
        RECT 111.765 126.810 112.095 127.310 ;
        RECT 110.700 126.250 111.200 126.630 ;
        RECT 111.425 126.470 112.120 126.640 ;
        RECT 109.180 125.910 110.530 126.080 ;
        RECT 110.110 125.870 110.530 125.910 ;
        RECT 108.820 125.400 109.240 125.740 ;
        RECT 109.530 125.410 109.940 125.740 ;
        RECT 107.060 124.980 107.910 125.150 ;
        RECT 108.470 124.760 108.790 125.220 ;
        RECT 108.990 124.970 109.240 125.400 ;
        RECT 109.530 124.760 109.940 125.200 ;
        RECT 110.110 125.140 110.280 125.870 ;
        RECT 110.450 125.320 110.800 125.690 ;
        RECT 110.980 125.380 111.200 126.250 ;
        RECT 111.370 125.680 111.780 126.300 ;
        RECT 111.950 125.500 112.120 126.470 ;
        RECT 111.425 125.310 112.120 125.500 ;
        RECT 110.110 124.940 111.125 125.140 ;
        RECT 111.425 124.980 111.595 125.310 ;
        RECT 111.765 124.760 112.095 125.140 ;
        RECT 112.310 125.020 112.535 127.140 ;
        RECT 112.705 126.810 113.035 127.310 ;
        RECT 113.205 126.640 113.375 127.140 ;
        RECT 112.710 126.470 113.375 126.640 ;
        RECT 112.710 125.480 112.940 126.470 ;
        RECT 113.110 125.650 113.460 126.300 ;
        RECT 114.555 126.220 115.765 127.310 ;
        RECT 114.555 125.680 115.075 126.220 ;
        RECT 115.245 125.510 115.765 126.050 ;
        RECT 112.710 125.310 113.375 125.480 ;
        RECT 112.705 124.760 113.035 125.140 ;
        RECT 113.205 125.020 113.375 125.310 ;
        RECT 114.555 124.760 115.765 125.510 ;
        RECT 10.510 124.590 115.850 124.760 ;
        RECT 10.595 123.840 11.805 124.590 ;
        RECT 11.975 123.840 13.185 124.590 ;
        RECT 10.595 123.300 11.115 123.840 ;
        RECT 11.285 123.130 11.805 123.670 ;
        RECT 10.595 122.040 11.805 123.130 ;
        RECT 11.975 123.130 12.495 123.670 ;
        RECT 12.665 123.300 13.185 123.840 ;
        RECT 13.415 123.770 13.625 124.590 ;
        RECT 13.795 123.790 14.125 124.420 ;
        RECT 13.795 123.190 14.045 123.790 ;
        RECT 14.295 123.770 14.525 124.590 ;
        RECT 14.735 123.915 14.995 124.420 ;
        RECT 15.175 124.210 15.505 124.590 ;
        RECT 15.685 124.040 15.855 124.420 ;
        RECT 16.205 124.110 16.505 124.590 ;
        RECT 14.215 123.350 14.545 123.600 ;
        RECT 11.975 122.040 13.185 123.130 ;
        RECT 13.415 122.040 13.625 123.180 ;
        RECT 13.795 122.210 14.125 123.190 ;
        RECT 14.295 122.040 14.525 123.180 ;
        RECT 14.735 123.115 14.905 123.915 ;
        RECT 15.190 123.870 15.855 124.040 ;
        RECT 16.675 123.940 16.935 124.395 ;
        RECT 17.105 124.110 17.365 124.590 ;
        RECT 17.545 123.940 17.805 124.395 ;
        RECT 17.975 124.110 18.225 124.590 ;
        RECT 18.405 123.940 18.665 124.395 ;
        RECT 18.835 124.110 19.085 124.590 ;
        RECT 19.265 123.940 19.525 124.395 ;
        RECT 19.695 124.110 19.940 124.590 ;
        RECT 20.110 123.940 20.385 124.395 ;
        RECT 20.555 124.110 20.800 124.590 ;
        RECT 20.970 123.940 21.230 124.395 ;
        RECT 21.400 124.110 21.660 124.590 ;
        RECT 21.830 123.940 22.090 124.395 ;
        RECT 22.260 124.110 22.520 124.590 ;
        RECT 22.690 123.940 22.950 124.395 ;
        RECT 23.120 124.030 23.380 124.590 ;
        RECT 15.190 123.615 15.360 123.870 ;
        RECT 16.205 123.770 22.950 123.940 ;
        RECT 15.075 123.285 15.360 123.615 ;
        RECT 15.595 123.320 15.925 123.690 ;
        RECT 15.190 123.140 15.360 123.285 ;
        RECT 16.205 123.180 17.370 123.770 ;
        RECT 23.550 123.600 23.800 124.410 ;
        RECT 23.980 124.065 24.240 124.590 ;
        RECT 24.410 123.600 24.660 124.410 ;
        RECT 24.840 124.080 25.145 124.590 ;
        RECT 17.540 123.350 24.660 123.600 ;
        RECT 24.830 123.350 25.145 123.910 ;
        RECT 25.315 123.865 25.605 124.590 ;
        RECT 26.970 123.780 27.215 124.385 ;
        RECT 27.435 124.055 27.945 124.590 ;
        RECT 26.695 123.610 27.925 123.780 ;
        RECT 14.735 122.210 15.005 123.115 ;
        RECT 15.190 122.970 15.855 123.140 ;
        RECT 15.175 122.040 15.505 122.800 ;
        RECT 15.685 122.210 15.855 122.970 ;
        RECT 16.205 122.955 22.950 123.180 ;
        RECT 16.205 122.040 16.475 122.785 ;
        RECT 16.645 122.215 16.935 122.955 ;
        RECT 17.545 122.940 22.950 122.955 ;
        RECT 17.105 122.045 17.360 122.770 ;
        RECT 17.545 122.215 17.805 122.940 ;
        RECT 17.975 122.045 18.220 122.770 ;
        RECT 18.405 122.215 18.665 122.940 ;
        RECT 18.835 122.045 19.080 122.770 ;
        RECT 19.265 122.215 19.525 122.940 ;
        RECT 19.695 122.045 19.940 122.770 ;
        RECT 20.110 122.215 20.370 122.940 ;
        RECT 20.540 122.045 20.800 122.770 ;
        RECT 20.970 122.215 21.230 122.940 ;
        RECT 21.400 122.045 21.660 122.770 ;
        RECT 21.830 122.215 22.090 122.940 ;
        RECT 22.260 122.045 22.520 122.770 ;
        RECT 22.690 122.215 22.950 122.940 ;
        RECT 23.120 122.045 23.380 122.840 ;
        RECT 23.550 122.215 23.800 123.350 ;
        RECT 17.105 122.040 23.380 122.045 ;
        RECT 23.980 122.040 24.240 122.850 ;
        RECT 24.415 122.210 24.660 123.350 ;
        RECT 24.840 122.040 25.135 122.850 ;
        RECT 25.315 122.040 25.605 123.205 ;
        RECT 26.695 122.800 27.035 123.610 ;
        RECT 27.205 123.045 27.955 123.235 ;
        RECT 26.695 122.390 27.210 122.800 ;
        RECT 27.445 122.040 27.615 122.800 ;
        RECT 27.785 122.380 27.955 123.045 ;
        RECT 28.125 123.060 28.315 124.420 ;
        RECT 28.485 123.570 28.760 124.420 ;
        RECT 28.950 124.055 29.480 124.420 ;
        RECT 29.905 124.190 30.235 124.590 ;
        RECT 29.305 124.020 29.480 124.055 ;
        RECT 28.485 123.400 28.765 123.570 ;
        RECT 28.485 123.260 28.760 123.400 ;
        RECT 28.965 123.060 29.135 123.860 ;
        RECT 28.125 122.890 29.135 123.060 ;
        RECT 29.305 123.850 30.235 124.020 ;
        RECT 30.405 123.850 30.660 124.420 ;
        RECT 29.305 122.720 29.475 123.850 ;
        RECT 30.065 123.680 30.235 123.850 ;
        RECT 28.350 122.550 29.475 122.720 ;
        RECT 29.645 123.350 29.840 123.680 ;
        RECT 30.065 123.350 30.320 123.680 ;
        RECT 29.645 122.380 29.815 123.350 ;
        RECT 30.490 123.180 30.660 123.850 ;
        RECT 31.210 123.880 31.465 124.410 ;
        RECT 31.645 124.130 31.930 124.590 ;
        RECT 31.210 123.570 31.390 123.880 ;
        RECT 32.110 123.680 32.360 124.330 ;
        RECT 31.125 123.400 31.390 123.570 ;
        RECT 27.785 122.210 29.815 122.380 ;
        RECT 29.985 122.040 30.155 123.180 ;
        RECT 30.325 122.210 30.660 123.180 ;
        RECT 31.210 123.020 31.390 123.400 ;
        RECT 31.560 123.350 32.360 123.680 ;
        RECT 31.210 122.350 31.465 123.020 ;
        RECT 31.645 122.040 31.930 122.840 ;
        RECT 32.110 122.760 32.360 123.350 ;
        RECT 32.560 123.995 32.880 124.325 ;
        RECT 33.060 124.110 33.720 124.590 ;
        RECT 33.920 124.200 34.770 124.370 ;
        RECT 32.560 123.100 32.750 123.995 ;
        RECT 33.070 123.670 33.730 123.940 ;
        RECT 33.400 123.610 33.730 123.670 ;
        RECT 32.920 123.440 33.250 123.500 ;
        RECT 33.920 123.440 34.090 124.200 ;
        RECT 35.330 124.130 35.650 124.590 ;
        RECT 35.850 123.950 36.100 124.380 ;
        RECT 36.390 124.150 36.800 124.590 ;
        RECT 36.970 124.210 37.985 124.410 ;
        RECT 34.260 123.780 35.510 123.950 ;
        RECT 34.260 123.660 34.590 123.780 ;
        RECT 32.920 123.270 34.820 123.440 ;
        RECT 32.560 122.930 34.480 123.100 ;
        RECT 32.560 122.910 32.880 122.930 ;
        RECT 32.110 122.250 32.440 122.760 ;
        RECT 32.710 122.300 32.880 122.910 ;
        RECT 34.650 122.760 34.820 123.270 ;
        RECT 34.990 123.200 35.170 123.610 ;
        RECT 35.340 123.020 35.510 123.780 ;
        RECT 33.050 122.040 33.380 122.730 ;
        RECT 33.610 122.590 34.820 122.760 ;
        RECT 34.990 122.710 35.510 123.020 ;
        RECT 35.680 123.610 36.100 123.950 ;
        RECT 36.390 123.610 36.800 123.940 ;
        RECT 35.680 122.840 35.870 123.610 ;
        RECT 36.970 123.480 37.140 124.210 ;
        RECT 38.285 124.040 38.455 124.370 ;
        RECT 38.625 124.210 38.955 124.590 ;
        RECT 37.310 123.660 37.660 124.030 ;
        RECT 36.970 123.440 37.390 123.480 ;
        RECT 36.040 123.270 37.390 123.440 ;
        RECT 36.040 123.110 36.290 123.270 ;
        RECT 36.800 122.840 37.050 123.100 ;
        RECT 35.680 122.590 37.050 122.840 ;
        RECT 33.610 122.300 33.850 122.590 ;
        RECT 34.650 122.510 34.820 122.590 ;
        RECT 34.050 122.040 34.470 122.420 ;
        RECT 34.650 122.260 35.280 122.510 ;
        RECT 35.750 122.040 36.080 122.420 ;
        RECT 36.250 122.300 36.420 122.590 ;
        RECT 37.220 122.425 37.390 123.270 ;
        RECT 37.840 123.100 38.060 123.970 ;
        RECT 38.285 123.850 38.980 124.040 ;
        RECT 37.560 122.720 38.060 123.100 ;
        RECT 38.230 123.050 38.640 123.670 ;
        RECT 38.810 122.880 38.980 123.850 ;
        RECT 38.285 122.710 38.980 122.880 ;
        RECT 36.600 122.040 36.980 122.420 ;
        RECT 37.220 122.255 38.050 122.425 ;
        RECT 38.285 122.210 38.455 122.710 ;
        RECT 38.625 122.040 38.955 122.540 ;
        RECT 39.170 122.210 39.395 124.330 ;
        RECT 39.565 124.210 39.895 124.590 ;
        RECT 40.065 124.040 40.235 124.330 ;
        RECT 39.570 123.870 40.235 124.040 ;
        RECT 40.870 123.880 41.125 124.410 ;
        RECT 41.305 124.130 41.590 124.590 ;
        RECT 39.570 122.880 39.800 123.870 ;
        RECT 39.970 123.050 40.320 123.700 ;
        RECT 40.870 123.020 41.050 123.880 ;
        RECT 41.770 123.680 42.020 124.330 ;
        RECT 41.220 123.350 42.020 123.680 ;
        RECT 39.570 122.710 40.235 122.880 ;
        RECT 39.565 122.040 39.895 122.540 ;
        RECT 40.065 122.210 40.235 122.710 ;
        RECT 40.870 122.550 41.125 123.020 ;
        RECT 40.785 122.380 41.125 122.550 ;
        RECT 40.870 122.350 41.125 122.380 ;
        RECT 41.305 122.040 41.590 122.840 ;
        RECT 41.770 122.760 42.020 123.350 ;
        RECT 42.220 123.995 42.540 124.325 ;
        RECT 42.720 124.110 43.380 124.590 ;
        RECT 43.580 124.200 44.430 124.370 ;
        RECT 42.220 123.100 42.410 123.995 ;
        RECT 42.730 123.670 43.390 123.940 ;
        RECT 43.060 123.610 43.390 123.670 ;
        RECT 42.580 123.440 42.910 123.500 ;
        RECT 43.580 123.440 43.750 124.200 ;
        RECT 44.990 124.130 45.310 124.590 ;
        RECT 45.510 123.950 45.760 124.380 ;
        RECT 46.050 124.150 46.460 124.590 ;
        RECT 46.630 124.210 47.645 124.410 ;
        RECT 43.920 123.780 45.170 123.950 ;
        RECT 43.920 123.660 44.250 123.780 ;
        RECT 42.580 123.270 44.480 123.440 ;
        RECT 42.220 122.930 44.140 123.100 ;
        RECT 42.220 122.910 42.540 122.930 ;
        RECT 41.770 122.250 42.100 122.760 ;
        RECT 42.370 122.300 42.540 122.910 ;
        RECT 44.310 122.760 44.480 123.270 ;
        RECT 44.650 123.200 44.830 123.610 ;
        RECT 45.000 123.020 45.170 123.780 ;
        RECT 42.710 122.040 43.040 122.730 ;
        RECT 43.270 122.590 44.480 122.760 ;
        RECT 44.650 122.710 45.170 123.020 ;
        RECT 45.340 123.610 45.760 123.950 ;
        RECT 46.050 123.610 46.460 123.940 ;
        RECT 45.340 122.840 45.530 123.610 ;
        RECT 46.630 123.480 46.800 124.210 ;
        RECT 47.945 124.040 48.115 124.370 ;
        RECT 48.285 124.210 48.615 124.590 ;
        RECT 46.970 123.660 47.320 124.030 ;
        RECT 46.630 123.440 47.050 123.480 ;
        RECT 45.700 123.270 47.050 123.440 ;
        RECT 45.700 123.110 45.950 123.270 ;
        RECT 46.460 122.840 46.710 123.100 ;
        RECT 45.340 122.590 46.710 122.840 ;
        RECT 43.270 122.300 43.510 122.590 ;
        RECT 44.310 122.510 44.480 122.590 ;
        RECT 43.710 122.040 44.130 122.420 ;
        RECT 44.310 122.260 44.940 122.510 ;
        RECT 45.410 122.040 45.740 122.420 ;
        RECT 45.910 122.300 46.080 122.590 ;
        RECT 46.880 122.425 47.050 123.270 ;
        RECT 47.500 123.100 47.720 123.970 ;
        RECT 47.945 123.850 48.640 124.040 ;
        RECT 47.220 122.720 47.720 123.100 ;
        RECT 47.890 123.050 48.300 123.670 ;
        RECT 48.470 122.880 48.640 123.850 ;
        RECT 47.945 122.710 48.640 122.880 ;
        RECT 46.260 122.040 46.640 122.420 ;
        RECT 46.880 122.255 47.710 122.425 ;
        RECT 47.945 122.210 48.115 122.710 ;
        RECT 48.285 122.040 48.615 122.540 ;
        RECT 48.830 122.210 49.055 124.330 ;
        RECT 49.225 124.210 49.555 124.590 ;
        RECT 49.725 124.040 49.895 124.330 ;
        RECT 49.230 123.870 49.895 124.040 ;
        RECT 49.230 122.880 49.460 123.870 ;
        RECT 51.075 123.865 51.365 124.590 ;
        RECT 51.625 124.040 51.795 124.420 ;
        RECT 51.975 124.210 52.305 124.590 ;
        RECT 51.625 123.870 52.290 124.040 ;
        RECT 52.485 123.915 52.745 124.420 ;
        RECT 49.630 123.050 49.980 123.700 ;
        RECT 51.555 123.320 51.885 123.690 ;
        RECT 52.120 123.615 52.290 123.870 ;
        RECT 52.120 123.285 52.405 123.615 ;
        RECT 49.230 122.710 49.895 122.880 ;
        RECT 49.225 122.040 49.555 122.540 ;
        RECT 49.725 122.210 49.895 122.710 ;
        RECT 51.075 122.040 51.365 123.205 ;
        RECT 52.120 123.140 52.290 123.285 ;
        RECT 51.625 122.970 52.290 123.140 ;
        RECT 52.575 123.115 52.745 123.915 ;
        RECT 51.625 122.210 51.795 122.970 ;
        RECT 51.975 122.040 52.305 122.800 ;
        RECT 52.475 122.210 52.745 123.115 ;
        RECT 53.840 123.850 54.095 124.420 ;
        RECT 54.265 124.190 54.595 124.590 ;
        RECT 55.020 124.055 55.550 124.420 ;
        RECT 55.740 124.250 56.015 124.420 ;
        RECT 55.735 124.080 56.015 124.250 ;
        RECT 55.020 124.020 55.195 124.055 ;
        RECT 54.265 123.850 55.195 124.020 ;
        RECT 53.840 123.180 54.010 123.850 ;
        RECT 54.265 123.680 54.435 123.850 ;
        RECT 54.180 123.350 54.435 123.680 ;
        RECT 54.660 123.350 54.855 123.680 ;
        RECT 53.840 122.210 54.175 123.180 ;
        RECT 54.345 122.040 54.515 123.180 ;
        RECT 54.685 122.380 54.855 123.350 ;
        RECT 55.025 122.720 55.195 123.850 ;
        RECT 55.365 123.060 55.535 123.860 ;
        RECT 55.740 123.260 56.015 124.080 ;
        RECT 56.185 123.060 56.375 124.420 ;
        RECT 56.555 124.055 57.065 124.590 ;
        RECT 57.285 123.780 57.530 124.385 ;
        RECT 58.250 123.780 58.495 124.385 ;
        RECT 58.715 124.055 59.225 124.590 ;
        RECT 56.575 123.610 57.805 123.780 ;
        RECT 55.365 122.890 56.375 123.060 ;
        RECT 56.545 123.045 57.295 123.235 ;
        RECT 55.025 122.550 56.150 122.720 ;
        RECT 56.545 122.380 56.715 123.045 ;
        RECT 57.465 122.800 57.805 123.610 ;
        RECT 54.685 122.210 56.715 122.380 ;
        RECT 56.885 122.040 57.055 122.800 ;
        RECT 57.290 122.390 57.805 122.800 ;
        RECT 57.975 123.610 59.205 123.780 ;
        RECT 57.975 122.800 58.315 123.610 ;
        RECT 58.485 123.045 59.235 123.235 ;
        RECT 57.975 122.390 58.490 122.800 ;
        RECT 58.725 122.040 58.895 122.800 ;
        RECT 59.065 122.380 59.235 123.045 ;
        RECT 59.405 123.060 59.595 124.420 ;
        RECT 59.765 123.570 60.040 124.420 ;
        RECT 60.230 124.055 60.760 124.420 ;
        RECT 61.185 124.190 61.515 124.590 ;
        RECT 60.585 124.020 60.760 124.055 ;
        RECT 59.765 123.400 60.045 123.570 ;
        RECT 59.765 123.260 60.040 123.400 ;
        RECT 60.245 123.060 60.415 123.860 ;
        RECT 59.405 122.890 60.415 123.060 ;
        RECT 60.585 123.850 61.515 124.020 ;
        RECT 61.685 123.850 61.940 124.420 ;
        RECT 60.585 122.720 60.755 123.850 ;
        RECT 61.345 123.680 61.515 123.850 ;
        RECT 59.630 122.550 60.755 122.720 ;
        RECT 60.925 123.350 61.120 123.680 ;
        RECT 61.345 123.350 61.600 123.680 ;
        RECT 60.925 122.380 61.095 123.350 ;
        RECT 61.770 123.180 61.940 123.850 ;
        RECT 62.115 123.820 65.625 124.590 ;
        RECT 66.170 124.250 66.425 124.410 ;
        RECT 66.085 124.080 66.425 124.250 ;
        RECT 66.605 124.130 66.890 124.590 ;
        RECT 59.065 122.210 61.095 122.380 ;
        RECT 61.265 122.040 61.435 123.180 ;
        RECT 61.605 122.210 61.940 123.180 ;
        RECT 62.115 123.130 63.805 123.650 ;
        RECT 63.975 123.300 65.625 123.820 ;
        RECT 66.170 123.880 66.425 124.080 ;
        RECT 62.115 122.040 65.625 123.130 ;
        RECT 66.170 123.020 66.350 123.880 ;
        RECT 67.070 123.680 67.320 124.330 ;
        RECT 66.520 123.350 67.320 123.680 ;
        RECT 66.170 122.350 66.425 123.020 ;
        RECT 66.605 122.040 66.890 122.840 ;
        RECT 67.070 122.760 67.320 123.350 ;
        RECT 67.520 123.995 67.840 124.325 ;
        RECT 68.020 124.110 68.680 124.590 ;
        RECT 68.880 124.200 69.730 124.370 ;
        RECT 67.520 123.100 67.710 123.995 ;
        RECT 68.030 123.670 68.690 123.940 ;
        RECT 68.360 123.610 68.690 123.670 ;
        RECT 67.880 123.440 68.210 123.500 ;
        RECT 68.880 123.440 69.050 124.200 ;
        RECT 70.290 124.130 70.610 124.590 ;
        RECT 70.810 123.950 71.060 124.380 ;
        RECT 71.350 124.150 71.760 124.590 ;
        RECT 71.930 124.210 72.945 124.410 ;
        RECT 69.220 123.780 70.470 123.950 ;
        RECT 69.220 123.660 69.550 123.780 ;
        RECT 67.880 123.270 69.780 123.440 ;
        RECT 67.520 122.930 69.440 123.100 ;
        RECT 67.520 122.910 67.840 122.930 ;
        RECT 67.070 122.250 67.400 122.760 ;
        RECT 67.670 122.300 67.840 122.910 ;
        RECT 69.610 122.760 69.780 123.270 ;
        RECT 69.950 123.200 70.130 123.610 ;
        RECT 70.300 123.020 70.470 123.780 ;
        RECT 68.010 122.040 68.340 122.730 ;
        RECT 68.570 122.590 69.780 122.760 ;
        RECT 69.950 122.710 70.470 123.020 ;
        RECT 70.640 123.610 71.060 123.950 ;
        RECT 71.350 123.610 71.760 123.940 ;
        RECT 70.640 122.840 70.830 123.610 ;
        RECT 71.930 123.480 72.100 124.210 ;
        RECT 73.245 124.040 73.415 124.370 ;
        RECT 73.585 124.210 73.915 124.590 ;
        RECT 72.270 123.660 72.620 124.030 ;
        RECT 71.930 123.440 72.350 123.480 ;
        RECT 71.000 123.270 72.350 123.440 ;
        RECT 71.000 123.110 71.250 123.270 ;
        RECT 71.760 122.840 72.010 123.100 ;
        RECT 70.640 122.590 72.010 122.840 ;
        RECT 68.570 122.300 68.810 122.590 ;
        RECT 69.610 122.510 69.780 122.590 ;
        RECT 69.010 122.040 69.430 122.420 ;
        RECT 69.610 122.260 70.240 122.510 ;
        RECT 70.710 122.040 71.040 122.420 ;
        RECT 71.210 122.300 71.380 122.590 ;
        RECT 72.180 122.425 72.350 123.270 ;
        RECT 72.800 123.100 73.020 123.970 ;
        RECT 73.245 123.850 73.940 124.040 ;
        RECT 72.520 122.720 73.020 123.100 ;
        RECT 73.190 123.050 73.600 123.670 ;
        RECT 73.770 122.880 73.940 123.850 ;
        RECT 73.245 122.710 73.940 122.880 ;
        RECT 71.560 122.040 71.940 122.420 ;
        RECT 72.180 122.255 73.010 122.425 ;
        RECT 73.245 122.210 73.415 122.710 ;
        RECT 73.585 122.040 73.915 122.540 ;
        RECT 74.130 122.210 74.355 124.330 ;
        RECT 74.525 124.210 74.855 124.590 ;
        RECT 75.025 124.040 75.195 124.330 ;
        RECT 74.530 123.870 75.195 124.040 ;
        RECT 75.455 123.915 75.715 124.420 ;
        RECT 75.895 124.210 76.225 124.590 ;
        RECT 76.405 124.040 76.575 124.420 ;
        RECT 74.530 122.880 74.760 123.870 ;
        RECT 74.930 123.050 75.280 123.700 ;
        RECT 75.455 123.115 75.625 123.915 ;
        RECT 75.910 123.870 76.575 124.040 ;
        RECT 75.910 123.615 76.080 123.870 ;
        RECT 76.835 123.865 77.125 124.590 ;
        RECT 77.385 124.110 77.685 124.590 ;
        RECT 77.855 123.940 78.115 124.395 ;
        RECT 78.285 124.110 78.545 124.590 ;
        RECT 78.725 123.940 78.985 124.395 ;
        RECT 79.155 124.110 79.405 124.590 ;
        RECT 79.585 123.940 79.845 124.395 ;
        RECT 80.015 124.110 80.265 124.590 ;
        RECT 80.445 123.940 80.705 124.395 ;
        RECT 80.875 124.110 81.120 124.590 ;
        RECT 81.290 123.940 81.565 124.395 ;
        RECT 81.735 124.110 81.980 124.590 ;
        RECT 82.150 123.940 82.410 124.395 ;
        RECT 82.580 124.110 82.840 124.590 ;
        RECT 83.010 123.940 83.270 124.395 ;
        RECT 83.440 124.110 83.700 124.590 ;
        RECT 83.870 123.940 84.130 124.395 ;
        RECT 84.300 124.030 84.560 124.590 ;
        RECT 77.385 123.770 84.130 123.940 ;
        RECT 75.795 123.285 76.080 123.615 ;
        RECT 76.315 123.320 76.645 123.690 ;
        RECT 75.910 123.140 76.080 123.285 ;
        RECT 74.530 122.710 75.195 122.880 ;
        RECT 74.525 122.040 74.855 122.540 ;
        RECT 75.025 122.210 75.195 122.710 ;
        RECT 75.455 122.210 75.725 123.115 ;
        RECT 75.910 122.970 76.575 123.140 ;
        RECT 75.895 122.040 76.225 122.800 ;
        RECT 76.405 122.210 76.575 122.970 ;
        RECT 76.835 122.040 77.125 123.205 ;
        RECT 77.385 123.180 78.550 123.770 ;
        RECT 84.730 123.600 84.980 124.410 ;
        RECT 85.160 124.065 85.420 124.590 ;
        RECT 85.590 123.600 85.840 124.410 ;
        RECT 86.020 124.080 86.325 124.590 ;
        RECT 78.720 123.350 85.840 123.600 ;
        RECT 86.010 123.350 86.325 123.910 ;
        RECT 87.230 123.780 87.475 124.385 ;
        RECT 87.695 124.055 88.205 124.590 ;
        RECT 86.955 123.610 88.185 123.780 ;
        RECT 77.385 122.955 84.130 123.180 ;
        RECT 77.385 122.040 77.655 122.785 ;
        RECT 77.825 122.215 78.115 122.955 ;
        RECT 78.725 122.940 84.130 122.955 ;
        RECT 78.285 122.045 78.540 122.770 ;
        RECT 78.725 122.215 78.985 122.940 ;
        RECT 79.155 122.045 79.400 122.770 ;
        RECT 79.585 122.215 79.845 122.940 ;
        RECT 80.015 122.045 80.260 122.770 ;
        RECT 80.445 122.215 80.705 122.940 ;
        RECT 80.875 122.045 81.120 122.770 ;
        RECT 81.290 122.215 81.550 122.940 ;
        RECT 81.720 122.045 81.980 122.770 ;
        RECT 82.150 122.215 82.410 122.940 ;
        RECT 82.580 122.045 82.840 122.770 ;
        RECT 83.010 122.215 83.270 122.940 ;
        RECT 83.440 122.045 83.700 122.770 ;
        RECT 83.870 122.215 84.130 122.940 ;
        RECT 84.300 122.045 84.560 122.840 ;
        RECT 84.730 122.215 84.980 123.350 ;
        RECT 78.285 122.040 84.560 122.045 ;
        RECT 85.160 122.040 85.420 122.850 ;
        RECT 85.595 122.210 85.840 123.350 ;
        RECT 86.020 122.040 86.315 122.850 ;
        RECT 86.955 122.800 87.295 123.610 ;
        RECT 87.465 123.045 88.215 123.235 ;
        RECT 86.955 122.390 87.470 122.800 ;
        RECT 87.705 122.040 87.875 122.800 ;
        RECT 88.045 122.380 88.215 123.045 ;
        RECT 88.385 123.060 88.575 124.420 ;
        RECT 88.745 123.570 89.020 124.420 ;
        RECT 89.210 124.055 89.740 124.420 ;
        RECT 90.165 124.190 90.495 124.590 ;
        RECT 89.565 124.020 89.740 124.055 ;
        RECT 88.745 123.400 89.025 123.570 ;
        RECT 88.745 123.260 89.020 123.400 ;
        RECT 89.225 123.060 89.395 123.860 ;
        RECT 88.385 122.890 89.395 123.060 ;
        RECT 89.565 123.850 90.495 124.020 ;
        RECT 90.665 123.850 90.920 124.420 ;
        RECT 89.565 122.720 89.735 123.850 ;
        RECT 90.325 123.680 90.495 123.850 ;
        RECT 88.610 122.550 89.735 122.720 ;
        RECT 89.905 123.350 90.100 123.680 ;
        RECT 90.325 123.350 90.580 123.680 ;
        RECT 89.905 122.380 90.075 123.350 ;
        RECT 90.750 123.180 90.920 123.850 ;
        RECT 91.155 123.770 91.365 124.590 ;
        RECT 91.535 123.790 91.865 124.420 ;
        RECT 91.535 123.190 91.785 123.790 ;
        RECT 92.035 123.770 92.265 124.590 ;
        RECT 93.395 124.080 93.700 124.590 ;
        RECT 91.955 123.350 92.285 123.600 ;
        RECT 93.395 123.350 93.710 123.910 ;
        RECT 93.880 123.600 94.130 124.410 ;
        RECT 94.300 124.065 94.560 124.590 ;
        RECT 94.740 123.600 94.990 124.410 ;
        RECT 95.160 124.030 95.420 124.590 ;
        RECT 95.590 123.940 95.850 124.395 ;
        RECT 96.020 124.110 96.280 124.590 ;
        RECT 96.450 123.940 96.710 124.395 ;
        RECT 96.880 124.110 97.140 124.590 ;
        RECT 97.310 123.940 97.570 124.395 ;
        RECT 97.740 124.110 97.985 124.590 ;
        RECT 98.155 123.940 98.430 124.395 ;
        RECT 98.600 124.110 98.845 124.590 ;
        RECT 99.015 123.940 99.275 124.395 ;
        RECT 99.455 124.110 99.705 124.590 ;
        RECT 99.875 123.940 100.135 124.395 ;
        RECT 100.315 124.110 100.565 124.590 ;
        RECT 100.735 123.940 100.995 124.395 ;
        RECT 101.175 124.110 101.435 124.590 ;
        RECT 101.605 123.940 101.865 124.395 ;
        RECT 102.035 124.110 102.335 124.590 ;
        RECT 95.590 123.770 102.335 123.940 ;
        RECT 102.595 123.865 102.885 124.590 ;
        RECT 103.890 123.880 104.145 124.410 ;
        RECT 104.325 124.130 104.610 124.590 ;
        RECT 93.880 123.350 101.000 123.600 ;
        RECT 88.045 122.210 90.075 122.380 ;
        RECT 90.245 122.040 90.415 123.180 ;
        RECT 90.585 122.210 90.920 123.180 ;
        RECT 91.155 122.040 91.365 123.180 ;
        RECT 91.535 122.210 91.865 123.190 ;
        RECT 92.035 122.040 92.265 123.180 ;
        RECT 93.405 122.040 93.700 122.850 ;
        RECT 93.880 122.210 94.125 123.350 ;
        RECT 94.300 122.040 94.560 122.850 ;
        RECT 94.740 122.215 94.990 123.350 ;
        RECT 101.170 123.180 102.335 123.770 ;
        RECT 95.590 122.955 102.335 123.180 ;
        RECT 95.590 122.940 100.995 122.955 ;
        RECT 95.160 122.045 95.420 122.840 ;
        RECT 95.590 122.215 95.850 122.940 ;
        RECT 96.020 122.045 96.280 122.770 ;
        RECT 96.450 122.215 96.710 122.940 ;
        RECT 96.880 122.045 97.140 122.770 ;
        RECT 97.310 122.215 97.570 122.940 ;
        RECT 97.740 122.045 98.000 122.770 ;
        RECT 98.170 122.215 98.430 122.940 ;
        RECT 98.600 122.045 98.845 122.770 ;
        RECT 99.015 122.215 99.275 122.940 ;
        RECT 99.460 122.045 99.705 122.770 ;
        RECT 99.875 122.215 100.135 122.940 ;
        RECT 100.320 122.045 100.565 122.770 ;
        RECT 100.735 122.215 100.995 122.940 ;
        RECT 101.180 122.045 101.435 122.770 ;
        RECT 101.605 122.215 101.895 122.955 ;
        RECT 95.160 122.040 101.435 122.045 ;
        RECT 102.065 122.040 102.335 122.785 ;
        RECT 102.595 122.040 102.885 123.205 ;
        RECT 103.890 123.020 104.070 123.880 ;
        RECT 104.790 123.680 105.040 124.330 ;
        RECT 104.240 123.350 105.040 123.680 ;
        RECT 103.890 122.550 104.145 123.020 ;
        RECT 103.805 122.380 104.145 122.550 ;
        RECT 103.890 122.350 104.145 122.380 ;
        RECT 104.325 122.040 104.610 122.840 ;
        RECT 104.790 122.760 105.040 123.350 ;
        RECT 105.240 123.995 105.560 124.325 ;
        RECT 105.740 124.110 106.400 124.590 ;
        RECT 106.600 124.200 107.450 124.370 ;
        RECT 105.240 123.100 105.430 123.995 ;
        RECT 105.750 123.670 106.410 123.940 ;
        RECT 106.080 123.610 106.410 123.670 ;
        RECT 105.600 123.440 105.930 123.500 ;
        RECT 106.600 123.440 106.770 124.200 ;
        RECT 108.010 124.130 108.330 124.590 ;
        RECT 108.530 123.950 108.780 124.380 ;
        RECT 109.070 124.150 109.480 124.590 ;
        RECT 109.650 124.210 110.665 124.410 ;
        RECT 106.940 123.780 108.190 123.950 ;
        RECT 106.940 123.660 107.270 123.780 ;
        RECT 105.600 123.270 107.500 123.440 ;
        RECT 105.240 122.930 107.160 123.100 ;
        RECT 105.240 122.910 105.560 122.930 ;
        RECT 104.790 122.250 105.120 122.760 ;
        RECT 105.390 122.300 105.560 122.910 ;
        RECT 107.330 122.760 107.500 123.270 ;
        RECT 107.670 123.200 107.850 123.610 ;
        RECT 108.020 123.020 108.190 123.780 ;
        RECT 105.730 122.040 106.060 122.730 ;
        RECT 106.290 122.590 107.500 122.760 ;
        RECT 107.670 122.710 108.190 123.020 ;
        RECT 108.360 123.610 108.780 123.950 ;
        RECT 109.070 123.610 109.480 123.940 ;
        RECT 108.360 122.840 108.550 123.610 ;
        RECT 109.650 123.480 109.820 124.210 ;
        RECT 110.965 124.040 111.135 124.370 ;
        RECT 111.305 124.210 111.635 124.590 ;
        RECT 109.990 123.660 110.340 124.030 ;
        RECT 109.650 123.440 110.070 123.480 ;
        RECT 108.720 123.270 110.070 123.440 ;
        RECT 108.720 123.110 108.970 123.270 ;
        RECT 109.480 122.840 109.730 123.100 ;
        RECT 108.360 122.590 109.730 122.840 ;
        RECT 106.290 122.300 106.530 122.590 ;
        RECT 107.330 122.510 107.500 122.590 ;
        RECT 106.730 122.040 107.150 122.420 ;
        RECT 107.330 122.260 107.960 122.510 ;
        RECT 108.430 122.040 108.760 122.420 ;
        RECT 108.930 122.300 109.100 122.590 ;
        RECT 109.900 122.425 110.070 123.270 ;
        RECT 110.520 123.100 110.740 123.970 ;
        RECT 110.965 123.850 111.660 124.040 ;
        RECT 110.240 122.720 110.740 123.100 ;
        RECT 110.910 123.050 111.320 123.670 ;
        RECT 111.490 122.880 111.660 123.850 ;
        RECT 110.965 122.710 111.660 122.880 ;
        RECT 109.280 122.040 109.660 122.420 ;
        RECT 109.900 122.255 110.730 122.425 ;
        RECT 110.965 122.210 111.135 122.710 ;
        RECT 111.305 122.040 111.635 122.540 ;
        RECT 111.850 122.210 112.075 124.330 ;
        RECT 112.245 124.210 112.575 124.590 ;
        RECT 112.745 124.040 112.915 124.330 ;
        RECT 112.250 123.870 112.915 124.040 ;
        RECT 113.175 123.915 113.435 124.420 ;
        RECT 113.615 124.210 113.945 124.590 ;
        RECT 114.125 124.040 114.295 124.420 ;
        RECT 112.250 122.880 112.480 123.870 ;
        RECT 112.650 123.050 113.000 123.700 ;
        RECT 113.175 123.115 113.345 123.915 ;
        RECT 113.630 123.870 114.295 124.040 ;
        RECT 113.630 123.615 113.800 123.870 ;
        RECT 114.555 123.840 115.765 124.590 ;
        RECT 113.515 123.285 113.800 123.615 ;
        RECT 114.035 123.320 114.365 123.690 ;
        RECT 113.630 123.140 113.800 123.285 ;
        RECT 112.250 122.710 112.915 122.880 ;
        RECT 112.245 122.040 112.575 122.540 ;
        RECT 112.745 122.210 112.915 122.710 ;
        RECT 113.175 122.210 113.445 123.115 ;
        RECT 113.630 122.970 114.295 123.140 ;
        RECT 113.615 122.040 113.945 122.800 ;
        RECT 114.125 122.210 114.295 122.970 ;
        RECT 114.555 123.130 115.075 123.670 ;
        RECT 115.245 123.300 115.765 123.840 ;
        RECT 114.555 122.040 115.765 123.130 ;
        RECT 10.510 121.870 115.850 122.040 ;
        RECT 10.595 120.780 11.805 121.870 ;
        RECT 10.595 120.070 11.115 120.610 ;
        RECT 11.285 120.240 11.805 120.780 ;
        RECT 12.435 120.705 12.725 121.870 ;
        RECT 13.445 121.200 13.615 121.700 ;
        RECT 13.785 121.370 14.115 121.870 ;
        RECT 13.445 121.030 14.110 121.200 ;
        RECT 13.360 120.210 13.710 120.860 ;
        RECT 10.595 119.320 11.805 120.070 ;
        RECT 12.435 119.320 12.725 120.045 ;
        RECT 13.880 120.040 14.110 121.030 ;
        RECT 13.445 119.870 14.110 120.040 ;
        RECT 13.445 119.580 13.615 119.870 ;
        RECT 13.785 119.320 14.115 119.700 ;
        RECT 14.285 119.580 14.510 121.700 ;
        RECT 14.725 121.370 15.055 121.870 ;
        RECT 15.225 121.200 15.395 121.700 ;
        RECT 15.630 121.485 16.460 121.655 ;
        RECT 16.700 121.490 17.080 121.870 ;
        RECT 14.700 121.030 15.395 121.200 ;
        RECT 14.700 120.060 14.870 121.030 ;
        RECT 15.040 120.240 15.450 120.860 ;
        RECT 15.620 120.810 16.120 121.190 ;
        RECT 14.700 119.870 15.395 120.060 ;
        RECT 15.620 119.940 15.840 120.810 ;
        RECT 16.290 120.640 16.460 121.485 ;
        RECT 17.260 121.320 17.430 121.610 ;
        RECT 17.600 121.490 17.930 121.870 ;
        RECT 18.400 121.400 19.030 121.650 ;
        RECT 19.210 121.490 19.630 121.870 ;
        RECT 18.860 121.320 19.030 121.400 ;
        RECT 19.830 121.320 20.070 121.610 ;
        RECT 16.630 121.070 18.000 121.320 ;
        RECT 16.630 120.810 16.880 121.070 ;
        RECT 17.390 120.640 17.640 120.800 ;
        RECT 16.290 120.470 17.640 120.640 ;
        RECT 16.290 120.430 16.710 120.470 ;
        RECT 16.020 119.880 16.370 120.250 ;
        RECT 14.725 119.320 15.055 119.700 ;
        RECT 15.225 119.540 15.395 119.870 ;
        RECT 16.540 119.700 16.710 120.430 ;
        RECT 17.810 120.300 18.000 121.070 ;
        RECT 16.880 119.970 17.290 120.300 ;
        RECT 17.580 119.960 18.000 120.300 ;
        RECT 18.170 120.890 18.690 121.200 ;
        RECT 18.860 121.150 20.070 121.320 ;
        RECT 20.300 121.180 20.630 121.870 ;
        RECT 18.170 120.130 18.340 120.890 ;
        RECT 18.510 120.300 18.690 120.710 ;
        RECT 18.860 120.640 19.030 121.150 ;
        RECT 20.800 121.000 20.970 121.610 ;
        RECT 21.240 121.150 21.570 121.660 ;
        RECT 20.800 120.980 21.120 121.000 ;
        RECT 19.200 120.810 21.120 120.980 ;
        RECT 18.860 120.470 20.760 120.640 ;
        RECT 19.090 120.130 19.420 120.250 ;
        RECT 18.170 119.960 19.420 120.130 ;
        RECT 15.695 119.500 16.710 119.700 ;
        RECT 16.880 119.320 17.290 119.760 ;
        RECT 17.580 119.530 17.830 119.960 ;
        RECT 18.030 119.320 18.350 119.780 ;
        RECT 19.590 119.710 19.760 120.470 ;
        RECT 20.430 120.410 20.760 120.470 ;
        RECT 19.950 120.240 20.280 120.300 ;
        RECT 19.950 119.970 20.610 120.240 ;
        RECT 20.930 119.915 21.120 120.810 ;
        RECT 18.910 119.540 19.760 119.710 ;
        RECT 19.960 119.320 20.620 119.800 ;
        RECT 20.800 119.585 21.120 119.915 ;
        RECT 21.320 120.560 21.570 121.150 ;
        RECT 21.750 121.070 22.035 121.870 ;
        RECT 22.215 121.190 22.470 121.560 ;
        RECT 22.215 121.020 22.555 121.190 ;
        RECT 22.215 120.890 22.470 121.020 ;
        RECT 21.320 120.230 22.120 120.560 ;
        RECT 21.320 119.580 21.570 120.230 ;
        RECT 22.290 120.030 22.470 120.890 ;
        RECT 21.750 119.320 22.035 119.780 ;
        RECT 22.215 119.500 22.470 120.030 ;
        RECT 23.020 120.730 23.355 121.700 ;
        RECT 23.525 120.730 23.695 121.870 ;
        RECT 23.865 121.530 25.895 121.700 ;
        RECT 23.020 120.060 23.190 120.730 ;
        RECT 23.865 120.560 24.035 121.530 ;
        RECT 23.360 120.230 23.615 120.560 ;
        RECT 23.840 120.230 24.035 120.560 ;
        RECT 24.205 121.190 25.330 121.360 ;
        RECT 23.445 120.060 23.615 120.230 ;
        RECT 24.205 120.060 24.375 121.190 ;
        RECT 23.020 119.490 23.275 120.060 ;
        RECT 23.445 119.890 24.375 120.060 ;
        RECT 24.545 120.850 25.555 121.020 ;
        RECT 24.545 120.050 24.715 120.850 ;
        RECT 24.200 119.855 24.375 119.890 ;
        RECT 23.445 119.320 23.775 119.720 ;
        RECT 24.200 119.490 24.730 119.855 ;
        RECT 24.920 119.830 25.195 120.650 ;
        RECT 24.915 119.660 25.195 119.830 ;
        RECT 24.920 119.490 25.195 119.660 ;
        RECT 25.365 119.490 25.555 120.850 ;
        RECT 25.725 120.865 25.895 121.530 ;
        RECT 26.065 121.110 26.235 121.870 ;
        RECT 27.990 121.530 28.245 121.560 ;
        RECT 26.470 121.110 26.985 121.520 ;
        RECT 27.905 121.360 28.245 121.530 ;
        RECT 25.725 120.675 26.475 120.865 ;
        RECT 26.645 120.300 26.985 121.110 ;
        RECT 25.755 120.130 26.985 120.300 ;
        RECT 27.990 120.890 28.245 121.360 ;
        RECT 28.425 121.070 28.710 121.870 ;
        RECT 28.890 121.150 29.220 121.660 ;
        RECT 25.735 119.320 26.245 119.855 ;
        RECT 26.465 119.525 26.710 120.130 ;
        RECT 27.990 120.030 28.170 120.890 ;
        RECT 28.890 120.560 29.140 121.150 ;
        RECT 29.490 121.000 29.660 121.610 ;
        RECT 29.830 121.180 30.160 121.870 ;
        RECT 30.390 121.320 30.630 121.610 ;
        RECT 30.830 121.490 31.250 121.870 ;
        RECT 31.430 121.400 32.060 121.650 ;
        RECT 32.530 121.490 32.860 121.870 ;
        RECT 31.430 121.320 31.600 121.400 ;
        RECT 33.030 121.320 33.200 121.610 ;
        RECT 33.380 121.490 33.760 121.870 ;
        RECT 34.000 121.485 34.830 121.655 ;
        RECT 30.390 121.150 31.600 121.320 ;
        RECT 28.340 120.230 29.140 120.560 ;
        RECT 27.990 119.500 28.245 120.030 ;
        RECT 28.425 119.320 28.710 119.780 ;
        RECT 28.890 119.580 29.140 120.230 ;
        RECT 29.340 120.980 29.660 121.000 ;
        RECT 29.340 120.810 31.260 120.980 ;
        RECT 29.340 119.915 29.530 120.810 ;
        RECT 31.430 120.640 31.600 121.150 ;
        RECT 31.770 120.890 32.290 121.200 ;
        RECT 29.700 120.470 31.600 120.640 ;
        RECT 29.700 120.410 30.030 120.470 ;
        RECT 30.180 120.240 30.510 120.300 ;
        RECT 29.850 119.970 30.510 120.240 ;
        RECT 29.340 119.585 29.660 119.915 ;
        RECT 29.840 119.320 30.500 119.800 ;
        RECT 30.700 119.710 30.870 120.470 ;
        RECT 31.770 120.300 31.950 120.710 ;
        RECT 31.040 120.130 31.370 120.250 ;
        RECT 32.120 120.130 32.290 120.890 ;
        RECT 31.040 119.960 32.290 120.130 ;
        RECT 32.460 121.070 33.830 121.320 ;
        RECT 32.460 120.300 32.650 121.070 ;
        RECT 33.580 120.810 33.830 121.070 ;
        RECT 32.820 120.640 33.070 120.800 ;
        RECT 34.000 120.640 34.170 121.485 ;
        RECT 35.065 121.200 35.235 121.700 ;
        RECT 35.405 121.370 35.735 121.870 ;
        RECT 34.340 120.810 34.840 121.190 ;
        RECT 35.065 121.030 35.760 121.200 ;
        RECT 32.820 120.470 34.170 120.640 ;
        RECT 33.750 120.430 34.170 120.470 ;
        RECT 32.460 119.960 32.880 120.300 ;
        RECT 33.170 119.970 33.580 120.300 ;
        RECT 30.700 119.540 31.550 119.710 ;
        RECT 32.110 119.320 32.430 119.780 ;
        RECT 32.630 119.530 32.880 119.960 ;
        RECT 33.170 119.320 33.580 119.760 ;
        RECT 33.750 119.700 33.920 120.430 ;
        RECT 34.090 119.880 34.440 120.250 ;
        RECT 34.620 119.940 34.840 120.810 ;
        RECT 35.010 120.240 35.420 120.860 ;
        RECT 35.590 120.060 35.760 121.030 ;
        RECT 35.065 119.870 35.760 120.060 ;
        RECT 33.750 119.500 34.765 119.700 ;
        RECT 35.065 119.540 35.235 119.870 ;
        RECT 35.405 119.320 35.735 119.700 ;
        RECT 35.950 119.580 36.175 121.700 ;
        RECT 36.345 121.370 36.675 121.870 ;
        RECT 36.845 121.200 37.015 121.700 ;
        RECT 36.350 121.030 37.015 121.200 ;
        RECT 36.350 120.040 36.580 121.030 ;
        RECT 36.750 120.210 37.100 120.860 ;
        RECT 38.195 120.705 38.485 121.870 ;
        RECT 39.115 120.795 39.385 121.700 ;
        RECT 39.555 121.110 39.885 121.870 ;
        RECT 40.065 120.940 40.235 121.700 ;
        RECT 36.350 119.870 37.015 120.040 ;
        RECT 36.345 119.320 36.675 119.700 ;
        RECT 36.845 119.580 37.015 119.870 ;
        RECT 38.195 119.320 38.485 120.045 ;
        RECT 39.115 119.995 39.285 120.795 ;
        RECT 39.570 120.770 40.235 120.940 ;
        RECT 40.495 120.780 41.705 121.870 ;
        RECT 41.985 121.070 42.155 121.870 ;
        RECT 42.325 120.850 42.655 121.700 ;
        RECT 42.825 121.070 42.995 121.870 ;
        RECT 43.165 120.850 43.495 121.700 ;
        RECT 43.665 121.070 43.835 121.870 ;
        RECT 44.005 120.850 44.335 121.700 ;
        RECT 44.505 121.070 44.675 121.870 ;
        RECT 44.845 120.850 45.175 121.700 ;
        RECT 45.345 121.070 45.515 121.870 ;
        RECT 45.685 120.850 46.015 121.700 ;
        RECT 46.185 121.070 46.355 121.870 ;
        RECT 46.525 120.850 46.855 121.700 ;
        RECT 47.025 121.070 47.195 121.870 ;
        RECT 47.365 120.850 47.695 121.700 ;
        RECT 47.865 121.070 48.035 121.870 ;
        RECT 48.205 120.850 48.535 121.700 ;
        RECT 48.705 121.070 48.875 121.870 ;
        RECT 49.045 120.850 49.375 121.700 ;
        RECT 49.545 121.070 49.715 121.870 ;
        RECT 49.885 120.850 50.215 121.700 ;
        RECT 50.385 121.070 50.555 121.870 ;
        RECT 50.725 120.850 51.055 121.700 ;
        RECT 51.225 121.020 51.395 121.870 ;
        RECT 51.565 120.850 51.895 121.700 ;
        RECT 52.065 121.020 52.235 121.870 ;
        RECT 52.405 120.850 52.735 121.700 ;
        RECT 39.570 120.625 39.740 120.770 ;
        RECT 39.455 120.295 39.740 120.625 ;
        RECT 39.570 120.040 39.740 120.295 ;
        RECT 39.975 120.220 40.305 120.590 ;
        RECT 40.495 120.240 41.015 120.780 ;
        RECT 41.875 120.680 48.535 120.850 ;
        RECT 48.705 120.680 51.055 120.850 ;
        RECT 51.225 120.680 52.735 120.850 ;
        RECT 52.955 120.730 53.185 121.870 ;
        RECT 53.355 120.720 53.685 121.700 ;
        RECT 53.855 120.730 54.065 121.870 ;
        RECT 54.670 121.530 54.925 121.560 ;
        RECT 54.585 121.360 54.925 121.530 ;
        RECT 54.670 120.890 54.925 121.360 ;
        RECT 55.105 121.070 55.390 121.870 ;
        RECT 55.570 121.150 55.900 121.660 ;
        RECT 41.185 120.070 41.705 120.610 ;
        RECT 39.115 119.490 39.375 119.995 ;
        RECT 39.570 119.870 40.235 120.040 ;
        RECT 39.555 119.320 39.885 119.700 ;
        RECT 40.065 119.490 40.235 119.870 ;
        RECT 40.495 119.320 41.705 120.070 ;
        RECT 41.875 120.140 42.150 120.680 ;
        RECT 48.705 120.510 48.880 120.680 ;
        RECT 51.225 120.510 51.395 120.680 ;
        RECT 42.320 120.310 48.880 120.510 ;
        RECT 49.085 120.310 51.395 120.510 ;
        RECT 51.565 120.310 52.740 120.510 ;
        RECT 52.935 120.310 53.265 120.560 ;
        RECT 48.705 120.140 48.880 120.310 ;
        RECT 51.225 120.140 51.395 120.310 ;
        RECT 41.875 119.970 48.535 120.140 ;
        RECT 48.705 119.970 51.055 120.140 ;
        RECT 51.225 119.970 52.735 120.140 ;
        RECT 41.985 119.320 42.155 119.800 ;
        RECT 42.325 119.495 42.655 119.970 ;
        RECT 42.825 119.320 42.995 119.800 ;
        RECT 43.165 119.495 43.495 119.970 ;
        RECT 43.665 119.320 43.835 119.800 ;
        RECT 44.005 119.495 44.335 119.970 ;
        RECT 44.505 119.320 44.675 119.800 ;
        RECT 44.845 119.495 45.175 119.970 ;
        RECT 45.345 119.320 45.515 119.800 ;
        RECT 45.685 119.495 46.015 119.970 ;
        RECT 46.185 119.320 46.355 119.800 ;
        RECT 46.525 119.495 46.855 119.970 ;
        RECT 46.605 119.490 46.775 119.495 ;
        RECT 47.025 119.320 47.195 119.800 ;
        RECT 47.365 119.495 47.695 119.970 ;
        RECT 47.445 119.490 47.615 119.495 ;
        RECT 47.865 119.320 48.035 119.800 ;
        RECT 48.205 119.495 48.535 119.970 ;
        RECT 48.285 119.490 48.535 119.495 ;
        RECT 48.705 119.320 48.875 119.800 ;
        RECT 49.045 119.495 49.375 119.970 ;
        RECT 49.545 119.320 49.715 119.800 ;
        RECT 49.885 119.495 50.215 119.970 ;
        RECT 50.385 119.320 50.555 119.800 ;
        RECT 50.725 119.495 51.055 119.970 ;
        RECT 51.225 119.320 51.395 119.800 ;
        RECT 51.565 119.495 51.895 119.970 ;
        RECT 52.065 119.320 52.235 119.800 ;
        RECT 52.405 119.495 52.735 119.970 ;
        RECT 52.955 119.320 53.185 120.140 ;
        RECT 53.435 120.120 53.685 120.720 ;
        RECT 53.355 119.490 53.685 120.120 ;
        RECT 53.855 119.320 54.065 120.140 ;
        RECT 54.670 120.030 54.850 120.890 ;
        RECT 55.570 120.560 55.820 121.150 ;
        RECT 56.170 121.000 56.340 121.610 ;
        RECT 56.510 121.180 56.840 121.870 ;
        RECT 57.070 121.320 57.310 121.610 ;
        RECT 57.510 121.490 57.930 121.870 ;
        RECT 58.110 121.400 58.740 121.650 ;
        RECT 59.210 121.490 59.540 121.870 ;
        RECT 58.110 121.320 58.280 121.400 ;
        RECT 59.710 121.320 59.880 121.610 ;
        RECT 60.060 121.490 60.440 121.870 ;
        RECT 60.680 121.485 61.510 121.655 ;
        RECT 57.070 121.150 58.280 121.320 ;
        RECT 55.020 120.230 55.820 120.560 ;
        RECT 54.670 119.500 54.925 120.030 ;
        RECT 55.105 119.320 55.390 119.780 ;
        RECT 55.570 119.580 55.820 120.230 ;
        RECT 56.020 120.980 56.340 121.000 ;
        RECT 56.020 120.810 57.940 120.980 ;
        RECT 56.020 119.915 56.210 120.810 ;
        RECT 58.110 120.640 58.280 121.150 ;
        RECT 58.450 120.890 58.970 121.200 ;
        RECT 56.380 120.470 58.280 120.640 ;
        RECT 56.380 120.410 56.710 120.470 ;
        RECT 56.860 120.240 57.190 120.300 ;
        RECT 56.530 119.970 57.190 120.240 ;
        RECT 56.020 119.585 56.340 119.915 ;
        RECT 56.520 119.320 57.180 119.800 ;
        RECT 57.380 119.710 57.550 120.470 ;
        RECT 58.450 120.300 58.630 120.710 ;
        RECT 57.720 120.130 58.050 120.250 ;
        RECT 58.800 120.130 58.970 120.890 ;
        RECT 57.720 119.960 58.970 120.130 ;
        RECT 59.140 121.070 60.510 121.320 ;
        RECT 59.140 120.300 59.330 121.070 ;
        RECT 60.260 120.810 60.510 121.070 ;
        RECT 59.500 120.640 59.750 120.800 ;
        RECT 60.680 120.640 60.850 121.485 ;
        RECT 61.745 121.200 61.915 121.700 ;
        RECT 62.085 121.370 62.415 121.870 ;
        RECT 61.020 120.810 61.520 121.190 ;
        RECT 61.745 121.030 62.440 121.200 ;
        RECT 59.500 120.470 60.850 120.640 ;
        RECT 60.430 120.430 60.850 120.470 ;
        RECT 59.140 119.960 59.560 120.300 ;
        RECT 59.850 119.970 60.260 120.300 ;
        RECT 57.380 119.540 58.230 119.710 ;
        RECT 58.790 119.320 59.110 119.780 ;
        RECT 59.310 119.530 59.560 119.960 ;
        RECT 59.850 119.320 60.260 119.760 ;
        RECT 60.430 119.700 60.600 120.430 ;
        RECT 60.770 119.880 61.120 120.250 ;
        RECT 61.300 119.940 61.520 120.810 ;
        RECT 61.690 120.240 62.100 120.860 ;
        RECT 62.270 120.060 62.440 121.030 ;
        RECT 61.745 119.870 62.440 120.060 ;
        RECT 60.430 119.500 61.445 119.700 ;
        RECT 61.745 119.540 61.915 119.870 ;
        RECT 62.085 119.320 62.415 119.700 ;
        RECT 62.630 119.580 62.855 121.700 ;
        RECT 63.025 121.370 63.355 121.870 ;
        RECT 63.525 121.200 63.695 121.700 ;
        RECT 63.030 121.030 63.695 121.200 ;
        RECT 63.030 120.040 63.260 121.030 ;
        RECT 63.430 120.210 63.780 120.860 ;
        RECT 63.955 120.705 64.245 121.870 ;
        RECT 64.415 120.795 64.685 121.700 ;
        RECT 64.855 121.110 65.185 121.870 ;
        RECT 65.365 120.940 65.535 121.700 ;
        RECT 63.030 119.870 63.695 120.040 ;
        RECT 63.025 119.320 63.355 119.700 ;
        RECT 63.525 119.580 63.695 119.870 ;
        RECT 63.955 119.320 64.245 120.045 ;
        RECT 64.415 119.995 64.585 120.795 ;
        RECT 64.870 120.770 65.535 120.940 ;
        RECT 65.795 120.780 68.385 121.870 ;
        RECT 64.870 120.625 65.040 120.770 ;
        RECT 64.755 120.295 65.040 120.625 ;
        RECT 64.870 120.040 65.040 120.295 ;
        RECT 65.275 120.220 65.605 120.590 ;
        RECT 65.795 120.260 67.005 120.780 ;
        RECT 68.595 120.730 68.825 121.870 ;
        RECT 68.995 120.720 69.325 121.700 ;
        RECT 69.495 120.730 69.705 121.870 ;
        RECT 69.935 121.110 70.450 121.520 ;
        RECT 70.685 121.110 70.855 121.870 ;
        RECT 71.025 121.530 73.055 121.700 ;
        RECT 67.175 120.090 68.385 120.610 ;
        RECT 68.575 120.310 68.905 120.560 ;
        RECT 64.415 119.490 64.675 119.995 ;
        RECT 64.870 119.870 65.535 120.040 ;
        RECT 64.855 119.320 65.185 119.700 ;
        RECT 65.365 119.490 65.535 119.870 ;
        RECT 65.795 119.320 68.385 120.090 ;
        RECT 68.595 119.320 68.825 120.140 ;
        RECT 69.075 120.120 69.325 120.720 ;
        RECT 69.935 120.300 70.275 121.110 ;
        RECT 71.025 120.865 71.195 121.530 ;
        RECT 71.590 121.190 72.715 121.360 ;
        RECT 70.445 120.675 71.195 120.865 ;
        RECT 71.365 120.850 72.375 121.020 ;
        RECT 68.995 119.490 69.325 120.120 ;
        RECT 69.495 119.320 69.705 120.140 ;
        RECT 69.935 120.130 71.165 120.300 ;
        RECT 70.210 119.525 70.455 120.130 ;
        RECT 70.675 119.320 71.185 119.855 ;
        RECT 71.365 119.490 71.555 120.850 ;
        RECT 71.725 119.830 72.000 120.650 ;
        RECT 72.205 120.050 72.375 120.850 ;
        RECT 72.545 120.060 72.715 121.190 ;
        RECT 72.885 120.560 73.055 121.530 ;
        RECT 73.225 120.730 73.395 121.870 ;
        RECT 73.565 120.730 73.900 121.700 ;
        RECT 72.885 120.230 73.080 120.560 ;
        RECT 73.305 120.230 73.560 120.560 ;
        RECT 73.305 120.060 73.475 120.230 ;
        RECT 73.730 120.060 73.900 120.730 ;
        RECT 74.075 120.780 75.745 121.870 ;
        RECT 75.915 121.110 76.430 121.520 ;
        RECT 76.665 121.110 76.835 121.870 ;
        RECT 77.005 121.530 79.035 121.700 ;
        RECT 74.075 120.260 74.825 120.780 ;
        RECT 74.995 120.090 75.745 120.610 ;
        RECT 75.915 120.300 76.255 121.110 ;
        RECT 77.005 120.865 77.175 121.530 ;
        RECT 77.570 121.190 78.695 121.360 ;
        RECT 76.425 120.675 77.175 120.865 ;
        RECT 77.345 120.850 78.355 121.020 ;
        RECT 75.915 120.130 77.145 120.300 ;
        RECT 72.545 119.890 73.475 120.060 ;
        RECT 72.545 119.855 72.720 119.890 ;
        RECT 71.725 119.660 72.005 119.830 ;
        RECT 71.725 119.490 72.000 119.660 ;
        RECT 72.190 119.490 72.720 119.855 ;
        RECT 73.145 119.320 73.475 119.720 ;
        RECT 73.645 119.490 73.900 120.060 ;
        RECT 74.075 119.320 75.745 120.090 ;
        RECT 76.190 119.525 76.435 120.130 ;
        RECT 76.655 119.320 77.165 119.855 ;
        RECT 77.345 119.490 77.535 120.850 ;
        RECT 77.705 120.510 77.980 120.650 ;
        RECT 77.705 120.340 77.985 120.510 ;
        RECT 77.705 119.490 77.980 120.340 ;
        RECT 78.185 120.050 78.355 120.850 ;
        RECT 78.525 120.060 78.695 121.190 ;
        RECT 78.865 120.560 79.035 121.530 ;
        RECT 79.205 120.730 79.375 121.870 ;
        RECT 79.545 120.730 79.880 121.700 ;
        RECT 78.865 120.230 79.060 120.560 ;
        RECT 79.285 120.230 79.540 120.560 ;
        RECT 79.285 120.060 79.455 120.230 ;
        RECT 79.710 120.060 79.880 120.730 ;
        RECT 80.430 120.890 80.685 121.560 ;
        RECT 80.865 121.070 81.150 121.870 ;
        RECT 81.330 121.150 81.660 121.660 ;
        RECT 80.430 120.170 80.610 120.890 ;
        RECT 81.330 120.560 81.580 121.150 ;
        RECT 81.930 121.000 82.100 121.610 ;
        RECT 82.270 121.180 82.600 121.870 ;
        RECT 82.830 121.320 83.070 121.610 ;
        RECT 83.270 121.490 83.690 121.870 ;
        RECT 83.870 121.400 84.500 121.650 ;
        RECT 84.970 121.490 85.300 121.870 ;
        RECT 83.870 121.320 84.040 121.400 ;
        RECT 85.470 121.320 85.640 121.610 ;
        RECT 85.820 121.490 86.200 121.870 ;
        RECT 86.440 121.485 87.270 121.655 ;
        RECT 82.830 121.150 84.040 121.320 ;
        RECT 80.780 120.230 81.580 120.560 ;
        RECT 78.525 119.890 79.455 120.060 ;
        RECT 78.525 119.855 78.700 119.890 ;
        RECT 78.170 119.490 78.700 119.855 ;
        RECT 79.125 119.320 79.455 119.720 ;
        RECT 79.625 119.490 79.880 120.060 ;
        RECT 80.345 120.030 80.610 120.170 ;
        RECT 80.345 120.000 80.685 120.030 ;
        RECT 80.430 119.500 80.685 120.000 ;
        RECT 80.865 119.320 81.150 119.780 ;
        RECT 81.330 119.580 81.580 120.230 ;
        RECT 81.780 120.980 82.100 121.000 ;
        RECT 81.780 120.810 83.700 120.980 ;
        RECT 81.780 119.915 81.970 120.810 ;
        RECT 83.870 120.640 84.040 121.150 ;
        RECT 84.210 120.890 84.730 121.200 ;
        RECT 82.140 120.470 84.040 120.640 ;
        RECT 82.140 120.410 82.470 120.470 ;
        RECT 82.620 120.240 82.950 120.300 ;
        RECT 82.290 119.970 82.950 120.240 ;
        RECT 81.780 119.585 82.100 119.915 ;
        RECT 82.280 119.320 82.940 119.800 ;
        RECT 83.140 119.710 83.310 120.470 ;
        RECT 84.210 120.300 84.390 120.710 ;
        RECT 83.480 120.130 83.810 120.250 ;
        RECT 84.560 120.130 84.730 120.890 ;
        RECT 83.480 119.960 84.730 120.130 ;
        RECT 84.900 121.070 86.270 121.320 ;
        RECT 84.900 120.300 85.090 121.070 ;
        RECT 86.020 120.810 86.270 121.070 ;
        RECT 85.260 120.640 85.510 120.800 ;
        RECT 86.440 120.640 86.610 121.485 ;
        RECT 87.505 121.200 87.675 121.700 ;
        RECT 87.845 121.370 88.175 121.870 ;
        RECT 86.780 120.810 87.280 121.190 ;
        RECT 87.505 121.030 88.200 121.200 ;
        RECT 85.260 120.470 86.610 120.640 ;
        RECT 86.190 120.430 86.610 120.470 ;
        RECT 84.900 119.960 85.320 120.300 ;
        RECT 85.610 119.970 86.020 120.300 ;
        RECT 83.140 119.540 83.990 119.710 ;
        RECT 84.550 119.320 84.870 119.780 ;
        RECT 85.070 119.530 85.320 119.960 ;
        RECT 85.610 119.320 86.020 119.760 ;
        RECT 86.190 119.700 86.360 120.430 ;
        RECT 86.530 119.880 86.880 120.250 ;
        RECT 87.060 119.940 87.280 120.810 ;
        RECT 87.450 120.240 87.860 120.860 ;
        RECT 88.030 120.060 88.200 121.030 ;
        RECT 87.505 119.870 88.200 120.060 ;
        RECT 86.190 119.500 87.205 119.700 ;
        RECT 87.505 119.540 87.675 119.870 ;
        RECT 87.845 119.320 88.175 119.700 ;
        RECT 88.390 119.580 88.615 121.700 ;
        RECT 88.785 121.370 89.115 121.870 ;
        RECT 89.285 121.200 89.455 121.700 ;
        RECT 88.790 121.030 89.455 121.200 ;
        RECT 88.790 120.040 89.020 121.030 ;
        RECT 89.190 120.210 89.540 120.860 ;
        RECT 89.715 120.705 90.005 121.870 ;
        RECT 90.550 121.530 90.805 121.560 ;
        RECT 90.465 121.360 90.805 121.530 ;
        RECT 90.550 120.890 90.805 121.360 ;
        RECT 90.985 121.070 91.270 121.870 ;
        RECT 91.450 121.150 91.780 121.660 ;
        RECT 88.790 119.870 89.455 120.040 ;
        RECT 88.785 119.320 89.115 119.700 ;
        RECT 89.285 119.580 89.455 119.870 ;
        RECT 89.715 119.320 90.005 120.045 ;
        RECT 90.550 120.030 90.730 120.890 ;
        RECT 91.450 120.560 91.700 121.150 ;
        RECT 92.050 121.000 92.220 121.610 ;
        RECT 92.390 121.180 92.720 121.870 ;
        RECT 92.950 121.320 93.190 121.610 ;
        RECT 93.390 121.490 93.810 121.870 ;
        RECT 93.990 121.400 94.620 121.650 ;
        RECT 95.090 121.490 95.420 121.870 ;
        RECT 93.990 121.320 94.160 121.400 ;
        RECT 95.590 121.320 95.760 121.610 ;
        RECT 95.940 121.490 96.320 121.870 ;
        RECT 96.560 121.485 97.390 121.655 ;
        RECT 92.950 121.150 94.160 121.320 ;
        RECT 90.900 120.230 91.700 120.560 ;
        RECT 90.550 119.500 90.805 120.030 ;
        RECT 90.985 119.320 91.270 119.780 ;
        RECT 91.450 119.580 91.700 120.230 ;
        RECT 91.900 120.980 92.220 121.000 ;
        RECT 91.900 120.810 93.820 120.980 ;
        RECT 91.900 119.915 92.090 120.810 ;
        RECT 93.990 120.640 94.160 121.150 ;
        RECT 94.330 120.890 94.850 121.200 ;
        RECT 92.260 120.470 94.160 120.640 ;
        RECT 92.260 120.410 92.590 120.470 ;
        RECT 92.740 120.240 93.070 120.300 ;
        RECT 92.410 119.970 93.070 120.240 ;
        RECT 91.900 119.585 92.220 119.915 ;
        RECT 92.400 119.320 93.060 119.800 ;
        RECT 93.260 119.710 93.430 120.470 ;
        RECT 94.330 120.300 94.510 120.710 ;
        RECT 93.600 120.130 93.930 120.250 ;
        RECT 94.680 120.130 94.850 120.890 ;
        RECT 93.600 119.960 94.850 120.130 ;
        RECT 95.020 121.070 96.390 121.320 ;
        RECT 95.020 120.300 95.210 121.070 ;
        RECT 96.140 120.810 96.390 121.070 ;
        RECT 95.380 120.640 95.630 120.800 ;
        RECT 96.560 120.640 96.730 121.485 ;
        RECT 97.625 121.200 97.795 121.700 ;
        RECT 97.965 121.370 98.295 121.870 ;
        RECT 96.900 120.810 97.400 121.190 ;
        RECT 97.625 121.030 98.320 121.200 ;
        RECT 95.380 120.470 96.730 120.640 ;
        RECT 96.310 120.430 96.730 120.470 ;
        RECT 95.020 119.960 95.440 120.300 ;
        RECT 95.730 119.970 96.140 120.300 ;
        RECT 93.260 119.540 94.110 119.710 ;
        RECT 94.670 119.320 94.990 119.780 ;
        RECT 95.190 119.530 95.440 119.960 ;
        RECT 95.730 119.320 96.140 119.760 ;
        RECT 96.310 119.700 96.480 120.430 ;
        RECT 96.650 119.880 97.000 120.250 ;
        RECT 97.180 119.940 97.400 120.810 ;
        RECT 97.570 120.240 97.980 120.860 ;
        RECT 98.150 120.060 98.320 121.030 ;
        RECT 97.625 119.870 98.320 120.060 ;
        RECT 96.310 119.500 97.325 119.700 ;
        RECT 97.625 119.540 97.795 119.870 ;
        RECT 97.965 119.320 98.295 119.700 ;
        RECT 98.510 119.580 98.735 121.700 ;
        RECT 98.905 121.370 99.235 121.870 ;
        RECT 99.405 121.200 99.575 121.700 ;
        RECT 98.910 121.030 99.575 121.200 ;
        RECT 98.910 120.040 99.140 121.030 ;
        RECT 100.210 120.890 100.465 121.560 ;
        RECT 100.645 121.070 100.930 121.870 ;
        RECT 101.110 121.150 101.440 121.660 ;
        RECT 99.310 120.210 99.660 120.860 ;
        RECT 98.910 119.870 99.575 120.040 ;
        RECT 98.905 119.320 99.235 119.700 ;
        RECT 99.405 119.580 99.575 119.870 ;
        RECT 100.210 120.030 100.390 120.890 ;
        RECT 101.110 120.560 101.360 121.150 ;
        RECT 101.710 121.000 101.880 121.610 ;
        RECT 102.050 121.180 102.380 121.870 ;
        RECT 102.610 121.320 102.850 121.610 ;
        RECT 103.050 121.490 103.470 121.870 ;
        RECT 103.650 121.400 104.280 121.650 ;
        RECT 104.750 121.490 105.080 121.870 ;
        RECT 103.650 121.320 103.820 121.400 ;
        RECT 105.250 121.320 105.420 121.610 ;
        RECT 105.600 121.490 105.980 121.870 ;
        RECT 106.220 121.485 107.050 121.655 ;
        RECT 102.610 121.150 103.820 121.320 ;
        RECT 100.560 120.230 101.360 120.560 ;
        RECT 100.210 119.830 100.465 120.030 ;
        RECT 100.125 119.660 100.465 119.830 ;
        RECT 100.210 119.500 100.465 119.660 ;
        RECT 100.645 119.320 100.930 119.780 ;
        RECT 101.110 119.580 101.360 120.230 ;
        RECT 101.560 120.980 101.880 121.000 ;
        RECT 101.560 120.810 103.480 120.980 ;
        RECT 101.560 119.915 101.750 120.810 ;
        RECT 103.650 120.640 103.820 121.150 ;
        RECT 103.990 120.890 104.510 121.200 ;
        RECT 101.920 120.470 103.820 120.640 ;
        RECT 101.920 120.410 102.250 120.470 ;
        RECT 102.400 120.240 102.730 120.300 ;
        RECT 102.070 119.970 102.730 120.240 ;
        RECT 101.560 119.585 101.880 119.915 ;
        RECT 102.060 119.320 102.720 119.800 ;
        RECT 102.920 119.710 103.090 120.470 ;
        RECT 103.990 120.300 104.170 120.710 ;
        RECT 103.260 120.130 103.590 120.250 ;
        RECT 104.340 120.130 104.510 120.890 ;
        RECT 103.260 119.960 104.510 120.130 ;
        RECT 104.680 121.070 106.050 121.320 ;
        RECT 104.680 120.300 104.870 121.070 ;
        RECT 105.800 120.810 106.050 121.070 ;
        RECT 105.040 120.640 105.290 120.800 ;
        RECT 106.220 120.640 106.390 121.485 ;
        RECT 107.285 121.200 107.455 121.700 ;
        RECT 107.625 121.370 107.955 121.870 ;
        RECT 106.560 120.810 107.060 121.190 ;
        RECT 107.285 121.030 107.980 121.200 ;
        RECT 105.040 120.470 106.390 120.640 ;
        RECT 105.970 120.430 106.390 120.470 ;
        RECT 104.680 119.960 105.100 120.300 ;
        RECT 105.390 119.970 105.800 120.300 ;
        RECT 102.920 119.540 103.770 119.710 ;
        RECT 104.330 119.320 104.650 119.780 ;
        RECT 104.850 119.530 105.100 119.960 ;
        RECT 105.390 119.320 105.800 119.760 ;
        RECT 105.970 119.700 106.140 120.430 ;
        RECT 106.310 119.880 106.660 120.250 ;
        RECT 106.840 119.940 107.060 120.810 ;
        RECT 107.230 120.240 107.640 120.860 ;
        RECT 107.810 120.060 107.980 121.030 ;
        RECT 107.285 119.870 107.980 120.060 ;
        RECT 105.970 119.500 106.985 119.700 ;
        RECT 107.285 119.540 107.455 119.870 ;
        RECT 107.625 119.320 107.955 119.700 ;
        RECT 108.170 119.580 108.395 121.700 ;
        RECT 108.565 121.370 108.895 121.870 ;
        RECT 109.065 121.200 109.235 121.700 ;
        RECT 108.570 121.030 109.235 121.200 ;
        RECT 108.570 120.040 108.800 121.030 ;
        RECT 108.970 120.210 109.320 120.860 ;
        RECT 109.495 120.780 110.705 121.870 ;
        RECT 110.875 120.780 114.385 121.870 ;
        RECT 114.555 120.780 115.765 121.870 ;
        RECT 109.495 120.240 110.015 120.780 ;
        RECT 110.185 120.070 110.705 120.610 ;
        RECT 110.875 120.260 112.565 120.780 ;
        RECT 112.735 120.090 114.385 120.610 ;
        RECT 114.555 120.240 115.075 120.780 ;
        RECT 108.570 119.870 109.235 120.040 ;
        RECT 108.565 119.320 108.895 119.700 ;
        RECT 109.065 119.580 109.235 119.870 ;
        RECT 109.495 119.320 110.705 120.070 ;
        RECT 110.875 119.320 114.385 120.090 ;
        RECT 115.245 120.070 115.765 120.610 ;
        RECT 114.555 119.320 115.765 120.070 ;
        RECT 10.510 119.150 115.850 119.320 ;
        RECT 10.595 118.400 11.805 119.150 ;
        RECT 10.595 117.860 11.115 118.400 ;
        RECT 11.975 118.380 13.645 119.150 ;
        RECT 13.905 118.600 14.075 118.890 ;
        RECT 14.245 118.770 14.575 119.150 ;
        RECT 13.905 118.430 14.570 118.600 ;
        RECT 11.285 117.690 11.805 118.230 ;
        RECT 10.595 116.600 11.805 117.690 ;
        RECT 11.975 117.690 12.725 118.210 ;
        RECT 12.895 117.860 13.645 118.380 ;
        RECT 11.975 116.600 13.645 117.690 ;
        RECT 13.820 117.610 14.170 118.260 ;
        RECT 14.340 117.440 14.570 118.430 ;
        RECT 13.905 117.270 14.570 117.440 ;
        RECT 13.905 116.770 14.075 117.270 ;
        RECT 14.245 116.600 14.575 117.100 ;
        RECT 14.745 116.770 14.970 118.890 ;
        RECT 15.185 118.770 15.515 119.150 ;
        RECT 15.685 118.600 15.855 118.930 ;
        RECT 16.155 118.770 17.170 118.970 ;
        RECT 15.160 118.410 15.855 118.600 ;
        RECT 15.160 117.440 15.330 118.410 ;
        RECT 15.500 117.610 15.910 118.230 ;
        RECT 16.080 117.660 16.300 118.530 ;
        RECT 16.480 118.220 16.830 118.590 ;
        RECT 17.000 118.040 17.170 118.770 ;
        RECT 17.340 118.710 17.750 119.150 ;
        RECT 18.040 118.510 18.290 118.940 ;
        RECT 18.490 118.690 18.810 119.150 ;
        RECT 19.370 118.760 20.220 118.930 ;
        RECT 17.340 118.170 17.750 118.500 ;
        RECT 18.040 118.170 18.460 118.510 ;
        RECT 16.750 118.000 17.170 118.040 ;
        RECT 16.750 117.830 18.100 118.000 ;
        RECT 15.160 117.270 15.855 117.440 ;
        RECT 16.080 117.280 16.580 117.660 ;
        RECT 15.185 116.600 15.515 117.100 ;
        RECT 15.685 116.770 15.855 117.270 ;
        RECT 16.750 116.985 16.920 117.830 ;
        RECT 17.850 117.670 18.100 117.830 ;
        RECT 17.090 117.400 17.340 117.660 ;
        RECT 18.270 117.400 18.460 118.170 ;
        RECT 17.090 117.150 18.460 117.400 ;
        RECT 18.630 118.340 19.880 118.510 ;
        RECT 18.630 117.580 18.800 118.340 ;
        RECT 19.550 118.220 19.880 118.340 ;
        RECT 18.970 117.760 19.150 118.170 ;
        RECT 20.050 118.000 20.220 118.760 ;
        RECT 20.420 118.670 21.080 119.150 ;
        RECT 21.260 118.555 21.580 118.885 ;
        RECT 20.410 118.230 21.070 118.500 ;
        RECT 20.410 118.170 20.740 118.230 ;
        RECT 20.890 118.000 21.220 118.060 ;
        RECT 19.320 117.830 21.220 118.000 ;
        RECT 18.630 117.270 19.150 117.580 ;
        RECT 19.320 117.320 19.490 117.830 ;
        RECT 21.390 117.660 21.580 118.555 ;
        RECT 19.660 117.490 21.580 117.660 ;
        RECT 21.260 117.470 21.580 117.490 ;
        RECT 21.780 118.240 22.030 118.890 ;
        RECT 22.210 118.690 22.495 119.150 ;
        RECT 22.675 118.810 22.930 118.970 ;
        RECT 22.675 118.640 23.015 118.810 ;
        RECT 22.675 118.440 22.930 118.640 ;
        RECT 21.780 117.910 22.580 118.240 ;
        RECT 19.320 117.150 20.530 117.320 ;
        RECT 16.090 116.815 16.920 116.985 ;
        RECT 17.160 116.600 17.540 116.980 ;
        RECT 17.720 116.860 17.890 117.150 ;
        RECT 19.320 117.070 19.490 117.150 ;
        RECT 18.060 116.600 18.390 116.980 ;
        RECT 18.860 116.820 19.490 117.070 ;
        RECT 19.670 116.600 20.090 116.980 ;
        RECT 20.290 116.860 20.530 117.150 ;
        RECT 20.760 116.600 21.090 117.290 ;
        RECT 21.260 116.860 21.430 117.470 ;
        RECT 21.780 117.320 22.030 117.910 ;
        RECT 22.750 117.580 22.930 118.440 ;
        RECT 23.475 118.380 25.145 119.150 ;
        RECT 25.315 118.425 25.605 119.150 ;
        RECT 26.150 118.810 26.405 118.970 ;
        RECT 26.065 118.640 26.405 118.810 ;
        RECT 26.585 118.690 26.870 119.150 ;
        RECT 26.150 118.440 26.405 118.640 ;
        RECT 21.700 116.810 22.030 117.320 ;
        RECT 22.210 116.600 22.495 117.400 ;
        RECT 22.675 116.910 22.930 117.580 ;
        RECT 23.475 117.690 24.225 118.210 ;
        RECT 24.395 117.860 25.145 118.380 ;
        RECT 23.475 116.600 25.145 117.690 ;
        RECT 25.315 116.600 25.605 117.765 ;
        RECT 26.150 117.580 26.330 118.440 ;
        RECT 27.050 118.240 27.300 118.890 ;
        RECT 26.500 117.910 27.300 118.240 ;
        RECT 26.150 116.910 26.405 117.580 ;
        RECT 26.585 116.600 26.870 117.400 ;
        RECT 27.050 117.320 27.300 117.910 ;
        RECT 27.500 118.555 27.820 118.885 ;
        RECT 28.000 118.670 28.660 119.150 ;
        RECT 28.860 118.760 29.710 118.930 ;
        RECT 27.500 117.660 27.690 118.555 ;
        RECT 28.010 118.230 28.670 118.500 ;
        RECT 28.340 118.170 28.670 118.230 ;
        RECT 27.860 118.000 28.190 118.060 ;
        RECT 28.860 118.000 29.030 118.760 ;
        RECT 30.270 118.690 30.590 119.150 ;
        RECT 30.790 118.510 31.040 118.940 ;
        RECT 31.330 118.710 31.740 119.150 ;
        RECT 31.910 118.770 32.925 118.970 ;
        RECT 29.200 118.340 30.450 118.510 ;
        RECT 29.200 118.220 29.530 118.340 ;
        RECT 27.860 117.830 29.760 118.000 ;
        RECT 27.500 117.490 29.420 117.660 ;
        RECT 27.500 117.470 27.820 117.490 ;
        RECT 27.050 116.810 27.380 117.320 ;
        RECT 27.650 116.860 27.820 117.470 ;
        RECT 29.590 117.320 29.760 117.830 ;
        RECT 29.930 117.760 30.110 118.170 ;
        RECT 30.280 117.580 30.450 118.340 ;
        RECT 27.990 116.600 28.320 117.290 ;
        RECT 28.550 117.150 29.760 117.320 ;
        RECT 29.930 117.270 30.450 117.580 ;
        RECT 30.620 118.170 31.040 118.510 ;
        RECT 31.330 118.170 31.740 118.500 ;
        RECT 30.620 117.400 30.810 118.170 ;
        RECT 31.910 118.040 32.080 118.770 ;
        RECT 33.225 118.600 33.395 118.930 ;
        RECT 33.565 118.770 33.895 119.150 ;
        RECT 32.250 118.220 32.600 118.590 ;
        RECT 31.910 118.000 32.330 118.040 ;
        RECT 30.980 117.830 32.330 118.000 ;
        RECT 30.980 117.670 31.230 117.830 ;
        RECT 31.740 117.400 31.990 117.660 ;
        RECT 30.620 117.150 31.990 117.400 ;
        RECT 28.550 116.860 28.790 117.150 ;
        RECT 29.590 117.070 29.760 117.150 ;
        RECT 28.990 116.600 29.410 116.980 ;
        RECT 29.590 116.820 30.220 117.070 ;
        RECT 30.690 116.600 31.020 116.980 ;
        RECT 31.190 116.860 31.360 117.150 ;
        RECT 32.160 116.985 32.330 117.830 ;
        RECT 32.780 117.660 33.000 118.530 ;
        RECT 33.225 118.410 33.920 118.600 ;
        RECT 32.500 117.280 33.000 117.660 ;
        RECT 33.170 117.610 33.580 118.230 ;
        RECT 33.750 117.440 33.920 118.410 ;
        RECT 33.225 117.270 33.920 117.440 ;
        RECT 31.540 116.600 31.920 116.980 ;
        RECT 32.160 116.815 32.990 116.985 ;
        RECT 33.225 116.770 33.395 117.270 ;
        RECT 33.565 116.600 33.895 117.100 ;
        RECT 34.110 116.770 34.335 118.890 ;
        RECT 34.505 118.770 34.835 119.150 ;
        RECT 35.005 118.600 35.175 118.890 ;
        RECT 34.510 118.430 35.175 118.600 ;
        RECT 35.435 118.475 35.695 118.980 ;
        RECT 35.875 118.770 36.205 119.150 ;
        RECT 36.385 118.600 36.555 118.980 ;
        RECT 34.510 117.440 34.740 118.430 ;
        RECT 34.910 117.610 35.260 118.260 ;
        RECT 35.435 117.675 35.605 118.475 ;
        RECT 35.890 118.430 36.555 118.600 ;
        RECT 35.890 118.175 36.060 118.430 ;
        RECT 38.010 118.340 38.255 118.945 ;
        RECT 38.475 118.615 38.985 119.150 ;
        RECT 35.775 117.845 36.060 118.175 ;
        RECT 36.295 117.880 36.625 118.250 ;
        RECT 37.735 118.170 38.965 118.340 ;
        RECT 35.890 117.700 36.060 117.845 ;
        RECT 34.510 117.270 35.175 117.440 ;
        RECT 34.505 116.600 34.835 117.100 ;
        RECT 35.005 116.770 35.175 117.270 ;
        RECT 35.435 116.770 35.705 117.675 ;
        RECT 35.890 117.530 36.555 117.700 ;
        RECT 35.875 116.600 36.205 117.360 ;
        RECT 36.385 116.770 36.555 117.530 ;
        RECT 37.735 117.360 38.075 118.170 ;
        RECT 38.245 117.605 38.995 117.795 ;
        RECT 37.735 116.950 38.250 117.360 ;
        RECT 38.485 116.600 38.655 117.360 ;
        RECT 38.825 116.940 38.995 117.605 ;
        RECT 39.165 117.620 39.355 118.980 ;
        RECT 39.525 118.130 39.800 118.980 ;
        RECT 39.990 118.615 40.520 118.980 ;
        RECT 40.945 118.750 41.275 119.150 ;
        RECT 40.345 118.580 40.520 118.615 ;
        RECT 39.525 117.960 39.805 118.130 ;
        RECT 39.525 117.820 39.800 117.960 ;
        RECT 40.005 117.620 40.175 118.420 ;
        RECT 39.165 117.450 40.175 117.620 ;
        RECT 40.345 118.410 41.275 118.580 ;
        RECT 41.445 118.410 41.700 118.980 ;
        RECT 41.875 118.640 42.180 119.150 ;
        RECT 40.345 117.280 40.515 118.410 ;
        RECT 41.105 118.240 41.275 118.410 ;
        RECT 39.390 117.110 40.515 117.280 ;
        RECT 40.685 117.910 40.880 118.240 ;
        RECT 41.105 117.910 41.360 118.240 ;
        RECT 40.685 116.940 40.855 117.910 ;
        RECT 41.530 117.740 41.700 118.410 ;
        RECT 41.875 117.910 42.190 118.470 ;
        RECT 42.360 118.160 42.610 118.970 ;
        RECT 42.780 118.625 43.040 119.150 ;
        RECT 43.220 118.160 43.470 118.970 ;
        RECT 43.640 118.590 43.900 119.150 ;
        RECT 44.070 118.500 44.330 118.955 ;
        RECT 44.500 118.670 44.760 119.150 ;
        RECT 44.930 118.500 45.190 118.955 ;
        RECT 45.360 118.670 45.620 119.150 ;
        RECT 45.790 118.500 46.050 118.955 ;
        RECT 46.220 118.670 46.465 119.150 ;
        RECT 46.635 118.500 46.910 118.955 ;
        RECT 47.080 118.670 47.325 119.150 ;
        RECT 47.495 118.500 47.755 118.955 ;
        RECT 47.935 118.670 48.185 119.150 ;
        RECT 48.355 118.500 48.615 118.955 ;
        RECT 48.795 118.670 49.045 119.150 ;
        RECT 49.215 118.500 49.475 118.955 ;
        RECT 49.655 118.670 49.915 119.150 ;
        RECT 50.085 118.500 50.345 118.955 ;
        RECT 50.515 118.670 50.815 119.150 ;
        RECT 44.070 118.330 50.815 118.500 ;
        RECT 51.075 118.425 51.365 119.150 ;
        RECT 51.535 118.475 51.795 118.980 ;
        RECT 51.975 118.770 52.305 119.150 ;
        RECT 52.485 118.600 52.655 118.980 ;
        RECT 42.360 117.910 49.480 118.160 ;
        RECT 38.825 116.770 40.855 116.940 ;
        RECT 41.025 116.600 41.195 117.740 ;
        RECT 41.365 116.770 41.700 117.740 ;
        RECT 41.885 116.600 42.180 117.410 ;
        RECT 42.360 116.770 42.605 117.910 ;
        RECT 42.780 116.600 43.040 117.410 ;
        RECT 43.220 116.775 43.470 117.910 ;
        RECT 49.650 117.740 50.815 118.330 ;
        RECT 44.070 117.515 50.815 117.740 ;
        RECT 44.070 117.500 49.475 117.515 ;
        RECT 43.640 116.605 43.900 117.400 ;
        RECT 44.070 116.775 44.330 117.500 ;
        RECT 44.500 116.605 44.760 117.330 ;
        RECT 44.930 116.775 45.190 117.500 ;
        RECT 45.360 116.605 45.620 117.330 ;
        RECT 45.790 116.775 46.050 117.500 ;
        RECT 46.220 116.605 46.480 117.330 ;
        RECT 46.650 116.775 46.910 117.500 ;
        RECT 47.080 116.605 47.325 117.330 ;
        RECT 47.495 116.775 47.755 117.500 ;
        RECT 47.940 116.605 48.185 117.330 ;
        RECT 48.355 116.775 48.615 117.500 ;
        RECT 48.800 116.605 49.045 117.330 ;
        RECT 49.215 116.775 49.475 117.500 ;
        RECT 49.660 116.605 49.915 117.330 ;
        RECT 50.085 116.775 50.375 117.515 ;
        RECT 43.640 116.600 49.915 116.605 ;
        RECT 50.545 116.600 50.815 117.345 ;
        RECT 51.075 116.600 51.365 117.765 ;
        RECT 51.535 117.675 51.705 118.475 ;
        RECT 51.990 118.430 52.655 118.600 ;
        RECT 53.465 118.600 53.635 118.890 ;
        RECT 53.805 118.770 54.135 119.150 ;
        RECT 53.465 118.430 54.130 118.600 ;
        RECT 51.990 118.175 52.160 118.430 ;
        RECT 51.875 117.845 52.160 118.175 ;
        RECT 52.395 117.880 52.725 118.250 ;
        RECT 51.990 117.700 52.160 117.845 ;
        RECT 51.535 116.770 51.805 117.675 ;
        RECT 51.990 117.530 52.655 117.700 ;
        RECT 53.380 117.610 53.730 118.260 ;
        RECT 51.975 116.600 52.305 117.360 ;
        RECT 52.485 116.770 52.655 117.530 ;
        RECT 53.900 117.440 54.130 118.430 ;
        RECT 53.465 117.270 54.130 117.440 ;
        RECT 53.465 116.770 53.635 117.270 ;
        RECT 53.805 116.600 54.135 117.100 ;
        RECT 54.305 116.770 54.530 118.890 ;
        RECT 54.745 118.770 55.075 119.150 ;
        RECT 55.245 118.600 55.415 118.930 ;
        RECT 55.715 118.770 56.730 118.970 ;
        RECT 54.720 118.410 55.415 118.600 ;
        RECT 54.720 117.440 54.890 118.410 ;
        RECT 55.060 117.610 55.470 118.230 ;
        RECT 55.640 117.660 55.860 118.530 ;
        RECT 56.040 118.220 56.390 118.590 ;
        RECT 56.560 118.040 56.730 118.770 ;
        RECT 56.900 118.710 57.310 119.150 ;
        RECT 57.600 118.510 57.850 118.940 ;
        RECT 58.050 118.690 58.370 119.150 ;
        RECT 58.930 118.760 59.780 118.930 ;
        RECT 56.900 118.170 57.310 118.500 ;
        RECT 57.600 118.170 58.020 118.510 ;
        RECT 56.310 118.000 56.730 118.040 ;
        RECT 56.310 117.830 57.660 118.000 ;
        RECT 54.720 117.270 55.415 117.440 ;
        RECT 55.640 117.280 56.140 117.660 ;
        RECT 54.745 116.600 55.075 117.100 ;
        RECT 55.245 116.770 55.415 117.270 ;
        RECT 56.310 116.985 56.480 117.830 ;
        RECT 57.410 117.670 57.660 117.830 ;
        RECT 56.650 117.400 56.900 117.660 ;
        RECT 57.830 117.400 58.020 118.170 ;
        RECT 56.650 117.150 58.020 117.400 ;
        RECT 58.190 118.340 59.440 118.510 ;
        RECT 58.190 117.580 58.360 118.340 ;
        RECT 59.110 118.220 59.440 118.340 ;
        RECT 58.530 117.760 58.710 118.170 ;
        RECT 59.610 118.000 59.780 118.760 ;
        RECT 59.980 118.670 60.640 119.150 ;
        RECT 60.820 118.555 61.140 118.885 ;
        RECT 59.970 118.230 60.630 118.500 ;
        RECT 59.970 118.170 60.300 118.230 ;
        RECT 60.450 118.000 60.780 118.060 ;
        RECT 58.880 117.830 60.780 118.000 ;
        RECT 58.190 117.270 58.710 117.580 ;
        RECT 58.880 117.320 59.050 117.830 ;
        RECT 60.950 117.660 61.140 118.555 ;
        RECT 59.220 117.490 61.140 117.660 ;
        RECT 60.820 117.470 61.140 117.490 ;
        RECT 61.340 118.240 61.590 118.890 ;
        RECT 61.770 118.690 62.055 119.150 ;
        RECT 62.235 118.810 62.490 118.970 ;
        RECT 62.235 118.640 62.575 118.810 ;
        RECT 62.235 118.440 62.490 118.640 ;
        RECT 61.340 117.910 62.140 118.240 ;
        RECT 58.880 117.150 60.090 117.320 ;
        RECT 55.650 116.815 56.480 116.985 ;
        RECT 56.720 116.600 57.100 116.980 ;
        RECT 57.280 116.860 57.450 117.150 ;
        RECT 58.880 117.070 59.050 117.150 ;
        RECT 57.620 116.600 57.950 116.980 ;
        RECT 58.420 116.820 59.050 117.070 ;
        RECT 59.230 116.600 59.650 116.980 ;
        RECT 59.850 116.860 60.090 117.150 ;
        RECT 60.320 116.600 60.650 117.290 ;
        RECT 60.820 116.860 60.990 117.470 ;
        RECT 61.340 117.320 61.590 117.910 ;
        RECT 62.310 117.580 62.490 118.440 ;
        RECT 63.035 118.380 65.625 119.150 ;
        RECT 66.170 118.810 66.425 118.970 ;
        RECT 66.085 118.640 66.425 118.810 ;
        RECT 66.605 118.690 66.890 119.150 ;
        RECT 61.260 116.810 61.590 117.320 ;
        RECT 61.770 116.600 62.055 117.400 ;
        RECT 62.235 116.910 62.490 117.580 ;
        RECT 63.035 117.690 64.245 118.210 ;
        RECT 64.415 117.860 65.625 118.380 ;
        RECT 66.170 118.440 66.425 118.640 ;
        RECT 63.035 116.600 65.625 117.690 ;
        RECT 66.170 117.580 66.350 118.440 ;
        RECT 67.070 118.240 67.320 118.890 ;
        RECT 66.520 117.910 67.320 118.240 ;
        RECT 66.170 116.910 66.425 117.580 ;
        RECT 66.605 116.600 66.890 117.400 ;
        RECT 67.070 117.320 67.320 117.910 ;
        RECT 67.520 118.555 67.840 118.885 ;
        RECT 68.020 118.670 68.680 119.150 ;
        RECT 68.880 118.760 69.730 118.930 ;
        RECT 67.520 117.660 67.710 118.555 ;
        RECT 68.030 118.230 68.690 118.500 ;
        RECT 68.360 118.170 68.690 118.230 ;
        RECT 67.880 118.000 68.210 118.060 ;
        RECT 68.880 118.000 69.050 118.760 ;
        RECT 70.290 118.690 70.610 119.150 ;
        RECT 70.810 118.510 71.060 118.940 ;
        RECT 71.350 118.710 71.760 119.150 ;
        RECT 71.930 118.770 72.945 118.970 ;
        RECT 69.220 118.340 70.470 118.510 ;
        RECT 69.220 118.220 69.550 118.340 ;
        RECT 67.880 117.830 69.780 118.000 ;
        RECT 67.520 117.490 69.440 117.660 ;
        RECT 67.520 117.470 67.840 117.490 ;
        RECT 67.070 116.810 67.400 117.320 ;
        RECT 67.670 116.860 67.840 117.470 ;
        RECT 69.610 117.320 69.780 117.830 ;
        RECT 69.950 117.760 70.130 118.170 ;
        RECT 70.300 117.580 70.470 118.340 ;
        RECT 68.010 116.600 68.340 117.290 ;
        RECT 68.570 117.150 69.780 117.320 ;
        RECT 69.950 117.270 70.470 117.580 ;
        RECT 70.640 118.170 71.060 118.510 ;
        RECT 71.350 118.170 71.760 118.500 ;
        RECT 70.640 117.400 70.830 118.170 ;
        RECT 71.930 118.040 72.100 118.770 ;
        RECT 73.245 118.600 73.415 118.930 ;
        RECT 73.585 118.770 73.915 119.150 ;
        RECT 72.270 118.220 72.620 118.590 ;
        RECT 71.930 118.000 72.350 118.040 ;
        RECT 71.000 117.830 72.350 118.000 ;
        RECT 71.000 117.670 71.250 117.830 ;
        RECT 71.760 117.400 72.010 117.660 ;
        RECT 70.640 117.150 72.010 117.400 ;
        RECT 68.570 116.860 68.810 117.150 ;
        RECT 69.610 117.070 69.780 117.150 ;
        RECT 69.010 116.600 69.430 116.980 ;
        RECT 69.610 116.820 70.240 117.070 ;
        RECT 70.710 116.600 71.040 116.980 ;
        RECT 71.210 116.860 71.380 117.150 ;
        RECT 72.180 116.985 72.350 117.830 ;
        RECT 72.800 117.660 73.020 118.530 ;
        RECT 73.245 118.410 73.940 118.600 ;
        RECT 72.520 117.280 73.020 117.660 ;
        RECT 73.190 117.610 73.600 118.230 ;
        RECT 73.770 117.440 73.940 118.410 ;
        RECT 73.245 117.270 73.940 117.440 ;
        RECT 71.560 116.600 71.940 116.980 ;
        RECT 72.180 116.815 73.010 116.985 ;
        RECT 73.245 116.770 73.415 117.270 ;
        RECT 73.585 116.600 73.915 117.100 ;
        RECT 74.130 116.770 74.355 118.890 ;
        RECT 74.525 118.770 74.855 119.150 ;
        RECT 75.025 118.600 75.195 118.890 ;
        RECT 74.530 118.430 75.195 118.600 ;
        RECT 74.530 117.440 74.760 118.430 ;
        RECT 75.495 118.330 75.725 119.150 ;
        RECT 75.895 118.350 76.225 118.980 ;
        RECT 74.930 117.610 75.280 118.260 ;
        RECT 75.475 117.910 75.805 118.160 ;
        RECT 75.975 117.750 76.225 118.350 ;
        RECT 76.395 118.330 76.605 119.150 ;
        RECT 76.835 118.425 77.125 119.150 ;
        RECT 77.670 118.440 77.925 118.970 ;
        RECT 78.105 118.690 78.390 119.150 ;
        RECT 74.530 117.270 75.195 117.440 ;
        RECT 74.525 116.600 74.855 117.100 ;
        RECT 75.025 116.770 75.195 117.270 ;
        RECT 75.495 116.600 75.725 117.740 ;
        RECT 75.895 116.770 76.225 117.750 ;
        RECT 76.395 116.600 76.605 117.740 ;
        RECT 76.835 116.600 77.125 117.765 ;
        RECT 77.670 117.580 77.850 118.440 ;
        RECT 78.570 118.240 78.820 118.890 ;
        RECT 78.020 117.910 78.820 118.240 ;
        RECT 77.670 117.110 77.925 117.580 ;
        RECT 77.585 116.940 77.925 117.110 ;
        RECT 77.670 116.910 77.925 116.940 ;
        RECT 78.105 116.600 78.390 117.400 ;
        RECT 78.570 117.320 78.820 117.910 ;
        RECT 79.020 118.555 79.340 118.885 ;
        RECT 79.520 118.670 80.180 119.150 ;
        RECT 80.380 118.760 81.230 118.930 ;
        RECT 79.020 117.660 79.210 118.555 ;
        RECT 79.530 118.230 80.190 118.500 ;
        RECT 79.860 118.170 80.190 118.230 ;
        RECT 79.380 118.000 79.710 118.060 ;
        RECT 80.380 118.000 80.550 118.760 ;
        RECT 81.790 118.690 82.110 119.150 ;
        RECT 82.310 118.510 82.560 118.940 ;
        RECT 82.850 118.710 83.260 119.150 ;
        RECT 83.430 118.770 84.445 118.970 ;
        RECT 80.720 118.340 81.970 118.510 ;
        RECT 80.720 118.220 81.050 118.340 ;
        RECT 79.380 117.830 81.280 118.000 ;
        RECT 79.020 117.490 80.940 117.660 ;
        RECT 79.020 117.470 79.340 117.490 ;
        RECT 78.570 116.810 78.900 117.320 ;
        RECT 79.170 116.860 79.340 117.470 ;
        RECT 81.110 117.320 81.280 117.830 ;
        RECT 81.450 117.760 81.630 118.170 ;
        RECT 81.800 117.580 81.970 118.340 ;
        RECT 79.510 116.600 79.840 117.290 ;
        RECT 80.070 117.150 81.280 117.320 ;
        RECT 81.450 117.270 81.970 117.580 ;
        RECT 82.140 118.170 82.560 118.510 ;
        RECT 82.850 118.170 83.260 118.500 ;
        RECT 82.140 117.400 82.330 118.170 ;
        RECT 83.430 118.040 83.600 118.770 ;
        RECT 84.745 118.600 84.915 118.930 ;
        RECT 85.085 118.770 85.415 119.150 ;
        RECT 83.770 118.220 84.120 118.590 ;
        RECT 83.430 118.000 83.850 118.040 ;
        RECT 82.500 117.830 83.850 118.000 ;
        RECT 82.500 117.670 82.750 117.830 ;
        RECT 83.260 117.400 83.510 117.660 ;
        RECT 82.140 117.150 83.510 117.400 ;
        RECT 80.070 116.860 80.310 117.150 ;
        RECT 81.110 117.070 81.280 117.150 ;
        RECT 80.510 116.600 80.930 116.980 ;
        RECT 81.110 116.820 81.740 117.070 ;
        RECT 82.210 116.600 82.540 116.980 ;
        RECT 82.710 116.860 82.880 117.150 ;
        RECT 83.680 116.985 83.850 117.830 ;
        RECT 84.300 117.660 84.520 118.530 ;
        RECT 84.745 118.410 85.440 118.600 ;
        RECT 84.020 117.280 84.520 117.660 ;
        RECT 84.690 117.610 85.100 118.230 ;
        RECT 85.270 117.440 85.440 118.410 ;
        RECT 84.745 117.270 85.440 117.440 ;
        RECT 83.060 116.600 83.440 116.980 ;
        RECT 83.680 116.815 84.510 116.985 ;
        RECT 84.745 116.770 84.915 117.270 ;
        RECT 85.085 116.600 85.415 117.100 ;
        RECT 85.630 116.770 85.855 118.890 ;
        RECT 86.025 118.770 86.355 119.150 ;
        RECT 86.525 118.600 86.695 118.890 ;
        RECT 86.030 118.430 86.695 118.600 ;
        RECT 86.955 118.475 87.215 118.980 ;
        RECT 87.395 118.770 87.725 119.150 ;
        RECT 87.905 118.600 88.075 118.980 ;
        RECT 86.030 117.440 86.260 118.430 ;
        RECT 86.430 117.610 86.780 118.260 ;
        RECT 86.955 117.675 87.125 118.475 ;
        RECT 87.410 118.430 88.075 118.600 ;
        RECT 88.795 118.475 89.055 118.980 ;
        RECT 89.235 118.770 89.565 119.150 ;
        RECT 89.745 118.600 89.915 118.980 ;
        RECT 87.410 118.175 87.580 118.430 ;
        RECT 87.295 117.845 87.580 118.175 ;
        RECT 87.815 117.880 88.145 118.250 ;
        RECT 87.410 117.700 87.580 117.845 ;
        RECT 86.030 117.270 86.695 117.440 ;
        RECT 86.025 116.600 86.355 117.100 ;
        RECT 86.525 116.770 86.695 117.270 ;
        RECT 86.955 116.770 87.225 117.675 ;
        RECT 87.410 117.530 88.075 117.700 ;
        RECT 87.395 116.600 87.725 117.360 ;
        RECT 87.905 116.770 88.075 117.530 ;
        RECT 88.795 117.675 88.965 118.475 ;
        RECT 89.250 118.430 89.915 118.600 ;
        RECT 89.250 118.175 89.420 118.430 ;
        RECT 91.095 118.380 94.605 119.150 ;
        RECT 89.135 117.845 89.420 118.175 ;
        RECT 89.655 117.880 89.985 118.250 ;
        RECT 89.250 117.700 89.420 117.845 ;
        RECT 88.795 116.770 89.065 117.675 ;
        RECT 89.250 117.530 89.915 117.700 ;
        RECT 89.235 116.600 89.565 117.360 ;
        RECT 89.745 116.770 89.915 117.530 ;
        RECT 91.095 117.690 92.785 118.210 ;
        RECT 92.955 117.860 94.605 118.380 ;
        RECT 94.815 118.330 95.045 119.150 ;
        RECT 95.215 118.350 95.545 118.980 ;
        RECT 94.795 117.910 95.125 118.160 ;
        RECT 95.295 117.750 95.545 118.350 ;
        RECT 95.715 118.330 95.925 119.150 ;
        RECT 96.245 118.600 96.415 118.980 ;
        RECT 96.595 118.770 96.925 119.150 ;
        RECT 96.245 118.430 96.910 118.600 ;
        RECT 97.105 118.475 97.365 118.980 ;
        RECT 96.175 117.880 96.505 118.250 ;
        RECT 96.740 118.175 96.910 118.430 ;
        RECT 91.095 116.600 94.605 117.690 ;
        RECT 94.815 116.600 95.045 117.740 ;
        RECT 95.215 116.770 95.545 117.750 ;
        RECT 96.740 117.845 97.025 118.175 ;
        RECT 95.715 116.600 95.925 117.740 ;
        RECT 96.740 117.700 96.910 117.845 ;
        RECT 96.245 117.530 96.910 117.700 ;
        RECT 97.195 117.675 97.365 118.475 ;
        RECT 98.730 118.340 98.975 118.945 ;
        RECT 99.195 118.615 99.705 119.150 ;
        RECT 96.245 116.770 96.415 117.530 ;
        RECT 96.595 116.600 96.925 117.360 ;
        RECT 97.095 116.770 97.365 117.675 ;
        RECT 98.455 118.170 99.685 118.340 ;
        RECT 98.455 117.360 98.795 118.170 ;
        RECT 98.965 117.605 99.715 117.795 ;
        RECT 98.455 116.950 98.970 117.360 ;
        RECT 99.205 116.600 99.375 117.360 ;
        RECT 99.545 116.940 99.715 117.605 ;
        RECT 99.885 117.620 100.075 118.980 ;
        RECT 100.245 118.810 100.520 118.980 ;
        RECT 100.245 118.640 100.525 118.810 ;
        RECT 100.245 117.820 100.520 118.640 ;
        RECT 100.710 118.615 101.240 118.980 ;
        RECT 101.665 118.750 101.995 119.150 ;
        RECT 101.065 118.580 101.240 118.615 ;
        RECT 100.725 117.620 100.895 118.420 ;
        RECT 99.885 117.450 100.895 117.620 ;
        RECT 101.065 118.410 101.995 118.580 ;
        RECT 102.165 118.410 102.420 118.980 ;
        RECT 102.595 118.425 102.885 119.150 ;
        RECT 103.055 118.645 103.340 119.150 ;
        RECT 103.510 118.475 103.835 118.980 ;
        RECT 101.065 117.280 101.235 118.410 ;
        RECT 101.825 118.240 101.995 118.410 ;
        RECT 100.110 117.110 101.235 117.280 ;
        RECT 101.405 117.910 101.600 118.240 ;
        RECT 101.825 117.910 102.080 118.240 ;
        RECT 101.405 116.940 101.575 117.910 ;
        RECT 102.250 117.740 102.420 118.410 ;
        RECT 103.055 117.945 103.835 118.475 ;
        RECT 99.545 116.770 101.575 116.940 ;
        RECT 101.745 116.600 101.915 117.740 ;
        RECT 102.085 116.770 102.420 117.740 ;
        RECT 102.595 116.600 102.885 117.765 ;
        RECT 103.055 116.600 103.335 117.570 ;
        RECT 103.505 116.770 103.835 117.945 ;
        RECT 104.025 117.910 104.265 118.860 ;
        RECT 104.435 118.380 106.105 119.150 ;
        RECT 104.435 117.690 105.185 118.210 ;
        RECT 105.355 117.860 106.105 118.380 ;
        RECT 106.315 118.330 106.545 119.150 ;
        RECT 106.715 118.350 107.045 118.980 ;
        RECT 106.295 117.910 106.625 118.160 ;
        RECT 106.795 117.750 107.045 118.350 ;
        RECT 107.215 118.330 107.425 119.150 ;
        RECT 107.655 118.400 108.865 119.150 ;
        RECT 109.040 118.605 114.385 119.150 ;
        RECT 104.005 116.600 104.265 117.570 ;
        RECT 104.435 116.600 106.105 117.690 ;
        RECT 106.315 116.600 106.545 117.740 ;
        RECT 106.715 116.770 107.045 117.750 ;
        RECT 107.215 116.600 107.425 117.740 ;
        RECT 107.655 117.690 108.175 118.230 ;
        RECT 108.345 117.860 108.865 118.400 ;
        RECT 107.655 116.600 108.865 117.690 ;
        RECT 110.630 117.035 110.980 118.285 ;
        RECT 112.460 117.775 112.800 118.605 ;
        RECT 114.555 118.400 115.765 119.150 ;
        RECT 114.555 117.690 115.075 118.230 ;
        RECT 115.245 117.860 115.765 118.400 ;
        RECT 109.040 116.600 114.385 117.035 ;
        RECT 114.555 116.600 115.765 117.690 ;
        RECT 10.510 116.430 115.850 116.600 ;
        RECT 10.595 115.340 11.805 116.430 ;
        RECT 10.595 114.630 11.115 115.170 ;
        RECT 11.285 114.800 11.805 115.340 ;
        RECT 12.435 115.265 12.725 116.430 ;
        RECT 13.815 115.340 17.325 116.430 ;
        RECT 13.815 114.820 15.505 115.340 ;
        RECT 17.555 115.290 17.765 116.430 ;
        RECT 17.935 115.280 18.265 116.260 ;
        RECT 18.435 115.290 18.665 116.430 ;
        RECT 19.795 115.340 23.305 116.430 ;
        RECT 23.480 115.995 28.825 116.430 ;
        RECT 15.675 114.650 17.325 115.170 ;
        RECT 10.595 113.880 11.805 114.630 ;
        RECT 12.435 113.880 12.725 114.605 ;
        RECT 13.815 113.880 17.325 114.650 ;
        RECT 17.555 113.880 17.765 114.700 ;
        RECT 17.935 114.680 18.185 115.280 ;
        RECT 18.355 114.870 18.685 115.120 ;
        RECT 19.795 114.820 21.485 115.340 ;
        RECT 17.935 114.050 18.265 114.680 ;
        RECT 18.435 113.880 18.665 114.700 ;
        RECT 21.655 114.650 23.305 115.170 ;
        RECT 25.070 114.745 25.420 115.995 ;
        RECT 29.035 115.290 29.265 116.430 ;
        RECT 29.435 115.280 29.765 116.260 ;
        RECT 29.935 115.290 30.145 116.430 ;
        RECT 30.375 115.340 32.045 116.430 ;
        RECT 32.305 115.500 32.475 116.260 ;
        RECT 32.655 115.670 32.985 116.430 ;
        RECT 19.795 113.880 23.305 114.650 ;
        RECT 26.900 114.425 27.240 115.255 ;
        RECT 29.015 114.870 29.345 115.120 ;
        RECT 23.480 113.880 28.825 114.425 ;
        RECT 29.035 113.880 29.265 114.700 ;
        RECT 29.515 114.680 29.765 115.280 ;
        RECT 30.375 114.820 31.125 115.340 ;
        RECT 32.305 115.330 32.970 115.500 ;
        RECT 33.155 115.355 33.425 116.260 ;
        RECT 32.800 115.185 32.970 115.330 ;
        RECT 29.435 114.050 29.765 114.680 ;
        RECT 29.935 113.880 30.145 114.700 ;
        RECT 31.295 114.650 32.045 115.170 ;
        RECT 32.235 114.780 32.565 115.150 ;
        RECT 32.800 114.855 33.085 115.185 ;
        RECT 30.375 113.880 32.045 114.650 ;
        RECT 32.800 114.600 32.970 114.855 ;
        RECT 32.305 114.430 32.970 114.600 ;
        RECT 33.255 114.555 33.425 115.355 ;
        RECT 34.055 115.670 34.570 116.080 ;
        RECT 34.805 115.670 34.975 116.430 ;
        RECT 35.145 116.090 37.175 116.260 ;
        RECT 34.055 114.860 34.395 115.670 ;
        RECT 35.145 115.425 35.315 116.090 ;
        RECT 35.710 115.750 36.835 115.920 ;
        RECT 34.565 115.235 35.315 115.425 ;
        RECT 35.485 115.410 36.495 115.580 ;
        RECT 34.055 114.690 35.285 114.860 ;
        RECT 32.305 114.050 32.475 114.430 ;
        RECT 32.655 113.880 32.985 114.260 ;
        RECT 33.165 114.050 33.425 114.555 ;
        RECT 34.330 114.085 34.575 114.690 ;
        RECT 34.795 113.880 35.305 114.415 ;
        RECT 35.485 114.050 35.675 115.410 ;
        RECT 35.845 115.070 36.120 115.210 ;
        RECT 35.845 114.900 36.125 115.070 ;
        RECT 35.845 114.050 36.120 114.900 ;
        RECT 36.325 114.610 36.495 115.410 ;
        RECT 36.665 114.620 36.835 115.750 ;
        RECT 37.005 115.120 37.175 116.090 ;
        RECT 37.345 115.290 37.515 116.430 ;
        RECT 37.685 115.290 38.020 116.260 ;
        RECT 37.005 114.790 37.200 115.120 ;
        RECT 37.425 114.790 37.680 115.120 ;
        RECT 37.425 114.620 37.595 114.790 ;
        RECT 37.850 114.620 38.020 115.290 ;
        RECT 38.195 115.265 38.485 116.430 ;
        RECT 38.655 115.340 41.245 116.430 ;
        RECT 38.655 114.820 39.865 115.340 ;
        RECT 41.475 115.290 41.685 116.430 ;
        RECT 41.855 115.280 42.185 116.260 ;
        RECT 42.355 115.290 42.585 116.430 ;
        RECT 43.255 115.340 44.925 116.430 ;
        RECT 40.035 114.650 41.245 115.170 ;
        RECT 36.665 114.450 37.595 114.620 ;
        RECT 36.665 114.415 36.840 114.450 ;
        RECT 36.310 114.050 36.840 114.415 ;
        RECT 37.265 113.880 37.595 114.280 ;
        RECT 37.765 114.050 38.020 114.620 ;
        RECT 38.195 113.880 38.485 114.605 ;
        RECT 38.655 113.880 41.245 114.650 ;
        RECT 41.475 113.880 41.685 114.700 ;
        RECT 41.855 114.680 42.105 115.280 ;
        RECT 42.275 114.870 42.605 115.120 ;
        RECT 43.255 114.820 44.005 115.340 ;
        RECT 45.245 115.280 45.575 116.430 ;
        RECT 45.745 115.410 45.915 116.260 ;
        RECT 46.085 115.630 46.415 116.430 ;
        RECT 46.585 115.410 46.755 116.260 ;
        RECT 46.935 115.630 47.175 116.430 ;
        RECT 47.345 115.450 47.675 116.260 ;
        RECT 45.745 115.240 46.755 115.410 ;
        RECT 46.960 115.280 47.675 115.450 ;
        RECT 47.855 115.340 51.365 116.430 ;
        RECT 51.540 115.995 56.885 116.430 ;
        RECT 41.855 114.050 42.185 114.680 ;
        RECT 42.355 113.880 42.585 114.700 ;
        RECT 44.175 114.650 44.925 115.170 ;
        RECT 45.745 115.070 46.240 115.240 ;
        RECT 45.745 114.900 46.245 115.070 ;
        RECT 46.960 115.040 47.130 115.280 ;
        RECT 45.745 114.700 46.240 114.900 ;
        RECT 46.630 114.870 47.130 115.040 ;
        RECT 47.300 114.870 47.680 115.110 ;
        RECT 46.960 114.700 47.130 114.870 ;
        RECT 47.855 114.820 49.545 115.340 ;
        RECT 43.255 113.880 44.925 114.650 ;
        RECT 45.245 113.880 45.575 114.680 ;
        RECT 45.745 114.530 46.755 114.700 ;
        RECT 46.960 114.530 47.595 114.700 ;
        RECT 49.715 114.650 51.365 115.170 ;
        RECT 53.130 114.745 53.480 115.995 ;
        RECT 57.095 115.290 57.325 116.430 ;
        RECT 57.495 115.280 57.825 116.260 ;
        RECT 57.995 115.290 58.205 116.430 ;
        RECT 58.440 115.995 63.785 116.430 ;
        RECT 45.745 114.050 45.915 114.530 ;
        RECT 46.085 113.880 46.415 114.360 ;
        RECT 46.585 114.050 46.755 114.530 ;
        RECT 47.005 113.880 47.245 114.360 ;
        RECT 47.425 114.050 47.595 114.530 ;
        RECT 47.855 113.880 51.365 114.650 ;
        RECT 54.960 114.425 55.300 115.255 ;
        RECT 57.075 114.870 57.405 115.120 ;
        RECT 51.540 113.880 56.885 114.425 ;
        RECT 57.095 113.880 57.325 114.700 ;
        RECT 57.575 114.680 57.825 115.280 ;
        RECT 60.030 114.745 60.380 115.995 ;
        RECT 63.955 115.265 64.245 116.430 ;
        RECT 65.335 115.340 68.845 116.430 ;
        RECT 57.495 114.050 57.825 114.680 ;
        RECT 57.995 113.880 58.205 114.700 ;
        RECT 61.860 114.425 62.200 115.255 ;
        RECT 65.335 114.820 67.025 115.340 ;
        RECT 69.055 115.290 69.285 116.430 ;
        RECT 69.455 115.280 69.785 116.260 ;
        RECT 69.955 115.290 70.165 116.430 ;
        RECT 70.855 115.340 72.525 116.430 ;
        RECT 72.695 115.355 72.965 116.260 ;
        RECT 73.135 115.670 73.465 116.430 ;
        RECT 73.645 115.500 73.815 116.260 ;
        RECT 67.195 114.650 68.845 115.170 ;
        RECT 69.035 114.870 69.365 115.120 ;
        RECT 58.440 113.880 63.785 114.425 ;
        RECT 63.955 113.880 64.245 114.605 ;
        RECT 65.335 113.880 68.845 114.650 ;
        RECT 69.055 113.880 69.285 114.700 ;
        RECT 69.535 114.680 69.785 115.280 ;
        RECT 70.855 114.820 71.605 115.340 ;
        RECT 69.455 114.050 69.785 114.680 ;
        RECT 69.955 113.880 70.165 114.700 ;
        RECT 71.775 114.650 72.525 115.170 ;
        RECT 70.855 113.880 72.525 114.650 ;
        RECT 72.695 114.555 72.865 115.355 ;
        RECT 73.150 115.330 73.815 115.500 ;
        RECT 74.075 115.340 75.745 116.430 ;
        RECT 75.920 115.995 81.265 116.430 ;
        RECT 73.150 115.185 73.320 115.330 ;
        RECT 73.035 114.855 73.320 115.185 ;
        RECT 73.150 114.600 73.320 114.855 ;
        RECT 73.555 114.780 73.885 115.150 ;
        RECT 74.075 114.820 74.825 115.340 ;
        RECT 74.995 114.650 75.745 115.170 ;
        RECT 77.510 114.745 77.860 115.995 ;
        RECT 81.475 115.290 81.705 116.430 ;
        RECT 81.875 115.280 82.205 116.260 ;
        RECT 82.375 115.290 82.585 116.430 ;
        RECT 82.815 115.340 84.025 116.430 ;
        RECT 84.200 115.995 89.545 116.430 ;
        RECT 72.695 114.050 72.955 114.555 ;
        RECT 73.150 114.430 73.815 114.600 ;
        RECT 73.135 113.880 73.465 114.260 ;
        RECT 73.645 114.050 73.815 114.430 ;
        RECT 74.075 113.880 75.745 114.650 ;
        RECT 79.340 114.425 79.680 115.255 ;
        RECT 81.455 114.870 81.785 115.120 ;
        RECT 75.920 113.880 81.265 114.425 ;
        RECT 81.475 113.880 81.705 114.700 ;
        RECT 81.955 114.680 82.205 115.280 ;
        RECT 82.815 114.800 83.335 115.340 ;
        RECT 81.875 114.050 82.205 114.680 ;
        RECT 82.375 113.880 82.585 114.700 ;
        RECT 83.505 114.630 84.025 115.170 ;
        RECT 85.790 114.745 86.140 115.995 ;
        RECT 89.715 115.265 90.005 116.430 ;
        RECT 90.180 115.995 95.525 116.430 ;
        RECT 95.700 115.995 101.045 116.430 ;
        RECT 82.815 113.880 84.025 114.630 ;
        RECT 87.620 114.425 87.960 115.255 ;
        RECT 91.770 114.745 92.120 115.995 ;
        RECT 84.200 113.880 89.545 114.425 ;
        RECT 89.715 113.880 90.005 114.605 ;
        RECT 93.600 114.425 93.940 115.255 ;
        RECT 97.290 114.745 97.640 115.995 ;
        RECT 101.305 115.500 101.475 116.260 ;
        RECT 101.655 115.670 101.985 116.430 ;
        RECT 101.305 115.330 101.970 115.500 ;
        RECT 102.155 115.355 102.425 116.260 ;
        RECT 99.120 114.425 99.460 115.255 ;
        RECT 101.800 115.185 101.970 115.330 ;
        RECT 101.235 114.780 101.565 115.150 ;
        RECT 101.800 114.855 102.085 115.185 ;
        RECT 101.800 114.600 101.970 114.855 ;
        RECT 101.305 114.430 101.970 114.600 ;
        RECT 102.255 114.555 102.425 115.355 ;
        RECT 103.055 115.340 106.565 116.430 ;
        RECT 106.735 115.355 107.005 116.260 ;
        RECT 107.175 115.670 107.505 116.430 ;
        RECT 107.685 115.500 107.855 116.260 ;
        RECT 103.055 114.820 104.745 115.340 ;
        RECT 104.915 114.650 106.565 115.170 ;
        RECT 90.180 113.880 95.525 114.425 ;
        RECT 95.700 113.880 101.045 114.425 ;
        RECT 101.305 114.050 101.475 114.430 ;
        RECT 101.655 113.880 101.985 114.260 ;
        RECT 102.165 114.050 102.425 114.555 ;
        RECT 103.055 113.880 106.565 114.650 ;
        RECT 106.735 114.555 106.905 115.355 ;
        RECT 107.190 115.330 107.855 115.500 ;
        RECT 107.190 115.185 107.360 115.330 ;
        RECT 108.155 115.290 108.385 116.430 ;
        RECT 108.555 115.280 108.885 116.260 ;
        RECT 109.055 115.290 109.265 116.430 ;
        RECT 110.415 115.355 110.685 116.260 ;
        RECT 110.855 115.670 111.185 116.430 ;
        RECT 111.365 115.500 111.535 116.260 ;
        RECT 107.075 114.855 107.360 115.185 ;
        RECT 107.190 114.600 107.360 114.855 ;
        RECT 107.595 114.780 107.925 115.150 ;
        RECT 108.135 114.870 108.465 115.120 ;
        RECT 106.735 114.050 106.995 114.555 ;
        RECT 107.190 114.430 107.855 114.600 ;
        RECT 107.175 113.880 107.505 114.260 ;
        RECT 107.685 114.050 107.855 114.430 ;
        RECT 108.155 113.880 108.385 114.700 ;
        RECT 108.635 114.680 108.885 115.280 ;
        RECT 108.555 114.050 108.885 114.680 ;
        RECT 109.055 113.880 109.265 114.700 ;
        RECT 110.415 114.555 110.585 115.355 ;
        RECT 110.870 115.330 111.535 115.500 ;
        RECT 111.795 115.340 114.385 116.430 ;
        RECT 114.555 115.340 115.765 116.430 ;
        RECT 110.870 115.185 111.040 115.330 ;
        RECT 110.755 114.855 111.040 115.185 ;
        RECT 110.870 114.600 111.040 114.855 ;
        RECT 111.275 114.780 111.605 115.150 ;
        RECT 111.795 114.820 113.005 115.340 ;
        RECT 113.175 114.650 114.385 115.170 ;
        RECT 114.555 114.800 115.075 115.340 ;
        RECT 110.415 114.050 110.675 114.555 ;
        RECT 110.870 114.430 111.535 114.600 ;
        RECT 110.855 113.880 111.185 114.260 ;
        RECT 111.365 114.050 111.535 114.430 ;
        RECT 111.795 113.880 114.385 114.650 ;
        RECT 115.245 114.630 115.765 115.170 ;
        RECT 114.555 113.880 115.765 114.630 ;
        RECT 10.510 113.710 115.850 113.880 ;
        RECT 10.595 112.960 11.805 113.710 ;
        RECT 11.975 112.960 13.185 113.710 ;
        RECT 10.595 112.420 11.115 112.960 ;
        RECT 11.285 112.250 11.805 112.790 ;
        RECT 10.595 111.160 11.805 112.250 ;
        RECT 11.975 112.250 12.495 112.790 ;
        RECT 12.665 112.420 13.185 112.960 ;
        RECT 13.355 112.940 16.865 113.710 ;
        RECT 17.040 113.165 22.385 113.710 ;
        RECT 13.355 112.250 15.045 112.770 ;
        RECT 15.215 112.420 16.865 112.940 ;
        RECT 11.975 111.160 13.185 112.250 ;
        RECT 13.355 111.160 16.865 112.250 ;
        RECT 18.630 111.595 18.980 112.845 ;
        RECT 20.460 112.335 20.800 113.165 ;
        RECT 22.555 113.035 22.815 113.540 ;
        RECT 22.995 113.330 23.325 113.710 ;
        RECT 23.505 113.160 23.675 113.540 ;
        RECT 22.555 112.235 22.725 113.035 ;
        RECT 23.010 112.990 23.675 113.160 ;
        RECT 23.010 112.735 23.180 112.990 ;
        RECT 23.935 112.960 25.145 113.710 ;
        RECT 25.315 112.985 25.605 113.710 ;
        RECT 26.240 113.165 31.585 113.710 ;
        RECT 22.895 112.405 23.180 112.735 ;
        RECT 23.415 112.440 23.745 112.810 ;
        RECT 23.010 112.260 23.180 112.405 ;
        RECT 17.040 111.160 22.385 111.595 ;
        RECT 22.555 111.330 22.825 112.235 ;
        RECT 23.010 112.090 23.675 112.260 ;
        RECT 22.995 111.160 23.325 111.920 ;
        RECT 23.505 111.330 23.675 112.090 ;
        RECT 23.935 112.250 24.455 112.790 ;
        RECT 24.625 112.420 25.145 112.960 ;
        RECT 23.935 111.160 25.145 112.250 ;
        RECT 25.315 111.160 25.605 112.325 ;
        RECT 27.830 111.595 28.180 112.845 ;
        RECT 29.660 112.335 30.000 113.165 ;
        RECT 31.845 113.160 32.015 113.540 ;
        RECT 32.195 113.330 32.525 113.710 ;
        RECT 31.845 112.990 32.510 113.160 ;
        RECT 32.705 113.035 32.965 113.540 ;
        RECT 31.775 112.440 32.105 112.810 ;
        RECT 32.340 112.735 32.510 112.990 ;
        RECT 32.340 112.405 32.625 112.735 ;
        RECT 32.340 112.260 32.510 112.405 ;
        RECT 31.845 112.090 32.510 112.260 ;
        RECT 32.795 112.235 32.965 113.035 ;
        RECT 33.595 112.940 37.105 113.710 ;
        RECT 26.240 111.160 31.585 111.595 ;
        RECT 31.845 111.330 32.015 112.090 ;
        RECT 32.195 111.160 32.525 111.920 ;
        RECT 32.695 111.330 32.965 112.235 ;
        RECT 33.595 112.250 35.285 112.770 ;
        RECT 35.455 112.420 37.105 112.940 ;
        RECT 37.275 113.035 37.535 113.540 ;
        RECT 37.715 113.330 38.045 113.710 ;
        RECT 38.225 113.160 38.395 113.540 ;
        RECT 38.660 113.165 44.005 113.710 ;
        RECT 44.180 113.165 49.525 113.710 ;
        RECT 33.595 111.160 37.105 112.250 ;
        RECT 37.275 112.235 37.445 113.035 ;
        RECT 37.730 112.990 38.395 113.160 ;
        RECT 37.730 112.735 37.900 112.990 ;
        RECT 37.615 112.405 37.900 112.735 ;
        RECT 38.135 112.440 38.465 112.810 ;
        RECT 37.730 112.260 37.900 112.405 ;
        RECT 37.275 111.330 37.545 112.235 ;
        RECT 37.730 112.090 38.395 112.260 ;
        RECT 37.715 111.160 38.045 111.920 ;
        RECT 38.225 111.330 38.395 112.090 ;
        RECT 40.250 111.595 40.600 112.845 ;
        RECT 42.080 112.335 42.420 113.165 ;
        RECT 45.770 111.595 46.120 112.845 ;
        RECT 47.600 112.335 47.940 113.165 ;
        RECT 49.785 113.160 49.955 113.540 ;
        RECT 50.135 113.330 50.465 113.710 ;
        RECT 49.785 112.990 50.450 113.160 ;
        RECT 50.645 113.035 50.905 113.540 ;
        RECT 49.715 112.440 50.045 112.810 ;
        RECT 50.280 112.735 50.450 112.990 ;
        RECT 50.280 112.405 50.565 112.735 ;
        RECT 50.280 112.260 50.450 112.405 ;
        RECT 49.785 112.090 50.450 112.260 ;
        RECT 50.735 112.235 50.905 113.035 ;
        RECT 51.075 112.985 51.365 113.710 ;
        RECT 51.535 112.960 52.745 113.710 ;
        RECT 38.660 111.160 44.005 111.595 ;
        RECT 44.180 111.160 49.525 111.595 ;
        RECT 49.785 111.330 49.955 112.090 ;
        RECT 50.135 111.160 50.465 111.920 ;
        RECT 50.635 111.330 50.905 112.235 ;
        RECT 51.075 111.160 51.365 112.325 ;
        RECT 51.535 112.250 52.055 112.790 ;
        RECT 52.225 112.420 52.745 112.960 ;
        RECT 53.005 113.060 53.175 113.540 ;
        RECT 53.355 113.230 53.595 113.710 ;
        RECT 53.845 113.060 54.015 113.540 ;
        RECT 54.185 113.230 54.515 113.710 ;
        RECT 54.685 113.060 54.855 113.540 ;
        RECT 53.005 112.890 53.640 113.060 ;
        RECT 53.845 112.890 54.855 113.060 ;
        RECT 55.025 112.910 55.355 113.710 ;
        RECT 55.675 112.940 57.345 113.710 ;
        RECT 57.520 113.165 62.865 113.710 ;
        RECT 63.040 113.165 68.385 113.710 ;
        RECT 53.470 112.720 53.640 112.890 ;
        RECT 52.920 112.480 53.300 112.720 ;
        RECT 53.470 112.550 53.970 112.720 ;
        RECT 53.470 112.310 53.640 112.550 ;
        RECT 54.360 112.350 54.855 112.890 ;
        RECT 51.535 111.160 52.745 112.250 ;
        RECT 52.925 112.140 53.640 112.310 ;
        RECT 53.845 112.180 54.855 112.350 ;
        RECT 52.925 111.330 53.255 112.140 ;
        RECT 53.425 111.160 53.665 111.960 ;
        RECT 53.845 111.330 54.015 112.180 ;
        RECT 54.185 111.160 54.515 111.960 ;
        RECT 54.685 111.330 54.855 112.180 ;
        RECT 55.025 111.160 55.355 112.310 ;
        RECT 55.675 112.250 56.425 112.770 ;
        RECT 56.595 112.420 57.345 112.940 ;
        RECT 55.675 111.160 57.345 112.250 ;
        RECT 59.110 111.595 59.460 112.845 ;
        RECT 60.940 112.335 61.280 113.165 ;
        RECT 64.630 111.595 64.980 112.845 ;
        RECT 66.460 112.335 66.800 113.165 ;
        RECT 68.645 113.160 68.815 113.540 ;
        RECT 68.995 113.330 69.325 113.710 ;
        RECT 68.645 112.990 69.310 113.160 ;
        RECT 69.505 113.035 69.765 113.540 ;
        RECT 68.575 112.440 68.905 112.810 ;
        RECT 69.140 112.735 69.310 112.990 ;
        RECT 69.140 112.405 69.425 112.735 ;
        RECT 69.140 112.260 69.310 112.405 ;
        RECT 68.645 112.090 69.310 112.260 ;
        RECT 69.595 112.235 69.765 113.035 ;
        RECT 70.025 113.160 70.195 113.540 ;
        RECT 70.375 113.330 70.705 113.710 ;
        RECT 70.025 112.990 70.690 113.160 ;
        RECT 70.885 113.035 71.145 113.540 ;
        RECT 69.955 112.440 70.285 112.810 ;
        RECT 70.520 112.735 70.690 112.990 ;
        RECT 70.520 112.405 70.805 112.735 ;
        RECT 70.520 112.260 70.690 112.405 ;
        RECT 57.520 111.160 62.865 111.595 ;
        RECT 63.040 111.160 68.385 111.595 ;
        RECT 68.645 111.330 68.815 112.090 ;
        RECT 68.995 111.160 69.325 111.920 ;
        RECT 69.495 111.330 69.765 112.235 ;
        RECT 70.025 112.090 70.690 112.260 ;
        RECT 70.975 112.235 71.145 113.035 ;
        RECT 71.405 113.060 71.575 113.540 ;
        RECT 71.755 113.230 71.995 113.710 ;
        RECT 72.245 113.060 72.415 113.540 ;
        RECT 72.585 113.230 72.915 113.710 ;
        RECT 73.085 113.060 73.255 113.540 ;
        RECT 71.405 112.890 72.040 113.060 ;
        RECT 72.245 112.890 73.255 113.060 ;
        RECT 73.425 112.910 73.755 113.710 ;
        RECT 74.075 112.940 76.665 113.710 ;
        RECT 76.835 112.985 77.125 113.710 ;
        RECT 77.755 112.940 79.425 113.710 ;
        RECT 79.600 113.165 84.945 113.710 ;
        RECT 71.870 112.720 72.040 112.890 ;
        RECT 71.320 112.480 71.700 112.720 ;
        RECT 71.870 112.550 72.370 112.720 ;
        RECT 71.870 112.310 72.040 112.550 ;
        RECT 72.760 112.350 73.255 112.890 ;
        RECT 70.025 111.330 70.195 112.090 ;
        RECT 70.375 111.160 70.705 111.920 ;
        RECT 70.875 111.330 71.145 112.235 ;
        RECT 71.325 112.140 72.040 112.310 ;
        RECT 72.245 112.180 73.255 112.350 ;
        RECT 71.325 111.330 71.655 112.140 ;
        RECT 71.825 111.160 72.065 111.960 ;
        RECT 72.245 111.330 72.415 112.180 ;
        RECT 72.585 111.160 72.915 111.960 ;
        RECT 73.085 111.330 73.255 112.180 ;
        RECT 73.425 111.160 73.755 112.310 ;
        RECT 74.075 112.250 75.285 112.770 ;
        RECT 75.455 112.420 76.665 112.940 ;
        RECT 74.075 111.160 76.665 112.250 ;
        RECT 76.835 111.160 77.125 112.325 ;
        RECT 77.755 112.250 78.505 112.770 ;
        RECT 78.675 112.420 79.425 112.940 ;
        RECT 77.755 111.160 79.425 112.250 ;
        RECT 81.190 111.595 81.540 112.845 ;
        RECT 83.020 112.335 83.360 113.165 ;
        RECT 85.205 113.160 85.375 113.540 ;
        RECT 85.555 113.330 85.885 113.710 ;
        RECT 85.205 112.990 85.870 113.160 ;
        RECT 86.065 113.035 86.325 113.540 ;
        RECT 85.135 112.440 85.465 112.810 ;
        RECT 85.700 112.735 85.870 112.990 ;
        RECT 85.700 112.405 85.985 112.735 ;
        RECT 85.700 112.260 85.870 112.405 ;
        RECT 85.205 112.090 85.870 112.260 ;
        RECT 86.155 112.235 86.325 113.035 ;
        RECT 86.495 112.940 90.005 113.710 ;
        RECT 90.265 113.160 90.435 113.540 ;
        RECT 90.615 113.330 90.945 113.710 ;
        RECT 90.265 112.990 90.930 113.160 ;
        RECT 91.125 113.035 91.385 113.540 ;
        RECT 79.600 111.160 84.945 111.595 ;
        RECT 85.205 111.330 85.375 112.090 ;
        RECT 85.555 111.160 85.885 111.920 ;
        RECT 86.055 111.330 86.325 112.235 ;
        RECT 86.495 112.250 88.185 112.770 ;
        RECT 88.355 112.420 90.005 112.940 ;
        RECT 90.195 112.440 90.525 112.810 ;
        RECT 90.760 112.735 90.930 112.990 ;
        RECT 90.760 112.405 91.045 112.735 ;
        RECT 90.760 112.260 90.930 112.405 ;
        RECT 86.495 111.160 90.005 112.250 ;
        RECT 90.265 112.090 90.930 112.260 ;
        RECT 91.215 112.235 91.385 113.035 ;
        RECT 92.015 112.940 95.525 113.710 ;
        RECT 95.785 113.160 95.955 113.540 ;
        RECT 96.135 113.330 96.465 113.710 ;
        RECT 95.785 112.990 96.450 113.160 ;
        RECT 96.645 113.035 96.905 113.540 ;
        RECT 90.265 111.330 90.435 112.090 ;
        RECT 90.615 111.160 90.945 111.920 ;
        RECT 91.115 111.330 91.385 112.235 ;
        RECT 92.015 112.250 93.705 112.770 ;
        RECT 93.875 112.420 95.525 112.940 ;
        RECT 95.715 112.440 96.045 112.810 ;
        RECT 96.280 112.735 96.450 112.990 ;
        RECT 96.280 112.405 96.565 112.735 ;
        RECT 96.280 112.260 96.450 112.405 ;
        RECT 92.015 111.160 95.525 112.250 ;
        RECT 95.785 112.090 96.450 112.260 ;
        RECT 96.735 112.235 96.905 113.035 ;
        RECT 97.075 112.940 99.665 113.710 ;
        RECT 99.925 113.160 100.095 113.540 ;
        RECT 100.275 113.330 100.605 113.710 ;
        RECT 99.925 112.990 100.590 113.160 ;
        RECT 100.785 113.035 101.045 113.540 ;
        RECT 95.785 111.330 95.955 112.090 ;
        RECT 96.135 111.160 96.465 111.920 ;
        RECT 96.635 111.330 96.905 112.235 ;
        RECT 97.075 112.250 98.285 112.770 ;
        RECT 98.455 112.420 99.665 112.940 ;
        RECT 99.855 112.440 100.185 112.810 ;
        RECT 100.420 112.735 100.590 112.990 ;
        RECT 100.420 112.405 100.705 112.735 ;
        RECT 100.420 112.260 100.590 112.405 ;
        RECT 97.075 111.160 99.665 112.250 ;
        RECT 99.925 112.090 100.590 112.260 ;
        RECT 100.875 112.235 101.045 113.035 ;
        RECT 101.305 113.160 101.475 113.540 ;
        RECT 101.655 113.330 101.985 113.710 ;
        RECT 101.305 112.990 101.970 113.160 ;
        RECT 102.165 113.035 102.425 113.540 ;
        RECT 101.235 112.440 101.565 112.810 ;
        RECT 101.800 112.735 101.970 112.990 ;
        RECT 101.800 112.405 102.085 112.735 ;
        RECT 101.800 112.260 101.970 112.405 ;
        RECT 99.925 111.330 100.095 112.090 ;
        RECT 100.275 111.160 100.605 111.920 ;
        RECT 100.775 111.330 101.045 112.235 ;
        RECT 101.305 112.090 101.970 112.260 ;
        RECT 102.255 112.235 102.425 113.035 ;
        RECT 102.595 112.985 102.885 113.710 ;
        RECT 103.980 113.160 104.235 113.450 ;
        RECT 104.405 113.330 104.735 113.710 ;
        RECT 103.980 112.990 104.730 113.160 ;
        RECT 101.305 111.330 101.475 112.090 ;
        RECT 101.655 111.160 101.985 111.920 ;
        RECT 102.155 111.330 102.425 112.235 ;
        RECT 102.595 111.160 102.885 112.325 ;
        RECT 103.980 112.170 104.330 112.820 ;
        RECT 104.500 112.000 104.730 112.990 ;
        RECT 103.980 111.830 104.730 112.000 ;
        RECT 103.980 111.330 104.235 111.830 ;
        RECT 104.405 111.160 104.735 111.660 ;
        RECT 104.905 111.330 105.075 113.450 ;
        RECT 105.435 113.350 105.765 113.710 ;
        RECT 105.935 113.320 106.430 113.490 ;
        RECT 106.635 113.320 107.490 113.490 ;
        RECT 105.305 112.130 105.765 113.180 ;
        RECT 105.245 111.345 105.570 112.130 ;
        RECT 105.935 111.960 106.105 113.320 ;
        RECT 106.275 112.410 106.625 113.030 ;
        RECT 106.795 112.810 107.150 113.030 ;
        RECT 106.795 112.220 106.965 112.810 ;
        RECT 107.320 112.610 107.490 113.320 ;
        RECT 108.365 113.250 108.695 113.710 ;
        RECT 108.905 113.350 109.255 113.520 ;
        RECT 107.695 112.780 108.485 113.030 ;
        RECT 108.905 112.960 109.165 113.350 ;
        RECT 109.475 113.260 110.425 113.540 ;
        RECT 110.595 113.270 110.785 113.710 ;
        RECT 110.955 113.330 112.025 113.500 ;
        RECT 108.655 112.610 108.825 112.790 ;
        RECT 105.935 111.790 106.330 111.960 ;
        RECT 106.500 111.830 106.965 112.220 ;
        RECT 107.135 112.440 108.825 112.610 ;
        RECT 106.160 111.660 106.330 111.790 ;
        RECT 107.135 111.660 107.305 112.440 ;
        RECT 108.995 112.270 109.165 112.960 ;
        RECT 107.665 112.100 109.165 112.270 ;
        RECT 109.355 112.300 109.565 113.090 ;
        RECT 109.735 112.470 110.085 113.090 ;
        RECT 110.255 112.480 110.425 113.260 ;
        RECT 110.955 113.100 111.125 113.330 ;
        RECT 110.595 112.930 111.125 113.100 ;
        RECT 110.595 112.650 110.815 112.930 ;
        RECT 111.295 112.760 111.535 113.160 ;
        RECT 110.255 112.310 110.660 112.480 ;
        RECT 110.995 112.390 111.535 112.760 ;
        RECT 111.705 112.975 112.025 113.330 ;
        RECT 111.705 112.720 112.030 112.975 ;
        RECT 112.225 112.900 112.395 113.710 ;
        RECT 112.565 113.060 112.895 113.540 ;
        RECT 113.065 113.240 113.235 113.710 ;
        RECT 113.405 113.060 113.735 113.540 ;
        RECT 113.905 113.240 114.075 113.710 ;
        RECT 112.565 112.890 114.330 113.060 ;
        RECT 114.555 112.960 115.765 113.710 ;
        RECT 111.705 112.510 113.735 112.720 ;
        RECT 111.705 112.500 112.050 112.510 ;
        RECT 109.355 112.140 110.030 112.300 ;
        RECT 110.490 112.220 110.660 112.310 ;
        RECT 109.355 112.130 110.320 112.140 ;
        RECT 108.995 111.960 109.165 112.100 ;
        RECT 105.740 111.160 105.990 111.620 ;
        RECT 106.160 111.330 106.410 111.660 ;
        RECT 106.625 111.330 107.305 111.660 ;
        RECT 107.475 111.760 108.550 111.930 ;
        RECT 108.995 111.790 109.555 111.960 ;
        RECT 109.860 111.840 110.320 112.130 ;
        RECT 110.490 112.050 111.710 112.220 ;
        RECT 107.475 111.420 107.645 111.760 ;
        RECT 107.880 111.160 108.210 111.590 ;
        RECT 108.380 111.420 108.550 111.760 ;
        RECT 108.845 111.160 109.215 111.620 ;
        RECT 109.385 111.330 109.555 111.790 ;
        RECT 110.490 111.670 110.660 112.050 ;
        RECT 111.880 111.880 112.050 112.500 ;
        RECT 113.920 112.340 114.330 112.890 ;
        RECT 109.790 111.330 110.660 111.670 ;
        RECT 111.250 111.710 112.050 111.880 ;
        RECT 110.830 111.160 111.080 111.620 ;
        RECT 111.250 111.420 111.420 111.710 ;
        RECT 111.600 111.160 111.930 111.540 ;
        RECT 112.225 111.160 112.395 112.220 ;
        RECT 112.605 112.170 114.330 112.340 ;
        RECT 114.555 112.250 115.075 112.790 ;
        RECT 115.245 112.420 115.765 112.960 ;
        RECT 112.605 111.330 112.895 112.170 ;
        RECT 113.065 111.160 113.235 112.000 ;
        RECT 113.445 111.330 113.695 112.170 ;
        RECT 113.905 111.160 114.075 112.000 ;
        RECT 114.555 111.160 115.765 112.250 ;
        RECT 10.510 110.990 115.850 111.160 ;
        RECT 10.595 109.900 11.805 110.990 ;
        RECT 10.595 109.190 11.115 109.730 ;
        RECT 11.285 109.360 11.805 109.900 ;
        RECT 12.435 109.825 12.725 110.990 ;
        RECT 12.895 109.900 14.105 110.990 ;
        RECT 14.585 110.150 14.755 110.990 ;
        RECT 14.965 109.980 15.215 110.820 ;
        RECT 15.425 110.150 15.595 110.990 ;
        RECT 15.765 109.980 16.055 110.820 ;
        RECT 12.895 109.360 13.415 109.900 ;
        RECT 14.330 109.810 16.055 109.980 ;
        RECT 16.265 109.930 16.435 110.990 ;
        RECT 16.730 110.610 17.060 110.990 ;
        RECT 17.240 110.440 17.410 110.730 ;
        RECT 17.580 110.530 17.830 110.990 ;
        RECT 16.610 110.270 17.410 110.440 ;
        RECT 18.000 110.480 18.870 110.820 ;
        RECT 13.585 109.190 14.105 109.730 ;
        RECT 10.595 108.440 11.805 109.190 ;
        RECT 12.435 108.440 12.725 109.165 ;
        RECT 12.895 108.440 14.105 109.190 ;
        RECT 14.330 109.260 14.740 109.810 ;
        RECT 16.610 109.650 16.780 110.270 ;
        RECT 18.000 110.100 18.170 110.480 ;
        RECT 19.105 110.360 19.275 110.820 ;
        RECT 19.445 110.530 19.815 110.990 ;
        RECT 20.110 110.390 20.280 110.730 ;
        RECT 20.450 110.560 20.780 110.990 ;
        RECT 21.015 110.390 21.185 110.730 ;
        RECT 16.950 109.930 18.170 110.100 ;
        RECT 18.340 110.020 18.800 110.310 ;
        RECT 19.105 110.190 19.665 110.360 ;
        RECT 20.110 110.220 21.185 110.390 ;
        RECT 21.355 110.490 22.035 110.820 ;
        RECT 22.250 110.490 22.500 110.820 ;
        RECT 22.670 110.530 22.920 110.990 ;
        RECT 19.495 110.050 19.665 110.190 ;
        RECT 18.340 110.010 19.305 110.020 ;
        RECT 18.000 109.840 18.170 109.930 ;
        RECT 18.630 109.850 19.305 110.010 ;
        RECT 16.610 109.640 16.955 109.650 ;
        RECT 14.925 109.430 16.955 109.640 ;
        RECT 14.330 109.090 16.095 109.260 ;
        RECT 14.585 108.440 14.755 108.910 ;
        RECT 14.925 108.610 15.255 109.090 ;
        RECT 15.425 108.440 15.595 108.910 ;
        RECT 15.765 108.610 16.095 109.090 ;
        RECT 16.265 108.440 16.435 109.250 ;
        RECT 16.630 109.175 16.955 109.430 ;
        RECT 16.635 108.820 16.955 109.175 ;
        RECT 17.125 109.390 17.665 109.760 ;
        RECT 18.000 109.670 18.405 109.840 ;
        RECT 17.125 108.990 17.365 109.390 ;
        RECT 17.845 109.220 18.065 109.500 ;
        RECT 17.535 109.050 18.065 109.220 ;
        RECT 17.535 108.820 17.705 109.050 ;
        RECT 18.235 108.890 18.405 109.670 ;
        RECT 18.575 109.060 18.925 109.680 ;
        RECT 19.095 109.060 19.305 109.850 ;
        RECT 19.495 109.880 20.995 110.050 ;
        RECT 19.495 109.190 19.665 109.880 ;
        RECT 21.355 109.710 21.525 110.490 ;
        RECT 22.330 110.360 22.500 110.490 ;
        RECT 19.835 109.540 21.525 109.710 ;
        RECT 21.695 109.930 22.160 110.320 ;
        RECT 22.330 110.190 22.725 110.360 ;
        RECT 19.835 109.360 20.005 109.540 ;
        RECT 16.635 108.650 17.705 108.820 ;
        RECT 17.875 108.440 18.065 108.880 ;
        RECT 18.235 108.610 19.185 108.890 ;
        RECT 19.495 108.800 19.755 109.190 ;
        RECT 20.175 109.120 20.965 109.370 ;
        RECT 19.405 108.630 19.755 108.800 ;
        RECT 19.965 108.440 20.295 108.900 ;
        RECT 21.170 108.830 21.340 109.540 ;
        RECT 21.695 109.340 21.865 109.930 ;
        RECT 21.510 109.120 21.865 109.340 ;
        RECT 22.035 109.120 22.385 109.740 ;
        RECT 22.555 108.830 22.725 110.190 ;
        RECT 23.090 110.020 23.415 110.805 ;
        RECT 22.895 108.970 23.355 110.020 ;
        RECT 21.170 108.660 22.025 108.830 ;
        RECT 22.230 108.660 22.725 108.830 ;
        RECT 22.895 108.440 23.225 108.800 ;
        RECT 23.585 108.700 23.755 110.820 ;
        RECT 23.925 110.490 24.255 110.990 ;
        RECT 24.425 110.320 24.680 110.820 ;
        RECT 23.930 110.150 24.680 110.320 ;
        RECT 23.930 109.160 24.160 110.150 ;
        RECT 24.330 109.330 24.680 109.980 ;
        RECT 24.855 109.915 25.125 110.820 ;
        RECT 25.295 110.230 25.625 110.990 ;
        RECT 25.805 110.060 25.975 110.820 ;
        RECT 23.930 108.990 24.680 109.160 ;
        RECT 23.925 108.440 24.255 108.820 ;
        RECT 24.425 108.700 24.680 108.990 ;
        RECT 24.855 109.115 25.025 109.915 ;
        RECT 25.310 109.890 25.975 110.060 ;
        RECT 26.235 109.915 26.505 110.820 ;
        RECT 26.675 110.230 27.005 110.990 ;
        RECT 27.185 110.060 27.355 110.820 ;
        RECT 27.925 110.150 28.095 110.990 ;
        RECT 25.310 109.745 25.480 109.890 ;
        RECT 25.195 109.415 25.480 109.745 ;
        RECT 25.310 109.160 25.480 109.415 ;
        RECT 25.715 109.340 26.045 109.710 ;
        RECT 24.855 108.610 25.115 109.115 ;
        RECT 25.310 108.990 25.975 109.160 ;
        RECT 25.295 108.440 25.625 108.820 ;
        RECT 25.805 108.610 25.975 108.990 ;
        RECT 26.235 109.115 26.405 109.915 ;
        RECT 26.690 109.890 27.355 110.060 ;
        RECT 28.305 109.980 28.555 110.820 ;
        RECT 28.765 110.150 28.935 110.990 ;
        RECT 29.105 109.980 29.395 110.820 ;
        RECT 26.690 109.745 26.860 109.890 ;
        RECT 26.575 109.415 26.860 109.745 ;
        RECT 27.670 109.810 29.395 109.980 ;
        RECT 29.605 109.930 29.775 110.990 ;
        RECT 30.070 110.610 30.400 110.990 ;
        RECT 30.580 110.440 30.750 110.730 ;
        RECT 30.920 110.530 31.170 110.990 ;
        RECT 29.950 110.270 30.750 110.440 ;
        RECT 31.340 110.480 32.210 110.820 ;
        RECT 26.690 109.160 26.860 109.415 ;
        RECT 27.095 109.340 27.425 109.710 ;
        RECT 27.670 109.260 28.080 109.810 ;
        RECT 29.950 109.650 30.120 110.270 ;
        RECT 31.340 110.100 31.510 110.480 ;
        RECT 32.445 110.360 32.615 110.820 ;
        RECT 32.785 110.530 33.155 110.990 ;
        RECT 33.450 110.390 33.620 110.730 ;
        RECT 33.790 110.560 34.120 110.990 ;
        RECT 34.355 110.390 34.525 110.730 ;
        RECT 30.290 109.930 31.510 110.100 ;
        RECT 31.680 110.020 32.140 110.310 ;
        RECT 32.445 110.190 33.005 110.360 ;
        RECT 33.450 110.220 34.525 110.390 ;
        RECT 34.695 110.490 35.375 110.820 ;
        RECT 35.590 110.490 35.840 110.820 ;
        RECT 36.010 110.530 36.260 110.990 ;
        RECT 32.835 110.050 33.005 110.190 ;
        RECT 31.680 110.010 32.645 110.020 ;
        RECT 31.340 109.840 31.510 109.930 ;
        RECT 31.970 109.850 32.645 110.010 ;
        RECT 29.950 109.640 30.295 109.650 ;
        RECT 28.265 109.430 30.295 109.640 ;
        RECT 26.235 108.610 26.495 109.115 ;
        RECT 26.690 108.990 27.355 109.160 ;
        RECT 27.670 109.090 29.435 109.260 ;
        RECT 26.675 108.440 27.005 108.820 ;
        RECT 27.185 108.610 27.355 108.990 ;
        RECT 27.925 108.440 28.095 108.910 ;
        RECT 28.265 108.610 28.595 109.090 ;
        RECT 28.765 108.440 28.935 108.910 ;
        RECT 29.105 108.610 29.435 109.090 ;
        RECT 29.605 108.440 29.775 109.250 ;
        RECT 29.970 109.175 30.295 109.430 ;
        RECT 29.975 108.820 30.295 109.175 ;
        RECT 30.465 109.390 31.005 109.760 ;
        RECT 31.340 109.670 31.745 109.840 ;
        RECT 30.465 108.990 30.705 109.390 ;
        RECT 31.185 109.220 31.405 109.500 ;
        RECT 30.875 109.050 31.405 109.220 ;
        RECT 30.875 108.820 31.045 109.050 ;
        RECT 31.575 108.890 31.745 109.670 ;
        RECT 31.915 109.060 32.265 109.680 ;
        RECT 32.435 109.060 32.645 109.850 ;
        RECT 32.835 109.880 34.335 110.050 ;
        RECT 32.835 109.190 33.005 109.880 ;
        RECT 34.695 109.710 34.865 110.490 ;
        RECT 35.670 110.360 35.840 110.490 ;
        RECT 33.175 109.540 34.865 109.710 ;
        RECT 35.035 109.930 35.500 110.320 ;
        RECT 35.670 110.190 36.065 110.360 ;
        RECT 33.175 109.360 33.345 109.540 ;
        RECT 29.975 108.650 31.045 108.820 ;
        RECT 31.215 108.440 31.405 108.880 ;
        RECT 31.575 108.610 32.525 108.890 ;
        RECT 32.835 108.800 33.095 109.190 ;
        RECT 33.515 109.120 34.305 109.370 ;
        RECT 32.745 108.630 33.095 108.800 ;
        RECT 33.305 108.440 33.635 108.900 ;
        RECT 34.510 108.830 34.680 109.540 ;
        RECT 35.035 109.340 35.205 109.930 ;
        RECT 34.850 109.120 35.205 109.340 ;
        RECT 35.375 109.120 35.725 109.740 ;
        RECT 35.895 108.830 36.065 110.190 ;
        RECT 36.430 110.020 36.755 110.805 ;
        RECT 36.235 108.970 36.695 110.020 ;
        RECT 34.510 108.660 35.365 108.830 ;
        RECT 35.570 108.660 36.065 108.830 ;
        RECT 36.235 108.440 36.565 108.800 ;
        RECT 36.925 108.700 37.095 110.820 ;
        RECT 37.265 110.490 37.595 110.990 ;
        RECT 37.765 110.320 38.020 110.820 ;
        RECT 37.270 110.150 38.020 110.320 ;
        RECT 37.270 109.160 37.500 110.150 ;
        RECT 37.670 109.330 38.020 109.980 ;
        RECT 38.195 109.825 38.485 110.990 ;
        RECT 39.635 109.850 39.845 110.990 ;
        RECT 40.015 109.840 40.345 110.820 ;
        RECT 40.515 109.850 40.745 110.990 ;
        RECT 41.415 109.915 41.685 110.820 ;
        RECT 41.855 110.230 42.185 110.990 ;
        RECT 42.365 110.060 42.535 110.820 ;
        RECT 37.270 108.990 38.020 109.160 ;
        RECT 37.265 108.440 37.595 108.820 ;
        RECT 37.765 108.700 38.020 108.990 ;
        RECT 38.195 108.440 38.485 109.165 ;
        RECT 39.635 108.440 39.845 109.260 ;
        RECT 40.015 109.240 40.265 109.840 ;
        RECT 40.435 109.430 40.765 109.680 ;
        RECT 40.015 108.610 40.345 109.240 ;
        RECT 40.515 108.440 40.745 109.260 ;
        RECT 41.415 109.115 41.585 109.915 ;
        RECT 41.870 109.890 42.535 110.060 ;
        RECT 42.795 109.900 44.465 110.990 ;
        RECT 44.725 110.060 44.895 110.820 ;
        RECT 45.075 110.230 45.405 110.990 ;
        RECT 41.870 109.745 42.040 109.890 ;
        RECT 41.755 109.415 42.040 109.745 ;
        RECT 41.870 109.160 42.040 109.415 ;
        RECT 42.275 109.340 42.605 109.710 ;
        RECT 42.795 109.380 43.545 109.900 ;
        RECT 44.725 109.890 45.390 110.060 ;
        RECT 45.575 109.915 45.845 110.820 ;
        RECT 46.325 110.150 46.495 110.990 ;
        RECT 46.705 109.980 46.955 110.820 ;
        RECT 47.165 110.150 47.335 110.990 ;
        RECT 47.505 109.980 47.795 110.820 ;
        RECT 45.220 109.745 45.390 109.890 ;
        RECT 43.715 109.210 44.465 109.730 ;
        RECT 44.655 109.340 44.985 109.710 ;
        RECT 45.220 109.415 45.505 109.745 ;
        RECT 41.415 108.610 41.675 109.115 ;
        RECT 41.870 108.990 42.535 109.160 ;
        RECT 41.855 108.440 42.185 108.820 ;
        RECT 42.365 108.610 42.535 108.990 ;
        RECT 42.795 108.440 44.465 109.210 ;
        RECT 45.220 109.160 45.390 109.415 ;
        RECT 44.725 108.990 45.390 109.160 ;
        RECT 45.675 109.115 45.845 109.915 ;
        RECT 44.725 108.610 44.895 108.990 ;
        RECT 45.075 108.440 45.405 108.820 ;
        RECT 45.585 108.610 45.845 109.115 ;
        RECT 46.070 109.810 47.795 109.980 ;
        RECT 48.005 109.930 48.175 110.990 ;
        RECT 48.470 110.610 48.800 110.990 ;
        RECT 48.980 110.440 49.150 110.730 ;
        RECT 49.320 110.530 49.570 110.990 ;
        RECT 48.350 110.270 49.150 110.440 ;
        RECT 49.740 110.480 50.610 110.820 ;
        RECT 46.070 109.260 46.480 109.810 ;
        RECT 48.350 109.650 48.520 110.270 ;
        RECT 49.740 110.100 49.910 110.480 ;
        RECT 50.845 110.360 51.015 110.820 ;
        RECT 51.185 110.530 51.555 110.990 ;
        RECT 51.850 110.390 52.020 110.730 ;
        RECT 52.190 110.560 52.520 110.990 ;
        RECT 52.755 110.390 52.925 110.730 ;
        RECT 48.690 109.930 49.910 110.100 ;
        RECT 50.080 110.020 50.540 110.310 ;
        RECT 50.845 110.190 51.405 110.360 ;
        RECT 51.850 110.220 52.925 110.390 ;
        RECT 53.095 110.490 53.775 110.820 ;
        RECT 53.990 110.490 54.240 110.820 ;
        RECT 54.410 110.530 54.660 110.990 ;
        RECT 51.235 110.050 51.405 110.190 ;
        RECT 50.080 110.010 51.045 110.020 ;
        RECT 49.740 109.840 49.910 109.930 ;
        RECT 50.370 109.850 51.045 110.010 ;
        RECT 48.350 109.640 48.695 109.650 ;
        RECT 46.665 109.430 48.695 109.640 ;
        RECT 46.070 109.090 47.835 109.260 ;
        RECT 46.325 108.440 46.495 108.910 ;
        RECT 46.665 108.610 46.995 109.090 ;
        RECT 47.165 108.440 47.335 108.910 ;
        RECT 47.505 108.610 47.835 109.090 ;
        RECT 48.005 108.440 48.175 109.250 ;
        RECT 48.370 109.175 48.695 109.430 ;
        RECT 48.375 108.820 48.695 109.175 ;
        RECT 48.865 109.390 49.405 109.760 ;
        RECT 49.740 109.670 50.145 109.840 ;
        RECT 48.865 108.990 49.105 109.390 ;
        RECT 49.585 109.220 49.805 109.500 ;
        RECT 49.275 109.050 49.805 109.220 ;
        RECT 49.275 108.820 49.445 109.050 ;
        RECT 49.975 108.890 50.145 109.670 ;
        RECT 50.315 109.060 50.665 109.680 ;
        RECT 50.835 109.060 51.045 109.850 ;
        RECT 51.235 109.880 52.735 110.050 ;
        RECT 51.235 109.190 51.405 109.880 ;
        RECT 53.095 109.710 53.265 110.490 ;
        RECT 54.070 110.360 54.240 110.490 ;
        RECT 51.575 109.540 53.265 109.710 ;
        RECT 53.435 109.930 53.900 110.320 ;
        RECT 54.070 110.190 54.465 110.360 ;
        RECT 51.575 109.360 51.745 109.540 ;
        RECT 48.375 108.650 49.445 108.820 ;
        RECT 49.615 108.440 49.805 108.880 ;
        RECT 49.975 108.610 50.925 108.890 ;
        RECT 51.235 108.800 51.495 109.190 ;
        RECT 51.915 109.120 52.705 109.370 ;
        RECT 51.145 108.630 51.495 108.800 ;
        RECT 51.705 108.440 52.035 108.900 ;
        RECT 52.910 108.830 53.080 109.540 ;
        RECT 53.435 109.340 53.605 109.930 ;
        RECT 53.250 109.120 53.605 109.340 ;
        RECT 53.775 109.120 54.125 109.740 ;
        RECT 54.295 108.830 54.465 110.190 ;
        RECT 54.830 110.020 55.155 110.805 ;
        RECT 54.635 108.970 55.095 110.020 ;
        RECT 52.910 108.660 53.765 108.830 ;
        RECT 53.970 108.660 54.465 108.830 ;
        RECT 54.635 108.440 54.965 108.800 ;
        RECT 55.325 108.700 55.495 110.820 ;
        RECT 55.665 110.490 55.995 110.990 ;
        RECT 56.165 110.320 56.420 110.820 ;
        RECT 55.670 110.150 56.420 110.320 ;
        RECT 55.670 109.160 55.900 110.150 ;
        RECT 57.145 110.060 57.315 110.820 ;
        RECT 57.495 110.230 57.825 110.990 ;
        RECT 56.070 109.330 56.420 109.980 ;
        RECT 57.145 109.890 57.810 110.060 ;
        RECT 57.995 109.915 58.265 110.820 ;
        RECT 57.640 109.745 57.810 109.890 ;
        RECT 57.075 109.340 57.405 109.710 ;
        RECT 57.640 109.415 57.925 109.745 ;
        RECT 57.640 109.160 57.810 109.415 ;
        RECT 55.670 108.990 56.420 109.160 ;
        RECT 55.665 108.440 55.995 108.820 ;
        RECT 56.165 108.700 56.420 108.990 ;
        RECT 57.145 108.990 57.810 109.160 ;
        RECT 58.095 109.115 58.265 109.915 ;
        RECT 58.475 109.850 58.705 110.990 ;
        RECT 58.875 109.840 59.205 110.820 ;
        RECT 59.375 109.850 59.585 110.990 ;
        RECT 59.815 109.900 61.025 110.990 ;
        RECT 61.285 110.060 61.455 110.820 ;
        RECT 61.635 110.230 61.965 110.990 ;
        RECT 58.455 109.430 58.785 109.680 ;
        RECT 57.145 108.610 57.315 108.990 ;
        RECT 57.495 108.440 57.825 108.820 ;
        RECT 58.005 108.610 58.265 109.115 ;
        RECT 58.475 108.440 58.705 109.260 ;
        RECT 58.955 109.240 59.205 109.840 ;
        RECT 59.815 109.360 60.335 109.900 ;
        RECT 61.285 109.890 61.950 110.060 ;
        RECT 62.135 109.915 62.405 110.820 ;
        RECT 61.780 109.745 61.950 109.890 ;
        RECT 58.875 108.610 59.205 109.240 ;
        RECT 59.375 108.440 59.585 109.260 ;
        RECT 60.505 109.190 61.025 109.730 ;
        RECT 61.215 109.340 61.545 109.710 ;
        RECT 61.780 109.415 62.065 109.745 ;
        RECT 59.815 108.440 61.025 109.190 ;
        RECT 61.780 109.160 61.950 109.415 ;
        RECT 61.285 108.990 61.950 109.160 ;
        RECT 62.235 109.115 62.405 109.915 ;
        RECT 62.575 109.900 63.785 110.990 ;
        RECT 62.575 109.360 63.095 109.900 ;
        RECT 63.955 109.825 64.245 110.990 ;
        RECT 64.965 110.060 65.135 110.820 ;
        RECT 65.315 110.230 65.645 110.990 ;
        RECT 64.965 109.890 65.630 110.060 ;
        RECT 65.815 109.915 66.085 110.820 ;
        RECT 65.460 109.745 65.630 109.890 ;
        RECT 63.265 109.190 63.785 109.730 ;
        RECT 64.895 109.340 65.225 109.710 ;
        RECT 65.460 109.415 65.745 109.745 ;
        RECT 61.285 108.610 61.455 108.990 ;
        RECT 61.635 108.440 61.965 108.820 ;
        RECT 62.145 108.610 62.405 109.115 ;
        RECT 62.575 108.440 63.785 109.190 ;
        RECT 63.955 108.440 64.245 109.165 ;
        RECT 65.460 109.160 65.630 109.415 ;
        RECT 64.965 108.990 65.630 109.160 ;
        RECT 65.915 109.115 66.085 109.915 ;
        RECT 66.315 109.850 66.525 110.990 ;
        RECT 66.695 109.840 67.025 110.820 ;
        RECT 67.195 109.850 67.425 110.990 ;
        RECT 67.640 110.320 67.895 110.820 ;
        RECT 68.065 110.490 68.395 110.990 ;
        RECT 67.640 110.150 68.390 110.320 ;
        RECT 64.965 108.610 65.135 108.990 ;
        RECT 65.315 108.440 65.645 108.820 ;
        RECT 65.825 108.610 66.085 109.115 ;
        RECT 66.315 108.440 66.525 109.260 ;
        RECT 66.695 109.240 66.945 109.840 ;
        RECT 67.115 109.430 67.445 109.680 ;
        RECT 67.640 109.330 67.990 109.980 ;
        RECT 66.695 108.610 67.025 109.240 ;
        RECT 67.195 108.440 67.425 109.260 ;
        RECT 68.160 109.160 68.390 110.150 ;
        RECT 67.640 108.990 68.390 109.160 ;
        RECT 67.640 108.700 67.895 108.990 ;
        RECT 68.065 108.440 68.395 108.820 ;
        RECT 68.565 108.700 68.735 110.820 ;
        RECT 68.905 110.020 69.230 110.805 ;
        RECT 69.400 110.530 69.650 110.990 ;
        RECT 69.820 110.490 70.070 110.820 ;
        RECT 70.285 110.490 70.965 110.820 ;
        RECT 69.820 110.360 69.990 110.490 ;
        RECT 69.595 110.190 69.990 110.360 ;
        RECT 68.965 108.970 69.425 110.020 ;
        RECT 69.595 108.830 69.765 110.190 ;
        RECT 70.160 109.930 70.625 110.320 ;
        RECT 69.935 109.120 70.285 109.740 ;
        RECT 70.455 109.340 70.625 109.930 ;
        RECT 70.795 109.710 70.965 110.490 ;
        RECT 71.135 110.390 71.305 110.730 ;
        RECT 71.540 110.560 71.870 110.990 ;
        RECT 72.040 110.390 72.210 110.730 ;
        RECT 72.505 110.530 72.875 110.990 ;
        RECT 71.135 110.220 72.210 110.390 ;
        RECT 73.045 110.360 73.215 110.820 ;
        RECT 73.450 110.480 74.320 110.820 ;
        RECT 74.490 110.530 74.740 110.990 ;
        RECT 72.655 110.190 73.215 110.360 ;
        RECT 72.655 110.050 72.825 110.190 ;
        RECT 71.325 109.880 72.825 110.050 ;
        RECT 73.520 110.020 73.980 110.310 ;
        RECT 70.795 109.540 72.485 109.710 ;
        RECT 70.455 109.120 70.810 109.340 ;
        RECT 70.980 108.830 71.150 109.540 ;
        RECT 71.355 109.120 72.145 109.370 ;
        RECT 72.315 109.360 72.485 109.540 ;
        RECT 72.655 109.190 72.825 109.880 ;
        RECT 69.095 108.440 69.425 108.800 ;
        RECT 69.595 108.660 70.090 108.830 ;
        RECT 70.295 108.660 71.150 108.830 ;
        RECT 72.025 108.440 72.355 108.900 ;
        RECT 72.565 108.800 72.825 109.190 ;
        RECT 73.015 110.010 73.980 110.020 ;
        RECT 74.150 110.100 74.320 110.480 ;
        RECT 74.910 110.440 75.080 110.730 ;
        RECT 75.260 110.610 75.590 110.990 ;
        RECT 74.910 110.270 75.710 110.440 ;
        RECT 73.015 109.850 73.690 110.010 ;
        RECT 74.150 109.930 75.370 110.100 ;
        RECT 73.015 109.060 73.225 109.850 ;
        RECT 74.150 109.840 74.320 109.930 ;
        RECT 73.395 109.060 73.745 109.680 ;
        RECT 73.915 109.670 74.320 109.840 ;
        RECT 73.915 108.890 74.085 109.670 ;
        RECT 74.255 109.220 74.475 109.500 ;
        RECT 74.655 109.390 75.195 109.760 ;
        RECT 75.540 109.650 75.710 110.270 ;
        RECT 75.885 109.930 76.055 110.990 ;
        RECT 76.265 109.980 76.555 110.820 ;
        RECT 76.725 110.150 76.895 110.990 ;
        RECT 77.105 109.980 77.355 110.820 ;
        RECT 77.565 110.150 77.735 110.990 ;
        RECT 79.445 110.150 79.615 110.990 ;
        RECT 79.825 109.980 80.075 110.820 ;
        RECT 80.285 110.150 80.455 110.990 ;
        RECT 80.625 109.980 80.915 110.820 ;
        RECT 76.265 109.810 77.990 109.980 ;
        RECT 74.255 109.050 74.785 109.220 ;
        RECT 72.565 108.630 72.915 108.800 ;
        RECT 73.135 108.610 74.085 108.890 ;
        RECT 74.255 108.440 74.445 108.880 ;
        RECT 74.615 108.820 74.785 109.050 ;
        RECT 74.955 108.990 75.195 109.390 ;
        RECT 75.365 109.640 75.710 109.650 ;
        RECT 75.365 109.430 77.395 109.640 ;
        RECT 75.365 109.175 75.690 109.430 ;
        RECT 77.580 109.260 77.990 109.810 ;
        RECT 75.365 108.820 75.685 109.175 ;
        RECT 74.615 108.650 75.685 108.820 ;
        RECT 75.885 108.440 76.055 109.250 ;
        RECT 76.225 109.090 77.990 109.260 ;
        RECT 79.190 109.810 80.915 109.980 ;
        RECT 81.125 109.930 81.295 110.990 ;
        RECT 81.590 110.610 81.920 110.990 ;
        RECT 82.100 110.440 82.270 110.730 ;
        RECT 82.440 110.530 82.690 110.990 ;
        RECT 81.470 110.270 82.270 110.440 ;
        RECT 82.860 110.480 83.730 110.820 ;
        RECT 79.190 109.260 79.600 109.810 ;
        RECT 81.470 109.650 81.640 110.270 ;
        RECT 82.860 110.100 83.030 110.480 ;
        RECT 83.965 110.360 84.135 110.820 ;
        RECT 84.305 110.530 84.675 110.990 ;
        RECT 84.970 110.390 85.140 110.730 ;
        RECT 85.310 110.560 85.640 110.990 ;
        RECT 85.875 110.390 86.045 110.730 ;
        RECT 81.810 109.930 83.030 110.100 ;
        RECT 83.200 110.020 83.660 110.310 ;
        RECT 83.965 110.190 84.525 110.360 ;
        RECT 84.970 110.220 86.045 110.390 ;
        RECT 86.215 110.490 86.895 110.820 ;
        RECT 87.110 110.490 87.360 110.820 ;
        RECT 87.530 110.530 87.780 110.990 ;
        RECT 84.355 110.050 84.525 110.190 ;
        RECT 83.200 110.010 84.165 110.020 ;
        RECT 82.860 109.840 83.030 109.930 ;
        RECT 83.490 109.850 84.165 110.010 ;
        RECT 81.470 109.640 81.815 109.650 ;
        RECT 79.785 109.430 81.815 109.640 ;
        RECT 79.190 109.090 80.955 109.260 ;
        RECT 76.225 108.610 76.555 109.090 ;
        RECT 76.725 108.440 76.895 108.910 ;
        RECT 77.065 108.610 77.395 109.090 ;
        RECT 77.565 108.440 77.735 108.910 ;
        RECT 79.445 108.440 79.615 108.910 ;
        RECT 79.785 108.610 80.115 109.090 ;
        RECT 80.285 108.440 80.455 108.910 ;
        RECT 80.625 108.610 80.955 109.090 ;
        RECT 81.125 108.440 81.295 109.250 ;
        RECT 81.490 109.175 81.815 109.430 ;
        RECT 81.495 108.820 81.815 109.175 ;
        RECT 81.985 109.390 82.525 109.760 ;
        RECT 82.860 109.670 83.265 109.840 ;
        RECT 81.985 108.990 82.225 109.390 ;
        RECT 82.705 109.220 82.925 109.500 ;
        RECT 82.395 109.050 82.925 109.220 ;
        RECT 82.395 108.820 82.565 109.050 ;
        RECT 83.095 108.890 83.265 109.670 ;
        RECT 83.435 109.060 83.785 109.680 ;
        RECT 83.955 109.060 84.165 109.850 ;
        RECT 84.355 109.880 85.855 110.050 ;
        RECT 84.355 109.190 84.525 109.880 ;
        RECT 86.215 109.710 86.385 110.490 ;
        RECT 87.190 110.360 87.360 110.490 ;
        RECT 84.695 109.540 86.385 109.710 ;
        RECT 86.555 109.930 87.020 110.320 ;
        RECT 87.190 110.190 87.585 110.360 ;
        RECT 84.695 109.360 84.865 109.540 ;
        RECT 81.495 108.650 82.565 108.820 ;
        RECT 82.735 108.440 82.925 108.880 ;
        RECT 83.095 108.610 84.045 108.890 ;
        RECT 84.355 108.800 84.615 109.190 ;
        RECT 85.035 109.120 85.825 109.370 ;
        RECT 84.265 108.630 84.615 108.800 ;
        RECT 84.825 108.440 85.155 108.900 ;
        RECT 86.030 108.830 86.200 109.540 ;
        RECT 86.555 109.340 86.725 109.930 ;
        RECT 86.370 109.120 86.725 109.340 ;
        RECT 86.895 109.120 87.245 109.740 ;
        RECT 87.415 108.830 87.585 110.190 ;
        RECT 87.950 110.020 88.275 110.805 ;
        RECT 87.755 108.970 88.215 110.020 ;
        RECT 86.030 108.660 86.885 108.830 ;
        RECT 87.090 108.660 87.585 108.830 ;
        RECT 87.755 108.440 88.085 108.800 ;
        RECT 88.445 108.700 88.615 110.820 ;
        RECT 88.785 110.490 89.115 110.990 ;
        RECT 89.285 110.320 89.540 110.820 ;
        RECT 88.790 110.150 89.540 110.320 ;
        RECT 88.790 109.160 89.020 110.150 ;
        RECT 89.190 109.330 89.540 109.980 ;
        RECT 89.715 109.825 90.005 110.990 ;
        RECT 90.485 110.150 90.655 110.990 ;
        RECT 90.865 109.980 91.115 110.820 ;
        RECT 91.325 110.150 91.495 110.990 ;
        RECT 91.665 109.980 91.955 110.820 ;
        RECT 90.230 109.810 91.955 109.980 ;
        RECT 92.165 109.930 92.335 110.990 ;
        RECT 92.630 110.610 92.960 110.990 ;
        RECT 93.140 110.440 93.310 110.730 ;
        RECT 93.480 110.530 93.730 110.990 ;
        RECT 92.510 110.270 93.310 110.440 ;
        RECT 93.900 110.480 94.770 110.820 ;
        RECT 90.230 109.260 90.640 109.810 ;
        RECT 92.510 109.650 92.680 110.270 ;
        RECT 93.900 110.100 94.070 110.480 ;
        RECT 95.005 110.360 95.175 110.820 ;
        RECT 95.345 110.530 95.715 110.990 ;
        RECT 96.010 110.390 96.180 110.730 ;
        RECT 96.350 110.560 96.680 110.990 ;
        RECT 96.915 110.390 97.085 110.730 ;
        RECT 92.850 109.930 94.070 110.100 ;
        RECT 94.240 110.020 94.700 110.310 ;
        RECT 95.005 110.190 95.565 110.360 ;
        RECT 96.010 110.220 97.085 110.390 ;
        RECT 97.255 110.490 97.935 110.820 ;
        RECT 98.150 110.490 98.400 110.820 ;
        RECT 98.570 110.530 98.820 110.990 ;
        RECT 95.395 110.050 95.565 110.190 ;
        RECT 94.240 110.010 95.205 110.020 ;
        RECT 93.900 109.840 94.070 109.930 ;
        RECT 94.530 109.850 95.205 110.010 ;
        RECT 92.510 109.640 92.855 109.650 ;
        RECT 90.825 109.430 92.855 109.640 ;
        RECT 88.790 108.990 89.540 109.160 ;
        RECT 88.785 108.440 89.115 108.820 ;
        RECT 89.285 108.700 89.540 108.990 ;
        RECT 89.715 108.440 90.005 109.165 ;
        RECT 90.230 109.090 91.995 109.260 ;
        RECT 90.485 108.440 90.655 108.910 ;
        RECT 90.825 108.610 91.155 109.090 ;
        RECT 91.325 108.440 91.495 108.910 ;
        RECT 91.665 108.610 91.995 109.090 ;
        RECT 92.165 108.440 92.335 109.250 ;
        RECT 92.530 109.175 92.855 109.430 ;
        RECT 92.535 108.820 92.855 109.175 ;
        RECT 93.025 109.390 93.565 109.760 ;
        RECT 93.900 109.670 94.305 109.840 ;
        RECT 93.025 108.990 93.265 109.390 ;
        RECT 93.745 109.220 93.965 109.500 ;
        RECT 93.435 109.050 93.965 109.220 ;
        RECT 93.435 108.820 93.605 109.050 ;
        RECT 94.135 108.890 94.305 109.670 ;
        RECT 94.475 109.060 94.825 109.680 ;
        RECT 94.995 109.060 95.205 109.850 ;
        RECT 95.395 109.880 96.895 110.050 ;
        RECT 95.395 109.190 95.565 109.880 ;
        RECT 97.255 109.710 97.425 110.490 ;
        RECT 98.230 110.360 98.400 110.490 ;
        RECT 95.735 109.540 97.425 109.710 ;
        RECT 97.595 109.930 98.060 110.320 ;
        RECT 98.230 110.190 98.625 110.360 ;
        RECT 95.735 109.360 95.905 109.540 ;
        RECT 92.535 108.650 93.605 108.820 ;
        RECT 93.775 108.440 93.965 108.880 ;
        RECT 94.135 108.610 95.085 108.890 ;
        RECT 95.395 108.800 95.655 109.190 ;
        RECT 96.075 109.120 96.865 109.370 ;
        RECT 95.305 108.630 95.655 108.800 ;
        RECT 95.865 108.440 96.195 108.900 ;
        RECT 97.070 108.830 97.240 109.540 ;
        RECT 97.595 109.340 97.765 109.930 ;
        RECT 97.410 109.120 97.765 109.340 ;
        RECT 97.935 109.120 98.285 109.740 ;
        RECT 98.455 108.830 98.625 110.190 ;
        RECT 98.990 110.020 99.315 110.805 ;
        RECT 98.795 108.970 99.255 110.020 ;
        RECT 97.070 108.660 97.925 108.830 ;
        RECT 98.130 108.660 98.625 108.830 ;
        RECT 98.795 108.440 99.125 108.800 ;
        RECT 99.485 108.700 99.655 110.820 ;
        RECT 99.825 110.490 100.155 110.990 ;
        RECT 100.325 110.320 100.580 110.820 ;
        RECT 99.830 110.150 100.580 110.320 ;
        RECT 99.830 109.160 100.060 110.150 ;
        RECT 100.230 109.330 100.580 109.980 ;
        RECT 101.215 109.900 103.805 110.990 ;
        RECT 103.980 110.320 104.235 110.820 ;
        RECT 104.405 110.490 104.735 110.990 ;
        RECT 103.980 110.150 104.730 110.320 ;
        RECT 101.215 109.380 102.425 109.900 ;
        RECT 102.595 109.210 103.805 109.730 ;
        RECT 103.980 109.330 104.330 109.980 ;
        RECT 99.830 108.990 100.580 109.160 ;
        RECT 99.825 108.440 100.155 108.820 ;
        RECT 100.325 108.700 100.580 108.990 ;
        RECT 101.215 108.440 103.805 109.210 ;
        RECT 104.500 109.160 104.730 110.150 ;
        RECT 103.980 108.990 104.730 109.160 ;
        RECT 103.980 108.700 104.235 108.990 ;
        RECT 104.405 108.440 104.735 108.820 ;
        RECT 104.905 108.700 105.075 110.820 ;
        RECT 105.245 110.020 105.570 110.805 ;
        RECT 105.740 110.530 105.990 110.990 ;
        RECT 106.160 110.490 106.410 110.820 ;
        RECT 106.625 110.490 107.305 110.820 ;
        RECT 106.160 110.360 106.330 110.490 ;
        RECT 105.935 110.190 106.330 110.360 ;
        RECT 105.305 108.970 105.765 110.020 ;
        RECT 105.935 108.830 106.105 110.190 ;
        RECT 106.500 109.930 106.965 110.320 ;
        RECT 106.275 109.120 106.625 109.740 ;
        RECT 106.795 109.340 106.965 109.930 ;
        RECT 107.135 109.710 107.305 110.490 ;
        RECT 107.475 110.390 107.645 110.730 ;
        RECT 107.880 110.560 108.210 110.990 ;
        RECT 108.380 110.390 108.550 110.730 ;
        RECT 108.845 110.530 109.215 110.990 ;
        RECT 107.475 110.220 108.550 110.390 ;
        RECT 109.385 110.360 109.555 110.820 ;
        RECT 109.790 110.480 110.660 110.820 ;
        RECT 110.830 110.530 111.080 110.990 ;
        RECT 108.995 110.190 109.555 110.360 ;
        RECT 108.995 110.050 109.165 110.190 ;
        RECT 107.665 109.880 109.165 110.050 ;
        RECT 109.860 110.020 110.320 110.310 ;
        RECT 107.135 109.540 108.825 109.710 ;
        RECT 106.795 109.120 107.150 109.340 ;
        RECT 107.320 108.830 107.490 109.540 ;
        RECT 107.695 109.120 108.485 109.370 ;
        RECT 108.655 109.360 108.825 109.540 ;
        RECT 108.995 109.190 109.165 109.880 ;
        RECT 105.435 108.440 105.765 108.800 ;
        RECT 105.935 108.660 106.430 108.830 ;
        RECT 106.635 108.660 107.490 108.830 ;
        RECT 108.365 108.440 108.695 108.900 ;
        RECT 108.905 108.800 109.165 109.190 ;
        RECT 109.355 110.010 110.320 110.020 ;
        RECT 110.490 110.100 110.660 110.480 ;
        RECT 111.250 110.440 111.420 110.730 ;
        RECT 111.600 110.610 111.930 110.990 ;
        RECT 111.250 110.270 112.050 110.440 ;
        RECT 109.355 109.850 110.030 110.010 ;
        RECT 110.490 109.930 111.710 110.100 ;
        RECT 109.355 109.060 109.565 109.850 ;
        RECT 110.490 109.840 110.660 109.930 ;
        RECT 109.735 109.060 110.085 109.680 ;
        RECT 110.255 109.670 110.660 109.840 ;
        RECT 110.255 108.890 110.425 109.670 ;
        RECT 110.595 109.220 110.815 109.500 ;
        RECT 110.995 109.390 111.535 109.760 ;
        RECT 111.880 109.650 112.050 110.270 ;
        RECT 112.225 109.930 112.395 110.990 ;
        RECT 112.605 109.980 112.895 110.820 ;
        RECT 113.065 110.150 113.235 110.990 ;
        RECT 113.445 109.980 113.695 110.820 ;
        RECT 113.905 110.150 114.075 110.990 ;
        RECT 112.605 109.810 114.330 109.980 ;
        RECT 110.595 109.050 111.125 109.220 ;
        RECT 108.905 108.630 109.255 108.800 ;
        RECT 109.475 108.610 110.425 108.890 ;
        RECT 110.595 108.440 110.785 108.880 ;
        RECT 110.955 108.820 111.125 109.050 ;
        RECT 111.295 108.990 111.535 109.390 ;
        RECT 111.705 109.640 112.050 109.650 ;
        RECT 111.705 109.430 113.735 109.640 ;
        RECT 111.705 109.175 112.030 109.430 ;
        RECT 113.920 109.260 114.330 109.810 ;
        RECT 114.555 109.900 115.765 110.990 ;
        RECT 114.555 109.360 115.075 109.900 ;
        RECT 111.705 108.820 112.025 109.175 ;
        RECT 110.955 108.650 112.025 108.820 ;
        RECT 112.225 108.440 112.395 109.250 ;
        RECT 112.565 109.090 114.330 109.260 ;
        RECT 115.245 109.190 115.765 109.730 ;
        RECT 112.565 108.610 112.895 109.090 ;
        RECT 113.065 108.440 113.235 108.910 ;
        RECT 113.405 108.610 113.735 109.090 ;
        RECT 113.905 108.440 114.075 108.910 ;
        RECT 114.555 108.440 115.765 109.190 ;
        RECT 10.510 108.270 115.850 108.440 ;
        RECT 10.595 107.520 11.805 108.270 ;
        RECT 10.595 106.980 11.115 107.520 ;
        RECT 12.035 107.450 12.245 108.270 ;
        RECT 12.415 107.470 12.745 108.100 ;
        RECT 11.285 106.810 11.805 107.350 ;
        RECT 12.415 106.870 12.665 107.470 ;
        RECT 12.915 107.450 13.145 108.270 ;
        RECT 13.395 107.450 13.625 108.270 ;
        RECT 13.795 107.470 14.125 108.100 ;
        RECT 12.835 107.030 13.165 107.280 ;
        RECT 13.375 107.030 13.705 107.280 ;
        RECT 13.875 106.870 14.125 107.470 ;
        RECT 14.295 107.450 14.505 108.270 ;
        RECT 15.045 107.800 15.215 108.270 ;
        RECT 15.385 107.620 15.715 108.100 ;
        RECT 15.885 107.800 16.055 108.270 ;
        RECT 16.225 107.620 16.555 108.100 ;
        RECT 14.790 107.450 16.555 107.620 ;
        RECT 16.725 107.460 16.895 108.270 ;
        RECT 17.095 107.890 18.165 108.060 ;
        RECT 17.095 107.535 17.415 107.890 ;
        RECT 10.595 105.720 11.805 106.810 ;
        RECT 12.035 105.720 12.245 106.860 ;
        RECT 12.415 105.890 12.745 106.870 ;
        RECT 12.915 105.720 13.145 106.860 ;
        RECT 13.395 105.720 13.625 106.860 ;
        RECT 13.795 105.890 14.125 106.870 ;
        RECT 14.790 106.900 15.200 107.450 ;
        RECT 17.090 107.280 17.415 107.535 ;
        RECT 15.385 107.070 17.415 107.280 ;
        RECT 17.070 107.060 17.415 107.070 ;
        RECT 17.585 107.320 17.825 107.720 ;
        RECT 17.995 107.660 18.165 107.890 ;
        RECT 18.335 107.830 18.525 108.270 ;
        RECT 18.695 107.820 19.645 108.100 ;
        RECT 19.865 107.910 20.215 108.080 ;
        RECT 17.995 107.490 18.525 107.660 ;
        RECT 14.295 105.720 14.505 106.860 ;
        RECT 14.790 106.730 16.515 106.900 ;
        RECT 15.045 105.720 15.215 106.560 ;
        RECT 15.425 105.890 15.675 106.730 ;
        RECT 15.885 105.720 16.055 106.560 ;
        RECT 16.225 105.890 16.515 106.730 ;
        RECT 16.725 105.720 16.895 106.780 ;
        RECT 17.070 106.440 17.240 107.060 ;
        RECT 17.585 106.950 18.125 107.320 ;
        RECT 18.305 107.210 18.525 107.490 ;
        RECT 18.695 107.040 18.865 107.820 ;
        RECT 18.460 106.870 18.865 107.040 ;
        RECT 19.035 107.030 19.385 107.650 ;
        RECT 18.460 106.780 18.630 106.870 ;
        RECT 19.555 106.860 19.765 107.650 ;
        RECT 17.410 106.610 18.630 106.780 ;
        RECT 19.090 106.700 19.765 106.860 ;
        RECT 17.070 106.270 17.870 106.440 ;
        RECT 17.190 105.720 17.520 106.100 ;
        RECT 17.700 105.980 17.870 106.270 ;
        RECT 18.460 106.230 18.630 106.610 ;
        RECT 18.800 106.690 19.765 106.700 ;
        RECT 19.955 107.520 20.215 107.910 ;
        RECT 20.425 107.810 20.755 108.270 ;
        RECT 21.630 107.880 22.485 108.050 ;
        RECT 22.690 107.880 23.185 108.050 ;
        RECT 23.355 107.910 23.685 108.270 ;
        RECT 19.955 106.830 20.125 107.520 ;
        RECT 20.295 107.170 20.465 107.350 ;
        RECT 20.635 107.340 21.425 107.590 ;
        RECT 21.630 107.170 21.800 107.880 ;
        RECT 21.970 107.370 22.325 107.590 ;
        RECT 20.295 107.000 21.985 107.170 ;
        RECT 18.800 106.400 19.260 106.690 ;
        RECT 19.955 106.660 21.455 106.830 ;
        RECT 19.955 106.520 20.125 106.660 ;
        RECT 19.565 106.350 20.125 106.520 ;
        RECT 18.040 105.720 18.290 106.180 ;
        RECT 18.460 105.890 19.330 106.230 ;
        RECT 19.565 105.890 19.735 106.350 ;
        RECT 20.570 106.320 21.645 106.490 ;
        RECT 19.905 105.720 20.275 106.180 ;
        RECT 20.570 105.980 20.740 106.320 ;
        RECT 20.910 105.720 21.240 106.150 ;
        RECT 21.475 105.980 21.645 106.320 ;
        RECT 21.815 106.220 21.985 107.000 ;
        RECT 22.155 106.780 22.325 107.370 ;
        RECT 22.495 106.970 22.845 107.590 ;
        RECT 22.155 106.390 22.620 106.780 ;
        RECT 23.015 106.520 23.185 107.880 ;
        RECT 23.355 106.690 23.815 107.740 ;
        RECT 22.790 106.350 23.185 106.520 ;
        RECT 22.790 106.220 22.960 106.350 ;
        RECT 21.815 105.890 22.495 106.220 ;
        RECT 22.710 105.890 22.960 106.220 ;
        RECT 23.130 105.720 23.380 106.180 ;
        RECT 23.550 105.905 23.875 106.690 ;
        RECT 24.045 105.890 24.215 108.010 ;
        RECT 24.385 107.890 24.715 108.270 ;
        RECT 24.885 107.720 25.140 108.010 ;
        RECT 24.390 107.550 25.140 107.720 ;
        RECT 24.390 106.560 24.620 107.550 ;
        RECT 25.315 107.545 25.605 108.270 ;
        RECT 25.835 107.450 26.045 108.270 ;
        RECT 26.215 107.470 26.545 108.100 ;
        RECT 24.790 106.730 25.140 107.380 ;
        RECT 24.390 106.390 25.140 106.560 ;
        RECT 24.385 105.720 24.715 106.220 ;
        RECT 24.885 105.890 25.140 106.390 ;
        RECT 25.315 105.720 25.605 106.885 ;
        RECT 26.215 106.870 26.465 107.470 ;
        RECT 26.715 107.450 26.945 108.270 ;
        RECT 27.195 107.450 27.425 108.270 ;
        RECT 27.595 107.470 27.925 108.100 ;
        RECT 26.635 107.030 26.965 107.280 ;
        RECT 27.175 107.030 27.505 107.280 ;
        RECT 27.675 106.870 27.925 107.470 ;
        RECT 28.095 107.450 28.305 108.270 ;
        RECT 28.575 107.450 28.805 108.270 ;
        RECT 28.975 107.470 29.305 108.100 ;
        RECT 28.555 107.030 28.885 107.280 ;
        RECT 29.055 106.870 29.305 107.470 ;
        RECT 29.475 107.450 29.685 108.270 ;
        RECT 29.920 107.720 30.175 108.010 ;
        RECT 30.345 107.890 30.675 108.270 ;
        RECT 29.920 107.550 30.670 107.720 ;
        RECT 25.835 105.720 26.045 106.860 ;
        RECT 26.215 105.890 26.545 106.870 ;
        RECT 26.715 105.720 26.945 106.860 ;
        RECT 27.195 105.720 27.425 106.860 ;
        RECT 27.595 105.890 27.925 106.870 ;
        RECT 28.095 105.720 28.305 106.860 ;
        RECT 28.575 105.720 28.805 106.860 ;
        RECT 28.975 105.890 29.305 106.870 ;
        RECT 29.475 105.720 29.685 106.860 ;
        RECT 29.920 106.730 30.270 107.380 ;
        RECT 30.440 106.560 30.670 107.550 ;
        RECT 29.920 106.390 30.670 106.560 ;
        RECT 29.920 105.890 30.175 106.390 ;
        RECT 30.345 105.720 30.675 106.220 ;
        RECT 30.845 105.890 31.015 108.010 ;
        RECT 31.375 107.910 31.705 108.270 ;
        RECT 31.875 107.880 32.370 108.050 ;
        RECT 32.575 107.880 33.430 108.050 ;
        RECT 31.245 106.690 31.705 107.740 ;
        RECT 31.185 105.905 31.510 106.690 ;
        RECT 31.875 106.520 32.045 107.880 ;
        RECT 32.215 106.970 32.565 107.590 ;
        RECT 32.735 107.370 33.090 107.590 ;
        RECT 32.735 106.780 32.905 107.370 ;
        RECT 33.260 107.170 33.430 107.880 ;
        RECT 34.305 107.810 34.635 108.270 ;
        RECT 34.845 107.910 35.195 108.080 ;
        RECT 33.635 107.340 34.425 107.590 ;
        RECT 34.845 107.520 35.105 107.910 ;
        RECT 35.415 107.820 36.365 108.100 ;
        RECT 36.535 107.830 36.725 108.270 ;
        RECT 36.895 107.890 37.965 108.060 ;
        RECT 34.595 107.170 34.765 107.350 ;
        RECT 31.875 106.350 32.270 106.520 ;
        RECT 32.440 106.390 32.905 106.780 ;
        RECT 33.075 107.000 34.765 107.170 ;
        RECT 32.100 106.220 32.270 106.350 ;
        RECT 33.075 106.220 33.245 107.000 ;
        RECT 34.935 106.830 35.105 107.520 ;
        RECT 33.605 106.660 35.105 106.830 ;
        RECT 35.295 106.860 35.505 107.650 ;
        RECT 35.675 107.030 36.025 107.650 ;
        RECT 36.195 107.040 36.365 107.820 ;
        RECT 36.895 107.660 37.065 107.890 ;
        RECT 36.535 107.490 37.065 107.660 ;
        RECT 36.535 107.210 36.755 107.490 ;
        RECT 37.235 107.320 37.475 107.720 ;
        RECT 36.195 106.870 36.600 107.040 ;
        RECT 36.935 106.950 37.475 107.320 ;
        RECT 37.645 107.535 37.965 107.890 ;
        RECT 37.645 107.280 37.970 107.535 ;
        RECT 38.165 107.460 38.335 108.270 ;
        RECT 38.505 107.620 38.835 108.100 ;
        RECT 39.005 107.800 39.175 108.270 ;
        RECT 39.345 107.620 39.675 108.100 ;
        RECT 39.845 107.800 40.015 108.270 ;
        RECT 40.805 107.800 40.975 108.270 ;
        RECT 41.145 107.620 41.475 108.100 ;
        RECT 41.645 107.800 41.815 108.270 ;
        RECT 41.985 107.620 42.315 108.100 ;
        RECT 38.505 107.450 40.270 107.620 ;
        RECT 37.645 107.070 39.675 107.280 ;
        RECT 37.645 107.060 37.990 107.070 ;
        RECT 35.295 106.700 35.970 106.860 ;
        RECT 36.430 106.780 36.600 106.870 ;
        RECT 35.295 106.690 36.260 106.700 ;
        RECT 34.935 106.520 35.105 106.660 ;
        RECT 31.680 105.720 31.930 106.180 ;
        RECT 32.100 105.890 32.350 106.220 ;
        RECT 32.565 105.890 33.245 106.220 ;
        RECT 33.415 106.320 34.490 106.490 ;
        RECT 34.935 106.350 35.495 106.520 ;
        RECT 35.800 106.400 36.260 106.690 ;
        RECT 36.430 106.610 37.650 106.780 ;
        RECT 33.415 105.980 33.585 106.320 ;
        RECT 33.820 105.720 34.150 106.150 ;
        RECT 34.320 105.980 34.490 106.320 ;
        RECT 34.785 105.720 35.155 106.180 ;
        RECT 35.325 105.890 35.495 106.350 ;
        RECT 36.430 106.230 36.600 106.610 ;
        RECT 37.820 106.440 37.990 107.060 ;
        RECT 39.860 106.900 40.270 107.450 ;
        RECT 35.730 105.890 36.600 106.230 ;
        RECT 37.190 106.270 37.990 106.440 ;
        RECT 36.770 105.720 37.020 106.180 ;
        RECT 37.190 105.980 37.360 106.270 ;
        RECT 37.540 105.720 37.870 106.100 ;
        RECT 38.165 105.720 38.335 106.780 ;
        RECT 38.545 106.730 40.270 106.900 ;
        RECT 40.550 107.450 42.315 107.620 ;
        RECT 42.485 107.460 42.655 108.270 ;
        RECT 42.855 107.890 43.925 108.060 ;
        RECT 42.855 107.535 43.175 107.890 ;
        RECT 40.550 106.900 40.960 107.450 ;
        RECT 42.850 107.280 43.175 107.535 ;
        RECT 41.145 107.070 43.175 107.280 ;
        RECT 42.830 107.060 43.175 107.070 ;
        RECT 43.345 107.320 43.585 107.720 ;
        RECT 43.755 107.660 43.925 107.890 ;
        RECT 44.095 107.830 44.285 108.270 ;
        RECT 44.455 107.820 45.405 108.100 ;
        RECT 45.625 107.910 45.975 108.080 ;
        RECT 43.755 107.490 44.285 107.660 ;
        RECT 40.550 106.730 42.275 106.900 ;
        RECT 38.545 105.890 38.835 106.730 ;
        RECT 39.005 105.720 39.175 106.560 ;
        RECT 39.385 105.890 39.635 106.730 ;
        RECT 39.845 105.720 40.015 106.560 ;
        RECT 40.805 105.720 40.975 106.560 ;
        RECT 41.185 105.890 41.435 106.730 ;
        RECT 41.645 105.720 41.815 106.560 ;
        RECT 41.985 105.890 42.275 106.730 ;
        RECT 42.485 105.720 42.655 106.780 ;
        RECT 42.830 106.440 43.000 107.060 ;
        RECT 43.345 106.950 43.885 107.320 ;
        RECT 44.065 107.210 44.285 107.490 ;
        RECT 44.455 107.040 44.625 107.820 ;
        RECT 44.220 106.870 44.625 107.040 ;
        RECT 44.795 107.030 45.145 107.650 ;
        RECT 44.220 106.780 44.390 106.870 ;
        RECT 45.315 106.860 45.525 107.650 ;
        RECT 43.170 106.610 44.390 106.780 ;
        RECT 44.850 106.700 45.525 106.860 ;
        RECT 42.830 106.270 43.630 106.440 ;
        RECT 42.950 105.720 43.280 106.100 ;
        RECT 43.460 105.980 43.630 106.270 ;
        RECT 44.220 106.230 44.390 106.610 ;
        RECT 44.560 106.690 45.525 106.700 ;
        RECT 45.715 107.520 45.975 107.910 ;
        RECT 46.185 107.810 46.515 108.270 ;
        RECT 47.390 107.880 48.245 108.050 ;
        RECT 48.450 107.880 48.945 108.050 ;
        RECT 49.115 107.910 49.445 108.270 ;
        RECT 45.715 106.830 45.885 107.520 ;
        RECT 46.055 107.170 46.225 107.350 ;
        RECT 46.395 107.340 47.185 107.590 ;
        RECT 47.390 107.170 47.560 107.880 ;
        RECT 47.730 107.370 48.085 107.590 ;
        RECT 46.055 107.000 47.745 107.170 ;
        RECT 44.560 106.400 45.020 106.690 ;
        RECT 45.715 106.660 47.215 106.830 ;
        RECT 45.715 106.520 45.885 106.660 ;
        RECT 45.325 106.350 45.885 106.520 ;
        RECT 43.800 105.720 44.050 106.180 ;
        RECT 44.220 105.890 45.090 106.230 ;
        RECT 45.325 105.890 45.495 106.350 ;
        RECT 46.330 106.320 47.405 106.490 ;
        RECT 45.665 105.720 46.035 106.180 ;
        RECT 46.330 105.980 46.500 106.320 ;
        RECT 46.670 105.720 47.000 106.150 ;
        RECT 47.235 105.980 47.405 106.320 ;
        RECT 47.575 106.220 47.745 107.000 ;
        RECT 47.915 106.780 48.085 107.370 ;
        RECT 48.255 106.970 48.605 107.590 ;
        RECT 47.915 106.390 48.380 106.780 ;
        RECT 48.775 106.520 48.945 107.880 ;
        RECT 49.115 106.690 49.575 107.740 ;
        RECT 48.550 106.350 48.945 106.520 ;
        RECT 48.550 106.220 48.720 106.350 ;
        RECT 47.575 105.890 48.255 106.220 ;
        RECT 48.470 105.890 48.720 106.220 ;
        RECT 48.890 105.720 49.140 106.180 ;
        RECT 49.310 105.905 49.635 106.690 ;
        RECT 49.805 105.890 49.975 108.010 ;
        RECT 50.145 107.890 50.475 108.270 ;
        RECT 50.645 107.720 50.900 108.010 ;
        RECT 50.150 107.550 50.900 107.720 ;
        RECT 50.150 106.560 50.380 107.550 ;
        RECT 51.075 107.545 51.365 108.270 ;
        RECT 52.305 107.800 52.475 108.270 ;
        RECT 52.645 107.620 52.975 108.100 ;
        RECT 53.145 107.800 53.315 108.270 ;
        RECT 53.485 107.620 53.815 108.100 ;
        RECT 52.050 107.450 53.815 107.620 ;
        RECT 53.985 107.460 54.155 108.270 ;
        RECT 54.355 107.890 55.425 108.060 ;
        RECT 54.355 107.535 54.675 107.890 ;
        RECT 50.550 106.730 50.900 107.380 ;
        RECT 52.050 106.900 52.460 107.450 ;
        RECT 54.350 107.280 54.675 107.535 ;
        RECT 52.645 107.070 54.675 107.280 ;
        RECT 54.330 107.060 54.675 107.070 ;
        RECT 54.845 107.320 55.085 107.720 ;
        RECT 55.255 107.660 55.425 107.890 ;
        RECT 55.595 107.830 55.785 108.270 ;
        RECT 55.955 107.820 56.905 108.100 ;
        RECT 57.125 107.910 57.475 108.080 ;
        RECT 55.255 107.490 55.785 107.660 ;
        RECT 50.150 106.390 50.900 106.560 ;
        RECT 50.145 105.720 50.475 106.220 ;
        RECT 50.645 105.890 50.900 106.390 ;
        RECT 51.075 105.720 51.365 106.885 ;
        RECT 52.050 106.730 53.775 106.900 ;
        RECT 52.305 105.720 52.475 106.560 ;
        RECT 52.685 105.890 52.935 106.730 ;
        RECT 53.145 105.720 53.315 106.560 ;
        RECT 53.485 105.890 53.775 106.730 ;
        RECT 53.985 105.720 54.155 106.780 ;
        RECT 54.330 106.440 54.500 107.060 ;
        RECT 54.845 106.950 55.385 107.320 ;
        RECT 55.565 107.210 55.785 107.490 ;
        RECT 55.955 107.040 56.125 107.820 ;
        RECT 55.720 106.870 56.125 107.040 ;
        RECT 56.295 107.030 56.645 107.650 ;
        RECT 55.720 106.780 55.890 106.870 ;
        RECT 56.815 106.860 57.025 107.650 ;
        RECT 54.670 106.610 55.890 106.780 ;
        RECT 56.350 106.700 57.025 106.860 ;
        RECT 54.330 106.270 55.130 106.440 ;
        RECT 54.450 105.720 54.780 106.100 ;
        RECT 54.960 105.980 55.130 106.270 ;
        RECT 55.720 106.230 55.890 106.610 ;
        RECT 56.060 106.690 57.025 106.700 ;
        RECT 57.215 107.520 57.475 107.910 ;
        RECT 57.685 107.810 58.015 108.270 ;
        RECT 58.890 107.880 59.745 108.050 ;
        RECT 59.950 107.880 60.445 108.050 ;
        RECT 60.615 107.910 60.945 108.270 ;
        RECT 57.215 106.830 57.385 107.520 ;
        RECT 57.555 107.170 57.725 107.350 ;
        RECT 57.895 107.340 58.685 107.590 ;
        RECT 58.890 107.170 59.060 107.880 ;
        RECT 59.230 107.370 59.585 107.590 ;
        RECT 57.555 107.000 59.245 107.170 ;
        RECT 56.060 106.400 56.520 106.690 ;
        RECT 57.215 106.660 58.715 106.830 ;
        RECT 57.215 106.520 57.385 106.660 ;
        RECT 56.825 106.350 57.385 106.520 ;
        RECT 55.300 105.720 55.550 106.180 ;
        RECT 55.720 105.890 56.590 106.230 ;
        RECT 56.825 105.890 56.995 106.350 ;
        RECT 57.830 106.320 58.905 106.490 ;
        RECT 57.165 105.720 57.535 106.180 ;
        RECT 57.830 105.980 58.000 106.320 ;
        RECT 58.170 105.720 58.500 106.150 ;
        RECT 58.735 105.980 58.905 106.320 ;
        RECT 59.075 106.220 59.245 107.000 ;
        RECT 59.415 106.780 59.585 107.370 ;
        RECT 59.755 106.970 60.105 107.590 ;
        RECT 59.415 106.390 59.880 106.780 ;
        RECT 60.275 106.520 60.445 107.880 ;
        RECT 60.615 106.690 61.075 107.740 ;
        RECT 60.050 106.350 60.445 106.520 ;
        RECT 60.050 106.220 60.220 106.350 ;
        RECT 59.075 105.890 59.755 106.220 ;
        RECT 59.970 105.890 60.220 106.220 ;
        RECT 60.390 105.720 60.640 106.180 ;
        RECT 60.810 105.905 61.135 106.690 ;
        RECT 61.305 105.890 61.475 108.010 ;
        RECT 61.645 107.890 61.975 108.270 ;
        RECT 62.145 107.720 62.400 108.010 ;
        RECT 63.805 107.800 63.975 108.270 ;
        RECT 61.650 107.550 62.400 107.720 ;
        RECT 64.145 107.620 64.475 108.100 ;
        RECT 64.645 107.800 64.815 108.270 ;
        RECT 64.985 107.620 65.315 108.100 ;
        RECT 61.650 106.560 61.880 107.550 ;
        RECT 63.550 107.450 65.315 107.620 ;
        RECT 65.485 107.460 65.655 108.270 ;
        RECT 65.855 107.890 66.925 108.060 ;
        RECT 65.855 107.535 66.175 107.890 ;
        RECT 62.050 106.730 62.400 107.380 ;
        RECT 63.550 106.900 63.960 107.450 ;
        RECT 65.850 107.280 66.175 107.535 ;
        RECT 64.145 107.070 66.175 107.280 ;
        RECT 65.830 107.060 66.175 107.070 ;
        RECT 66.345 107.320 66.585 107.720 ;
        RECT 66.755 107.660 66.925 107.890 ;
        RECT 67.095 107.830 67.285 108.270 ;
        RECT 67.455 107.820 68.405 108.100 ;
        RECT 68.625 107.910 68.975 108.080 ;
        RECT 66.755 107.490 67.285 107.660 ;
        RECT 63.550 106.730 65.275 106.900 ;
        RECT 61.650 106.390 62.400 106.560 ;
        RECT 61.645 105.720 61.975 106.220 ;
        RECT 62.145 105.890 62.400 106.390 ;
        RECT 63.805 105.720 63.975 106.560 ;
        RECT 64.185 105.890 64.435 106.730 ;
        RECT 64.645 105.720 64.815 106.560 ;
        RECT 64.985 105.890 65.275 106.730 ;
        RECT 65.485 105.720 65.655 106.780 ;
        RECT 65.830 106.440 66.000 107.060 ;
        RECT 66.345 106.950 66.885 107.320 ;
        RECT 67.065 107.210 67.285 107.490 ;
        RECT 67.455 107.040 67.625 107.820 ;
        RECT 67.220 106.870 67.625 107.040 ;
        RECT 67.795 107.030 68.145 107.650 ;
        RECT 67.220 106.780 67.390 106.870 ;
        RECT 68.315 106.860 68.525 107.650 ;
        RECT 66.170 106.610 67.390 106.780 ;
        RECT 67.850 106.700 68.525 106.860 ;
        RECT 65.830 106.270 66.630 106.440 ;
        RECT 65.950 105.720 66.280 106.100 ;
        RECT 66.460 105.980 66.630 106.270 ;
        RECT 67.220 106.230 67.390 106.610 ;
        RECT 67.560 106.690 68.525 106.700 ;
        RECT 68.715 107.520 68.975 107.910 ;
        RECT 69.185 107.810 69.515 108.270 ;
        RECT 70.390 107.880 71.245 108.050 ;
        RECT 71.450 107.880 71.945 108.050 ;
        RECT 72.115 107.910 72.445 108.270 ;
        RECT 68.715 106.830 68.885 107.520 ;
        RECT 69.055 107.170 69.225 107.350 ;
        RECT 69.395 107.340 70.185 107.590 ;
        RECT 70.390 107.170 70.560 107.880 ;
        RECT 70.730 107.370 71.085 107.590 ;
        RECT 69.055 107.000 70.745 107.170 ;
        RECT 67.560 106.400 68.020 106.690 ;
        RECT 68.715 106.660 70.215 106.830 ;
        RECT 68.715 106.520 68.885 106.660 ;
        RECT 68.325 106.350 68.885 106.520 ;
        RECT 66.800 105.720 67.050 106.180 ;
        RECT 67.220 105.890 68.090 106.230 ;
        RECT 68.325 105.890 68.495 106.350 ;
        RECT 69.330 106.320 70.405 106.490 ;
        RECT 68.665 105.720 69.035 106.180 ;
        RECT 69.330 105.980 69.500 106.320 ;
        RECT 69.670 105.720 70.000 106.150 ;
        RECT 70.235 105.980 70.405 106.320 ;
        RECT 70.575 106.220 70.745 107.000 ;
        RECT 70.915 106.780 71.085 107.370 ;
        RECT 71.255 106.970 71.605 107.590 ;
        RECT 70.915 106.390 71.380 106.780 ;
        RECT 71.775 106.520 71.945 107.880 ;
        RECT 72.115 106.690 72.575 107.740 ;
        RECT 71.550 106.350 71.945 106.520 ;
        RECT 71.550 106.220 71.720 106.350 ;
        RECT 70.575 105.890 71.255 106.220 ;
        RECT 71.470 105.890 71.720 106.220 ;
        RECT 71.890 105.720 72.140 106.180 ;
        RECT 72.310 105.905 72.635 106.690 ;
        RECT 72.805 105.890 72.975 108.010 ;
        RECT 73.145 107.890 73.475 108.270 ;
        RECT 73.645 107.720 73.900 108.010 ;
        RECT 73.150 107.550 73.900 107.720 ;
        RECT 73.150 106.560 73.380 107.550 ;
        RECT 74.135 107.450 74.345 108.270 ;
        RECT 74.515 107.470 74.845 108.100 ;
        RECT 73.550 106.730 73.900 107.380 ;
        RECT 74.515 106.870 74.765 107.470 ;
        RECT 75.015 107.450 75.245 108.270 ;
        RECT 75.495 107.450 75.725 108.270 ;
        RECT 75.895 107.470 76.225 108.100 ;
        RECT 74.935 107.030 75.265 107.280 ;
        RECT 75.475 107.030 75.805 107.280 ;
        RECT 75.975 106.870 76.225 107.470 ;
        RECT 76.395 107.450 76.605 108.270 ;
        RECT 76.835 107.545 77.125 108.270 ;
        RECT 77.605 107.800 77.775 108.270 ;
        RECT 77.945 107.620 78.275 108.100 ;
        RECT 78.445 107.800 78.615 108.270 ;
        RECT 78.785 107.620 79.115 108.100 ;
        RECT 77.350 107.450 79.115 107.620 ;
        RECT 79.285 107.460 79.455 108.270 ;
        RECT 79.655 107.890 80.725 108.060 ;
        RECT 79.655 107.535 79.975 107.890 ;
        RECT 77.350 106.900 77.760 107.450 ;
        RECT 79.650 107.280 79.975 107.535 ;
        RECT 77.945 107.070 79.975 107.280 ;
        RECT 79.630 107.060 79.975 107.070 ;
        RECT 80.145 107.320 80.385 107.720 ;
        RECT 80.555 107.660 80.725 107.890 ;
        RECT 80.895 107.830 81.085 108.270 ;
        RECT 81.255 107.820 82.205 108.100 ;
        RECT 82.425 107.910 82.775 108.080 ;
        RECT 80.555 107.490 81.085 107.660 ;
        RECT 73.150 106.390 73.900 106.560 ;
        RECT 73.145 105.720 73.475 106.220 ;
        RECT 73.645 105.890 73.900 106.390 ;
        RECT 74.135 105.720 74.345 106.860 ;
        RECT 74.515 105.890 74.845 106.870 ;
        RECT 75.015 105.720 75.245 106.860 ;
        RECT 75.495 105.720 75.725 106.860 ;
        RECT 75.895 105.890 76.225 106.870 ;
        RECT 76.395 105.720 76.605 106.860 ;
        RECT 76.835 105.720 77.125 106.885 ;
        RECT 77.350 106.730 79.075 106.900 ;
        RECT 77.605 105.720 77.775 106.560 ;
        RECT 77.985 105.890 78.235 106.730 ;
        RECT 78.445 105.720 78.615 106.560 ;
        RECT 78.785 105.890 79.075 106.730 ;
        RECT 79.285 105.720 79.455 106.780 ;
        RECT 79.630 106.440 79.800 107.060 ;
        RECT 80.145 106.950 80.685 107.320 ;
        RECT 80.865 107.210 81.085 107.490 ;
        RECT 81.255 107.040 81.425 107.820 ;
        RECT 81.020 106.870 81.425 107.040 ;
        RECT 81.595 107.030 81.945 107.650 ;
        RECT 81.020 106.780 81.190 106.870 ;
        RECT 82.115 106.860 82.325 107.650 ;
        RECT 79.970 106.610 81.190 106.780 ;
        RECT 81.650 106.700 82.325 106.860 ;
        RECT 79.630 106.270 80.430 106.440 ;
        RECT 79.750 105.720 80.080 106.100 ;
        RECT 80.260 105.980 80.430 106.270 ;
        RECT 81.020 106.230 81.190 106.610 ;
        RECT 81.360 106.690 82.325 106.700 ;
        RECT 82.515 107.520 82.775 107.910 ;
        RECT 82.985 107.810 83.315 108.270 ;
        RECT 84.190 107.880 85.045 108.050 ;
        RECT 85.250 107.880 85.745 108.050 ;
        RECT 85.915 107.910 86.245 108.270 ;
        RECT 82.515 106.830 82.685 107.520 ;
        RECT 82.855 107.170 83.025 107.350 ;
        RECT 83.195 107.340 83.985 107.590 ;
        RECT 84.190 107.170 84.360 107.880 ;
        RECT 84.530 107.370 84.885 107.590 ;
        RECT 82.855 107.000 84.545 107.170 ;
        RECT 81.360 106.400 81.820 106.690 ;
        RECT 82.515 106.660 84.015 106.830 ;
        RECT 82.515 106.520 82.685 106.660 ;
        RECT 82.125 106.350 82.685 106.520 ;
        RECT 80.600 105.720 80.850 106.180 ;
        RECT 81.020 105.890 81.890 106.230 ;
        RECT 82.125 105.890 82.295 106.350 ;
        RECT 83.130 106.320 84.205 106.490 ;
        RECT 82.465 105.720 82.835 106.180 ;
        RECT 83.130 105.980 83.300 106.320 ;
        RECT 83.470 105.720 83.800 106.150 ;
        RECT 84.035 105.980 84.205 106.320 ;
        RECT 84.375 106.220 84.545 107.000 ;
        RECT 84.715 106.780 84.885 107.370 ;
        RECT 85.055 106.970 85.405 107.590 ;
        RECT 84.715 106.390 85.180 106.780 ;
        RECT 85.575 106.520 85.745 107.880 ;
        RECT 85.915 106.690 86.375 107.740 ;
        RECT 85.350 106.350 85.745 106.520 ;
        RECT 85.350 106.220 85.520 106.350 ;
        RECT 84.375 105.890 85.055 106.220 ;
        RECT 85.270 105.890 85.520 106.220 ;
        RECT 85.690 105.720 85.940 106.180 ;
        RECT 86.110 105.905 86.435 106.690 ;
        RECT 86.605 105.890 86.775 108.010 ;
        RECT 86.945 107.890 87.275 108.270 ;
        RECT 87.445 107.720 87.700 108.010 ;
        RECT 88.185 107.800 88.355 108.270 ;
        RECT 86.950 107.550 87.700 107.720 ;
        RECT 88.525 107.620 88.855 108.100 ;
        RECT 89.025 107.800 89.195 108.270 ;
        RECT 89.365 107.620 89.695 108.100 ;
        RECT 86.950 106.560 87.180 107.550 ;
        RECT 87.930 107.450 89.695 107.620 ;
        RECT 89.865 107.460 90.035 108.270 ;
        RECT 90.235 107.890 91.305 108.060 ;
        RECT 90.235 107.535 90.555 107.890 ;
        RECT 87.350 106.730 87.700 107.380 ;
        RECT 87.930 106.900 88.340 107.450 ;
        RECT 90.230 107.280 90.555 107.535 ;
        RECT 88.525 107.070 90.555 107.280 ;
        RECT 90.210 107.060 90.555 107.070 ;
        RECT 90.725 107.320 90.965 107.720 ;
        RECT 91.135 107.660 91.305 107.890 ;
        RECT 91.475 107.830 91.665 108.270 ;
        RECT 91.835 107.820 92.785 108.100 ;
        RECT 93.005 107.910 93.355 108.080 ;
        RECT 91.135 107.490 91.665 107.660 ;
        RECT 87.930 106.730 89.655 106.900 ;
        RECT 86.950 106.390 87.700 106.560 ;
        RECT 86.945 105.720 87.275 106.220 ;
        RECT 87.445 105.890 87.700 106.390 ;
        RECT 88.185 105.720 88.355 106.560 ;
        RECT 88.565 105.890 88.815 106.730 ;
        RECT 89.025 105.720 89.195 106.560 ;
        RECT 89.365 105.890 89.655 106.730 ;
        RECT 89.865 105.720 90.035 106.780 ;
        RECT 90.210 106.440 90.380 107.060 ;
        RECT 90.725 106.950 91.265 107.320 ;
        RECT 91.445 107.210 91.665 107.490 ;
        RECT 91.835 107.040 92.005 107.820 ;
        RECT 91.600 106.870 92.005 107.040 ;
        RECT 92.175 107.030 92.525 107.650 ;
        RECT 91.600 106.780 91.770 106.870 ;
        RECT 92.695 106.860 92.905 107.650 ;
        RECT 90.550 106.610 91.770 106.780 ;
        RECT 92.230 106.700 92.905 106.860 ;
        RECT 90.210 106.270 91.010 106.440 ;
        RECT 90.330 105.720 90.660 106.100 ;
        RECT 90.840 105.980 91.010 106.270 ;
        RECT 91.600 106.230 91.770 106.610 ;
        RECT 91.940 106.690 92.905 106.700 ;
        RECT 93.095 107.520 93.355 107.910 ;
        RECT 93.565 107.810 93.895 108.270 ;
        RECT 94.770 107.880 95.625 108.050 ;
        RECT 95.830 107.880 96.325 108.050 ;
        RECT 96.495 107.910 96.825 108.270 ;
        RECT 93.095 106.830 93.265 107.520 ;
        RECT 93.435 107.170 93.605 107.350 ;
        RECT 93.775 107.340 94.565 107.590 ;
        RECT 94.770 107.170 94.940 107.880 ;
        RECT 95.110 107.370 95.465 107.590 ;
        RECT 93.435 107.000 95.125 107.170 ;
        RECT 91.940 106.400 92.400 106.690 ;
        RECT 93.095 106.660 94.595 106.830 ;
        RECT 93.095 106.520 93.265 106.660 ;
        RECT 92.705 106.350 93.265 106.520 ;
        RECT 91.180 105.720 91.430 106.180 ;
        RECT 91.600 105.890 92.470 106.230 ;
        RECT 92.705 105.890 92.875 106.350 ;
        RECT 93.710 106.320 94.785 106.490 ;
        RECT 93.045 105.720 93.415 106.180 ;
        RECT 93.710 105.980 93.880 106.320 ;
        RECT 94.050 105.720 94.380 106.150 ;
        RECT 94.615 105.980 94.785 106.320 ;
        RECT 94.955 106.220 95.125 107.000 ;
        RECT 95.295 106.780 95.465 107.370 ;
        RECT 95.635 106.970 95.985 107.590 ;
        RECT 95.295 106.390 95.760 106.780 ;
        RECT 96.155 106.520 96.325 107.880 ;
        RECT 96.495 106.690 96.955 107.740 ;
        RECT 95.930 106.350 96.325 106.520 ;
        RECT 95.930 106.220 96.100 106.350 ;
        RECT 94.955 105.890 95.635 106.220 ;
        RECT 95.850 105.890 96.100 106.220 ;
        RECT 96.270 105.720 96.520 106.180 ;
        RECT 96.690 105.905 97.015 106.690 ;
        RECT 97.185 105.890 97.355 108.010 ;
        RECT 97.525 107.890 97.855 108.270 ;
        RECT 98.025 107.720 98.280 108.010 ;
        RECT 97.530 107.550 98.280 107.720 ;
        RECT 97.530 106.560 97.760 107.550 ;
        RECT 98.515 107.450 98.725 108.270 ;
        RECT 98.895 107.470 99.225 108.100 ;
        RECT 97.930 106.730 98.280 107.380 ;
        RECT 98.895 106.870 99.145 107.470 ;
        RECT 99.395 107.450 99.625 108.270 ;
        RECT 99.895 107.450 100.105 108.270 ;
        RECT 100.275 107.470 100.605 108.100 ;
        RECT 99.315 107.030 99.645 107.280 ;
        RECT 100.275 106.870 100.525 107.470 ;
        RECT 100.775 107.450 101.005 108.270 ;
        RECT 101.255 107.450 101.485 108.270 ;
        RECT 101.655 107.470 101.985 108.100 ;
        RECT 100.695 107.030 101.025 107.280 ;
        RECT 101.235 107.030 101.565 107.280 ;
        RECT 101.735 106.870 101.985 107.470 ;
        RECT 102.155 107.450 102.365 108.270 ;
        RECT 102.595 107.545 102.885 108.270 ;
        RECT 103.365 107.800 103.535 108.270 ;
        RECT 103.705 107.620 104.035 108.100 ;
        RECT 104.205 107.800 104.375 108.270 ;
        RECT 104.545 107.620 104.875 108.100 ;
        RECT 103.110 107.450 104.875 107.620 ;
        RECT 105.045 107.460 105.215 108.270 ;
        RECT 105.415 107.890 106.485 108.060 ;
        RECT 105.415 107.535 105.735 107.890 ;
        RECT 103.110 106.900 103.520 107.450 ;
        RECT 105.410 107.280 105.735 107.535 ;
        RECT 103.705 107.070 105.735 107.280 ;
        RECT 105.390 107.060 105.735 107.070 ;
        RECT 105.905 107.320 106.145 107.720 ;
        RECT 106.315 107.660 106.485 107.890 ;
        RECT 106.655 107.830 106.845 108.270 ;
        RECT 107.015 107.820 107.965 108.100 ;
        RECT 108.185 107.910 108.535 108.080 ;
        RECT 106.315 107.490 106.845 107.660 ;
        RECT 97.530 106.390 98.280 106.560 ;
        RECT 97.525 105.720 97.855 106.220 ;
        RECT 98.025 105.890 98.280 106.390 ;
        RECT 98.515 105.720 98.725 106.860 ;
        RECT 98.895 105.890 99.225 106.870 ;
        RECT 99.395 105.720 99.625 106.860 ;
        RECT 99.895 105.720 100.105 106.860 ;
        RECT 100.275 105.890 100.605 106.870 ;
        RECT 100.775 105.720 101.005 106.860 ;
        RECT 101.255 105.720 101.485 106.860 ;
        RECT 101.655 105.890 101.985 106.870 ;
        RECT 102.155 105.720 102.365 106.860 ;
        RECT 102.595 105.720 102.885 106.885 ;
        RECT 103.110 106.730 104.835 106.900 ;
        RECT 103.365 105.720 103.535 106.560 ;
        RECT 103.745 105.890 103.995 106.730 ;
        RECT 104.205 105.720 104.375 106.560 ;
        RECT 104.545 105.890 104.835 106.730 ;
        RECT 105.045 105.720 105.215 106.780 ;
        RECT 105.390 106.440 105.560 107.060 ;
        RECT 105.905 106.950 106.445 107.320 ;
        RECT 106.625 107.210 106.845 107.490 ;
        RECT 107.015 107.040 107.185 107.820 ;
        RECT 106.780 106.870 107.185 107.040 ;
        RECT 107.355 107.030 107.705 107.650 ;
        RECT 106.780 106.780 106.950 106.870 ;
        RECT 107.875 106.860 108.085 107.650 ;
        RECT 105.730 106.610 106.950 106.780 ;
        RECT 107.410 106.700 108.085 106.860 ;
        RECT 105.390 106.270 106.190 106.440 ;
        RECT 105.510 105.720 105.840 106.100 ;
        RECT 106.020 105.980 106.190 106.270 ;
        RECT 106.780 106.230 106.950 106.610 ;
        RECT 107.120 106.690 108.085 106.700 ;
        RECT 108.275 107.520 108.535 107.910 ;
        RECT 108.745 107.810 109.075 108.270 ;
        RECT 109.950 107.880 110.805 108.050 ;
        RECT 111.010 107.880 111.505 108.050 ;
        RECT 111.675 107.910 112.005 108.270 ;
        RECT 108.275 106.830 108.445 107.520 ;
        RECT 108.615 107.170 108.785 107.350 ;
        RECT 108.955 107.340 109.745 107.590 ;
        RECT 109.950 107.170 110.120 107.880 ;
        RECT 110.290 107.370 110.645 107.590 ;
        RECT 108.615 107.000 110.305 107.170 ;
        RECT 107.120 106.400 107.580 106.690 ;
        RECT 108.275 106.660 109.775 106.830 ;
        RECT 108.275 106.520 108.445 106.660 ;
        RECT 107.885 106.350 108.445 106.520 ;
        RECT 106.360 105.720 106.610 106.180 ;
        RECT 106.780 105.890 107.650 106.230 ;
        RECT 107.885 105.890 108.055 106.350 ;
        RECT 108.890 106.320 109.965 106.490 ;
        RECT 108.225 105.720 108.595 106.180 ;
        RECT 108.890 105.980 109.060 106.320 ;
        RECT 109.230 105.720 109.560 106.150 ;
        RECT 109.795 105.980 109.965 106.320 ;
        RECT 110.135 106.220 110.305 107.000 ;
        RECT 110.475 106.780 110.645 107.370 ;
        RECT 110.815 106.970 111.165 107.590 ;
        RECT 110.475 106.390 110.940 106.780 ;
        RECT 111.335 106.520 111.505 107.880 ;
        RECT 111.675 106.690 112.135 107.740 ;
        RECT 111.110 106.350 111.505 106.520 ;
        RECT 111.110 106.220 111.280 106.350 ;
        RECT 110.135 105.890 110.815 106.220 ;
        RECT 111.030 105.890 111.280 106.220 ;
        RECT 111.450 105.720 111.700 106.180 ;
        RECT 111.870 105.905 112.195 106.690 ;
        RECT 112.365 105.890 112.535 108.010 ;
        RECT 112.705 107.890 113.035 108.270 ;
        RECT 113.205 107.720 113.460 108.010 ;
        RECT 112.710 107.550 113.460 107.720 ;
        RECT 112.710 106.560 112.940 107.550 ;
        RECT 114.555 107.520 115.765 108.270 ;
        RECT 113.110 106.730 113.460 107.380 ;
        RECT 114.555 106.810 115.075 107.350 ;
        RECT 115.245 106.980 115.765 107.520 ;
        RECT 112.710 106.390 113.460 106.560 ;
        RECT 112.705 105.720 113.035 106.220 ;
        RECT 113.205 105.890 113.460 106.390 ;
        RECT 114.555 105.720 115.765 106.810 ;
        RECT 10.510 105.550 115.850 105.720 ;
        RECT 10.595 104.460 11.805 105.550 ;
        RECT 10.595 103.750 11.115 104.290 ;
        RECT 11.285 103.920 11.805 104.460 ;
        RECT 12.435 104.385 12.725 105.550 ;
        RECT 13.205 104.710 13.375 105.550 ;
        RECT 13.585 104.540 13.835 105.380 ;
        RECT 14.045 104.710 14.215 105.550 ;
        RECT 14.385 104.540 14.675 105.380 ;
        RECT 12.950 104.370 14.675 104.540 ;
        RECT 14.885 104.490 15.055 105.550 ;
        RECT 15.350 105.170 15.680 105.550 ;
        RECT 15.860 105.000 16.030 105.290 ;
        RECT 16.200 105.090 16.450 105.550 ;
        RECT 15.230 104.830 16.030 105.000 ;
        RECT 16.620 105.040 17.490 105.380 ;
        RECT 12.950 103.820 13.360 104.370 ;
        RECT 15.230 104.210 15.400 104.830 ;
        RECT 16.620 104.660 16.790 105.040 ;
        RECT 17.725 104.920 17.895 105.380 ;
        RECT 18.065 105.090 18.435 105.550 ;
        RECT 18.730 104.950 18.900 105.290 ;
        RECT 19.070 105.120 19.400 105.550 ;
        RECT 19.635 104.950 19.805 105.290 ;
        RECT 15.570 104.490 16.790 104.660 ;
        RECT 16.960 104.580 17.420 104.870 ;
        RECT 17.725 104.750 18.285 104.920 ;
        RECT 18.730 104.780 19.805 104.950 ;
        RECT 19.975 105.050 20.655 105.380 ;
        RECT 20.870 105.050 21.120 105.380 ;
        RECT 21.290 105.090 21.540 105.550 ;
        RECT 18.115 104.610 18.285 104.750 ;
        RECT 16.960 104.570 17.925 104.580 ;
        RECT 16.620 104.400 16.790 104.490 ;
        RECT 17.250 104.410 17.925 104.570 ;
        RECT 15.230 104.200 15.575 104.210 ;
        RECT 13.545 103.990 15.575 104.200 ;
        RECT 10.595 103.000 11.805 103.750 ;
        RECT 12.435 103.000 12.725 103.725 ;
        RECT 12.950 103.650 14.715 103.820 ;
        RECT 13.205 103.000 13.375 103.470 ;
        RECT 13.545 103.170 13.875 103.650 ;
        RECT 14.045 103.000 14.215 103.470 ;
        RECT 14.385 103.170 14.715 103.650 ;
        RECT 14.885 103.000 15.055 103.810 ;
        RECT 15.250 103.735 15.575 103.990 ;
        RECT 15.255 103.380 15.575 103.735 ;
        RECT 15.745 103.950 16.285 104.320 ;
        RECT 16.620 104.230 17.025 104.400 ;
        RECT 15.745 103.550 15.985 103.950 ;
        RECT 16.465 103.780 16.685 104.060 ;
        RECT 16.155 103.610 16.685 103.780 ;
        RECT 16.155 103.380 16.325 103.610 ;
        RECT 16.855 103.450 17.025 104.230 ;
        RECT 17.195 103.620 17.545 104.240 ;
        RECT 17.715 103.620 17.925 104.410 ;
        RECT 18.115 104.440 19.615 104.610 ;
        RECT 18.115 103.750 18.285 104.440 ;
        RECT 19.975 104.270 20.145 105.050 ;
        RECT 20.950 104.920 21.120 105.050 ;
        RECT 18.455 104.100 20.145 104.270 ;
        RECT 20.315 104.490 20.780 104.880 ;
        RECT 20.950 104.750 21.345 104.920 ;
        RECT 18.455 103.920 18.625 104.100 ;
        RECT 15.255 103.210 16.325 103.380 ;
        RECT 16.495 103.000 16.685 103.440 ;
        RECT 16.855 103.170 17.805 103.450 ;
        RECT 18.115 103.360 18.375 103.750 ;
        RECT 18.795 103.680 19.585 103.930 ;
        RECT 18.025 103.190 18.375 103.360 ;
        RECT 18.585 103.000 18.915 103.460 ;
        RECT 19.790 103.390 19.960 104.100 ;
        RECT 20.315 103.900 20.485 104.490 ;
        RECT 20.130 103.680 20.485 103.900 ;
        RECT 20.655 103.680 21.005 104.300 ;
        RECT 21.175 103.390 21.345 104.750 ;
        RECT 21.710 104.580 22.035 105.365 ;
        RECT 21.515 103.530 21.975 104.580 ;
        RECT 19.790 103.220 20.645 103.390 ;
        RECT 20.850 103.220 21.345 103.390 ;
        RECT 21.515 103.000 21.845 103.360 ;
        RECT 22.205 103.260 22.375 105.380 ;
        RECT 22.545 105.050 22.875 105.550 ;
        RECT 23.045 104.880 23.300 105.380 ;
        RECT 22.550 104.710 23.300 104.880 ;
        RECT 22.550 103.720 22.780 104.710 ;
        RECT 22.950 103.890 23.300 104.540 ;
        RECT 23.475 104.460 25.145 105.550 ;
        RECT 23.475 103.940 24.225 104.460 ;
        RECT 25.315 104.385 25.605 105.550 ;
        RECT 26.085 104.710 26.255 105.550 ;
        RECT 26.465 104.540 26.715 105.380 ;
        RECT 26.925 104.710 27.095 105.550 ;
        RECT 27.265 104.540 27.555 105.380 ;
        RECT 25.830 104.370 27.555 104.540 ;
        RECT 27.765 104.490 27.935 105.550 ;
        RECT 28.230 105.170 28.560 105.550 ;
        RECT 28.740 105.000 28.910 105.290 ;
        RECT 29.080 105.090 29.330 105.550 ;
        RECT 28.110 104.830 28.910 105.000 ;
        RECT 29.500 105.040 30.370 105.380 ;
        RECT 24.395 103.770 25.145 104.290 ;
        RECT 22.550 103.550 23.300 103.720 ;
        RECT 22.545 103.000 22.875 103.380 ;
        RECT 23.045 103.260 23.300 103.550 ;
        RECT 23.475 103.000 25.145 103.770 ;
        RECT 25.830 103.820 26.240 104.370 ;
        RECT 28.110 104.210 28.280 104.830 ;
        RECT 29.500 104.660 29.670 105.040 ;
        RECT 30.605 104.920 30.775 105.380 ;
        RECT 30.945 105.090 31.315 105.550 ;
        RECT 31.610 104.950 31.780 105.290 ;
        RECT 31.950 105.120 32.280 105.550 ;
        RECT 32.515 104.950 32.685 105.290 ;
        RECT 28.450 104.490 29.670 104.660 ;
        RECT 29.840 104.580 30.300 104.870 ;
        RECT 30.605 104.750 31.165 104.920 ;
        RECT 31.610 104.780 32.685 104.950 ;
        RECT 32.855 105.050 33.535 105.380 ;
        RECT 33.750 105.050 34.000 105.380 ;
        RECT 34.170 105.090 34.420 105.550 ;
        RECT 30.995 104.610 31.165 104.750 ;
        RECT 29.840 104.570 30.805 104.580 ;
        RECT 29.500 104.400 29.670 104.490 ;
        RECT 30.130 104.410 30.805 104.570 ;
        RECT 28.110 104.200 28.455 104.210 ;
        RECT 26.425 103.990 28.455 104.200 ;
        RECT 25.315 103.000 25.605 103.725 ;
        RECT 25.830 103.650 27.595 103.820 ;
        RECT 26.085 103.000 26.255 103.470 ;
        RECT 26.425 103.170 26.755 103.650 ;
        RECT 26.925 103.000 27.095 103.470 ;
        RECT 27.265 103.170 27.595 103.650 ;
        RECT 27.765 103.000 27.935 103.810 ;
        RECT 28.130 103.735 28.455 103.990 ;
        RECT 28.135 103.380 28.455 103.735 ;
        RECT 28.625 103.950 29.165 104.320 ;
        RECT 29.500 104.230 29.905 104.400 ;
        RECT 28.625 103.550 28.865 103.950 ;
        RECT 29.345 103.780 29.565 104.060 ;
        RECT 29.035 103.610 29.565 103.780 ;
        RECT 29.035 103.380 29.205 103.610 ;
        RECT 29.735 103.450 29.905 104.230 ;
        RECT 30.075 103.620 30.425 104.240 ;
        RECT 30.595 103.620 30.805 104.410 ;
        RECT 30.995 104.440 32.495 104.610 ;
        RECT 30.995 103.750 31.165 104.440 ;
        RECT 32.855 104.270 33.025 105.050 ;
        RECT 33.830 104.920 34.000 105.050 ;
        RECT 31.335 104.100 33.025 104.270 ;
        RECT 33.195 104.490 33.660 104.880 ;
        RECT 33.830 104.750 34.225 104.920 ;
        RECT 31.335 103.920 31.505 104.100 ;
        RECT 28.135 103.210 29.205 103.380 ;
        RECT 29.375 103.000 29.565 103.440 ;
        RECT 29.735 103.170 30.685 103.450 ;
        RECT 30.995 103.360 31.255 103.750 ;
        RECT 31.675 103.680 32.465 103.930 ;
        RECT 30.905 103.190 31.255 103.360 ;
        RECT 31.465 103.000 31.795 103.460 ;
        RECT 32.670 103.390 32.840 104.100 ;
        RECT 33.195 103.900 33.365 104.490 ;
        RECT 33.010 103.680 33.365 103.900 ;
        RECT 33.535 103.680 33.885 104.300 ;
        RECT 34.055 103.390 34.225 104.750 ;
        RECT 34.590 104.580 34.915 105.365 ;
        RECT 34.395 103.530 34.855 104.580 ;
        RECT 32.670 103.220 33.525 103.390 ;
        RECT 33.730 103.220 34.225 103.390 ;
        RECT 34.395 103.000 34.725 103.360 ;
        RECT 35.085 103.260 35.255 105.380 ;
        RECT 35.425 105.050 35.755 105.550 ;
        RECT 35.925 104.880 36.180 105.380 ;
        RECT 35.430 104.710 36.180 104.880 ;
        RECT 35.430 103.720 35.660 104.710 ;
        RECT 35.830 103.890 36.180 104.540 ;
        RECT 36.355 104.460 38.025 105.550 ;
        RECT 36.355 103.940 37.105 104.460 ;
        RECT 38.195 104.385 38.485 105.550 ;
        RECT 39.580 105.115 44.925 105.550 ;
        RECT 37.275 103.770 38.025 104.290 ;
        RECT 41.170 103.865 41.520 105.115 ;
        RECT 45.155 104.410 45.365 105.550 ;
        RECT 45.535 104.400 45.865 105.380 ;
        RECT 46.035 104.410 46.265 105.550 ;
        RECT 46.935 104.460 49.525 105.550 ;
        RECT 35.430 103.550 36.180 103.720 ;
        RECT 35.425 103.000 35.755 103.380 ;
        RECT 35.925 103.260 36.180 103.550 ;
        RECT 36.355 103.000 38.025 103.770 ;
        RECT 38.195 103.000 38.485 103.725 ;
        RECT 43.000 103.545 43.340 104.375 ;
        RECT 39.580 103.000 44.925 103.545 ;
        RECT 45.155 103.000 45.365 103.820 ;
        RECT 45.535 103.800 45.785 104.400 ;
        RECT 45.955 103.990 46.285 104.240 ;
        RECT 46.935 103.940 48.145 104.460 ;
        RECT 49.735 104.410 49.965 105.550 ;
        RECT 50.135 104.400 50.465 105.380 ;
        RECT 50.635 104.410 50.845 105.550 ;
        RECT 45.535 103.170 45.865 103.800 ;
        RECT 46.035 103.000 46.265 103.820 ;
        RECT 48.315 103.770 49.525 104.290 ;
        RECT 49.715 103.990 50.045 104.240 ;
        RECT 46.935 103.000 49.525 103.770 ;
        RECT 49.735 103.000 49.965 103.820 ;
        RECT 50.215 103.800 50.465 104.400 ;
        RECT 51.075 104.385 51.365 105.550 ;
        RECT 52.035 104.410 52.265 105.550 ;
        RECT 52.435 104.400 52.765 105.380 ;
        RECT 52.935 104.410 53.145 105.550 ;
        RECT 53.685 104.710 53.855 105.550 ;
        RECT 54.065 104.540 54.315 105.380 ;
        RECT 54.525 104.710 54.695 105.550 ;
        RECT 54.865 104.540 55.155 105.380 ;
        RECT 52.015 103.990 52.345 104.240 ;
        RECT 50.135 103.170 50.465 103.800 ;
        RECT 50.635 103.000 50.845 103.820 ;
        RECT 51.075 103.000 51.365 103.725 ;
        RECT 52.035 103.000 52.265 103.820 ;
        RECT 52.515 103.800 52.765 104.400 ;
        RECT 53.430 104.370 55.155 104.540 ;
        RECT 55.365 104.490 55.535 105.550 ;
        RECT 55.830 105.170 56.160 105.550 ;
        RECT 56.340 105.000 56.510 105.290 ;
        RECT 56.680 105.090 56.930 105.550 ;
        RECT 55.710 104.830 56.510 105.000 ;
        RECT 57.100 105.040 57.970 105.380 ;
        RECT 53.430 103.820 53.840 104.370 ;
        RECT 55.710 104.210 55.880 104.830 ;
        RECT 57.100 104.660 57.270 105.040 ;
        RECT 58.205 104.920 58.375 105.380 ;
        RECT 58.545 105.090 58.915 105.550 ;
        RECT 59.210 104.950 59.380 105.290 ;
        RECT 59.550 105.120 59.880 105.550 ;
        RECT 60.115 104.950 60.285 105.290 ;
        RECT 56.050 104.490 57.270 104.660 ;
        RECT 57.440 104.580 57.900 104.870 ;
        RECT 58.205 104.750 58.765 104.920 ;
        RECT 59.210 104.780 60.285 104.950 ;
        RECT 60.455 105.050 61.135 105.380 ;
        RECT 61.350 105.050 61.600 105.380 ;
        RECT 61.770 105.090 62.020 105.550 ;
        RECT 58.595 104.610 58.765 104.750 ;
        RECT 57.440 104.570 58.405 104.580 ;
        RECT 57.100 104.400 57.270 104.490 ;
        RECT 57.730 104.410 58.405 104.570 ;
        RECT 55.710 104.200 56.055 104.210 ;
        RECT 54.025 103.990 56.055 104.200 ;
        RECT 52.435 103.170 52.765 103.800 ;
        RECT 52.935 103.000 53.145 103.820 ;
        RECT 53.430 103.650 55.195 103.820 ;
        RECT 53.685 103.000 53.855 103.470 ;
        RECT 54.025 103.170 54.355 103.650 ;
        RECT 54.525 103.000 54.695 103.470 ;
        RECT 54.865 103.170 55.195 103.650 ;
        RECT 55.365 103.000 55.535 103.810 ;
        RECT 55.730 103.735 56.055 103.990 ;
        RECT 55.735 103.380 56.055 103.735 ;
        RECT 56.225 103.950 56.765 104.320 ;
        RECT 57.100 104.230 57.505 104.400 ;
        RECT 56.225 103.550 56.465 103.950 ;
        RECT 56.945 103.780 57.165 104.060 ;
        RECT 56.635 103.610 57.165 103.780 ;
        RECT 56.635 103.380 56.805 103.610 ;
        RECT 57.335 103.450 57.505 104.230 ;
        RECT 57.675 103.620 58.025 104.240 ;
        RECT 58.195 103.620 58.405 104.410 ;
        RECT 58.595 104.440 60.095 104.610 ;
        RECT 58.595 103.750 58.765 104.440 ;
        RECT 60.455 104.270 60.625 105.050 ;
        RECT 61.430 104.920 61.600 105.050 ;
        RECT 58.935 104.100 60.625 104.270 ;
        RECT 60.795 104.490 61.260 104.880 ;
        RECT 61.430 104.750 61.825 104.920 ;
        RECT 58.935 103.920 59.105 104.100 ;
        RECT 55.735 103.210 56.805 103.380 ;
        RECT 56.975 103.000 57.165 103.440 ;
        RECT 57.335 103.170 58.285 103.450 ;
        RECT 58.595 103.360 58.855 103.750 ;
        RECT 59.275 103.680 60.065 103.930 ;
        RECT 58.505 103.190 58.855 103.360 ;
        RECT 59.065 103.000 59.395 103.460 ;
        RECT 60.270 103.390 60.440 104.100 ;
        RECT 60.795 103.900 60.965 104.490 ;
        RECT 60.610 103.680 60.965 103.900 ;
        RECT 61.135 103.680 61.485 104.300 ;
        RECT 61.655 103.390 61.825 104.750 ;
        RECT 62.190 104.580 62.515 105.365 ;
        RECT 61.995 103.530 62.455 104.580 ;
        RECT 60.270 103.220 61.125 103.390 ;
        RECT 61.330 103.220 61.825 103.390 ;
        RECT 61.995 103.000 62.325 103.360 ;
        RECT 62.685 103.260 62.855 105.380 ;
        RECT 63.025 105.050 63.355 105.550 ;
        RECT 63.525 104.880 63.780 105.380 ;
        RECT 63.030 104.710 63.780 104.880 ;
        RECT 63.030 103.720 63.260 104.710 ;
        RECT 63.430 103.890 63.780 104.540 ;
        RECT 63.955 104.385 64.245 105.550 ;
        RECT 64.420 105.115 69.765 105.550 ;
        RECT 66.010 103.865 66.360 105.115 ;
        RECT 69.995 104.410 70.205 105.550 ;
        RECT 70.375 104.400 70.705 105.380 ;
        RECT 70.875 104.410 71.105 105.550 ;
        RECT 71.320 105.115 76.665 105.550 ;
        RECT 63.030 103.550 63.780 103.720 ;
        RECT 63.025 103.000 63.355 103.380 ;
        RECT 63.525 103.260 63.780 103.550 ;
        RECT 63.955 103.000 64.245 103.725 ;
        RECT 67.840 103.545 68.180 104.375 ;
        RECT 64.420 103.000 69.765 103.545 ;
        RECT 69.995 103.000 70.205 103.820 ;
        RECT 70.375 103.800 70.625 104.400 ;
        RECT 70.795 103.990 71.125 104.240 ;
        RECT 72.910 103.865 73.260 105.115 ;
        RECT 76.835 104.385 77.125 105.550 ;
        RECT 78.220 105.115 83.565 105.550 ;
        RECT 70.375 103.170 70.705 103.800 ;
        RECT 70.875 103.000 71.105 103.820 ;
        RECT 74.740 103.545 75.080 104.375 ;
        RECT 79.810 103.865 80.160 105.115 ;
        RECT 83.795 104.410 84.005 105.550 ;
        RECT 84.175 104.400 84.505 105.380 ;
        RECT 84.675 104.410 84.905 105.550 ;
        RECT 85.575 104.460 88.165 105.550 ;
        RECT 71.320 103.000 76.665 103.545 ;
        RECT 76.835 103.000 77.125 103.725 ;
        RECT 81.640 103.545 81.980 104.375 ;
        RECT 78.220 103.000 83.565 103.545 ;
        RECT 83.795 103.000 84.005 103.820 ;
        RECT 84.175 103.800 84.425 104.400 ;
        RECT 84.595 103.990 84.925 104.240 ;
        RECT 85.575 103.940 86.785 104.460 ;
        RECT 88.375 104.410 88.605 105.550 ;
        RECT 88.775 104.400 89.105 105.380 ;
        RECT 89.275 104.410 89.485 105.550 ;
        RECT 84.175 103.170 84.505 103.800 ;
        RECT 84.675 103.000 84.905 103.820 ;
        RECT 86.955 103.770 88.165 104.290 ;
        RECT 88.355 103.990 88.685 104.240 ;
        RECT 85.575 103.000 88.165 103.770 ;
        RECT 88.375 103.000 88.605 103.820 ;
        RECT 88.855 103.800 89.105 104.400 ;
        RECT 89.715 104.385 90.005 105.550 ;
        RECT 90.175 104.460 91.845 105.550 ;
        RECT 92.325 104.710 92.495 105.550 ;
        RECT 92.705 104.540 92.955 105.380 ;
        RECT 93.165 104.710 93.335 105.550 ;
        RECT 93.505 104.540 93.795 105.380 ;
        RECT 90.175 103.940 90.925 104.460 ;
        RECT 92.070 104.370 93.795 104.540 ;
        RECT 94.005 104.490 94.175 105.550 ;
        RECT 94.470 105.170 94.800 105.550 ;
        RECT 94.980 105.000 95.150 105.290 ;
        RECT 95.320 105.090 95.570 105.550 ;
        RECT 94.350 104.830 95.150 105.000 ;
        RECT 95.740 105.040 96.610 105.380 ;
        RECT 88.775 103.170 89.105 103.800 ;
        RECT 89.275 103.000 89.485 103.820 ;
        RECT 91.095 103.770 91.845 104.290 ;
        RECT 89.715 103.000 90.005 103.725 ;
        RECT 90.175 103.000 91.845 103.770 ;
        RECT 92.070 103.820 92.480 104.370 ;
        RECT 94.350 104.210 94.520 104.830 ;
        RECT 95.740 104.660 95.910 105.040 ;
        RECT 96.845 104.920 97.015 105.380 ;
        RECT 97.185 105.090 97.555 105.550 ;
        RECT 97.850 104.950 98.020 105.290 ;
        RECT 98.190 105.120 98.520 105.550 ;
        RECT 98.755 104.950 98.925 105.290 ;
        RECT 94.690 104.490 95.910 104.660 ;
        RECT 96.080 104.580 96.540 104.870 ;
        RECT 96.845 104.750 97.405 104.920 ;
        RECT 97.850 104.780 98.925 104.950 ;
        RECT 99.095 105.050 99.775 105.380 ;
        RECT 99.990 105.050 100.240 105.380 ;
        RECT 100.410 105.090 100.660 105.550 ;
        RECT 97.235 104.610 97.405 104.750 ;
        RECT 96.080 104.570 97.045 104.580 ;
        RECT 95.740 104.400 95.910 104.490 ;
        RECT 96.370 104.410 97.045 104.570 ;
        RECT 94.350 104.200 94.695 104.210 ;
        RECT 92.665 103.990 94.695 104.200 ;
        RECT 92.070 103.650 93.835 103.820 ;
        RECT 92.325 103.000 92.495 103.470 ;
        RECT 92.665 103.170 92.995 103.650 ;
        RECT 93.165 103.000 93.335 103.470 ;
        RECT 93.505 103.170 93.835 103.650 ;
        RECT 94.005 103.000 94.175 103.810 ;
        RECT 94.370 103.735 94.695 103.990 ;
        RECT 94.375 103.380 94.695 103.735 ;
        RECT 94.865 103.950 95.405 104.320 ;
        RECT 95.740 104.230 96.145 104.400 ;
        RECT 94.865 103.550 95.105 103.950 ;
        RECT 95.585 103.780 95.805 104.060 ;
        RECT 95.275 103.610 95.805 103.780 ;
        RECT 95.275 103.380 95.445 103.610 ;
        RECT 95.975 103.450 96.145 104.230 ;
        RECT 96.315 103.620 96.665 104.240 ;
        RECT 96.835 103.620 97.045 104.410 ;
        RECT 97.235 104.440 98.735 104.610 ;
        RECT 97.235 103.750 97.405 104.440 ;
        RECT 99.095 104.270 99.265 105.050 ;
        RECT 100.070 104.920 100.240 105.050 ;
        RECT 97.575 104.100 99.265 104.270 ;
        RECT 99.435 104.490 99.900 104.880 ;
        RECT 100.070 104.750 100.465 104.920 ;
        RECT 97.575 103.920 97.745 104.100 ;
        RECT 94.375 103.210 95.445 103.380 ;
        RECT 95.615 103.000 95.805 103.440 ;
        RECT 95.975 103.170 96.925 103.450 ;
        RECT 97.235 103.360 97.495 103.750 ;
        RECT 97.915 103.680 98.705 103.930 ;
        RECT 97.145 103.190 97.495 103.360 ;
        RECT 97.705 103.000 98.035 103.460 ;
        RECT 98.910 103.390 99.080 104.100 ;
        RECT 99.435 103.900 99.605 104.490 ;
        RECT 99.250 103.680 99.605 103.900 ;
        RECT 99.775 103.680 100.125 104.300 ;
        RECT 100.295 103.390 100.465 104.750 ;
        RECT 100.830 104.580 101.155 105.365 ;
        RECT 100.635 103.530 101.095 104.580 ;
        RECT 98.910 103.220 99.765 103.390 ;
        RECT 99.970 103.220 100.465 103.390 ;
        RECT 100.635 103.000 100.965 103.360 ;
        RECT 101.325 103.260 101.495 105.380 ;
        RECT 101.665 105.050 101.995 105.550 ;
        RECT 102.165 104.880 102.420 105.380 ;
        RECT 101.670 104.710 102.420 104.880 ;
        RECT 101.670 103.720 101.900 104.710 ;
        RECT 102.070 103.890 102.420 104.540 ;
        RECT 102.595 104.385 102.885 105.550 ;
        RECT 103.055 104.460 104.265 105.550 ;
        RECT 104.435 104.460 107.945 105.550 ;
        RECT 103.055 103.920 103.575 104.460 ;
        RECT 103.745 103.750 104.265 104.290 ;
        RECT 104.435 103.940 106.125 104.460 ;
        RECT 108.155 104.410 108.385 105.550 ;
        RECT 108.555 104.400 108.885 105.380 ;
        RECT 109.055 104.410 109.265 105.550 ;
        RECT 109.495 104.460 113.005 105.550 ;
        RECT 113.175 104.475 113.445 105.380 ;
        RECT 113.615 104.790 113.945 105.550 ;
        RECT 114.125 104.620 114.305 105.380 ;
        RECT 106.295 103.770 107.945 104.290 ;
        RECT 108.135 103.990 108.465 104.240 ;
        RECT 101.670 103.550 102.420 103.720 ;
        RECT 101.665 103.000 101.995 103.380 ;
        RECT 102.165 103.260 102.420 103.550 ;
        RECT 102.595 103.000 102.885 103.725 ;
        RECT 103.055 103.000 104.265 103.750 ;
        RECT 104.435 103.000 107.945 103.770 ;
        RECT 108.155 103.000 108.385 103.820 ;
        RECT 108.635 103.800 108.885 104.400 ;
        RECT 109.495 103.940 111.185 104.460 ;
        RECT 108.555 103.170 108.885 103.800 ;
        RECT 109.055 103.000 109.265 103.820 ;
        RECT 111.355 103.770 113.005 104.290 ;
        RECT 109.495 103.000 113.005 103.770 ;
        RECT 113.175 103.675 113.355 104.475 ;
        RECT 113.630 104.450 114.305 104.620 ;
        RECT 114.555 104.460 115.765 105.550 ;
        RECT 113.630 104.305 113.800 104.450 ;
        RECT 113.525 103.975 113.800 104.305 ;
        RECT 113.630 103.720 113.800 103.975 ;
        RECT 114.025 103.900 114.365 104.270 ;
        RECT 114.555 103.920 115.075 104.460 ;
        RECT 115.245 103.750 115.765 104.290 ;
        RECT 113.175 103.170 113.435 103.675 ;
        RECT 113.630 103.550 114.295 103.720 ;
        RECT 113.615 103.000 113.945 103.380 ;
        RECT 114.125 103.170 114.295 103.550 ;
        RECT 114.555 103.000 115.765 103.750 ;
        RECT 10.510 102.830 115.850 103.000 ;
        RECT 19.165 66.070 30.165 66.940 ;
        RECT 19.165 54.930 20.835 66.070 ;
        RECT 21.465 65.555 26.465 65.725 ;
        RECT 21.235 55.300 21.405 65.340 ;
        RECT 26.525 55.300 26.695 65.340 ;
        RECT 27.095 54.930 27.265 66.070 ;
        RECT 27.895 65.555 28.895 65.725 ;
        RECT 27.665 55.300 27.835 65.340 ;
        RECT 28.955 55.300 29.125 65.340 ;
        RECT 29.525 54.930 30.165 66.070 ;
        RECT 19.165 52.860 30.165 54.930 ;
        RECT 19.165 49.370 21.005 52.860 ;
        RECT 22.765 52.780 30.165 52.860 ;
        RECT 21.635 52.350 22.135 52.520 ;
        RECT 21.405 50.095 21.575 52.135 ;
        RECT 22.195 50.095 22.365 52.135 ;
        RECT 21.635 49.710 22.135 49.880 ;
        RECT 22.765 49.370 25.085 52.780 ;
        RECT 25.715 52.270 26.215 52.440 ;
        RECT 19.165 48.650 25.085 49.370 ;
        RECT 19.135 48.040 23.045 48.260 ;
        RECT 19.135 45.640 20.855 48.040 ;
        RECT 21.485 47.530 21.985 47.700 ;
        RECT 21.255 46.320 21.425 47.360 ;
        RECT 22.045 46.320 22.215 47.360 ;
        RECT 21.485 45.980 21.985 46.150 ;
        RECT 22.615 45.640 23.045 48.040 ;
        RECT 24.025 46.290 25.085 48.650 ;
        RECT 25.485 47.015 25.655 52.055 ;
        RECT 26.275 47.015 26.445 52.055 ;
        RECT 25.715 46.630 26.215 46.800 ;
        RECT 26.845 46.290 27.015 52.780 ;
        RECT 27.645 52.270 28.145 52.440 ;
        RECT 27.415 47.015 27.585 52.055 ;
        RECT 28.205 47.015 28.375 52.055 ;
        RECT 27.645 46.630 28.145 46.800 ;
        RECT 28.775 46.290 30.165 52.780 ;
        RECT 30.365 66.080 41.365 66.950 ;
        RECT 30.365 54.940 32.035 66.080 ;
        RECT 32.665 65.565 37.665 65.735 ;
        RECT 32.435 55.310 32.605 65.350 ;
        RECT 37.725 55.310 37.895 65.350 ;
        RECT 38.295 54.940 38.465 66.080 ;
        RECT 39.095 65.565 40.095 65.735 ;
        RECT 38.865 55.310 39.035 65.350 ;
        RECT 40.155 55.310 40.325 65.350 ;
        RECT 40.725 54.940 41.365 66.080 ;
        RECT 30.365 52.870 41.365 54.940 ;
        RECT 30.365 49.380 32.205 52.870 ;
        RECT 33.965 52.790 41.365 52.870 ;
        RECT 32.835 52.360 33.335 52.530 ;
        RECT 32.605 50.105 32.775 52.145 ;
        RECT 33.395 50.105 33.565 52.145 ;
        RECT 32.835 49.720 33.335 49.890 ;
        RECT 33.965 49.380 36.285 52.790 ;
        RECT 36.915 52.280 37.415 52.450 ;
        RECT 30.365 48.660 36.285 49.380 ;
        RECT 24.025 45.800 30.165 46.290 ;
        RECT 30.335 48.050 34.245 48.270 ;
        RECT 19.135 45.370 23.045 45.640 ;
        RECT 30.335 45.650 32.055 48.050 ;
        RECT 32.685 47.540 33.185 47.710 ;
        RECT 32.455 46.330 32.625 47.370 ;
        RECT 33.245 46.330 33.415 47.370 ;
        RECT 32.685 45.990 33.185 46.160 ;
        RECT 33.815 45.650 34.245 48.050 ;
        RECT 35.225 46.300 36.285 48.660 ;
        RECT 36.685 47.025 36.855 52.065 ;
        RECT 37.475 47.025 37.645 52.065 ;
        RECT 36.915 46.640 37.415 46.810 ;
        RECT 38.045 46.300 38.215 52.790 ;
        RECT 38.845 52.280 39.345 52.450 ;
        RECT 38.615 47.025 38.785 52.065 ;
        RECT 39.405 47.025 39.575 52.065 ;
        RECT 38.845 46.640 39.345 46.810 ;
        RECT 39.975 46.300 41.365 52.790 ;
        RECT 41.585 66.050 52.585 66.920 ;
        RECT 41.585 54.910 43.255 66.050 ;
        RECT 43.885 65.535 48.885 65.705 ;
        RECT 43.655 55.280 43.825 65.320 ;
        RECT 48.945 55.280 49.115 65.320 ;
        RECT 49.515 54.910 49.685 66.050 ;
        RECT 50.315 65.535 51.315 65.705 ;
        RECT 50.085 55.280 50.255 65.320 ;
        RECT 51.375 55.280 51.545 65.320 ;
        RECT 51.945 54.910 52.585 66.050 ;
        RECT 41.585 52.840 52.585 54.910 ;
        RECT 41.585 49.350 43.425 52.840 ;
        RECT 45.185 52.760 52.585 52.840 ;
        RECT 44.055 52.330 44.555 52.500 ;
        RECT 43.825 50.075 43.995 52.115 ;
        RECT 44.615 50.075 44.785 52.115 ;
        RECT 44.055 49.690 44.555 49.860 ;
        RECT 45.185 49.350 47.505 52.760 ;
        RECT 48.135 52.250 48.635 52.420 ;
        RECT 41.585 48.630 47.505 49.350 ;
        RECT 35.225 45.810 41.365 46.300 ;
        RECT 41.555 48.020 45.465 48.240 ;
        RECT 30.335 45.380 34.245 45.650 ;
        RECT 41.555 45.620 43.275 48.020 ;
        RECT 43.905 47.510 44.405 47.680 ;
        RECT 43.675 46.300 43.845 47.340 ;
        RECT 44.465 46.300 44.635 47.340 ;
        RECT 43.905 45.960 44.405 46.130 ;
        RECT 45.035 45.620 45.465 48.020 ;
        RECT 46.445 46.270 47.505 48.630 ;
        RECT 47.905 46.995 48.075 52.035 ;
        RECT 48.695 46.995 48.865 52.035 ;
        RECT 48.135 46.610 48.635 46.780 ;
        RECT 49.265 46.270 49.435 52.760 ;
        RECT 50.065 52.250 50.565 52.420 ;
        RECT 49.835 46.995 50.005 52.035 ;
        RECT 50.625 46.995 50.795 52.035 ;
        RECT 50.065 46.610 50.565 46.780 ;
        RECT 51.195 46.270 52.585 52.760 ;
        RECT 52.835 66.030 63.835 66.900 ;
        RECT 52.835 54.890 54.505 66.030 ;
        RECT 55.135 65.515 60.135 65.685 ;
        RECT 54.905 55.260 55.075 65.300 ;
        RECT 60.195 55.260 60.365 65.300 ;
        RECT 60.765 54.890 60.935 66.030 ;
        RECT 61.565 65.515 62.565 65.685 ;
        RECT 61.335 55.260 61.505 65.300 ;
        RECT 62.625 55.260 62.795 65.300 ;
        RECT 63.195 54.890 63.835 66.030 ;
        RECT 52.835 52.820 63.835 54.890 ;
        RECT 52.835 49.330 54.675 52.820 ;
        RECT 56.435 52.740 63.835 52.820 ;
        RECT 55.305 52.310 55.805 52.480 ;
        RECT 55.075 50.055 55.245 52.095 ;
        RECT 55.865 50.055 56.035 52.095 ;
        RECT 55.305 49.670 55.805 49.840 ;
        RECT 56.435 49.330 58.755 52.740 ;
        RECT 59.385 52.230 59.885 52.400 ;
        RECT 52.835 48.610 58.755 49.330 ;
        RECT 46.445 45.780 52.585 46.270 ;
        RECT 52.805 48.000 56.715 48.220 ;
        RECT 41.555 45.350 45.465 45.620 ;
        RECT 52.805 45.600 54.525 48.000 ;
        RECT 55.155 47.490 55.655 47.660 ;
        RECT 54.925 46.280 55.095 47.320 ;
        RECT 55.715 46.280 55.885 47.320 ;
        RECT 55.155 45.940 55.655 46.110 ;
        RECT 56.285 45.600 56.715 48.000 ;
        RECT 57.695 46.250 58.755 48.610 ;
        RECT 59.155 46.975 59.325 52.015 ;
        RECT 59.945 46.975 60.115 52.015 ;
        RECT 59.385 46.590 59.885 46.760 ;
        RECT 60.515 46.250 60.685 52.740 ;
        RECT 61.315 52.230 61.815 52.400 ;
        RECT 61.085 46.975 61.255 52.015 ;
        RECT 61.875 46.975 62.045 52.015 ;
        RECT 61.315 46.590 61.815 46.760 ;
        RECT 62.445 46.250 63.835 52.740 ;
        RECT 64.055 66.020 75.055 66.890 ;
        RECT 64.055 54.880 65.725 66.020 ;
        RECT 66.355 65.505 71.355 65.675 ;
        RECT 66.125 55.250 66.295 65.290 ;
        RECT 71.415 55.250 71.585 65.290 ;
        RECT 71.985 54.880 72.155 66.020 ;
        RECT 72.785 65.505 73.785 65.675 ;
        RECT 72.555 55.250 72.725 65.290 ;
        RECT 73.845 55.250 74.015 65.290 ;
        RECT 74.415 54.880 75.055 66.020 ;
        RECT 64.055 52.810 75.055 54.880 ;
        RECT 64.055 49.320 65.895 52.810 ;
        RECT 67.655 52.730 75.055 52.810 ;
        RECT 66.525 52.300 67.025 52.470 ;
        RECT 66.295 50.045 66.465 52.085 ;
        RECT 67.085 50.045 67.255 52.085 ;
        RECT 66.525 49.660 67.025 49.830 ;
        RECT 67.655 49.320 69.975 52.730 ;
        RECT 70.605 52.220 71.105 52.390 ;
        RECT 64.055 48.600 69.975 49.320 ;
        RECT 57.695 45.760 63.835 46.250 ;
        RECT 64.025 47.990 67.935 48.210 ;
        RECT 52.805 45.330 56.715 45.600 ;
        RECT 64.025 45.590 65.745 47.990 ;
        RECT 66.375 47.480 66.875 47.650 ;
        RECT 66.145 46.270 66.315 47.310 ;
        RECT 66.935 46.270 67.105 47.310 ;
        RECT 66.375 45.930 66.875 46.100 ;
        RECT 67.505 45.590 67.935 47.990 ;
        RECT 68.915 46.240 69.975 48.600 ;
        RECT 70.375 46.965 70.545 52.005 ;
        RECT 71.165 46.965 71.335 52.005 ;
        RECT 70.605 46.580 71.105 46.750 ;
        RECT 71.735 46.240 71.905 52.730 ;
        RECT 72.535 52.220 73.035 52.390 ;
        RECT 72.305 46.965 72.475 52.005 ;
        RECT 73.095 46.965 73.265 52.005 ;
        RECT 72.535 46.580 73.035 46.750 ;
        RECT 73.665 46.240 75.055 52.730 ;
        RECT 75.295 66.010 86.295 66.880 ;
        RECT 75.295 54.870 76.965 66.010 ;
        RECT 77.595 65.495 82.595 65.665 ;
        RECT 77.365 55.240 77.535 65.280 ;
        RECT 82.655 55.240 82.825 65.280 ;
        RECT 83.225 54.870 83.395 66.010 ;
        RECT 84.025 65.495 85.025 65.665 ;
        RECT 83.795 55.240 83.965 65.280 ;
        RECT 85.085 55.240 85.255 65.280 ;
        RECT 85.655 54.870 86.295 66.010 ;
        RECT 75.295 52.800 86.295 54.870 ;
        RECT 75.295 49.310 77.135 52.800 ;
        RECT 78.895 52.720 86.295 52.800 ;
        RECT 77.765 52.290 78.265 52.460 ;
        RECT 77.535 50.035 77.705 52.075 ;
        RECT 78.325 50.035 78.495 52.075 ;
        RECT 77.765 49.650 78.265 49.820 ;
        RECT 78.895 49.310 81.215 52.720 ;
        RECT 81.845 52.210 82.345 52.380 ;
        RECT 75.295 48.590 81.215 49.310 ;
        RECT 68.915 45.750 75.055 46.240 ;
        RECT 75.265 47.980 79.175 48.200 ;
        RECT 64.025 45.320 67.935 45.590 ;
        RECT 75.265 45.580 76.985 47.980 ;
        RECT 77.615 47.470 78.115 47.640 ;
        RECT 77.385 46.260 77.555 47.300 ;
        RECT 78.175 46.260 78.345 47.300 ;
        RECT 77.615 45.920 78.115 46.090 ;
        RECT 78.745 45.580 79.175 47.980 ;
        RECT 80.155 46.230 81.215 48.590 ;
        RECT 81.615 46.955 81.785 51.995 ;
        RECT 82.405 46.955 82.575 51.995 ;
        RECT 81.845 46.570 82.345 46.740 ;
        RECT 82.975 46.230 83.145 52.720 ;
        RECT 83.775 52.210 84.275 52.380 ;
        RECT 83.545 46.955 83.715 51.995 ;
        RECT 84.335 46.955 84.505 51.995 ;
        RECT 83.775 46.570 84.275 46.740 ;
        RECT 84.905 46.230 86.295 52.720 ;
        RECT 86.545 66.020 97.545 66.890 ;
        RECT 131.125 66.880 140.025 66.890 ;
        RECT 86.545 54.880 88.215 66.020 ;
        RECT 88.845 65.505 93.845 65.675 ;
        RECT 88.615 55.250 88.785 65.290 ;
        RECT 93.905 55.250 94.075 65.290 ;
        RECT 94.475 54.880 94.645 66.020 ;
        RECT 95.275 65.505 96.275 65.675 ;
        RECT 95.045 55.250 95.215 65.290 ;
        RECT 96.335 55.250 96.505 65.290 ;
        RECT 96.905 54.880 97.545 66.020 ;
        RECT 86.545 52.810 97.545 54.880 ;
        RECT 86.545 49.320 88.385 52.810 ;
        RECT 90.145 52.730 97.545 52.810 ;
        RECT 89.015 52.300 89.515 52.470 ;
        RECT 88.785 50.045 88.955 52.085 ;
        RECT 89.575 50.045 89.745 52.085 ;
        RECT 89.015 49.660 89.515 49.830 ;
        RECT 90.145 49.320 92.465 52.730 ;
        RECT 93.095 52.220 93.595 52.390 ;
        RECT 86.545 48.600 92.465 49.320 ;
        RECT 80.155 45.740 86.295 46.230 ;
        RECT 86.515 47.990 90.425 48.210 ;
        RECT 75.265 45.310 79.175 45.580 ;
        RECT 86.515 45.590 88.235 47.990 ;
        RECT 88.865 47.480 89.365 47.650 ;
        RECT 88.635 46.270 88.805 47.310 ;
        RECT 89.425 46.270 89.595 47.310 ;
        RECT 88.865 45.930 89.365 46.100 ;
        RECT 89.995 45.590 90.425 47.990 ;
        RECT 91.405 46.240 92.465 48.600 ;
        RECT 92.865 46.965 93.035 52.005 ;
        RECT 93.655 46.965 93.825 52.005 ;
        RECT 93.095 46.580 93.595 46.750 ;
        RECT 94.225 46.240 94.395 52.730 ;
        RECT 95.025 52.220 95.525 52.390 ;
        RECT 94.795 46.965 94.965 52.005 ;
        RECT 95.585 46.965 95.755 52.005 ;
        RECT 95.025 46.580 95.525 46.750 ;
        RECT 96.155 46.240 97.545 52.730 ;
        RECT 97.825 66.010 108.825 66.880 ;
        RECT 97.825 54.870 99.495 66.010 ;
        RECT 100.125 65.495 105.125 65.665 ;
        RECT 99.895 55.240 100.065 65.280 ;
        RECT 105.185 55.240 105.355 65.280 ;
        RECT 105.755 54.870 105.925 66.010 ;
        RECT 106.555 65.495 107.555 65.665 ;
        RECT 106.325 55.240 106.495 65.280 ;
        RECT 107.615 55.240 107.785 65.280 ;
        RECT 108.185 54.870 108.825 66.010 ;
        RECT 97.825 52.800 108.825 54.870 ;
        RECT 97.825 49.310 99.665 52.800 ;
        RECT 101.425 52.720 108.825 52.800 ;
        RECT 100.295 52.290 100.795 52.460 ;
        RECT 100.065 50.035 100.235 52.075 ;
        RECT 100.855 50.035 101.025 52.075 ;
        RECT 100.295 49.650 100.795 49.820 ;
        RECT 101.425 49.310 103.745 52.720 ;
        RECT 104.375 52.210 104.875 52.380 ;
        RECT 97.825 48.590 103.745 49.310 ;
        RECT 91.405 45.750 97.545 46.240 ;
        RECT 97.795 47.980 101.705 48.200 ;
        RECT 86.515 45.320 90.425 45.590 ;
        RECT 97.795 45.580 99.515 47.980 ;
        RECT 100.145 47.470 100.645 47.640 ;
        RECT 99.915 46.260 100.085 47.300 ;
        RECT 100.705 46.260 100.875 47.300 ;
        RECT 100.145 45.920 100.645 46.090 ;
        RECT 101.275 45.580 101.705 47.980 ;
        RECT 102.685 46.230 103.745 48.590 ;
        RECT 104.145 46.955 104.315 51.995 ;
        RECT 104.935 46.955 105.105 51.995 ;
        RECT 104.375 46.570 104.875 46.740 ;
        RECT 105.505 46.230 105.675 52.720 ;
        RECT 106.305 52.210 106.805 52.380 ;
        RECT 106.075 46.955 106.245 51.995 ;
        RECT 106.865 46.955 107.035 51.995 ;
        RECT 106.305 46.570 106.805 46.740 ;
        RECT 107.435 46.230 108.825 52.720 ;
        RECT 109.095 66.010 120.095 66.880 ;
        RECT 109.095 54.870 110.765 66.010 ;
        RECT 111.395 65.495 116.395 65.665 ;
        RECT 111.165 55.240 111.335 65.280 ;
        RECT 116.455 55.240 116.625 65.280 ;
        RECT 117.025 54.870 117.195 66.010 ;
        RECT 117.825 65.495 118.825 65.665 ;
        RECT 117.595 55.240 117.765 65.280 ;
        RECT 118.885 55.240 119.055 65.280 ;
        RECT 119.455 54.870 120.095 66.010 ;
        RECT 109.095 52.800 120.095 54.870 ;
        RECT 109.095 49.310 110.935 52.800 ;
        RECT 112.695 52.720 120.095 52.800 ;
        RECT 111.565 52.290 112.065 52.460 ;
        RECT 111.335 50.035 111.505 52.075 ;
        RECT 112.125 50.035 112.295 52.075 ;
        RECT 111.565 49.650 112.065 49.820 ;
        RECT 112.695 49.310 115.015 52.720 ;
        RECT 115.645 52.210 116.145 52.380 ;
        RECT 109.095 48.590 115.015 49.310 ;
        RECT 102.685 45.740 108.825 46.230 ;
        RECT 109.065 47.980 112.975 48.200 ;
        RECT 97.795 45.310 101.705 45.580 ;
        RECT 109.065 45.580 110.785 47.980 ;
        RECT 111.415 47.470 111.915 47.640 ;
        RECT 111.185 46.260 111.355 47.300 ;
        RECT 111.975 46.260 112.145 47.300 ;
        RECT 111.415 45.920 111.915 46.090 ;
        RECT 112.545 45.580 112.975 47.980 ;
        RECT 113.955 46.230 115.015 48.590 ;
        RECT 115.415 46.955 115.585 51.995 ;
        RECT 116.205 46.955 116.375 51.995 ;
        RECT 115.645 46.570 116.145 46.740 ;
        RECT 116.775 46.230 116.945 52.720 ;
        RECT 117.575 52.210 118.075 52.380 ;
        RECT 117.345 46.955 117.515 51.995 ;
        RECT 118.135 46.955 118.305 51.995 ;
        RECT 117.575 46.570 118.075 46.740 ;
        RECT 118.705 46.230 120.095 52.720 ;
        RECT 120.345 66.010 140.025 66.880 ;
        RECT 120.345 54.870 122.015 66.010 ;
        RECT 122.645 65.495 127.645 65.665 ;
        RECT 122.415 55.240 122.585 65.280 ;
        RECT 127.705 55.240 127.875 65.280 ;
        RECT 128.275 54.870 128.445 66.010 ;
        RECT 130.705 65.980 140.025 66.010 ;
        RECT 129.075 65.495 130.075 65.665 ;
        RECT 128.845 55.240 129.015 65.280 ;
        RECT 130.135 55.240 130.305 65.280 ;
        RECT 130.705 54.870 132.765 65.980 ;
        RECT 133.395 65.465 138.395 65.635 ;
        RECT 133.165 55.210 133.335 65.250 ;
        RECT 138.455 55.210 138.625 65.250 ;
        RECT 120.345 54.840 132.765 54.870 ;
        RECT 139.025 54.840 140.025 65.980 ;
        RECT 120.345 54.720 140.025 54.840 ;
        RECT 120.345 53.550 140.035 54.720 ;
        RECT 120.345 52.800 131.345 53.550 ;
        RECT 120.345 49.310 122.185 52.800 ;
        RECT 123.945 52.720 131.345 52.800 ;
        RECT 122.815 52.290 123.315 52.460 ;
        RECT 122.585 50.035 122.755 52.075 ;
        RECT 123.375 50.035 123.545 52.075 ;
        RECT 122.815 49.650 123.315 49.820 ;
        RECT 123.945 49.310 126.265 52.720 ;
        RECT 126.895 52.210 127.395 52.380 ;
        RECT 120.345 48.590 126.265 49.310 ;
        RECT 113.955 45.740 120.095 46.230 ;
        RECT 120.315 47.980 124.225 48.200 ;
        RECT 109.065 45.310 112.975 45.580 ;
        RECT 120.315 45.580 122.035 47.980 ;
        RECT 122.665 47.470 123.165 47.640 ;
        RECT 122.435 46.260 122.605 47.300 ;
        RECT 123.225 46.260 123.395 47.300 ;
        RECT 122.665 45.920 123.165 46.090 ;
        RECT 123.795 45.580 124.225 47.980 ;
        RECT 125.205 46.230 126.265 48.590 ;
        RECT 126.665 46.955 126.835 51.995 ;
        RECT 127.455 46.955 127.625 51.995 ;
        RECT 126.895 46.570 127.395 46.740 ;
        RECT 128.025 46.230 128.195 52.720 ;
        RECT 128.825 52.210 129.325 52.380 ;
        RECT 128.595 46.955 128.765 51.995 ;
        RECT 129.385 46.955 129.555 51.995 ;
        RECT 128.825 46.570 129.325 46.740 ;
        RECT 129.955 46.230 131.345 52.720 ;
        RECT 125.205 45.740 131.345 46.230 ;
        RECT 120.315 45.310 124.225 45.580 ;
        RECT 25.695 39.770 29.605 40.040 ;
        RECT 18.575 39.120 24.715 39.610 ;
        RECT 18.575 32.630 19.965 39.120 ;
        RECT 20.595 38.610 21.095 38.780 ;
        RECT 20.365 33.355 20.535 38.395 ;
        RECT 21.155 33.355 21.325 38.395 ;
        RECT 20.595 32.970 21.095 33.140 ;
        RECT 21.725 32.630 21.895 39.120 ;
        RECT 22.525 38.610 23.025 38.780 ;
        RECT 22.295 33.355 22.465 38.395 ;
        RECT 23.085 33.355 23.255 38.395 ;
        RECT 23.655 36.760 24.715 39.120 ;
        RECT 25.695 37.370 26.125 39.770 ;
        RECT 26.755 39.260 27.255 39.430 ;
        RECT 26.525 38.050 26.695 39.090 ;
        RECT 27.315 38.050 27.485 39.090 ;
        RECT 26.755 37.710 27.255 37.880 ;
        RECT 27.885 37.370 29.605 39.770 ;
        RECT 36.975 39.770 40.885 40.040 ;
        RECT 25.695 37.150 29.605 37.370 ;
        RECT 29.855 39.120 35.995 39.610 ;
        RECT 23.655 36.040 29.575 36.760 ;
        RECT 22.525 32.970 23.025 33.140 ;
        RECT 23.655 32.630 25.975 36.040 ;
        RECT 26.605 35.530 27.105 35.700 ;
        RECT 26.375 33.275 26.545 35.315 ;
        RECT 27.165 33.275 27.335 35.315 ;
        RECT 26.605 32.890 27.105 33.060 ;
        RECT 18.575 32.550 25.975 32.630 ;
        RECT 27.735 32.550 29.575 36.040 ;
        RECT 18.575 30.480 29.575 32.550 ;
        RECT 18.575 19.340 19.215 30.480 ;
        RECT 19.615 20.070 19.785 30.110 ;
        RECT 20.905 20.070 21.075 30.110 ;
        RECT 19.845 19.685 20.845 19.855 ;
        RECT 21.475 19.340 21.645 30.480 ;
        RECT 22.045 20.070 22.215 30.110 ;
        RECT 27.335 20.070 27.505 30.110 ;
        RECT 22.275 19.685 27.275 19.855 ;
        RECT 27.905 19.340 29.575 30.480 ;
        RECT 18.575 18.470 29.575 19.340 ;
        RECT 29.855 32.630 31.245 39.120 ;
        RECT 31.875 38.610 32.375 38.780 ;
        RECT 31.645 33.355 31.815 38.395 ;
        RECT 32.435 33.355 32.605 38.395 ;
        RECT 31.875 32.970 32.375 33.140 ;
        RECT 33.005 32.630 33.175 39.120 ;
        RECT 33.805 38.610 34.305 38.780 ;
        RECT 33.575 33.355 33.745 38.395 ;
        RECT 34.365 33.355 34.535 38.395 ;
        RECT 34.935 36.760 35.995 39.120 ;
        RECT 36.975 37.370 37.405 39.770 ;
        RECT 38.035 39.260 38.535 39.430 ;
        RECT 37.805 38.050 37.975 39.090 ;
        RECT 38.595 38.050 38.765 39.090 ;
        RECT 38.035 37.710 38.535 37.880 ;
        RECT 39.165 37.370 40.885 39.770 ;
        RECT 48.265 39.750 52.175 40.020 ;
        RECT 36.975 37.150 40.885 37.370 ;
        RECT 41.145 39.100 47.285 39.590 ;
        RECT 34.935 36.040 40.855 36.760 ;
        RECT 33.805 32.970 34.305 33.140 ;
        RECT 34.935 32.630 37.255 36.040 ;
        RECT 37.885 35.530 38.385 35.700 ;
        RECT 37.655 33.275 37.825 35.315 ;
        RECT 38.445 33.275 38.615 35.315 ;
        RECT 37.885 32.890 38.385 33.060 ;
        RECT 29.855 32.550 37.255 32.630 ;
        RECT 39.015 32.550 40.855 36.040 ;
        RECT 29.855 30.480 40.855 32.550 ;
        RECT 29.855 19.340 30.495 30.480 ;
        RECT 30.895 20.070 31.065 30.110 ;
        RECT 32.185 20.070 32.355 30.110 ;
        RECT 31.125 19.685 32.125 19.855 ;
        RECT 32.755 19.340 32.925 30.480 ;
        RECT 33.325 20.070 33.495 30.110 ;
        RECT 38.615 20.070 38.785 30.110 ;
        RECT 33.555 19.685 38.555 19.855 ;
        RECT 39.185 19.340 40.855 30.480 ;
        RECT 29.855 18.470 40.855 19.340 ;
        RECT 41.145 32.610 42.535 39.100 ;
        RECT 43.165 38.590 43.665 38.760 ;
        RECT 42.935 33.335 43.105 38.375 ;
        RECT 43.725 33.335 43.895 38.375 ;
        RECT 43.165 32.950 43.665 33.120 ;
        RECT 44.295 32.610 44.465 39.100 ;
        RECT 45.095 38.590 45.595 38.760 ;
        RECT 44.865 33.335 45.035 38.375 ;
        RECT 45.655 33.335 45.825 38.375 ;
        RECT 46.225 36.740 47.285 39.100 ;
        RECT 48.265 37.350 48.695 39.750 ;
        RECT 49.325 39.240 49.825 39.410 ;
        RECT 49.095 38.030 49.265 39.070 ;
        RECT 49.885 38.030 50.055 39.070 ;
        RECT 49.325 37.690 49.825 37.860 ;
        RECT 50.455 37.350 52.175 39.750 ;
        RECT 59.485 39.750 63.395 40.020 ;
        RECT 48.265 37.130 52.175 37.350 ;
        RECT 52.365 39.100 58.505 39.590 ;
        RECT 46.225 36.020 52.145 36.740 ;
        RECT 45.095 32.950 45.595 33.120 ;
        RECT 46.225 32.610 48.545 36.020 ;
        RECT 49.175 35.510 49.675 35.680 ;
        RECT 48.945 33.255 49.115 35.295 ;
        RECT 49.735 33.255 49.905 35.295 ;
        RECT 49.175 32.870 49.675 33.040 ;
        RECT 41.145 32.530 48.545 32.610 ;
        RECT 50.305 32.530 52.145 36.020 ;
        RECT 41.145 30.460 52.145 32.530 ;
        RECT 41.145 19.320 41.785 30.460 ;
        RECT 42.185 20.050 42.355 30.090 ;
        RECT 43.475 20.050 43.645 30.090 ;
        RECT 42.415 19.665 43.415 19.835 ;
        RECT 44.045 19.320 44.215 30.460 ;
        RECT 44.615 20.050 44.785 30.090 ;
        RECT 49.905 20.050 50.075 30.090 ;
        RECT 44.845 19.665 49.845 19.835 ;
        RECT 50.475 19.320 52.145 30.460 ;
        RECT 41.145 18.450 52.145 19.320 ;
        RECT 52.365 32.610 53.755 39.100 ;
        RECT 54.385 38.590 54.885 38.760 ;
        RECT 54.155 33.335 54.325 38.375 ;
        RECT 54.945 33.335 55.115 38.375 ;
        RECT 54.385 32.950 54.885 33.120 ;
        RECT 55.515 32.610 55.685 39.100 ;
        RECT 56.315 38.590 56.815 38.760 ;
        RECT 56.085 33.335 56.255 38.375 ;
        RECT 56.875 33.335 57.045 38.375 ;
        RECT 57.445 36.740 58.505 39.100 ;
        RECT 59.485 37.350 59.915 39.750 ;
        RECT 60.545 39.240 61.045 39.410 ;
        RECT 60.315 38.030 60.485 39.070 ;
        RECT 61.105 38.030 61.275 39.070 ;
        RECT 60.545 37.690 61.045 37.860 ;
        RECT 61.675 37.350 63.395 39.750 ;
        RECT 70.685 39.750 74.595 40.020 ;
        RECT 59.485 37.130 63.395 37.350 ;
        RECT 63.565 39.100 69.705 39.590 ;
        RECT 57.445 36.020 63.365 36.740 ;
        RECT 56.315 32.950 56.815 33.120 ;
        RECT 57.445 32.610 59.765 36.020 ;
        RECT 60.395 35.510 60.895 35.680 ;
        RECT 60.165 33.255 60.335 35.295 ;
        RECT 60.955 33.255 61.125 35.295 ;
        RECT 60.395 32.870 60.895 33.040 ;
        RECT 52.365 32.530 59.765 32.610 ;
        RECT 61.525 32.530 63.365 36.020 ;
        RECT 52.365 30.460 63.365 32.530 ;
        RECT 52.365 19.320 53.005 30.460 ;
        RECT 53.405 20.050 53.575 30.090 ;
        RECT 54.695 20.050 54.865 30.090 ;
        RECT 53.635 19.665 54.635 19.835 ;
        RECT 55.265 19.320 55.435 30.460 ;
        RECT 55.835 20.050 56.005 30.090 ;
        RECT 61.125 20.050 61.295 30.090 ;
        RECT 56.065 19.665 61.065 19.835 ;
        RECT 61.695 19.320 63.365 30.460 ;
        RECT 52.365 18.450 63.365 19.320 ;
        RECT 63.565 32.610 64.955 39.100 ;
        RECT 65.585 38.590 66.085 38.760 ;
        RECT 65.355 33.335 65.525 38.375 ;
        RECT 66.145 33.335 66.315 38.375 ;
        RECT 65.585 32.950 66.085 33.120 ;
        RECT 66.715 32.610 66.885 39.100 ;
        RECT 67.515 38.590 68.015 38.760 ;
        RECT 67.285 33.335 67.455 38.375 ;
        RECT 68.075 33.335 68.245 38.375 ;
        RECT 68.645 36.740 69.705 39.100 ;
        RECT 70.685 37.350 71.115 39.750 ;
        RECT 71.745 39.240 72.245 39.410 ;
        RECT 71.515 38.030 71.685 39.070 ;
        RECT 72.305 38.030 72.475 39.070 ;
        RECT 71.745 37.690 72.245 37.860 ;
        RECT 72.875 37.350 74.595 39.750 ;
        RECT 81.975 39.740 85.885 40.010 ;
        RECT 70.685 37.130 74.595 37.350 ;
        RECT 74.855 39.090 80.995 39.580 ;
        RECT 68.645 36.020 74.565 36.740 ;
        RECT 67.515 32.950 68.015 33.120 ;
        RECT 68.645 32.610 70.965 36.020 ;
        RECT 71.595 35.510 72.095 35.680 ;
        RECT 71.365 33.255 71.535 35.295 ;
        RECT 72.155 33.255 72.325 35.295 ;
        RECT 71.595 32.870 72.095 33.040 ;
        RECT 63.565 32.530 70.965 32.610 ;
        RECT 72.725 32.530 74.565 36.020 ;
        RECT 63.565 30.460 74.565 32.530 ;
        RECT 63.565 19.320 64.205 30.460 ;
        RECT 64.605 20.050 64.775 30.090 ;
        RECT 65.895 20.050 66.065 30.090 ;
        RECT 64.835 19.665 65.835 19.835 ;
        RECT 66.465 19.320 66.635 30.460 ;
        RECT 67.035 20.050 67.205 30.090 ;
        RECT 72.325 20.050 72.495 30.090 ;
        RECT 67.265 19.665 72.265 19.835 ;
        RECT 72.895 19.320 74.565 30.460 ;
        RECT 63.565 18.450 74.565 19.320 ;
        RECT 74.855 32.600 76.245 39.090 ;
        RECT 76.875 38.580 77.375 38.750 ;
        RECT 76.645 33.325 76.815 38.365 ;
        RECT 77.435 33.325 77.605 38.365 ;
        RECT 76.875 32.940 77.375 33.110 ;
        RECT 78.005 32.600 78.175 39.090 ;
        RECT 78.805 38.580 79.305 38.750 ;
        RECT 78.575 33.325 78.745 38.365 ;
        RECT 79.365 33.325 79.535 38.365 ;
        RECT 79.935 36.730 80.995 39.090 ;
        RECT 81.975 37.340 82.405 39.740 ;
        RECT 83.035 39.230 83.535 39.400 ;
        RECT 82.805 38.020 82.975 39.060 ;
        RECT 83.595 38.020 83.765 39.060 ;
        RECT 83.035 37.680 83.535 37.850 ;
        RECT 84.165 37.340 85.885 39.740 ;
        RECT 93.215 39.760 97.125 40.030 ;
        RECT 81.975 37.120 85.885 37.340 ;
        RECT 86.095 39.110 92.235 39.600 ;
        RECT 79.935 36.010 85.855 36.730 ;
        RECT 78.805 32.940 79.305 33.110 ;
        RECT 79.935 32.600 82.255 36.010 ;
        RECT 82.885 35.500 83.385 35.670 ;
        RECT 82.655 33.245 82.825 35.285 ;
        RECT 83.445 33.245 83.615 35.285 ;
        RECT 82.885 32.860 83.385 33.030 ;
        RECT 74.855 32.520 82.255 32.600 ;
        RECT 84.015 32.520 85.855 36.010 ;
        RECT 74.855 30.450 85.855 32.520 ;
        RECT 74.855 19.310 75.495 30.450 ;
        RECT 75.895 20.040 76.065 30.080 ;
        RECT 77.185 20.040 77.355 30.080 ;
        RECT 76.125 19.655 77.125 19.825 ;
        RECT 77.755 19.310 77.925 30.450 ;
        RECT 78.325 20.040 78.495 30.080 ;
        RECT 83.615 20.040 83.785 30.080 ;
        RECT 78.555 19.655 83.555 19.825 ;
        RECT 84.185 19.310 85.855 30.450 ;
        RECT 74.855 18.440 85.855 19.310 ;
        RECT 86.095 32.620 87.485 39.110 ;
        RECT 88.115 38.600 88.615 38.770 ;
        RECT 87.885 33.345 88.055 38.385 ;
        RECT 88.675 33.345 88.845 38.385 ;
        RECT 88.115 32.960 88.615 33.130 ;
        RECT 89.245 32.620 89.415 39.110 ;
        RECT 90.045 38.600 90.545 38.770 ;
        RECT 89.815 33.345 89.985 38.385 ;
        RECT 90.605 33.345 90.775 38.385 ;
        RECT 91.175 36.750 92.235 39.110 ;
        RECT 93.215 37.360 93.645 39.760 ;
        RECT 94.275 39.250 94.775 39.420 ;
        RECT 94.045 38.040 94.215 39.080 ;
        RECT 94.835 38.040 95.005 39.080 ;
        RECT 94.275 37.700 94.775 37.870 ;
        RECT 95.405 37.360 97.125 39.760 ;
        RECT 104.425 39.780 108.335 40.050 ;
        RECT 93.215 37.140 97.125 37.360 ;
        RECT 97.305 39.130 103.445 39.620 ;
        RECT 91.175 36.030 97.095 36.750 ;
        RECT 90.045 32.960 90.545 33.130 ;
        RECT 91.175 32.620 93.495 36.030 ;
        RECT 94.125 35.520 94.625 35.690 ;
        RECT 93.895 33.265 94.065 35.305 ;
        RECT 94.685 33.265 94.855 35.305 ;
        RECT 94.125 32.880 94.625 33.050 ;
        RECT 86.095 32.540 93.495 32.620 ;
        RECT 95.255 32.540 97.095 36.030 ;
        RECT 86.095 30.470 97.095 32.540 ;
        RECT 86.095 19.330 86.735 30.470 ;
        RECT 87.135 20.060 87.305 30.100 ;
        RECT 88.425 20.060 88.595 30.100 ;
        RECT 87.365 19.675 88.365 19.845 ;
        RECT 88.995 19.330 89.165 30.470 ;
        RECT 89.565 20.060 89.735 30.100 ;
        RECT 94.855 20.060 95.025 30.100 ;
        RECT 89.795 19.675 94.795 19.845 ;
        RECT 95.425 19.330 97.095 30.470 ;
        RECT 86.095 18.460 97.095 19.330 ;
        RECT 97.305 32.640 98.695 39.130 ;
        RECT 99.325 38.620 99.825 38.790 ;
        RECT 99.095 33.365 99.265 38.405 ;
        RECT 99.885 33.365 100.055 38.405 ;
        RECT 99.325 32.980 99.825 33.150 ;
        RECT 100.455 32.640 100.625 39.130 ;
        RECT 101.255 38.620 101.755 38.790 ;
        RECT 101.025 33.365 101.195 38.405 ;
        RECT 101.815 33.365 101.985 38.405 ;
        RECT 102.385 36.770 103.445 39.130 ;
        RECT 104.425 37.380 104.855 39.780 ;
        RECT 105.485 39.270 105.985 39.440 ;
        RECT 105.255 38.060 105.425 39.100 ;
        RECT 106.045 38.060 106.215 39.100 ;
        RECT 105.485 37.720 105.985 37.890 ;
        RECT 106.615 37.380 108.335 39.780 ;
        RECT 115.625 39.820 119.535 40.090 ;
        RECT 104.425 37.160 108.335 37.380 ;
        RECT 108.505 39.170 114.645 39.660 ;
        RECT 102.385 36.050 108.305 36.770 ;
        RECT 101.255 32.980 101.755 33.150 ;
        RECT 102.385 32.640 104.705 36.050 ;
        RECT 105.335 35.540 105.835 35.710 ;
        RECT 105.105 33.285 105.275 35.325 ;
        RECT 105.895 33.285 106.065 35.325 ;
        RECT 105.335 32.900 105.835 33.070 ;
        RECT 97.305 32.560 104.705 32.640 ;
        RECT 106.465 32.560 108.305 36.050 ;
        RECT 97.305 30.490 108.305 32.560 ;
        RECT 97.305 19.350 97.945 30.490 ;
        RECT 98.345 20.080 98.515 30.120 ;
        RECT 99.635 20.080 99.805 30.120 ;
        RECT 98.575 19.695 99.575 19.865 ;
        RECT 100.205 19.350 100.375 30.490 ;
        RECT 100.775 20.080 100.945 30.120 ;
        RECT 106.065 20.080 106.235 30.120 ;
        RECT 101.005 19.695 106.005 19.865 ;
        RECT 106.635 19.350 108.305 30.490 ;
        RECT 97.305 18.480 108.305 19.350 ;
        RECT 108.505 32.680 109.895 39.170 ;
        RECT 110.525 38.660 111.025 38.830 ;
        RECT 110.295 33.405 110.465 38.445 ;
        RECT 111.085 33.405 111.255 38.445 ;
        RECT 110.525 33.020 111.025 33.190 ;
        RECT 111.655 32.680 111.825 39.170 ;
        RECT 112.455 38.660 112.955 38.830 ;
        RECT 112.225 33.405 112.395 38.445 ;
        RECT 113.015 33.405 113.185 38.445 ;
        RECT 113.585 36.810 114.645 39.170 ;
        RECT 115.625 37.420 116.055 39.820 ;
        RECT 116.685 39.310 117.185 39.480 ;
        RECT 116.455 38.100 116.625 39.140 ;
        RECT 117.245 38.100 117.415 39.140 ;
        RECT 116.685 37.760 117.185 37.930 ;
        RECT 117.815 37.420 119.535 39.820 ;
        RECT 126.835 39.840 130.745 40.110 ;
        RECT 115.625 37.200 119.535 37.420 ;
        RECT 119.715 39.190 125.855 39.680 ;
        RECT 113.585 36.090 119.505 36.810 ;
        RECT 112.455 33.020 112.955 33.190 ;
        RECT 113.585 32.680 115.905 36.090 ;
        RECT 116.535 35.580 117.035 35.750 ;
        RECT 116.305 33.325 116.475 35.365 ;
        RECT 117.095 33.325 117.265 35.365 ;
        RECT 116.535 32.940 117.035 33.110 ;
        RECT 108.505 32.600 115.905 32.680 ;
        RECT 117.665 32.600 119.505 36.090 ;
        RECT 108.505 30.530 119.505 32.600 ;
        RECT 108.505 19.390 109.145 30.530 ;
        RECT 109.545 20.120 109.715 30.160 ;
        RECT 110.835 20.120 111.005 30.160 ;
        RECT 109.775 19.735 110.775 19.905 ;
        RECT 111.405 19.390 111.575 30.530 ;
        RECT 111.975 20.120 112.145 30.160 ;
        RECT 117.265 20.120 117.435 30.160 ;
        RECT 112.205 19.735 117.205 19.905 ;
        RECT 117.835 19.390 119.505 30.530 ;
        RECT 108.505 18.520 119.505 19.390 ;
        RECT 119.715 32.700 121.105 39.190 ;
        RECT 121.735 38.680 122.235 38.850 ;
        RECT 121.505 33.425 121.675 38.465 ;
        RECT 122.295 33.425 122.465 38.465 ;
        RECT 121.735 33.040 122.235 33.210 ;
        RECT 122.865 32.700 123.035 39.190 ;
        RECT 123.665 38.680 124.165 38.850 ;
        RECT 123.435 33.425 123.605 38.465 ;
        RECT 124.225 33.425 124.395 38.465 ;
        RECT 124.795 36.830 125.855 39.190 ;
        RECT 126.835 37.440 127.265 39.840 ;
        RECT 127.895 39.330 128.395 39.500 ;
        RECT 127.665 38.120 127.835 39.160 ;
        RECT 128.455 38.120 128.625 39.160 ;
        RECT 127.895 37.780 128.395 37.950 ;
        RECT 129.025 37.440 130.745 39.840 ;
        RECT 126.835 37.220 130.745 37.440 ;
        RECT 124.795 36.110 130.715 36.830 ;
        RECT 123.665 33.040 124.165 33.210 ;
        RECT 124.795 32.700 127.115 36.110 ;
        RECT 127.745 35.600 128.245 35.770 ;
        RECT 127.515 33.345 127.685 35.385 ;
        RECT 128.305 33.345 128.475 35.385 ;
        RECT 127.745 32.960 128.245 33.130 ;
        RECT 119.715 32.620 127.115 32.700 ;
        RECT 128.875 32.620 130.715 36.110 ;
        RECT 119.715 31.140 130.715 32.620 ;
        RECT 119.715 30.550 139.465 31.140 ;
        RECT 119.715 19.410 120.355 30.550 ;
        RECT 120.755 20.140 120.925 30.180 ;
        RECT 122.045 20.140 122.215 30.180 ;
        RECT 120.985 19.755 121.985 19.925 ;
        RECT 122.615 19.410 122.785 30.550 ;
        RECT 129.045 30.520 139.465 30.550 ;
        RECT 123.185 20.140 123.355 30.180 ;
        RECT 128.475 20.140 128.645 30.180 ;
        RECT 123.415 19.755 128.415 19.925 ;
        RECT 129.045 19.410 132.075 30.520 ;
        RECT 132.475 20.110 132.645 30.150 ;
        RECT 137.765 20.110 137.935 30.150 ;
        RECT 132.705 19.725 137.705 19.895 ;
        RECT 119.715 19.380 132.075 19.410 ;
        RECT 138.335 19.380 139.465 30.520 ;
        RECT 119.715 18.540 139.465 19.380 ;
        RECT 131.925 18.520 139.465 18.540 ;
      LAYER met1 ;
        RECT 135.340 223.880 136.790 225.180 ;
        RECT 10.510 206.035 115.850 206.515 ;
        RECT 59.340 205.155 59.660 205.215 ;
        RECT 66.255 205.155 66.545 205.200 ;
        RECT 59.340 205.015 66.545 205.155 ;
        RECT 59.340 204.955 59.660 205.015 ;
        RECT 66.255 204.970 66.545 205.015 ;
        RECT 66.700 203.935 67.020 204.195 ;
        RECT 10.510 203.315 115.850 203.795 ;
        RECT 60.720 203.115 61.040 203.175 ;
        RECT 62.575 203.115 62.865 203.160 ;
        RECT 60.720 202.975 62.865 203.115 ;
        RECT 60.720 202.915 61.040 202.975 ;
        RECT 62.575 202.930 62.865 202.975 ;
        RECT 61.655 202.590 61.945 202.820 ;
        RECT 67.275 202.775 67.565 202.820 ;
        RECT 70.395 202.775 70.685 202.820 ;
        RECT 72.285 202.775 72.575 202.820 ;
        RECT 67.275 202.635 72.575 202.775 ;
        RECT 67.275 202.590 67.565 202.635 ;
        RECT 70.395 202.590 70.685 202.635 ;
        RECT 72.285 202.590 72.575 202.635 ;
        RECT 57.055 202.095 57.345 202.140 ;
        RECT 59.340 202.095 59.660 202.155 ;
        RECT 57.055 201.955 59.660 202.095 ;
        RECT 57.055 201.910 57.345 201.955 ;
        RECT 59.340 201.895 59.660 201.955 ;
        RECT 61.195 202.095 61.485 202.140 ;
        RECT 61.730 202.095 61.870 202.590 ;
        RECT 63.940 202.435 64.260 202.495 ;
        RECT 64.415 202.435 64.705 202.480 ;
        RECT 63.940 202.295 64.705 202.435 ;
        RECT 63.940 202.235 64.260 202.295 ;
        RECT 64.415 202.250 64.705 202.295 ;
        RECT 61.195 201.955 61.870 202.095 ;
        RECT 61.195 201.910 61.485 201.955 ;
        RECT 63.480 201.555 63.800 201.815 ;
        RECT 66.195 201.800 66.485 202.115 ;
        RECT 67.275 202.095 67.565 202.140 ;
        RECT 70.855 202.095 71.145 202.140 ;
        RECT 72.690 202.095 72.980 202.140 ;
        RECT 67.275 201.955 72.980 202.095 ;
        RECT 67.275 201.910 67.565 201.955 ;
        RECT 70.855 201.910 71.145 201.955 ;
        RECT 72.690 201.910 72.980 201.955 ;
        RECT 73.155 202.095 73.445 202.140 ;
        RECT 76.360 202.095 76.680 202.155 ;
        RECT 73.155 201.955 76.680 202.095 ;
        RECT 73.155 201.910 73.445 201.955 ;
        RECT 76.360 201.895 76.680 201.955 ;
        RECT 76.835 201.910 77.125 202.140 ;
        RECT 65.895 201.755 66.485 201.800 ;
        RECT 66.700 201.755 67.020 201.815 ;
        RECT 69.135 201.755 69.785 201.800 ;
        RECT 65.895 201.615 69.785 201.755 ;
        RECT 65.895 201.570 66.185 201.615 ;
        RECT 66.700 201.555 67.020 201.615 ;
        RECT 69.135 201.570 69.785 201.615 ;
        RECT 71.300 201.755 71.620 201.815 ;
        RECT 71.775 201.755 72.065 201.800 ;
        RECT 71.300 201.615 72.065 201.755 ;
        RECT 71.300 201.555 71.620 201.615 ;
        RECT 71.775 201.570 72.065 201.615 ;
        RECT 73.600 201.755 73.920 201.815 ;
        RECT 76.910 201.755 77.050 201.910 ;
        RECT 73.600 201.615 77.050 201.755 ;
        RECT 73.600 201.555 73.920 201.615 ;
        RECT 56.580 201.215 56.900 201.475 ;
        RECT 60.260 201.215 60.580 201.475 ;
        RECT 62.495 201.415 62.785 201.460 ;
        RECT 64.400 201.415 64.720 201.475 ;
        RECT 62.495 201.275 64.720 201.415 ;
        RECT 62.495 201.230 62.785 201.275 ;
        RECT 64.400 201.215 64.720 201.275 ;
        RECT 74.980 201.415 75.300 201.475 ;
        RECT 75.915 201.415 76.205 201.460 ;
        RECT 74.980 201.275 76.205 201.415 ;
        RECT 74.980 201.215 75.300 201.275 ;
        RECT 75.915 201.230 76.205 201.275 ;
        RECT 10.510 200.595 115.850 201.075 ;
        RECT 58.880 200.395 59.200 200.455 ;
        RECT 63.480 200.395 63.800 200.455 ;
        RECT 65.320 200.395 65.640 200.455 ;
        RECT 77.755 200.395 78.045 200.440 ;
        RECT 53.910 200.255 62.790 200.395 ;
        RECT 51.535 200.055 51.825 200.100 ;
        RECT 53.910 200.055 54.050 200.255 ;
        RECT 58.880 200.195 59.200 200.255 ;
        RECT 51.535 199.915 54.050 200.055 ;
        RECT 54.395 200.055 54.685 200.100 ;
        RECT 56.580 200.055 56.900 200.115 ;
        RECT 57.635 200.055 58.285 200.100 ;
        RECT 54.395 199.915 58.285 200.055 ;
        RECT 51.535 199.870 51.825 199.915 ;
        RECT 54.395 199.870 54.985 199.915 ;
        RECT 54.695 199.555 54.985 199.870 ;
        RECT 56.580 199.855 56.900 199.915 ;
        RECT 57.635 199.870 58.285 199.915 ;
        RECT 60.260 199.855 60.580 200.115 ;
        RECT 62.650 199.760 62.790 200.255 ;
        RECT 63.480 200.255 65.640 200.395 ;
        RECT 63.480 200.195 63.800 200.255 ;
        RECT 65.320 200.195 65.640 200.255 ;
        RECT 74.610 200.255 78.045 200.395 ;
        RECT 63.940 200.055 64.260 200.115 ;
        RECT 69.115 200.055 69.405 200.100 ;
        RECT 72.355 200.055 73.005 200.100 ;
        RECT 74.610 200.055 74.750 200.255 ;
        RECT 77.755 200.210 78.045 200.255 ;
        RECT 63.940 199.915 65.090 200.055 ;
        RECT 63.940 199.855 64.260 199.915 ;
        RECT 64.950 199.775 65.090 199.915 ;
        RECT 69.115 199.915 74.750 200.055 ;
        RECT 69.115 199.870 69.705 199.915 ;
        RECT 72.355 199.870 73.005 199.915 ;
        RECT 55.775 199.715 56.065 199.760 ;
        RECT 59.355 199.715 59.645 199.760 ;
        RECT 61.190 199.715 61.480 199.760 ;
        RECT 55.775 199.575 61.480 199.715 ;
        RECT 55.775 199.530 56.065 199.575 ;
        RECT 59.355 199.530 59.645 199.575 ;
        RECT 61.190 199.530 61.480 199.575 ;
        RECT 62.575 199.715 62.865 199.760 ;
        RECT 64.860 199.715 65.180 199.775 ;
        RECT 65.795 199.715 66.085 199.760 ;
        RECT 62.575 199.575 64.630 199.715 ;
        RECT 62.575 199.530 62.865 199.575 ;
        RECT 52.900 199.375 53.220 199.435 ;
        RECT 61.655 199.375 61.945 199.420 ;
        RECT 52.900 199.235 61.945 199.375 ;
        RECT 52.900 199.175 53.220 199.235 ;
        RECT 61.655 199.190 61.945 199.235 ;
        RECT 63.940 199.175 64.260 199.435 ;
        RECT 64.490 199.375 64.630 199.575 ;
        RECT 64.860 199.575 66.085 199.715 ;
        RECT 64.860 199.515 65.180 199.575 ;
        RECT 65.795 199.530 66.085 199.575 ;
        RECT 69.415 199.555 69.705 199.870 ;
        RECT 74.980 199.855 75.300 200.115 ;
        RECT 70.495 199.715 70.785 199.760 ;
        RECT 74.075 199.715 74.365 199.760 ;
        RECT 75.910 199.715 76.200 199.760 ;
        RECT 70.495 199.575 76.200 199.715 ;
        RECT 70.495 199.530 70.785 199.575 ;
        RECT 74.075 199.530 74.365 199.575 ;
        RECT 75.910 199.530 76.200 199.575 ;
        RECT 76.360 199.515 76.680 199.775 ;
        RECT 78.200 199.515 78.520 199.775 ;
        RECT 68.080 199.375 68.400 199.435 ;
        RECT 64.490 199.235 68.400 199.375 ;
        RECT 68.080 199.175 68.400 199.235 ;
        RECT 55.775 199.035 56.065 199.080 ;
        RECT 58.895 199.035 59.185 199.080 ;
        RECT 60.785 199.035 61.075 199.080 ;
        RECT 55.775 198.895 61.075 199.035 ;
        RECT 55.775 198.850 56.065 198.895 ;
        RECT 58.895 198.850 59.185 198.895 ;
        RECT 60.785 198.850 61.075 198.895 ;
        RECT 66.715 199.035 67.005 199.080 ;
        RECT 69.460 199.035 69.780 199.095 ;
        RECT 66.715 198.895 69.780 199.035 ;
        RECT 66.715 198.850 67.005 198.895 ;
        RECT 63.020 198.695 63.340 198.755 ;
        RECT 64.415 198.695 64.705 198.740 ;
        RECT 66.790 198.695 66.930 198.850 ;
        RECT 69.460 198.835 69.780 198.895 ;
        RECT 70.495 199.035 70.785 199.080 ;
        RECT 73.615 199.035 73.905 199.080 ;
        RECT 75.505 199.035 75.795 199.080 ;
        RECT 70.495 198.895 75.795 199.035 ;
        RECT 70.495 198.850 70.785 198.895 ;
        RECT 73.615 198.850 73.905 198.895 ;
        RECT 75.505 198.850 75.795 198.895 ;
        RECT 63.020 198.555 66.930 198.695 ;
        RECT 67.160 198.695 67.480 198.755 ;
        RECT 67.635 198.695 67.925 198.740 ;
        RECT 67.160 198.555 67.925 198.695 ;
        RECT 63.020 198.495 63.340 198.555 ;
        RECT 64.415 198.510 64.705 198.555 ;
        RECT 67.160 198.495 67.480 198.555 ;
        RECT 67.635 198.510 67.925 198.555 ;
        RECT 10.510 197.875 115.850 198.355 ;
        RECT 52.900 197.675 53.220 197.735 ;
        RECT 50.230 197.535 53.220 197.675 ;
        RECT 49.695 196.995 49.985 197.040 ;
        RECT 50.230 196.995 50.370 197.535 ;
        RECT 52.900 197.475 53.220 197.535 ;
        RECT 64.400 197.475 64.720 197.735 ;
        RECT 70.855 197.675 71.145 197.720 ;
        RECT 71.300 197.675 71.620 197.735 ;
        RECT 70.855 197.535 71.620 197.675 ;
        RECT 70.855 197.490 71.145 197.535 ;
        RECT 71.300 197.475 71.620 197.535 ;
        RECT 50.565 197.335 50.855 197.380 ;
        RECT 52.455 197.335 52.745 197.380 ;
        RECT 55.575 197.335 55.865 197.380 ;
        RECT 50.565 197.195 55.865 197.335 ;
        RECT 50.565 197.150 50.855 197.195 ;
        RECT 52.455 197.150 52.745 197.195 ;
        RECT 55.575 197.150 55.865 197.195 ;
        RECT 59.355 197.150 59.645 197.380 ;
        RECT 63.035 197.335 63.325 197.380 ;
        RECT 74.635 197.335 74.925 197.380 ;
        RECT 77.755 197.335 78.045 197.380 ;
        RECT 79.645 197.335 79.935 197.380 ;
        RECT 63.035 197.195 69.230 197.335 ;
        RECT 63.035 197.150 63.325 197.195 ;
        RECT 49.695 196.855 50.370 196.995 ;
        RECT 51.075 196.995 51.365 197.040 ;
        RECT 59.430 196.995 59.570 197.150 ;
        RECT 51.075 196.855 59.570 196.995 ;
        RECT 60.260 196.995 60.580 197.055 ;
        RECT 60.735 196.995 61.025 197.040 ;
        RECT 65.780 196.995 66.100 197.055 ;
        RECT 69.090 197.040 69.230 197.195 ;
        RECT 74.635 197.195 79.935 197.335 ;
        RECT 74.635 197.150 74.925 197.195 ;
        RECT 77.755 197.150 78.045 197.195 ;
        RECT 79.645 197.150 79.935 197.195 ;
        RECT 60.260 196.855 61.025 196.995 ;
        RECT 49.695 196.810 49.985 196.855 ;
        RECT 51.075 196.810 51.365 196.855 ;
        RECT 60.260 196.795 60.580 196.855 ;
        RECT 60.735 196.810 61.025 196.855 ;
        RECT 63.110 196.855 64.630 196.995 ;
        RECT 65.590 196.855 66.100 196.995 ;
        RECT 63.110 196.715 63.250 196.855 ;
        RECT 50.160 196.655 50.450 196.700 ;
        RECT 51.995 196.655 52.285 196.700 ;
        RECT 55.575 196.655 55.865 196.700 ;
        RECT 50.160 196.515 55.865 196.655 ;
        RECT 50.160 196.470 50.450 196.515 ;
        RECT 51.995 196.470 52.285 196.515 ;
        RECT 55.575 196.470 55.865 196.515 ;
        RECT 53.355 196.315 54.005 196.360 ;
        RECT 54.740 196.315 55.060 196.375 ;
        RECT 56.655 196.360 56.945 196.675 ;
        RECT 61.180 196.455 61.500 196.715 ;
        RECT 62.575 196.470 62.865 196.700 ;
        RECT 56.655 196.315 57.245 196.360 ;
        RECT 53.355 196.175 57.245 196.315 ;
        RECT 53.355 196.130 54.005 196.175 ;
        RECT 54.740 196.115 55.060 196.175 ;
        RECT 56.955 196.130 57.245 196.175 ;
        RECT 60.720 196.315 61.040 196.375 ;
        RECT 62.650 196.315 62.790 196.470 ;
        RECT 63.020 196.455 63.340 196.715 ;
        RECT 63.480 196.455 63.800 196.715 ;
        RECT 64.490 196.605 64.630 196.855 ;
        RECT 65.780 196.795 66.100 196.855 ;
        RECT 69.015 196.995 69.305 197.040 ;
        RECT 71.300 196.995 71.620 197.055 ;
        RECT 69.015 196.855 71.620 196.995 ;
        RECT 69.015 196.810 69.305 196.855 ;
        RECT 71.300 196.795 71.620 196.855 ;
        RECT 76.360 196.995 76.680 197.055 ;
        RECT 80.500 196.995 80.820 197.055 ;
        RECT 76.360 196.855 80.820 196.995 ;
        RECT 76.360 196.795 76.680 196.855 ;
        RECT 80.500 196.795 80.820 196.855 ;
        RECT 65.340 196.605 65.630 196.700 ;
        RECT 64.490 196.470 65.630 196.605 ;
        RECT 64.490 196.465 65.550 196.470 ;
        RECT 66.240 196.455 66.560 196.715 ;
        RECT 66.715 196.655 67.005 196.700 ;
        RECT 68.080 196.655 68.400 196.715 ;
        RECT 66.715 196.515 68.400 196.655 ;
        RECT 66.715 196.470 67.005 196.515 ;
        RECT 68.080 196.455 68.400 196.515 ;
        RECT 69.460 196.455 69.780 196.715 ;
        RECT 65.780 196.315 66.100 196.375 ;
        RECT 69.000 196.315 69.320 196.375 ;
        RECT 73.555 196.360 73.845 196.675 ;
        RECT 74.635 196.655 74.925 196.700 ;
        RECT 78.215 196.655 78.505 196.700 ;
        RECT 80.050 196.655 80.340 196.700 ;
        RECT 74.635 196.515 80.340 196.655 ;
        RECT 74.635 196.470 74.925 196.515 ;
        RECT 78.215 196.470 78.505 196.515 ;
        RECT 80.050 196.470 80.340 196.515 ;
        RECT 60.720 196.175 69.320 196.315 ;
        RECT 60.720 196.115 61.040 196.175 ;
        RECT 65.780 196.115 66.100 196.175 ;
        RECT 69.000 196.115 69.320 196.175 ;
        RECT 73.255 196.315 73.845 196.360 ;
        RECT 74.060 196.315 74.380 196.375 ;
        RECT 76.495 196.315 77.145 196.360 ;
        RECT 73.255 196.175 77.145 196.315 ;
        RECT 73.255 196.130 73.545 196.175 ;
        RECT 74.060 196.115 74.380 196.175 ;
        RECT 76.495 196.130 77.145 196.175 ;
        RECT 79.120 196.115 79.440 196.375 ;
        RECT 58.420 195.775 58.740 196.035 ;
        RECT 65.320 195.975 65.640 196.035 ;
        RECT 67.620 195.975 67.940 196.035 ;
        RECT 65.320 195.835 67.940 195.975 ;
        RECT 65.320 195.775 65.640 195.835 ;
        RECT 67.620 195.775 67.940 195.835 ;
        RECT 71.760 195.775 72.080 196.035 ;
        RECT 10.510 195.155 115.850 195.635 ;
        RECT 54.740 194.755 55.060 195.015 ;
        RECT 59.355 194.955 59.645 195.000 ;
        RECT 61.180 194.955 61.500 195.015 ;
        RECT 59.355 194.815 61.500 194.955 ;
        RECT 59.355 194.770 59.645 194.815 ;
        RECT 61.180 194.755 61.500 194.815 ;
        RECT 63.940 194.755 64.260 195.015 ;
        RECT 67.620 194.955 67.940 195.015 ;
        RECT 72.315 194.955 72.605 195.000 ;
        RECT 67.620 194.815 72.605 194.955 ;
        RECT 67.620 194.755 67.940 194.815 ;
        RECT 72.315 194.770 72.605 194.815 ;
        RECT 73.155 194.955 73.445 195.000 ;
        RECT 73.600 194.955 73.920 195.015 ;
        RECT 73.155 194.815 73.920 194.955 ;
        RECT 73.155 194.770 73.445 194.815 ;
        RECT 73.600 194.755 73.920 194.815 ;
        RECT 74.060 194.955 74.380 195.015 ;
        RECT 74.535 194.955 74.825 195.000 ;
        RECT 74.060 194.815 74.825 194.955 ;
        RECT 74.060 194.755 74.380 194.815 ;
        RECT 74.535 194.770 74.825 194.815 ;
        RECT 75.915 194.955 76.205 195.000 ;
        RECT 79.120 194.955 79.440 195.015 ;
        RECT 75.915 194.815 79.440 194.955 ;
        RECT 75.915 194.770 76.205 194.815 ;
        RECT 79.120 194.755 79.440 194.815 ;
        RECT 65.210 194.615 65.500 194.660 ;
        RECT 67.160 194.615 67.480 194.675 ;
        RECT 55.290 194.475 64.170 194.615 ;
        RECT 42.320 194.075 42.640 194.335 ;
        RECT 55.290 194.320 55.430 194.475 ;
        RECT 59.430 194.335 59.570 194.475 ;
        RECT 64.030 194.335 64.170 194.475 ;
        RECT 65.210 194.475 67.480 194.615 ;
        RECT 65.210 194.430 65.500 194.475 ;
        RECT 67.160 194.415 67.480 194.475 ;
        RECT 69.000 194.415 69.320 194.675 ;
        RECT 71.300 194.415 71.620 194.675 ;
        RECT 89.240 194.615 89.560 194.675 ;
        RECT 91.075 194.615 91.725 194.660 ;
        RECT 94.675 194.615 94.965 194.660 ;
        RECT 89.240 194.475 94.965 194.615 ;
        RECT 89.240 194.415 89.560 194.475 ;
        RECT 91.075 194.430 91.725 194.475 ;
        RECT 94.375 194.430 94.965 194.475 ;
        RECT 55.215 194.090 55.505 194.320 ;
        RECT 59.340 194.075 59.660 194.335 ;
        RECT 60.720 194.275 61.040 194.335 ;
        RECT 61.195 194.275 61.485 194.320 ;
        RECT 60.720 194.135 61.485 194.275 ;
        RECT 60.720 194.075 61.040 194.135 ;
        RECT 61.195 194.090 61.485 194.135 ;
        RECT 61.640 194.275 61.960 194.335 ;
        RECT 62.575 194.275 62.865 194.320 ;
        RECT 63.480 194.275 63.800 194.335 ;
        RECT 61.640 194.135 63.800 194.275 ;
        RECT 61.640 194.075 61.960 194.135 ;
        RECT 62.575 194.090 62.865 194.135 ;
        RECT 63.480 194.075 63.800 194.135 ;
        RECT 63.940 194.075 64.260 194.335 ;
        RECT 64.400 194.275 64.720 194.335 ;
        RECT 66.255 194.275 66.545 194.320 ;
        RECT 64.400 194.135 66.545 194.275 ;
        RECT 64.400 194.075 64.720 194.135 ;
        RECT 66.255 194.090 66.545 194.135 ;
        RECT 56.595 193.935 56.885 193.980 ;
        RECT 58.420 193.935 58.740 193.995 ;
        RECT 56.595 193.795 59.340 193.935 ;
        RECT 56.595 193.750 56.885 193.795 ;
        RECT 58.420 193.735 58.740 193.795 ;
        RECT 42.780 193.055 43.100 193.315 ;
        RECT 59.200 193.255 59.340 193.795 ;
        RECT 65.795 193.750 66.085 193.980 ;
        RECT 62.560 193.595 62.880 193.655 ;
        RECT 64.415 193.595 64.705 193.640 ;
        RECT 62.560 193.455 64.705 193.595 ;
        RECT 65.870 193.595 66.010 193.750 ;
        RECT 67.620 193.735 67.940 193.995 ;
        RECT 69.090 193.935 69.230 194.415 ;
        RECT 69.920 194.075 70.240 194.335 ;
        RECT 74.060 194.075 74.380 194.335 ;
        RECT 75.455 194.090 75.745 194.320 ;
        RECT 80.500 194.275 80.820 194.335 ;
        RECT 86.480 194.275 86.800 194.335 ;
        RECT 87.415 194.275 87.705 194.320 ;
        RECT 80.500 194.135 87.705 194.275 ;
        RECT 70.840 193.935 71.160 193.995 ;
        RECT 75.530 193.935 75.670 194.090 ;
        RECT 80.500 194.075 80.820 194.135 ;
        RECT 86.480 194.075 86.800 194.135 ;
        RECT 87.415 194.090 87.705 194.135 ;
        RECT 87.880 194.275 88.170 194.320 ;
        RECT 89.715 194.275 90.005 194.320 ;
        RECT 93.295 194.275 93.585 194.320 ;
        RECT 87.880 194.135 93.585 194.275 ;
        RECT 87.880 194.090 88.170 194.135 ;
        RECT 89.715 194.090 90.005 194.135 ;
        RECT 93.295 194.090 93.585 194.135 ;
        RECT 94.375 194.115 94.665 194.430 ;
        RECT 102.135 194.275 102.425 194.320 ;
        RECT 102.580 194.275 102.900 194.335 ;
        RECT 102.135 194.135 102.900 194.275 ;
        RECT 102.135 194.090 102.425 194.135 ;
        RECT 102.580 194.075 102.900 194.135 ;
        RECT 103.500 194.275 103.820 194.335 ;
        RECT 103.975 194.275 104.265 194.320 ;
        RECT 103.500 194.135 104.265 194.275 ;
        RECT 103.500 194.075 103.820 194.135 ;
        RECT 103.975 194.090 104.265 194.135 ;
        RECT 69.090 193.795 75.670 193.935 ;
        RECT 88.795 193.935 89.085 193.980 ;
        RECT 92.460 193.935 92.780 193.995 ;
        RECT 88.795 193.795 92.780 193.935 ;
        RECT 70.840 193.735 71.160 193.795 ;
        RECT 88.795 193.750 89.085 193.795 ;
        RECT 92.460 193.735 92.780 193.795 ;
        RECT 66.240 193.595 66.560 193.655 ;
        RECT 65.870 193.455 66.560 193.595 ;
        RECT 62.560 193.395 62.880 193.455 ;
        RECT 64.415 193.410 64.705 193.455 ;
        RECT 66.240 193.395 66.560 193.455 ;
        RECT 88.285 193.595 88.575 193.640 ;
        RECT 90.175 193.595 90.465 193.640 ;
        RECT 93.295 193.595 93.585 193.640 ;
        RECT 88.285 193.455 93.585 193.595 ;
        RECT 88.285 193.410 88.575 193.455 ;
        RECT 90.175 193.410 90.465 193.455 ;
        RECT 93.295 193.410 93.585 193.455 ;
        RECT 63.020 193.255 63.340 193.315 ;
        RECT 59.200 193.115 63.340 193.255 ;
        RECT 63.020 193.055 63.340 193.115 ;
        RECT 70.855 193.255 71.145 193.300 ;
        RECT 72.235 193.255 72.525 193.300 ;
        RECT 70.855 193.115 72.525 193.255 ;
        RECT 70.855 193.070 71.145 193.115 ;
        RECT 72.235 193.070 72.525 193.115 ;
        RECT 96.155 193.255 96.445 193.300 ;
        RECT 97.520 193.255 97.840 193.315 ;
        RECT 96.155 193.115 97.840 193.255 ;
        RECT 96.155 193.070 96.445 193.115 ;
        RECT 97.520 193.055 97.840 193.115 ;
        RECT 101.675 193.255 101.965 193.300 ;
        RECT 102.120 193.255 102.440 193.315 ;
        RECT 101.675 193.115 102.440 193.255 ;
        RECT 101.675 193.070 101.965 193.115 ;
        RECT 102.120 193.055 102.440 193.115 ;
        RECT 104.895 193.255 105.185 193.300 ;
        RECT 105.800 193.255 106.120 193.315 ;
        RECT 104.895 193.115 106.120 193.255 ;
        RECT 104.895 193.070 105.185 193.115 ;
        RECT 105.800 193.055 106.120 193.115 ;
        RECT 10.510 192.435 115.850 192.915 ;
        RECT 60.260 192.035 60.580 192.295 ;
        RECT 63.940 192.235 64.260 192.295 ;
        RECT 74.060 192.235 74.380 192.295 ;
        RECT 63.940 192.095 74.380 192.235 ;
        RECT 63.940 192.035 64.260 192.095 ;
        RECT 74.060 192.035 74.380 192.095 ;
        RECT 88.795 192.235 89.085 192.280 ;
        RECT 89.240 192.235 89.560 192.295 ;
        RECT 102.580 192.235 102.900 192.295 ;
        RECT 88.795 192.095 89.560 192.235 ;
        RECT 88.795 192.050 89.085 192.095 ;
        RECT 89.240 192.035 89.560 192.095 ;
        RECT 89.790 192.095 102.900 192.235 ;
        RECT 27.110 191.895 27.400 191.940 ;
        RECT 29.890 191.895 30.180 191.940 ;
        RECT 31.750 191.895 32.040 191.940 ;
        RECT 69.015 191.895 69.305 191.940 ;
        RECT 69.460 191.895 69.780 191.955 ;
        RECT 27.110 191.755 32.040 191.895 ;
        RECT 27.110 191.710 27.400 191.755 ;
        RECT 29.890 191.710 30.180 191.755 ;
        RECT 31.750 191.710 32.040 191.755 ;
        RECT 60.350 191.755 69.780 191.895 ;
        RECT 29.440 191.555 29.760 191.615 ;
        RECT 30.375 191.555 30.665 191.600 ;
        RECT 29.440 191.415 30.665 191.555 ;
        RECT 29.440 191.355 29.760 191.415 ;
        RECT 30.375 191.370 30.665 191.415 ;
        RECT 27.110 191.215 27.400 191.260 ;
        RECT 29.900 191.215 30.220 191.275 ;
        RECT 32.215 191.215 32.505 191.260 ;
        RECT 27.110 191.075 29.645 191.215 ;
        RECT 27.110 191.030 27.400 191.075 ;
        RECT 24.380 190.875 24.700 190.935 ;
        RECT 29.430 190.920 29.645 191.075 ;
        RECT 29.900 191.075 32.505 191.215 ;
        RECT 29.900 191.015 30.220 191.075 ;
        RECT 32.215 191.030 32.505 191.075 ;
        RECT 40.495 191.030 40.785 191.260 ;
        RECT 25.250 190.875 25.540 190.920 ;
        RECT 28.510 190.875 28.800 190.920 ;
        RECT 24.380 190.735 28.800 190.875 ;
        RECT 24.380 190.675 24.700 190.735 ;
        RECT 25.250 190.690 25.540 190.735 ;
        RECT 28.510 190.690 28.800 190.735 ;
        RECT 29.430 190.875 29.720 190.920 ;
        RECT 31.290 190.875 31.580 190.920 ;
        RECT 29.430 190.735 31.580 190.875 ;
        RECT 40.570 190.875 40.710 191.030 ;
        RECT 40.940 191.015 41.260 191.275 ;
        RECT 45.555 191.215 45.845 191.260 ;
        RECT 46.000 191.215 46.320 191.275 ;
        RECT 45.555 191.075 46.320 191.215 ;
        RECT 45.555 191.030 45.845 191.075 ;
        RECT 46.000 191.015 46.320 191.075 ;
        RECT 58.880 191.015 59.200 191.275 ;
        RECT 60.350 190.935 60.490 191.755 ;
        RECT 69.015 191.710 69.305 191.755 ;
        RECT 69.460 191.695 69.780 191.755 ;
        RECT 66.715 191.555 67.005 191.600 ;
        RECT 67.160 191.555 67.480 191.615 ;
        RECT 66.715 191.415 67.480 191.555 ;
        RECT 66.715 191.370 67.005 191.415 ;
        RECT 67.160 191.355 67.480 191.415 ;
        RECT 71.760 191.555 72.080 191.615 ;
        RECT 72.695 191.555 72.985 191.600 ;
        RECT 71.760 191.415 72.985 191.555 ;
        RECT 71.760 191.355 72.080 191.415 ;
        RECT 72.695 191.370 72.985 191.415 ;
        RECT 74.060 191.555 74.380 191.615 ;
        RECT 78.200 191.555 78.520 191.615 ;
        RECT 74.060 191.415 88.550 191.555 ;
        RECT 74.060 191.355 74.380 191.415 ;
        RECT 78.200 191.355 78.520 191.415 ;
        RECT 60.735 191.215 61.025 191.260 ;
        RECT 61.640 191.215 61.960 191.275 ;
        RECT 60.735 191.075 61.960 191.215 ;
        RECT 60.735 191.030 61.025 191.075 ;
        RECT 61.640 191.015 61.960 191.075 ;
        RECT 66.240 191.215 66.560 191.275 ;
        RECT 71.850 191.215 71.990 191.355 ;
        RECT 66.240 191.075 71.990 191.215 ;
        RECT 80.515 191.215 80.805 191.260 ;
        RECT 81.420 191.215 81.740 191.275 ;
        RECT 88.410 191.260 88.550 191.415 ;
        RECT 80.515 191.075 81.740 191.215 ;
        RECT 66.240 191.015 66.560 191.075 ;
        RECT 80.515 191.030 80.805 191.075 ;
        RECT 81.420 191.015 81.740 191.075 ;
        RECT 81.895 191.030 82.185 191.260 ;
        RECT 88.335 191.215 88.625 191.260 ;
        RECT 89.790 191.215 89.930 192.095 ;
        RECT 102.580 192.035 102.900 192.095 ;
        RECT 101.315 191.895 101.605 191.940 ;
        RECT 104.435 191.895 104.725 191.940 ;
        RECT 106.325 191.895 106.615 191.940 ;
        RECT 101.315 191.755 106.615 191.895 ;
        RECT 101.315 191.710 101.605 191.755 ;
        RECT 104.435 191.710 104.725 191.755 ;
        RECT 106.325 191.710 106.615 191.755 ;
        RECT 95.235 191.555 95.525 191.600 ;
        RECT 98.440 191.555 98.760 191.615 ;
        RECT 95.235 191.415 98.760 191.555 ;
        RECT 95.235 191.370 95.525 191.415 ;
        RECT 98.440 191.355 98.760 191.415 ;
        RECT 105.800 191.355 106.120 191.615 ;
        RECT 88.335 191.075 89.930 191.215 ;
        RECT 93.395 191.215 93.685 191.260 ;
        RECT 97.520 191.215 97.840 191.275 ;
        RECT 93.395 191.075 97.840 191.215 ;
        RECT 88.335 191.030 88.625 191.075 ;
        RECT 93.395 191.030 93.685 191.075 ;
        RECT 42.320 190.875 42.640 190.935 ;
        RECT 44.620 190.875 44.940 190.935 ;
        RECT 40.570 190.735 44.940 190.875 ;
        RECT 29.430 190.690 29.720 190.735 ;
        RECT 31.290 190.690 31.580 190.735 ;
        RECT 42.320 190.675 42.640 190.735 ;
        RECT 44.620 190.675 44.940 190.735 ;
        RECT 59.355 190.875 59.645 190.920 ;
        RECT 60.260 190.875 60.580 190.935 ;
        RECT 59.355 190.735 60.580 190.875 ;
        RECT 59.355 190.690 59.645 190.735 ;
        RECT 60.260 190.675 60.580 190.735 ;
        RECT 67.620 190.875 67.940 190.935 ;
        RECT 69.000 190.875 69.320 190.935 ;
        RECT 67.620 190.735 69.320 190.875 ;
        RECT 67.620 190.675 67.940 190.735 ;
        RECT 69.000 190.675 69.320 190.735 ;
        RECT 76.360 190.875 76.680 190.935 ;
        RECT 81.970 190.875 82.110 191.030 ;
        RECT 97.520 191.015 97.840 191.075 ;
        RECT 100.235 190.920 100.525 191.235 ;
        RECT 101.315 191.215 101.605 191.260 ;
        RECT 104.895 191.215 105.185 191.260 ;
        RECT 106.730 191.215 107.020 191.260 ;
        RECT 101.315 191.075 107.020 191.215 ;
        RECT 101.315 191.030 101.605 191.075 ;
        RECT 104.895 191.030 105.185 191.075 ;
        RECT 106.730 191.030 107.020 191.075 ;
        RECT 107.195 191.215 107.485 191.260 ;
        RECT 107.640 191.215 107.960 191.275 ;
        RECT 107.195 191.075 107.960 191.215 ;
        RECT 107.195 191.030 107.485 191.075 ;
        RECT 107.640 191.015 107.960 191.075 ;
        RECT 109.495 191.030 109.785 191.260 ;
        RECT 76.360 190.735 82.110 190.875 ;
        RECT 99.935 190.875 100.525 190.920 ;
        RECT 102.120 190.875 102.440 190.935 ;
        RECT 103.175 190.875 103.825 190.920 ;
        RECT 99.935 190.735 103.825 190.875 ;
        RECT 76.360 190.675 76.680 190.735 ;
        RECT 99.935 190.690 100.225 190.735 ;
        RECT 102.120 190.675 102.440 190.735 ;
        RECT 103.175 190.690 103.825 190.735 ;
        RECT 106.260 190.875 106.580 190.935 ;
        RECT 109.570 190.875 109.710 191.030 ;
        RECT 106.260 190.735 109.710 190.875 ;
        RECT 106.260 190.675 106.580 190.735 ;
        RECT 23.245 190.535 23.535 190.580 ;
        RECT 28.060 190.535 28.380 190.595 ;
        RECT 23.245 190.395 28.380 190.535 ;
        RECT 23.245 190.350 23.535 190.395 ;
        RECT 28.060 190.335 28.380 190.395 ;
        RECT 40.020 190.335 40.340 190.595 ;
        RECT 43.700 190.535 44.020 190.595 ;
        RECT 44.175 190.535 44.465 190.580 ;
        RECT 43.700 190.395 44.465 190.535 ;
        RECT 43.700 190.335 44.020 190.395 ;
        RECT 44.175 190.350 44.465 190.395 ;
        RECT 46.460 190.335 46.780 190.595 ;
        RECT 59.815 190.535 60.105 190.580 ;
        RECT 60.720 190.535 61.040 190.595 ;
        RECT 59.815 190.395 61.040 190.535 ;
        RECT 59.815 190.350 60.105 190.395 ;
        RECT 60.720 190.335 61.040 190.395 ;
        RECT 61.180 190.535 61.500 190.595 ;
        RECT 65.335 190.535 65.625 190.580 ;
        RECT 61.180 190.395 65.625 190.535 ;
        RECT 61.180 190.335 61.500 190.395 ;
        RECT 65.335 190.350 65.625 190.395 ;
        RECT 69.935 190.535 70.225 190.580 ;
        RECT 70.380 190.535 70.700 190.595 ;
        RECT 69.935 190.395 70.700 190.535 ;
        RECT 69.935 190.350 70.225 190.395 ;
        RECT 70.380 190.335 70.700 190.395 ;
        RECT 80.960 190.335 81.280 190.595 ;
        RECT 82.815 190.535 83.105 190.580 ;
        RECT 84.640 190.535 84.960 190.595 ;
        RECT 82.815 190.395 84.960 190.535 ;
        RECT 82.815 190.350 83.105 190.395 ;
        RECT 84.640 190.335 84.960 190.395 ;
        RECT 90.175 190.535 90.465 190.580 ;
        RECT 90.620 190.535 90.940 190.595 ;
        RECT 90.175 190.395 90.940 190.535 ;
        RECT 90.175 190.350 90.465 190.395 ;
        RECT 90.620 190.335 90.940 190.395 ;
        RECT 97.995 190.535 98.285 190.580 ;
        RECT 99.360 190.535 99.680 190.595 ;
        RECT 97.995 190.395 99.680 190.535 ;
        RECT 97.995 190.350 98.285 190.395 ;
        RECT 99.360 190.335 99.680 190.395 ;
        RECT 110.415 190.535 110.705 190.580 ;
        RECT 112.240 190.535 112.560 190.595 ;
        RECT 110.415 190.395 112.560 190.535 ;
        RECT 110.415 190.350 110.705 190.395 ;
        RECT 112.240 190.335 112.560 190.395 ;
        RECT 10.510 189.715 115.850 190.195 ;
        RECT 24.380 189.315 24.700 189.575 ;
        RECT 49.695 189.515 49.985 189.560 ;
        RECT 47.930 189.375 49.985 189.515 ;
        RECT 34.040 189.175 34.360 189.235 ;
        RECT 38.655 189.175 38.945 189.220 ;
        RECT 24.010 189.035 31.510 189.175 ;
        RECT 24.010 188.895 24.150 189.035 ;
        RECT 23.920 188.635 24.240 188.895 ;
        RECT 28.520 188.635 28.840 188.895 ;
        RECT 31.370 188.880 31.510 189.035 ;
        RECT 34.040 189.035 38.945 189.175 ;
        RECT 34.040 188.975 34.360 189.035 ;
        RECT 38.655 188.990 38.945 189.035 ;
        RECT 41.975 189.175 42.265 189.220 ;
        RECT 42.780 189.175 43.100 189.235 ;
        RECT 47.930 189.220 48.070 189.375 ;
        RECT 49.695 189.330 49.985 189.375 ;
        RECT 70.840 189.315 71.160 189.575 ;
        RECT 76.360 189.315 76.680 189.575 ;
        RECT 92.460 189.315 92.780 189.575 ;
        RECT 102.135 189.515 102.425 189.560 ;
        RECT 103.500 189.515 103.820 189.575 ;
        RECT 102.135 189.375 103.820 189.515 ;
        RECT 102.135 189.330 102.425 189.375 ;
        RECT 103.500 189.315 103.820 189.375 ;
        RECT 45.215 189.175 45.865 189.220 ;
        RECT 41.975 189.035 45.865 189.175 ;
        RECT 41.975 188.990 42.565 189.035 ;
        RECT 31.295 188.650 31.585 188.880 ;
        RECT 38.180 188.635 38.500 188.895 ;
        RECT 42.275 188.675 42.565 188.990 ;
        RECT 42.780 188.975 43.100 189.035 ;
        RECT 45.215 188.990 45.865 189.035 ;
        RECT 47.855 188.990 48.145 189.220 ;
        RECT 67.160 188.975 67.480 189.235 ;
        RECT 70.380 188.975 70.700 189.235 ;
        RECT 73.600 189.175 73.920 189.235 ;
        RECT 74.535 189.175 74.825 189.220 ;
        RECT 73.600 189.035 74.825 189.175 ;
        RECT 73.600 188.975 73.920 189.035 ;
        RECT 74.535 188.990 74.825 189.035 ;
        RECT 79.530 189.175 79.820 189.220 ;
        RECT 80.960 189.175 81.280 189.235 ;
        RECT 82.790 189.175 83.080 189.220 ;
        RECT 79.530 189.035 83.080 189.175 ;
        RECT 79.530 188.990 79.820 189.035 ;
        RECT 80.960 188.975 81.280 189.035 ;
        RECT 82.790 188.990 83.080 189.035 ;
        RECT 83.710 189.175 84.000 189.220 ;
        RECT 85.570 189.175 85.860 189.220 ;
        RECT 83.710 189.035 85.860 189.175 ;
        RECT 83.710 188.990 84.000 189.035 ;
        RECT 85.570 188.990 85.860 189.035 ;
        RECT 89.715 189.175 90.005 189.220 ;
        RECT 90.620 189.175 90.940 189.235 ;
        RECT 100.295 189.175 100.585 189.220 ;
        RECT 89.715 189.035 100.585 189.175 ;
        RECT 89.715 188.990 90.005 189.035 ;
        RECT 43.355 188.835 43.645 188.880 ;
        RECT 46.935 188.835 47.225 188.880 ;
        RECT 48.770 188.835 49.060 188.880 ;
        RECT 43.355 188.695 49.060 188.835 ;
        RECT 43.355 188.650 43.645 188.695 ;
        RECT 46.935 188.650 47.225 188.695 ;
        RECT 48.770 188.650 49.060 188.695 ;
        RECT 49.680 188.835 50.000 188.895 ;
        RECT 50.615 188.835 50.905 188.880 ;
        RECT 49.680 188.695 50.905 188.835 ;
        RECT 49.680 188.635 50.000 188.695 ;
        RECT 50.615 188.650 50.905 188.695 ;
        RECT 54.740 188.635 55.060 188.895 ;
        RECT 78.200 188.835 78.520 188.895 ;
        RECT 73.690 188.695 78.520 188.835 ;
        RECT 26.680 188.495 27.000 188.555 ;
        RECT 27.155 188.495 27.445 188.540 ;
        RECT 26.680 188.355 27.445 188.495 ;
        RECT 26.680 188.295 27.000 188.355 ;
        RECT 27.155 188.310 27.445 188.355 ;
        RECT 28.060 188.295 28.380 188.555 ;
        RECT 35.895 188.310 36.185 188.540 ;
        RECT 28.150 188.155 28.290 188.295 ;
        RECT 31.280 188.155 31.600 188.215 ;
        RECT 28.150 188.015 31.600 188.155 ;
        RECT 35.970 188.155 36.110 188.310 ;
        RECT 39.100 188.295 39.420 188.555 ;
        RECT 49.235 188.495 49.525 188.540 ;
        RECT 52.900 188.495 53.220 188.555 ;
        RECT 58.420 188.495 58.740 188.555 ;
        RECT 49.235 188.355 58.740 188.495 ;
        RECT 49.235 188.310 49.525 188.355 ;
        RECT 52.900 188.295 53.220 188.355 ;
        RECT 58.420 188.295 58.740 188.355 ;
        RECT 73.140 188.495 73.460 188.555 ;
        RECT 73.690 188.540 73.830 188.695 ;
        RECT 78.200 188.635 78.520 188.695 ;
        RECT 81.390 188.835 81.680 188.880 ;
        RECT 83.710 188.835 83.925 188.990 ;
        RECT 90.620 188.975 90.940 189.035 ;
        RECT 100.295 188.990 100.585 189.035 ;
        RECT 103.975 189.175 104.265 189.220 ;
        RECT 106.375 189.175 106.665 189.220 ;
        RECT 109.615 189.175 110.265 189.220 ;
        RECT 103.975 189.035 110.265 189.175 ;
        RECT 103.975 188.990 104.265 189.035 ;
        RECT 106.375 188.990 106.965 189.035 ;
        RECT 109.615 188.990 110.265 189.035 ;
        RECT 81.390 188.695 83.925 188.835 ;
        RECT 81.390 188.650 81.680 188.695 ;
        RECT 84.640 188.635 84.960 188.895 ;
        RECT 86.480 188.635 86.800 188.895 ;
        RECT 90.175 188.835 90.465 188.880 ;
        RECT 93.395 188.835 93.685 188.880 ;
        RECT 87.030 188.695 90.465 188.835 ;
        RECT 73.615 188.495 73.905 188.540 ;
        RECT 73.140 188.355 73.905 188.495 ;
        RECT 73.140 188.295 73.460 188.355 ;
        RECT 73.615 188.310 73.905 188.355 ;
        RECT 74.075 188.495 74.365 188.540 ;
        RECT 87.030 188.495 87.170 188.695 ;
        RECT 90.175 188.650 90.465 188.695 ;
        RECT 92.090 188.695 93.685 188.835 ;
        RECT 74.075 188.355 87.170 188.495 ;
        RECT 74.075 188.310 74.365 188.355 ;
        RECT 36.355 188.155 36.645 188.200 ;
        RECT 35.970 188.015 36.645 188.155 ;
        RECT 31.280 187.955 31.600 188.015 ;
        RECT 36.355 187.970 36.645 188.015 ;
        RECT 43.355 188.155 43.645 188.200 ;
        RECT 46.475 188.155 46.765 188.200 ;
        RECT 48.365 188.155 48.655 188.200 ;
        RECT 43.355 188.015 48.655 188.155 ;
        RECT 43.355 187.970 43.645 188.015 ;
        RECT 46.475 187.970 46.765 188.015 ;
        RECT 48.365 187.970 48.655 188.015 ;
        RECT 75.990 187.875 76.130 188.355 ;
        RECT 89.255 188.310 89.545 188.540 ;
        RECT 81.390 188.155 81.680 188.200 ;
        RECT 84.170 188.155 84.460 188.200 ;
        RECT 86.030 188.155 86.320 188.200 ;
        RECT 81.390 188.015 86.320 188.155 ;
        RECT 81.390 187.970 81.680 188.015 ;
        RECT 84.170 187.970 84.460 188.015 ;
        RECT 86.030 187.970 86.320 188.015 ;
        RECT 30.360 187.615 30.680 187.875 ;
        RECT 30.820 187.815 31.140 187.875 ;
        RECT 31.755 187.815 32.045 187.860 ;
        RECT 30.820 187.675 32.045 187.815 ;
        RECT 30.820 187.615 31.140 187.675 ;
        RECT 31.755 187.630 32.045 187.675 ;
        RECT 32.660 187.615 32.980 187.875 ;
        RECT 40.480 187.615 40.800 187.875 ;
        RECT 55.675 187.815 55.965 187.860 ;
        RECT 57.040 187.815 57.360 187.875 ;
        RECT 55.675 187.675 57.360 187.815 ;
        RECT 55.675 187.630 55.965 187.675 ;
        RECT 57.040 187.615 57.360 187.675 ;
        RECT 67.160 187.815 67.480 187.875 ;
        RECT 67.635 187.815 67.925 187.860 ;
        RECT 69.920 187.815 70.240 187.875 ;
        RECT 67.160 187.675 70.240 187.815 ;
        RECT 67.160 187.615 67.480 187.675 ;
        RECT 67.635 187.630 67.925 187.675 ;
        RECT 69.920 187.615 70.240 187.675 ;
        RECT 75.900 187.815 76.220 187.875 ;
        RECT 77.525 187.815 77.815 187.860 ;
        RECT 75.900 187.675 77.815 187.815 ;
        RECT 75.900 187.615 76.220 187.675 ;
        RECT 77.525 187.630 77.815 187.675 ;
        RECT 78.200 187.815 78.520 187.875 ;
        RECT 89.330 187.815 89.470 188.310 ;
        RECT 92.090 188.200 92.230 188.695 ;
        RECT 93.395 188.650 93.685 188.695 ;
        RECT 95.235 188.835 95.525 188.880 ;
        RECT 100.740 188.835 101.060 188.895 ;
        RECT 95.235 188.695 101.060 188.835 ;
        RECT 95.235 188.650 95.525 188.695 ;
        RECT 100.740 188.635 101.060 188.695 ;
        RECT 102.580 188.835 102.900 188.895 ;
        RECT 103.515 188.835 103.805 188.880 ;
        RECT 104.880 188.835 105.200 188.895 ;
        RECT 102.580 188.695 105.200 188.835 ;
        RECT 102.580 188.635 102.900 188.695 ;
        RECT 103.515 188.650 103.805 188.695 ;
        RECT 104.880 188.635 105.200 188.695 ;
        RECT 106.675 188.675 106.965 188.990 ;
        RECT 112.240 188.975 112.560 189.235 ;
        RECT 107.755 188.835 108.045 188.880 ;
        RECT 111.335 188.835 111.625 188.880 ;
        RECT 113.170 188.835 113.460 188.880 ;
        RECT 107.755 188.695 113.460 188.835 ;
        RECT 107.755 188.650 108.045 188.695 ;
        RECT 111.335 188.650 111.625 188.695 ;
        RECT 113.170 188.650 113.460 188.695 ;
        RECT 99.375 188.310 99.665 188.540 ;
        RECT 92.015 187.970 92.305 188.200 ;
        RECT 99.450 188.155 99.590 188.310 ;
        RECT 99.820 188.295 100.140 188.555 ;
        RECT 113.635 188.495 113.925 188.540 ;
        RECT 114.080 188.495 114.400 188.555 ;
        RECT 113.635 188.355 114.400 188.495 ;
        RECT 113.635 188.310 113.925 188.355 ;
        RECT 114.080 188.295 114.400 188.355 ;
        RECT 104.420 188.155 104.740 188.215 ;
        RECT 99.450 188.015 104.740 188.155 ;
        RECT 104.420 187.955 104.740 188.015 ;
        RECT 107.755 188.155 108.045 188.200 ;
        RECT 110.875 188.155 111.165 188.200 ;
        RECT 112.765 188.155 113.055 188.200 ;
        RECT 107.755 188.015 113.055 188.155 ;
        RECT 107.755 187.970 108.045 188.015 ;
        RECT 110.875 187.970 111.165 188.015 ;
        RECT 112.765 187.970 113.055 188.015 ;
        RECT 92.460 187.815 92.780 187.875 ;
        RECT 78.200 187.675 92.780 187.815 ;
        RECT 78.200 187.615 78.520 187.675 ;
        RECT 92.460 187.615 92.780 187.675 ;
        RECT 97.995 187.815 98.285 187.860 ;
        RECT 100.280 187.815 100.600 187.875 ;
        RECT 97.995 187.675 100.600 187.815 ;
        RECT 97.995 187.630 98.285 187.675 ;
        RECT 100.280 187.615 100.600 187.675 ;
        RECT 104.895 187.815 105.185 187.860 ;
        RECT 109.480 187.815 109.800 187.875 ;
        RECT 104.895 187.675 109.800 187.815 ;
        RECT 104.895 187.630 105.185 187.675 ;
        RECT 109.480 187.615 109.800 187.675 ;
        RECT 10.510 186.995 115.850 187.475 ;
        RECT 28.995 186.795 29.285 186.840 ;
        RECT 34.040 186.795 34.360 186.855 ;
        RECT 28.995 186.655 34.360 186.795 ;
        RECT 28.995 186.610 29.285 186.655 ;
        RECT 34.040 186.595 34.360 186.655 ;
        RECT 37.810 186.655 48.070 186.795 ;
        RECT 22.655 186.455 22.945 186.500 ;
        RECT 25.775 186.455 26.065 186.500 ;
        RECT 27.665 186.455 27.955 186.500 ;
        RECT 22.655 186.315 27.955 186.455 ;
        RECT 22.655 186.270 22.945 186.315 ;
        RECT 25.775 186.270 26.065 186.315 ;
        RECT 27.665 186.270 27.955 186.315 ;
        RECT 31.855 186.455 32.145 186.500 ;
        RECT 34.975 186.455 35.265 186.500 ;
        RECT 36.865 186.455 37.155 186.500 ;
        RECT 31.855 186.315 37.155 186.455 ;
        RECT 31.855 186.270 32.145 186.315 ;
        RECT 34.975 186.270 35.265 186.315 ;
        RECT 36.865 186.270 37.155 186.315 ;
        RECT 28.535 186.115 28.825 186.160 ;
        RECT 29.900 186.115 30.220 186.175 ;
        RECT 37.810 186.160 37.950 186.655 ;
        RECT 41.975 186.455 42.265 186.500 ;
        RECT 45.095 186.455 45.385 186.500 ;
        RECT 46.985 186.455 47.275 186.500 ;
        RECT 41.975 186.315 47.275 186.455 ;
        RECT 41.975 186.270 42.265 186.315 ;
        RECT 45.095 186.270 45.385 186.315 ;
        RECT 46.985 186.270 47.275 186.315 ;
        RECT 28.535 185.975 30.220 186.115 ;
        RECT 28.535 185.930 28.825 185.975 ;
        RECT 29.900 185.915 30.220 185.975 ;
        RECT 37.735 185.930 38.025 186.160 ;
        RECT 46.460 185.915 46.780 186.175 ;
        RECT 47.930 186.160 48.070 186.655 ;
        RECT 106.260 186.595 106.580 186.855 ;
        RECT 52.555 186.455 52.845 186.500 ;
        RECT 55.675 186.455 55.965 186.500 ;
        RECT 57.565 186.455 57.855 186.500 ;
        RECT 52.555 186.315 57.855 186.455 ;
        RECT 52.555 186.270 52.845 186.315 ;
        RECT 55.675 186.270 55.965 186.315 ;
        RECT 57.565 186.270 57.855 186.315 ;
        RECT 59.800 186.455 60.120 186.515 ;
        RECT 60.720 186.455 61.040 186.515 ;
        RECT 77.250 186.455 77.540 186.500 ;
        RECT 80.030 186.455 80.320 186.500 ;
        RECT 81.890 186.455 82.180 186.500 ;
        RECT 59.800 186.315 62.790 186.455 ;
        RECT 59.800 186.255 60.120 186.315 ;
        RECT 60.720 186.255 61.040 186.315 ;
        RECT 47.855 186.115 48.145 186.160 ;
        RECT 53.360 186.115 53.680 186.175 ;
        RECT 47.855 185.975 53.680 186.115 ;
        RECT 47.855 185.930 48.145 185.975 ;
        RECT 53.360 185.915 53.680 185.975 ;
        RECT 57.040 185.915 57.360 186.175 ;
        RECT 58.420 185.915 58.740 186.175 ;
        RECT 58.880 186.115 59.200 186.175 ;
        RECT 62.650 186.160 62.790 186.315 ;
        RECT 77.250 186.315 82.180 186.455 ;
        RECT 77.250 186.270 77.540 186.315 ;
        RECT 80.030 186.270 80.320 186.315 ;
        RECT 81.890 186.270 82.180 186.315 ;
        RECT 91.045 186.455 91.335 186.500 ;
        RECT 92.935 186.455 93.225 186.500 ;
        RECT 96.055 186.455 96.345 186.500 ;
        RECT 91.045 186.315 96.345 186.455 ;
        RECT 91.045 186.270 91.335 186.315 ;
        RECT 92.935 186.270 93.225 186.315 ;
        RECT 96.055 186.270 96.345 186.315 ;
        RECT 61.655 186.115 61.945 186.160 ;
        RECT 58.880 185.975 61.945 186.115 ;
        RECT 58.880 185.915 59.200 185.975 ;
        RECT 61.655 185.930 61.945 185.975 ;
        RECT 62.575 185.930 62.865 186.160 ;
        RECT 81.420 186.115 81.740 186.175 ;
        RECT 72.770 185.975 81.740 186.115 ;
        RECT 21.575 185.480 21.865 185.795 ;
        RECT 22.655 185.775 22.945 185.820 ;
        RECT 26.235 185.775 26.525 185.820 ;
        RECT 28.070 185.775 28.360 185.820 ;
        RECT 30.820 185.795 31.140 185.835 ;
        RECT 22.655 185.635 28.360 185.775 ;
        RECT 22.655 185.590 22.945 185.635 ;
        RECT 26.235 185.590 26.525 185.635 ;
        RECT 28.070 185.590 28.360 185.635 ;
        RECT 30.775 185.575 31.140 185.795 ;
        RECT 31.855 185.775 32.145 185.820 ;
        RECT 35.435 185.775 35.725 185.820 ;
        RECT 37.270 185.775 37.560 185.820 ;
        RECT 31.855 185.635 37.560 185.775 ;
        RECT 31.855 185.590 32.145 185.635 ;
        RECT 35.435 185.590 35.725 185.635 ;
        RECT 37.270 185.590 37.560 185.635 ;
        RECT 24.840 185.480 25.160 185.495 ;
        RECT 21.275 185.435 21.865 185.480 ;
        RECT 24.515 185.435 25.165 185.480 ;
        RECT 21.275 185.295 25.165 185.435 ;
        RECT 21.275 185.250 21.565 185.295 ;
        RECT 24.515 185.250 25.165 185.295 ;
        RECT 24.840 185.235 25.160 185.250 ;
        RECT 27.140 185.235 27.460 185.495 ;
        RECT 30.775 185.480 31.065 185.575 ;
        RECT 30.475 185.435 31.065 185.480 ;
        RECT 33.715 185.435 34.365 185.480 ;
        RECT 36.355 185.435 36.645 185.480 ;
        RECT 30.475 185.295 34.365 185.435 ;
        RECT 30.475 185.250 30.765 185.295 ;
        RECT 33.715 185.250 34.365 185.295 ;
        RECT 34.590 185.295 36.645 185.435 ;
        RECT 34.590 185.155 34.730 185.295 ;
        RECT 36.355 185.250 36.645 185.295 ;
        RECT 40.020 185.435 40.340 185.495 ;
        RECT 40.895 185.480 41.185 185.795 ;
        RECT 41.975 185.775 42.265 185.820 ;
        RECT 45.555 185.775 45.845 185.820 ;
        RECT 47.390 185.775 47.680 185.820 ;
        RECT 41.975 185.635 47.680 185.775 ;
        RECT 41.975 185.590 42.265 185.635 ;
        RECT 45.555 185.590 45.845 185.635 ;
        RECT 47.390 185.590 47.680 185.635 ;
        RECT 48.315 185.775 48.605 185.820 ;
        RECT 50.600 185.775 50.920 185.835 ;
        RECT 48.315 185.635 50.920 185.775 ;
        RECT 48.315 185.590 48.605 185.635 ;
        RECT 40.595 185.435 41.185 185.480 ;
        RECT 43.835 185.435 44.485 185.480 ;
        RECT 40.020 185.295 44.485 185.435 ;
        RECT 40.020 185.235 40.340 185.295 ;
        RECT 40.595 185.250 40.885 185.295 ;
        RECT 43.835 185.250 44.485 185.295 ;
        RECT 45.080 185.435 45.400 185.495 ;
        RECT 48.390 185.435 48.530 185.590 ;
        RECT 50.600 185.575 50.920 185.635 ;
        RECT 51.475 185.480 51.765 185.795 ;
        RECT 52.555 185.775 52.845 185.820 ;
        RECT 56.135 185.775 56.425 185.820 ;
        RECT 57.970 185.775 58.260 185.820 ;
        RECT 52.555 185.635 58.260 185.775 ;
        RECT 52.555 185.590 52.845 185.635 ;
        RECT 56.135 185.590 56.425 185.635 ;
        RECT 57.970 185.590 58.260 185.635 ;
        RECT 60.260 185.775 60.580 185.835 ;
        RECT 72.770 185.820 72.910 185.975 ;
        RECT 81.420 185.915 81.740 185.975 ;
        RECT 82.355 186.115 82.645 186.160 ;
        RECT 83.260 186.115 83.580 186.175 ;
        RECT 86.480 186.115 86.800 186.175 ;
        RECT 90.175 186.115 90.465 186.160 ;
        RECT 82.355 185.975 90.465 186.115 ;
        RECT 82.355 185.930 82.645 185.975 ;
        RECT 83.260 185.915 83.580 185.975 ;
        RECT 86.480 185.915 86.800 185.975 ;
        RECT 90.175 185.930 90.465 185.975 ;
        RECT 103.515 186.115 103.805 186.160 ;
        RECT 104.420 186.115 104.740 186.175 ;
        RECT 103.515 185.975 104.740 186.115 ;
        RECT 103.515 185.930 103.805 185.975 ;
        RECT 104.420 185.915 104.740 185.975 ;
        RECT 109.480 185.915 109.800 186.175 ;
        RECT 62.115 185.775 62.405 185.820 ;
        RECT 60.260 185.635 62.405 185.775 ;
        RECT 60.260 185.575 60.580 185.635 ;
        RECT 62.115 185.590 62.405 185.635 ;
        RECT 63.035 185.590 63.325 185.820 ;
        RECT 72.695 185.590 72.985 185.820 ;
        RECT 77.250 185.775 77.540 185.820 ;
        RECT 77.250 185.635 79.785 185.775 ;
        RECT 77.250 185.590 77.540 185.635 ;
        RECT 45.080 185.295 48.530 185.435 ;
        RECT 48.775 185.435 49.065 185.480 ;
        RECT 51.175 185.435 51.765 185.480 ;
        RECT 54.415 185.435 55.065 185.480 ;
        RECT 48.775 185.295 55.065 185.435 ;
        RECT 45.080 185.235 45.400 185.295 ;
        RECT 48.775 185.250 49.065 185.295 ;
        RECT 51.175 185.250 51.465 185.295 ;
        RECT 54.415 185.250 55.065 185.295 ;
        RECT 60.720 185.235 61.040 185.495 ;
        RECT 61.640 185.435 61.960 185.495 ;
        RECT 63.110 185.435 63.250 185.590 ;
        RECT 79.570 185.480 79.785 185.635 ;
        RECT 80.500 185.575 80.820 185.835 ;
        RECT 88.335 185.590 88.625 185.820 ;
        RECT 90.640 185.775 90.930 185.820 ;
        RECT 92.475 185.775 92.765 185.820 ;
        RECT 96.055 185.775 96.345 185.820 ;
        RECT 90.640 185.635 96.345 185.775 ;
        RECT 90.640 185.590 90.930 185.635 ;
        RECT 92.475 185.590 92.765 185.635 ;
        RECT 96.055 185.590 96.345 185.635 ;
        RECT 61.640 185.295 63.250 185.435 ;
        RECT 72.235 185.435 72.525 185.480 ;
        RECT 75.390 185.435 75.680 185.480 ;
        RECT 78.650 185.435 78.940 185.480 ;
        RECT 72.235 185.295 78.940 185.435 ;
        RECT 61.640 185.235 61.960 185.295 ;
        RECT 72.235 185.250 72.525 185.295 ;
        RECT 75.390 185.250 75.680 185.295 ;
        RECT 78.650 185.250 78.940 185.295 ;
        RECT 79.570 185.435 79.860 185.480 ;
        RECT 81.430 185.435 81.720 185.480 ;
        RECT 79.570 185.295 81.720 185.435 ;
        RECT 88.410 185.435 88.550 185.590 ;
        RECT 91.080 185.435 91.400 185.495 ;
        RECT 88.410 185.295 91.400 185.435 ;
        RECT 79.570 185.250 79.860 185.295 ;
        RECT 81.430 185.250 81.720 185.295 ;
        RECT 91.080 185.235 91.400 185.295 ;
        RECT 91.540 185.235 91.860 185.495 ;
        RECT 97.135 185.480 97.425 185.795 ;
        RECT 101.200 185.575 101.520 185.835 ;
        RECT 93.835 185.435 94.485 185.480 ;
        RECT 97.135 185.435 97.725 185.480 ;
        RECT 93.010 185.295 97.725 185.435 ;
        RECT 19.795 185.095 20.085 185.140 ;
        RECT 22.080 185.095 22.400 185.155 ;
        RECT 19.795 184.955 22.400 185.095 ;
        RECT 19.795 184.910 20.085 184.955 ;
        RECT 22.080 184.895 22.400 184.955 ;
        RECT 34.500 184.895 34.820 185.155 ;
        RECT 37.260 185.095 37.580 185.155 ;
        RECT 39.115 185.095 39.405 185.140 ;
        RECT 37.260 184.955 39.405 185.095 ;
        RECT 37.260 184.895 37.580 184.955 ;
        RECT 39.115 184.910 39.405 184.955 ;
        RECT 43.240 185.095 43.560 185.155 ;
        RECT 73.600 185.140 73.920 185.155 ;
        RECT 49.695 185.095 49.985 185.140 ;
        RECT 43.240 184.955 49.985 185.095 ;
        RECT 43.240 184.895 43.560 184.955 ;
        RECT 49.695 184.910 49.985 184.955 ;
        RECT 73.385 184.910 73.920 185.140 ;
        RECT 88.795 185.095 89.085 185.140 ;
        RECT 93.010 185.095 93.150 185.295 ;
        RECT 93.835 185.250 94.485 185.295 ;
        RECT 97.435 185.250 97.725 185.295 ;
        RECT 99.820 185.435 100.140 185.495 ;
        RECT 104.435 185.435 104.725 185.480 ;
        RECT 99.820 185.295 104.725 185.435 ;
        RECT 99.820 185.235 100.140 185.295 ;
        RECT 104.435 185.250 104.725 185.295 ;
        RECT 88.795 184.955 93.150 185.095 ;
        RECT 93.380 185.095 93.700 185.155 ;
        RECT 98.915 185.095 99.205 185.140 ;
        RECT 93.380 184.955 99.205 185.095 ;
        RECT 88.795 184.910 89.085 184.955 ;
        RECT 73.600 184.895 73.920 184.910 ;
        RECT 93.380 184.895 93.700 184.955 ;
        RECT 98.915 184.910 99.205 184.955 ;
        RECT 102.135 185.095 102.425 185.140 ;
        RECT 102.580 185.095 102.900 185.155 ;
        RECT 102.135 184.955 102.900 185.095 ;
        RECT 102.135 184.910 102.425 184.955 ;
        RECT 102.580 184.895 102.900 184.955 ;
        RECT 103.975 185.095 104.265 185.140 ;
        RECT 105.800 185.095 106.120 185.155 ;
        RECT 106.735 185.095 107.025 185.140 ;
        RECT 103.975 184.955 107.025 185.095 ;
        RECT 103.975 184.910 104.265 184.955 ;
        RECT 105.800 184.895 106.120 184.955 ;
        RECT 106.735 184.910 107.025 184.955 ;
        RECT 10.510 184.275 115.850 184.755 ;
        RECT 24.840 184.075 25.160 184.135 ;
        RECT 26.235 184.075 26.525 184.120 ;
        RECT 24.840 183.935 26.525 184.075 ;
        RECT 24.840 183.875 25.160 183.935 ;
        RECT 26.235 183.890 26.525 183.935 ;
        RECT 29.440 183.875 29.760 184.135 ;
        RECT 29.915 183.890 30.205 184.120 ;
        RECT 34.055 184.075 34.345 184.120 ;
        RECT 34.500 184.075 34.820 184.135 ;
        RECT 40.035 184.075 40.325 184.120 ;
        RECT 34.055 183.935 34.820 184.075 ;
        RECT 34.055 183.890 34.345 183.935 ;
        RECT 27.140 183.735 27.460 183.795 ;
        RECT 29.990 183.735 30.130 183.890 ;
        RECT 34.500 183.875 34.820 183.935 ;
        RECT 35.050 183.935 40.325 184.075 ;
        RECT 27.140 183.595 30.130 183.735 ;
        RECT 31.280 183.735 31.600 183.795 ;
        RECT 35.050 183.735 35.190 183.935 ;
        RECT 40.035 183.890 40.325 183.935 ;
        RECT 41.875 184.075 42.165 184.120 ;
        RECT 41.875 183.935 45.770 184.075 ;
        RECT 41.875 183.890 42.165 183.935 ;
        RECT 31.280 183.595 35.190 183.735 ;
        RECT 37.735 183.735 38.025 183.780 ;
        RECT 38.180 183.735 38.500 183.795 ;
        RECT 43.715 183.735 44.005 183.780 ;
        RECT 37.735 183.595 44.005 183.735 ;
        RECT 45.630 183.735 45.770 183.935 ;
        RECT 46.000 183.875 46.320 184.135 ;
        RECT 50.615 184.075 50.905 184.120 ;
        RECT 54.740 184.075 55.060 184.135 ;
        RECT 50.615 183.935 55.060 184.075 ;
        RECT 50.615 183.890 50.905 183.935 ;
        RECT 54.740 183.875 55.060 183.935 ;
        RECT 58.880 184.075 59.200 184.135 ;
        RECT 73.600 184.075 73.920 184.135 ;
        RECT 74.075 184.075 74.365 184.120 ;
        RECT 58.880 183.935 63.710 184.075 ;
        RECT 58.880 183.875 59.200 183.935 ;
        RECT 49.220 183.735 49.540 183.795 ;
        RECT 45.630 183.595 49.540 183.735 ;
        RECT 27.140 183.535 27.460 183.595 ;
        RECT 31.280 183.535 31.600 183.595 ;
        RECT 37.735 183.550 38.025 183.595 ;
        RECT 38.180 183.535 38.500 183.595 ;
        RECT 43.715 183.550 44.005 183.595 ;
        RECT 49.220 183.535 49.540 183.595 ;
        RECT 57.960 183.735 58.280 183.795 ;
        RECT 57.960 183.595 62.790 183.735 ;
        RECT 57.960 183.535 58.280 183.595 ;
        RECT 19.320 183.395 19.640 183.455 ;
        RECT 23.920 183.395 24.240 183.455 ;
        RECT 26.695 183.395 26.985 183.440 ;
        RECT 19.320 183.255 26.985 183.395 ;
        RECT 19.320 183.195 19.640 183.255 ;
        RECT 23.920 183.195 24.240 183.255 ;
        RECT 26.695 183.210 26.985 183.255 ;
        RECT 28.535 183.395 28.825 183.440 ;
        RECT 30.360 183.395 30.680 183.455 ;
        RECT 28.535 183.255 30.680 183.395 ;
        RECT 28.535 183.210 28.825 183.255 ;
        RECT 30.360 183.195 30.680 183.255 ;
        RECT 30.820 183.195 31.140 183.455 ;
        RECT 27.600 183.055 27.920 183.115 ;
        RECT 31.370 183.055 31.510 183.535 ;
        RECT 32.660 183.395 32.980 183.455 ;
        RECT 33.135 183.395 33.425 183.440 ;
        RECT 32.660 183.255 33.425 183.395 ;
        RECT 32.660 183.195 32.980 183.255 ;
        RECT 33.135 183.210 33.425 183.255 ;
        RECT 34.975 183.395 35.265 183.440 ;
        RECT 37.260 183.395 37.580 183.455 ;
        RECT 34.975 183.255 37.580 183.395 ;
        RECT 34.975 183.210 35.265 183.255 ;
        RECT 37.260 183.195 37.580 183.255 ;
        RECT 39.575 183.395 39.865 183.440 ;
        RECT 44.175 183.395 44.465 183.440 ;
        RECT 44.620 183.395 44.940 183.455 ;
        RECT 39.575 183.255 43.930 183.395 ;
        RECT 39.575 183.210 39.865 183.255 ;
        RECT 43.790 183.115 43.930 183.255 ;
        RECT 44.175 183.255 44.940 183.395 ;
        RECT 44.175 183.210 44.465 183.255 ;
        RECT 44.620 183.195 44.940 183.255 ;
        RECT 46.460 183.395 46.780 183.455 ;
        RECT 48.315 183.395 48.605 183.440 ;
        RECT 46.460 183.255 48.605 183.395 ;
        RECT 46.460 183.195 46.780 183.255 ;
        RECT 48.315 183.210 48.605 183.255 ;
        RECT 48.775 183.210 49.065 183.440 ;
        RECT 51.535 183.395 51.825 183.440 ;
        RECT 51.980 183.395 52.300 183.455 ;
        RECT 51.535 183.255 52.300 183.395 ;
        RECT 51.535 183.210 51.825 183.255 ;
        RECT 38.655 183.055 38.945 183.100 ;
        RECT 39.100 183.055 39.420 183.115 ;
        RECT 42.795 183.055 43.085 183.100 ;
        RECT 43.700 183.055 44.020 183.115 ;
        RECT 27.600 182.915 31.510 183.055 ;
        RECT 38.270 182.915 43.470 183.055 ;
        RECT 27.600 182.855 27.920 182.915 ;
        RECT 27.140 182.715 27.460 182.775 ;
        RECT 38.270 182.715 38.410 182.915 ;
        RECT 38.655 182.870 38.945 182.915 ;
        RECT 39.100 182.855 39.420 182.915 ;
        RECT 42.795 182.870 43.085 182.915 ;
        RECT 27.140 182.575 38.410 182.715 ;
        RECT 43.330 182.715 43.470 182.915 ;
        RECT 43.700 182.915 47.610 183.055 ;
        RECT 43.700 182.855 44.020 182.915 ;
        RECT 47.470 182.715 47.610 182.915 ;
        RECT 47.840 182.855 48.160 183.115 ;
        RECT 48.850 183.055 48.990 183.210 ;
        RECT 51.980 183.195 52.300 183.255 ;
        RECT 58.420 183.195 58.740 183.455 ;
        RECT 59.800 183.195 60.120 183.455 ;
        RECT 48.390 182.915 48.990 183.055 ;
        RECT 48.390 182.715 48.530 182.915 ;
        RECT 58.895 182.870 59.185 183.100 ;
        RECT 59.355 183.055 59.645 183.100 ;
        RECT 61.640 183.055 61.960 183.115 ;
        RECT 59.355 182.915 61.960 183.055 ;
        RECT 59.355 182.870 59.645 182.915 ;
        RECT 43.330 182.575 47.150 182.715 ;
        RECT 47.470 182.575 48.530 182.715 ;
        RECT 58.970 182.715 59.110 182.870 ;
        RECT 61.640 182.855 61.960 182.915 ;
        RECT 62.100 182.855 62.420 183.115 ;
        RECT 62.650 183.055 62.790 183.595 ;
        RECT 63.020 183.195 63.340 183.455 ;
        RECT 63.570 183.440 63.710 183.935 ;
        RECT 73.600 183.935 74.365 184.075 ;
        RECT 73.600 183.875 73.920 183.935 ;
        RECT 74.075 183.890 74.365 183.935 ;
        RECT 76.375 184.075 76.665 184.120 ;
        RECT 80.500 184.075 80.820 184.135 ;
        RECT 80.975 184.075 81.265 184.120 ;
        RECT 76.375 183.935 80.270 184.075 ;
        RECT 76.375 183.890 76.665 183.935 ;
        RECT 63.940 183.735 64.260 183.795 ;
        RECT 66.255 183.735 66.545 183.780 ;
        RECT 63.940 183.595 66.545 183.735 ;
        RECT 63.940 183.535 64.260 183.595 ;
        RECT 66.255 183.550 66.545 183.595 ;
        RECT 69.000 183.735 69.320 183.795 ;
        RECT 69.935 183.735 70.225 183.780 ;
        RECT 69.000 183.595 70.225 183.735 ;
        RECT 69.000 183.535 69.320 183.595 ;
        RECT 69.935 183.550 70.225 183.595 ;
        RECT 70.470 183.595 77.510 183.735 ;
        RECT 63.495 183.210 63.785 183.440 ;
        RECT 64.860 183.395 65.180 183.455 ;
        RECT 67.160 183.395 67.480 183.455 ;
        RECT 64.860 183.255 67.480 183.395 ;
        RECT 64.860 183.195 65.180 183.255 ;
        RECT 67.160 183.195 67.480 183.255 ;
        RECT 67.620 183.195 67.940 183.455 ;
        RECT 70.470 183.055 70.610 183.595 ;
        RECT 74.060 183.395 74.380 183.455 ;
        RECT 77.370 183.440 77.510 183.595 ;
        RECT 80.130 183.440 80.270 183.935 ;
        RECT 80.500 183.935 81.265 184.075 ;
        RECT 80.500 183.875 80.820 183.935 ;
        RECT 80.975 183.890 81.265 183.935 ;
        RECT 93.380 184.075 93.700 184.135 ;
        RECT 94.775 184.075 95.065 184.120 ;
        RECT 93.380 183.935 95.065 184.075 ;
        RECT 93.380 183.875 93.700 183.935 ;
        RECT 94.775 183.890 95.065 183.935 ;
        RECT 100.280 183.875 100.600 184.135 ;
        RECT 101.200 184.075 101.520 184.135 ;
        RECT 102.135 184.075 102.425 184.120 ;
        RECT 101.200 183.935 102.425 184.075 ;
        RECT 101.200 183.875 101.520 183.935 ;
        RECT 102.135 183.890 102.425 183.935 ;
        RECT 83.260 183.535 83.580 183.795 ;
        RECT 85.675 183.735 85.965 183.780 ;
        RECT 88.915 183.735 89.565 183.780 ;
        RECT 85.675 183.595 89.565 183.735 ;
        RECT 85.675 183.550 86.265 183.595 ;
        RECT 88.915 183.550 89.565 183.595 ;
        RECT 94.300 183.735 94.620 183.795 ;
        RECT 95.235 183.735 95.525 183.780 ;
        RECT 99.835 183.735 100.125 183.780 ;
        RECT 94.300 183.595 100.125 183.735 ;
        RECT 85.975 183.455 86.265 183.550 ;
        RECT 94.300 183.535 94.620 183.595 ;
        RECT 95.235 183.550 95.525 183.595 ;
        RECT 99.835 183.550 100.125 183.595 ;
        RECT 106.835 183.735 107.125 183.780 ;
        RECT 110.075 183.735 110.725 183.780 ;
        RECT 106.835 183.595 110.725 183.735 ;
        RECT 106.835 183.550 107.425 183.595 ;
        RECT 110.075 183.550 110.725 183.595 ;
        RECT 107.135 183.455 107.425 183.550 ;
        RECT 74.535 183.395 74.825 183.440 ;
        RECT 74.060 183.255 74.825 183.395 ;
        RECT 74.060 183.195 74.380 183.255 ;
        RECT 74.535 183.210 74.825 183.255 ;
        RECT 77.295 183.210 77.585 183.440 ;
        RECT 80.055 183.210 80.345 183.440 ;
        RECT 85.975 183.235 86.340 183.455 ;
        RECT 86.020 183.195 86.340 183.235 ;
        RECT 87.055 183.395 87.345 183.440 ;
        RECT 90.635 183.395 90.925 183.440 ;
        RECT 92.470 183.395 92.760 183.440 ;
        RECT 87.055 183.255 92.760 183.395 ;
        RECT 87.055 183.210 87.345 183.255 ;
        RECT 90.635 183.210 90.925 183.255 ;
        RECT 92.470 183.210 92.760 183.255 ;
        RECT 103.975 183.395 104.265 183.440 ;
        RECT 104.880 183.395 105.200 183.455 ;
        RECT 103.975 183.255 105.200 183.395 ;
        RECT 103.975 183.210 104.265 183.255 ;
        RECT 104.880 183.195 105.200 183.255 ;
        RECT 107.135 183.235 107.500 183.455 ;
        RECT 107.180 183.195 107.500 183.235 ;
        RECT 108.215 183.395 108.505 183.440 ;
        RECT 111.795 183.395 112.085 183.440 ;
        RECT 113.630 183.395 113.920 183.440 ;
        RECT 108.215 183.255 113.920 183.395 ;
        RECT 108.215 183.210 108.505 183.255 ;
        RECT 111.795 183.210 112.085 183.255 ;
        RECT 113.630 183.210 113.920 183.255 ;
        RECT 62.650 182.915 70.610 183.055 ;
        RECT 73.140 183.055 73.460 183.115 ;
        RECT 74.980 183.055 75.300 183.115 ;
        RECT 73.140 182.915 75.300 183.055 ;
        RECT 73.140 182.855 73.460 182.915 ;
        RECT 74.980 182.855 75.300 182.915 ;
        RECT 78.675 183.055 78.965 183.100 ;
        RECT 81.880 183.055 82.200 183.115 ;
        RECT 78.675 182.915 82.200 183.055 ;
        RECT 78.675 182.870 78.965 182.915 ;
        RECT 81.880 182.855 82.200 182.915 ;
        RECT 86.480 183.055 86.800 183.115 ;
        RECT 92.935 183.055 93.225 183.100 ;
        RECT 86.480 182.915 93.225 183.055 ;
        RECT 86.480 182.855 86.800 182.915 ;
        RECT 92.935 182.870 93.225 182.915 ;
        RECT 94.315 183.055 94.605 183.100 ;
        RECT 99.375 183.055 99.665 183.100 ;
        RECT 94.315 182.915 99.665 183.055 ;
        RECT 94.315 182.870 94.605 182.915 ;
        RECT 99.375 182.870 99.665 182.915 ;
        RECT 60.260 182.715 60.580 182.775 ;
        RECT 60.735 182.715 61.025 182.760 ;
        RECT 58.970 182.575 61.025 182.715 ;
        RECT 61.730 182.715 61.870 182.855 ;
        RECT 64.860 182.715 65.180 182.775 ;
        RECT 61.730 182.575 65.180 182.715 ;
        RECT 27.140 182.515 27.460 182.575 ;
        RECT 47.010 182.375 47.150 182.575 ;
        RECT 60.260 182.515 60.580 182.575 ;
        RECT 60.735 182.530 61.025 182.575 ;
        RECT 64.860 182.515 65.180 182.575 ;
        RECT 69.935 182.715 70.225 182.760 ;
        RECT 70.840 182.715 71.160 182.775 ;
        RECT 69.935 182.575 71.160 182.715 ;
        RECT 69.935 182.530 70.225 182.575 ;
        RECT 70.840 182.515 71.160 182.575 ;
        RECT 87.055 182.715 87.345 182.760 ;
        RECT 90.175 182.715 90.465 182.760 ;
        RECT 92.065 182.715 92.355 182.760 ;
        RECT 87.055 182.575 92.355 182.715 ;
        RECT 87.055 182.530 87.345 182.575 ;
        RECT 90.175 182.530 90.465 182.575 ;
        RECT 92.065 182.530 92.355 182.575 ;
        RECT 47.840 182.375 48.160 182.435 ;
        RECT 47.010 182.235 48.160 182.375 ;
        RECT 47.840 182.175 48.160 182.235 ;
        RECT 52.455 182.375 52.745 182.420 ;
        RECT 52.900 182.375 53.220 182.435 ;
        RECT 52.455 182.235 53.220 182.375 ;
        RECT 52.455 182.190 52.745 182.235 ;
        RECT 52.900 182.175 53.220 182.235 ;
        RECT 57.515 182.375 57.805 182.420 ;
        RECT 58.420 182.375 58.740 182.435 ;
        RECT 57.515 182.235 58.740 182.375 ;
        RECT 57.515 182.190 57.805 182.235 ;
        RECT 58.420 182.175 58.740 182.235 ;
        RECT 73.140 182.375 73.460 182.435 ;
        RECT 84.195 182.375 84.485 182.420 ;
        RECT 85.560 182.375 85.880 182.435 ;
        RECT 73.140 182.235 85.880 182.375 ;
        RECT 73.140 182.175 73.460 182.235 ;
        RECT 84.195 182.190 84.485 182.235 ;
        RECT 85.560 182.175 85.880 182.235 ;
        RECT 89.240 182.375 89.560 182.435 ;
        RECT 91.620 182.375 91.910 182.420 ;
        RECT 89.240 182.235 91.910 182.375 ;
        RECT 89.240 182.175 89.560 182.235 ;
        RECT 91.620 182.190 91.910 182.235 ;
        RECT 92.460 182.375 92.780 182.435 ;
        RECT 94.390 182.375 94.530 182.870 ;
        RECT 99.450 182.715 99.590 182.870 ;
        RECT 103.500 182.855 103.820 183.115 ;
        RECT 107.640 183.055 107.960 183.115 ;
        RECT 114.080 183.055 114.400 183.115 ;
        RECT 107.640 182.915 114.400 183.055 ;
        RECT 107.640 182.855 107.960 182.915 ;
        RECT 114.080 182.855 114.400 182.915 ;
        RECT 104.420 182.715 104.740 182.775 ;
        RECT 99.450 182.575 104.740 182.715 ;
        RECT 104.420 182.515 104.740 182.575 ;
        RECT 108.215 182.715 108.505 182.760 ;
        RECT 111.335 182.715 111.625 182.760 ;
        RECT 113.225 182.715 113.515 182.760 ;
        RECT 108.215 182.575 113.515 182.715 ;
        RECT 108.215 182.530 108.505 182.575 ;
        RECT 111.335 182.530 111.625 182.575 ;
        RECT 113.225 182.530 113.515 182.575 ;
        RECT 92.460 182.235 94.530 182.375 ;
        RECT 96.140 182.375 96.460 182.435 ;
        RECT 97.075 182.375 97.365 182.420 ;
        RECT 96.140 182.235 97.365 182.375 ;
        RECT 92.460 182.175 92.780 182.235 ;
        RECT 96.140 182.175 96.460 182.235 ;
        RECT 97.075 182.190 97.365 182.235 ;
        RECT 100.740 182.375 101.060 182.435 ;
        RECT 112.700 182.420 113.020 182.435 ;
        RECT 105.355 182.375 105.645 182.420 ;
        RECT 100.740 182.235 105.645 182.375 ;
        RECT 100.740 182.175 101.060 182.235 ;
        RECT 105.355 182.190 105.645 182.235 ;
        RECT 112.700 182.190 113.070 182.420 ;
        RECT 112.700 182.175 113.020 182.190 ;
        RECT 10.510 181.555 115.850 182.035 ;
        RECT 30.820 181.155 31.140 181.415 ;
        RECT 44.620 181.155 44.940 181.415 ;
        RECT 53.820 181.355 54.140 181.415 ;
        RECT 45.170 181.215 54.140 181.355 ;
        RECT 29.440 181.015 29.760 181.075 ;
        RECT 31.280 181.015 31.600 181.075 ;
        RECT 45.170 181.015 45.310 181.215 ;
        RECT 53.820 181.155 54.140 181.215 ;
        RECT 59.800 181.355 60.120 181.415 ;
        RECT 62.100 181.355 62.420 181.415 ;
        RECT 67.620 181.355 67.940 181.415 ;
        RECT 59.800 181.215 62.420 181.355 ;
        RECT 59.800 181.155 60.120 181.215 ;
        RECT 62.100 181.155 62.420 181.215 ;
        RECT 62.650 181.215 67.940 181.355 ;
        RECT 29.440 180.875 45.310 181.015 ;
        RECT 48.415 181.015 48.705 181.060 ;
        RECT 51.535 181.015 51.825 181.060 ;
        RECT 53.425 181.015 53.715 181.060 ;
        RECT 48.415 180.875 53.715 181.015 ;
        RECT 29.440 180.815 29.760 180.875 ;
        RECT 31.280 180.815 31.600 180.875 ;
        RECT 27.140 180.675 27.460 180.735 ;
        RECT 27.615 180.675 27.905 180.720 ;
        RECT 27.140 180.535 27.905 180.675 ;
        RECT 27.140 180.475 27.460 180.535 ;
        RECT 27.615 180.490 27.905 180.535 ;
        RECT 34.040 180.675 34.360 180.735 ;
        RECT 34.040 180.535 35.650 180.675 ;
        RECT 34.040 180.475 34.360 180.535 ;
        RECT 20.255 180.335 20.545 180.380 ;
        RECT 22.080 180.335 22.400 180.395 ;
        RECT 20.255 180.195 22.400 180.335 ;
        RECT 20.255 180.150 20.545 180.195 ;
        RECT 22.080 180.135 22.400 180.195 ;
        RECT 23.935 180.335 24.225 180.380 ;
        RECT 30.360 180.335 30.680 180.395 ;
        RECT 23.935 180.195 30.680 180.335 ;
        RECT 23.935 180.150 24.225 180.195 ;
        RECT 30.360 180.135 30.680 180.195 ;
        RECT 31.295 180.150 31.585 180.380 ;
        RECT 26.695 179.995 26.985 180.040 ;
        RECT 31.370 179.995 31.510 180.150 ;
        RECT 34.500 180.135 34.820 180.395 ;
        RECT 35.510 180.380 35.650 180.535 ;
        RECT 36.430 180.380 36.570 180.875 ;
        RECT 48.415 180.830 48.705 180.875 ;
        RECT 51.535 180.830 51.825 180.875 ;
        RECT 53.425 180.830 53.715 180.875 ;
        RECT 60.260 181.015 60.580 181.075 ;
        RECT 62.650 181.015 62.790 181.215 ;
        RECT 67.620 181.155 67.940 181.215 ;
        RECT 86.480 181.355 86.800 181.415 ;
        RECT 90.635 181.355 90.925 181.400 ;
        RECT 86.480 181.215 90.925 181.355 ;
        RECT 86.480 181.155 86.800 181.215 ;
        RECT 90.635 181.170 90.925 181.215 ;
        RECT 91.540 181.155 91.860 181.415 ;
        RECT 107.180 181.355 107.500 181.415 ;
        RECT 108.575 181.355 108.865 181.400 ;
        RECT 107.180 181.215 108.865 181.355 ;
        RECT 107.180 181.155 107.500 181.215 ;
        RECT 108.575 181.170 108.865 181.215 ;
        RECT 111.335 181.355 111.625 181.400 ;
        RECT 112.700 181.355 113.020 181.415 ;
        RECT 111.335 181.215 113.020 181.355 ;
        RECT 111.335 181.170 111.625 181.215 ;
        RECT 112.700 181.155 113.020 181.215 ;
        RECT 60.260 180.875 62.790 181.015 ;
        RECT 60.260 180.815 60.580 180.875 ;
        RECT 39.560 180.675 39.880 180.735 ;
        RECT 41.415 180.675 41.705 180.720 ;
        RECT 45.080 180.675 45.400 180.735 ;
        RECT 45.555 180.675 45.845 180.720 ;
        RECT 39.560 180.535 45.845 180.675 ;
        RECT 39.560 180.475 39.880 180.535 ;
        RECT 41.415 180.490 41.705 180.535 ;
        RECT 45.080 180.475 45.400 180.535 ;
        RECT 45.555 180.490 45.845 180.535 ;
        RECT 52.900 180.475 53.220 180.735 ;
        RECT 58.880 180.675 59.200 180.735 ;
        RECT 61.195 180.675 61.485 180.720 ;
        RECT 58.880 180.535 61.485 180.675 ;
        RECT 58.880 180.475 59.200 180.535 ;
        RECT 61.195 180.490 61.485 180.535 ;
        RECT 61.640 180.475 61.960 180.735 ;
        RECT 62.100 180.475 62.420 180.735 ;
        RECT 62.650 180.720 62.790 180.875 ;
        RECT 63.020 180.815 63.340 181.075 ;
        RECT 77.395 181.015 77.685 181.060 ;
        RECT 80.515 181.015 80.805 181.060 ;
        RECT 82.405 181.015 82.695 181.060 ;
        RECT 77.395 180.875 82.695 181.015 ;
        RECT 77.395 180.830 77.685 180.875 ;
        RECT 80.515 180.830 80.805 180.875 ;
        RECT 82.405 180.830 82.695 180.875 ;
        RECT 101.775 181.015 102.065 181.060 ;
        RECT 104.895 181.015 105.185 181.060 ;
        RECT 106.785 181.015 107.075 181.060 ;
        RECT 101.775 180.875 107.075 181.015 ;
        RECT 101.775 180.830 102.065 180.875 ;
        RECT 104.895 180.830 105.185 180.875 ;
        RECT 106.785 180.830 107.075 180.875 ;
        RECT 62.575 180.490 62.865 180.720 ;
        RECT 35.435 180.150 35.725 180.380 ;
        RECT 35.895 180.150 36.185 180.380 ;
        RECT 36.355 180.150 36.645 180.380 ;
        RECT 40.955 180.335 41.245 180.380 ;
        RECT 44.160 180.335 44.480 180.395 ;
        RECT 40.955 180.195 44.480 180.335 ;
        RECT 40.955 180.150 41.245 180.195 ;
        RECT 26.695 179.855 31.510 179.995 ;
        RECT 33.580 179.995 33.900 180.055 ;
        RECT 35.970 179.995 36.110 180.150 ;
        RECT 44.160 180.135 44.480 180.195 ;
        RECT 47.335 180.040 47.625 180.355 ;
        RECT 48.415 180.335 48.705 180.380 ;
        RECT 51.995 180.335 52.285 180.380 ;
        RECT 53.830 180.335 54.120 180.380 ;
        RECT 48.415 180.195 54.120 180.335 ;
        RECT 48.415 180.150 48.705 180.195 ;
        RECT 51.995 180.150 52.285 180.195 ;
        RECT 53.830 180.150 54.120 180.195 ;
        RECT 54.295 180.150 54.585 180.380 ;
        RECT 59.355 180.335 59.645 180.380 ;
        RECT 63.110 180.335 63.250 180.815 ;
        RECT 63.480 180.475 63.800 180.735 ;
        RECT 79.120 180.675 79.440 180.735 ;
        RECT 69.550 180.535 79.440 180.675 ;
        RECT 59.355 180.195 63.250 180.335 ;
        RECT 59.355 180.150 59.645 180.195 ;
        RECT 33.580 179.855 36.110 179.995 ;
        RECT 40.495 179.995 40.785 180.040 ;
        RECT 47.035 179.995 47.625 180.040 ;
        RECT 50.275 179.995 50.925 180.040 ;
        RECT 40.495 179.855 50.925 179.995 ;
        RECT 26.695 179.810 26.985 179.855 ;
        RECT 33.580 179.795 33.900 179.855 ;
        RECT 40.495 179.810 40.785 179.855 ;
        RECT 47.035 179.810 47.325 179.855 ;
        RECT 50.275 179.810 50.925 179.855 ;
        RECT 53.360 179.995 53.680 180.055 ;
        RECT 54.370 179.995 54.510 180.150 ;
        RECT 53.360 179.855 54.510 179.995 ;
        RECT 61.640 179.995 61.960 180.055 ;
        RECT 69.550 179.995 69.690 180.535 ;
        RECT 79.120 180.475 79.440 180.535 ;
        RECT 83.260 180.475 83.580 180.735 ;
        RECT 89.255 180.675 89.545 180.720 ;
        RECT 93.380 180.675 93.700 180.735 ;
        RECT 89.255 180.535 93.700 180.675 ;
        RECT 89.255 180.490 89.545 180.535 ;
        RECT 93.380 180.475 93.700 180.535 ;
        RECT 96.140 180.475 96.460 180.735 ;
        RECT 102.580 180.675 102.900 180.735 ;
        RECT 106.275 180.675 106.565 180.720 ;
        RECT 102.580 180.535 106.565 180.675 ;
        RECT 102.580 180.475 102.900 180.535 ;
        RECT 106.275 180.490 106.565 180.535 ;
        RECT 71.775 180.335 72.065 180.380 ;
        RECT 74.980 180.335 75.300 180.395 ;
        RECT 71.775 180.195 75.300 180.335 ;
        RECT 71.775 180.150 72.065 180.195 ;
        RECT 74.980 180.135 75.300 180.195 ;
        RECT 61.640 179.855 69.690 179.995 ;
        RECT 53.360 179.795 53.680 179.855 ;
        RECT 61.640 179.795 61.960 179.855 ;
        RECT 69.920 179.795 70.240 180.055 ;
        RECT 76.315 180.040 76.605 180.355 ;
        RECT 77.395 180.335 77.685 180.380 ;
        RECT 80.975 180.335 81.265 180.380 ;
        RECT 82.810 180.335 83.100 180.380 ;
        RECT 77.395 180.195 83.100 180.335 ;
        RECT 77.395 180.150 77.685 180.195 ;
        RECT 80.975 180.150 81.265 180.195 ;
        RECT 82.810 180.150 83.100 180.195 ;
        RECT 84.640 180.135 84.960 180.395 ;
        RECT 91.080 180.135 91.400 180.395 ;
        RECT 92.475 180.335 92.765 180.380 ;
        RECT 92.935 180.335 93.225 180.380 ;
        RECT 92.475 180.195 93.225 180.335 ;
        RECT 92.475 180.150 92.765 180.195 ;
        RECT 92.935 180.150 93.225 180.195 ;
        RECT 76.015 179.995 76.605 180.040 ;
        RECT 79.255 179.995 79.905 180.040 ;
        RECT 81.420 179.995 81.740 180.055 ;
        RECT 100.695 180.040 100.985 180.355 ;
        RECT 101.775 180.335 102.065 180.380 ;
        RECT 105.355 180.335 105.645 180.380 ;
        RECT 107.190 180.335 107.480 180.380 ;
        RECT 101.775 180.195 107.480 180.335 ;
        RECT 101.775 180.150 102.065 180.195 ;
        RECT 105.355 180.150 105.645 180.195 ;
        RECT 107.190 180.150 107.480 180.195 ;
        RECT 107.640 180.135 107.960 180.395 ;
        RECT 108.115 180.150 108.405 180.380 ;
        RECT 76.015 179.855 81.740 179.995 ;
        RECT 76.015 179.810 76.305 179.855 ;
        RECT 79.255 179.810 79.905 179.855 ;
        RECT 81.420 179.795 81.740 179.855 ;
        RECT 81.895 179.810 82.185 180.040 ;
        RECT 100.395 179.995 100.985 180.040 ;
        RECT 103.500 180.040 103.820 180.055 ;
        RECT 103.500 179.995 104.285 180.040 ;
        RECT 100.395 179.855 104.285 179.995 ;
        RECT 100.395 179.810 100.685 179.855 ;
        RECT 103.500 179.810 104.285 179.855 ;
        RECT 104.880 179.995 105.200 180.055 ;
        RECT 108.190 179.995 108.330 180.150 ;
        RECT 110.400 180.135 110.720 180.395 ;
        RECT 104.880 179.855 108.330 179.995 ;
        RECT 23.015 179.655 23.305 179.700 ;
        RECT 28.520 179.655 28.840 179.715 ;
        RECT 23.015 179.515 28.840 179.655 ;
        RECT 23.015 179.470 23.305 179.515 ;
        RECT 28.520 179.455 28.840 179.515 ;
        RECT 28.980 179.455 29.300 179.715 ;
        RECT 31.740 179.655 32.060 179.715 ;
        RECT 32.215 179.655 32.505 179.700 ;
        RECT 31.740 179.515 32.505 179.655 ;
        RECT 31.740 179.455 32.060 179.515 ;
        RECT 32.215 179.470 32.505 179.515 ;
        RECT 37.260 179.655 37.580 179.715 ;
        RECT 37.735 179.655 38.025 179.700 ;
        RECT 37.260 179.515 38.025 179.655 ;
        RECT 37.260 179.455 37.580 179.515 ;
        RECT 37.735 179.470 38.025 179.515 ;
        RECT 59.815 179.655 60.105 179.700 ;
        RECT 64.400 179.655 64.720 179.715 ;
        RECT 67.160 179.655 67.480 179.715 ;
        RECT 59.815 179.515 67.480 179.655 ;
        RECT 59.815 179.470 60.105 179.515 ;
        RECT 64.400 179.455 64.720 179.515 ;
        RECT 67.160 179.455 67.480 179.515 ;
        RECT 69.460 179.655 69.780 179.715 ;
        RECT 72.220 179.655 72.540 179.715 ;
        RECT 74.535 179.655 74.825 179.700 ;
        RECT 69.460 179.515 74.825 179.655 ;
        RECT 81.970 179.655 82.110 179.810 ;
        RECT 103.500 179.795 103.820 179.810 ;
        RECT 104.880 179.795 105.200 179.855 ;
        RECT 83.735 179.655 84.025 179.700 ;
        RECT 81.970 179.515 84.025 179.655 ;
        RECT 69.460 179.455 69.780 179.515 ;
        RECT 72.220 179.455 72.540 179.515 ;
        RECT 74.535 179.470 74.825 179.515 ;
        RECT 83.735 179.470 84.025 179.515 ;
        RECT 86.020 179.455 86.340 179.715 ;
        RECT 97.060 179.655 97.380 179.715 ;
        RECT 98.915 179.655 99.205 179.700 ;
        RECT 97.060 179.515 99.205 179.655 ;
        RECT 97.060 179.455 97.380 179.515 ;
        RECT 98.915 179.470 99.205 179.515 ;
        RECT 10.510 178.835 115.850 179.315 ;
        RECT 27.140 178.635 27.460 178.695 ;
        RECT 22.170 178.495 30.130 178.635 ;
        RECT 19.320 177.955 19.640 178.015 ;
        RECT 20.715 177.955 21.005 178.000 ;
        RECT 19.320 177.815 21.005 177.955 ;
        RECT 19.320 177.755 19.640 177.815 ;
        RECT 20.715 177.770 21.005 177.815 ;
        RECT 15.180 177.615 15.500 177.675 ;
        RECT 22.170 177.660 22.310 178.495 ;
        RECT 27.140 178.435 27.460 178.495 ;
        RECT 23.000 178.095 23.320 178.355 ;
        RECT 28.980 178.295 29.300 178.355 ;
        RECT 24.700 178.155 29.300 178.295 ;
        RECT 24.700 177.955 24.840 178.155 ;
        RECT 28.980 178.095 29.300 178.155 ;
        RECT 22.630 177.815 24.840 177.955 ;
        RECT 22.630 177.675 22.770 177.815 ;
        RECT 26.680 177.755 27.000 178.015 ;
        RECT 27.600 177.755 27.920 178.015 ;
        RECT 28.060 177.755 28.380 178.015 ;
        RECT 28.535 177.955 28.825 178.000 ;
        RECT 29.440 177.955 29.760 178.015 ;
        RECT 28.535 177.815 29.760 177.955 ;
        RECT 29.990 177.955 30.130 178.495 ;
        RECT 30.360 178.435 30.680 178.695 ;
        RECT 32.215 178.635 32.505 178.680 ;
        RECT 34.040 178.635 34.360 178.695 ;
        RECT 32.215 178.495 34.360 178.635 ;
        RECT 32.215 178.450 32.505 178.495 ;
        RECT 34.040 178.435 34.360 178.495 ;
        RECT 37.720 178.435 38.040 178.695 ;
        RECT 45.080 178.635 45.400 178.695 ;
        RECT 48.315 178.635 48.605 178.680 ;
        RECT 45.080 178.495 48.605 178.635 ;
        RECT 45.080 178.435 45.400 178.495 ;
        RECT 48.315 178.450 48.605 178.495 ;
        RECT 51.535 178.635 51.825 178.680 ;
        RECT 51.980 178.635 52.300 178.695 ;
        RECT 51.535 178.495 52.300 178.635 ;
        RECT 51.535 178.450 51.825 178.495 ;
        RECT 51.980 178.435 52.300 178.495 ;
        RECT 53.820 178.635 54.140 178.695 ;
        RECT 61.640 178.635 61.960 178.695 ;
        RECT 63.495 178.635 63.785 178.680 ;
        RECT 64.860 178.635 65.180 178.695 ;
        RECT 53.820 178.495 61.960 178.635 ;
        RECT 53.820 178.435 54.140 178.495 ;
        RECT 61.640 178.435 61.960 178.495 ;
        RECT 62.180 178.495 65.180 178.635 ;
        RECT 37.810 178.295 37.950 178.435 ;
        RECT 44.160 178.295 44.480 178.355 ;
        RECT 62.180 178.295 62.320 178.495 ;
        RECT 63.495 178.450 63.785 178.495 ;
        RECT 64.860 178.435 65.180 178.495 ;
        RECT 67.160 178.435 67.480 178.695 ;
        RECT 72.235 178.635 72.525 178.680 ;
        RECT 74.060 178.635 74.380 178.695 ;
        RECT 72.235 178.495 74.380 178.635 ;
        RECT 72.235 178.450 72.525 178.495 ;
        RECT 74.060 178.435 74.380 178.495 ;
        RECT 81.420 178.435 81.740 178.695 ;
        RECT 86.020 178.635 86.340 178.695 ;
        RECT 88.795 178.635 89.085 178.680 ;
        RECT 86.020 178.495 89.085 178.635 ;
        RECT 86.020 178.435 86.340 178.495 ;
        RECT 88.795 178.450 89.085 178.495 ;
        RECT 94.300 178.435 94.620 178.695 ;
        RECT 100.280 178.635 100.600 178.695 ;
        RECT 96.690 178.495 100.600 178.635 ;
        RECT 36.890 178.155 37.950 178.295 ;
        RECT 39.190 178.155 62.320 178.295 ;
        RECT 63.020 178.295 63.340 178.355 ;
        RECT 67.250 178.295 67.390 178.435 ;
        RECT 63.020 178.155 65.090 178.295 ;
        RECT 34.500 177.955 34.820 178.015 ;
        RECT 36.890 178.000 37.030 178.155 ;
        RECT 35.895 177.955 36.185 178.000 ;
        RECT 29.990 177.815 33.350 177.955 ;
        RECT 28.535 177.770 28.825 177.815 ;
        RECT 29.440 177.755 29.760 177.815 ;
        RECT 15.655 177.615 15.945 177.660 ;
        RECT 15.180 177.475 15.945 177.615 ;
        RECT 15.180 177.415 15.500 177.475 ;
        RECT 15.655 177.430 15.945 177.475 ;
        RECT 22.095 177.430 22.385 177.660 ;
        RECT 22.540 177.415 22.860 177.675 ;
        RECT 23.920 177.615 24.240 177.675 ;
        RECT 33.210 177.660 33.350 177.815 ;
        RECT 34.500 177.815 36.185 177.955 ;
        RECT 34.500 177.755 34.820 177.815 ;
        RECT 32.675 177.615 32.965 177.660 ;
        RECT 23.920 177.475 32.965 177.615 ;
        RECT 23.920 177.415 24.240 177.475 ;
        RECT 32.675 177.430 32.965 177.475 ;
        RECT 33.135 177.430 33.425 177.660 ;
        RECT 20.255 177.275 20.545 177.320 ;
        RECT 25.300 177.275 25.620 177.335 ;
        RECT 20.255 177.135 25.620 177.275 ;
        RECT 20.255 177.090 20.545 177.135 ;
        RECT 25.300 177.075 25.620 177.135 ;
        RECT 26.680 177.275 27.000 177.335 ;
        RECT 29.440 177.275 29.760 177.335 ;
        RECT 26.680 177.135 29.760 177.275 ;
        RECT 26.680 177.075 27.000 177.135 ;
        RECT 29.440 177.075 29.760 177.135 ;
        RECT 18.875 176.935 19.165 176.980 ;
        RECT 22.540 176.935 22.860 176.995 ;
        RECT 18.875 176.795 22.860 176.935 ;
        RECT 18.875 176.750 19.165 176.795 ;
        RECT 22.540 176.735 22.860 176.795 ;
        RECT 24.855 176.935 25.145 176.980 ;
        RECT 28.060 176.935 28.380 176.995 ;
        RECT 24.855 176.795 28.380 176.935 ;
        RECT 24.855 176.750 25.145 176.795 ;
        RECT 28.060 176.735 28.380 176.795 ;
        RECT 29.915 176.935 30.205 176.980 ;
        RECT 30.820 176.935 31.140 176.995 ;
        RECT 29.915 176.795 31.140 176.935 ;
        RECT 35.510 176.935 35.650 177.815 ;
        RECT 35.895 177.770 36.185 177.815 ;
        RECT 36.815 177.770 37.105 178.000 ;
        RECT 37.275 177.770 37.565 178.000 ;
        RECT 37.735 177.955 38.025 178.000 ;
        RECT 39.190 177.955 39.330 178.155 ;
        RECT 37.735 177.815 39.330 177.955 ;
        RECT 39.575 177.955 39.865 178.000 ;
        RECT 40.020 177.955 40.340 178.015 ;
        RECT 39.575 177.815 40.340 177.955 ;
        RECT 37.735 177.770 38.025 177.815 ;
        RECT 39.575 177.770 39.865 177.815 ;
        RECT 37.350 177.615 37.490 177.770 ;
        RECT 40.020 177.755 40.340 177.815 ;
        RECT 40.480 177.755 40.800 178.015 ;
        RECT 40.940 177.755 41.260 178.015 ;
        RECT 41.490 178.000 41.630 178.155 ;
        RECT 44.160 178.095 44.480 178.155 ;
        RECT 63.020 178.095 63.340 178.155 ;
        RECT 41.415 177.770 41.705 178.000 ;
        RECT 43.240 177.755 43.560 178.015 ;
        RECT 48.760 177.755 49.080 178.015 ;
        RECT 55.215 177.955 55.505 178.000 ;
        RECT 52.530 177.815 55.505 177.955 ;
        RECT 41.030 177.615 41.170 177.755 ;
        RECT 52.530 177.675 52.670 177.815 ;
        RECT 55.215 177.770 55.505 177.815 ;
        RECT 57.055 177.955 57.345 178.000 ;
        RECT 57.055 177.815 57.730 177.955 ;
        RECT 57.055 177.770 57.345 177.815 ;
        RECT 37.350 177.475 41.170 177.615 ;
        RECT 47.840 177.615 48.160 177.675 ;
        RECT 52.440 177.615 52.760 177.675 ;
        RECT 47.840 177.475 52.760 177.615 ;
        RECT 35.880 177.275 36.200 177.335 ;
        RECT 37.350 177.275 37.490 177.475 ;
        RECT 47.840 177.415 48.160 177.475 ;
        RECT 52.440 177.415 52.760 177.475 ;
        RECT 54.295 177.430 54.585 177.660 ;
        RECT 40.020 177.275 40.340 177.335 ;
        RECT 35.880 177.135 37.490 177.275 ;
        RECT 37.810 177.135 40.340 177.275 ;
        RECT 35.880 177.075 36.200 177.135 ;
        RECT 37.810 176.935 37.950 177.135 ;
        RECT 40.020 177.075 40.340 177.135 ;
        RECT 50.615 177.275 50.905 177.320 ;
        RECT 54.370 177.275 54.510 177.430 ;
        RECT 50.615 177.135 54.510 177.275 ;
        RECT 57.590 177.275 57.730 177.815 ;
        RECT 57.960 177.755 58.280 178.015 ;
        RECT 58.420 177.955 58.740 178.015 ;
        RECT 60.735 177.955 61.025 178.000 ;
        RECT 62.575 177.955 62.865 178.000 ;
        RECT 64.415 177.955 64.705 178.000 ;
        RECT 58.420 177.815 64.705 177.955 ;
        RECT 64.950 177.955 65.090 178.155 ;
        RECT 66.330 178.155 67.390 178.295 ;
        RECT 80.515 178.295 80.805 178.340 ;
        RECT 84.640 178.295 84.960 178.355 ;
        RECT 80.515 178.155 84.960 178.295 ;
        RECT 66.330 178.000 66.470 178.155 ;
        RECT 80.515 178.110 80.805 178.155 ;
        RECT 84.640 178.095 84.960 178.155 ;
        RECT 85.560 178.295 85.880 178.355 ;
        RECT 89.255 178.295 89.545 178.340 ;
        RECT 91.080 178.295 91.400 178.355 ;
        RECT 85.560 178.155 89.545 178.295 ;
        RECT 85.560 178.095 85.880 178.155 ;
        RECT 89.255 178.110 89.545 178.155 ;
        RECT 89.790 178.155 91.400 178.295 ;
        RECT 64.950 177.945 65.550 177.955 ;
        RECT 65.795 177.945 66.085 178.000 ;
        RECT 64.950 177.815 66.085 177.945 ;
        RECT 58.420 177.755 58.740 177.815 ;
        RECT 60.735 177.770 61.025 177.815 ;
        RECT 62.575 177.770 62.865 177.815 ;
        RECT 64.415 177.770 64.705 177.815 ;
        RECT 65.410 177.805 66.085 177.815 ;
        RECT 65.795 177.770 66.085 177.805 ;
        RECT 66.255 177.770 66.545 178.000 ;
        RECT 67.175 177.770 67.465 178.000 ;
        RECT 59.340 177.415 59.660 177.675 ;
        RECT 63.480 177.615 63.800 177.675 ;
        RECT 67.250 177.615 67.390 177.770 ;
        RECT 69.460 177.755 69.780 178.015 ;
        RECT 73.140 177.955 73.460 178.015 ;
        RECT 74.535 177.955 74.825 178.000 ;
        RECT 73.140 177.815 74.825 177.955 ;
        RECT 73.140 177.755 73.460 177.815 ;
        RECT 74.535 177.770 74.825 177.815 ;
        RECT 81.880 177.955 82.200 178.015 ;
        RECT 89.790 177.955 89.930 178.155 ;
        RECT 91.080 178.095 91.400 178.155 ;
        RECT 96.690 178.015 96.830 178.495 ;
        RECT 100.280 178.435 100.600 178.495 ;
        RECT 100.740 178.635 101.060 178.695 ;
        RECT 105.355 178.635 105.645 178.680 ;
        RECT 100.740 178.495 105.645 178.635 ;
        RECT 100.740 178.435 101.060 178.495 ;
        RECT 105.355 178.450 105.645 178.495 ;
        RECT 105.800 178.435 106.120 178.695 ;
        RECT 110.400 178.635 110.720 178.695 ;
        RECT 111.335 178.635 111.625 178.680 ;
        RECT 110.400 178.495 111.625 178.635 ;
        RECT 110.400 178.435 110.720 178.495 ;
        RECT 111.335 178.450 111.625 178.495 ;
        RECT 97.520 178.295 97.840 178.355 ;
        RECT 108.100 178.295 108.420 178.355 ;
        RECT 97.520 178.155 100.970 178.295 ;
        RECT 97.520 178.095 97.840 178.155 ;
        RECT 92.460 177.955 92.780 178.015 ;
        RECT 81.880 177.815 89.930 177.955 ;
        RECT 90.250 177.815 92.780 177.955 ;
        RECT 81.880 177.755 82.200 177.815 ;
        RECT 63.480 177.475 67.390 177.615 ;
        RECT 73.615 177.615 73.905 177.660 ;
        RECT 74.980 177.615 75.300 177.675 ;
        RECT 90.250 177.660 90.390 177.815 ;
        RECT 92.460 177.755 92.780 177.815 ;
        RECT 93.840 177.955 94.160 178.015 ;
        RECT 96.155 177.955 96.445 178.000 ;
        RECT 93.840 177.815 96.445 177.955 ;
        RECT 93.840 177.755 94.160 177.815 ;
        RECT 96.155 177.770 96.445 177.815 ;
        RECT 96.600 177.755 96.920 178.015 ;
        RECT 97.060 177.755 97.380 178.015 ;
        RECT 97.980 177.755 98.300 178.015 ;
        RECT 99.820 177.755 100.140 178.015 ;
        RECT 100.280 177.755 100.600 178.015 ;
        RECT 100.830 178.000 100.970 178.155 ;
        RECT 101.750 178.155 108.420 178.295 ;
        RECT 101.750 178.000 101.890 178.155 ;
        RECT 108.100 178.095 108.420 178.155 ;
        RECT 100.755 177.770 101.045 178.000 ;
        RECT 101.675 177.770 101.965 178.000 ;
        RECT 73.615 177.475 75.300 177.615 ;
        RECT 63.480 177.415 63.800 177.475 ;
        RECT 73.615 177.430 73.905 177.475 ;
        RECT 74.980 177.415 75.300 177.475 ;
        RECT 77.295 177.430 77.585 177.660 ;
        RECT 83.735 177.430 84.025 177.660 ;
        RECT 90.175 177.430 90.465 177.660 ;
        RECT 91.555 177.615 91.845 177.660 ;
        RECT 97.150 177.615 97.290 177.755 ;
        RECT 91.555 177.475 97.290 177.615 ;
        RECT 98.070 177.615 98.210 177.755 ;
        RECT 101.750 177.615 101.890 177.770 ;
        RECT 98.070 177.475 101.890 177.615 ;
        RECT 91.555 177.430 91.845 177.475 ;
        RECT 65.335 177.275 65.625 177.320 ;
        RECT 69.920 177.275 70.240 177.335 ;
        RECT 57.590 177.135 70.240 177.275 ;
        RECT 50.615 177.090 50.905 177.135 ;
        RECT 65.335 177.090 65.625 177.135 ;
        RECT 69.920 177.075 70.240 177.135 ;
        RECT 76.375 177.275 76.665 177.320 ;
        RECT 77.370 177.275 77.510 177.430 ;
        RECT 76.375 177.135 77.510 177.275 ;
        RECT 83.810 177.275 83.950 177.430 ;
        RECT 104.420 177.415 104.740 177.675 ;
        RECT 108.115 177.430 108.405 177.660 ;
        RECT 86.955 177.275 87.245 177.320 ;
        RECT 83.810 177.135 87.245 177.275 ;
        RECT 76.375 177.090 76.665 177.135 ;
        RECT 86.955 177.090 87.245 177.135 ;
        RECT 107.655 177.275 107.945 177.320 ;
        RECT 108.190 177.275 108.330 177.430 ;
        RECT 107.655 177.135 108.330 177.275 ;
        RECT 107.655 177.090 107.945 177.135 ;
        RECT 35.510 176.795 37.950 176.935 ;
        RECT 29.915 176.750 30.205 176.795 ;
        RECT 30.820 176.735 31.140 176.795 ;
        RECT 39.100 176.735 39.420 176.995 ;
        RECT 41.400 176.935 41.720 176.995 ;
        RECT 42.795 176.935 43.085 176.980 ;
        RECT 41.400 176.795 43.085 176.935 ;
        RECT 41.400 176.735 41.720 176.795 ;
        RECT 42.795 176.750 43.085 176.795 ;
        RECT 46.460 176.735 46.780 176.995 ;
        RECT 61.640 176.935 61.960 176.995 ;
        RECT 63.480 176.935 63.800 176.995 ;
        RECT 64.875 176.935 65.165 176.980 ;
        RECT 61.640 176.795 65.165 176.935 ;
        RECT 61.640 176.735 61.960 176.795 ;
        RECT 63.480 176.735 63.800 176.795 ;
        RECT 64.875 176.750 65.165 176.795 ;
        RECT 68.080 176.735 68.400 176.995 ;
        RECT 86.480 176.735 86.800 176.995 ;
        RECT 94.775 176.935 95.065 176.980 ;
        RECT 97.520 176.935 97.840 176.995 ;
        RECT 94.775 176.795 97.840 176.935 ;
        RECT 94.775 176.750 95.065 176.795 ;
        RECT 97.520 176.735 97.840 176.795 ;
        RECT 98.455 176.935 98.745 176.980 ;
        RECT 98.900 176.935 99.220 176.995 ;
        RECT 98.455 176.795 99.220 176.935 ;
        RECT 98.455 176.750 98.745 176.795 ;
        RECT 98.900 176.735 99.220 176.795 ;
        RECT 100.280 176.935 100.600 176.995 ;
        RECT 106.720 176.935 107.040 176.995 ;
        RECT 109.020 176.935 109.340 176.995 ;
        RECT 100.280 176.795 109.340 176.935 ;
        RECT 100.280 176.735 100.600 176.795 ;
        RECT 106.720 176.735 107.040 176.795 ;
        RECT 109.020 176.735 109.340 176.795 ;
        RECT 10.510 176.115 115.850 176.595 ;
        RECT 43.240 175.915 43.560 175.975 ;
        RECT 68.080 175.915 68.400 175.975 ;
        RECT 71.760 175.915 72.080 175.975 ;
        RECT 83.260 175.915 83.580 175.975 ;
        RECT 84.655 175.915 84.945 175.960 ;
        RECT 40.110 175.775 43.560 175.915 ;
        RECT 18.055 175.575 18.345 175.620 ;
        RECT 21.175 175.575 21.465 175.620 ;
        RECT 23.065 175.575 23.355 175.620 ;
        RECT 18.055 175.435 23.355 175.575 ;
        RECT 18.055 175.390 18.345 175.435 ;
        RECT 21.175 175.390 21.465 175.435 ;
        RECT 23.065 175.390 23.355 175.435 ;
        RECT 27.255 175.575 27.545 175.620 ;
        RECT 30.375 175.575 30.665 175.620 ;
        RECT 32.265 175.575 32.555 175.620 ;
        RECT 39.100 175.575 39.420 175.635 ;
        RECT 27.255 175.435 32.555 175.575 ;
        RECT 27.255 175.390 27.545 175.435 ;
        RECT 30.375 175.390 30.665 175.435 ;
        RECT 32.265 175.390 32.555 175.435 ;
        RECT 34.590 175.435 39.420 175.575 ;
        RECT 23.935 175.235 24.225 175.280 ;
        RECT 24.840 175.235 25.160 175.295 ;
        RECT 29.900 175.235 30.220 175.295 ;
        RECT 23.935 175.095 30.220 175.235 ;
        RECT 23.935 175.050 24.225 175.095 ;
        RECT 24.840 175.035 25.160 175.095 ;
        RECT 29.900 175.035 30.220 175.095 ;
        RECT 31.740 175.035 32.060 175.295 ;
        RECT 34.590 174.940 34.730 175.435 ;
        RECT 39.100 175.375 39.420 175.435 ;
        RECT 39.560 175.235 39.880 175.295 ;
        RECT 35.510 175.095 39.880 175.235 ;
        RECT 35.510 174.940 35.650 175.095 ;
        RECT 39.560 175.035 39.880 175.095 ;
        RECT 16.975 174.600 17.265 174.915 ;
        RECT 18.055 174.895 18.345 174.940 ;
        RECT 21.635 174.895 21.925 174.940 ;
        RECT 23.470 174.895 23.760 174.940 ;
        RECT 18.055 174.755 23.760 174.895 ;
        RECT 18.055 174.710 18.345 174.755 ;
        RECT 21.635 174.710 21.925 174.755 ;
        RECT 23.470 174.710 23.760 174.755 ;
        RECT 20.240 174.600 20.560 174.615 ;
        RECT 16.675 174.555 17.265 174.600 ;
        RECT 19.915 174.555 20.565 174.600 ;
        RECT 16.675 174.415 20.565 174.555 ;
        RECT 16.675 174.370 16.965 174.415 ;
        RECT 19.915 174.370 20.565 174.415 ;
        RECT 20.240 174.355 20.560 174.370 ;
        RECT 22.540 174.355 22.860 174.615 ;
        RECT 25.300 174.555 25.620 174.615 ;
        RECT 26.175 174.600 26.465 174.915 ;
        RECT 27.255 174.895 27.545 174.940 ;
        RECT 30.835 174.895 31.125 174.940 ;
        RECT 32.670 174.895 32.960 174.940 ;
        RECT 27.255 174.755 32.960 174.895 ;
        RECT 27.255 174.710 27.545 174.755 ;
        RECT 30.835 174.710 31.125 174.755 ;
        RECT 32.670 174.710 32.960 174.755 ;
        RECT 33.135 174.710 33.425 174.940 ;
        RECT 34.515 174.710 34.805 174.940 ;
        RECT 35.435 174.710 35.725 174.940 ;
        RECT 25.875 174.555 26.465 174.600 ;
        RECT 29.115 174.555 29.765 174.600 ;
        RECT 25.300 174.415 29.765 174.555 ;
        RECT 25.300 174.355 25.620 174.415 ;
        RECT 25.875 174.370 26.165 174.415 ;
        RECT 29.115 174.370 29.765 174.415 ;
        RECT 30.360 174.555 30.680 174.615 ;
        RECT 33.210 174.555 33.350 174.710 ;
        RECT 35.880 174.695 36.200 174.955 ;
        RECT 36.355 174.895 36.645 174.940 ;
        RECT 36.355 174.755 38.870 174.895 ;
        RECT 36.355 174.710 36.645 174.755 ;
        RECT 38.730 174.615 38.870 174.755 ;
        RECT 39.100 174.695 39.420 174.955 ;
        RECT 40.110 174.940 40.250 175.775 ;
        RECT 43.240 175.715 43.560 175.775 ;
        RECT 44.710 175.775 60.490 175.915 ;
        RECT 40.940 175.375 41.260 175.635 ;
        RECT 41.030 175.235 41.170 175.375 ;
        RECT 44.710 175.235 44.850 175.775 ;
        RECT 52.440 175.375 52.760 175.635 ;
        RECT 54.755 175.390 55.045 175.620 ;
        RECT 60.350 175.575 60.490 175.775 ;
        RECT 61.270 175.775 75.670 175.915 ;
        RECT 61.270 175.575 61.410 175.775 ;
        RECT 68.080 175.715 68.400 175.775 ;
        RECT 71.760 175.715 72.080 175.775 ;
        RECT 60.350 175.435 61.410 175.575 ;
        RECT 64.860 175.575 65.180 175.635 ;
        RECT 71.300 175.575 71.620 175.635 ;
        RECT 64.860 175.435 75.210 175.575 ;
        RECT 51.995 175.235 52.285 175.280 ;
        RECT 52.530 175.235 52.670 175.375 ;
        RECT 40.570 175.095 44.850 175.235 ;
        RECT 40.570 174.940 40.710 175.095 ;
        RECT 40.035 174.710 40.325 174.940 ;
        RECT 40.495 174.710 40.785 174.940 ;
        RECT 40.955 174.895 41.245 174.940 ;
        RECT 44.160 174.895 44.480 174.955 ;
        RECT 44.710 174.940 44.850 175.095 ;
        RECT 45.170 175.095 47.150 175.235 ;
        RECT 45.170 174.940 45.310 175.095 ;
        RECT 47.010 174.955 47.150 175.095 ;
        RECT 51.995 175.095 52.670 175.235 ;
        RECT 51.995 175.050 52.285 175.095 ;
        RECT 52.900 175.035 53.220 175.295 ;
        RECT 54.830 175.235 54.970 175.390 ;
        RECT 64.860 175.375 65.180 175.435 ;
        RECT 54.830 175.095 56.810 175.235 ;
        RECT 40.955 174.755 44.480 174.895 ;
        RECT 40.955 174.710 41.245 174.755 ;
        RECT 30.360 174.415 33.350 174.555 ;
        RECT 38.640 174.555 38.960 174.615 ;
        RECT 41.030 174.555 41.170 174.710 ;
        RECT 44.160 174.695 44.480 174.755 ;
        RECT 44.635 174.710 44.925 174.940 ;
        RECT 45.095 174.710 45.385 174.940 ;
        RECT 46.015 174.710 46.305 174.940 ;
        RECT 46.090 174.555 46.230 174.710 ;
        RECT 46.920 174.695 47.240 174.955 ;
        RECT 48.760 174.895 49.080 174.955 ;
        RECT 49.695 174.895 49.985 174.940 ;
        RECT 52.455 174.895 52.745 174.940 ;
        RECT 48.760 174.755 52.745 174.895 ;
        RECT 52.990 174.895 53.130 175.035 ;
        RECT 56.120 174.895 56.440 174.955 ;
        RECT 56.670 174.940 56.810 175.095 ;
        RECT 52.990 174.755 56.440 174.895 ;
        RECT 48.760 174.695 49.080 174.755 ;
        RECT 49.695 174.710 49.985 174.755 ;
        RECT 52.455 174.710 52.745 174.755 ;
        RECT 56.120 174.695 56.440 174.755 ;
        RECT 56.595 174.710 56.885 174.940 ;
        RECT 61.640 174.695 61.960 174.955 ;
        RECT 63.480 174.895 63.800 174.955 ;
        RECT 64.400 174.895 64.720 174.955 ;
        RECT 67.710 174.940 67.850 175.435 ;
        RECT 71.300 175.375 71.620 175.435 ;
        RECT 72.680 175.235 73.000 175.295 ;
        RECT 73.600 175.235 73.920 175.295 ;
        RECT 72.680 175.095 73.920 175.235 ;
        RECT 72.680 175.035 73.000 175.095 ;
        RECT 73.600 175.035 73.920 175.095 ;
        RECT 63.480 174.755 64.720 174.895 ;
        RECT 63.480 174.695 63.800 174.755 ;
        RECT 64.400 174.695 64.720 174.755 ;
        RECT 67.635 174.710 67.925 174.940 ;
        RECT 68.080 174.695 68.400 174.955 ;
        RECT 68.540 174.695 68.860 174.955 ;
        RECT 69.475 174.710 69.765 174.940 ;
        RECT 38.640 174.415 41.170 174.555 ;
        RECT 41.490 174.415 46.230 174.555 ;
        RECT 30.360 174.355 30.680 174.415 ;
        RECT 38.640 174.355 38.960 174.415 ;
        RECT 15.180 174.015 15.500 174.275 ;
        RECT 24.380 174.215 24.700 174.275 ;
        RECT 34.500 174.215 34.820 174.275 ;
        RECT 24.380 174.075 34.820 174.215 ;
        RECT 24.380 174.015 24.700 174.075 ;
        RECT 34.500 174.015 34.820 174.075 ;
        RECT 37.720 174.015 38.040 174.275 ;
        RECT 39.100 174.215 39.420 174.275 ;
        RECT 40.020 174.215 40.340 174.275 ;
        RECT 41.490 174.215 41.630 174.415 ;
        RECT 39.100 174.075 41.630 174.215 ;
        RECT 39.100 174.015 39.420 174.075 ;
        RECT 40.020 174.015 40.340 174.075 ;
        RECT 42.320 174.015 42.640 174.275 ;
        RECT 42.795 174.215 43.085 174.260 ;
        RECT 44.620 174.215 44.940 174.275 ;
        RECT 42.795 174.075 44.940 174.215 ;
        RECT 46.090 174.215 46.230 174.415 ;
        RECT 46.460 174.555 46.780 174.615 ;
        RECT 52.915 174.555 53.205 174.600 ;
        RECT 69.550 174.555 69.690 174.710 ;
        RECT 71.300 174.695 71.620 174.955 ;
        RECT 71.760 174.695 72.080 174.955 ;
        RECT 72.220 174.695 72.540 174.955 ;
        RECT 75.070 174.940 75.210 175.435 ;
        RECT 75.530 174.940 75.670 175.775 ;
        RECT 83.260 175.775 84.945 175.915 ;
        RECT 83.260 175.715 83.580 175.775 ;
        RECT 84.655 175.730 84.945 175.775 ;
        RECT 89.240 175.715 89.560 175.975 ;
        RECT 98.440 175.915 98.760 175.975 ;
        RECT 107.180 175.915 107.500 175.975 ;
        RECT 98.440 175.775 107.500 175.915 ;
        RECT 98.440 175.715 98.760 175.775 ;
        RECT 107.180 175.715 107.500 175.775 ;
        RECT 108.100 175.715 108.420 175.975 ;
        RECT 83.720 175.575 84.040 175.635 ;
        RECT 97.980 175.575 98.300 175.635 ;
        RECT 83.720 175.435 98.300 175.575 ;
        RECT 83.720 175.375 84.040 175.435 ;
        RECT 79.120 175.235 79.440 175.295 ;
        RECT 93.840 175.235 94.160 175.295 ;
        RECT 79.120 175.095 94.160 175.235 ;
        RECT 79.120 175.035 79.440 175.095 ;
        RECT 73.155 174.710 73.445 174.940 ;
        RECT 74.995 174.710 75.285 174.940 ;
        RECT 75.455 174.710 75.745 174.940 ;
        RECT 73.230 174.555 73.370 174.710 ;
        RECT 75.900 174.695 76.220 174.955 ;
        RECT 76.835 174.710 77.125 174.940 ;
        RECT 86.480 174.895 86.800 174.955 ;
        RECT 91.630 174.940 91.770 175.095 ;
        RECT 93.840 175.035 94.160 175.095 ;
        RECT 88.335 174.895 88.625 174.940 ;
        RECT 86.480 174.755 88.625 174.895 ;
        RECT 74.060 174.555 74.380 174.615 ;
        RECT 76.910 174.555 77.050 174.710 ;
        RECT 86.480 174.695 86.800 174.755 ;
        RECT 88.335 174.710 88.625 174.755 ;
        RECT 91.555 174.710 91.845 174.940 ;
        RECT 92.015 174.710 92.305 174.940 ;
        RECT 92.475 174.895 92.765 174.940 ;
        RECT 92.920 174.895 93.240 174.955 ;
        RECT 92.475 174.755 93.240 174.895 ;
        RECT 92.475 174.710 92.765 174.755 ;
        RECT 46.460 174.415 53.205 174.555 ;
        RECT 46.460 174.355 46.780 174.415 ;
        RECT 52.915 174.370 53.205 174.415 ;
        RECT 53.450 174.415 60.950 174.555 ;
        RECT 51.980 174.215 52.300 174.275 ;
        RECT 46.090 174.075 52.300 174.215 ;
        RECT 42.795 174.030 43.085 174.075 ;
        RECT 44.620 174.015 44.940 174.075 ;
        RECT 51.980 174.015 52.300 174.075 ;
        RECT 52.440 174.215 52.760 174.275 ;
        RECT 53.450 174.215 53.590 174.415 ;
        RECT 52.440 174.075 53.590 174.215 ;
        RECT 52.440 174.015 52.760 174.075 ;
        RECT 55.660 174.015 55.980 174.275 ;
        RECT 57.500 174.015 57.820 174.275 ;
        RECT 60.810 174.260 60.950 174.415 ;
        RECT 62.650 174.415 77.050 174.555 ;
        RECT 62.650 174.275 62.790 174.415 ;
        RECT 74.060 174.355 74.380 174.415 ;
        RECT 78.200 174.355 78.520 174.615 ;
        RECT 81.420 174.555 81.740 174.615 ;
        RECT 92.090 174.555 92.230 174.710 ;
        RECT 92.920 174.695 93.240 174.755 ;
        RECT 93.395 174.895 93.685 174.940 ;
        RECT 94.390 174.895 94.530 175.435 ;
        RECT 97.980 175.375 98.300 175.435 ;
        RECT 104.435 175.575 104.725 175.620 ;
        RECT 105.340 175.575 105.660 175.635 ;
        RECT 104.435 175.435 105.660 175.575 ;
        RECT 104.435 175.390 104.725 175.435 ;
        RECT 105.340 175.375 105.660 175.435 ;
        RECT 100.740 175.235 101.060 175.295 ;
        RECT 95.770 175.095 101.060 175.235 ;
        RECT 95.770 174.940 95.910 175.095 ;
        RECT 100.740 175.035 101.060 175.095 ;
        RECT 94.775 174.895 95.065 174.940 ;
        RECT 93.395 174.755 95.065 174.895 ;
        RECT 93.395 174.710 93.685 174.755 ;
        RECT 94.775 174.710 95.065 174.755 ;
        RECT 95.695 174.710 95.985 174.940 ;
        RECT 96.140 174.695 96.460 174.955 ;
        RECT 96.615 174.895 96.905 174.940 ;
        RECT 99.820 174.895 100.140 174.955 ;
        RECT 96.615 174.755 100.140 174.895 ;
        RECT 96.615 174.710 96.905 174.755 ;
        RECT 96.230 174.555 96.370 174.695 ;
        RECT 81.420 174.415 96.370 174.555 ;
        RECT 81.420 174.355 81.740 174.415 ;
        RECT 60.735 174.215 61.025 174.260 ;
        RECT 61.640 174.215 61.960 174.275 ;
        RECT 60.735 174.075 61.960 174.215 ;
        RECT 60.735 174.030 61.025 174.075 ;
        RECT 61.640 174.015 61.960 174.075 ;
        RECT 62.560 174.015 62.880 174.275 ;
        RECT 64.400 174.215 64.720 174.275 ;
        RECT 66.255 174.215 66.545 174.260 ;
        RECT 64.400 174.075 66.545 174.215 ;
        RECT 64.400 174.015 64.720 174.075 ;
        RECT 66.255 174.030 66.545 174.075 ;
        RECT 69.460 174.215 69.780 174.275 ;
        RECT 69.935 174.215 70.225 174.260 ;
        RECT 69.460 174.075 70.225 174.215 ;
        RECT 69.460 174.015 69.780 174.075 ;
        RECT 69.935 174.030 70.225 174.075 ;
        RECT 72.220 174.215 72.540 174.275 ;
        RECT 73.615 174.215 73.905 174.260 ;
        RECT 72.220 174.075 73.905 174.215 ;
        RECT 72.220 174.015 72.540 174.075 ;
        RECT 73.615 174.030 73.905 174.075 ;
        RECT 90.175 174.215 90.465 174.260 ;
        RECT 90.620 174.215 90.940 174.275 ;
        RECT 90.175 174.075 90.940 174.215 ;
        RECT 90.175 174.030 90.465 174.075 ;
        RECT 90.620 174.015 90.940 174.075 ;
        RECT 93.840 174.215 94.160 174.275 ;
        RECT 96.690 174.215 96.830 174.710 ;
        RECT 99.820 174.695 100.140 174.755 ;
        RECT 101.675 174.895 101.965 174.940 ;
        RECT 103.960 174.895 104.280 174.955 ;
        RECT 101.675 174.755 104.280 174.895 ;
        RECT 101.675 174.710 101.965 174.755 ;
        RECT 103.960 174.695 104.280 174.755 ;
        RECT 105.800 174.940 106.120 174.955 ;
        RECT 105.800 174.710 106.335 174.940 ;
        RECT 106.720 174.880 107.040 174.955 ;
        RECT 108.190 174.940 108.330 175.715 ;
        RECT 108.560 175.575 108.880 175.635 ;
        RECT 111.795 175.575 112.085 175.620 ;
        RECT 108.560 175.435 112.085 175.575 ;
        RECT 108.560 175.375 108.880 175.435 ;
        RECT 111.795 175.390 112.085 175.435 ;
        RECT 109.020 175.235 109.340 175.295 ;
        RECT 109.020 175.095 110.170 175.235 ;
        RECT 109.020 175.035 109.340 175.095 ;
        RECT 106.540 174.740 107.040 174.880 ;
        RECT 105.800 174.695 106.120 174.710 ;
        RECT 106.720 174.695 107.040 174.740 ;
        RECT 107.180 174.680 107.500 174.940 ;
        RECT 108.115 174.895 108.405 174.940 ;
        RECT 108.575 174.895 108.865 174.940 ;
        RECT 108.115 174.755 108.865 174.895 ;
        RECT 108.115 174.710 108.405 174.755 ;
        RECT 108.575 174.710 108.865 174.755 ;
        RECT 109.480 174.695 109.800 174.955 ;
        RECT 110.030 174.940 110.170 175.095 ;
        RECT 109.955 174.710 110.245 174.940 ;
        RECT 110.400 174.695 110.720 174.955 ;
        RECT 111.780 174.895 112.100 174.955 ;
        RECT 113.175 174.895 113.465 174.940 ;
        RECT 111.780 174.755 113.465 174.895 ;
        RECT 111.780 174.695 112.100 174.755 ;
        RECT 113.175 174.710 113.465 174.755 ;
        RECT 97.995 174.555 98.285 174.600 ;
        RECT 100.740 174.555 101.060 174.615 ;
        RECT 97.995 174.415 101.060 174.555 ;
        RECT 135.635 174.550 136.775 223.880 ;
        RECT 138.130 223.810 139.580 225.110 ;
        RECT 143.180 223.840 144.630 225.140 ;
        RECT 97.995 174.370 98.285 174.415 ;
        RECT 100.740 174.355 101.060 174.415 ;
        RECT 93.840 174.075 96.830 174.215 ;
        RECT 93.840 174.015 94.160 174.075 ;
        RECT 104.880 174.015 105.200 174.275 ;
        RECT 112.240 174.015 112.560 174.275 ;
        RECT 10.510 173.395 115.850 173.875 ;
        RECT 135.580 173.430 136.830 174.550 ;
        RECT 135.635 173.420 136.775 173.430 ;
        RECT 20.240 173.195 20.560 173.255 ;
        RECT 20.715 173.195 21.005 173.240 ;
        RECT 20.240 173.055 21.005 173.195 ;
        RECT 20.240 172.995 20.560 173.055 ;
        RECT 20.715 173.010 21.005 173.055 ;
        RECT 22.540 173.195 22.860 173.255 ;
        RECT 27.155 173.195 27.445 173.240 ;
        RECT 22.540 173.055 27.445 173.195 ;
        RECT 22.540 172.995 22.860 173.055 ;
        RECT 27.155 173.010 27.445 173.055 ;
        RECT 28.060 172.995 28.380 173.255 ;
        RECT 29.440 173.195 29.760 173.255 ;
        RECT 35.880 173.195 36.200 173.255 ;
        RECT 29.440 173.055 36.200 173.195 ;
        RECT 29.440 172.995 29.760 173.055 ;
        RECT 35.880 172.995 36.200 173.055 ;
        RECT 46.920 173.195 47.240 173.255 ;
        RECT 51.535 173.195 51.825 173.240 ;
        RECT 46.920 173.055 51.825 173.195 ;
        RECT 46.920 172.995 47.240 173.055 ;
        RECT 51.535 173.010 51.825 173.055 ;
        RECT 51.980 173.195 52.300 173.255 ;
        RECT 62.560 173.195 62.880 173.255 ;
        RECT 81.420 173.195 81.740 173.255 ;
        RECT 51.980 173.055 62.880 173.195 ;
        RECT 51.980 172.995 52.300 173.055 ;
        RECT 62.560 172.995 62.880 173.055 ;
        RECT 63.110 173.055 81.740 173.195 ;
        RECT 21.635 172.855 21.925 172.900 ;
        RECT 23.460 172.855 23.780 172.915 ;
        RECT 21.635 172.715 23.780 172.855 ;
        RECT 21.635 172.670 21.925 172.715 ;
        RECT 23.460 172.655 23.780 172.715 ;
        RECT 19.320 172.515 19.640 172.575 ;
        RECT 21.175 172.515 21.465 172.560 ;
        RECT 22.540 172.515 22.860 172.575 ;
        RECT 19.320 172.375 22.860 172.515 ;
        RECT 19.320 172.315 19.640 172.375 ;
        RECT 21.175 172.330 21.465 172.375 ;
        RECT 22.540 172.315 22.860 172.375 ;
        RECT 24.380 172.315 24.700 172.575 ;
        RECT 28.150 172.560 28.290 172.995 ;
        RECT 29.530 172.855 29.670 172.995 ;
        RECT 53.015 172.855 53.305 172.900 ;
        RECT 55.660 172.855 55.980 172.915 ;
        RECT 56.255 172.855 56.905 172.900 ;
        RECT 29.070 172.715 29.670 172.855 ;
        RECT 49.770 172.715 52.670 172.855 ;
        RECT 29.070 172.560 29.210 172.715 ;
        RECT 28.075 172.330 28.365 172.560 ;
        RECT 28.995 172.330 29.285 172.560 ;
        RECT 29.915 172.330 30.205 172.560 ;
        RECT 15.180 171.495 15.500 171.555 ;
        RECT 29.990 171.495 30.130 172.330 ;
        RECT 30.360 172.315 30.680 172.575 ;
        RECT 30.835 172.515 31.125 172.560 ;
        RECT 31.280 172.515 31.600 172.575 ;
        RECT 34.055 172.515 34.345 172.560 ;
        RECT 30.835 172.375 34.345 172.515 ;
        RECT 30.835 172.330 31.125 172.375 ;
        RECT 31.280 172.315 31.600 172.375 ;
        RECT 34.055 172.330 34.345 172.375 ;
        RECT 34.515 172.330 34.805 172.560 ;
        RECT 30.450 172.175 30.590 172.315 ;
        RECT 33.580 172.175 33.900 172.235 ;
        RECT 34.590 172.175 34.730 172.330 ;
        RECT 34.960 172.315 35.280 172.575 ;
        RECT 35.880 172.315 36.200 172.575 ;
        RECT 38.640 172.515 38.960 172.575 ;
        RECT 39.115 172.515 39.405 172.560 ;
        RECT 38.640 172.375 39.405 172.515 ;
        RECT 38.640 172.315 38.960 172.375 ;
        RECT 39.115 172.330 39.405 172.375 ;
        RECT 39.560 172.315 39.880 172.575 ;
        RECT 40.020 172.315 40.340 172.575 ;
        RECT 40.955 172.515 41.245 172.560 ;
        RECT 49.770 172.515 49.910 172.715 ;
        RECT 40.955 172.375 49.910 172.515 ;
        RECT 40.955 172.330 41.245 172.375 ;
        RECT 50.140 172.315 50.460 172.575 ;
        RECT 52.530 172.515 52.670 172.715 ;
        RECT 53.015 172.715 56.905 172.855 ;
        RECT 53.015 172.670 53.605 172.715 ;
        RECT 52.530 172.375 53.130 172.515 ;
        RECT 52.440 172.175 52.760 172.235 ;
        RECT 30.450 172.035 52.760 172.175 ;
        RECT 33.580 171.975 33.900 172.035 ;
        RECT 52.440 171.975 52.760 172.035 ;
        RECT 15.180 171.355 30.130 171.495 ;
        RECT 31.740 171.495 32.060 171.555 ;
        RECT 32.215 171.495 32.505 171.540 ;
        RECT 31.740 171.355 32.505 171.495 ;
        RECT 15.180 171.295 15.500 171.355 ;
        RECT 31.740 171.295 32.060 171.355 ;
        RECT 32.215 171.310 32.505 171.355 ;
        RECT 32.660 171.295 32.980 171.555 ;
        RECT 34.040 171.495 34.360 171.555 ;
        RECT 37.735 171.495 38.025 171.540 ;
        RECT 34.040 171.355 38.025 171.495 ;
        RECT 34.040 171.295 34.360 171.355 ;
        RECT 37.735 171.310 38.025 171.355 ;
        RECT 43.715 171.495 44.005 171.540 ;
        RECT 46.460 171.495 46.780 171.555 ;
        RECT 43.715 171.355 46.780 171.495 ;
        RECT 52.990 171.495 53.130 172.375 ;
        RECT 53.315 172.355 53.605 172.670 ;
        RECT 55.660 172.655 55.980 172.715 ;
        RECT 56.255 172.670 56.905 172.715 ;
        RECT 57.500 172.855 57.820 172.915 ;
        RECT 58.895 172.855 59.185 172.900 ;
        RECT 57.500 172.715 59.185 172.855 ;
        RECT 57.500 172.655 57.820 172.715 ;
        RECT 58.895 172.670 59.185 172.715 ;
        RECT 61.640 172.855 61.960 172.915 ;
        RECT 63.110 172.855 63.250 173.055 ;
        RECT 81.420 172.995 81.740 173.055 ;
        RECT 81.895 173.195 82.185 173.240 ;
        RECT 99.835 173.195 100.125 173.240 ;
        RECT 105.340 173.195 105.660 173.255 ;
        RECT 81.895 173.055 86.250 173.195 ;
        RECT 81.895 173.010 82.185 173.055 ;
        RECT 61.640 172.715 63.250 172.855 ;
        RECT 71.760 172.855 72.080 172.915 ;
        RECT 86.110 172.855 86.250 173.055 ;
        RECT 99.835 173.055 105.660 173.195 ;
        RECT 99.835 173.010 100.125 173.055 ;
        RECT 105.340 172.995 105.660 173.055 ;
        RECT 86.475 172.855 87.125 172.900 ;
        RECT 90.075 172.855 90.365 172.900 ;
        RECT 71.760 172.715 72.910 172.855 ;
        RECT 86.110 172.715 90.365 172.855 ;
        RECT 61.640 172.655 61.960 172.715 ;
        RECT 71.760 172.655 72.080 172.715 ;
        RECT 54.395 172.515 54.685 172.560 ;
        RECT 57.975 172.515 58.265 172.560 ;
        RECT 59.810 172.515 60.100 172.560 ;
        RECT 54.395 172.375 60.100 172.515 ;
        RECT 54.395 172.330 54.685 172.375 ;
        RECT 57.975 172.330 58.265 172.375 ;
        RECT 59.810 172.330 60.100 172.375 ;
        RECT 71.300 172.515 71.620 172.575 ;
        RECT 72.770 172.560 72.910 172.715 ;
        RECT 86.475 172.670 87.125 172.715 ;
        RECT 89.775 172.670 90.365 172.715 ;
        RECT 103.515 172.855 103.805 172.900 ;
        RECT 105.915 172.855 106.205 172.900 ;
        RECT 109.155 172.855 109.805 172.900 ;
        RECT 103.515 172.715 109.805 172.855 ;
        RECT 103.515 172.670 103.805 172.715 ;
        RECT 105.915 172.670 106.505 172.715 ;
        RECT 109.155 172.670 109.805 172.715 ;
        RECT 111.795 172.855 112.085 172.900 ;
        RECT 112.240 172.855 112.560 172.915 ;
        RECT 111.795 172.715 112.560 172.855 ;
        RECT 111.795 172.670 112.085 172.715 ;
        RECT 72.235 172.515 72.525 172.560 ;
        RECT 71.300 172.375 72.525 172.515 ;
        RECT 71.300 172.315 71.620 172.375 ;
        RECT 72.235 172.330 72.525 172.375 ;
        RECT 72.695 172.330 72.985 172.560 ;
        RECT 73.140 172.315 73.460 172.575 ;
        RECT 74.060 172.315 74.380 172.575 ;
        RECT 81.435 172.515 81.725 172.560 ;
        RECT 81.880 172.515 82.200 172.575 ;
        RECT 81.435 172.375 82.200 172.515 ;
        RECT 81.435 172.330 81.725 172.375 ;
        RECT 81.880 172.315 82.200 172.375 ;
        RECT 82.800 172.315 83.120 172.575 ;
        RECT 83.280 172.515 83.570 172.560 ;
        RECT 85.115 172.515 85.405 172.560 ;
        RECT 88.695 172.515 88.985 172.560 ;
        RECT 83.280 172.375 88.985 172.515 ;
        RECT 83.280 172.330 83.570 172.375 ;
        RECT 85.115 172.330 85.405 172.375 ;
        RECT 88.695 172.330 88.985 172.375 ;
        RECT 89.775 172.355 90.065 172.670 ;
        RECT 100.295 172.330 100.585 172.560 ;
        RECT 53.820 172.175 54.140 172.235 ;
        RECT 56.120 172.175 56.440 172.235 ;
        RECT 60.275 172.175 60.565 172.220 ;
        RECT 53.820 172.035 60.565 172.175 ;
        RECT 53.820 171.975 54.140 172.035 ;
        RECT 56.120 171.975 56.440 172.035 ;
        RECT 60.275 171.990 60.565 172.035 ;
        RECT 84.180 171.975 84.500 172.235 ;
        RECT 91.555 172.175 91.845 172.220 ;
        RECT 95.235 172.175 95.525 172.220 ;
        RECT 97.060 172.175 97.380 172.235 ;
        RECT 91.555 172.035 97.380 172.175 ;
        RECT 91.555 171.990 91.845 172.035 ;
        RECT 95.235 171.990 95.525 172.035 ;
        RECT 97.060 171.975 97.380 172.035 ;
        RECT 98.440 172.175 98.760 172.235 ;
        RECT 98.915 172.175 99.205 172.220 ;
        RECT 98.440 172.035 99.205 172.175 ;
        RECT 98.440 171.975 98.760 172.035 ;
        RECT 98.915 171.990 99.205 172.035 ;
        RECT 54.395 171.835 54.685 171.880 ;
        RECT 57.515 171.835 57.805 171.880 ;
        RECT 59.405 171.835 59.695 171.880 ;
        RECT 54.395 171.695 59.695 171.835 ;
        RECT 54.395 171.650 54.685 171.695 ;
        RECT 57.515 171.650 57.805 171.695 ;
        RECT 59.405 171.650 59.695 171.695 ;
        RECT 83.685 171.835 83.975 171.880 ;
        RECT 85.575 171.835 85.865 171.880 ;
        RECT 88.695 171.835 88.985 171.880 ;
        RECT 100.370 171.835 100.510 172.330 ;
        RECT 103.040 172.315 103.360 172.575 ;
        RECT 106.215 172.355 106.505 172.670 ;
        RECT 112.240 172.655 112.560 172.715 ;
        RECT 107.295 172.515 107.585 172.560 ;
        RECT 110.875 172.515 111.165 172.560 ;
        RECT 112.710 172.515 113.000 172.560 ;
        RECT 107.295 172.375 113.000 172.515 ;
        RECT 107.295 172.330 107.585 172.375 ;
        RECT 110.875 172.330 111.165 172.375 ;
        RECT 112.710 172.330 113.000 172.375 ;
        RECT 111.780 172.175 112.100 172.235 ;
        RECT 102.210 172.035 112.100 172.175 ;
        RECT 102.210 171.880 102.350 172.035 ;
        RECT 111.780 171.975 112.100 172.035 ;
        RECT 113.175 172.175 113.465 172.220 ;
        RECT 113.620 172.175 113.940 172.235 ;
        RECT 113.175 172.035 113.940 172.175 ;
        RECT 113.175 171.990 113.465 172.035 ;
        RECT 113.620 171.975 113.940 172.035 ;
        RECT 133.700 172.190 134.930 172.680 ;
        RECT 133.700 171.930 136.690 172.190 ;
        RECT 138.330 171.930 139.470 223.810 ;
        RECT 83.685 171.695 88.985 171.835 ;
        RECT 83.685 171.650 83.975 171.695 ;
        RECT 85.575 171.650 85.865 171.695 ;
        RECT 88.695 171.650 88.985 171.695 ;
        RECT 92.090 171.695 100.510 171.835 ;
        RECT 55.200 171.495 55.520 171.555 ;
        RECT 52.990 171.355 55.520 171.495 ;
        RECT 43.715 171.310 44.005 171.355 ;
        RECT 46.460 171.295 46.780 171.355 ;
        RECT 55.200 171.295 55.520 171.355 ;
        RECT 70.855 171.495 71.145 171.540 ;
        RECT 71.300 171.495 71.620 171.555 ;
        RECT 70.855 171.355 71.620 171.495 ;
        RECT 70.855 171.310 71.145 171.355 ;
        RECT 71.300 171.295 71.620 171.355 ;
        RECT 84.640 171.495 84.960 171.555 ;
        RECT 92.090 171.540 92.230 171.695 ;
        RECT 102.135 171.650 102.425 171.880 ;
        RECT 107.295 171.835 107.585 171.880 ;
        RECT 110.415 171.835 110.705 171.880 ;
        RECT 112.305 171.835 112.595 171.880 ;
        RECT 107.295 171.695 112.595 171.835 ;
        RECT 107.295 171.650 107.585 171.695 ;
        RECT 110.415 171.650 110.705 171.695 ;
        RECT 112.305 171.650 112.595 171.695 ;
        RECT 92.015 171.495 92.305 171.540 ;
        RECT 84.640 171.355 92.305 171.495 ;
        RECT 84.640 171.295 84.960 171.355 ;
        RECT 92.015 171.310 92.305 171.355 ;
        RECT 104.420 171.295 104.740 171.555 ;
        RECT 10.510 170.675 115.850 171.155 ;
        RECT 133.700 170.790 139.470 171.930 ;
        RECT 133.700 170.600 136.690 170.790 ;
        RECT 23.935 170.475 24.225 170.520 ;
        RECT 24.840 170.475 25.160 170.535 ;
        RECT 23.935 170.335 25.160 170.475 ;
        RECT 23.935 170.290 24.225 170.335 ;
        RECT 24.840 170.275 25.160 170.335 ;
        RECT 34.500 170.475 34.820 170.535 ;
        RECT 35.880 170.475 36.200 170.535 ;
        RECT 60.735 170.475 61.025 170.520 ;
        RECT 83.720 170.475 84.040 170.535 ;
        RECT 34.500 170.335 84.040 170.475 ;
        RECT 34.500 170.275 34.820 170.335 ;
        RECT 35.880 170.275 36.200 170.335 ;
        RECT 60.735 170.290 61.025 170.335 ;
        RECT 83.720 170.275 84.040 170.335 ;
        RECT 84.180 170.475 84.500 170.535 ;
        RECT 87.875 170.475 88.165 170.520 ;
        RECT 84.180 170.335 88.165 170.475 ;
        RECT 84.180 170.275 84.500 170.335 ;
        RECT 87.875 170.290 88.165 170.335 ;
        RECT 22.080 170.135 22.400 170.195 ;
        RECT 40.020 170.135 40.340 170.195 ;
        RECT 22.080 169.995 40.340 170.135 ;
        RECT 22.080 169.935 22.400 169.995 ;
        RECT 40.020 169.935 40.340 169.995 ;
        RECT 50.255 170.135 50.545 170.180 ;
        RECT 53.375 170.135 53.665 170.180 ;
        RECT 55.265 170.135 55.555 170.180 ;
        RECT 50.255 169.995 55.555 170.135 ;
        RECT 50.255 169.950 50.545 169.995 ;
        RECT 53.375 169.950 53.665 169.995 ;
        RECT 55.265 169.950 55.555 169.995 ;
        RECT 74.950 170.135 75.240 170.180 ;
        RECT 77.730 170.135 78.020 170.180 ;
        RECT 79.590 170.135 79.880 170.180 ;
        RECT 74.950 169.995 79.880 170.135 ;
        RECT 74.950 169.950 75.240 169.995 ;
        RECT 77.730 169.950 78.020 169.995 ;
        RECT 79.590 169.950 79.880 169.995 ;
        RECT 86.955 169.950 87.245 170.180 ;
        RECT 133.700 170.120 134.930 170.600 ;
        RECT 45.095 169.795 45.385 169.840 ;
        RECT 47.380 169.795 47.700 169.855 ;
        RECT 45.095 169.655 47.700 169.795 ;
        RECT 45.095 169.610 45.385 169.655 ;
        RECT 47.380 169.595 47.700 169.655 ;
        RECT 56.120 169.595 56.440 169.855 ;
        RECT 67.620 169.795 67.940 169.855 ;
        RECT 71.085 169.795 71.375 169.840 ;
        RECT 80.055 169.795 80.345 169.840 ;
        RECT 83.260 169.795 83.580 169.855 ;
        RECT 67.620 169.655 78.890 169.795 ;
        RECT 67.620 169.595 67.940 169.655 ;
        RECT 71.085 169.610 71.375 169.655 ;
        RECT 30.360 169.255 30.680 169.515 ;
        RECT 32.675 169.455 32.965 169.500 ;
        RECT 36.355 169.455 36.645 169.500 ;
        RECT 38.180 169.455 38.500 169.515 ;
        RECT 30.910 169.315 38.500 169.455 ;
        RECT 22.540 169.115 22.860 169.175 ;
        RECT 30.910 169.115 31.050 169.315 ;
        RECT 32.675 169.270 32.965 169.315 ;
        RECT 36.355 169.270 36.645 169.315 ;
        RECT 38.180 169.255 38.500 169.315 ;
        RECT 46.935 169.270 47.225 169.500 ;
        RECT 22.540 168.975 31.050 169.115 ;
        RECT 31.280 169.115 31.600 169.175 ;
        RECT 32.215 169.115 32.505 169.160 ;
        RECT 31.280 168.975 32.505 169.115 ;
        RECT 22.540 168.915 22.860 168.975 ;
        RECT 31.280 168.915 31.600 168.975 ;
        RECT 32.215 168.930 32.505 168.975 ;
        RECT 36.815 169.115 37.105 169.160 ;
        RECT 38.640 169.115 38.960 169.175 ;
        RECT 36.815 168.975 38.960 169.115 ;
        RECT 36.815 168.930 37.105 168.975 ;
        RECT 38.640 168.915 38.960 168.975 ;
        RECT 41.875 168.775 42.165 168.820 ;
        RECT 43.700 168.775 44.020 168.835 ;
        RECT 41.875 168.635 44.020 168.775 ;
        RECT 41.875 168.590 42.165 168.635 ;
        RECT 43.700 168.575 44.020 168.635 ;
        RECT 46.460 168.775 46.780 168.835 ;
        RECT 47.010 168.775 47.150 169.270 ;
        RECT 49.175 169.160 49.465 169.475 ;
        RECT 50.255 169.455 50.545 169.500 ;
        RECT 53.835 169.455 54.125 169.500 ;
        RECT 55.670 169.455 55.960 169.500 ;
        RECT 50.255 169.315 55.960 169.455 ;
        RECT 50.255 169.270 50.545 169.315 ;
        RECT 53.835 169.270 54.125 169.315 ;
        RECT 55.670 169.270 55.960 169.315 ;
        RECT 61.655 169.455 61.945 169.500 ;
        RECT 63.480 169.455 63.800 169.515 ;
        RECT 61.655 169.315 63.800 169.455 ;
        RECT 61.655 169.270 61.945 169.315 ;
        RECT 63.480 169.255 63.800 169.315 ;
        RECT 74.950 169.455 75.240 169.500 ;
        RECT 74.950 169.315 77.485 169.455 ;
        RECT 74.950 169.270 75.240 169.315 ;
        RECT 48.875 169.115 49.465 169.160 ;
        RECT 49.680 169.115 50.000 169.175 ;
        RECT 52.115 169.115 52.765 169.160 ;
        RECT 48.875 168.975 52.765 169.115 ;
        RECT 48.875 168.930 49.165 168.975 ;
        RECT 49.680 168.915 50.000 168.975 ;
        RECT 52.115 168.930 52.765 168.975 ;
        RECT 54.740 168.915 55.060 169.175 ;
        RECT 55.200 169.115 55.520 169.175 ;
        RECT 57.500 169.115 57.820 169.175 ;
        RECT 73.090 169.115 73.380 169.160 ;
        RECT 75.440 169.115 75.760 169.175 ;
        RECT 77.270 169.160 77.485 169.315 ;
        RECT 78.200 169.255 78.520 169.515 ;
        RECT 78.750 169.455 78.890 169.655 ;
        RECT 80.055 169.655 83.580 169.795 ;
        RECT 80.055 169.610 80.345 169.655 ;
        RECT 83.260 169.595 83.580 169.655 ;
        RECT 84.180 169.595 84.500 169.855 ;
        RECT 84.640 169.595 84.960 169.855 ;
        RECT 87.030 169.795 87.170 169.950 ;
        RECT 91.080 169.795 91.400 169.855 ;
        RECT 103.500 169.795 103.820 169.855 ;
        RECT 87.030 169.655 89.010 169.795 ;
        RECT 88.870 169.500 89.010 169.655 ;
        RECT 91.080 169.655 103.820 169.795 ;
        RECT 91.080 169.595 91.400 169.655 ;
        RECT 93.010 169.500 93.150 169.655 ;
        RECT 103.500 169.595 103.820 169.655 ;
        RECT 85.115 169.455 85.405 169.500 ;
        RECT 78.750 169.315 85.405 169.455 ;
        RECT 85.115 169.270 85.405 169.315 ;
        RECT 88.795 169.270 89.085 169.500 ;
        RECT 92.935 169.270 93.225 169.500 ;
        RECT 94.315 169.270 94.605 169.500 ;
        RECT 76.350 169.115 76.640 169.160 ;
        RECT 55.200 168.975 62.790 169.115 ;
        RECT 55.200 168.915 55.520 168.975 ;
        RECT 57.500 168.915 57.820 168.975 ;
        RECT 56.120 168.775 56.440 168.835 ;
        RECT 62.650 168.820 62.790 168.975 ;
        RECT 73.090 168.975 76.640 169.115 ;
        RECT 73.090 168.930 73.380 168.975 ;
        RECT 75.440 168.915 75.760 168.975 ;
        RECT 76.350 168.930 76.640 168.975 ;
        RECT 77.270 169.115 77.560 169.160 ;
        RECT 79.130 169.115 79.420 169.160 ;
        RECT 77.270 168.975 79.420 169.115 ;
        RECT 77.270 168.930 77.560 168.975 ;
        RECT 79.130 168.930 79.420 168.975 ;
        RECT 93.380 168.915 93.700 169.175 ;
        RECT 46.460 168.635 56.440 168.775 ;
        RECT 46.460 168.575 46.780 168.635 ;
        RECT 56.120 168.575 56.440 168.635 ;
        RECT 62.575 168.590 62.865 168.820 ;
        RECT 86.940 168.775 87.260 168.835 ;
        RECT 94.390 168.775 94.530 169.270 ;
        RECT 97.980 169.255 98.300 169.515 ;
        RECT 100.740 169.455 101.060 169.515 ;
        RECT 105.800 169.455 106.120 169.515 ;
        RECT 100.740 169.315 106.120 169.455 ;
        RECT 100.740 169.255 101.060 169.315 ;
        RECT 105.800 169.255 106.120 169.315 ;
        RECT 108.560 169.455 108.880 169.515 ;
        RECT 109.955 169.455 110.245 169.500 ;
        RECT 108.560 169.315 110.245 169.455 ;
        RECT 108.560 169.255 108.880 169.315 ;
        RECT 109.955 169.270 110.245 169.315 ;
        RECT 110.875 169.455 111.165 169.500 ;
        RECT 115.920 169.455 116.240 169.515 ;
        RECT 110.875 169.315 116.240 169.455 ;
        RECT 110.875 169.270 111.165 169.315 ;
        RECT 115.920 169.255 116.240 169.315 ;
        RECT 97.535 169.115 97.825 169.160 ;
        RECT 100.280 169.115 100.600 169.175 ;
        RECT 107.640 169.115 107.960 169.175 ;
        RECT 109.480 169.160 109.800 169.175 ;
        RECT 109.385 169.115 109.800 169.160 ;
        RECT 97.535 168.975 100.600 169.115 ;
        RECT 97.535 168.930 97.825 168.975 ;
        RECT 100.280 168.915 100.600 168.975 ;
        RECT 104.510 168.975 109.800 169.115 ;
        RECT 99.820 168.775 100.140 168.835 ;
        RECT 86.940 168.635 100.140 168.775 ;
        RECT 86.940 168.575 87.260 168.635 ;
        RECT 99.820 168.575 100.140 168.635 ;
        RECT 101.200 168.775 101.520 168.835 ;
        RECT 104.510 168.820 104.650 168.975 ;
        RECT 107.640 168.915 107.960 168.975 ;
        RECT 109.385 168.930 109.800 168.975 ;
        RECT 109.480 168.915 109.800 168.930 ;
        RECT 104.435 168.775 104.725 168.820 ;
        RECT 101.200 168.635 104.725 168.775 ;
        RECT 101.200 168.575 101.520 168.635 ;
        RECT 104.435 168.590 104.725 168.635 ;
        RECT 10.510 167.955 115.850 168.435 ;
        RECT 38.180 167.755 38.500 167.815 ;
        RECT 49.680 167.755 50.000 167.815 ;
        RECT 50.155 167.755 50.445 167.800 ;
        RECT 38.180 167.615 43.470 167.755 ;
        RECT 38.180 167.555 38.500 167.615 ;
        RECT 23.460 167.415 23.780 167.475 ;
        RECT 29.915 167.415 30.205 167.460 ;
        RECT 38.640 167.415 38.960 167.475 ;
        RECT 39.215 167.415 39.505 167.460 ;
        RECT 42.455 167.415 43.105 167.460 ;
        RECT 20.790 167.275 22.770 167.415 ;
        RECT 20.790 167.120 20.930 167.275 ;
        RECT 22.630 167.135 22.770 167.275 ;
        RECT 23.460 167.275 35.190 167.415 ;
        RECT 23.460 167.215 23.780 167.275 ;
        RECT 29.915 167.230 30.205 167.275 ;
        RECT 20.715 166.890 21.005 167.120 ;
        RECT 21.175 167.075 21.465 167.120 ;
        RECT 22.080 167.075 22.400 167.135 ;
        RECT 21.175 166.935 22.400 167.075 ;
        RECT 21.175 166.890 21.465 166.935 ;
        RECT 22.080 166.875 22.400 166.935 ;
        RECT 22.540 166.875 22.860 167.135 ;
        RECT 23.000 167.075 23.320 167.135 ;
        RECT 23.935 167.075 24.225 167.120 ;
        RECT 23.000 166.935 24.225 167.075 ;
        RECT 23.000 166.875 23.320 166.935 ;
        RECT 23.935 166.890 24.225 166.935 ;
        RECT 27.155 166.735 27.445 166.780 ;
        RECT 27.600 166.735 27.920 166.795 ;
        RECT 27.155 166.595 27.920 166.735 ;
        RECT 27.155 166.550 27.445 166.595 ;
        RECT 27.600 166.535 27.920 166.595 ;
        RECT 30.835 166.735 31.125 166.780 ;
        RECT 30.835 166.595 34.270 166.735 ;
        RECT 30.835 166.550 31.125 166.595 ;
        RECT 23.015 166.395 23.305 166.440 ;
        RECT 32.200 166.395 32.520 166.455 ;
        RECT 23.015 166.255 32.520 166.395 ;
        RECT 34.130 166.395 34.270 166.595 ;
        RECT 34.500 166.535 34.820 166.795 ;
        RECT 35.050 166.735 35.190 167.275 ;
        RECT 38.640 167.275 43.105 167.415 ;
        RECT 43.330 167.415 43.470 167.615 ;
        RECT 49.680 167.615 50.445 167.755 ;
        RECT 49.680 167.555 50.000 167.615 ;
        RECT 50.155 167.570 50.445 167.615 ;
        RECT 62.575 167.755 62.865 167.800 ;
        RECT 62.575 167.615 66.930 167.755 ;
        RECT 62.575 167.570 62.865 167.615 ;
        RECT 61.195 167.415 61.485 167.460 ;
        RECT 61.640 167.415 61.960 167.475 ;
        RECT 65.795 167.415 66.085 167.460 ;
        RECT 43.330 167.275 49.910 167.415 ;
        RECT 38.640 167.215 38.960 167.275 ;
        RECT 39.215 167.230 39.805 167.275 ;
        RECT 42.455 167.230 43.105 167.275 ;
        RECT 39.515 166.915 39.805 167.230 ;
        RECT 40.595 167.075 40.885 167.120 ;
        RECT 44.175 167.075 44.465 167.120 ;
        RECT 46.010 167.075 46.300 167.120 ;
        RECT 40.595 166.935 46.300 167.075 ;
        RECT 40.595 166.890 40.885 166.935 ;
        RECT 44.175 166.890 44.465 166.935 ;
        RECT 46.010 166.890 46.300 166.935 ;
        RECT 46.460 166.875 46.780 167.135 ;
        RECT 49.770 167.120 49.910 167.275 ;
        RECT 61.195 167.275 66.085 167.415 ;
        RECT 61.195 167.230 61.485 167.275 ;
        RECT 61.640 167.215 61.960 167.275 ;
        RECT 65.795 167.230 66.085 167.275 ;
        RECT 49.695 167.075 49.985 167.120 ;
        RECT 54.295 167.075 54.585 167.120 ;
        RECT 49.695 166.935 54.585 167.075 ;
        RECT 49.695 166.890 49.985 166.935 ;
        RECT 54.295 166.890 54.585 166.935 ;
        RECT 55.660 166.875 55.980 167.135 ;
        RECT 60.720 167.075 61.040 167.135 ;
        RECT 63.495 167.075 63.785 167.120 ;
        RECT 60.720 166.935 63.785 167.075 ;
        RECT 60.720 166.875 61.040 166.935 ;
        RECT 63.495 166.890 63.785 166.935 ;
        RECT 35.050 166.595 40.250 166.735 ;
        RECT 37.735 166.395 38.025 166.440 ;
        RECT 38.180 166.395 38.500 166.455 ;
        RECT 34.130 166.255 38.500 166.395 ;
        RECT 23.015 166.210 23.305 166.255 ;
        RECT 32.200 166.195 32.520 166.255 ;
        RECT 37.735 166.210 38.025 166.255 ;
        RECT 38.180 166.195 38.500 166.255 ;
        RECT 18.860 166.055 19.180 166.115 ;
        RECT 20.255 166.055 20.545 166.100 ;
        RECT 18.860 165.915 20.545 166.055 ;
        RECT 18.860 165.855 19.180 165.915 ;
        RECT 20.255 165.870 20.545 165.915 ;
        RECT 22.095 166.055 22.385 166.100 ;
        RECT 23.920 166.055 24.240 166.115 ;
        RECT 22.095 165.915 24.240 166.055 ;
        RECT 22.095 165.870 22.385 165.915 ;
        RECT 23.920 165.855 24.240 165.915 ;
        RECT 24.855 166.055 25.145 166.100 ;
        RECT 27.140 166.055 27.460 166.115 ;
        RECT 24.855 165.915 27.460 166.055 ;
        RECT 24.855 165.870 25.145 165.915 ;
        RECT 27.140 165.855 27.460 165.915 ;
        RECT 33.580 165.855 33.900 166.115 ;
        RECT 37.275 166.055 37.565 166.100 ;
        RECT 39.560 166.055 39.880 166.115 ;
        RECT 37.275 165.915 39.880 166.055 ;
        RECT 40.110 166.055 40.250 166.595 ;
        RECT 45.080 166.535 45.400 166.795 ;
        RECT 63.020 166.735 63.340 166.795 ;
        RECT 66.790 166.780 66.930 167.615 ;
        RECT 67.620 167.555 67.940 167.815 ;
        RECT 75.440 167.555 75.760 167.815 ;
        RECT 78.200 167.555 78.520 167.815 ;
        RECT 99.820 167.755 100.140 167.815 ;
        RECT 104.895 167.755 105.185 167.800 ;
        RECT 99.820 167.615 105.185 167.755 ;
        RECT 99.820 167.555 100.140 167.615 ;
        RECT 104.895 167.570 105.185 167.615 ;
        RECT 93.380 167.415 93.700 167.475 ;
        RECT 93.955 167.415 94.245 167.460 ;
        RECT 97.195 167.415 97.845 167.460 ;
        RECT 93.380 167.275 97.845 167.415 ;
        RECT 93.380 167.215 93.700 167.275 ;
        RECT 93.955 167.230 94.545 167.275 ;
        RECT 97.195 167.230 97.845 167.275 ;
        RECT 102.120 167.415 102.440 167.475 ;
        RECT 106.375 167.415 106.665 167.460 ;
        RECT 109.615 167.415 110.265 167.460 ;
        RECT 102.120 167.275 110.265 167.415 ;
        RECT 68.095 167.075 68.385 167.120 ;
        RECT 69.920 167.075 70.240 167.135 ;
        RECT 71.775 167.075 72.065 167.120 ;
        RECT 68.095 166.935 72.065 167.075 ;
        RECT 68.095 166.890 68.385 166.935 ;
        RECT 69.920 166.875 70.240 166.935 ;
        RECT 71.775 166.890 72.065 166.935 ;
        RECT 72.235 167.075 72.525 167.120 ;
        RECT 72.680 167.075 73.000 167.135 ;
        RECT 72.235 166.935 73.000 167.075 ;
        RECT 72.235 166.890 72.525 166.935 ;
        RECT 72.680 166.875 73.000 166.935 ;
        RECT 75.900 166.875 76.220 167.135 ;
        RECT 77.295 167.075 77.585 167.120 ;
        RECT 76.450 166.935 77.585 167.075 ;
        RECT 64.875 166.735 65.165 166.780 ;
        RECT 63.020 166.595 65.165 166.735 ;
        RECT 63.020 166.535 63.340 166.595 ;
        RECT 64.875 166.550 65.165 166.595 ;
        RECT 65.335 166.550 65.625 166.780 ;
        RECT 66.715 166.735 67.005 166.780 ;
        RECT 70.855 166.735 71.145 166.780 ;
        RECT 73.140 166.735 73.460 166.795 ;
        RECT 66.715 166.595 73.460 166.735 ;
        RECT 66.715 166.550 67.005 166.595 ;
        RECT 70.855 166.550 71.145 166.595 ;
        RECT 40.595 166.395 40.885 166.440 ;
        RECT 43.715 166.395 44.005 166.440 ;
        RECT 45.605 166.395 45.895 166.440 ;
        RECT 40.595 166.255 45.895 166.395 ;
        RECT 40.595 166.210 40.885 166.255 ;
        RECT 43.715 166.210 44.005 166.255 ;
        RECT 45.605 166.210 45.895 166.255 ;
        RECT 62.100 166.395 62.420 166.455 ;
        RECT 63.955 166.395 64.245 166.440 ;
        RECT 62.100 166.255 64.245 166.395 ;
        RECT 62.100 166.195 62.420 166.255 ;
        RECT 63.955 166.210 64.245 166.255 ;
        RECT 47.840 166.055 48.160 166.115 ;
        RECT 40.110 165.915 48.160 166.055 ;
        RECT 37.275 165.870 37.565 165.915 ;
        RECT 39.560 165.855 39.880 165.915 ;
        RECT 47.840 165.855 48.160 165.915 ;
        RECT 63.480 166.055 63.800 166.115 ;
        RECT 65.410 166.055 65.550 166.550 ;
        RECT 73.140 166.535 73.460 166.595 ;
        RECT 69.935 166.395 70.225 166.440 ;
        RECT 76.450 166.395 76.590 166.935 ;
        RECT 77.295 166.890 77.585 166.935 ;
        RECT 87.400 166.875 87.720 167.135 ;
        RECT 94.255 166.915 94.545 167.230 ;
        RECT 102.120 167.215 102.440 167.275 ;
        RECT 106.375 167.230 106.965 167.275 ;
        RECT 109.615 167.230 110.265 167.275 ;
        RECT 95.335 167.075 95.625 167.120 ;
        RECT 98.915 167.075 99.205 167.120 ;
        RECT 100.750 167.075 101.040 167.120 ;
        RECT 95.335 166.935 101.040 167.075 ;
        RECT 95.335 166.890 95.625 166.935 ;
        RECT 98.915 166.890 99.205 166.935 ;
        RECT 100.750 166.890 101.040 166.935 ;
        RECT 103.500 166.875 103.820 167.135 ;
        RECT 106.675 166.915 106.965 167.230 ;
        RECT 112.240 167.215 112.560 167.475 ;
        RECT 107.755 167.075 108.045 167.120 ;
        RECT 111.335 167.075 111.625 167.120 ;
        RECT 113.170 167.075 113.460 167.120 ;
        RECT 107.755 166.935 113.460 167.075 ;
        RECT 107.755 166.890 108.045 166.935 ;
        RECT 111.335 166.890 111.625 166.935 ;
        RECT 113.170 166.890 113.460 166.935 ;
        RECT 89.255 166.735 89.545 166.780 ;
        RECT 92.475 166.735 92.765 166.780 ;
        RECT 99.360 166.735 99.680 166.795 ;
        RECT 89.255 166.595 99.680 166.735 ;
        RECT 89.255 166.550 89.545 166.595 ;
        RECT 92.475 166.550 92.765 166.595 ;
        RECT 99.360 166.535 99.680 166.595 ;
        RECT 99.820 166.535 100.140 166.795 ;
        RECT 101.200 166.535 101.520 166.795 ;
        RECT 109.480 166.735 109.800 166.795 ;
        RECT 113.620 166.735 113.940 166.795 ;
        RECT 109.480 166.595 113.940 166.735 ;
        RECT 109.480 166.535 109.800 166.595 ;
        RECT 113.620 166.535 113.940 166.595 ;
        RECT 69.935 166.255 76.590 166.395 ;
        RECT 87.875 166.395 88.165 166.440 ;
        RECT 93.840 166.395 94.160 166.455 ;
        RECT 87.875 166.255 94.160 166.395 ;
        RECT 69.935 166.210 70.225 166.255 ;
        RECT 87.875 166.210 88.165 166.255 ;
        RECT 93.840 166.195 94.160 166.255 ;
        RECT 95.335 166.395 95.625 166.440 ;
        RECT 98.455 166.395 98.745 166.440 ;
        RECT 100.345 166.395 100.635 166.440 ;
        RECT 95.335 166.255 100.635 166.395 ;
        RECT 95.335 166.210 95.625 166.255 ;
        RECT 98.455 166.210 98.745 166.255 ;
        RECT 100.345 166.210 100.635 166.255 ;
        RECT 107.755 166.395 108.045 166.440 ;
        RECT 110.875 166.395 111.165 166.440 ;
        RECT 112.765 166.395 113.055 166.440 ;
        RECT 107.755 166.255 113.055 166.395 ;
        RECT 107.755 166.210 108.045 166.255 ;
        RECT 110.875 166.210 111.165 166.255 ;
        RECT 112.765 166.210 113.055 166.255 ;
        RECT 63.480 165.915 65.550 166.055 ;
        RECT 74.075 166.055 74.365 166.100 ;
        RECT 78.660 166.055 78.980 166.115 ;
        RECT 74.075 165.915 78.980 166.055 ;
        RECT 63.480 165.855 63.800 165.915 ;
        RECT 74.075 165.870 74.365 165.915 ;
        RECT 78.660 165.855 78.980 165.915 ;
        RECT 92.015 166.055 92.305 166.100 ;
        RECT 92.920 166.055 93.240 166.115 ;
        RECT 92.015 165.915 93.240 166.055 ;
        RECT 92.015 165.870 92.305 165.915 ;
        RECT 92.920 165.855 93.240 165.915 ;
        RECT 103.960 165.855 104.280 166.115 ;
        RECT 10.510 165.235 115.850 165.715 ;
        RECT 135.580 165.470 136.830 166.590 ;
        RECT 16.575 165.035 16.865 165.080 ;
        RECT 27.600 165.035 27.920 165.095 ;
        RECT 40.940 165.035 41.260 165.095 ;
        RECT 16.575 164.895 41.260 165.035 ;
        RECT 16.575 164.850 16.865 164.895 ;
        RECT 27.600 164.835 27.920 164.895 ;
        RECT 40.940 164.835 41.260 164.895 ;
        RECT 52.915 165.035 53.205 165.080 ;
        RECT 54.740 165.035 55.060 165.095 ;
        RECT 52.915 164.895 55.060 165.035 ;
        RECT 52.915 164.850 53.205 164.895 ;
        RECT 54.740 164.835 55.060 164.895 ;
        RECT 73.140 165.035 73.460 165.095 ;
        RECT 84.180 165.035 84.500 165.095 ;
        RECT 96.155 165.035 96.445 165.080 ;
        RECT 99.820 165.035 100.140 165.095 ;
        RECT 73.140 164.895 84.870 165.035 ;
        RECT 73.140 164.835 73.460 164.895 ;
        RECT 84.180 164.835 84.500 164.895 ;
        RECT 19.435 164.695 19.725 164.740 ;
        RECT 22.555 164.695 22.845 164.740 ;
        RECT 24.445 164.695 24.735 164.740 ;
        RECT 19.435 164.555 24.735 164.695 ;
        RECT 19.435 164.510 19.725 164.555 ;
        RECT 22.555 164.510 22.845 164.555 ;
        RECT 24.445 164.510 24.735 164.555 ;
        RECT 31.855 164.695 32.145 164.740 ;
        RECT 34.975 164.695 35.265 164.740 ;
        RECT 36.865 164.695 37.155 164.740 ;
        RECT 31.855 164.555 37.155 164.695 ;
        RECT 31.855 164.510 32.145 164.555 ;
        RECT 34.975 164.510 35.265 164.555 ;
        RECT 36.865 164.510 37.155 164.555 ;
        RECT 38.655 164.510 38.945 164.740 ;
        RECT 72.190 164.695 72.480 164.740 ;
        RECT 74.970 164.695 75.260 164.740 ;
        RECT 76.830 164.695 77.120 164.740 ;
        RECT 72.190 164.555 77.120 164.695 ;
        RECT 72.190 164.510 72.480 164.555 ;
        RECT 74.970 164.510 75.260 164.555 ;
        RECT 76.830 164.510 77.120 164.555 ;
        RECT 23.920 164.155 24.240 164.415 ;
        RECT 25.300 164.355 25.620 164.415 ;
        RECT 25.300 164.215 28.750 164.355 ;
        RECT 25.300 164.155 25.620 164.215 ;
        RECT 28.610 164.060 28.750 164.215 ;
        RECT 28.980 164.155 29.300 164.415 ;
        RECT 36.355 164.355 36.645 164.400 ;
        RECT 38.730 164.355 38.870 164.510 ;
        RECT 36.355 164.215 38.870 164.355 ;
        RECT 39.100 164.355 39.420 164.415 ;
        RECT 42.795 164.355 43.085 164.400 ;
        RECT 46.935 164.355 47.225 164.400 ;
        RECT 56.580 164.355 56.900 164.415 ;
        RECT 58.435 164.355 58.725 164.400 ;
        RECT 68.325 164.355 68.615 164.400 ;
        RECT 69.920 164.355 70.240 164.415 ;
        RECT 39.100 164.215 52.670 164.355 ;
        RECT 36.355 164.170 36.645 164.215 ;
        RECT 39.100 164.155 39.420 164.215 ;
        RECT 42.795 164.170 43.085 164.215 ;
        RECT 46.935 164.170 47.225 164.215 ;
        RECT 18.355 163.720 18.645 164.035 ;
        RECT 19.435 164.015 19.725 164.060 ;
        RECT 23.015 164.015 23.305 164.060 ;
        RECT 24.850 164.015 25.140 164.060 ;
        RECT 19.435 163.875 25.140 164.015 ;
        RECT 19.435 163.830 19.725 163.875 ;
        RECT 23.015 163.830 23.305 163.875 ;
        RECT 24.850 163.830 25.140 163.875 ;
        RECT 28.535 163.830 28.825 164.060 ;
        RECT 18.055 163.675 18.645 163.720 ;
        RECT 18.860 163.675 19.180 163.735 ;
        RECT 21.295 163.675 21.945 163.720 ;
        RECT 18.055 163.535 21.945 163.675 ;
        RECT 18.055 163.490 18.345 163.535 ;
        RECT 18.860 163.475 19.180 163.535 ;
        RECT 21.295 163.490 21.945 163.535 ;
        RECT 28.610 163.335 28.750 163.830 ;
        RECT 30.775 163.720 31.065 164.035 ;
        RECT 31.855 164.015 32.145 164.060 ;
        RECT 35.435 164.015 35.725 164.060 ;
        RECT 37.270 164.015 37.560 164.060 ;
        RECT 31.855 163.875 37.560 164.015 ;
        RECT 31.855 163.830 32.145 163.875 ;
        RECT 35.435 163.830 35.725 163.875 ;
        RECT 37.270 163.830 37.560 163.875 ;
        RECT 37.735 163.830 38.025 164.060 ;
        RECT 30.475 163.675 31.065 163.720 ;
        RECT 31.280 163.675 31.600 163.735 ;
        RECT 33.715 163.675 34.365 163.720 ;
        RECT 37.810 163.675 37.950 163.830 ;
        RECT 39.560 163.815 39.880 164.075 ;
        RECT 43.700 164.015 44.020 164.075 ;
        RECT 47.395 164.015 47.685 164.060 ;
        RECT 43.700 163.875 47.685 164.015 ;
        RECT 43.700 163.815 44.020 163.875 ;
        RECT 47.395 163.830 47.685 163.875 ;
        RECT 47.840 163.815 48.160 164.075 ;
        RECT 51.995 164.015 52.285 164.060 ;
        RECT 49.770 163.875 52.285 164.015 ;
        RECT 30.475 163.535 34.365 163.675 ;
        RECT 30.475 163.490 30.765 163.535 ;
        RECT 31.280 163.475 31.600 163.535 ;
        RECT 33.715 163.490 34.365 163.535 ;
        RECT 37.350 163.535 37.950 163.675 ;
        RECT 37.350 163.335 37.490 163.535 ;
        RECT 28.610 163.195 37.490 163.335 ;
        RECT 38.180 163.335 38.500 163.395 ;
        RECT 43.255 163.335 43.545 163.380 ;
        RECT 38.180 163.195 43.545 163.335 ;
        RECT 38.180 163.135 38.500 163.195 ;
        RECT 43.255 163.150 43.545 163.195 ;
        RECT 45.555 163.335 45.845 163.380 ;
        RECT 46.000 163.335 46.320 163.395 ;
        RECT 49.770 163.380 49.910 163.875 ;
        RECT 51.995 163.830 52.285 163.875 ;
        RECT 52.530 163.675 52.670 164.215 ;
        RECT 56.580 164.215 67.850 164.355 ;
        RECT 56.580 164.155 56.900 164.215 ;
        RECT 58.435 164.170 58.725 164.215 ;
        RECT 55.660 164.015 55.980 164.075 ;
        RECT 56.135 164.015 56.425 164.060 ;
        RECT 59.340 164.015 59.660 164.075 ;
        RECT 55.660 163.875 59.660 164.015 ;
        RECT 55.660 163.815 55.980 163.875 ;
        RECT 56.135 163.830 56.425 163.875 ;
        RECT 59.340 163.815 59.660 163.875 ;
        RECT 61.640 163.815 61.960 164.075 ;
        RECT 59.815 163.675 60.105 163.720 ;
        RECT 52.530 163.535 60.105 163.675 ;
        RECT 59.815 163.490 60.105 163.535 ;
        RECT 45.555 163.195 46.320 163.335 ;
        RECT 45.555 163.150 45.845 163.195 ;
        RECT 46.000 163.135 46.320 163.195 ;
        RECT 49.695 163.150 49.985 163.380 ;
        RECT 55.675 163.335 55.965 163.380 ;
        RECT 58.420 163.335 58.740 163.395 ;
        RECT 55.675 163.195 58.740 163.335 ;
        RECT 67.710 163.335 67.850 164.215 ;
        RECT 68.325 164.215 70.240 164.355 ;
        RECT 68.325 164.170 68.615 164.215 ;
        RECT 69.920 164.155 70.240 164.215 ;
        RECT 77.295 164.355 77.585 164.400 ;
        RECT 83.260 164.355 83.580 164.415 ;
        RECT 77.295 164.215 83.580 164.355 ;
        RECT 84.730 164.355 84.870 164.895 ;
        RECT 96.155 164.895 100.140 165.035 ;
        RECT 96.155 164.850 96.445 164.895 ;
        RECT 99.820 164.835 100.140 164.895 ;
        RECT 102.120 164.835 102.440 165.095 ;
        RECT 105.915 164.695 106.205 164.740 ;
        RECT 109.035 164.695 109.325 164.740 ;
        RECT 110.925 164.695 111.215 164.740 ;
        RECT 105.915 164.555 111.215 164.695 ;
        RECT 105.915 164.510 106.205 164.555 ;
        RECT 109.035 164.510 109.325 164.555 ;
        RECT 110.925 164.510 111.215 164.555 ;
        RECT 85.115 164.355 85.405 164.400 ;
        RECT 91.555 164.355 91.845 164.400 ;
        RECT 98.440 164.355 98.760 164.415 ;
        RECT 99.375 164.355 99.665 164.400 ;
        RECT 84.730 164.215 99.665 164.355 ;
        RECT 77.295 164.170 77.585 164.215 ;
        RECT 83.260 164.155 83.580 164.215 ;
        RECT 85.115 164.170 85.405 164.215 ;
        RECT 91.555 164.170 91.845 164.215 ;
        RECT 98.440 164.155 98.760 164.215 ;
        RECT 99.375 164.170 99.665 164.215 ;
        RECT 109.940 164.355 110.260 164.415 ;
        RECT 111.795 164.355 112.085 164.400 ;
        RECT 109.940 164.215 112.085 164.355 ;
        RECT 72.190 164.015 72.480 164.060 ;
        RECT 75.455 164.015 75.745 164.060 ;
        RECT 72.190 163.875 74.725 164.015 ;
        RECT 72.190 163.830 72.480 163.875 ;
        RECT 70.330 163.675 70.620 163.720 ;
        RECT 71.760 163.675 72.080 163.735 ;
        RECT 74.510 163.720 74.725 163.875 ;
        RECT 75.455 163.875 77.970 164.015 ;
        RECT 75.455 163.830 75.745 163.875 ;
        RECT 73.590 163.675 73.880 163.720 ;
        RECT 70.330 163.535 73.880 163.675 ;
        RECT 70.330 163.490 70.620 163.535 ;
        RECT 71.760 163.475 72.080 163.535 ;
        RECT 73.590 163.490 73.880 163.535 ;
        RECT 74.510 163.675 74.800 163.720 ;
        RECT 76.370 163.675 76.660 163.720 ;
        RECT 74.510 163.535 76.660 163.675 ;
        RECT 74.510 163.490 74.800 163.535 ;
        RECT 76.370 163.490 76.660 163.535 ;
        RECT 75.440 163.335 75.760 163.395 ;
        RECT 77.830 163.380 77.970 163.875 ;
        RECT 78.660 163.815 78.980 164.075 ;
        RECT 92.920 163.815 93.240 164.075 ;
        RECT 93.380 164.015 93.700 164.075 ;
        RECT 95.235 164.015 95.525 164.060 ;
        RECT 93.380 163.875 95.525 164.015 ;
        RECT 93.380 163.815 93.700 163.875 ;
        RECT 95.235 163.830 95.525 163.875 ;
        RECT 86.495 163.675 86.785 163.720 ;
        RECT 89.700 163.675 90.020 163.735 ;
        RECT 92.475 163.675 92.765 163.720 ;
        RECT 86.495 163.535 92.765 163.675 ;
        RECT 99.450 163.675 99.590 164.170 ;
        RECT 109.940 164.155 110.260 164.215 ;
        RECT 111.795 164.170 112.085 164.215 ;
        RECT 101.675 164.015 101.965 164.060 ;
        RECT 103.500 164.015 103.820 164.075 ;
        RECT 101.675 163.875 103.820 164.015 ;
        RECT 101.675 163.830 101.965 163.875 ;
        RECT 103.500 163.815 103.820 163.875 ;
        RECT 103.960 163.675 104.280 163.735 ;
        RECT 104.835 163.720 105.125 164.035 ;
        RECT 105.915 164.015 106.205 164.060 ;
        RECT 109.495 164.015 109.785 164.060 ;
        RECT 111.330 164.015 111.620 164.060 ;
        RECT 105.915 163.875 111.620 164.015 ;
        RECT 105.915 163.830 106.205 163.875 ;
        RECT 109.495 163.830 109.785 163.875 ;
        RECT 111.330 163.830 111.620 163.875 ;
        RECT 113.160 163.815 113.480 164.075 ;
        RECT 104.535 163.675 105.125 163.720 ;
        RECT 107.775 163.675 108.425 163.720 ;
        RECT 99.450 163.535 100.510 163.675 ;
        RECT 86.495 163.490 86.785 163.535 ;
        RECT 89.700 163.475 90.020 163.535 ;
        RECT 92.475 163.490 92.765 163.535 ;
        RECT 67.710 163.195 75.760 163.335 ;
        RECT 55.675 163.150 55.965 163.195 ;
        RECT 58.420 163.135 58.740 163.195 ;
        RECT 75.440 163.135 75.760 163.195 ;
        RECT 77.755 163.150 78.045 163.380 ;
        RECT 79.580 163.335 79.900 163.395 ;
        RECT 86.035 163.335 86.325 163.380 ;
        RECT 79.580 163.195 86.325 163.335 ;
        RECT 79.580 163.135 79.900 163.195 ;
        RECT 86.035 163.150 86.325 163.195 ;
        RECT 88.335 163.335 88.625 163.380 ;
        RECT 91.080 163.335 91.400 163.395 ;
        RECT 88.335 163.195 91.400 163.335 ;
        RECT 88.335 163.150 88.625 163.195 ;
        RECT 91.080 163.135 91.400 163.195 ;
        RECT 94.300 163.335 94.620 163.395 ;
        RECT 94.775 163.335 95.065 163.380 ;
        RECT 94.300 163.195 95.065 163.335 ;
        RECT 94.300 163.135 94.620 163.195 ;
        RECT 94.775 163.150 95.065 163.195 ;
        RECT 96.615 163.335 96.905 163.380 ;
        RECT 97.060 163.335 97.380 163.395 ;
        RECT 96.615 163.195 97.380 163.335 ;
        RECT 96.615 163.150 96.905 163.195 ;
        RECT 97.060 163.135 97.380 163.195 ;
        RECT 98.440 163.135 98.760 163.395 ;
        RECT 98.915 163.335 99.205 163.380 ;
        RECT 99.820 163.335 100.140 163.395 ;
        RECT 98.915 163.195 100.140 163.335 ;
        RECT 100.370 163.335 100.510 163.535 ;
        RECT 103.960 163.535 108.425 163.675 ;
        RECT 103.960 163.475 104.280 163.535 ;
        RECT 104.535 163.490 104.825 163.535 ;
        RECT 107.775 163.490 108.425 163.535 ;
        RECT 110.415 163.675 110.705 163.720 ;
        RECT 110.415 163.535 112.470 163.675 ;
        RECT 110.415 163.490 110.705 163.535 ;
        RECT 101.660 163.335 101.980 163.395 ;
        RECT 100.370 163.195 101.980 163.335 ;
        RECT 98.915 163.150 99.205 163.195 ;
        RECT 99.820 163.135 100.140 163.195 ;
        RECT 101.660 163.135 101.980 163.195 ;
        RECT 103.055 163.335 103.345 163.380 ;
        RECT 103.500 163.335 103.820 163.395 ;
        RECT 112.330 163.380 112.470 163.535 ;
        RECT 103.055 163.195 103.820 163.335 ;
        RECT 103.055 163.150 103.345 163.195 ;
        RECT 103.500 163.135 103.820 163.195 ;
        RECT 112.255 163.150 112.545 163.380 ;
        RECT 10.510 162.515 115.850 162.995 ;
        RECT 17.955 162.130 18.245 162.360 ;
        RECT 20.715 162.315 21.005 162.360 ;
        RECT 22.080 162.315 22.400 162.375 ;
        RECT 20.715 162.175 22.400 162.315 ;
        RECT 20.715 162.130 21.005 162.175 ;
        RECT 18.030 161.975 18.170 162.130 ;
        RECT 22.080 162.115 22.400 162.175 ;
        RECT 30.360 162.315 30.680 162.375 ;
        RECT 34.515 162.315 34.805 162.360 ;
        RECT 30.360 162.175 34.805 162.315 ;
        RECT 30.360 162.115 30.680 162.175 ;
        RECT 34.515 162.130 34.805 162.175 ;
        RECT 39.560 162.315 39.880 162.375 ;
        RECT 39.560 162.175 42.550 162.315 ;
        RECT 39.560 162.115 39.880 162.175 ;
        RECT 23.015 161.975 23.305 162.020 ;
        RECT 23.460 161.975 23.780 162.035 ;
        RECT 18.030 161.835 22.770 161.975 ;
        RECT 22.630 161.695 22.770 161.835 ;
        RECT 23.015 161.835 23.780 161.975 ;
        RECT 23.015 161.790 23.305 161.835 ;
        RECT 23.460 161.775 23.780 161.835 ;
        RECT 27.140 161.775 27.460 162.035 ;
        RECT 29.435 161.975 30.085 162.020 ;
        RECT 32.200 161.975 32.520 162.035 ;
        RECT 33.035 161.975 33.325 162.020 ;
        RECT 37.275 161.975 37.565 162.020 ;
        RECT 38.180 161.975 38.500 162.035 ;
        RECT 29.435 161.835 33.325 161.975 ;
        RECT 29.435 161.790 30.085 161.835 ;
        RECT 32.200 161.775 32.520 161.835 ;
        RECT 32.735 161.790 33.325 161.835 ;
        RECT 35.510 161.835 38.500 161.975 ;
        RECT 15.195 161.635 15.485 161.680 ;
        RECT 17.940 161.635 18.260 161.695 ;
        RECT 15.195 161.495 18.260 161.635 ;
        RECT 15.195 161.450 15.485 161.495 ;
        RECT 17.940 161.435 18.260 161.495 ;
        RECT 18.400 161.435 18.720 161.695 ;
        RECT 22.540 161.435 22.860 161.695 ;
        RECT 25.300 161.635 25.620 161.695 ;
        RECT 25.775 161.635 26.065 161.680 ;
        RECT 25.300 161.495 26.065 161.635 ;
        RECT 25.300 161.435 25.620 161.495 ;
        RECT 25.775 161.450 26.065 161.495 ;
        RECT 26.240 161.635 26.530 161.680 ;
        RECT 28.075 161.635 28.365 161.680 ;
        RECT 31.655 161.635 31.945 161.680 ;
        RECT 26.240 161.495 31.945 161.635 ;
        RECT 26.240 161.450 26.530 161.495 ;
        RECT 28.075 161.450 28.365 161.495 ;
        RECT 31.655 161.450 31.945 161.495 ;
        RECT 32.735 161.475 33.025 161.790 ;
        RECT 17.495 161.295 17.785 161.340 ;
        RECT 23.935 161.295 24.225 161.340 ;
        RECT 24.840 161.295 25.160 161.355 ;
        RECT 17.495 161.155 25.160 161.295 ;
        RECT 17.495 161.110 17.785 161.155 ;
        RECT 23.935 161.110 24.225 161.155 ;
        RECT 24.840 161.095 25.160 161.155 ;
        RECT 33.580 161.295 33.900 161.355 ;
        RECT 35.510 161.295 35.650 161.835 ;
        RECT 37.275 161.790 37.565 161.835 ;
        RECT 38.180 161.775 38.500 161.835 ;
        RECT 38.640 161.975 38.960 162.035 ;
        RECT 42.410 161.975 42.550 162.175 ;
        RECT 45.080 162.115 45.400 162.375 ;
        RECT 59.815 162.315 60.105 162.360 ;
        RECT 70.840 162.315 71.160 162.375 ;
        RECT 59.815 162.175 71.160 162.315 ;
        RECT 59.815 162.130 60.105 162.175 ;
        RECT 59.890 161.975 60.030 162.130 ;
        RECT 70.840 162.115 71.160 162.175 ;
        RECT 71.760 162.115 72.080 162.375 ;
        RECT 75.900 162.315 76.220 162.375 ;
        RECT 73.230 162.175 76.220 162.315 ;
        RECT 73.230 161.975 73.370 162.175 ;
        RECT 75.900 162.115 76.220 162.175 ;
        RECT 95.220 162.315 95.540 162.375 ;
        RECT 97.060 162.315 97.380 162.375 ;
        RECT 95.220 162.175 97.380 162.315 ;
        RECT 95.220 162.115 95.540 162.175 ;
        RECT 97.060 162.115 97.380 162.175 ;
        RECT 113.160 162.315 113.480 162.375 ;
        RECT 114.095 162.315 114.385 162.360 ;
        RECT 113.160 162.175 114.385 162.315 ;
        RECT 113.160 162.115 113.480 162.175 ;
        RECT 114.095 162.130 114.385 162.175 ;
        RECT 79.580 161.975 79.900 162.035 ;
        RECT 80.745 161.975 81.035 162.020 ;
        RECT 38.640 161.835 42.090 161.975 ;
        RECT 42.410 161.835 60.030 161.975 ;
        RECT 60.810 161.835 62.330 161.975 ;
        RECT 38.640 161.775 38.960 161.835 ;
        RECT 40.020 161.635 40.340 161.695 ;
        RECT 41.950 161.680 42.090 161.835 ;
        RECT 40.955 161.635 41.245 161.680 ;
        RECT 40.020 161.495 41.245 161.635 ;
        RECT 40.020 161.435 40.340 161.495 ;
        RECT 40.955 161.450 41.245 161.495 ;
        RECT 41.875 161.450 42.165 161.680 ;
        RECT 42.335 161.450 42.625 161.680 ;
        RECT 42.795 161.635 43.085 161.680 ;
        RECT 45.080 161.635 45.400 161.695 ;
        RECT 42.795 161.495 45.400 161.635 ;
        RECT 42.795 161.450 43.085 161.495 ;
        RECT 37.735 161.295 38.025 161.340 ;
        RECT 33.580 161.155 35.650 161.295 ;
        RECT 35.970 161.155 38.025 161.295 ;
        RECT 33.580 161.095 33.900 161.155 ;
        RECT 26.645 160.955 26.935 161.000 ;
        RECT 28.535 160.955 28.825 161.000 ;
        RECT 31.655 160.955 31.945 161.000 ;
        RECT 26.645 160.815 31.945 160.955 ;
        RECT 26.645 160.770 26.935 160.815 ;
        RECT 28.535 160.770 28.825 160.815 ;
        RECT 31.655 160.770 31.945 160.815 ;
        RECT 34.500 160.955 34.820 161.015 ;
        RECT 35.435 160.955 35.725 161.000 ;
        RECT 34.500 160.815 35.725 160.955 ;
        RECT 34.500 160.755 34.820 160.815 ;
        RECT 35.435 160.770 35.725 160.815 ;
        RECT 15.640 160.415 15.960 160.675 ;
        RECT 20.255 160.615 20.545 160.660 ;
        RECT 23.460 160.615 23.780 160.675 ;
        RECT 20.255 160.475 23.780 160.615 ;
        RECT 20.255 160.430 20.545 160.475 ;
        RECT 23.460 160.415 23.780 160.475 ;
        RECT 28.980 160.615 29.300 160.675 ;
        RECT 35.970 160.615 36.110 161.155 ;
        RECT 37.735 161.110 38.025 161.155 ;
        RECT 38.195 161.295 38.485 161.340 ;
        RECT 39.100 161.295 39.420 161.355 ;
        RECT 38.195 161.155 39.420 161.295 ;
        RECT 42.410 161.295 42.550 161.450 ;
        RECT 45.080 161.435 45.400 161.495 ;
        RECT 46.000 161.435 46.320 161.695 ;
        RECT 47.840 161.635 48.160 161.695 ;
        RECT 49.695 161.635 49.985 161.680 ;
        RECT 57.960 161.635 58.280 161.695 ;
        RECT 47.840 161.495 58.280 161.635 ;
        RECT 47.840 161.435 48.160 161.495 ;
        RECT 49.695 161.450 49.985 161.495 ;
        RECT 57.960 161.435 58.280 161.495 ;
        RECT 58.895 161.635 59.185 161.680 ;
        RECT 60.260 161.635 60.580 161.695 ;
        RECT 60.810 161.680 60.950 161.835 ;
        RECT 62.190 161.695 62.330 161.835 ;
        RECT 72.310 161.835 73.370 161.975 ;
        RECT 74.610 161.835 81.035 161.975 ;
        RECT 58.895 161.495 60.580 161.635 ;
        RECT 58.895 161.450 59.185 161.495 ;
        RECT 60.260 161.435 60.580 161.495 ;
        RECT 60.735 161.450 61.025 161.680 ;
        RECT 61.180 161.435 61.500 161.695 ;
        RECT 62.100 161.635 62.420 161.695 ;
        RECT 72.310 161.680 72.450 161.835 ;
        RECT 74.610 161.695 74.750 161.835 ;
        RECT 79.580 161.775 79.900 161.835 ;
        RECT 80.745 161.790 81.035 161.835 ;
        RECT 82.750 161.975 83.040 162.020 ;
        RECT 85.100 161.975 85.420 162.035 ;
        RECT 86.010 161.975 86.300 162.020 ;
        RECT 82.750 161.835 86.300 161.975 ;
        RECT 82.750 161.790 83.040 161.835 ;
        RECT 85.100 161.775 85.420 161.835 ;
        RECT 86.010 161.790 86.300 161.835 ;
        RECT 86.930 161.975 87.220 162.020 ;
        RECT 88.790 161.975 89.080 162.020 ;
        RECT 86.930 161.835 89.080 161.975 ;
        RECT 86.930 161.790 87.220 161.835 ;
        RECT 88.790 161.790 89.080 161.835 ;
        RECT 92.410 161.975 92.700 162.020 ;
        RECT 93.840 161.975 94.160 162.035 ;
        RECT 95.670 161.975 95.960 162.020 ;
        RECT 92.410 161.835 95.960 161.975 ;
        RECT 92.410 161.790 92.700 161.835 ;
        RECT 63.035 161.635 63.325 161.680 ;
        RECT 62.100 161.495 63.325 161.635 ;
        RECT 62.100 161.435 62.420 161.495 ;
        RECT 63.035 161.450 63.325 161.495 ;
        RECT 72.235 161.450 72.525 161.680 ;
        RECT 72.680 161.635 73.000 161.695 ;
        RECT 74.075 161.635 74.365 161.680 ;
        RECT 72.680 161.495 74.365 161.635 ;
        RECT 72.680 161.435 73.000 161.495 ;
        RECT 74.075 161.450 74.365 161.495 ;
        RECT 74.520 161.435 74.840 161.695 ;
        RECT 75.900 161.635 76.220 161.695 ;
        RECT 78.215 161.635 78.505 161.680 ;
        RECT 78.660 161.635 78.980 161.695 ;
        RECT 75.900 161.495 78.980 161.635 ;
        RECT 75.900 161.435 76.220 161.495 ;
        RECT 78.215 161.450 78.505 161.495 ;
        RECT 78.660 161.435 78.980 161.495 ;
        RECT 79.135 161.450 79.425 161.680 ;
        RECT 84.610 161.635 84.900 161.680 ;
        RECT 86.930 161.635 87.145 161.790 ;
        RECT 93.840 161.775 94.160 161.835 ;
        RECT 95.670 161.790 95.960 161.835 ;
        RECT 96.590 161.975 96.880 162.020 ;
        RECT 98.450 161.975 98.740 162.020 ;
        RECT 104.895 161.975 105.185 162.020 ;
        RECT 96.590 161.835 98.740 161.975 ;
        RECT 96.590 161.790 96.880 161.835 ;
        RECT 98.450 161.790 98.740 161.835 ;
        RECT 101.750 161.835 105.185 161.975 ;
        RECT 84.610 161.495 87.145 161.635 ;
        RECT 87.875 161.635 88.165 161.680 ;
        RECT 90.160 161.635 90.480 161.695 ;
        RECT 87.875 161.495 90.480 161.635 ;
        RECT 84.610 161.450 84.900 161.495 ;
        RECT 87.875 161.450 88.165 161.495 ;
        RECT 43.240 161.295 43.560 161.355 ;
        RECT 69.000 161.295 69.320 161.355 ;
        RECT 42.410 161.155 43.560 161.295 ;
        RECT 38.195 161.110 38.485 161.155 ;
        RECT 36.340 160.955 36.660 161.015 ;
        RECT 38.270 160.955 38.410 161.110 ;
        RECT 39.100 161.095 39.420 161.155 ;
        RECT 43.240 161.095 43.560 161.155 ;
        RECT 58.050 161.155 69.320 161.295 ;
        RECT 58.050 161.000 58.190 161.155 ;
        RECT 69.000 161.095 69.320 161.155 ;
        RECT 73.140 161.095 73.460 161.355 ;
        RECT 79.210 161.295 79.350 161.450 ;
        RECT 90.160 161.435 90.480 161.495 ;
        RECT 94.270 161.635 94.560 161.680 ;
        RECT 96.590 161.635 96.805 161.790 ;
        RECT 94.270 161.495 96.805 161.635 ;
        RECT 100.280 161.635 100.600 161.695 ;
        RECT 101.750 161.635 101.890 161.835 ;
        RECT 104.895 161.790 105.185 161.835 ;
        RECT 100.280 161.495 101.890 161.635 ;
        RECT 94.270 161.450 94.560 161.495 ;
        RECT 100.280 161.435 100.600 161.495 ;
        RECT 102.120 161.435 102.440 161.695 ;
        RECT 103.500 161.635 103.820 161.695 ;
        RECT 104.435 161.635 104.725 161.680 ;
        RECT 109.955 161.635 110.245 161.680 ;
        RECT 103.500 161.495 110.245 161.635 ;
        RECT 103.500 161.435 103.820 161.495 ;
        RECT 104.435 161.450 104.725 161.495 ;
        RECT 109.955 161.450 110.245 161.495 ;
        RECT 76.450 161.155 79.350 161.295 ;
        RECT 83.260 161.295 83.580 161.355 ;
        RECT 86.480 161.295 86.800 161.355 ;
        RECT 89.715 161.295 90.005 161.340 ;
        RECT 83.260 161.155 90.005 161.295 ;
        RECT 57.975 160.955 58.265 161.000 ;
        RECT 36.340 160.815 38.410 160.955 ;
        RECT 49.770 160.815 58.265 160.955 ;
        RECT 36.340 160.755 36.660 160.815 ;
        RECT 28.980 160.475 36.110 160.615 ;
        RECT 28.980 160.415 29.300 160.475 ;
        RECT 44.160 160.415 44.480 160.675 ;
        RECT 45.080 160.615 45.400 160.675 ;
        RECT 49.770 160.615 49.910 160.815 ;
        RECT 57.975 160.770 58.265 160.815 ;
        RECT 60.260 160.955 60.580 161.015 ;
        RECT 76.450 161.000 76.590 161.155 ;
        RECT 83.260 161.095 83.580 161.155 ;
        RECT 86.480 161.095 86.800 161.155 ;
        RECT 89.715 161.110 90.005 161.155 ;
        RECT 96.140 161.295 96.460 161.355 ;
        RECT 97.535 161.295 97.825 161.340 ;
        RECT 96.140 161.155 97.825 161.295 ;
        RECT 96.140 161.095 96.460 161.155 ;
        RECT 97.535 161.110 97.825 161.155 ;
        RECT 99.375 161.295 99.665 161.340 ;
        RECT 100.740 161.295 101.060 161.355 ;
        RECT 99.375 161.155 101.060 161.295 ;
        RECT 99.375 161.110 99.665 161.155 ;
        RECT 100.740 161.095 101.060 161.155 ;
        RECT 101.215 161.295 101.505 161.340 ;
        RECT 103.040 161.295 103.360 161.355 ;
        RECT 101.215 161.155 103.360 161.295 ;
        RECT 101.215 161.110 101.505 161.155 ;
        RECT 103.040 161.095 103.360 161.155 ;
        RECT 103.975 161.110 104.265 161.340 ;
        RECT 110.875 161.110 111.165 161.340 ;
        RECT 62.115 160.955 62.405 161.000 ;
        RECT 60.260 160.815 76.130 160.955 ;
        RECT 60.260 160.755 60.580 160.815 ;
        RECT 62.115 160.770 62.405 160.815 ;
        RECT 45.080 160.475 49.910 160.615 ;
        RECT 50.155 160.615 50.445 160.660 ;
        RECT 51.980 160.615 52.300 160.675 ;
        RECT 50.155 160.475 52.300 160.615 ;
        RECT 45.080 160.415 45.400 160.475 ;
        RECT 50.155 160.430 50.445 160.475 ;
        RECT 51.980 160.415 52.300 160.475 ;
        RECT 52.440 160.615 52.760 160.675 ;
        RECT 63.955 160.615 64.245 160.660 ;
        RECT 70.380 160.615 70.700 160.675 ;
        RECT 52.440 160.475 70.700 160.615 ;
        RECT 52.440 160.415 52.760 160.475 ;
        RECT 63.955 160.430 64.245 160.475 ;
        RECT 70.380 160.415 70.700 160.475 ;
        RECT 70.840 160.615 71.160 160.675 ;
        RECT 74.980 160.615 75.300 160.675 ;
        RECT 70.840 160.475 75.300 160.615 ;
        RECT 75.990 160.615 76.130 160.815 ;
        RECT 76.375 160.770 76.665 161.000 ;
        RECT 84.610 160.955 84.900 161.000 ;
        RECT 87.390 160.955 87.680 161.000 ;
        RECT 89.250 160.955 89.540 161.000 ;
        RECT 77.370 160.815 84.410 160.955 ;
        RECT 77.370 160.615 77.510 160.815 ;
        RECT 75.990 160.475 77.510 160.615 ;
        RECT 77.755 160.615 78.045 160.660 ;
        RECT 78.200 160.615 78.520 160.675 ;
        RECT 77.755 160.475 78.520 160.615 ;
        RECT 70.840 160.415 71.160 160.475 ;
        RECT 74.980 160.415 75.300 160.475 ;
        RECT 77.755 160.430 78.045 160.475 ;
        RECT 78.200 160.415 78.520 160.475 ;
        RECT 80.055 160.615 80.345 160.660 ;
        RECT 81.880 160.615 82.200 160.675 ;
        RECT 80.055 160.475 82.200 160.615 ;
        RECT 84.270 160.615 84.410 160.815 ;
        RECT 84.610 160.815 89.540 160.955 ;
        RECT 84.610 160.770 84.900 160.815 ;
        RECT 87.390 160.770 87.680 160.815 ;
        RECT 89.250 160.770 89.540 160.815 ;
        RECT 94.270 160.955 94.560 161.000 ;
        RECT 97.050 160.955 97.340 161.000 ;
        RECT 98.910 160.955 99.200 161.000 ;
        RECT 94.270 160.815 99.200 160.955 ;
        RECT 94.270 160.770 94.560 160.815 ;
        RECT 97.050 160.770 97.340 160.815 ;
        RECT 98.910 160.770 99.200 160.815 ;
        RECT 101.660 160.955 101.980 161.015 ;
        RECT 104.050 160.955 104.190 161.110 ;
        RECT 101.660 160.815 104.190 160.955 ;
        RECT 106.735 160.955 107.025 161.000 ;
        RECT 110.950 160.955 111.090 161.110 ;
        RECT 106.735 160.815 111.090 160.955 ;
        RECT 101.660 160.755 101.980 160.815 ;
        RECT 106.735 160.770 107.025 160.815 ;
        RECT 87.860 160.615 88.180 160.675 ;
        RECT 84.270 160.475 88.180 160.615 ;
        RECT 80.055 160.430 80.345 160.475 ;
        RECT 81.880 160.415 82.200 160.475 ;
        RECT 87.860 160.415 88.180 160.475 ;
        RECT 89.700 160.615 90.020 160.675 ;
        RECT 90.405 160.615 90.695 160.660 ;
        RECT 89.700 160.475 90.695 160.615 ;
        RECT 89.700 160.415 90.020 160.475 ;
        RECT 90.405 160.430 90.695 160.475 ;
        RECT 98.440 160.615 98.760 160.675 ;
        RECT 107.195 160.615 107.485 160.660 ;
        RECT 98.440 160.475 107.485 160.615 ;
        RECT 98.440 160.415 98.760 160.475 ;
        RECT 107.195 160.430 107.485 160.475 ;
        RECT 10.510 159.795 115.850 160.275 ;
        RECT 13.125 159.595 13.415 159.640 ;
        RECT 24.840 159.595 25.160 159.655 ;
        RECT 30.820 159.595 31.140 159.655 ;
        RECT 36.340 159.595 36.660 159.655 ;
        RECT 52.440 159.595 52.760 159.655 ;
        RECT 13.125 159.455 22.770 159.595 ;
        RECT 13.125 159.410 13.415 159.455 ;
        RECT 22.630 159.315 22.770 159.455 ;
        RECT 24.840 159.455 36.660 159.595 ;
        RECT 24.840 159.395 25.160 159.455 ;
        RECT 30.820 159.395 31.140 159.455 ;
        RECT 16.990 159.255 17.280 159.300 ;
        RECT 19.770 159.255 20.060 159.300 ;
        RECT 21.630 159.255 21.920 159.300 ;
        RECT 16.990 159.115 21.920 159.255 ;
        RECT 16.990 159.070 17.280 159.115 ;
        RECT 19.770 159.070 20.060 159.115 ;
        RECT 21.630 159.070 21.920 159.115 ;
        RECT 22.540 159.255 22.860 159.315 ;
        RECT 31.740 159.255 32.060 159.315 ;
        RECT 22.540 159.115 32.060 159.255 ;
        RECT 22.540 159.055 22.860 159.115 ;
        RECT 31.740 159.055 32.060 159.115 ;
        RECT 22.080 158.915 22.400 158.975 ;
        RECT 25.300 158.915 25.620 158.975 ;
        RECT 22.080 158.775 25.620 158.915 ;
        RECT 22.080 158.715 22.400 158.775 ;
        RECT 25.300 158.715 25.620 158.775 ;
        RECT 25.775 158.915 26.065 158.960 ;
        RECT 28.980 158.915 29.300 158.975 ;
        RECT 25.775 158.775 29.300 158.915 ;
        RECT 25.775 158.730 26.065 158.775 ;
        RECT 28.980 158.715 29.300 158.775 ;
        RECT 32.215 158.915 32.505 158.960 ;
        RECT 32.750 158.915 32.890 159.455 ;
        RECT 36.340 159.395 36.660 159.455 ;
        RECT 45.630 159.455 52.760 159.595 ;
        RECT 45.080 159.255 45.400 159.315 ;
        RECT 32.215 158.775 32.890 158.915 ;
        RECT 42.410 159.115 45.400 159.255 ;
        RECT 32.215 158.730 32.505 158.775 ;
        RECT 16.990 158.575 17.280 158.620 ;
        RECT 20.255 158.575 20.545 158.620 ;
        RECT 16.990 158.435 19.525 158.575 ;
        RECT 16.990 158.390 17.280 158.435 ;
        RECT 15.130 158.235 15.420 158.280 ;
        RECT 15.640 158.235 15.960 158.295 ;
        RECT 19.310 158.280 19.525 158.435 ;
        RECT 20.255 158.435 22.770 158.575 ;
        RECT 20.255 158.390 20.545 158.435 ;
        RECT 18.390 158.235 18.680 158.280 ;
        RECT 15.130 158.095 18.680 158.235 ;
        RECT 15.130 158.050 15.420 158.095 ;
        RECT 15.640 158.035 15.960 158.095 ;
        RECT 18.390 158.050 18.680 158.095 ;
        RECT 19.310 158.235 19.600 158.280 ;
        RECT 21.170 158.235 21.460 158.280 ;
        RECT 19.310 158.095 21.460 158.235 ;
        RECT 19.310 158.050 19.600 158.095 ;
        RECT 21.170 158.050 21.460 158.095 ;
        RECT 22.630 157.940 22.770 158.435 ;
        RECT 23.460 158.375 23.780 158.635 ;
        RECT 28.535 158.575 28.825 158.620 ;
        RECT 30.835 158.575 31.125 158.620 ;
        RECT 35.420 158.575 35.740 158.635 ;
        RECT 28.535 158.435 31.125 158.575 ;
        RECT 28.535 158.390 28.825 158.435 ;
        RECT 30.835 158.390 31.125 158.435 ;
        RECT 31.370 158.435 35.740 158.575 ;
        RECT 23.920 158.235 24.240 158.295 ;
        RECT 31.370 158.235 31.510 158.435 ;
        RECT 35.420 158.375 35.740 158.435 ;
        RECT 35.880 158.375 36.200 158.635 ;
        RECT 36.340 158.360 36.630 158.590 ;
        RECT 36.800 158.375 37.120 158.635 ;
        RECT 37.735 158.575 38.025 158.620 ;
        RECT 38.180 158.575 38.500 158.635 ;
        RECT 37.735 158.435 38.500 158.575 ;
        RECT 37.735 158.390 38.025 158.435 ;
        RECT 38.180 158.375 38.500 158.435 ;
        RECT 40.020 158.375 40.340 158.635 ;
        RECT 40.940 158.375 41.260 158.635 ;
        RECT 41.415 158.390 41.705 158.620 ;
        RECT 41.860 158.575 42.180 158.635 ;
        RECT 42.410 158.575 42.550 159.115 ;
        RECT 45.080 159.055 45.400 159.115 ;
        RECT 42.780 158.915 43.100 158.975 ;
        RECT 43.715 158.915 44.005 158.960 ;
        RECT 42.780 158.775 44.005 158.915 ;
        RECT 42.780 158.715 43.100 158.775 ;
        RECT 43.715 158.730 44.005 158.775 ;
        RECT 41.860 158.435 42.550 158.575 ;
        RECT 23.920 158.095 31.510 158.235 ;
        RECT 23.920 158.035 24.240 158.095 ;
        RECT 22.555 157.710 22.845 157.940 ;
        RECT 24.840 157.895 25.160 157.955 ;
        RECT 28.995 157.895 29.285 157.940 ;
        RECT 24.840 157.755 29.285 157.895 ;
        RECT 24.840 157.695 25.160 157.755 ;
        RECT 28.995 157.710 29.285 157.755 ;
        RECT 29.900 157.895 30.220 157.955 ;
        RECT 31.295 157.895 31.585 157.940 ;
        RECT 29.900 157.755 31.585 157.895 ;
        RECT 29.900 157.695 30.220 157.755 ;
        RECT 31.295 157.710 31.585 157.755 ;
        RECT 34.500 157.695 34.820 157.955 ;
        RECT 36.415 157.895 36.555 158.360 ;
        RECT 38.640 158.235 38.960 158.295 ;
        RECT 41.490 158.235 41.630 158.390 ;
        RECT 41.860 158.375 42.180 158.435 ;
        RECT 43.240 158.375 43.560 158.635 ;
        RECT 45.080 158.375 45.400 158.635 ;
        RECT 45.630 158.620 45.770 159.455 ;
        RECT 52.440 159.395 52.760 159.455 ;
        RECT 59.340 159.595 59.660 159.655 ;
        RECT 84.655 159.595 84.945 159.640 ;
        RECT 85.100 159.595 85.420 159.655 ;
        RECT 59.340 159.455 71.070 159.595 ;
        RECT 59.340 159.395 59.660 159.455 ;
        RECT 51.490 159.255 51.780 159.300 ;
        RECT 54.270 159.255 54.560 159.300 ;
        RECT 56.130 159.255 56.420 159.300 ;
        RECT 51.490 159.115 56.420 159.255 ;
        RECT 51.490 159.070 51.780 159.115 ;
        RECT 54.270 159.070 54.560 159.115 ;
        RECT 56.130 159.070 56.420 159.115 ;
        RECT 56.670 159.115 61.870 159.255 ;
        RECT 47.380 158.915 47.700 158.975 ;
        RECT 56.670 158.915 56.810 159.115 ;
        RECT 46.090 158.775 47.700 158.915 ;
        RECT 46.090 158.620 46.230 158.775 ;
        RECT 47.380 158.715 47.700 158.775 ;
        RECT 51.150 158.775 56.810 158.915 ;
        RECT 45.555 158.390 45.845 158.620 ;
        RECT 46.015 158.390 46.305 158.620 ;
        RECT 46.920 158.575 47.240 158.635 ;
        RECT 51.150 158.575 51.290 158.775 ;
        RECT 57.960 158.715 58.280 158.975 ;
        RECT 46.920 158.435 51.290 158.575 ;
        RECT 51.490 158.575 51.780 158.620 ;
        RECT 51.490 158.435 54.025 158.575 ;
        RECT 43.330 158.235 43.470 158.375 ;
        RECT 45.630 158.235 45.770 158.390 ;
        RECT 46.920 158.375 47.240 158.435 ;
        RECT 51.490 158.390 51.780 158.435 ;
        RECT 36.890 158.095 45.770 158.235 ;
        RECT 49.630 158.235 49.920 158.280 ;
        RECT 51.980 158.235 52.300 158.295 ;
        RECT 53.810 158.280 54.025 158.435 ;
        RECT 54.740 158.375 55.060 158.635 ;
        RECT 56.120 158.575 56.440 158.635 ;
        RECT 56.595 158.575 56.885 158.620 ;
        RECT 56.120 158.435 56.885 158.575 ;
        RECT 56.120 158.375 56.440 158.435 ;
        RECT 56.595 158.390 56.885 158.435 ;
        RECT 52.890 158.235 53.180 158.280 ;
        RECT 49.630 158.095 53.180 158.235 ;
        RECT 36.890 157.895 37.030 158.095 ;
        RECT 38.640 158.035 38.960 158.095 ;
        RECT 49.630 158.050 49.920 158.095 ;
        RECT 51.980 158.035 52.300 158.095 ;
        RECT 52.890 158.050 53.180 158.095 ;
        RECT 53.810 158.235 54.100 158.280 ;
        RECT 55.670 158.235 55.960 158.280 ;
        RECT 53.810 158.095 55.960 158.235 ;
        RECT 56.670 158.235 56.810 158.390 ;
        RECT 59.340 158.375 59.660 158.635 ;
        RECT 61.180 158.235 61.500 158.295 ;
        RECT 56.670 158.095 61.500 158.235 ;
        RECT 61.730 158.235 61.870 159.115 ;
        RECT 70.380 158.915 70.700 158.975 ;
        RECT 69.550 158.775 70.700 158.915 ;
        RECT 70.930 158.915 71.070 159.455 ;
        RECT 77.370 159.455 84.410 159.595 ;
        RECT 71.760 159.255 72.080 159.315 ;
        RECT 71.760 159.115 74.290 159.255 ;
        RECT 71.760 159.055 72.080 159.115 ;
        RECT 74.150 158.915 74.290 159.115 ;
        RECT 77.370 158.915 77.510 159.455 ;
        RECT 77.710 159.255 78.000 159.300 ;
        RECT 80.490 159.255 80.780 159.300 ;
        RECT 82.350 159.255 82.640 159.300 ;
        RECT 77.710 159.115 82.640 159.255 ;
        RECT 77.710 159.070 78.000 159.115 ;
        RECT 80.490 159.070 80.780 159.115 ;
        RECT 82.350 159.070 82.640 159.115 ;
        RECT 70.930 158.775 73.140 158.915 ;
        RECT 74.150 158.775 77.510 158.915 ;
        RECT 78.660 158.915 78.980 158.975 ;
        RECT 80.975 158.915 81.265 158.960 ;
        RECT 81.880 158.915 82.200 158.975 ;
        RECT 78.660 158.775 80.730 158.915 ;
        RECT 62.560 158.575 62.880 158.635 ;
        RECT 63.480 158.575 63.800 158.635 ;
        RECT 62.560 158.435 63.800 158.575 ;
        RECT 62.560 158.375 62.880 158.435 ;
        RECT 63.480 158.375 63.800 158.435 ;
        RECT 69.000 158.375 69.320 158.635 ;
        RECT 69.550 158.620 69.690 158.775 ;
        RECT 70.380 158.715 70.700 158.775 ;
        RECT 69.475 158.390 69.765 158.620 ;
        RECT 69.920 158.375 70.240 158.635 ;
        RECT 70.855 158.390 71.145 158.620 ;
        RECT 73.000 158.575 73.140 158.775 ;
        RECT 78.660 158.715 78.980 158.775 ;
        RECT 77.710 158.575 78.000 158.620 ;
        RECT 80.590 158.575 80.730 158.775 ;
        RECT 80.975 158.775 82.200 158.915 ;
        RECT 80.975 158.730 81.265 158.775 ;
        RECT 81.880 158.715 82.200 158.775 ;
        RECT 82.815 158.915 83.105 158.960 ;
        RECT 83.260 158.915 83.580 158.975 ;
        RECT 82.815 158.775 83.580 158.915 ;
        RECT 84.270 158.915 84.410 159.455 ;
        RECT 84.655 159.455 85.420 159.595 ;
        RECT 84.655 159.410 84.945 159.455 ;
        RECT 85.100 159.395 85.420 159.455 ;
        RECT 90.160 159.395 90.480 159.655 ;
        RECT 92.475 159.595 92.765 159.640 ;
        RECT 93.380 159.595 93.700 159.655 ;
        RECT 102.120 159.595 102.440 159.655 ;
        RECT 108.560 159.595 108.880 159.655 ;
        RECT 92.475 159.455 93.700 159.595 ;
        RECT 92.475 159.410 92.765 159.455 ;
        RECT 93.380 159.395 93.700 159.455 ;
        RECT 93.930 159.455 108.880 159.595 ;
        RECT 85.560 159.255 85.880 159.315 ;
        RECT 93.930 159.255 94.070 159.455 ;
        RECT 102.120 159.395 102.440 159.455 ;
        RECT 108.560 159.395 108.880 159.455 ;
        RECT 110.875 159.595 111.165 159.640 ;
        RECT 112.240 159.595 112.560 159.655 ;
        RECT 110.875 159.455 112.560 159.595 ;
        RECT 110.875 159.410 111.165 159.455 ;
        RECT 112.240 159.395 112.560 159.455 ;
        RECT 85.560 159.115 94.070 159.255 ;
        RECT 85.560 159.055 85.880 159.115 ;
        RECT 96.140 159.055 96.460 159.315 ;
        RECT 97.075 159.070 97.365 159.300 ;
        RECT 97.520 159.255 97.840 159.315 ;
        RECT 98.440 159.255 98.760 159.315 ;
        RECT 97.520 159.115 98.760 159.255 ;
        RECT 84.270 158.775 86.250 158.915 ;
        RECT 82.815 158.730 83.105 158.775 ;
        RECT 83.260 158.715 83.580 158.775 ;
        RECT 86.110 158.635 86.250 158.775 ;
        RECT 95.220 158.715 95.540 158.975 ;
        RECT 96.230 158.915 96.370 159.055 ;
        RECT 97.150 158.915 97.290 159.070 ;
        RECT 97.520 159.055 97.840 159.115 ;
        RECT 98.440 159.055 98.760 159.115 ;
        RECT 101.660 159.255 101.980 159.315 ;
        RECT 101.660 159.115 104.190 159.255 ;
        RECT 101.660 159.055 101.980 159.115 ;
        RECT 103.500 158.915 103.820 158.975 ;
        RECT 104.050 158.960 104.190 159.115 ;
        RECT 96.230 158.775 97.290 158.915 ;
        RECT 98.530 158.775 103.820 158.915 ;
        RECT 85.115 158.575 85.405 158.620 ;
        RECT 73.000 158.435 74.750 158.575 ;
        RECT 70.930 158.235 71.070 158.390 ;
        RECT 71.760 158.235 72.080 158.295 ;
        RECT 61.730 158.095 72.080 158.235 ;
        RECT 53.810 158.050 54.100 158.095 ;
        RECT 55.670 158.050 55.960 158.095 ;
        RECT 61.180 158.035 61.500 158.095 ;
        RECT 36.415 157.755 37.030 157.895 ;
        RECT 43.255 157.895 43.545 157.940 ;
        RECT 43.700 157.895 44.020 157.955 ;
        RECT 43.255 157.755 44.020 157.895 ;
        RECT 43.255 157.710 43.545 157.755 ;
        RECT 43.700 157.695 44.020 157.755 ;
        RECT 46.460 157.895 46.780 157.955 ;
        RECT 62.650 157.940 62.790 158.095 ;
        RECT 71.760 158.035 72.080 158.095 ;
        RECT 47.625 157.895 47.915 157.940 ;
        RECT 46.460 157.755 47.915 157.895 ;
        RECT 46.460 157.695 46.780 157.755 ;
        RECT 47.625 157.710 47.915 157.755 ;
        RECT 62.575 157.895 62.865 157.940 ;
        RECT 63.480 157.895 63.800 157.955 ;
        RECT 62.575 157.755 63.800 157.895 ;
        RECT 62.575 157.710 62.865 157.755 ;
        RECT 63.480 157.695 63.800 157.755 ;
        RECT 67.160 157.895 67.480 157.955 ;
        RECT 67.635 157.895 67.925 157.940 ;
        RECT 67.160 157.755 67.925 157.895 ;
        RECT 67.160 157.695 67.480 157.755 ;
        RECT 67.635 157.710 67.925 157.755 ;
        RECT 68.540 157.895 68.860 157.955 ;
        RECT 72.680 157.895 73.000 157.955 ;
        RECT 73.845 157.895 74.135 157.940 ;
        RECT 68.540 157.755 74.135 157.895 ;
        RECT 74.610 157.895 74.750 158.435 ;
        RECT 77.710 158.435 80.245 158.575 ;
        RECT 80.590 158.435 85.405 158.575 ;
        RECT 77.710 158.390 78.000 158.435 ;
        RECT 75.850 158.235 76.140 158.280 ;
        RECT 78.200 158.235 78.520 158.295 ;
        RECT 80.030 158.280 80.245 158.435 ;
        RECT 85.115 158.390 85.405 158.435 ;
        RECT 79.110 158.235 79.400 158.280 ;
        RECT 75.850 158.095 79.400 158.235 ;
        RECT 75.850 158.050 76.140 158.095 ;
        RECT 78.200 158.035 78.520 158.095 ;
        RECT 79.110 158.050 79.400 158.095 ;
        RECT 80.030 158.235 80.320 158.280 ;
        RECT 81.890 158.235 82.180 158.280 ;
        RECT 80.030 158.095 82.180 158.235 ;
        RECT 85.190 158.235 85.330 158.390 ;
        RECT 86.020 158.375 86.340 158.635 ;
        RECT 86.940 158.375 87.260 158.635 ;
        RECT 87.415 158.390 87.705 158.620 ;
        RECT 87.490 158.235 87.630 158.390 ;
        RECT 87.860 158.375 88.180 158.635 ;
        RECT 91.080 158.375 91.400 158.635 ;
        RECT 94.300 158.575 94.620 158.635 ;
        RECT 96.155 158.575 96.445 158.620 ;
        RECT 94.300 158.435 96.445 158.575 ;
        RECT 94.300 158.375 94.620 158.435 ;
        RECT 96.155 158.390 96.445 158.435 ;
        RECT 97.060 158.575 97.380 158.635 ;
        RECT 98.530 158.620 98.670 158.775 ;
        RECT 103.500 158.715 103.820 158.775 ;
        RECT 103.975 158.730 104.265 158.960 ;
        RECT 97.535 158.575 97.825 158.620 ;
        RECT 97.060 158.435 97.825 158.575 ;
        RECT 97.060 158.375 97.380 158.435 ;
        RECT 97.535 158.390 97.825 158.435 ;
        RECT 98.455 158.390 98.745 158.620 ;
        RECT 98.915 158.390 99.205 158.620 ;
        RECT 88.320 158.235 88.640 158.295 ;
        RECT 93.840 158.235 94.160 158.295 ;
        RECT 98.990 158.235 99.130 158.390 ;
        RECT 99.360 158.375 99.680 158.635 ;
        RECT 100.280 158.575 100.600 158.635 ;
        RECT 104.895 158.575 105.185 158.620 ;
        RECT 100.280 158.435 105.185 158.575 ;
        RECT 100.280 158.375 100.600 158.435 ;
        RECT 104.895 158.390 105.185 158.435 ;
        RECT 105.340 158.375 105.660 158.635 ;
        RECT 109.955 158.575 110.245 158.620 ;
        RECT 107.270 158.435 110.245 158.575 ;
        RECT 85.190 158.095 86.250 158.235 ;
        RECT 87.490 158.095 99.130 158.235 ;
        RECT 80.030 158.050 80.320 158.095 ;
        RECT 81.890 158.050 82.180 158.095 ;
        RECT 85.560 157.895 85.880 157.955 ;
        RECT 74.610 157.755 85.880 157.895 ;
        RECT 86.110 157.895 86.250 158.095 ;
        RECT 88.320 158.035 88.640 158.095 ;
        RECT 93.840 158.035 94.160 158.095 ;
        RECT 86.940 157.895 87.260 157.955 ;
        RECT 86.110 157.755 87.260 157.895 ;
        RECT 68.540 157.695 68.860 157.755 ;
        RECT 72.680 157.695 73.000 157.755 ;
        RECT 73.845 157.710 74.135 157.755 ;
        RECT 85.560 157.695 85.880 157.755 ;
        RECT 86.940 157.695 87.260 157.755 ;
        RECT 89.255 157.895 89.545 157.940 ;
        RECT 97.520 157.895 97.840 157.955 ;
        RECT 89.255 157.755 97.840 157.895 ;
        RECT 98.990 157.895 99.130 158.095 ;
        RECT 100.280 157.895 100.600 157.955 ;
        RECT 98.990 157.755 100.600 157.895 ;
        RECT 89.255 157.710 89.545 157.755 ;
        RECT 97.520 157.695 97.840 157.755 ;
        RECT 100.280 157.695 100.600 157.755 ;
        RECT 100.755 157.895 101.045 157.940 ;
        RECT 101.660 157.895 101.980 157.955 ;
        RECT 107.270 157.940 107.410 158.435 ;
        RECT 109.955 158.390 110.245 158.435 ;
        RECT 100.755 157.755 101.980 157.895 ;
        RECT 100.755 157.710 101.045 157.755 ;
        RECT 101.660 157.695 101.980 157.755 ;
        RECT 107.195 157.710 107.485 157.940 ;
        RECT 10.510 157.075 115.850 157.555 ;
        RECT 17.955 156.690 18.245 156.920 ;
        RECT 21.635 156.875 21.925 156.920 ;
        RECT 23.000 156.875 23.320 156.935 ;
        RECT 21.635 156.735 23.320 156.875 ;
        RECT 21.635 156.690 21.925 156.735 ;
        RECT 17.480 156.535 17.800 156.595 ;
        RECT 18.030 156.535 18.170 156.690 ;
        RECT 23.000 156.675 23.320 156.735 ;
        RECT 28.980 156.875 29.300 156.935 ;
        RECT 38.640 156.875 38.960 156.935 ;
        RECT 28.980 156.735 34.270 156.875 ;
        RECT 28.980 156.675 29.300 156.735 ;
        RECT 23.920 156.535 24.240 156.595 ;
        RECT 33.120 156.535 33.440 156.595 ;
        RECT 17.480 156.395 24.240 156.535 ;
        RECT 17.480 156.335 17.800 156.395 ;
        RECT 23.920 156.335 24.240 156.395 ;
        RECT 30.910 156.395 33.440 156.535 ;
        RECT 15.180 156.195 15.500 156.255 ;
        RECT 17.940 156.195 18.260 156.255 ;
        RECT 15.180 156.055 18.260 156.195 ;
        RECT 15.180 155.995 15.500 156.055 ;
        RECT 17.940 155.995 18.260 156.055 ;
        RECT 18.400 155.995 18.720 156.255 ;
        RECT 24.840 155.995 25.160 156.255 ;
        RECT 26.235 156.195 26.525 156.240 ;
        RECT 29.900 156.195 30.220 156.255 ;
        RECT 30.910 156.240 31.050 156.395 ;
        RECT 33.120 156.335 33.440 156.395 ;
        RECT 26.235 156.055 30.220 156.195 ;
        RECT 26.235 156.010 26.525 156.055 ;
        RECT 29.900 155.995 30.220 156.055 ;
        RECT 30.835 156.010 31.125 156.240 ;
        RECT 31.295 156.010 31.585 156.240 ;
        RECT 17.495 155.855 17.785 155.900 ;
        RECT 31.370 155.855 31.510 156.010 ;
        RECT 31.740 155.995 32.060 156.255 ;
        RECT 32.200 156.195 32.520 156.255 ;
        RECT 32.675 156.195 32.965 156.240 ;
        RECT 32.200 156.055 32.965 156.195 ;
        RECT 32.200 155.995 32.520 156.055 ;
        RECT 32.675 156.010 32.965 156.055 ;
        RECT 33.595 156.010 33.885 156.240 ;
        RECT 34.130 156.195 34.270 156.735 ;
        RECT 35.050 156.735 38.960 156.875 ;
        RECT 35.050 156.240 35.190 156.735 ;
        RECT 38.640 156.675 38.960 156.735 ;
        RECT 50.615 156.875 50.905 156.920 ;
        RECT 54.740 156.875 55.060 156.935 ;
        RECT 50.615 156.735 55.060 156.875 ;
        RECT 50.615 156.690 50.905 156.735 ;
        RECT 54.740 156.675 55.060 156.735 ;
        RECT 55.200 156.875 55.520 156.935 ;
        RECT 61.655 156.875 61.945 156.920 ;
        RECT 62.100 156.875 62.420 156.935 ;
        RECT 55.200 156.735 62.420 156.875 ;
        RECT 55.200 156.675 55.520 156.735 ;
        RECT 61.655 156.690 61.945 156.735 ;
        RECT 62.100 156.675 62.420 156.735 ;
        RECT 67.620 156.875 67.940 156.935 ;
        RECT 87.860 156.875 88.180 156.935 ;
        RECT 67.620 156.735 71.070 156.875 ;
        RECT 67.620 156.675 67.940 156.735 ;
        RECT 52.440 156.535 52.760 156.595 ;
        RECT 53.770 156.535 54.060 156.580 ;
        RECT 57.030 156.535 57.320 156.580 ;
        RECT 52.440 156.395 57.320 156.535 ;
        RECT 52.440 156.335 52.760 156.395 ;
        RECT 53.770 156.350 54.060 156.395 ;
        RECT 57.030 156.350 57.320 156.395 ;
        RECT 57.950 156.535 58.240 156.580 ;
        RECT 59.810 156.535 60.100 156.580 ;
        RECT 57.950 156.395 60.100 156.535 ;
        RECT 57.950 156.350 58.240 156.395 ;
        RECT 59.810 156.350 60.100 156.395 ;
        RECT 63.480 156.535 63.800 156.595 ;
        RECT 68.540 156.535 68.860 156.595 ;
        RECT 63.480 156.395 65.090 156.535 ;
        RECT 34.515 156.195 34.805 156.240 ;
        RECT 34.130 156.055 34.805 156.195 ;
        RECT 34.515 156.010 34.805 156.055 ;
        RECT 34.975 156.010 35.265 156.240 ;
        RECT 17.495 155.715 26.450 155.855 ;
        RECT 31.370 155.715 31.970 155.855 ;
        RECT 17.495 155.670 17.785 155.715 ;
        RECT 26.310 155.575 26.450 155.715 ;
        RECT 31.830 155.575 31.970 155.715 ;
        RECT 26.220 155.315 26.540 155.575 ;
        RECT 28.995 155.515 29.285 155.560 ;
        RECT 29.900 155.515 30.220 155.575 ;
        RECT 28.995 155.375 30.220 155.515 ;
        RECT 28.995 155.330 29.285 155.375 ;
        RECT 29.900 155.315 30.220 155.375 ;
        RECT 31.740 155.315 32.060 155.575 ;
        RECT 33.670 155.515 33.810 156.010 ;
        RECT 35.420 155.995 35.740 156.255 ;
        RECT 37.275 156.195 37.565 156.240 ;
        RECT 37.275 156.055 37.950 156.195 ;
        RECT 37.275 156.010 37.565 156.055 ;
        RECT 37.810 155.855 37.950 156.055 ;
        RECT 38.180 155.995 38.500 156.255 ;
        RECT 38.640 155.995 38.960 156.255 ;
        RECT 39.100 156.195 39.420 156.255 ;
        RECT 41.860 156.195 42.180 156.255 ;
        RECT 39.100 156.055 42.180 156.195 ;
        RECT 39.100 155.995 39.420 156.055 ;
        RECT 41.860 155.995 42.180 156.055 ;
        RECT 48.760 156.195 49.080 156.255 ;
        RECT 49.695 156.195 49.985 156.240 ;
        RECT 48.760 156.055 49.985 156.195 ;
        RECT 48.760 155.995 49.080 156.055 ;
        RECT 49.695 156.010 49.985 156.055 ;
        RECT 55.630 156.195 55.920 156.240 ;
        RECT 57.950 156.195 58.165 156.350 ;
        RECT 63.480 156.335 63.800 156.395 ;
        RECT 55.630 156.055 58.165 156.195 ;
        RECT 55.630 156.010 55.920 156.055 ;
        RECT 62.560 155.995 62.880 156.255 ;
        RECT 63.035 156.195 63.325 156.240 ;
        RECT 63.940 156.195 64.260 156.255 ;
        RECT 64.950 156.240 65.090 156.395 ;
        RECT 65.870 156.395 68.860 156.535 ;
        RECT 65.870 156.240 66.010 156.395 ;
        RECT 68.540 156.335 68.860 156.395 ;
        RECT 63.035 156.055 64.260 156.195 ;
        RECT 63.035 156.010 63.325 156.055 ;
        RECT 63.940 155.995 64.260 156.055 ;
        RECT 64.875 156.010 65.165 156.240 ;
        RECT 65.795 156.010 66.085 156.240 ;
        RECT 66.255 156.010 66.545 156.240 ;
        RECT 66.715 156.195 67.005 156.240 ;
        RECT 69.000 156.195 69.320 156.255 ;
        RECT 69.920 156.195 70.240 156.255 ;
        RECT 66.715 156.055 70.240 156.195 ;
        RECT 66.715 156.010 67.005 156.055 ;
        RECT 40.020 155.855 40.340 155.915 ;
        RECT 37.810 155.715 40.340 155.855 ;
        RECT 37.810 155.515 37.950 155.715 ;
        RECT 40.020 155.655 40.340 155.715 ;
        RECT 54.280 155.855 54.600 155.915 ;
        RECT 58.895 155.855 59.185 155.900 ;
        RECT 54.280 155.715 59.185 155.855 ;
        RECT 54.280 155.655 54.600 155.715 ;
        RECT 58.895 155.670 59.185 155.715 ;
        RECT 60.735 155.855 61.025 155.900 ;
        RECT 61.180 155.855 61.500 155.915 ;
        RECT 60.735 155.715 61.500 155.855 ;
        RECT 66.330 155.855 66.470 156.010 ;
        RECT 69.000 155.995 69.320 156.055 ;
        RECT 69.920 155.995 70.240 156.055 ;
        RECT 70.380 155.995 70.700 156.255 ;
        RECT 70.930 156.240 71.070 156.735 ;
        RECT 87.860 156.735 91.310 156.875 ;
        RECT 87.860 156.675 88.180 156.735 ;
        RECT 86.020 156.535 86.340 156.595 ;
        RECT 86.020 156.395 90.850 156.535 ;
        RECT 86.020 156.335 86.340 156.395 ;
        RECT 70.855 156.010 71.145 156.240 ;
        RECT 71.760 155.995 72.080 156.255 ;
        RECT 87.860 156.195 88.180 156.255 ;
        RECT 88.795 156.195 89.085 156.240 ;
        RECT 87.860 156.055 89.085 156.195 ;
        RECT 87.860 155.995 88.180 156.055 ;
        RECT 88.795 156.010 89.085 156.055 ;
        RECT 89.255 156.010 89.545 156.240 ;
        RECT 70.470 155.855 70.610 155.995 ;
        RECT 66.330 155.715 70.610 155.855 ;
        RECT 74.980 155.855 75.300 155.915 ;
        RECT 88.320 155.855 88.640 155.915 ;
        RECT 89.330 155.855 89.470 156.010 ;
        RECT 89.700 155.995 90.020 156.255 ;
        RECT 90.710 156.240 90.850 156.395 ;
        RECT 90.635 156.010 90.925 156.240 ;
        RECT 91.170 156.195 91.310 156.735 ;
        RECT 100.280 156.675 100.600 156.935 ;
        RECT 93.840 156.535 94.160 156.595 ;
        RECT 99.820 156.535 100.140 156.595 ;
        RECT 93.840 156.395 95.910 156.535 ;
        RECT 93.840 156.335 94.160 156.395 ;
        RECT 95.220 156.195 95.540 156.255 ;
        RECT 95.770 156.240 95.910 156.395 ;
        RECT 96.230 156.395 100.140 156.535 ;
        RECT 100.370 156.535 100.510 156.675 ;
        RECT 104.420 156.535 104.740 156.595 ;
        RECT 100.370 156.395 100.970 156.535 ;
        RECT 96.230 156.240 96.370 156.395 ;
        RECT 99.820 156.335 100.140 156.395 ;
        RECT 91.170 156.055 95.540 156.195 ;
        RECT 74.980 155.715 89.470 155.855 ;
        RECT 90.710 155.855 90.850 156.010 ;
        RECT 95.220 155.995 95.540 156.055 ;
        RECT 95.695 156.010 95.985 156.240 ;
        RECT 96.155 156.010 96.445 156.240 ;
        RECT 97.060 155.995 97.380 156.255 ;
        RECT 99.360 156.195 99.680 156.255 ;
        RECT 100.830 156.240 100.970 156.395 ;
        RECT 101.290 156.395 104.740 156.535 ;
        RECT 101.290 156.240 101.430 156.395 ;
        RECT 104.420 156.335 104.740 156.395 ;
        RECT 100.295 156.195 100.585 156.240 ;
        RECT 99.360 156.055 100.585 156.195 ;
        RECT 99.360 155.995 99.680 156.055 ;
        RECT 100.295 156.010 100.585 156.055 ;
        RECT 100.755 156.010 101.045 156.240 ;
        RECT 101.215 156.010 101.505 156.240 ;
        RECT 102.135 156.010 102.425 156.240 ;
        RECT 97.150 155.855 97.290 155.995 ;
        RECT 102.210 155.855 102.350 156.010 ;
        RECT 108.560 155.995 108.880 156.255 ;
        RECT 90.710 155.715 102.350 155.855 ;
        RECT 105.355 155.855 105.645 155.900 ;
        RECT 107.180 155.855 107.500 155.915 ;
        RECT 105.355 155.715 107.500 155.855 ;
        RECT 60.735 155.670 61.025 155.715 ;
        RECT 61.180 155.655 61.500 155.715 ;
        RECT 74.980 155.655 75.300 155.715 ;
        RECT 88.320 155.655 88.640 155.715 ;
        RECT 105.355 155.670 105.645 155.715 ;
        RECT 107.180 155.655 107.500 155.715 ;
        RECT 109.495 155.670 109.785 155.900 ;
        RECT 33.670 155.375 37.950 155.515 ;
        RECT 55.630 155.515 55.920 155.560 ;
        RECT 58.410 155.515 58.700 155.560 ;
        RECT 60.270 155.515 60.560 155.560 ;
        RECT 55.630 155.375 60.560 155.515 ;
        RECT 55.630 155.330 55.920 155.375 ;
        RECT 58.410 155.330 58.700 155.375 ;
        RECT 60.270 155.330 60.560 155.375 ;
        RECT 63.955 155.515 64.245 155.560 ;
        RECT 72.680 155.515 73.000 155.575 ;
        RECT 63.955 155.375 73.000 155.515 ;
        RECT 63.955 155.330 64.245 155.375 ;
        RECT 72.680 155.315 73.000 155.375 ;
        RECT 86.940 155.515 87.260 155.575 ;
        RECT 103.040 155.515 103.360 155.575 ;
        RECT 86.940 155.375 103.360 155.515 ;
        RECT 86.940 155.315 87.260 155.375 ;
        RECT 103.040 155.315 103.360 155.375 ;
        RECT 106.260 155.515 106.580 155.575 ;
        RECT 109.570 155.515 109.710 155.670 ;
        RECT 106.260 155.375 109.710 155.515 ;
        RECT 106.260 155.315 106.580 155.375 ;
        RECT 15.640 154.975 15.960 155.235 ;
        RECT 20.255 155.175 20.545 155.220 ;
        RECT 23.460 155.175 23.780 155.235 ;
        RECT 20.255 155.035 23.780 155.175 ;
        RECT 20.255 154.990 20.545 155.035 ;
        RECT 23.460 154.975 23.780 155.035 ;
        RECT 29.440 154.975 29.760 155.235 ;
        RECT 36.815 155.175 37.105 155.220 ;
        RECT 38.180 155.175 38.500 155.235 ;
        RECT 36.815 155.035 38.500 155.175 ;
        RECT 36.815 154.990 37.105 155.035 ;
        RECT 38.180 154.975 38.500 155.035 ;
        RECT 39.100 155.175 39.420 155.235 ;
        RECT 51.980 155.220 52.300 155.235 ;
        RECT 40.495 155.175 40.785 155.220 ;
        RECT 39.100 155.035 40.785 155.175 ;
        RECT 39.100 154.975 39.420 155.035 ;
        RECT 40.495 154.990 40.785 155.035 ;
        RECT 51.765 154.990 52.300 155.220 ;
        RECT 51.980 154.975 52.300 154.990 ;
        RECT 68.080 154.975 68.400 155.235 ;
        RECT 68.555 155.175 68.845 155.220 ;
        RECT 69.000 155.175 69.320 155.235 ;
        RECT 68.555 155.035 69.320 155.175 ;
        RECT 68.555 154.990 68.845 155.035 ;
        RECT 69.000 154.975 69.320 155.035 ;
        RECT 87.415 155.175 87.705 155.220 ;
        RECT 87.860 155.175 88.180 155.235 ;
        RECT 87.415 155.035 88.180 155.175 ;
        RECT 87.415 154.990 87.705 155.035 ;
        RECT 87.860 154.975 88.180 155.035 ;
        RECT 93.840 154.975 94.160 155.235 ;
        RECT 97.060 155.175 97.380 155.235 ;
        RECT 98.915 155.175 99.205 155.220 ;
        RECT 97.060 155.035 99.205 155.175 ;
        RECT 97.060 154.975 97.380 155.035 ;
        RECT 98.915 154.990 99.205 155.035 ;
        RECT 108.115 155.175 108.405 155.220 ;
        RECT 109.480 155.175 109.800 155.235 ;
        RECT 108.115 155.035 109.800 155.175 ;
        RECT 108.115 154.990 108.405 155.035 ;
        RECT 109.480 154.975 109.800 155.035 ;
        RECT 10.510 154.355 115.850 154.835 ;
        RECT 13.125 154.155 13.415 154.200 ;
        RECT 17.480 154.155 17.800 154.215 ;
        RECT 13.125 154.015 17.800 154.155 ;
        RECT 13.125 153.970 13.415 154.015 ;
        RECT 17.480 153.955 17.800 154.015 ;
        RECT 26.220 154.155 26.540 154.215 ;
        RECT 30.820 154.155 31.140 154.215 ;
        RECT 26.220 154.015 31.140 154.155 ;
        RECT 26.220 153.955 26.540 154.015 ;
        RECT 30.820 153.955 31.140 154.015 ;
        RECT 31.740 154.155 32.060 154.215 ;
        RECT 39.560 154.155 39.880 154.215 ;
        RECT 31.740 154.015 39.880 154.155 ;
        RECT 31.740 153.955 32.060 154.015 ;
        RECT 39.560 153.955 39.880 154.015 ;
        RECT 48.760 153.955 49.080 154.215 ;
        RECT 64.875 154.155 65.165 154.200 ;
        RECT 70.380 154.155 70.700 154.215 ;
        RECT 64.875 154.015 70.700 154.155 ;
        RECT 64.875 153.970 65.165 154.015 ;
        RECT 70.380 153.955 70.700 154.015 ;
        RECT 95.220 154.155 95.540 154.215 ;
        RECT 99.360 154.155 99.680 154.215 ;
        RECT 95.220 154.015 99.680 154.155 ;
        RECT 95.220 153.955 95.540 154.015 ;
        RECT 99.360 153.955 99.680 154.015 ;
        RECT 107.180 153.955 107.500 154.215 ;
        RECT 16.990 153.815 17.280 153.860 ;
        RECT 19.770 153.815 20.060 153.860 ;
        RECT 21.630 153.815 21.920 153.860 ;
        RECT 16.990 153.675 21.920 153.815 ;
        RECT 16.990 153.630 17.280 153.675 ;
        RECT 19.770 153.630 20.060 153.675 ;
        RECT 21.630 153.630 21.920 153.675 ;
        RECT 22.555 153.630 22.845 153.860 ;
        RECT 20.255 153.475 20.545 153.520 ;
        RECT 22.630 153.475 22.770 153.630 ;
        RECT 30.910 153.520 31.050 153.955 ;
        RECT 55.200 153.815 55.520 153.875 ;
        RECT 61.655 153.815 61.945 153.860 ;
        RECT 55.200 153.675 61.945 153.815 ;
        RECT 55.200 153.615 55.520 153.675 ;
        RECT 61.655 153.630 61.945 153.675 ;
        RECT 62.100 153.815 62.420 153.875 ;
        RECT 65.780 153.815 66.100 153.875 ;
        RECT 62.100 153.675 66.100 153.815 ;
        RECT 62.100 153.615 62.420 153.675 ;
        RECT 65.780 153.615 66.100 153.675 ;
        RECT 66.240 153.815 66.560 153.875 ;
        RECT 66.240 153.675 67.850 153.815 ;
        RECT 66.240 153.615 66.560 153.675 ;
        RECT 20.255 153.335 22.770 153.475 ;
        RECT 20.255 153.290 20.545 153.335 ;
        RECT 30.835 153.290 31.125 153.520 ;
        RECT 46.460 153.475 46.780 153.535 ;
        RECT 51.075 153.475 51.365 153.520 ;
        RECT 46.460 153.335 51.365 153.475 ;
        RECT 46.460 153.275 46.780 153.335 ;
        RECT 51.075 153.290 51.365 153.335 ;
        RECT 51.520 153.475 51.840 153.535 ;
        RECT 55.675 153.475 55.965 153.520 ;
        RECT 63.480 153.475 63.800 153.535 ;
        RECT 67.710 153.520 67.850 153.675 ;
        RECT 66.715 153.475 67.005 153.520 ;
        RECT 51.520 153.335 55.965 153.475 ;
        RECT 51.520 153.275 51.840 153.335 ;
        RECT 55.675 153.290 55.965 153.335 ;
        RECT 62.650 153.335 67.005 153.475 ;
        RECT 16.990 153.135 17.280 153.180 ;
        RECT 16.990 152.995 19.525 153.135 ;
        RECT 16.990 152.950 17.280 152.995 ;
        RECT 15.130 152.795 15.420 152.840 ;
        RECT 15.640 152.795 15.960 152.855 ;
        RECT 19.310 152.840 19.525 152.995 ;
        RECT 22.080 152.935 22.400 153.195 ;
        RECT 23.460 152.935 23.780 153.195 ;
        RECT 29.900 152.935 30.220 153.195 ;
        RECT 57.960 152.935 58.280 153.195 ;
        RECT 62.650 153.180 62.790 153.335 ;
        RECT 63.480 153.275 63.800 153.335 ;
        RECT 66.715 153.290 67.005 153.335 ;
        RECT 67.635 153.290 67.925 153.520 ;
        RECT 74.520 153.475 74.840 153.535 ;
        RECT 99.820 153.475 100.140 153.535 ;
        RECT 71.390 153.335 74.840 153.475 ;
        RECT 60.735 152.950 61.025 153.180 ;
        RECT 62.575 152.950 62.865 153.180 ;
        RECT 65.780 153.135 66.100 153.195 ;
        RECT 66.255 153.135 66.545 153.180 ;
        RECT 68.095 153.135 68.385 153.180 ;
        RECT 65.780 152.995 66.545 153.135 ;
        RECT 18.390 152.795 18.680 152.840 ;
        RECT 15.130 152.655 18.680 152.795 ;
        RECT 15.130 152.610 15.420 152.655 ;
        RECT 15.640 152.595 15.960 152.655 ;
        RECT 18.390 152.610 18.680 152.655 ;
        RECT 19.310 152.795 19.600 152.840 ;
        RECT 21.170 152.795 21.460 152.840 ;
        RECT 19.310 152.655 21.460 152.795 ;
        RECT 19.310 152.610 19.600 152.655 ;
        RECT 21.170 152.610 21.460 152.655 ;
        RECT 25.760 152.795 26.080 152.855 ;
        RECT 30.375 152.795 30.665 152.840 ;
        RECT 30.820 152.795 31.140 152.855 ;
        RECT 55.215 152.795 55.505 152.840 ;
        RECT 25.760 152.655 31.140 152.795 ;
        RECT 25.760 152.595 26.080 152.655 ;
        RECT 30.375 152.610 30.665 152.655 ;
        RECT 30.820 152.595 31.140 152.655 ;
        RECT 52.070 152.655 55.505 152.795 ;
        RECT 60.810 152.795 60.950 152.950 ;
        RECT 65.780 152.935 66.100 152.995 ;
        RECT 66.255 152.950 66.545 152.995 ;
        RECT 66.790 152.995 68.385 153.135 ;
        RECT 66.790 152.795 66.930 152.995 ;
        RECT 68.095 152.950 68.385 152.995 ;
        RECT 69.920 153.135 70.240 153.195 ;
        RECT 70.395 153.135 70.685 153.180 ;
        RECT 69.920 152.995 70.685 153.135 ;
        RECT 69.920 152.935 70.240 152.995 ;
        RECT 70.395 152.950 70.685 152.995 ;
        RECT 70.840 152.935 71.160 153.195 ;
        RECT 71.390 153.180 71.530 153.335 ;
        RECT 74.520 153.275 74.840 153.335 ;
        RECT 97.610 153.335 100.140 153.475 ;
        RECT 71.315 152.950 71.605 153.180 ;
        RECT 71.760 153.135 72.080 153.195 ;
        RECT 72.235 153.135 72.525 153.180 ;
        RECT 71.760 152.995 72.525 153.135 ;
        RECT 71.760 152.935 72.080 152.995 ;
        RECT 72.235 152.950 72.525 152.995 ;
        RECT 82.355 152.950 82.645 153.180 ;
        RECT 60.810 152.655 66.930 152.795 ;
        RECT 67.620 152.795 67.940 152.855 ;
        RECT 69.015 152.795 69.305 152.840 ;
        RECT 67.620 152.655 69.305 152.795 ;
        RECT 82.430 152.795 82.570 152.950 ;
        RECT 82.800 152.935 83.120 153.195 ;
        RECT 86.940 153.135 87.260 153.195 ;
        RECT 88.335 153.135 88.625 153.180 ;
        RECT 86.940 152.995 88.625 153.135 ;
        RECT 86.940 152.935 87.260 152.995 ;
        RECT 88.335 152.950 88.625 152.995 ;
        RECT 95.220 153.135 95.540 153.195 ;
        RECT 97.610 153.180 97.750 153.335 ;
        RECT 99.820 153.275 100.140 153.335 ;
        RECT 104.420 153.275 104.740 153.535 ;
        RECT 97.075 153.135 97.365 153.180 ;
        RECT 95.220 152.995 97.365 153.135 ;
        RECT 95.220 152.935 95.540 152.995 ;
        RECT 97.075 152.950 97.365 152.995 ;
        RECT 97.535 152.950 97.825 153.180 ;
        RECT 97.995 153.135 98.285 153.180 ;
        RECT 98.440 153.135 98.760 153.195 ;
        RECT 97.995 152.995 98.760 153.135 ;
        RECT 97.995 152.950 98.285 152.995 ;
        RECT 98.440 152.935 98.760 152.995 ;
        RECT 98.915 152.950 99.205 153.180 ;
        RECT 83.260 152.795 83.580 152.855 ;
        RECT 96.600 152.795 96.920 152.855 ;
        RECT 98.990 152.795 99.130 152.950 ;
        RECT 100.280 152.935 100.600 153.195 ;
        RECT 109.480 152.935 109.800 153.195 ;
        RECT 106.260 152.795 106.580 152.855 ;
        RECT 82.430 152.655 96.370 152.795 ;
        RECT 52.070 152.515 52.210 152.655 ;
        RECT 55.215 152.610 55.505 152.655 ;
        RECT 62.650 152.515 62.790 152.655 ;
        RECT 67.620 152.595 67.940 152.655 ;
        RECT 69.015 152.610 69.305 152.655 ;
        RECT 83.260 152.595 83.580 152.655 ;
        RECT 28.075 152.455 28.365 152.500 ;
        RECT 28.980 152.455 29.300 152.515 ;
        RECT 28.075 152.315 29.300 152.455 ;
        RECT 28.075 152.270 28.365 152.315 ;
        RECT 28.980 152.255 29.300 152.315 ;
        RECT 48.760 152.455 49.080 152.515 ;
        RECT 50.615 152.455 50.905 152.500 ;
        RECT 51.980 152.455 52.300 152.515 ;
        RECT 48.760 152.315 52.300 152.455 ;
        RECT 48.760 152.255 49.080 152.315 ;
        RECT 50.615 152.270 50.905 152.315 ;
        RECT 51.980 152.255 52.300 152.315 ;
        RECT 52.900 152.255 53.220 152.515 ;
        RECT 54.755 152.455 55.045 152.500 ;
        RECT 56.120 152.455 56.440 152.515 ;
        RECT 54.755 152.315 56.440 152.455 ;
        RECT 54.755 152.270 55.045 152.315 ;
        RECT 56.120 152.255 56.440 152.315 ;
        RECT 58.880 152.255 59.200 152.515 ;
        RECT 59.800 152.255 60.120 152.515 ;
        RECT 62.560 152.255 62.880 152.515 ;
        RECT 63.020 152.455 63.340 152.515 ;
        RECT 66.240 152.455 66.560 152.515 ;
        RECT 63.020 152.315 66.560 152.455 ;
        RECT 63.020 152.255 63.340 152.315 ;
        RECT 66.240 152.255 66.560 152.315 ;
        RECT 68.540 152.255 68.860 152.515 ;
        RECT 81.880 152.255 82.200 152.515 ;
        RECT 83.735 152.455 84.025 152.500 ;
        RECT 84.640 152.455 84.960 152.515 ;
        RECT 83.735 152.315 84.960 152.455 ;
        RECT 83.735 152.270 84.025 152.315 ;
        RECT 84.640 152.255 84.960 152.315 ;
        RECT 88.780 152.255 89.100 152.515 ;
        RECT 94.300 152.455 94.620 152.515 ;
        RECT 95.695 152.455 95.985 152.500 ;
        RECT 94.300 152.315 95.985 152.455 ;
        RECT 96.230 152.455 96.370 152.655 ;
        RECT 96.600 152.655 99.130 152.795 ;
        RECT 99.450 152.655 106.580 152.795 ;
        RECT 96.600 152.595 96.920 152.655 ;
        RECT 99.450 152.455 99.590 152.655 ;
        RECT 106.260 152.595 106.580 152.655 ;
        RECT 96.230 152.315 99.590 152.455 ;
        RECT 99.820 152.455 100.140 152.515 ;
        RECT 100.740 152.455 101.060 152.515 ;
        RECT 99.820 152.315 101.060 152.455 ;
        RECT 94.300 152.255 94.620 152.315 ;
        RECT 95.695 152.270 95.985 152.315 ;
        RECT 99.820 152.255 100.140 152.315 ;
        RECT 100.740 152.255 101.060 152.315 ;
        RECT 102.580 152.455 102.900 152.515 ;
        RECT 103.055 152.455 103.345 152.500 ;
        RECT 104.895 152.455 105.185 152.500 ;
        RECT 102.580 152.315 105.185 152.455 ;
        RECT 102.580 152.255 102.900 152.315 ;
        RECT 103.055 152.270 103.345 152.315 ;
        RECT 104.895 152.270 105.185 152.315 ;
        RECT 105.340 152.255 105.660 152.515 ;
        RECT 110.415 152.455 110.705 152.500 ;
        RECT 112.240 152.455 112.560 152.515 ;
        RECT 110.415 152.315 112.560 152.455 ;
        RECT 110.415 152.270 110.705 152.315 ;
        RECT 112.240 152.255 112.560 152.315 ;
        RECT 10.510 151.635 115.850 152.115 ;
        RECT 15.180 151.435 15.500 151.495 ;
        RECT 22.540 151.435 22.860 151.495 ;
        RECT 30.820 151.435 31.140 151.495 ;
        RECT 43.255 151.435 43.545 151.480 ;
        RECT 47.380 151.435 47.700 151.495 ;
        RECT 15.180 151.295 24.150 151.435 ;
        RECT 15.180 151.235 15.500 151.295 ;
        RECT 22.540 151.235 22.860 151.295 ;
        RECT 17.940 151.095 18.260 151.155 ;
        RECT 18.875 151.095 19.165 151.140 ;
        RECT 17.940 150.955 19.165 151.095 ;
        RECT 17.940 150.895 18.260 150.955 ;
        RECT 18.875 150.910 19.165 150.955 ;
        RECT 18.400 150.755 18.720 150.815 ;
        RECT 23.000 150.755 23.320 150.815 ;
        RECT 24.010 150.800 24.150 151.295 ;
        RECT 30.820 151.295 37.950 151.435 ;
        RECT 30.820 151.235 31.140 151.295 ;
        RECT 24.395 151.095 24.685 151.140 ;
        RECT 28.010 151.095 28.300 151.140 ;
        RECT 31.270 151.095 31.560 151.140 ;
        RECT 24.395 150.955 31.560 151.095 ;
        RECT 24.395 150.910 24.685 150.955 ;
        RECT 28.010 150.910 28.300 150.955 ;
        RECT 31.270 150.910 31.560 150.955 ;
        RECT 32.190 151.095 32.480 151.140 ;
        RECT 34.050 151.095 34.340 151.140 ;
        RECT 32.190 150.955 34.340 151.095 ;
        RECT 32.190 150.910 32.480 150.955 ;
        RECT 34.050 150.910 34.340 150.955 ;
        RECT 25.760 150.800 26.080 150.815 ;
        RECT 18.400 150.615 23.320 150.755 ;
        RECT 18.400 150.555 18.720 150.615 ;
        RECT 23.000 150.555 23.320 150.615 ;
        RECT 23.935 150.570 24.225 150.800 ;
        RECT 25.760 150.570 26.295 150.800 ;
        RECT 29.870 150.755 30.160 150.800 ;
        RECT 32.190 150.755 32.405 150.910 ;
        RECT 29.870 150.615 32.405 150.755 ;
        RECT 29.870 150.570 30.160 150.615 ;
        RECT 25.760 150.555 26.080 150.570 ;
        RECT 33.120 150.555 33.440 150.815 ;
        RECT 36.800 150.555 37.120 150.815 ;
        RECT 37.810 150.800 37.950 151.295 ;
        RECT 43.255 151.295 47.700 151.435 ;
        RECT 43.255 151.250 43.545 151.295 ;
        RECT 47.380 151.235 47.700 151.295 ;
        RECT 52.440 151.235 52.760 151.495 ;
        RECT 54.280 151.235 54.600 151.495 ;
        RECT 99.820 151.435 100.140 151.495 ;
        RECT 95.770 151.295 100.140 151.435 ;
        RECT 38.180 151.095 38.500 151.155 ;
        RECT 45.555 151.095 45.845 151.140 ;
        RECT 46.475 151.095 46.765 151.140 ;
        RECT 38.180 150.955 42.090 151.095 ;
        RECT 38.180 150.895 38.500 150.955 ;
        RECT 37.275 150.570 37.565 150.800 ;
        RECT 37.735 150.570 38.025 150.800 ;
        RECT 38.655 150.755 38.945 150.800 ;
        RECT 40.020 150.755 40.340 150.815 ;
        RECT 41.950 150.800 42.090 150.955 ;
        RECT 45.555 150.955 46.765 151.095 ;
        RECT 45.555 150.910 45.845 150.955 ;
        RECT 46.475 150.910 46.765 150.955 ;
        RECT 49.220 151.095 49.540 151.155 ;
        RECT 51.520 151.095 51.840 151.155 ;
        RECT 63.955 151.095 64.245 151.140 ;
        RECT 49.220 150.955 64.245 151.095 ;
        RECT 49.220 150.895 49.540 150.955 ;
        RECT 51.520 150.895 51.840 150.955 ;
        RECT 63.955 150.910 64.245 150.955 ;
        RECT 65.795 151.095 66.085 151.140 ;
        RECT 68.540 151.095 68.860 151.155 ;
        RECT 71.315 151.095 71.605 151.140 ;
        RECT 65.795 150.955 71.605 151.095 ;
        RECT 65.795 150.910 66.085 150.955 ;
        RECT 68.540 150.895 68.860 150.955 ;
        RECT 71.315 150.910 71.605 150.955 ;
        RECT 79.530 151.095 79.820 151.140 ;
        RECT 81.880 151.095 82.200 151.155 ;
        RECT 82.790 151.095 83.080 151.140 ;
        RECT 79.530 150.955 83.080 151.095 ;
        RECT 79.530 150.910 79.820 150.955 ;
        RECT 81.880 150.895 82.200 150.955 ;
        RECT 82.790 150.910 83.080 150.955 ;
        RECT 83.710 151.095 84.000 151.140 ;
        RECT 85.570 151.095 85.860 151.140 ;
        RECT 83.710 150.955 85.860 151.095 ;
        RECT 83.710 150.910 84.000 150.955 ;
        RECT 85.570 150.910 85.860 150.955 ;
        RECT 88.435 151.095 88.725 151.140 ;
        RECT 91.675 151.095 92.325 151.140 ;
        RECT 88.435 150.955 92.325 151.095 ;
        RECT 88.435 150.910 89.025 150.955 ;
        RECT 91.675 150.910 92.325 150.955 ;
        RECT 92.920 151.095 93.240 151.155 ;
        RECT 94.315 151.095 94.605 151.140 ;
        RECT 92.920 150.955 94.605 151.095 ;
        RECT 38.655 150.615 40.340 150.755 ;
        RECT 38.655 150.570 38.945 150.615 ;
        RECT 17.955 150.230 18.245 150.460 ;
        RECT 22.080 150.415 22.400 150.475 ;
        RECT 34.975 150.415 35.265 150.460 ;
        RECT 22.080 150.275 35.265 150.415 ;
        RECT 18.030 150.075 18.170 150.230 ;
        RECT 22.080 150.215 22.400 150.275 ;
        RECT 34.975 150.230 35.265 150.275 ;
        RECT 26.220 150.075 26.540 150.135 ;
        RECT 18.030 149.935 26.540 150.075 ;
        RECT 26.220 149.875 26.540 149.935 ;
        RECT 29.870 150.075 30.160 150.120 ;
        RECT 32.650 150.075 32.940 150.120 ;
        RECT 34.510 150.075 34.800 150.120 ;
        RECT 29.870 149.935 34.800 150.075 ;
        RECT 37.350 150.075 37.490 150.570 ;
        RECT 40.020 150.555 40.340 150.615 ;
        RECT 40.495 150.755 40.785 150.800 ;
        RECT 40.495 150.615 41.630 150.755 ;
        RECT 40.495 150.570 40.785 150.615 ;
        RECT 38.180 150.415 38.500 150.475 ;
        RECT 40.955 150.415 41.245 150.460 ;
        RECT 38.180 150.275 41.245 150.415 ;
        RECT 41.490 150.415 41.630 150.615 ;
        RECT 41.875 150.570 42.165 150.800 ;
        RECT 44.160 150.555 44.480 150.815 ;
        RECT 44.620 150.555 44.940 150.815 ;
        RECT 47.855 150.570 48.145 150.800 ;
        RECT 45.080 150.415 45.400 150.475 ;
        RECT 41.490 150.275 45.400 150.415 ;
        RECT 38.180 150.215 38.500 150.275 ;
        RECT 40.955 150.230 41.245 150.275 ;
        RECT 45.080 150.215 45.400 150.275 ;
        RECT 45.540 150.415 45.860 150.475 ;
        RECT 47.930 150.415 48.070 150.570 ;
        RECT 48.300 150.555 48.620 150.815 ;
        RECT 48.760 150.555 49.080 150.815 ;
        RECT 49.695 150.570 49.985 150.800 ;
        RECT 51.995 150.755 52.285 150.800 ;
        RECT 52.440 150.755 52.760 150.815 ;
        RECT 51.995 150.615 52.760 150.755 ;
        RECT 51.995 150.570 52.285 150.615 ;
        RECT 49.770 150.415 49.910 150.570 ;
        RECT 52.440 150.555 52.760 150.615 ;
        RECT 52.900 150.755 53.220 150.815 ;
        RECT 53.375 150.755 53.665 150.800 ;
        RECT 52.900 150.615 53.665 150.755 ;
        RECT 52.900 150.555 53.220 150.615 ;
        RECT 53.375 150.570 53.665 150.615 ;
        RECT 63.480 150.555 63.800 150.815 ;
        RECT 69.000 150.555 69.320 150.815 ;
        RECT 70.380 150.555 70.700 150.815 ;
        RECT 81.390 150.755 81.680 150.800 ;
        RECT 83.710 150.755 83.925 150.910 ;
        RECT 88.735 150.815 89.025 150.910 ;
        RECT 92.920 150.895 93.240 150.955 ;
        RECT 94.315 150.910 94.605 150.955 ;
        RECT 81.390 150.615 83.925 150.755 ;
        RECT 81.390 150.570 81.680 150.615 ;
        RECT 84.640 150.555 84.960 150.815 ;
        RECT 86.480 150.555 86.800 150.815 ;
        RECT 88.735 150.595 89.100 150.815 ;
        RECT 95.770 150.800 95.910 151.295 ;
        RECT 99.820 151.235 100.140 151.295 ;
        RECT 100.280 151.435 100.600 151.495 ;
        RECT 104.895 151.435 105.185 151.480 ;
        RECT 100.280 151.295 105.185 151.435 ;
        RECT 100.280 151.235 100.600 151.295 ;
        RECT 98.455 151.095 98.745 151.140 ;
        RECT 98.915 151.095 99.205 151.140 ;
        RECT 98.455 150.955 99.205 151.095 ;
        RECT 98.455 150.910 98.745 150.955 ;
        RECT 98.915 150.910 99.205 150.955 ;
        RECT 101.290 150.830 101.430 151.295 ;
        RECT 104.895 151.250 105.185 151.295 ;
        RECT 103.975 151.095 104.265 151.140 ;
        RECT 106.375 151.095 106.665 151.140 ;
        RECT 109.615 151.095 110.265 151.140 ;
        RECT 103.975 150.955 110.265 151.095 ;
        RECT 103.975 150.910 104.265 150.955 ;
        RECT 106.375 150.910 106.965 150.955 ;
        RECT 109.615 150.910 110.265 150.955 ;
        RECT 88.780 150.555 89.100 150.595 ;
        RECT 89.815 150.755 90.105 150.800 ;
        RECT 93.395 150.755 93.685 150.800 ;
        RECT 95.230 150.755 95.520 150.800 ;
        RECT 89.815 150.615 95.520 150.755 ;
        RECT 89.815 150.570 90.105 150.615 ;
        RECT 93.395 150.570 93.685 150.615 ;
        RECT 95.230 150.570 95.520 150.615 ;
        RECT 95.695 150.570 95.985 150.800 ;
        RECT 97.060 150.555 97.380 150.815 ;
        RECT 99.820 150.800 100.140 150.815 ;
        RECT 99.820 150.570 100.355 150.800 ;
        RECT 100.755 150.570 101.045 150.800 ;
        RECT 101.215 150.600 101.505 150.830 ;
        RECT 99.820 150.555 100.140 150.570 ;
        RECT 69.935 150.415 70.225 150.460 ;
        RECT 72.220 150.415 72.540 150.475 ;
        RECT 45.540 150.275 48.990 150.415 ;
        RECT 49.770 150.275 52.210 150.415 ;
        RECT 45.540 150.215 45.860 150.275 ;
        RECT 48.850 150.135 48.990 150.275 ;
        RECT 52.070 150.135 52.210 150.275 ;
        RECT 69.935 150.275 72.540 150.415 ;
        RECT 69.935 150.230 70.225 150.275 ;
        RECT 72.220 150.215 72.540 150.275 ;
        RECT 97.995 150.415 98.285 150.460 ;
        RECT 97.995 150.275 99.590 150.415 ;
        RECT 97.995 150.230 98.285 150.275 ;
        RECT 39.560 150.075 39.880 150.135 ;
        RECT 37.350 149.935 39.880 150.075 ;
        RECT 29.870 149.890 30.160 149.935 ;
        RECT 32.650 149.890 32.940 149.935 ;
        RECT 34.510 149.890 34.800 149.935 ;
        RECT 39.560 149.875 39.880 149.935 ;
        RECT 41.030 149.935 45.310 150.075 ;
        RECT 41.030 149.795 41.170 149.935 ;
        RECT 18.400 149.735 18.720 149.795 ;
        RECT 20.715 149.735 21.005 149.780 ;
        RECT 18.400 149.595 21.005 149.735 ;
        RECT 18.400 149.535 18.720 149.595 ;
        RECT 20.715 149.550 21.005 149.595 ;
        RECT 34.040 149.735 34.360 149.795 ;
        RECT 35.435 149.735 35.725 149.780 ;
        RECT 34.040 149.595 35.725 149.735 ;
        RECT 34.040 149.535 34.360 149.595 ;
        RECT 35.435 149.550 35.725 149.595 ;
        RECT 40.940 149.535 41.260 149.795 ;
        RECT 41.860 149.535 42.180 149.795 ;
        RECT 42.795 149.735 43.085 149.780 ;
        RECT 44.620 149.735 44.940 149.795 ;
        RECT 45.170 149.780 45.310 149.935 ;
        RECT 48.760 149.875 49.080 150.135 ;
        RECT 51.980 150.075 52.300 150.135 ;
        RECT 59.800 150.075 60.120 150.135 ;
        RECT 51.980 149.935 60.120 150.075 ;
        RECT 51.980 149.875 52.300 149.935 ;
        RECT 59.800 149.875 60.120 149.935 ;
        RECT 81.390 150.075 81.680 150.120 ;
        RECT 84.170 150.075 84.460 150.120 ;
        RECT 86.030 150.075 86.320 150.120 ;
        RECT 81.390 149.935 86.320 150.075 ;
        RECT 81.390 149.890 81.680 149.935 ;
        RECT 84.170 149.890 84.460 149.935 ;
        RECT 86.030 149.890 86.320 149.935 ;
        RECT 89.815 150.075 90.105 150.120 ;
        RECT 92.935 150.075 93.225 150.120 ;
        RECT 94.825 150.075 95.115 150.120 ;
        RECT 89.815 149.935 95.115 150.075 ;
        RECT 89.815 149.890 90.105 149.935 ;
        RECT 92.935 149.890 93.225 149.935 ;
        RECT 94.825 149.890 95.115 149.935 ;
        RECT 96.600 150.075 96.920 150.135 ;
        RECT 98.900 150.075 99.220 150.135 ;
        RECT 96.600 149.935 99.220 150.075 ;
        RECT 99.450 150.075 99.590 150.275 ;
        RECT 100.830 150.135 100.970 150.570 ;
        RECT 102.120 150.555 102.440 150.815 ;
        RECT 103.040 150.755 103.360 150.815 ;
        RECT 103.515 150.755 103.805 150.800 ;
        RECT 103.040 150.615 103.805 150.755 ;
        RECT 103.040 150.555 103.360 150.615 ;
        RECT 103.515 150.570 103.805 150.615 ;
        RECT 106.675 150.595 106.965 150.910 ;
        RECT 112.240 150.895 112.560 151.155 ;
        RECT 107.755 150.755 108.045 150.800 ;
        RECT 111.335 150.755 111.625 150.800 ;
        RECT 113.170 150.755 113.460 150.800 ;
        RECT 107.755 150.615 113.460 150.755 ;
        RECT 107.755 150.570 108.045 150.615 ;
        RECT 111.335 150.570 111.625 150.615 ;
        RECT 113.170 150.570 113.460 150.615 ;
        RECT 113.635 150.415 113.925 150.460 ;
        RECT 101.290 150.275 113.925 150.415 ;
        RECT 101.290 150.135 101.430 150.275 ;
        RECT 113.635 150.230 113.925 150.275 ;
        RECT 99.450 149.935 100.050 150.075 ;
        RECT 96.600 149.875 96.920 149.935 ;
        RECT 98.900 149.875 99.220 149.935 ;
        RECT 42.795 149.595 44.940 149.735 ;
        RECT 42.795 149.550 43.085 149.595 ;
        RECT 44.620 149.535 44.940 149.595 ;
        RECT 45.095 149.550 45.385 149.780 ;
        RECT 57.040 149.535 57.360 149.795 ;
        RECT 68.095 149.735 68.385 149.780 ;
        RECT 68.540 149.735 68.860 149.795 ;
        RECT 68.095 149.595 68.860 149.735 ;
        RECT 68.095 149.550 68.385 149.595 ;
        RECT 68.540 149.535 68.860 149.595 ;
        RECT 69.920 149.535 70.240 149.795 ;
        RECT 72.695 149.735 72.985 149.780 ;
        RECT 73.600 149.735 73.920 149.795 ;
        RECT 72.695 149.595 73.920 149.735 ;
        RECT 72.695 149.550 72.985 149.595 ;
        RECT 73.600 149.535 73.920 149.595 ;
        RECT 77.525 149.735 77.815 149.780 ;
        RECT 79.120 149.735 79.440 149.795 ;
        RECT 77.525 149.595 79.440 149.735 ;
        RECT 77.525 149.550 77.815 149.595 ;
        RECT 79.120 149.535 79.440 149.595 ;
        RECT 86.940 149.535 87.260 149.795 ;
        RECT 96.155 149.735 96.445 149.780 ;
        RECT 97.980 149.735 98.300 149.795 ;
        RECT 96.155 149.595 98.300 149.735 ;
        RECT 96.155 149.550 96.445 149.595 ;
        RECT 97.980 149.535 98.300 149.595 ;
        RECT 98.455 149.735 98.745 149.780 ;
        RECT 99.360 149.735 99.680 149.795 ;
        RECT 98.455 149.595 99.680 149.735 ;
        RECT 99.910 149.735 100.050 149.935 ;
        RECT 100.740 149.875 101.060 150.135 ;
        RECT 101.200 149.875 101.520 150.135 ;
        RECT 107.755 150.075 108.045 150.120 ;
        RECT 110.875 150.075 111.165 150.120 ;
        RECT 112.765 150.075 113.055 150.120 ;
        RECT 107.755 149.935 113.055 150.075 ;
        RECT 107.755 149.890 108.045 149.935 ;
        RECT 110.875 149.890 111.165 149.935 ;
        RECT 112.765 149.890 113.055 149.935 ;
        RECT 104.880 149.735 105.200 149.795 ;
        RECT 99.910 149.595 105.200 149.735 ;
        RECT 98.455 149.550 98.745 149.595 ;
        RECT 99.360 149.535 99.680 149.595 ;
        RECT 104.880 149.535 105.200 149.595 ;
        RECT 10.510 148.915 115.850 149.395 ;
        RECT 18.860 148.715 19.180 148.775 ;
        RECT 28.520 148.715 28.840 148.775 ;
        RECT 16.650 148.575 19.180 148.715 ;
        RECT 13.125 148.035 13.415 148.080 ;
        RECT 16.650 148.035 16.790 148.575 ;
        RECT 18.860 148.515 19.180 148.575 ;
        RECT 24.700 148.575 28.840 148.715 ;
        RECT 16.990 148.375 17.280 148.420 ;
        RECT 19.770 148.375 20.060 148.420 ;
        RECT 21.630 148.375 21.920 148.420 ;
        RECT 16.990 148.235 21.920 148.375 ;
        RECT 16.990 148.190 17.280 148.235 ;
        RECT 19.770 148.190 20.060 148.235 ;
        RECT 21.630 148.190 21.920 148.235 ;
        RECT 13.125 147.895 16.790 148.035 ;
        RECT 18.860 148.035 19.180 148.095 ;
        RECT 20.255 148.035 20.545 148.080 ;
        RECT 18.860 147.895 20.545 148.035 ;
        RECT 13.125 147.850 13.415 147.895 ;
        RECT 18.860 147.835 19.180 147.895 ;
        RECT 20.255 147.850 20.545 147.895 ;
        RECT 22.080 147.835 22.400 148.095 ;
        RECT 22.540 148.035 22.860 148.095 ;
        RECT 24.700 148.035 24.840 148.575 ;
        RECT 28.520 148.515 28.840 148.575 ;
        RECT 29.915 148.715 30.205 148.760 ;
        RECT 33.120 148.715 33.440 148.775 ;
        RECT 42.320 148.715 42.640 148.775 ;
        RECT 29.915 148.575 33.440 148.715 ;
        RECT 29.915 148.530 30.205 148.575 ;
        RECT 33.120 148.515 33.440 148.575 ;
        RECT 41.950 148.575 42.640 148.715 ;
        RECT 26.220 148.375 26.540 148.435 ;
        RECT 32.200 148.375 32.520 148.435 ;
        RECT 38.180 148.375 38.500 148.435 ;
        RECT 26.220 148.235 26.910 148.375 ;
        RECT 26.220 148.175 26.540 148.235 ;
        RECT 26.770 148.080 26.910 148.235 ;
        RECT 32.200 148.235 38.500 148.375 ;
        RECT 32.200 148.175 32.520 148.235 ;
        RECT 38.180 148.175 38.500 148.235 ;
        RECT 22.540 147.895 24.840 148.035 ;
        RECT 22.540 147.835 22.860 147.895 ;
        RECT 26.695 147.850 26.985 148.080 ;
        RECT 32.290 148.035 32.430 148.175 ;
        RECT 41.950 148.080 42.090 148.575 ;
        RECT 42.320 148.515 42.640 148.575 ;
        RECT 42.795 148.715 43.085 148.760 ;
        RECT 43.240 148.715 43.560 148.775 ;
        RECT 42.795 148.575 43.560 148.715 ;
        RECT 42.795 148.530 43.085 148.575 ;
        RECT 43.240 148.515 43.560 148.575 ;
        RECT 59.800 148.715 60.120 148.775 ;
        RECT 66.715 148.715 67.005 148.760 ;
        RECT 67.160 148.715 67.480 148.775 ;
        RECT 59.800 148.575 66.010 148.715 ;
        RECT 59.800 148.515 60.120 148.575 ;
        RECT 44.175 148.375 44.465 148.420 ;
        RECT 45.080 148.375 45.400 148.435 ;
        RECT 47.840 148.375 48.160 148.435 ;
        RECT 52.440 148.375 52.760 148.435 ;
        RECT 44.175 148.235 45.400 148.375 ;
        RECT 44.175 148.190 44.465 148.235 ;
        RECT 45.080 148.175 45.400 148.235 ;
        RECT 45.630 148.235 52.760 148.375 ;
        RECT 30.450 147.895 32.430 148.035 ;
        RECT 16.990 147.695 17.280 147.740 ;
        RECT 16.990 147.555 19.525 147.695 ;
        RECT 16.990 147.510 17.280 147.555 ;
        RECT 15.180 147.400 15.500 147.415 ;
        RECT 19.310 147.400 19.525 147.555 ;
        RECT 25.760 147.495 26.080 147.755 ;
        RECT 28.980 147.495 29.300 147.755 ;
        RECT 30.450 147.740 30.590 147.895 ;
        RECT 41.875 147.850 42.165 148.080 ;
        RECT 45.630 148.035 45.770 148.235 ;
        RECT 47.840 148.175 48.160 148.235 ;
        RECT 52.440 148.175 52.760 148.235 ;
        RECT 57.470 148.375 57.760 148.420 ;
        RECT 60.250 148.375 60.540 148.420 ;
        RECT 62.110 148.375 62.400 148.420 ;
        RECT 57.470 148.235 62.400 148.375 ;
        RECT 65.870 148.375 66.010 148.575 ;
        RECT 66.715 148.575 67.480 148.715 ;
        RECT 66.715 148.530 67.005 148.575 ;
        RECT 67.160 148.515 67.480 148.575 ;
        RECT 70.380 148.515 70.700 148.775 ;
        RECT 92.920 148.515 93.240 148.775 ;
        RECT 96.615 148.715 96.905 148.760 ;
        RECT 97.060 148.715 97.380 148.775 ;
        RECT 96.615 148.575 97.380 148.715 ;
        RECT 96.615 148.530 96.905 148.575 ;
        RECT 97.060 148.515 97.380 148.575 ;
        RECT 97.980 148.715 98.300 148.775 ;
        RECT 107.640 148.715 107.960 148.775 ;
        RECT 97.980 148.575 107.960 148.715 ;
        RECT 97.980 148.515 98.300 148.575 ;
        RECT 107.640 148.515 107.960 148.575 ;
        RECT 71.760 148.375 72.080 148.435 ;
        RECT 65.870 148.235 72.080 148.375 ;
        RECT 57.470 148.190 57.760 148.235 ;
        RECT 60.250 148.190 60.540 148.235 ;
        RECT 62.110 148.190 62.400 148.235 ;
        RECT 48.300 148.035 48.620 148.095 ;
        RECT 53.605 148.035 53.895 148.080 ;
        RECT 56.120 148.035 56.440 148.095 ;
        RECT 42.410 147.895 45.770 148.035 ;
        RECT 46.090 147.895 50.830 148.035 ;
        RECT 30.375 147.510 30.665 147.740 ;
        RECT 31.295 147.510 31.585 147.740 ;
        RECT 15.130 147.355 15.500 147.400 ;
        RECT 18.390 147.355 18.680 147.400 ;
        RECT 15.130 147.215 18.680 147.355 ;
        RECT 15.130 147.170 15.500 147.215 ;
        RECT 18.390 147.170 18.680 147.215 ;
        RECT 19.310 147.355 19.600 147.400 ;
        RECT 21.170 147.355 21.460 147.400 ;
        RECT 26.235 147.355 26.525 147.400 ;
        RECT 31.370 147.355 31.510 147.510 ;
        RECT 31.740 147.495 32.060 147.755 ;
        RECT 32.215 147.695 32.505 147.740 ;
        RECT 36.340 147.695 36.660 147.755 ;
        RECT 32.215 147.555 36.660 147.695 ;
        RECT 32.215 147.510 32.505 147.555 ;
        RECT 36.340 147.495 36.660 147.555 ;
        RECT 36.815 147.695 37.105 147.740 ;
        RECT 42.410 147.695 42.550 147.895 ;
        RECT 36.815 147.555 42.550 147.695 ;
        RECT 36.815 147.510 37.105 147.555 ;
        RECT 36.890 147.355 37.030 147.510 ;
        RECT 42.780 147.495 43.100 147.755 ;
        RECT 45.540 147.495 45.860 147.755 ;
        RECT 46.090 147.740 46.230 147.895 ;
        RECT 48.300 147.835 48.620 147.895 ;
        RECT 50.690 147.755 50.830 147.895 ;
        RECT 51.150 147.895 56.440 148.035 ;
        RECT 46.015 147.510 46.305 147.740 ;
        RECT 46.460 147.495 46.780 147.755 ;
        RECT 47.395 147.695 47.685 147.740 ;
        RECT 47.395 147.555 49.910 147.695 ;
        RECT 47.395 147.510 47.685 147.555 ;
        RECT 19.310 147.215 21.460 147.355 ;
        RECT 19.310 147.170 19.600 147.215 ;
        RECT 21.170 147.170 21.460 147.215 ;
        RECT 23.090 147.215 31.510 147.355 ;
        RECT 32.290 147.215 37.030 147.355 ;
        RECT 15.180 147.155 15.500 147.170 ;
        RECT 17.940 147.015 18.260 147.075 ;
        RECT 23.090 147.015 23.230 147.215 ;
        RECT 26.235 147.170 26.525 147.215 ;
        RECT 17.940 146.875 23.230 147.015 ;
        RECT 23.935 147.015 24.225 147.060 ;
        RECT 26.680 147.015 27.000 147.075 ;
        RECT 23.935 146.875 27.000 147.015 ;
        RECT 17.940 146.815 18.260 146.875 ;
        RECT 23.935 146.830 24.225 146.875 ;
        RECT 26.680 146.815 27.000 146.875 ;
        RECT 28.520 147.015 28.840 147.075 ;
        RECT 32.290 147.015 32.430 147.215 ;
        RECT 41.415 147.170 41.705 147.400 ;
        RECT 48.775 147.355 49.065 147.400 ;
        RECT 43.330 147.215 49.065 147.355 ;
        RECT 49.770 147.355 49.910 147.555 ;
        RECT 50.140 147.495 50.460 147.755 ;
        RECT 50.600 147.495 50.920 147.755 ;
        RECT 51.150 147.740 51.290 147.895 ;
        RECT 53.605 147.850 53.895 147.895 ;
        RECT 56.120 147.835 56.440 147.895 ;
        RECT 58.880 148.035 59.200 148.095 ;
        RECT 60.735 148.035 61.025 148.080 ;
        RECT 58.880 147.895 61.025 148.035 ;
        RECT 58.880 147.835 59.200 147.895 ;
        RECT 60.735 147.850 61.025 147.895 ;
        RECT 61.180 148.035 61.500 148.095 ;
        RECT 62.575 148.035 62.865 148.080 ;
        RECT 61.180 147.895 62.865 148.035 ;
        RECT 61.180 147.835 61.500 147.895 ;
        RECT 62.575 147.850 62.865 147.895 ;
        RECT 64.400 148.035 64.720 148.095 ;
        RECT 65.795 148.035 66.085 148.080 ;
        RECT 64.400 147.895 66.085 148.035 ;
        RECT 64.400 147.835 64.720 147.895 ;
        RECT 65.795 147.850 66.085 147.895 ;
        RECT 66.700 147.835 67.020 148.095 ;
        RECT 51.075 147.510 51.365 147.740 ;
        RECT 51.980 147.495 52.300 147.755 ;
        RECT 57.470 147.695 57.760 147.740 ;
        RECT 65.335 147.695 65.625 147.740 ;
        RECT 66.790 147.695 66.930 147.835 ;
        RECT 67.250 147.740 67.390 148.235 ;
        RECT 71.760 148.175 72.080 148.235 ;
        RECT 76.380 148.375 76.670 148.420 ;
        RECT 78.240 148.375 78.530 148.420 ;
        RECT 81.020 148.375 81.310 148.420 ;
        RECT 76.380 148.235 81.310 148.375 ;
        RECT 76.380 148.190 76.670 148.235 ;
        RECT 78.240 148.190 78.530 148.235 ;
        RECT 81.020 148.190 81.310 148.235 ;
        RECT 86.940 148.375 87.260 148.435 ;
        RECT 105.340 148.375 105.660 148.435 ;
        RECT 86.940 148.235 105.660 148.375 ;
        RECT 86.940 148.175 87.260 148.235 ;
        RECT 79.120 148.035 79.440 148.095 ;
        RECT 84.180 148.035 84.500 148.095 ;
        RECT 86.495 148.035 86.785 148.080 ;
        RECT 92.920 148.035 93.240 148.095 ;
        RECT 68.170 147.895 81.650 148.035 ;
        RECT 68.170 147.740 68.310 147.895 ;
        RECT 79.120 147.835 79.440 147.895 ;
        RECT 57.470 147.555 60.005 147.695 ;
        RECT 57.470 147.510 57.760 147.555 ;
        RECT 52.070 147.355 52.210 147.495 ;
        RECT 49.770 147.215 52.210 147.355 ;
        RECT 53.820 147.355 54.140 147.415 ;
        RECT 59.790 147.400 60.005 147.555 ;
        RECT 65.335 147.555 66.930 147.695 ;
        RECT 65.335 147.510 65.625 147.555 ;
        RECT 67.175 147.510 67.465 147.740 ;
        RECT 68.095 147.510 68.385 147.740 ;
        RECT 68.540 147.495 68.860 147.755 ;
        RECT 69.015 147.695 69.305 147.740 ;
        RECT 70.380 147.695 70.700 147.755 ;
        RECT 72.235 147.695 72.525 147.740 ;
        RECT 69.015 147.555 72.525 147.695 ;
        RECT 69.015 147.510 69.305 147.555 ;
        RECT 70.380 147.495 70.700 147.555 ;
        RECT 72.235 147.510 72.525 147.555 ;
        RECT 72.680 147.495 73.000 147.755 ;
        RECT 73.140 147.495 73.460 147.755 ;
        RECT 74.075 147.510 74.365 147.740 ;
        RECT 74.535 147.695 74.825 147.740 ;
        RECT 74.980 147.695 75.300 147.755 ;
        RECT 74.535 147.555 75.300 147.695 ;
        RECT 74.535 147.510 74.825 147.555 ;
        RECT 55.610 147.355 55.900 147.400 ;
        RECT 58.870 147.355 59.160 147.400 ;
        RECT 53.820 147.215 59.160 147.355 ;
        RECT 28.520 146.875 32.430 147.015 ;
        RECT 32.660 147.015 32.980 147.075 ;
        RECT 33.595 147.015 33.885 147.060 ;
        RECT 32.660 146.875 33.885 147.015 ;
        RECT 28.520 146.815 28.840 146.875 ;
        RECT 32.660 146.815 32.980 146.875 ;
        RECT 33.595 146.830 33.885 146.875 ;
        RECT 37.275 147.015 37.565 147.060 ;
        RECT 37.720 147.015 38.040 147.075 ;
        RECT 37.275 146.875 38.040 147.015 ;
        RECT 41.490 147.015 41.630 147.170 ;
        RECT 43.330 147.015 43.470 147.215 ;
        RECT 48.775 147.170 49.065 147.215 ;
        RECT 53.820 147.155 54.140 147.215 ;
        RECT 55.610 147.170 55.900 147.215 ;
        RECT 58.870 147.170 59.160 147.215 ;
        RECT 59.790 147.355 60.080 147.400 ;
        RECT 61.650 147.355 61.940 147.400 ;
        RECT 59.790 147.215 61.940 147.355 ;
        RECT 59.790 147.170 60.080 147.215 ;
        RECT 61.650 147.170 61.940 147.215 ;
        RECT 66.715 147.355 67.005 147.400 ;
        RECT 70.855 147.355 71.145 147.400 ;
        RECT 66.715 147.215 71.145 147.355 ;
        RECT 66.715 147.170 67.005 147.215 ;
        RECT 70.855 147.170 71.145 147.215 ;
        RECT 71.760 147.355 72.080 147.415 ;
        RECT 74.150 147.355 74.290 147.510 ;
        RECT 74.980 147.495 75.300 147.555 ;
        RECT 75.900 147.495 76.220 147.755 ;
        RECT 77.755 147.695 78.045 147.740 ;
        RECT 81.020 147.695 81.310 147.740 ;
        RECT 76.450 147.555 78.045 147.695 ;
        RECT 76.450 147.355 76.590 147.555 ;
        RECT 77.755 147.510 78.045 147.555 ;
        RECT 78.775 147.555 81.310 147.695 ;
        RECT 81.510 147.695 81.650 147.895 ;
        RECT 84.180 147.895 93.240 148.035 ;
        RECT 84.180 147.835 84.500 147.895 ;
        RECT 86.495 147.850 86.785 147.895 ;
        RECT 92.920 147.835 93.240 147.895 ;
        RECT 96.155 148.035 96.445 148.080 ;
        RECT 96.600 148.035 96.920 148.095 ;
        RECT 96.155 147.895 96.920 148.035 ;
        RECT 96.155 147.850 96.445 147.895 ;
        RECT 96.600 147.835 96.920 147.895 ;
        RECT 87.415 147.695 87.705 147.740 ;
        RECT 92.015 147.695 92.305 147.740 ;
        RECT 81.510 147.555 87.705 147.695 ;
        RECT 78.775 147.400 78.990 147.555 ;
        RECT 81.020 147.510 81.310 147.555 ;
        RECT 87.415 147.510 87.705 147.555 ;
        RECT 89.330 147.555 92.305 147.695 ;
        RECT 71.760 147.215 74.290 147.355 ;
        RECT 75.530 147.215 76.590 147.355 ;
        RECT 76.840 147.355 77.130 147.400 ;
        RECT 78.700 147.355 78.990 147.400 ;
        RECT 76.840 147.215 78.990 147.355 ;
        RECT 71.760 147.155 72.080 147.215 ;
        RECT 41.490 146.875 43.470 147.015 ;
        RECT 43.715 147.015 44.005 147.060 ;
        RECT 57.040 147.015 57.360 147.075 ;
        RECT 43.715 146.875 57.360 147.015 ;
        RECT 37.275 146.830 37.565 146.875 ;
        RECT 37.720 146.815 38.040 146.875 ;
        RECT 43.715 146.830 44.005 146.875 ;
        RECT 57.040 146.815 57.360 146.875 ;
        RECT 63.940 147.015 64.260 147.075 ;
        RECT 64.415 147.015 64.705 147.060 ;
        RECT 63.940 146.875 64.705 147.015 ;
        RECT 63.940 146.815 64.260 146.875 ;
        RECT 64.415 146.830 64.705 146.875 ;
        RECT 68.540 147.015 68.860 147.075 ;
        RECT 72.680 147.015 73.000 147.075 ;
        RECT 75.530 147.060 75.670 147.215 ;
        RECT 76.840 147.170 77.130 147.215 ;
        RECT 78.700 147.170 78.990 147.215 ;
        RECT 79.620 147.355 79.910 147.400 ;
        RECT 82.340 147.355 82.660 147.415 ;
        RECT 82.880 147.355 83.170 147.400 ;
        RECT 79.620 147.215 83.170 147.355 ;
        RECT 79.620 147.170 79.910 147.215 ;
        RECT 82.340 147.155 82.660 147.215 ;
        RECT 82.880 147.170 83.170 147.215 ;
        RECT 68.540 146.875 73.000 147.015 ;
        RECT 68.540 146.815 68.860 146.875 ;
        RECT 72.680 146.815 73.000 146.875 ;
        RECT 75.455 146.830 75.745 147.060 ;
        RECT 80.040 147.015 80.360 147.075 ;
        RECT 84.885 147.015 85.175 147.060 ;
        RECT 80.040 146.875 85.175 147.015 ;
        RECT 80.040 146.815 80.360 146.875 ;
        RECT 84.885 146.830 85.175 146.875 ;
        RECT 86.940 146.815 87.260 147.075 ;
        RECT 89.330 147.060 89.470 147.555 ;
        RECT 92.015 147.510 92.305 147.555 ;
        RECT 94.300 147.695 94.620 147.755 ;
        RECT 95.235 147.695 95.525 147.740 ;
        RECT 94.300 147.555 95.525 147.695 ;
        RECT 94.300 147.495 94.620 147.555 ;
        RECT 95.235 147.510 95.525 147.555 ;
        RECT 97.980 147.695 98.300 147.755 ;
        RECT 99.450 147.740 99.590 148.235 ;
        RECT 105.340 148.175 105.660 148.235 ;
        RECT 108.990 148.375 109.280 148.420 ;
        RECT 111.770 148.375 112.060 148.420 ;
        RECT 113.630 148.375 113.920 148.420 ;
        RECT 108.990 148.235 113.920 148.375 ;
        RECT 108.990 148.190 109.280 148.235 ;
        RECT 111.770 148.190 112.060 148.235 ;
        RECT 113.630 148.190 113.920 148.235 ;
        RECT 101.675 148.035 101.965 148.080 ;
        RECT 104.880 148.035 105.200 148.095 ;
        RECT 112.700 148.035 113.020 148.095 ;
        RECT 101.675 147.895 105.200 148.035 ;
        RECT 101.675 147.850 101.965 147.895 ;
        RECT 104.880 147.835 105.200 147.895 ;
        RECT 107.500 147.895 113.020 148.035 ;
        RECT 98.455 147.695 98.745 147.740 ;
        RECT 97.980 147.555 98.745 147.695 ;
        RECT 97.980 147.495 98.300 147.555 ;
        RECT 98.455 147.510 98.745 147.555 ;
        RECT 98.915 147.510 99.205 147.740 ;
        RECT 99.375 147.510 99.665 147.740 ;
        RECT 99.820 147.680 100.140 147.755 ;
        RECT 100.295 147.680 100.585 147.740 ;
        RECT 107.500 147.695 107.640 147.895 ;
        RECT 112.700 147.835 113.020 147.895 ;
        RECT 99.820 147.540 100.585 147.680 ;
        RECT 96.615 147.355 96.905 147.400 ;
        RECT 97.075 147.355 97.365 147.400 ;
        RECT 96.615 147.215 97.365 147.355 ;
        RECT 98.990 147.355 99.130 147.510 ;
        RECT 99.820 147.495 100.140 147.540 ;
        RECT 100.295 147.510 100.585 147.540 ;
        RECT 101.750 147.555 107.640 147.695 ;
        RECT 108.990 147.695 109.280 147.740 ;
        RECT 108.990 147.555 111.525 147.695 ;
        RECT 100.740 147.355 101.060 147.415 ;
        RECT 98.990 147.215 101.060 147.355 ;
        RECT 96.615 147.170 96.905 147.215 ;
        RECT 97.075 147.170 97.365 147.215 ;
        RECT 100.740 147.155 101.060 147.215 ;
        RECT 89.255 146.830 89.545 147.060 ;
        RECT 94.315 147.015 94.605 147.060 ;
        RECT 101.750 147.015 101.890 147.555 ;
        RECT 108.990 147.510 109.280 147.555 ;
        RECT 102.135 147.170 102.425 147.400 ;
        RECT 94.315 146.875 101.890 147.015 ;
        RECT 102.210 147.015 102.350 147.170 ;
        RECT 102.580 147.155 102.900 147.415 ;
        RECT 105.125 147.355 105.415 147.400 ;
        RECT 106.260 147.355 106.580 147.415 ;
        RECT 104.050 147.215 106.580 147.355 ;
        RECT 104.050 147.015 104.190 147.215 ;
        RECT 105.125 147.170 105.415 147.215 ;
        RECT 106.260 147.155 106.580 147.215 ;
        RECT 107.130 147.355 107.420 147.400 ;
        RECT 108.560 147.355 108.880 147.415 ;
        RECT 111.310 147.400 111.525 147.555 ;
        RECT 112.240 147.495 112.560 147.755 ;
        RECT 114.080 147.495 114.400 147.755 ;
        RECT 110.390 147.355 110.680 147.400 ;
        RECT 107.130 147.215 110.680 147.355 ;
        RECT 107.130 147.170 107.420 147.215 ;
        RECT 108.560 147.155 108.880 147.215 ;
        RECT 110.390 147.170 110.680 147.215 ;
        RECT 111.310 147.355 111.600 147.400 ;
        RECT 113.170 147.355 113.460 147.400 ;
        RECT 111.310 147.215 113.460 147.355 ;
        RECT 111.310 147.170 111.600 147.215 ;
        RECT 113.170 147.170 113.460 147.215 ;
        RECT 102.210 146.875 104.190 147.015 ;
        RECT 104.435 147.015 104.725 147.060 ;
        RECT 109.940 147.015 110.260 147.075 ;
        RECT 104.435 146.875 110.260 147.015 ;
        RECT 94.315 146.830 94.605 146.875 ;
        RECT 104.435 146.830 104.725 146.875 ;
        RECT 109.940 146.815 110.260 146.875 ;
        RECT 10.510 146.195 115.850 146.675 ;
        RECT 14.735 145.995 15.025 146.040 ;
        RECT 15.180 145.995 15.500 146.055 ;
        RECT 14.735 145.855 15.500 145.995 ;
        RECT 14.735 145.810 15.025 145.855 ;
        RECT 15.180 145.795 15.500 145.855 ;
        RECT 23.000 145.995 23.320 146.055 ;
        RECT 46.015 145.995 46.305 146.040 ;
        RECT 46.460 145.995 46.780 146.055 ;
        RECT 23.000 145.855 32.430 145.995 ;
        RECT 23.000 145.795 23.320 145.855 ;
        RECT 17.890 145.655 18.180 145.700 ;
        RECT 19.320 145.655 19.640 145.715 ;
        RECT 21.150 145.655 21.440 145.700 ;
        RECT 17.890 145.515 21.440 145.655 ;
        RECT 17.890 145.470 18.180 145.515 ;
        RECT 19.320 145.455 19.640 145.515 ;
        RECT 21.150 145.470 21.440 145.515 ;
        RECT 22.070 145.655 22.360 145.700 ;
        RECT 23.930 145.655 24.220 145.700 ;
        RECT 22.070 145.515 24.220 145.655 ;
        RECT 22.070 145.470 22.360 145.515 ;
        RECT 23.930 145.470 24.220 145.515 ;
        RECT 14.720 145.315 15.040 145.375 ;
        RECT 15.195 145.315 15.485 145.360 ;
        RECT 14.720 145.175 15.485 145.315 ;
        RECT 14.720 145.115 15.040 145.175 ;
        RECT 15.195 145.130 15.485 145.175 ;
        RECT 19.750 145.315 20.040 145.360 ;
        RECT 22.070 145.315 22.285 145.470 ;
        RECT 19.750 145.175 22.285 145.315 ;
        RECT 23.015 145.315 23.305 145.360 ;
        RECT 25.760 145.315 26.080 145.375 ;
        RECT 23.015 145.175 26.080 145.315 ;
        RECT 19.750 145.130 20.040 145.175 ;
        RECT 23.015 145.130 23.305 145.175 ;
        RECT 25.760 145.115 26.080 145.175 ;
        RECT 26.680 145.115 27.000 145.375 ;
        RECT 30.820 145.360 31.140 145.375 ;
        RECT 30.820 145.130 31.355 145.360 ;
        RECT 31.740 145.315 32.060 145.375 ;
        RECT 32.290 145.360 32.430 145.855 ;
        RECT 46.015 145.855 46.780 145.995 ;
        RECT 46.015 145.810 46.305 145.855 ;
        RECT 46.460 145.795 46.780 145.855 ;
        RECT 53.820 145.795 54.140 146.055 ;
        RECT 56.120 145.795 56.440 146.055 ;
        RECT 57.960 145.995 58.280 146.055 ;
        RECT 58.435 145.995 58.725 146.040 ;
        RECT 57.960 145.855 58.725 145.995 ;
        RECT 57.960 145.795 58.280 145.855 ;
        RECT 58.435 145.810 58.725 145.855 ;
        RECT 73.140 145.995 73.460 146.055 ;
        RECT 74.075 145.995 74.365 146.040 ;
        RECT 73.140 145.855 74.365 145.995 ;
        RECT 73.140 145.795 73.460 145.855 ;
        RECT 74.075 145.810 74.365 145.855 ;
        RECT 74.980 145.995 75.300 146.055 ;
        RECT 76.375 145.995 76.665 146.040 ;
        RECT 74.980 145.855 76.665 145.995 ;
        RECT 37.720 145.700 38.040 145.715 ;
        RECT 34.980 145.655 35.270 145.700 ;
        RECT 36.840 145.655 37.130 145.700 ;
        RECT 34.980 145.515 37.130 145.655 ;
        RECT 34.980 145.470 35.270 145.515 ;
        RECT 36.840 145.470 37.130 145.515 ;
        RECT 31.545 145.175 32.060 145.315 ;
        RECT 30.820 145.115 31.140 145.130 ;
        RECT 31.740 145.115 32.060 145.175 ;
        RECT 32.215 145.130 32.505 145.360 ;
        RECT 33.135 145.315 33.425 145.360 ;
        RECT 36.915 145.315 37.130 145.470 ;
        RECT 37.720 145.655 38.050 145.700 ;
        RECT 41.020 145.655 41.310 145.700 ;
        RECT 37.720 145.515 41.310 145.655 ;
        RECT 37.720 145.470 38.050 145.515 ;
        RECT 41.020 145.470 41.310 145.515 ;
        RECT 48.760 145.655 49.080 145.715 ;
        RECT 50.140 145.655 50.460 145.715 ;
        RECT 70.380 145.655 70.700 145.715 ;
        RECT 48.760 145.515 70.700 145.655 ;
        RECT 74.150 145.655 74.290 145.810 ;
        RECT 74.980 145.795 75.300 145.855 ;
        RECT 76.375 145.810 76.665 145.855 ;
        RECT 79.120 145.795 79.440 146.055 ;
        RECT 79.595 145.995 79.885 146.040 ;
        RECT 80.040 145.995 80.360 146.055 ;
        RECT 79.595 145.855 80.360 145.995 ;
        RECT 79.595 145.810 79.885 145.855 ;
        RECT 79.670 145.655 79.810 145.810 ;
        RECT 80.040 145.795 80.360 145.855 ;
        RECT 82.340 145.795 82.660 146.055 ;
        RECT 86.940 145.795 87.260 146.055 ;
        RECT 108.100 145.995 108.420 146.055 ;
        RECT 98.070 145.855 108.420 145.995 ;
        RECT 74.150 145.515 79.810 145.655 ;
        RECT 37.720 145.455 38.040 145.470 ;
        RECT 48.760 145.455 49.080 145.515 ;
        RECT 50.140 145.455 50.460 145.515 ;
        RECT 70.380 145.455 70.700 145.515 ;
        RECT 39.160 145.315 39.450 145.360 ;
        RECT 33.135 145.175 36.570 145.315 ;
        RECT 36.915 145.175 39.450 145.315 ;
        RECT 33.135 145.130 33.425 145.175 ;
        RECT 15.885 144.975 16.175 145.020 ;
        RECT 17.940 144.975 18.260 145.035 ;
        RECT 15.885 144.835 18.260 144.975 ;
        RECT 15.885 144.790 16.175 144.835 ;
        RECT 17.940 144.775 18.260 144.835 ;
        RECT 23.920 144.975 24.240 145.035 ;
        RECT 24.855 144.975 25.145 145.020 ;
        RECT 23.920 144.835 31.510 144.975 ;
        RECT 23.920 144.775 24.240 144.835 ;
        RECT 24.855 144.790 25.145 144.835 ;
        RECT 19.750 144.635 20.040 144.680 ;
        RECT 22.530 144.635 22.820 144.680 ;
        RECT 24.390 144.635 24.680 144.680 ;
        RECT 19.750 144.495 24.680 144.635 ;
        RECT 19.750 144.450 20.040 144.495 ;
        RECT 22.530 144.450 22.820 144.495 ;
        RECT 24.390 144.450 24.680 144.495 ;
        RECT 25.760 144.435 26.080 144.695 ;
        RECT 29.915 144.295 30.205 144.340 ;
        RECT 30.820 144.295 31.140 144.355 ;
        RECT 29.915 144.155 31.140 144.295 ;
        RECT 31.370 144.295 31.510 144.835 ;
        RECT 34.055 144.790 34.345 145.020 ;
        RECT 34.130 144.295 34.270 144.790 ;
        RECT 35.880 144.775 36.200 145.035 ;
        RECT 36.430 144.975 36.570 145.175 ;
        RECT 39.160 145.130 39.450 145.175 ;
        RECT 49.220 145.115 49.540 145.375 ;
        RECT 52.440 145.315 52.760 145.375 ;
        RECT 53.375 145.315 53.665 145.360 ;
        RECT 52.440 145.175 53.665 145.315 ;
        RECT 52.440 145.115 52.760 145.175 ;
        RECT 53.375 145.130 53.665 145.175 ;
        RECT 56.580 145.115 56.900 145.375 ;
        RECT 62.100 145.315 62.420 145.375 ;
        RECT 65.795 145.315 66.085 145.360 ;
        RECT 62.100 145.175 66.085 145.315 ;
        RECT 62.100 145.115 62.420 145.175 ;
        RECT 65.795 145.130 66.085 145.175 ;
        RECT 74.060 145.315 74.380 145.375 ;
        RECT 74.535 145.315 74.825 145.360 ;
        RECT 74.060 145.175 74.825 145.315 ;
        RECT 74.060 145.115 74.380 145.175 ;
        RECT 74.535 145.130 74.825 145.175 ;
        RECT 82.815 145.315 83.105 145.360 ;
        RECT 83.260 145.315 83.580 145.375 ;
        RECT 82.815 145.175 83.580 145.315 ;
        RECT 82.815 145.130 83.105 145.175 ;
        RECT 83.260 145.115 83.580 145.175 ;
        RECT 84.195 145.315 84.485 145.360 ;
        RECT 86.480 145.315 86.800 145.375 ;
        RECT 84.195 145.175 86.800 145.315 ;
        RECT 84.195 145.130 84.485 145.175 ;
        RECT 86.480 145.115 86.800 145.175 ;
        RECT 97.075 145.315 97.365 145.360 ;
        RECT 97.520 145.315 97.840 145.375 ;
        RECT 97.075 145.175 97.840 145.315 ;
        RECT 97.075 145.130 97.365 145.175 ;
        RECT 97.520 145.115 97.840 145.175 ;
        RECT 38.180 144.975 38.500 145.035 ;
        RECT 43.025 144.975 43.315 145.020 ;
        RECT 46.000 144.975 46.320 145.035 ;
        RECT 46.475 144.975 46.765 145.020 ;
        RECT 36.430 144.835 39.790 144.975 ;
        RECT 38.180 144.775 38.500 144.835 ;
        RECT 34.520 144.635 34.810 144.680 ;
        RECT 36.380 144.635 36.670 144.680 ;
        RECT 39.160 144.635 39.450 144.680 ;
        RECT 34.520 144.495 39.450 144.635 ;
        RECT 39.650 144.635 39.790 144.835 ;
        RECT 43.025 144.835 46.765 144.975 ;
        RECT 43.025 144.790 43.315 144.835 ;
        RECT 46.000 144.775 46.320 144.835 ;
        RECT 46.475 144.790 46.765 144.835 ;
        RECT 47.395 144.975 47.685 145.020 ;
        RECT 47.840 144.975 48.160 145.035 ;
        RECT 49.310 144.975 49.450 145.115 ;
        RECT 55.215 144.975 55.505 145.020 ;
        RECT 47.395 144.835 55.505 144.975 ;
        RECT 47.395 144.790 47.685 144.835 ;
        RECT 47.840 144.775 48.160 144.835 ;
        RECT 55.215 144.790 55.505 144.835 ;
        RECT 73.600 144.975 73.920 145.035 ;
        RECT 78.675 144.975 78.965 145.020 ;
        RECT 83.720 144.975 84.040 145.035 ;
        RECT 98.070 145.020 98.210 145.855 ;
        RECT 108.100 145.795 108.420 145.855 ;
        RECT 108.560 145.795 108.880 146.055 ;
        RECT 110.875 145.995 111.165 146.040 ;
        RECT 112.240 145.995 112.560 146.055 ;
        RECT 110.875 145.855 112.560 145.995 ;
        RECT 110.875 145.810 111.165 145.855 ;
        RECT 112.240 145.795 112.560 145.855 ;
        RECT 98.455 145.655 98.745 145.700 ;
        RECT 98.915 145.655 99.205 145.700 ;
        RECT 106.260 145.655 106.580 145.715 ;
        RECT 98.455 145.515 99.205 145.655 ;
        RECT 98.455 145.470 98.745 145.515 ;
        RECT 98.915 145.470 99.205 145.515 ;
        RECT 101.290 145.515 106.580 145.655 ;
        RECT 100.280 145.115 100.600 145.375 ;
        RECT 100.740 145.115 101.060 145.375 ;
        RECT 101.290 145.360 101.430 145.515 ;
        RECT 106.260 145.455 106.580 145.515 ;
        RECT 101.215 145.130 101.505 145.360 ;
        RECT 102.120 145.115 102.440 145.375 ;
        RECT 103.040 145.315 103.360 145.375 ;
        RECT 107.180 145.315 107.500 145.375 ;
        RECT 108.115 145.315 108.405 145.360 ;
        RECT 103.040 145.175 108.405 145.315 ;
        RECT 103.040 145.115 103.360 145.175 ;
        RECT 107.180 145.115 107.500 145.175 ;
        RECT 108.115 145.130 108.405 145.175 ;
        RECT 109.940 145.115 110.260 145.375 ;
        RECT 73.600 144.835 84.040 144.975 ;
        RECT 73.600 144.775 73.920 144.835 ;
        RECT 78.675 144.790 78.965 144.835 ;
        RECT 83.720 144.775 84.040 144.835 ;
        RECT 97.995 144.790 98.285 145.020 ;
        RECT 98.900 144.975 99.220 145.035 ;
        RECT 99.820 144.975 100.140 145.035 ;
        RECT 102.210 144.975 102.350 145.115 ;
        RECT 98.900 144.835 102.350 144.975 ;
        RECT 98.900 144.775 99.220 144.835 ;
        RECT 99.820 144.775 100.140 144.835 ;
        RECT 81.435 144.635 81.725 144.680 ;
        RECT 82.800 144.635 83.120 144.695 ;
        RECT 39.650 144.495 44.850 144.635 ;
        RECT 34.520 144.450 34.810 144.495 ;
        RECT 36.380 144.450 36.670 144.495 ;
        RECT 39.160 144.450 39.450 144.495 ;
        RECT 31.370 144.155 34.270 144.295 ;
        RECT 42.780 144.295 43.100 144.355 ;
        RECT 44.175 144.295 44.465 144.340 ;
        RECT 42.780 144.155 44.465 144.295 ;
        RECT 44.710 144.295 44.850 144.495 ;
        RECT 81.435 144.495 83.120 144.635 ;
        RECT 81.435 144.450 81.725 144.495 ;
        RECT 82.800 144.435 83.120 144.495 ;
        RECT 96.155 144.635 96.445 144.680 ;
        RECT 102.580 144.635 102.900 144.695 ;
        RECT 96.155 144.495 102.900 144.635 ;
        RECT 96.155 144.450 96.445 144.495 ;
        RECT 102.580 144.435 102.900 144.495 ;
        RECT 54.740 144.295 55.060 144.355 ;
        RECT 44.710 144.155 55.060 144.295 ;
        RECT 29.915 144.110 30.205 144.155 ;
        RECT 30.820 144.095 31.140 144.155 ;
        RECT 42.780 144.095 43.100 144.155 ;
        RECT 44.175 144.110 44.465 144.155 ;
        RECT 54.740 144.095 55.060 144.155 ;
        RECT 66.715 144.295 67.005 144.340 ;
        RECT 69.000 144.295 69.320 144.355 ;
        RECT 66.715 144.155 69.320 144.295 ;
        RECT 66.715 144.110 67.005 144.155 ;
        RECT 69.000 144.095 69.320 144.155 ;
        RECT 98.440 144.095 98.760 144.355 ;
        RECT 10.510 143.475 115.850 143.955 ;
        RECT 18.860 143.275 19.180 143.335 ;
        RECT 20.255 143.275 20.545 143.320 ;
        RECT 18.860 143.135 20.545 143.275 ;
        RECT 18.860 143.075 19.180 143.135 ;
        RECT 20.255 143.090 20.545 143.135 ;
        RECT 35.880 143.275 36.200 143.335 ;
        RECT 41.875 143.275 42.165 143.320 ;
        RECT 35.880 143.135 42.165 143.275 ;
        RECT 35.880 143.075 36.200 143.135 ;
        RECT 41.875 143.090 42.165 143.135 ;
        RECT 68.540 143.075 68.860 143.335 ;
        RECT 19.320 142.935 19.640 142.995 ;
        RECT 21.175 142.935 21.465 142.980 ;
        RECT 19.320 142.795 21.465 142.935 ;
        RECT 19.320 142.735 19.640 142.795 ;
        RECT 21.175 142.750 21.465 142.795 ;
        RECT 57.615 142.935 57.905 142.980 ;
        RECT 60.735 142.935 61.025 142.980 ;
        RECT 62.625 142.935 62.915 142.980 ;
        RECT 57.615 142.795 62.915 142.935 ;
        RECT 57.615 142.750 57.905 142.795 ;
        RECT 60.735 142.750 61.025 142.795 ;
        RECT 62.625 142.750 62.915 142.795 ;
        RECT 71.760 142.735 72.080 142.995 ;
        RECT 77.710 142.935 78.000 142.980 ;
        RECT 80.490 142.935 80.780 142.980 ;
        RECT 82.350 142.935 82.640 142.980 ;
        RECT 77.710 142.795 82.640 142.935 ;
        RECT 77.710 142.750 78.000 142.795 ;
        RECT 80.490 142.750 80.780 142.795 ;
        RECT 82.350 142.750 82.640 142.795 ;
        RECT 69.015 142.595 69.305 142.640 ;
        RECT 69.460 142.595 69.780 142.655 ;
        RECT 46.550 142.455 51.750 142.595 ;
        RECT 46.550 142.315 46.690 142.455 ;
        RECT 18.400 142.255 18.720 142.315 ;
        RECT 19.335 142.255 19.625 142.300 ;
        RECT 18.400 142.115 19.625 142.255 ;
        RECT 18.400 142.055 18.720 142.115 ;
        RECT 19.335 142.070 19.625 142.115 ;
        RECT 21.635 142.255 21.925 142.300 ;
        RECT 22.540 142.255 22.860 142.315 ;
        RECT 21.635 142.115 22.860 142.255 ;
        RECT 21.635 142.070 21.925 142.115 ;
        RECT 22.540 142.055 22.860 142.115 ;
        RECT 42.780 142.055 43.100 142.315 ;
        RECT 44.535 142.255 44.825 142.300 ;
        RECT 44.535 142.070 44.850 142.255 ;
        RECT 44.710 141.915 44.850 142.070 ;
        RECT 45.080 142.055 45.400 142.315 ;
        RECT 45.555 142.255 45.845 142.300 ;
        RECT 46.000 142.255 46.320 142.315 ;
        RECT 45.555 142.115 46.320 142.255 ;
        RECT 45.555 142.070 45.845 142.115 ;
        RECT 46.000 142.055 46.320 142.115 ;
        RECT 46.460 142.055 46.780 142.315 ;
        RECT 48.760 142.255 49.080 142.315 ;
        RECT 51.610 142.300 51.750 142.455 ;
        RECT 69.015 142.455 69.780 142.595 ;
        RECT 71.850 142.595 71.990 142.735 ;
        RECT 75.900 142.595 76.220 142.655 ;
        RECT 78.660 142.595 78.980 142.655 ;
        RECT 71.850 142.455 73.370 142.595 ;
        RECT 69.015 142.410 69.305 142.455 ;
        RECT 69.460 142.395 69.780 142.455 ;
        RECT 49.695 142.255 49.985 142.300 ;
        RECT 48.760 142.115 49.985 142.255 ;
        RECT 48.760 142.055 49.080 142.115 ;
        RECT 49.695 142.070 49.985 142.115 ;
        RECT 50.155 142.070 50.445 142.300 ;
        RECT 50.615 142.070 50.905 142.300 ;
        RECT 51.535 142.255 51.825 142.300 ;
        RECT 51.980 142.255 52.300 142.315 ;
        RECT 51.535 142.115 52.300 142.255 ;
        RECT 51.535 142.070 51.825 142.115 ;
        RECT 48.850 141.915 48.990 142.055 ;
        RECT 44.710 141.775 48.990 141.915 ;
        RECT 49.220 141.915 49.540 141.975 ;
        RECT 50.230 141.915 50.370 142.070 ;
        RECT 49.220 141.775 50.370 141.915 ;
        RECT 49.220 141.715 49.540 141.775 ;
        RECT 37.720 141.575 38.040 141.635 ;
        RECT 43.255 141.575 43.545 141.620 ;
        RECT 37.720 141.435 43.545 141.575 ;
        RECT 37.720 141.375 38.040 141.435 ;
        RECT 43.255 141.390 43.545 141.435 ;
        RECT 44.160 141.575 44.480 141.635 ;
        RECT 48.315 141.575 48.605 141.620 ;
        RECT 44.160 141.435 48.605 141.575 ;
        RECT 50.690 141.575 50.830 142.070 ;
        RECT 51.980 142.055 52.300 142.115 ;
        RECT 52.440 142.255 52.760 142.315 ;
        RECT 53.375 142.255 53.665 142.300 ;
        RECT 52.440 142.115 53.665 142.255 ;
        RECT 52.440 142.055 52.760 142.115 ;
        RECT 53.375 142.070 53.665 142.115 ;
        RECT 56.535 141.960 56.825 142.275 ;
        RECT 57.615 142.255 57.905 142.300 ;
        RECT 61.195 142.255 61.485 142.300 ;
        RECT 63.030 142.255 63.320 142.300 ;
        RECT 57.615 142.115 63.320 142.255 ;
        RECT 57.615 142.070 57.905 142.115 ;
        RECT 61.195 142.070 61.485 142.115 ;
        RECT 63.030 142.070 63.320 142.115 ;
        RECT 63.480 142.055 63.800 142.315 ;
        RECT 68.080 142.055 68.400 142.315 ;
        RECT 70.380 142.255 70.700 142.315 ;
        RECT 73.230 142.300 73.370 142.455 ;
        RECT 75.900 142.455 80.730 142.595 ;
        RECT 75.900 142.395 76.220 142.455 ;
        RECT 78.660 142.395 78.980 142.455 ;
        RECT 71.315 142.255 71.605 142.300 ;
        RECT 70.380 142.115 71.605 142.255 ;
        RECT 70.380 142.055 70.700 142.115 ;
        RECT 71.315 142.070 71.605 142.115 ;
        RECT 71.775 142.070 72.065 142.300 ;
        RECT 72.235 142.070 72.525 142.300 ;
        RECT 73.155 142.070 73.445 142.300 ;
        RECT 77.710 142.255 78.000 142.300 ;
        RECT 80.590 142.255 80.730 142.455 ;
        RECT 80.960 142.395 81.280 142.655 ;
        RECT 105.340 142.395 105.660 142.655 ;
        RECT 82.815 142.255 83.105 142.300 ;
        RECT 77.710 142.115 80.245 142.255 ;
        RECT 80.590 142.115 83.105 142.255 ;
        RECT 77.710 142.070 78.000 142.115 ;
        RECT 53.835 141.915 54.125 141.960 ;
        RECT 56.235 141.915 56.825 141.960 ;
        RECT 59.475 141.915 60.125 141.960 ;
        RECT 53.835 141.775 60.125 141.915 ;
        RECT 53.835 141.730 54.125 141.775 ;
        RECT 56.235 141.730 56.525 141.775 ;
        RECT 59.475 141.730 60.125 141.775 ;
        RECT 62.115 141.915 62.405 141.960 ;
        RECT 62.560 141.915 62.880 141.975 ;
        RECT 62.115 141.775 62.880 141.915 ;
        RECT 62.115 141.730 62.405 141.775 ;
        RECT 62.560 141.715 62.880 141.775 ;
        RECT 69.475 141.915 69.765 141.960 ;
        RECT 69.935 141.915 70.225 141.960 ;
        RECT 69.475 141.775 70.225 141.915 ;
        RECT 69.475 141.730 69.765 141.775 ;
        RECT 69.935 141.730 70.225 141.775 ;
        RECT 70.840 141.915 71.160 141.975 ;
        RECT 71.850 141.915 71.990 142.070 ;
        RECT 70.840 141.775 71.990 141.915 ;
        RECT 72.310 141.915 72.450 142.070 ;
        RECT 74.060 141.960 74.380 141.975 ;
        RECT 79.120 141.960 79.440 141.975 ;
        RECT 73.845 141.915 74.380 141.960 ;
        RECT 72.310 141.775 74.380 141.915 ;
        RECT 70.840 141.715 71.160 141.775 ;
        RECT 54.740 141.575 55.060 141.635 ;
        RECT 50.690 141.435 55.060 141.575 ;
        RECT 44.160 141.375 44.480 141.435 ;
        RECT 48.315 141.390 48.605 141.435 ;
        RECT 54.740 141.375 55.060 141.435 ;
        RECT 67.175 141.575 67.465 141.620 ;
        RECT 68.080 141.575 68.400 141.635 ;
        RECT 67.175 141.435 68.400 141.575 ;
        RECT 71.850 141.575 71.990 141.775 ;
        RECT 73.845 141.730 74.380 141.775 ;
        RECT 75.850 141.915 76.140 141.960 ;
        RECT 79.110 141.915 79.440 141.960 ;
        RECT 75.850 141.775 79.440 141.915 ;
        RECT 75.850 141.730 76.140 141.775 ;
        RECT 79.110 141.730 79.440 141.775 ;
        RECT 80.030 141.960 80.245 142.115 ;
        RECT 82.815 142.070 83.105 142.115 ;
        RECT 106.260 142.255 106.580 142.315 ;
        RECT 106.735 142.255 107.025 142.300 ;
        RECT 106.260 142.115 107.025 142.255 ;
        RECT 106.260 142.055 106.580 142.115 ;
        RECT 106.735 142.070 107.025 142.115 ;
        RECT 107.180 142.255 107.500 142.315 ;
        RECT 109.035 142.255 109.325 142.300 ;
        RECT 107.180 142.115 109.325 142.255 ;
        RECT 107.180 142.055 107.500 142.115 ;
        RECT 109.035 142.070 109.325 142.115 ;
        RECT 80.030 141.915 80.320 141.960 ;
        RECT 81.890 141.915 82.180 141.960 ;
        RECT 80.030 141.775 82.180 141.915 ;
        RECT 80.030 141.730 80.320 141.775 ;
        RECT 81.890 141.730 82.180 141.775 ;
        RECT 74.060 141.715 74.380 141.730 ;
        RECT 79.120 141.715 79.440 141.730 ;
        RECT 72.680 141.575 73.000 141.635 ;
        RECT 71.850 141.435 73.000 141.575 ;
        RECT 67.175 141.390 67.465 141.435 ;
        RECT 68.080 141.375 68.400 141.435 ;
        RECT 72.680 141.375 73.000 141.435 ;
        RECT 104.880 141.575 105.200 141.635 ;
        RECT 106.275 141.575 106.565 141.620 ;
        RECT 104.880 141.435 106.565 141.575 ;
        RECT 104.880 141.375 105.200 141.435 ;
        RECT 106.275 141.390 106.565 141.435 ;
        RECT 108.575 141.575 108.865 141.620 ;
        RECT 109.020 141.575 109.340 141.635 ;
        RECT 108.575 141.435 109.340 141.575 ;
        RECT 108.575 141.390 108.865 141.435 ;
        RECT 109.020 141.375 109.340 141.435 ;
        RECT 109.480 141.375 109.800 141.635 ;
        RECT 10.510 140.755 115.850 141.235 ;
        RECT 135.635 141.220 136.775 165.470 ;
        RECT 56.580 140.555 56.900 140.615 ;
        RECT 58.895 140.555 59.185 140.600 ;
        RECT 56.580 140.415 59.185 140.555 ;
        RECT 56.580 140.355 56.900 140.415 ;
        RECT 58.895 140.370 59.185 140.415 ;
        RECT 62.560 140.355 62.880 140.615 ;
        RECT 74.060 140.355 74.380 140.615 ;
        RECT 76.375 140.370 76.665 140.600 ;
        RECT 79.120 140.555 79.440 140.615 ;
        RECT 79.595 140.555 79.885 140.600 ;
        RECT 79.120 140.415 79.885 140.555 ;
        RECT 37.720 140.015 38.040 140.275 ;
        RECT 40.495 140.215 40.785 140.260 ;
        RECT 44.160 140.215 44.480 140.275 ;
        RECT 48.760 140.215 49.080 140.275 ;
        RECT 40.495 140.075 44.480 140.215 ;
        RECT 40.495 140.030 40.785 140.075 ;
        RECT 44.160 140.015 44.480 140.075 ;
        RECT 44.710 140.075 49.080 140.215 ;
        RECT 14.260 139.875 14.580 139.935 ;
        RECT 16.115 139.875 16.405 139.920 ;
        RECT 14.260 139.735 16.405 139.875 ;
        RECT 14.260 139.675 14.580 139.735 ;
        RECT 16.115 139.690 16.405 139.735 ;
        RECT 29.440 139.875 29.760 139.935 ;
        RECT 29.915 139.875 30.205 139.920 ;
        RECT 29.440 139.735 30.205 139.875 ;
        RECT 29.440 139.675 29.760 139.735 ;
        RECT 29.915 139.690 30.205 139.735 ;
        RECT 30.360 139.675 30.680 139.935 ;
        RECT 31.295 139.690 31.585 139.920 ;
        RECT 34.040 139.875 34.360 139.935 ;
        RECT 35.895 139.875 36.185 139.920 ;
        RECT 34.040 139.735 36.185 139.875 ;
        RECT 31.370 139.195 31.510 139.690 ;
        RECT 34.040 139.675 34.360 139.735 ;
        RECT 35.895 139.690 36.185 139.735 ;
        RECT 37.275 139.690 37.565 139.920 ;
        RECT 36.800 139.335 37.120 139.595 ;
        RECT 37.350 139.535 37.490 139.690 ;
        RECT 38.640 139.675 38.960 139.935 ;
        RECT 39.100 139.675 39.420 139.935 ;
        RECT 41.400 139.675 41.720 139.935 ;
        RECT 41.875 139.875 42.165 139.920 ;
        RECT 43.700 139.875 44.020 139.935 ;
        RECT 44.710 139.920 44.850 140.075 ;
        RECT 48.760 140.015 49.080 140.075 ;
        RECT 68.555 140.215 68.845 140.260 ;
        RECT 69.015 140.215 69.305 140.260 ;
        RECT 68.555 140.075 69.305 140.215 ;
        RECT 68.555 140.030 68.845 140.075 ;
        RECT 69.015 140.030 69.305 140.075 ;
        RECT 71.390 140.075 74.750 140.215 ;
        RECT 41.875 139.735 44.020 139.875 ;
        RECT 41.875 139.690 42.165 139.735 ;
        RECT 43.700 139.675 44.020 139.735 ;
        RECT 44.635 139.690 44.925 139.920 ;
        RECT 45.080 139.675 45.400 139.935 ;
        RECT 45.540 139.675 45.860 139.935 ;
        RECT 46.460 139.675 46.780 139.935 ;
        RECT 49.220 139.875 49.540 139.935 ;
        RECT 47.010 139.735 49.540 139.875 ;
        RECT 43.255 139.535 43.545 139.580 ;
        RECT 37.350 139.395 43.545 139.535 ;
        RECT 45.170 139.535 45.310 139.675 ;
        RECT 47.010 139.535 47.150 139.735 ;
        RECT 49.220 139.675 49.540 139.735 ;
        RECT 53.835 139.875 54.125 139.920 ;
        RECT 54.740 139.875 55.060 139.935 ;
        RECT 53.835 139.735 55.060 139.875 ;
        RECT 53.835 139.690 54.125 139.735 ;
        RECT 54.740 139.675 55.060 139.735 ;
        RECT 55.660 139.875 55.980 139.935 ;
        RECT 59.355 139.875 59.645 139.920 ;
        RECT 61.655 139.875 61.945 139.920 ;
        RECT 55.660 139.735 59.645 139.875 ;
        RECT 55.660 139.675 55.980 139.735 ;
        RECT 59.355 139.690 59.645 139.735 ;
        RECT 61.270 139.735 61.945 139.875 ;
        RECT 45.170 139.395 47.150 139.535 ;
        RECT 47.840 139.535 48.160 139.595 ;
        RECT 57.975 139.535 58.265 139.580 ;
        RECT 60.720 139.535 61.040 139.595 ;
        RECT 47.840 139.395 61.040 139.535 ;
        RECT 43.255 139.350 43.545 139.395 ;
        RECT 47.840 139.335 48.160 139.395 ;
        RECT 57.975 139.350 58.265 139.395 ;
        RECT 60.720 139.335 61.040 139.395 ;
        RECT 53.360 139.195 53.680 139.255 ;
        RECT 61.270 139.240 61.410 139.735 ;
        RECT 61.655 139.690 61.945 139.735 ;
        RECT 67.175 139.875 67.465 139.920 ;
        RECT 67.620 139.875 67.940 139.935 ;
        RECT 67.175 139.735 67.940 139.875 ;
        RECT 67.175 139.690 67.465 139.735 ;
        RECT 67.620 139.675 67.940 139.735 ;
        RECT 70.380 139.675 70.700 139.935 ;
        RECT 70.840 139.675 71.160 139.935 ;
        RECT 71.390 139.920 71.530 140.075 ;
        RECT 71.315 139.690 71.605 139.920 ;
        RECT 71.760 139.875 72.080 139.935 ;
        RECT 74.610 139.920 74.750 140.075 ;
        RECT 72.235 139.875 72.525 139.920 ;
        RECT 71.760 139.735 72.525 139.875 ;
        RECT 71.760 139.675 72.080 139.735 ;
        RECT 72.235 139.690 72.525 139.735 ;
        RECT 74.535 139.690 74.825 139.920 ;
        RECT 76.450 139.875 76.590 140.370 ;
        RECT 79.120 140.355 79.440 140.415 ;
        RECT 79.595 140.370 79.885 140.415 ;
        RECT 92.460 140.555 92.780 140.615 ;
        RECT 105.340 140.555 105.660 140.615 ;
        RECT 92.460 140.415 99.130 140.555 ;
        RECT 92.460 140.355 92.780 140.415 ;
        RECT 85.115 140.215 85.405 140.260 ;
        RECT 89.700 140.215 90.020 140.275 ;
        RECT 94.315 140.215 94.605 140.260 ;
        RECT 85.115 140.075 94.605 140.215 ;
        RECT 85.115 140.030 85.405 140.075 ;
        RECT 89.700 140.015 90.020 140.075 ;
        RECT 77.755 139.875 78.045 139.920 ;
        RECT 76.450 139.735 78.045 139.875 ;
        RECT 77.755 139.690 78.045 139.735 ;
        RECT 80.055 139.875 80.345 139.920 ;
        RECT 83.260 139.875 83.580 139.935 ;
        RECT 90.405 139.875 90.695 139.920 ;
        RECT 80.055 139.735 83.580 139.875 ;
        RECT 80.055 139.690 80.345 139.735 ;
        RECT 68.095 139.535 68.385 139.580 ;
        RECT 68.095 139.395 71.530 139.535 ;
        RECT 68.095 139.350 68.385 139.395 ;
        RECT 71.390 139.255 71.530 139.395 ;
        RECT 73.600 139.335 73.920 139.595 ;
        RECT 74.610 139.535 74.750 139.690 ;
        RECT 83.260 139.675 83.580 139.735 ;
        RECT 86.570 139.735 90.695 139.875 ;
        RECT 74.610 139.395 80.270 139.535 ;
        RECT 31.370 139.055 53.680 139.195 ;
        RECT 53.360 138.995 53.680 139.055 ;
        RECT 61.195 139.010 61.485 139.240 ;
        RECT 69.000 139.195 69.320 139.255 ;
        RECT 69.000 139.055 71.070 139.195 ;
        RECT 69.000 138.995 69.320 139.055 ;
        RECT 16.560 138.655 16.880 138.915 ;
        RECT 23.460 138.855 23.780 138.915 ;
        RECT 28.995 138.855 29.285 138.900 ;
        RECT 23.460 138.715 29.285 138.855 ;
        RECT 23.460 138.655 23.780 138.715 ;
        RECT 28.995 138.670 29.285 138.715 ;
        RECT 29.440 138.855 29.760 138.915 ;
        RECT 29.915 138.855 30.205 138.900 ;
        RECT 29.440 138.715 30.205 138.855 ;
        RECT 29.440 138.655 29.760 138.715 ;
        RECT 29.915 138.670 30.205 138.715 ;
        RECT 32.200 138.855 32.520 138.915 ;
        RECT 34.975 138.855 35.265 138.900 ;
        RECT 32.200 138.715 35.265 138.855 ;
        RECT 32.200 138.655 32.520 138.715 ;
        RECT 34.975 138.670 35.265 138.715 ;
        RECT 37.260 138.655 37.580 138.915 ;
        RECT 38.180 138.655 38.500 138.915 ;
        RECT 40.035 138.855 40.325 138.900 ;
        RECT 40.940 138.855 41.260 138.915 ;
        RECT 40.035 138.715 41.260 138.855 ;
        RECT 40.035 138.670 40.325 138.715 ;
        RECT 40.940 138.655 41.260 138.715 ;
        RECT 41.860 138.655 42.180 138.915 ;
        RECT 42.795 138.855 43.085 138.900 ;
        RECT 60.260 138.855 60.580 138.915 ;
        RECT 42.795 138.715 60.580 138.855 ;
        RECT 42.795 138.670 43.085 138.715 ;
        RECT 60.260 138.655 60.580 138.715 ;
        RECT 66.255 138.855 66.545 138.900 ;
        RECT 67.620 138.855 67.940 138.915 ;
        RECT 66.255 138.715 67.940 138.855 ;
        RECT 66.255 138.670 66.545 138.715 ;
        RECT 67.620 138.655 67.940 138.715 ;
        RECT 68.555 138.855 68.845 138.900 ;
        RECT 70.380 138.855 70.700 138.915 ;
        RECT 68.555 138.715 70.700 138.855 ;
        RECT 70.930 138.855 71.070 139.055 ;
        RECT 71.300 138.995 71.620 139.255 ;
        RECT 78.675 139.195 78.965 139.240 ;
        RECT 79.580 139.195 79.900 139.255 ;
        RECT 78.675 139.055 79.900 139.195 ;
        RECT 80.130 139.195 80.270 139.395 ;
        RECT 84.180 139.335 84.500 139.595 ;
        RECT 84.640 139.335 84.960 139.595 ;
        RECT 84.730 139.195 84.870 139.335 ;
        RECT 80.130 139.055 84.870 139.195 ;
        RECT 78.675 139.010 78.965 139.055 ;
        RECT 79.580 138.995 79.900 139.055 ;
        RECT 86.570 138.855 86.710 139.735 ;
        RECT 90.405 139.690 90.695 139.735 ;
        RECT 87.400 139.535 87.720 139.595 ;
        RECT 89.255 139.535 89.545 139.580 ;
        RECT 87.400 139.395 89.545 139.535 ;
        RECT 87.400 139.335 87.720 139.395 ;
        RECT 89.255 139.350 89.545 139.395 ;
        RECT 90.480 139.195 90.620 139.690 ;
        RECT 91.080 139.675 91.400 139.935 ;
        RECT 91.630 139.920 91.770 140.075 ;
        RECT 94.315 140.030 94.605 140.075 ;
        RECT 98.990 139.935 99.130 140.415 ;
        RECT 99.450 140.415 105.660 140.555 ;
        RECT 91.630 139.735 91.950 139.920 ;
        RECT 91.660 139.690 91.950 139.735 ;
        RECT 92.460 139.675 92.780 139.935 ;
        RECT 94.775 139.875 95.065 139.920 ;
        RECT 97.980 139.875 98.300 139.935 ;
        RECT 94.775 139.735 98.300 139.875 ;
        RECT 94.775 139.690 95.065 139.735 ;
        RECT 97.980 139.675 98.300 139.735 ;
        RECT 98.900 139.675 99.220 139.935 ;
        RECT 92.920 139.535 93.240 139.595 ;
        RECT 93.855 139.535 94.145 139.580 ;
        RECT 99.450 139.535 99.590 140.415 ;
        RECT 105.340 140.355 105.660 140.415 ;
        RECT 101.660 140.215 101.980 140.275 ;
        RECT 100.370 140.075 101.980 140.215 ;
        RECT 100.370 139.920 100.510 140.075 ;
        RECT 101.660 140.015 101.980 140.075 ;
        RECT 107.130 140.215 107.420 140.260 ;
        RECT 109.480 140.215 109.800 140.275 ;
        RECT 110.390 140.215 110.680 140.260 ;
        RECT 107.130 140.075 110.680 140.215 ;
        RECT 107.130 140.030 107.420 140.075 ;
        RECT 109.480 140.015 109.800 140.075 ;
        RECT 110.390 140.030 110.680 140.075 ;
        RECT 111.310 140.215 111.600 140.260 ;
        RECT 113.170 140.215 113.460 140.260 ;
        RECT 135.580 140.230 136.830 141.220 ;
        RECT 111.310 140.075 113.460 140.215 ;
        RECT 135.635 140.155 136.775 140.230 ;
        RECT 111.310 140.030 111.600 140.075 ;
        RECT 113.170 140.030 113.460 140.075 ;
        RECT 99.835 139.690 100.125 139.920 ;
        RECT 100.295 139.690 100.585 139.920 ;
        RECT 92.920 139.395 99.590 139.535 ;
        RECT 99.910 139.535 100.050 139.690 ;
        RECT 100.740 139.675 101.060 139.935 ;
        RECT 103.040 139.875 103.360 139.935 ;
        RECT 103.515 139.875 103.805 139.920 ;
        RECT 103.040 139.735 103.805 139.875 ;
        RECT 103.040 139.675 103.360 139.735 ;
        RECT 103.515 139.690 103.805 139.735 ;
        RECT 108.990 139.875 109.280 139.920 ;
        RECT 111.310 139.875 111.525 140.030 ;
        RECT 108.990 139.735 111.525 139.875 ;
        RECT 108.990 139.690 109.280 139.735 ;
        RECT 104.880 139.580 105.200 139.595 ;
        RECT 104.880 139.535 105.415 139.580 ;
        RECT 99.910 139.395 105.415 139.535 ;
        RECT 92.920 139.335 93.240 139.395 ;
        RECT 93.855 139.350 94.145 139.395 ;
        RECT 104.880 139.350 105.415 139.395 ;
        RECT 104.880 139.335 105.200 139.350 ;
        RECT 112.240 139.335 112.560 139.595 ;
        RECT 114.080 139.335 114.400 139.595 ;
        RECT 100.280 139.195 100.600 139.255 ;
        RECT 90.480 139.055 100.600 139.195 ;
        RECT 100.280 138.995 100.600 139.055 ;
        RECT 108.990 139.195 109.280 139.240 ;
        RECT 111.770 139.195 112.060 139.240 ;
        RECT 113.630 139.195 113.920 139.240 ;
        RECT 108.990 139.055 113.920 139.195 ;
        RECT 108.990 139.010 109.280 139.055 ;
        RECT 111.770 139.010 112.060 139.055 ;
        RECT 113.630 139.010 113.920 139.055 ;
        RECT 132.510 139.190 135.210 140.010 ;
        RECT 143.370 139.390 144.510 223.840 ;
        RECT 137.240 139.380 144.510 139.390 ;
        RECT 136.210 139.190 144.510 139.380 ;
        RECT 70.930 138.715 86.710 138.855 ;
        RECT 86.955 138.855 87.245 138.900 ;
        RECT 89.240 138.855 89.560 138.915 ;
        RECT 86.955 138.715 89.560 138.855 ;
        RECT 68.555 138.670 68.845 138.715 ;
        RECT 70.380 138.655 70.700 138.715 ;
        RECT 86.955 138.670 87.245 138.715 ;
        RECT 89.240 138.655 89.560 138.715 ;
        RECT 96.615 138.855 96.905 138.900 ;
        RECT 100.740 138.855 101.060 138.915 ;
        RECT 96.615 138.715 101.060 138.855 ;
        RECT 96.615 138.670 96.905 138.715 ;
        RECT 100.740 138.655 101.060 138.715 ;
        RECT 102.120 138.655 102.440 138.915 ;
        RECT 103.975 138.855 104.265 138.900 ;
        RECT 104.420 138.855 104.740 138.915 ;
        RECT 103.975 138.715 104.740 138.855 ;
        RECT 103.975 138.670 104.265 138.715 ;
        RECT 104.420 138.655 104.740 138.715 ;
        RECT 132.510 138.530 144.510 139.190 ;
        RECT 10.510 138.035 115.850 138.515 ;
        RECT 132.510 138.190 135.210 138.530 ;
        RECT 136.210 138.250 144.510 138.530 ;
        RECT 136.210 138.240 138.350 138.250 ;
        RECT 29.440 137.635 29.760 137.895 ;
        RECT 30.360 137.835 30.680 137.895 ;
        RECT 31.755 137.835 32.045 137.880 ;
        RECT 30.360 137.695 32.045 137.835 ;
        RECT 30.360 137.635 30.680 137.695 ;
        RECT 31.755 137.650 32.045 137.695 ;
        RECT 34.500 137.635 34.820 137.895 ;
        RECT 49.695 137.835 49.985 137.880 ;
        RECT 45.170 137.695 49.985 137.835 ;
        RECT 13.360 137.495 13.650 137.540 ;
        RECT 15.220 137.495 15.510 137.540 ;
        RECT 18.000 137.495 18.290 137.540 ;
        RECT 45.170 137.495 45.310 137.695 ;
        RECT 49.695 137.650 49.985 137.695 ;
        RECT 13.360 137.355 18.290 137.495 ;
        RECT 13.360 137.310 13.650 137.355 ;
        RECT 15.220 137.310 15.510 137.355 ;
        RECT 18.000 137.310 18.290 137.355 ;
        RECT 33.210 137.355 45.310 137.495 ;
        RECT 13.800 137.155 14.120 137.215 ;
        RECT 14.735 137.155 15.025 137.200 ;
        RECT 23.920 137.155 24.240 137.215 ;
        RECT 13.800 137.015 15.025 137.155 ;
        RECT 13.800 136.955 14.120 137.015 ;
        RECT 14.735 136.970 15.025 137.015 ;
        RECT 15.270 137.015 24.240 137.155 ;
        RECT 12.895 136.815 13.185 136.860 ;
        RECT 15.270 136.815 15.410 137.015 ;
        RECT 23.920 136.955 24.240 137.015 ;
        RECT 24.380 137.155 24.700 137.215 ;
        RECT 27.615 137.155 27.905 137.200 ;
        RECT 24.380 137.015 27.905 137.155 ;
        RECT 24.380 136.955 24.700 137.015 ;
        RECT 27.615 136.970 27.905 137.015 ;
        RECT 31.280 136.955 31.600 137.215 ;
        RECT 18.000 136.815 18.290 136.860 ;
        RECT 12.895 136.675 15.410 136.815 ;
        RECT 15.755 136.675 18.290 136.815 ;
        RECT 12.895 136.630 13.185 136.675 ;
        RECT 15.755 136.520 15.970 136.675 ;
        RECT 18.000 136.630 18.290 136.675 ;
        RECT 26.220 136.615 26.540 136.875 ;
        RECT 28.520 136.615 28.840 136.875 ;
        RECT 30.820 136.615 31.140 136.875 ;
        RECT 33.210 136.815 33.350 137.355 ;
        RECT 45.555 137.310 45.845 137.540 ;
        RECT 49.770 137.495 49.910 137.650 ;
        RECT 53.360 137.635 53.680 137.895 ;
        RECT 55.200 137.835 55.520 137.895 ;
        RECT 78.200 137.835 78.520 137.895 ;
        RECT 55.200 137.695 78.520 137.835 ;
        RECT 55.200 137.635 55.520 137.695 ;
        RECT 78.200 137.635 78.520 137.695 ;
        RECT 78.905 137.835 79.195 137.880 ;
        RECT 84.640 137.835 84.960 137.895 ;
        RECT 78.905 137.695 84.960 137.835 ;
        RECT 78.905 137.650 79.195 137.695 ;
        RECT 84.640 137.635 84.960 137.695 ;
        RECT 89.700 137.835 90.020 137.895 ;
        RECT 90.405 137.835 90.695 137.880 ;
        RECT 89.700 137.695 90.695 137.835 ;
        RECT 89.700 137.635 90.020 137.695 ;
        RECT 90.405 137.650 90.695 137.695 ;
        RECT 97.980 137.835 98.300 137.895 ;
        RECT 102.365 137.835 102.655 137.880 ;
        RECT 103.960 137.835 104.280 137.895 ;
        RECT 97.980 137.695 104.280 137.835 ;
        RECT 97.980 137.635 98.300 137.695 ;
        RECT 102.365 137.650 102.655 137.695 ;
        RECT 103.960 137.635 104.280 137.695 ;
        RECT 112.240 137.835 112.560 137.895 ;
        RECT 112.715 137.835 113.005 137.880 ;
        RECT 112.240 137.695 113.005 137.835 ;
        RECT 112.240 137.635 112.560 137.695 ;
        RECT 112.715 137.650 113.005 137.695 ;
        RECT 54.740 137.495 55.060 137.555 ;
        RECT 69.000 137.495 69.320 137.555 ;
        RECT 49.770 137.355 54.510 137.495 ;
        RECT 33.580 137.155 33.900 137.215 ;
        RECT 33.580 137.015 34.730 137.155 ;
        RECT 33.580 136.955 33.900 137.015 ;
        RECT 34.055 136.815 34.345 136.860 ;
        RECT 33.210 136.675 34.345 136.815 ;
        RECT 34.590 136.815 34.730 137.015 ;
        RECT 34.960 136.955 35.280 137.215 ;
        RECT 35.435 136.815 35.725 136.860 ;
        RECT 34.590 136.675 35.725 136.815 ;
        RECT 34.055 136.630 34.345 136.675 ;
        RECT 35.435 136.630 35.725 136.675 ;
        RECT 45.095 136.815 45.385 136.860 ;
        RECT 45.630 136.815 45.770 137.310 ;
        RECT 47.840 137.155 48.160 137.215 ;
        RECT 48.315 137.155 48.605 137.200 ;
        RECT 47.840 137.015 48.605 137.155 ;
        RECT 54.370 137.155 54.510 137.355 ;
        RECT 54.740 137.355 69.320 137.495 ;
        RECT 54.740 137.295 55.060 137.355 ;
        RECT 69.000 137.295 69.320 137.355 ;
        RECT 82.770 137.495 83.060 137.540 ;
        RECT 85.550 137.495 85.840 137.540 ;
        RECT 87.410 137.495 87.700 137.540 ;
        RECT 82.770 137.355 87.700 137.495 ;
        RECT 82.770 137.310 83.060 137.355 ;
        RECT 85.550 137.310 85.840 137.355 ;
        RECT 87.410 137.310 87.700 137.355 ;
        RECT 88.335 137.310 88.625 137.540 ;
        RECT 94.270 137.495 94.560 137.540 ;
        RECT 97.050 137.495 97.340 137.540 ;
        RECT 98.910 137.495 99.200 137.540 ;
        RECT 94.270 137.355 99.200 137.495 ;
        RECT 94.270 137.310 94.560 137.355 ;
        RECT 97.050 137.310 97.340 137.355 ;
        RECT 98.910 137.310 99.200 137.355 ;
        RECT 106.230 137.495 106.520 137.540 ;
        RECT 109.010 137.495 109.300 137.540 ;
        RECT 110.870 137.495 111.160 137.540 ;
        RECT 106.230 137.355 111.160 137.495 ;
        RECT 106.230 137.310 106.520 137.355 ;
        RECT 109.010 137.310 109.300 137.355 ;
        RECT 110.870 137.310 111.160 137.355 ;
        RECT 78.660 137.155 78.980 137.215 ;
        RECT 86.035 137.155 86.325 137.200 ;
        RECT 88.410 137.155 88.550 137.310 ;
        RECT 54.370 137.015 62.330 137.155 ;
        RECT 47.840 136.955 48.160 137.015 ;
        RECT 48.315 136.970 48.605 137.015 ;
        RECT 45.095 136.675 45.770 136.815 ;
        RECT 46.000 136.815 46.320 136.875 ;
        RECT 47.395 136.815 47.685 136.860 ;
        RECT 46.000 136.675 47.685 136.815 ;
        RECT 45.095 136.630 45.385 136.675 ;
        RECT 46.000 136.615 46.320 136.675 ;
        RECT 47.395 136.630 47.685 136.675 ;
        RECT 51.075 136.630 51.365 136.860 ;
        RECT 13.820 136.475 14.110 136.520 ;
        RECT 15.680 136.475 15.970 136.520 ;
        RECT 13.820 136.335 15.970 136.475 ;
        RECT 13.820 136.290 14.110 136.335 ;
        RECT 15.680 136.290 15.970 136.335 ;
        RECT 16.560 136.520 16.880 136.535 ;
        RECT 16.560 136.475 16.890 136.520 ;
        RECT 19.860 136.475 20.150 136.520 ;
        RECT 16.560 136.335 20.150 136.475 ;
        RECT 16.560 136.290 16.890 136.335 ;
        RECT 19.860 136.290 20.150 136.335 ;
        RECT 32.215 136.475 32.505 136.520 ;
        RECT 42.780 136.475 43.100 136.535 ;
        RECT 32.215 136.335 43.100 136.475 ;
        RECT 32.215 136.290 32.505 136.335 ;
        RECT 16.560 136.275 16.880 136.290 ;
        RECT 42.780 136.275 43.100 136.335 ;
        RECT 45.540 136.475 45.860 136.535 ;
        RECT 47.855 136.475 48.145 136.520 ;
        RECT 48.760 136.475 49.080 136.535 ;
        RECT 45.540 136.335 49.080 136.475 ;
        RECT 45.540 136.275 45.860 136.335 ;
        RECT 47.855 136.290 48.145 136.335 ;
        RECT 48.760 136.275 49.080 136.335 ;
        RECT 51.150 136.195 51.290 136.630 ;
        RECT 51.520 136.615 51.840 136.875 ;
        RECT 51.995 136.815 52.285 136.860 ;
        RECT 52.440 136.815 52.760 136.875 ;
        RECT 51.995 136.675 52.760 136.815 ;
        RECT 51.995 136.630 52.285 136.675 ;
        RECT 52.440 136.615 52.760 136.675 ;
        RECT 52.915 136.815 53.205 136.860 ;
        RECT 54.280 136.815 54.600 136.875 ;
        RECT 52.915 136.675 54.600 136.815 ;
        RECT 52.915 136.630 53.205 136.675 ;
        RECT 54.280 136.615 54.600 136.675 ;
        RECT 54.740 136.615 55.060 136.875 ;
        RECT 55.200 136.615 55.520 136.875 ;
        RECT 55.660 136.615 55.980 136.875 ;
        RECT 56.595 136.815 56.885 136.860 ;
        RECT 57.500 136.815 57.820 136.875 ;
        RECT 56.210 136.675 57.820 136.815 ;
        RECT 54.830 136.475 54.970 136.615 ;
        RECT 51.840 136.335 54.970 136.475 ;
        RECT 21.865 136.135 22.155 136.180 ;
        RECT 22.540 136.135 22.860 136.195 ;
        RECT 21.865 135.995 22.860 136.135 ;
        RECT 21.865 135.950 22.155 135.995 ;
        RECT 22.540 135.935 22.860 135.995 ;
        RECT 23.000 136.135 23.320 136.195 ;
        RECT 25.315 136.135 25.605 136.180 ;
        RECT 23.000 135.995 25.605 136.135 ;
        RECT 23.000 135.935 23.320 135.995 ;
        RECT 25.315 135.950 25.605 135.995 ;
        RECT 29.900 135.935 30.220 136.195 ;
        RECT 31.280 136.135 31.600 136.195 ;
        RECT 33.135 136.135 33.425 136.180 ;
        RECT 31.280 135.995 33.425 136.135 ;
        RECT 31.280 135.935 31.600 135.995 ;
        RECT 33.135 135.950 33.425 135.995 ;
        RECT 44.175 136.135 44.465 136.180 ;
        RECT 45.080 136.135 45.400 136.195 ;
        RECT 44.175 135.995 45.400 136.135 ;
        RECT 44.175 135.950 44.465 135.995 ;
        RECT 45.080 135.935 45.400 135.995 ;
        RECT 51.060 136.135 51.380 136.195 ;
        RECT 51.840 136.135 51.980 136.335 ;
        RECT 51.060 135.995 51.980 136.135 ;
        RECT 52.900 136.135 53.220 136.195 ;
        RECT 56.210 136.135 56.350 136.675 ;
        RECT 56.595 136.630 56.885 136.675 ;
        RECT 57.500 136.615 57.820 136.675 ;
        RECT 58.420 136.815 58.740 136.875 ;
        RECT 58.895 136.815 59.185 136.860 ;
        RECT 58.420 136.675 59.185 136.815 ;
        RECT 58.420 136.615 58.740 136.675 ;
        RECT 58.895 136.630 59.185 136.675 ;
        RECT 60.275 136.630 60.565 136.860 ;
        RECT 60.720 136.815 61.040 136.875 ;
        RECT 62.190 136.860 62.330 137.015 ;
        RECT 78.660 137.015 85.790 137.155 ;
        RECT 78.660 136.955 78.980 137.015 ;
        RECT 61.195 136.815 61.485 136.860 ;
        RECT 60.720 136.675 61.485 136.815 ;
        RECT 60.350 136.475 60.490 136.630 ;
        RECT 60.720 136.615 61.040 136.675 ;
        RECT 61.195 136.630 61.485 136.675 ;
        RECT 62.115 136.630 62.405 136.860 ;
        RECT 63.020 136.615 63.340 136.875 ;
        RECT 82.770 136.815 83.060 136.860 ;
        RECT 85.650 136.815 85.790 137.015 ;
        RECT 86.035 137.015 88.550 137.155 ;
        RECT 99.375 137.155 99.665 137.200 ;
        RECT 99.375 137.015 109.250 137.155 ;
        RECT 86.035 136.970 86.325 137.015 ;
        RECT 99.375 136.970 99.665 137.015 ;
        RECT 87.875 136.815 88.165 136.860 ;
        RECT 82.770 136.675 85.305 136.815 ;
        RECT 85.650 136.675 88.165 136.815 ;
        RECT 82.770 136.630 83.060 136.675 ;
        RECT 56.670 136.335 60.490 136.475 ;
        RECT 61.640 136.475 61.960 136.535 ;
        RECT 63.110 136.475 63.250 136.615 ;
        RECT 61.640 136.335 63.250 136.475 ;
        RECT 80.910 136.475 81.200 136.520 ;
        RECT 83.260 136.475 83.580 136.535 ;
        RECT 85.090 136.520 85.305 136.675 ;
        RECT 87.875 136.630 88.165 136.675 ;
        RECT 89.240 136.615 89.560 136.875 ;
        RECT 94.270 136.815 94.560 136.860 ;
        RECT 97.535 136.815 97.825 136.860 ;
        RECT 94.270 136.675 96.805 136.815 ;
        RECT 94.270 136.630 94.560 136.675 ;
        RECT 84.170 136.475 84.460 136.520 ;
        RECT 80.910 136.335 84.460 136.475 ;
        RECT 56.670 136.195 56.810 136.335 ;
        RECT 61.640 136.275 61.960 136.335 ;
        RECT 80.910 136.290 81.200 136.335 ;
        RECT 83.260 136.275 83.580 136.335 ;
        RECT 84.170 136.290 84.460 136.335 ;
        RECT 85.090 136.475 85.380 136.520 ;
        RECT 86.950 136.475 87.240 136.520 ;
        RECT 85.090 136.335 87.240 136.475 ;
        RECT 85.090 136.290 85.380 136.335 ;
        RECT 86.950 136.290 87.240 136.335 ;
        RECT 91.540 136.475 91.860 136.535 ;
        RECT 96.590 136.520 96.805 136.675 ;
        RECT 97.535 136.675 100.050 136.815 ;
        RECT 97.535 136.630 97.825 136.675 ;
        RECT 92.410 136.475 92.700 136.520 ;
        RECT 95.670 136.475 95.960 136.520 ;
        RECT 91.540 136.335 95.960 136.475 ;
        RECT 91.540 136.275 91.860 136.335 ;
        RECT 92.410 136.290 92.700 136.335 ;
        RECT 95.670 136.290 95.960 136.335 ;
        RECT 96.590 136.475 96.880 136.520 ;
        RECT 98.450 136.475 98.740 136.520 ;
        RECT 96.590 136.335 98.740 136.475 ;
        RECT 96.590 136.290 96.880 136.335 ;
        RECT 98.450 136.290 98.740 136.335 ;
        RECT 52.900 135.995 56.350 136.135 ;
        RECT 51.060 135.935 51.380 135.995 ;
        RECT 52.900 135.935 53.220 135.995 ;
        RECT 56.580 135.935 56.900 136.195 ;
        RECT 59.340 135.935 59.660 136.195 ;
        RECT 63.035 136.135 63.325 136.180 ;
        RECT 64.400 136.135 64.720 136.195 ;
        RECT 99.910 136.180 100.050 136.675 ;
        RECT 100.740 136.615 101.060 136.875 ;
        RECT 106.230 136.815 106.520 136.860 ;
        RECT 109.110 136.815 109.250 137.015 ;
        RECT 109.480 136.955 109.800 137.215 ;
        RECT 114.080 137.155 114.400 137.215 ;
        RECT 111.410 137.015 114.400 137.155 ;
        RECT 111.410 136.860 111.550 137.015 ;
        RECT 114.080 136.955 114.400 137.015 ;
        RECT 111.335 136.815 111.625 136.860 ;
        RECT 106.230 136.675 108.765 136.815 ;
        RECT 109.110 136.675 111.625 136.815 ;
        RECT 106.230 136.630 106.520 136.675 ;
        RECT 104.420 136.520 104.740 136.535 ;
        RECT 108.550 136.520 108.765 136.675 ;
        RECT 111.335 136.630 111.625 136.675 ;
        RECT 111.795 136.630 112.085 136.860 ;
        RECT 104.370 136.475 104.740 136.520 ;
        RECT 107.630 136.475 107.920 136.520 ;
        RECT 104.370 136.335 107.920 136.475 ;
        RECT 104.370 136.290 104.740 136.335 ;
        RECT 107.630 136.290 107.920 136.335 ;
        RECT 108.550 136.475 108.840 136.520 ;
        RECT 110.410 136.475 110.700 136.520 ;
        RECT 108.550 136.335 110.700 136.475 ;
        RECT 108.550 136.290 108.840 136.335 ;
        RECT 110.410 136.290 110.700 136.335 ;
        RECT 104.420 136.275 104.740 136.290 ;
        RECT 63.035 135.995 64.720 136.135 ;
        RECT 63.035 135.950 63.325 135.995 ;
        RECT 64.400 135.935 64.720 135.995 ;
        RECT 99.835 135.950 100.125 136.180 ;
        RECT 109.020 136.135 109.340 136.195 ;
        RECT 111.870 136.135 112.010 136.630 ;
        RECT 109.020 135.995 112.010 136.135 ;
        RECT 109.020 135.935 109.340 135.995 ;
        RECT 10.510 135.315 115.850 135.795 ;
        RECT 13.800 134.915 14.120 135.175 ;
        RECT 25.775 135.115 26.065 135.160 ;
        RECT 26.220 135.115 26.540 135.175 ;
        RECT 25.775 134.975 26.540 135.115 ;
        RECT 25.775 134.930 26.065 134.975 ;
        RECT 26.220 134.915 26.540 134.975 ;
        RECT 31.740 134.915 32.060 135.175 ;
        RECT 34.500 135.115 34.820 135.175 ;
        RECT 36.355 135.115 36.645 135.160 ;
        RECT 34.500 134.975 36.645 135.115 ;
        RECT 34.500 134.915 34.820 134.975 ;
        RECT 36.355 134.930 36.645 134.975 ;
        RECT 41.860 135.115 42.180 135.175 ;
        RECT 42.335 135.115 42.625 135.160 ;
        RECT 41.860 134.975 42.625 135.115 ;
        RECT 41.860 134.915 42.180 134.975 ;
        RECT 42.335 134.930 42.625 134.975 ;
        RECT 42.780 135.115 43.100 135.175 ;
        RECT 47.395 135.115 47.685 135.160 ;
        RECT 51.060 135.115 51.380 135.175 ;
        RECT 42.780 134.975 47.685 135.115 ;
        RECT 42.780 134.915 43.100 134.975 ;
        RECT 47.395 134.930 47.685 134.975 ;
        RECT 49.310 134.975 51.380 135.115 ;
        RECT 14.735 134.775 15.025 134.820 ;
        RECT 17.890 134.775 18.180 134.820 ;
        RECT 21.150 134.775 21.440 134.820 ;
        RECT 14.735 134.635 21.440 134.775 ;
        RECT 14.735 134.590 15.025 134.635 ;
        RECT 17.890 134.590 18.180 134.635 ;
        RECT 21.150 134.590 21.440 134.635 ;
        RECT 22.070 134.775 22.360 134.820 ;
        RECT 23.930 134.775 24.220 134.820 ;
        RECT 22.070 134.635 24.220 134.775 ;
        RECT 22.070 134.590 22.360 134.635 ;
        RECT 23.930 134.590 24.220 134.635 ;
        RECT 28.075 134.775 28.365 134.820 ;
        RECT 34.055 134.775 34.345 134.820 ;
        RECT 43.715 134.775 44.005 134.820 ;
        RECT 49.310 134.775 49.450 134.975 ;
        RECT 51.060 134.915 51.380 134.975 ;
        RECT 56.580 134.915 56.900 135.175 ;
        RECT 57.960 135.115 58.280 135.175 ;
        RECT 57.960 134.975 70.150 135.115 ;
        RECT 57.960 134.915 58.280 134.975 ;
        RECT 51.980 134.775 52.300 134.835 ;
        RECT 28.075 134.635 33.810 134.775 ;
        RECT 28.075 134.590 28.365 134.635 ;
        RECT 12.880 134.235 13.200 134.495 ;
        RECT 14.260 134.235 14.580 134.495 ;
        RECT 19.750 134.435 20.040 134.480 ;
        RECT 22.070 134.435 22.285 134.590 ;
        RECT 19.750 134.295 22.285 134.435 ;
        RECT 19.750 134.250 20.040 134.295 ;
        RECT 23.000 134.235 23.320 134.495 ;
        RECT 24.380 134.435 24.700 134.495 ;
        RECT 27.615 134.435 27.905 134.480 ;
        RECT 23.550 134.295 27.905 134.435 ;
        RECT 23.550 134.095 23.690 134.295 ;
        RECT 24.380 134.235 24.700 134.295 ;
        RECT 27.615 134.250 27.905 134.295 ;
        RECT 32.660 134.235 32.980 134.495 ;
        RECT 33.120 134.235 33.440 134.495 ;
        RECT 33.670 134.435 33.810 134.635 ;
        RECT 34.055 134.635 44.005 134.775 ;
        RECT 34.055 134.590 34.345 134.635 ;
        RECT 43.715 134.590 44.005 134.635 ;
        RECT 45.170 134.635 49.450 134.775 ;
        RECT 49.770 134.635 52.300 134.775 ;
        RECT 45.170 134.480 45.310 134.635 ;
        RECT 35.435 134.435 35.725 134.480 ;
        RECT 33.670 134.295 34.270 134.435 ;
        RECT 19.410 133.955 23.690 134.095 ;
        RECT 23.920 134.095 24.240 134.155 ;
        RECT 24.855 134.095 25.145 134.140 ;
        RECT 23.920 133.955 25.145 134.095 ;
        RECT 19.410 133.475 19.550 133.955 ;
        RECT 23.920 133.895 24.240 133.955 ;
        RECT 24.855 133.910 25.145 133.955 ;
        RECT 27.140 134.095 27.460 134.155 ;
        RECT 28.535 134.095 28.825 134.140 ;
        RECT 33.580 134.095 33.900 134.155 ;
        RECT 27.140 133.955 33.900 134.095 ;
        RECT 34.130 134.095 34.270 134.295 ;
        RECT 35.435 134.295 36.110 134.435 ;
        RECT 35.435 134.250 35.725 134.295 ;
        RECT 35.970 134.155 36.110 134.295 ;
        RECT 41.415 134.250 41.705 134.480 ;
        RECT 45.095 134.250 45.385 134.480 ;
        RECT 45.555 134.250 45.845 134.480 ;
        RECT 46.015 134.250 46.305 134.480 ;
        RECT 34.500 134.095 34.820 134.155 ;
        RECT 34.130 133.955 34.820 134.095 ;
        RECT 27.140 133.895 27.460 133.955 ;
        RECT 28.535 133.910 28.825 133.955 ;
        RECT 33.580 133.895 33.900 133.955 ;
        RECT 34.500 133.895 34.820 133.955 ;
        RECT 35.880 133.895 36.200 134.155 ;
        RECT 40.480 133.895 40.800 134.155 ;
        RECT 41.490 134.095 41.630 134.250 ;
        RECT 41.860 134.095 42.180 134.155 ;
        RECT 41.490 133.955 42.180 134.095 ;
        RECT 41.860 133.895 42.180 133.955 ;
        RECT 19.750 133.755 20.040 133.800 ;
        RECT 22.530 133.755 22.820 133.800 ;
        RECT 24.390 133.755 24.680 133.800 ;
        RECT 19.750 133.615 24.680 133.755 ;
        RECT 19.750 133.570 20.040 133.615 ;
        RECT 22.530 133.570 22.820 133.615 ;
        RECT 24.390 133.570 24.680 133.615 ;
        RECT 33.120 133.755 33.440 133.815 ;
        RECT 45.630 133.755 45.770 134.250 ;
        RECT 46.090 134.095 46.230 134.250 ;
        RECT 46.920 134.235 47.240 134.495 ;
        RECT 48.850 134.480 48.990 134.635 ;
        RECT 48.775 134.250 49.065 134.480 ;
        RECT 49.220 134.235 49.540 134.495 ;
        RECT 49.770 134.480 49.910 134.635 ;
        RECT 51.980 134.575 52.300 134.635 ;
        RECT 55.660 134.775 55.980 134.835 ;
        RECT 59.340 134.820 59.660 134.835 ;
        RECT 57.285 134.775 57.575 134.820 ;
        RECT 55.660 134.635 57.575 134.775 ;
        RECT 55.660 134.575 55.980 134.635 ;
        RECT 57.285 134.590 57.575 134.635 ;
        RECT 59.290 134.775 59.660 134.820 ;
        RECT 62.550 134.775 62.840 134.820 ;
        RECT 59.290 134.635 62.840 134.775 ;
        RECT 59.290 134.590 59.660 134.635 ;
        RECT 62.550 134.590 62.840 134.635 ;
        RECT 63.470 134.775 63.760 134.820 ;
        RECT 65.330 134.775 65.620 134.820 ;
        RECT 63.470 134.635 65.620 134.775 ;
        RECT 70.010 134.775 70.150 134.975 ;
        RECT 70.380 134.915 70.700 135.175 ;
        RECT 82.815 135.115 83.105 135.160 ;
        RECT 83.260 135.115 83.580 135.175 ;
        RECT 89.715 135.115 90.005 135.160 ;
        RECT 90.160 135.115 90.480 135.175 ;
        RECT 82.815 134.975 83.580 135.115 ;
        RECT 82.815 134.930 83.105 134.975 ;
        RECT 83.260 134.915 83.580 134.975 ;
        RECT 87.030 134.975 89.470 135.115 ;
        RECT 87.030 134.775 87.170 134.975 ;
        RECT 70.010 134.635 87.170 134.775 ;
        RECT 63.470 134.590 63.760 134.635 ;
        RECT 65.330 134.590 65.620 134.635 ;
        RECT 59.340 134.575 59.660 134.590 ;
        RECT 49.695 134.250 49.985 134.480 ;
        RECT 50.615 134.435 50.905 134.480 ;
        RECT 52.900 134.435 53.220 134.495 ;
        RECT 50.615 134.295 53.220 134.435 ;
        RECT 50.615 134.250 50.905 134.295 ;
        RECT 48.300 134.095 48.620 134.155 ;
        RECT 46.090 133.955 48.620 134.095 ;
        RECT 48.300 133.895 48.620 133.955 ;
        RECT 49.310 133.755 49.450 134.235 ;
        RECT 33.120 133.615 33.810 133.755 ;
        RECT 45.630 133.615 49.450 133.755 ;
        RECT 33.120 133.555 33.440 133.615 ;
        RECT 15.885 133.415 16.175 133.460 ;
        RECT 19.320 133.415 19.640 133.475 ;
        RECT 33.670 133.460 33.810 133.615 ;
        RECT 15.885 133.275 19.640 133.415 ;
        RECT 15.885 133.230 16.175 133.275 ;
        RECT 19.320 133.215 19.640 133.275 ;
        RECT 33.595 133.230 33.885 133.460 ;
        RECT 46.920 133.415 47.240 133.475 ;
        RECT 50.690 133.415 50.830 134.250 ;
        RECT 52.900 134.235 53.220 134.295 ;
        RECT 53.835 134.435 54.125 134.480 ;
        RECT 55.750 134.435 55.890 134.575 ;
        RECT 53.835 134.295 55.890 134.435 ;
        RECT 61.150 134.435 61.440 134.480 ;
        RECT 63.470 134.435 63.685 134.590 ;
        RECT 87.400 134.575 87.720 134.835 ;
        RECT 87.860 134.775 88.180 134.835 ;
        RECT 89.330 134.775 89.470 134.975 ;
        RECT 89.715 134.975 90.480 135.115 ;
        RECT 89.715 134.930 90.005 134.975 ;
        RECT 90.160 134.915 90.480 134.975 ;
        RECT 91.540 134.915 91.860 135.175 ;
        RECT 94.760 135.115 95.080 135.175 ;
        RECT 95.235 135.115 95.525 135.160 ;
        RECT 94.760 134.975 95.525 135.115 ;
        RECT 94.760 134.915 95.080 134.975 ;
        RECT 95.235 134.930 95.525 134.975 ;
        RECT 99.375 135.115 99.665 135.160 ;
        RECT 99.820 135.115 100.140 135.175 ;
        RECT 99.375 134.975 100.140 135.115 ;
        RECT 99.375 134.930 99.665 134.975 ;
        RECT 99.820 134.915 100.140 134.975 ;
        RECT 100.280 134.915 100.600 135.175 ;
        RECT 103.960 135.115 104.280 135.175 ;
        RECT 104.435 135.115 104.725 135.160 ;
        RECT 103.960 134.975 104.725 135.115 ;
        RECT 103.960 134.915 104.280 134.975 ;
        RECT 104.435 134.930 104.725 134.975 ;
        RECT 104.880 134.915 105.200 135.175 ;
        RECT 106.735 135.115 107.025 135.160 ;
        RECT 108.575 135.115 108.865 135.160 ;
        RECT 109.480 135.115 109.800 135.175 ;
        RECT 106.735 134.975 107.870 135.115 ;
        RECT 106.735 134.930 107.025 134.975 ;
        RECT 92.460 134.775 92.780 134.835 ;
        RECT 87.860 134.635 89.010 134.775 ;
        RECT 89.330 134.635 92.780 134.775 ;
        RECT 87.860 134.575 88.180 134.635 ;
        RECT 61.150 134.295 63.685 134.435 ;
        RECT 53.835 134.250 54.125 134.295 ;
        RECT 61.150 134.250 61.440 134.295 ;
        RECT 64.400 134.235 64.720 134.495 ;
        RECT 69.015 134.435 69.305 134.480 ;
        RECT 69.015 134.295 70.610 134.435 ;
        RECT 69.015 134.250 69.305 134.295 ;
        RECT 63.480 134.095 63.800 134.155 ;
        RECT 66.255 134.095 66.545 134.140 ;
        RECT 63.480 133.955 66.545 134.095 ;
        RECT 63.480 133.895 63.800 133.955 ;
        RECT 66.255 133.910 66.545 133.955 ;
        RECT 68.095 133.910 68.385 134.140 ;
        RECT 61.150 133.755 61.440 133.800 ;
        RECT 63.930 133.755 64.220 133.800 ;
        RECT 65.790 133.755 66.080 133.800 ;
        RECT 61.150 133.615 66.080 133.755 ;
        RECT 68.170 133.755 68.310 133.910 ;
        RECT 69.920 133.895 70.240 134.155 ;
        RECT 70.470 134.095 70.610 134.295 ;
        RECT 71.315 134.250 71.605 134.480 ;
        RECT 83.275 134.435 83.565 134.480 ;
        RECT 83.720 134.435 84.040 134.495 ;
        RECT 88.870 134.480 89.010 134.635 ;
        RECT 92.460 134.575 92.780 134.635 ;
        RECT 92.935 134.775 93.225 134.820 ;
        RECT 95.695 134.775 95.985 134.820 ;
        RECT 100.370 134.775 100.510 134.915 ;
        RECT 92.935 134.635 95.985 134.775 ;
        RECT 92.935 134.590 93.225 134.635 ;
        RECT 95.695 134.590 95.985 134.635 ;
        RECT 97.150 134.635 100.510 134.775 ;
        RECT 83.275 134.295 84.040 134.435 ;
        RECT 83.275 134.250 83.565 134.295 ;
        RECT 70.840 134.095 71.160 134.155 ;
        RECT 71.390 134.095 71.530 134.250 ;
        RECT 83.720 134.235 84.040 134.295 ;
        RECT 88.795 134.250 89.085 134.480 ;
        RECT 91.095 134.250 91.385 134.480 ;
        RECT 70.470 133.955 71.530 134.095 ;
        RECT 70.840 133.895 71.160 133.955 ;
        RECT 72.220 133.895 72.540 134.155 ;
        RECT 73.600 133.755 73.920 133.815 ;
        RECT 68.170 133.615 73.920 133.755 ;
        RECT 83.810 133.755 83.950 134.235 ;
        RECT 88.335 134.095 88.625 134.140 ;
        RECT 90.620 134.095 90.940 134.155 ;
        RECT 88.335 133.955 90.940 134.095 ;
        RECT 88.335 133.910 88.625 133.955 ;
        RECT 90.620 133.895 90.940 133.955 ;
        RECT 86.020 133.755 86.340 133.815 ;
        RECT 91.170 133.755 91.310 134.250 ;
        RECT 94.300 134.235 94.620 134.495 ;
        RECT 97.150 134.480 97.290 134.635 ;
        RECT 101.200 134.575 101.520 134.835 ;
        RECT 101.675 134.775 101.965 134.820 ;
        RECT 102.120 134.775 102.440 134.835 ;
        RECT 101.675 134.635 102.440 134.775 ;
        RECT 101.675 134.590 101.965 134.635 ;
        RECT 102.120 134.575 102.440 134.635 ;
        RECT 97.075 134.250 97.365 134.480 ;
        RECT 97.535 134.250 97.825 134.480 ;
        RECT 93.855 133.910 94.145 134.140 ;
        RECT 97.610 134.095 97.750 134.250 ;
        RECT 97.980 134.235 98.300 134.495 ;
        RECT 98.900 134.235 99.220 134.495 ;
        RECT 100.295 134.435 100.585 134.480 ;
        RECT 101.290 134.435 101.430 134.575 ;
        RECT 107.730 134.480 107.870 134.975 ;
        RECT 108.575 134.975 109.800 135.115 ;
        RECT 108.575 134.930 108.865 134.975 ;
        RECT 109.480 134.915 109.800 134.975 ;
        RECT 135.660 134.480 136.800 134.510 ;
        RECT 100.295 134.295 101.430 134.435 ;
        RECT 100.295 134.250 100.585 134.295 ;
        RECT 107.655 134.250 107.945 134.480 ;
        RECT 100.740 134.095 101.060 134.155 ;
        RECT 97.610 133.955 101.060 134.095 ;
        RECT 83.810 133.615 91.310 133.755 ;
        RECT 93.930 133.755 94.070 133.910 ;
        RECT 100.740 133.895 101.060 133.955 ;
        RECT 101.215 133.910 101.505 134.140 ;
        RECT 103.975 134.095 104.265 134.140 ;
        RECT 105.340 134.095 105.660 134.155 ;
        RECT 103.975 133.955 105.660 134.095 ;
        RECT 103.975 133.910 104.265 133.955 ;
        RECT 97.520 133.755 97.840 133.815 ;
        RECT 93.930 133.615 97.840 133.755 ;
        RECT 101.290 133.755 101.430 133.910 ;
        RECT 105.340 133.895 105.660 133.955 ;
        RECT 105.800 133.755 106.120 133.815 ;
        RECT 101.290 133.615 106.120 133.755 ;
        RECT 61.150 133.570 61.440 133.615 ;
        RECT 63.930 133.570 64.220 133.615 ;
        RECT 65.790 133.570 66.080 133.615 ;
        RECT 73.600 133.555 73.920 133.615 ;
        RECT 86.020 133.555 86.340 133.615 ;
        RECT 97.520 133.555 97.840 133.615 ;
        RECT 105.800 133.555 106.120 133.615 ;
        RECT 46.920 133.275 50.830 133.415 ;
        RECT 46.920 133.215 47.240 133.275 ;
        RECT 88.780 133.215 89.100 133.475 ;
        RECT 93.380 133.215 93.700 133.475 ;
        RECT 98.900 133.415 99.220 133.475 ;
        RECT 100.295 133.415 100.585 133.460 ;
        RECT 98.900 133.275 100.585 133.415 ;
        RECT 135.590 133.400 136.850 134.480 ;
        RECT 98.900 133.215 99.220 133.275 ;
        RECT 100.295 133.230 100.585 133.275 ;
        RECT 10.510 132.595 115.850 133.075 ;
        RECT 12.880 132.395 13.200 132.455 ;
        RECT 17.035 132.395 17.325 132.440 ;
        RECT 27.140 132.395 27.460 132.455 ;
        RECT 12.880 132.255 17.325 132.395 ;
        RECT 12.880 132.195 13.200 132.255 ;
        RECT 17.035 132.210 17.325 132.255 ;
        RECT 19.870 132.255 27.460 132.395 ;
        RECT 18.860 132.055 19.180 132.115 ;
        RECT 19.870 132.055 20.010 132.255 ;
        RECT 27.140 132.195 27.460 132.255 ;
        RECT 28.535 132.395 28.825 132.440 ;
        RECT 30.360 132.395 30.680 132.455 ;
        RECT 28.535 132.255 30.680 132.395 ;
        RECT 28.535 132.210 28.825 132.255 ;
        RECT 30.360 132.195 30.680 132.255 ;
        RECT 30.820 132.395 31.140 132.455 ;
        RECT 35.880 132.395 36.200 132.455 ;
        RECT 42.795 132.395 43.085 132.440 ;
        RECT 43.240 132.395 43.560 132.455 ;
        RECT 30.820 132.255 41.630 132.395 ;
        RECT 30.820 132.195 31.140 132.255 ;
        RECT 35.880 132.195 36.200 132.255 ;
        RECT 13.890 131.915 20.010 132.055 ;
        RECT 13.890 131.760 14.030 131.915 ;
        RECT 18.860 131.855 19.180 131.915 ;
        RECT 13.815 131.530 14.105 131.760 ;
        RECT 19.320 131.515 19.640 131.775 ;
        RECT 19.870 131.760 20.010 131.915 ;
        RECT 22.080 132.055 22.400 132.115 ;
        RECT 22.080 131.915 41.170 132.055 ;
        RECT 22.080 131.855 22.400 131.915 ;
        RECT 19.795 131.530 20.085 131.760 ;
        RECT 28.520 131.715 28.840 131.775 ;
        RECT 30.360 131.715 30.680 131.775 ;
        RECT 27.690 131.575 30.680 131.715 ;
        RECT 14.275 131.375 14.565 131.420 ;
        RECT 17.940 131.375 18.260 131.435 ;
        RECT 14.275 131.235 18.260 131.375 ;
        RECT 14.275 131.190 14.565 131.235 ;
        RECT 17.940 131.175 18.260 131.235 ;
        RECT 26.680 131.175 27.000 131.435 ;
        RECT 27.690 131.420 27.830 131.575 ;
        RECT 28.520 131.515 28.840 131.575 ;
        RECT 30.360 131.515 30.680 131.575 ;
        RECT 32.215 131.715 32.505 131.760 ;
        RECT 33.580 131.715 33.900 131.775 ;
        RECT 41.030 131.760 41.170 131.915 ;
        RECT 32.215 131.575 33.900 131.715 ;
        RECT 32.215 131.530 32.505 131.575 ;
        RECT 33.580 131.515 33.900 131.575 ;
        RECT 40.955 131.530 41.245 131.760 ;
        RECT 41.490 131.715 41.630 132.255 ;
        RECT 42.795 132.255 43.560 132.395 ;
        RECT 42.795 132.210 43.085 132.255 ;
        RECT 43.240 132.195 43.560 132.255 ;
        RECT 48.760 132.395 49.080 132.455 ;
        RECT 52.225 132.395 52.515 132.440 ;
        RECT 48.760 132.255 52.515 132.395 ;
        RECT 48.760 132.195 49.080 132.255 ;
        RECT 52.225 132.210 52.515 132.255 ;
        RECT 66.255 132.395 66.545 132.440 ;
        RECT 67.160 132.395 67.480 132.455 ;
        RECT 66.255 132.255 67.480 132.395 ;
        RECT 66.255 132.210 66.545 132.255 ;
        RECT 67.160 132.195 67.480 132.255 ;
        RECT 68.540 132.195 68.860 132.455 ;
        RECT 98.900 132.195 99.220 132.455 ;
        RECT 99.360 132.195 99.680 132.455 ;
        RECT 43.720 132.055 44.010 132.100 ;
        RECT 45.580 132.055 45.870 132.100 ;
        RECT 48.360 132.055 48.650 132.100 ;
        RECT 87.860 132.055 88.180 132.115 ;
        RECT 43.720 131.915 48.650 132.055 ;
        RECT 43.720 131.870 44.010 131.915 ;
        RECT 45.580 131.870 45.870 131.915 ;
        RECT 48.360 131.870 48.650 131.915 ;
        RECT 59.890 131.915 88.180 132.055 ;
        RECT 41.490 131.575 43.930 131.715 ;
        RECT 27.615 131.190 27.905 131.420 ;
        RECT 40.480 131.375 40.800 131.435 ;
        RECT 28.150 131.235 40.800 131.375 ;
        RECT 14.735 131.035 15.025 131.080 ;
        RECT 22.080 131.035 22.400 131.095 ;
        RECT 14.735 130.895 22.400 131.035 ;
        RECT 14.735 130.850 15.025 130.895 ;
        RECT 22.080 130.835 22.400 130.895 ;
        RECT 16.575 130.695 16.865 130.740 ;
        RECT 17.020 130.695 17.340 130.755 ;
        RECT 16.575 130.555 17.340 130.695 ;
        RECT 16.575 130.510 16.865 130.555 ;
        RECT 17.020 130.495 17.340 130.555 ;
        RECT 17.940 130.695 18.260 130.755 ;
        RECT 18.875 130.695 19.165 130.740 ;
        RECT 22.540 130.695 22.860 130.755 ;
        RECT 28.150 130.695 28.290 131.235 ;
        RECT 40.480 131.175 40.800 131.235 ;
        RECT 41.875 131.190 42.165 131.420 ;
        RECT 28.520 131.035 28.840 131.095 ;
        RECT 31.295 131.035 31.585 131.080 ;
        RECT 28.520 130.895 31.585 131.035 ;
        RECT 28.520 130.835 28.840 130.895 ;
        RECT 31.295 130.850 31.585 130.895 ;
        RECT 41.950 130.755 42.090 131.190 ;
        RECT 43.240 131.175 43.560 131.435 ;
        RECT 43.790 131.375 43.930 131.575 ;
        RECT 45.080 131.515 45.400 131.775 ;
        RECT 59.890 131.760 60.030 131.915 ;
        RECT 87.860 131.855 88.180 131.915 ;
        RECT 59.815 131.715 60.105 131.760 ;
        RECT 45.630 131.575 60.105 131.715 ;
        RECT 45.630 131.375 45.770 131.575 ;
        RECT 59.815 131.530 60.105 131.575 ;
        RECT 61.640 131.515 61.960 131.775 ;
        RECT 70.395 131.715 70.685 131.760 ;
        RECT 71.760 131.715 72.080 131.775 ;
        RECT 67.250 131.575 69.690 131.715 ;
        RECT 48.360 131.375 48.650 131.420 ;
        RECT 43.790 131.235 45.770 131.375 ;
        RECT 46.115 131.235 48.650 131.375 ;
        RECT 46.115 131.080 46.330 131.235 ;
        RECT 48.360 131.190 48.650 131.235 ;
        RECT 60.735 131.375 61.025 131.420 ;
        RECT 62.575 131.375 62.865 131.420 ;
        RECT 64.860 131.375 65.180 131.435 ;
        RECT 67.250 131.420 67.390 131.575 ;
        RECT 69.550 131.420 69.690 131.575 ;
        RECT 70.395 131.575 72.080 131.715 ;
        RECT 70.395 131.530 70.685 131.575 ;
        RECT 71.760 131.515 72.080 131.575 ;
        RECT 72.235 131.530 72.525 131.760 ;
        RECT 87.950 131.715 88.090 131.855 ;
        RECT 87.950 131.575 98.210 131.715 ;
        RECT 67.175 131.375 67.465 131.420 ;
        RECT 60.735 131.235 65.180 131.375 ;
        RECT 60.735 131.190 61.025 131.235 ;
        RECT 62.575 131.190 62.865 131.235 ;
        RECT 64.860 131.175 65.180 131.235 ;
        RECT 65.870 131.235 67.465 131.375 ;
        RECT 44.180 131.035 44.470 131.080 ;
        RECT 46.040 131.035 46.330 131.080 ;
        RECT 44.180 130.895 46.330 131.035 ;
        RECT 44.180 130.850 44.470 130.895 ;
        RECT 46.040 130.850 46.330 130.895 ;
        RECT 46.920 131.080 47.240 131.095 ;
        RECT 65.870 131.080 66.010 131.235 ;
        RECT 67.175 131.190 67.465 131.235 ;
        RECT 68.095 131.190 68.385 131.420 ;
        RECT 69.475 131.375 69.765 131.420 ;
        RECT 70.840 131.375 71.160 131.435 ;
        RECT 69.475 131.235 71.160 131.375 ;
        RECT 69.475 131.190 69.765 131.235 ;
        RECT 46.920 131.035 47.250 131.080 ;
        RECT 50.220 131.035 50.510 131.080 ;
        RECT 65.795 131.035 66.085 131.080 ;
        RECT 46.920 130.895 50.510 131.035 ;
        RECT 46.920 130.850 47.250 130.895 ;
        RECT 50.220 130.850 50.510 130.895 ;
        RECT 59.200 130.895 66.085 131.035 ;
        RECT 68.170 131.035 68.310 131.190 ;
        RECT 70.840 131.175 71.160 131.235 ;
        RECT 71.300 131.375 71.620 131.435 ;
        RECT 72.310 131.375 72.450 131.530 ;
        RECT 71.300 131.235 72.450 131.375 ;
        RECT 71.300 131.175 71.620 131.235 ;
        RECT 97.520 131.175 97.840 131.435 ;
        RECT 98.070 131.420 98.210 131.575 ;
        RECT 97.995 131.375 98.285 131.420 ;
        RECT 100.295 131.375 100.585 131.420 ;
        RECT 97.995 131.235 100.585 131.375 ;
        RECT 97.995 131.190 98.285 131.235 ;
        RECT 100.295 131.190 100.585 131.235 ;
        RECT 101.215 131.375 101.505 131.420 ;
        RECT 101.660 131.375 101.980 131.435 ;
        RECT 101.215 131.235 101.980 131.375 ;
        RECT 101.215 131.190 101.505 131.235 ;
        RECT 101.660 131.175 101.980 131.235 ;
        RECT 70.380 131.035 70.700 131.095 ;
        RECT 73.155 131.035 73.445 131.080 ;
        RECT 68.170 130.895 73.445 131.035 ;
        RECT 46.920 130.835 47.240 130.850 ;
        RECT 17.940 130.555 28.290 130.695 ;
        RECT 28.995 130.695 29.285 130.740 ;
        RECT 30.360 130.695 30.680 130.755 ;
        RECT 28.995 130.555 30.680 130.695 ;
        RECT 17.940 130.495 18.260 130.555 ;
        RECT 18.875 130.510 19.165 130.555 ;
        RECT 22.540 130.495 22.860 130.555 ;
        RECT 28.995 130.510 29.285 130.555 ;
        RECT 30.360 130.495 30.680 130.555 ;
        RECT 30.835 130.695 31.125 130.740 ;
        RECT 34.500 130.695 34.820 130.755 ;
        RECT 30.835 130.555 34.820 130.695 ;
        RECT 30.835 130.510 31.125 130.555 ;
        RECT 34.500 130.495 34.820 130.555 ;
        RECT 41.860 130.695 42.180 130.755 ;
        RECT 59.200 130.695 59.340 130.895 ;
        RECT 65.795 130.850 66.085 130.895 ;
        RECT 70.380 130.835 70.700 130.895 ;
        RECT 73.155 130.850 73.445 130.895 ;
        RECT 73.600 131.035 73.920 131.095 ;
        RECT 82.340 131.035 82.660 131.095 ;
        RECT 73.600 130.895 82.660 131.035 ;
        RECT 73.600 130.835 73.920 130.895 ;
        RECT 82.340 130.835 82.660 130.895 ;
        RECT 41.860 130.555 59.340 130.695 ;
        RECT 63.020 130.695 63.340 130.755 ;
        RECT 63.495 130.695 63.785 130.740 ;
        RECT 63.020 130.555 63.785 130.695 ;
        RECT 41.860 130.495 42.180 130.555 ;
        RECT 63.020 130.495 63.340 130.555 ;
        RECT 63.495 130.510 63.785 130.555 ;
        RECT 75.455 130.695 75.745 130.740 ;
        RECT 78.200 130.695 78.520 130.755 ;
        RECT 75.455 130.555 78.520 130.695 ;
        RECT 75.455 130.510 75.745 130.555 ;
        RECT 78.200 130.495 78.520 130.555 ;
        RECT 86.020 130.695 86.340 130.755 ;
        RECT 106.720 130.695 107.040 130.755 ;
        RECT 86.020 130.555 107.040 130.695 ;
        RECT 86.020 130.495 86.340 130.555 ;
        RECT 106.720 130.495 107.040 130.555 ;
        RECT 10.510 129.875 115.850 130.355 ;
        RECT 22.080 129.720 22.400 129.735 ;
        RECT 21.865 129.490 22.400 129.720 ;
        RECT 22.080 129.475 22.400 129.490 ;
        RECT 34.500 129.720 34.820 129.735 ;
        RECT 34.500 129.490 35.035 129.720 ;
        RECT 37.260 129.675 37.580 129.735 ;
        RECT 37.735 129.675 38.025 129.720 ;
        RECT 37.260 129.535 38.025 129.675 ;
        RECT 34.500 129.475 34.820 129.490 ;
        RECT 37.260 129.475 37.580 129.535 ;
        RECT 37.735 129.490 38.025 129.535 ;
        RECT 38.180 129.475 38.500 129.735 ;
        RECT 41.400 129.675 41.720 129.735 ;
        RECT 42.335 129.675 42.625 129.720 ;
        RECT 41.400 129.535 42.625 129.675 ;
        RECT 41.400 129.475 41.720 129.535 ;
        RECT 42.335 129.490 42.625 129.535 ;
        RECT 46.015 129.675 46.305 129.720 ;
        RECT 46.920 129.675 47.240 129.735 ;
        RECT 46.015 129.535 47.240 129.675 ;
        RECT 46.015 129.490 46.305 129.535 ;
        RECT 46.920 129.475 47.240 129.535 ;
        RECT 48.760 129.475 49.080 129.735 ;
        RECT 53.820 129.675 54.140 129.735 ;
        RECT 58.420 129.675 58.740 129.735 ;
        RECT 53.820 129.535 58.740 129.675 ;
        RECT 53.820 129.475 54.140 129.535 ;
        RECT 58.420 129.475 58.740 129.535 ;
        RECT 66.255 129.675 66.545 129.720 ;
        RECT 71.300 129.675 71.620 129.735 ;
        RECT 66.255 129.535 71.620 129.675 ;
        RECT 66.255 129.490 66.545 129.535 ;
        RECT 71.300 129.475 71.620 129.535 ;
        RECT 77.295 129.490 77.585 129.720 ;
        RECT 16.560 129.380 16.880 129.395 ;
        RECT 29.440 129.380 29.760 129.395 ;
        RECT 13.820 129.335 14.110 129.380 ;
        RECT 15.680 129.335 15.970 129.380 ;
        RECT 13.820 129.195 15.970 129.335 ;
        RECT 13.820 129.150 14.110 129.195 ;
        RECT 15.680 129.150 15.970 129.195 ;
        RECT 14.720 128.795 15.040 129.055 ;
        RECT 15.755 128.995 15.970 129.150 ;
        RECT 16.560 129.335 16.890 129.380 ;
        RECT 19.860 129.335 20.150 129.380 ;
        RECT 16.560 129.195 20.150 129.335 ;
        RECT 16.560 129.150 16.890 129.195 ;
        RECT 19.860 129.150 20.150 129.195 ;
        RECT 26.700 129.335 26.990 129.380 ;
        RECT 28.560 129.335 28.850 129.380 ;
        RECT 26.700 129.195 28.850 129.335 ;
        RECT 26.700 129.150 26.990 129.195 ;
        RECT 28.560 129.150 28.850 129.195 ;
        RECT 16.560 129.135 16.880 129.150 ;
        RECT 18.000 128.995 18.290 129.040 ;
        RECT 15.755 128.855 18.290 128.995 ;
        RECT 18.000 128.810 18.290 128.855 ;
        RECT 23.920 128.995 24.240 129.055 ;
        RECT 25.775 128.995 26.065 129.040 ;
        RECT 23.920 128.855 26.065 128.995 ;
        RECT 28.635 128.995 28.850 129.150 ;
        RECT 29.440 129.335 29.770 129.380 ;
        RECT 32.740 129.335 33.030 129.380 ;
        RECT 29.440 129.195 33.030 129.335 ;
        RECT 29.440 129.150 29.770 129.195 ;
        RECT 32.740 129.150 33.030 129.195 ;
        RECT 34.040 129.335 34.360 129.395 ;
        RECT 42.795 129.335 43.085 129.380 ;
        RECT 34.040 129.195 43.085 129.335 ;
        RECT 29.440 129.135 29.760 129.150 ;
        RECT 34.040 129.135 34.360 129.195 ;
        RECT 42.795 129.150 43.085 129.195 ;
        RECT 44.635 129.335 44.925 129.380 ;
        RECT 63.020 129.335 63.340 129.395 ;
        RECT 72.680 129.380 73.000 129.395 ;
        RECT 64.875 129.335 65.165 129.380 ;
        RECT 44.635 129.195 65.165 129.335 ;
        RECT 44.635 129.150 44.925 129.195 ;
        RECT 63.020 129.135 63.340 129.195 ;
        RECT 64.875 129.150 65.165 129.195 ;
        RECT 69.410 129.335 69.700 129.380 ;
        RECT 72.670 129.335 73.000 129.380 ;
        RECT 69.410 129.195 73.000 129.335 ;
        RECT 69.410 129.150 69.700 129.195 ;
        RECT 72.670 129.150 73.000 129.195 ;
        RECT 72.680 129.135 73.000 129.150 ;
        RECT 73.590 129.335 73.880 129.380 ;
        RECT 75.450 129.335 75.740 129.380 ;
        RECT 73.590 129.195 75.740 129.335 ;
        RECT 73.590 129.150 73.880 129.195 ;
        RECT 75.450 129.150 75.740 129.195 ;
        RECT 30.880 128.995 31.170 129.040 ;
        RECT 28.635 128.855 31.170 128.995 ;
        RECT 23.920 128.795 24.240 128.855 ;
        RECT 25.775 128.810 26.065 128.855 ;
        RECT 30.880 128.810 31.170 128.855 ;
        RECT 36.815 128.995 37.105 129.040 ;
        RECT 39.115 128.995 39.405 129.040 ;
        RECT 41.415 128.995 41.705 129.040 ;
        RECT 41.860 128.995 42.180 129.055 ;
        RECT 36.815 128.855 42.180 128.995 ;
        RECT 36.815 128.810 37.105 128.855 ;
        RECT 39.115 128.810 39.405 128.855 ;
        RECT 41.415 128.810 41.705 128.855 ;
        RECT 41.860 128.795 42.180 128.855 ;
        RECT 46.475 128.995 46.765 129.040 ;
        RECT 53.820 128.995 54.140 129.055 ;
        RECT 46.475 128.855 54.140 128.995 ;
        RECT 46.475 128.810 46.765 128.855 ;
        RECT 53.820 128.795 54.140 128.855 ;
        RECT 55.675 128.810 55.965 129.040 ;
        RECT 71.270 128.995 71.560 129.040 ;
        RECT 73.590 128.995 73.805 129.150 ;
        RECT 71.270 128.855 73.805 128.995 ;
        RECT 74.535 128.995 74.825 129.040 ;
        RECT 77.370 128.995 77.510 129.490 ;
        RECT 82.340 129.475 82.660 129.735 ;
        RECT 84.655 129.490 84.945 129.720 ;
        RECT 82.815 129.335 83.105 129.380 ;
        RECT 84.180 129.335 84.500 129.395 ;
        RECT 82.815 129.195 84.500 129.335 ;
        RECT 82.815 129.150 83.105 129.195 ;
        RECT 84.180 129.135 84.500 129.195 ;
        RECT 74.535 128.855 77.510 128.995 ;
        RECT 71.270 128.810 71.560 128.855 ;
        RECT 74.535 128.810 74.825 128.855 ;
        RECT 12.895 128.655 13.185 128.700 ;
        RECT 24.010 128.655 24.150 128.795 ;
        RECT 12.895 128.515 24.150 128.655 ;
        RECT 27.615 128.655 27.905 128.700 ;
        RECT 29.440 128.655 29.760 128.715 ;
        RECT 27.615 128.515 29.760 128.655 ;
        RECT 12.895 128.470 13.185 128.515 ;
        RECT 27.615 128.470 27.905 128.515 ;
        RECT 29.440 128.455 29.760 128.515 ;
        RECT 33.580 128.655 33.900 128.715 ;
        RECT 35.895 128.655 36.185 128.700 ;
        RECT 33.580 128.515 36.185 128.655 ;
        RECT 33.580 128.455 33.900 128.515 ;
        RECT 35.895 128.470 36.185 128.515 ;
        RECT 40.020 128.455 40.340 128.715 ;
        RECT 40.495 128.470 40.785 128.700 ;
        RECT 13.360 128.315 13.650 128.360 ;
        RECT 15.220 128.315 15.510 128.360 ;
        RECT 18.000 128.315 18.290 128.360 ;
        RECT 13.360 128.175 18.290 128.315 ;
        RECT 13.360 128.130 13.650 128.175 ;
        RECT 15.220 128.130 15.510 128.175 ;
        RECT 18.000 128.130 18.290 128.175 ;
        RECT 26.240 128.315 26.530 128.360 ;
        RECT 28.100 128.315 28.390 128.360 ;
        RECT 30.880 128.315 31.170 128.360 ;
        RECT 26.240 128.175 31.170 128.315 ;
        RECT 26.240 128.130 26.530 128.175 ;
        RECT 28.100 128.130 28.390 128.175 ;
        RECT 30.880 128.130 31.170 128.175 ;
        RECT 32.660 128.315 32.980 128.375 ;
        RECT 40.570 128.315 40.710 128.470 ;
        RECT 47.840 128.455 48.160 128.715 ;
        RECT 48.300 128.455 48.620 128.715 ;
        RECT 55.750 128.655 55.890 128.810 ;
        RECT 78.200 128.795 78.520 129.055 ;
        RECT 84.730 128.995 84.870 129.490 ;
        RECT 88.780 129.475 89.100 129.735 ;
        RECT 93.380 129.475 93.700 129.735 ;
        RECT 96.155 129.675 96.445 129.720 ;
        RECT 97.060 129.675 97.380 129.735 ;
        RECT 96.155 129.535 97.380 129.675 ;
        RECT 96.155 129.490 96.445 129.535 ;
        RECT 97.060 129.475 97.380 129.535 ;
        RECT 98.440 129.675 98.760 129.735 ;
        RECT 103.055 129.675 103.345 129.720 ;
        RECT 98.440 129.535 103.345 129.675 ;
        RECT 98.440 129.475 98.760 129.535 ;
        RECT 103.055 129.490 103.345 129.535 ;
        RECT 100.370 129.195 104.650 129.335 ;
        RECT 100.370 129.055 100.510 129.195 ;
        RECT 86.495 128.995 86.785 129.040 ;
        RECT 84.730 128.855 86.785 128.995 ;
        RECT 86.495 128.810 86.785 128.855 ;
        RECT 87.860 128.995 88.180 129.055 ;
        RECT 94.315 128.995 94.605 129.040 ;
        RECT 97.075 128.995 97.365 129.040 ;
        RECT 87.860 128.855 97.365 128.995 ;
        RECT 87.860 128.795 88.180 128.855 ;
        RECT 94.315 128.810 94.605 128.855 ;
        RECT 97.075 128.810 97.365 128.855 ;
        RECT 50.690 128.515 55.890 128.655 ;
        RECT 67.405 128.655 67.695 128.700 ;
        RECT 73.600 128.655 73.920 128.715 ;
        RECT 67.405 128.515 73.920 128.655 ;
        RECT 50.690 128.360 50.830 128.515 ;
        RECT 67.405 128.470 67.695 128.515 ;
        RECT 73.600 128.455 73.920 128.515 ;
        RECT 76.375 128.655 76.665 128.700 ;
        RECT 78.660 128.655 78.980 128.715 ;
        RECT 76.375 128.515 78.980 128.655 ;
        RECT 76.375 128.470 76.665 128.515 ;
        RECT 78.660 128.455 78.980 128.515 ;
        RECT 81.895 128.655 82.185 128.700 ;
        RECT 81.895 128.515 86.250 128.655 ;
        RECT 81.895 128.470 82.185 128.515 ;
        RECT 32.660 128.175 40.710 128.315 ;
        RECT 32.660 128.115 32.980 128.175 ;
        RECT 50.615 128.130 50.905 128.360 ;
        RECT 71.270 128.315 71.560 128.360 ;
        RECT 74.050 128.315 74.340 128.360 ;
        RECT 75.910 128.315 76.200 128.360 ;
        RECT 71.270 128.175 76.200 128.315 ;
        RECT 71.270 128.130 71.560 128.175 ;
        RECT 74.050 128.130 74.340 128.175 ;
        RECT 75.910 128.130 76.200 128.175 ;
        RECT 76.820 128.315 77.140 128.375 ;
        RECT 81.970 128.315 82.110 128.470 ;
        RECT 76.820 128.175 82.110 128.315 ;
        RECT 76.820 128.115 77.140 128.175 ;
        RECT 54.280 127.775 54.600 128.035 ;
        RECT 56.595 127.975 56.885 128.020 ;
        RECT 57.960 127.975 58.280 128.035 ;
        RECT 56.595 127.835 58.280 127.975 ;
        RECT 56.595 127.790 56.885 127.835 ;
        RECT 57.960 127.775 58.280 127.835 ;
        RECT 81.880 127.975 82.200 128.035 ;
        RECT 85.575 127.975 85.865 128.020 ;
        RECT 81.880 127.835 85.865 127.975 ;
        RECT 86.110 127.975 86.250 128.515 ;
        RECT 86.955 128.470 87.245 128.700 ;
        RECT 86.480 128.315 86.800 128.375 ;
        RECT 87.030 128.315 87.170 128.470 ;
        RECT 95.220 128.455 95.540 128.715 ;
        RECT 86.480 128.175 87.170 128.315 ;
        RECT 97.150 128.315 97.290 128.810 ;
        RECT 100.280 128.795 100.600 129.055 ;
        RECT 104.510 129.040 104.650 129.195 ;
        RECT 103.975 128.995 104.265 129.040 ;
        RECT 102.210 128.855 104.265 128.995 ;
        RECT 97.980 128.455 98.300 128.715 ;
        RECT 98.440 128.655 98.760 128.715 ;
        RECT 99.375 128.655 99.665 128.700 ;
        RECT 98.440 128.515 99.665 128.655 ;
        RECT 98.440 128.455 98.760 128.515 ;
        RECT 99.375 128.470 99.665 128.515 ;
        RECT 99.835 128.655 100.125 128.700 ;
        RECT 101.660 128.655 101.980 128.715 ;
        RECT 99.835 128.515 101.980 128.655 ;
        RECT 99.835 128.470 100.125 128.515 ;
        RECT 101.660 128.455 101.980 128.515 ;
        RECT 102.210 128.315 102.350 128.855 ;
        RECT 103.975 128.810 104.265 128.855 ;
        RECT 104.435 128.810 104.725 129.040 ;
        RECT 106.720 128.795 107.040 129.055 ;
        RECT 108.575 128.810 108.865 129.040 ;
        RECT 103.500 128.655 103.820 128.715 ;
        RECT 108.650 128.655 108.790 128.810 ;
        RECT 103.500 128.515 108.790 128.655 ;
        RECT 103.500 128.455 103.820 128.515 ;
        RECT 97.150 128.175 102.350 128.315 ;
        RECT 86.480 128.115 86.800 128.175 ;
        RECT 94.760 127.975 95.080 128.035 ;
        RECT 86.110 127.835 95.080 127.975 ;
        RECT 81.880 127.775 82.200 127.835 ;
        RECT 85.575 127.790 85.865 127.835 ;
        RECT 94.760 127.775 95.080 127.835 ;
        RECT 102.135 127.975 102.425 128.020 ;
        RECT 104.880 127.975 105.200 128.035 ;
        RECT 102.135 127.835 105.200 127.975 ;
        RECT 102.135 127.790 102.425 127.835 ;
        RECT 104.880 127.775 105.200 127.835 ;
        RECT 107.180 127.775 107.500 128.035 ;
        RECT 109.480 127.775 109.800 128.035 ;
        RECT 10.510 127.155 115.850 127.635 ;
        RECT 15.195 126.955 15.485 127.000 ;
        RECT 16.560 126.955 16.880 127.015 ;
        RECT 15.195 126.815 16.880 126.955 ;
        RECT 15.195 126.770 15.485 126.815 ;
        RECT 16.560 126.755 16.880 126.815 ;
        RECT 28.535 126.955 28.825 127.000 ;
        RECT 28.980 126.955 29.300 127.015 ;
        RECT 28.535 126.815 29.300 126.955 ;
        RECT 28.535 126.770 28.825 126.815 ;
        RECT 28.980 126.755 29.300 126.815 ;
        RECT 29.440 126.755 29.760 127.015 ;
        RECT 32.675 126.955 32.965 127.000 ;
        RECT 33.120 126.955 33.440 127.015 ;
        RECT 32.675 126.815 33.440 126.955 ;
        RECT 32.675 126.770 32.965 126.815 ;
        RECT 33.120 126.755 33.440 126.815 ;
        RECT 42.320 126.755 42.640 127.015 ;
        RECT 48.300 126.955 48.620 127.015 ;
        RECT 50.845 126.955 51.135 127.000 ;
        RECT 48.300 126.815 51.135 126.955 ;
        RECT 48.300 126.755 48.620 126.815 ;
        RECT 50.845 126.770 51.135 126.815 ;
        RECT 72.680 126.955 73.000 127.015 ;
        RECT 74.995 126.955 75.285 127.000 ;
        RECT 72.680 126.815 75.285 126.955 ;
        RECT 72.680 126.755 73.000 126.815 ;
        RECT 74.995 126.770 75.285 126.815 ;
        RECT 84.180 126.955 84.500 127.015 ;
        RECT 89.025 126.955 89.315 127.000 ;
        RECT 97.980 126.955 98.300 127.015 ;
        RECT 84.180 126.815 98.300 126.955 ;
        RECT 84.180 126.755 84.500 126.815 ;
        RECT 89.025 126.770 89.315 126.815 ;
        RECT 97.980 126.755 98.300 126.815 ;
        RECT 103.500 126.755 103.820 127.015 ;
        RECT 14.720 126.615 15.040 126.675 ;
        RECT 16.115 126.615 16.405 126.660 ;
        RECT 54.710 126.615 55.000 126.660 ;
        RECT 57.490 126.615 57.780 126.660 ;
        RECT 59.350 126.615 59.640 126.660 ;
        RECT 14.720 126.475 16.405 126.615 ;
        RECT 14.720 126.415 15.040 126.475 ;
        RECT 16.115 126.430 16.405 126.475 ;
        RECT 16.650 126.475 24.610 126.615 ;
        RECT 14.260 125.935 14.580 125.995 ;
        RECT 14.735 125.935 15.025 125.980 ;
        RECT 16.650 125.935 16.790 126.475 ;
        RECT 18.860 126.275 19.180 126.335 ;
        RECT 20.240 126.275 20.560 126.335 ;
        RECT 18.860 126.135 20.560 126.275 ;
        RECT 18.860 126.075 19.180 126.135 ;
        RECT 20.240 126.075 20.560 126.135 ;
        RECT 24.470 125.995 24.610 126.475 ;
        RECT 54.710 126.475 59.640 126.615 ;
        RECT 54.710 126.430 55.000 126.475 ;
        RECT 57.490 126.430 57.780 126.475 ;
        RECT 59.350 126.430 59.640 126.475 ;
        RECT 80.520 126.615 80.810 126.660 ;
        RECT 82.380 126.615 82.670 126.660 ;
        RECT 85.160 126.615 85.450 126.660 ;
        RECT 80.520 126.475 85.450 126.615 ;
        RECT 98.070 126.615 98.210 126.755 ;
        RECT 108.070 126.615 108.360 126.660 ;
        RECT 110.850 126.615 111.140 126.660 ;
        RECT 112.710 126.615 113.000 126.660 ;
        RECT 98.070 126.475 100.970 126.615 ;
        RECT 80.520 126.430 80.810 126.475 ;
        RECT 82.380 126.430 82.670 126.475 ;
        RECT 85.160 126.430 85.450 126.475 ;
        RECT 28.520 126.275 28.840 126.335 ;
        RECT 30.835 126.275 31.125 126.320 ;
        RECT 28.520 126.135 32.430 126.275 ;
        RECT 28.520 126.075 28.840 126.135 ;
        RECT 30.835 126.090 31.125 126.135 ;
        RECT 14.260 125.795 16.790 125.935 ;
        RECT 14.260 125.735 14.580 125.795 ;
        RECT 14.735 125.750 15.025 125.795 ;
        RECT 17.020 125.735 17.340 125.995 ;
        RECT 19.795 125.935 20.085 125.980 ;
        RECT 22.080 125.935 22.400 125.995 ;
        RECT 19.795 125.795 22.400 125.935 ;
        RECT 19.795 125.750 20.085 125.795 ;
        RECT 22.080 125.735 22.400 125.795 ;
        RECT 22.555 125.935 22.845 125.980 ;
        RECT 23.000 125.935 23.320 125.995 ;
        RECT 22.555 125.795 23.320 125.935 ;
        RECT 22.555 125.750 22.845 125.795 ;
        RECT 23.000 125.735 23.320 125.795 ;
        RECT 24.380 125.935 24.700 125.995 ;
        RECT 26.695 125.935 26.985 125.980 ;
        RECT 28.075 125.935 28.365 125.980 ;
        RECT 24.380 125.795 28.365 125.935 ;
        RECT 24.380 125.735 24.700 125.795 ;
        RECT 26.695 125.750 26.985 125.795 ;
        RECT 28.075 125.750 28.365 125.795 ;
        RECT 30.360 125.735 30.680 125.995 ;
        RECT 31.755 125.935 32.045 125.980 ;
        RECT 30.910 125.795 32.045 125.935 ;
        RECT 32.290 125.935 32.430 126.135 ;
        RECT 34.040 126.075 34.360 126.335 ;
        RECT 57.960 126.075 58.280 126.335 ;
        RECT 59.815 126.275 60.105 126.320 ;
        RECT 63.480 126.275 63.800 126.335 ;
        RECT 59.815 126.135 63.800 126.275 ;
        RECT 59.815 126.090 60.105 126.135 ;
        RECT 63.480 126.075 63.800 126.135 ;
        RECT 69.475 126.275 69.765 126.320 ;
        RECT 71.300 126.275 71.620 126.335 ;
        RECT 76.820 126.275 77.140 126.335 ;
        RECT 69.475 126.135 77.140 126.275 ;
        RECT 69.475 126.090 69.765 126.135 ;
        RECT 71.300 126.075 71.620 126.135 ;
        RECT 76.820 126.075 77.140 126.135 ;
        RECT 78.660 126.275 78.980 126.335 ;
        RECT 80.055 126.275 80.345 126.320 ;
        RECT 78.660 126.135 80.345 126.275 ;
        RECT 78.660 126.075 78.980 126.135 ;
        RECT 34.975 125.935 35.265 125.980 ;
        RECT 32.290 125.795 35.265 125.935 ;
        RECT 30.910 125.655 31.050 125.795 ;
        RECT 31.755 125.750 32.045 125.795 ;
        RECT 34.975 125.750 35.265 125.795 ;
        RECT 40.480 125.735 40.800 125.995 ;
        RECT 41.415 125.935 41.705 125.980 ;
        RECT 41.860 125.935 42.180 125.995 ;
        RECT 41.415 125.795 42.180 125.935 ;
        RECT 41.415 125.750 41.705 125.795 ;
        RECT 41.860 125.735 42.180 125.795 ;
        RECT 43.700 125.735 44.020 125.995 ;
        RECT 54.710 125.935 55.000 125.980 ;
        RECT 54.710 125.795 57.245 125.935 ;
        RECT 54.710 125.750 55.000 125.795 ;
        RECT 19.320 125.395 19.640 125.655 ;
        RECT 30.820 125.395 31.140 125.655 ;
        RECT 52.850 125.595 53.140 125.640 ;
        RECT 54.280 125.595 54.600 125.655 ;
        RECT 57.030 125.640 57.245 125.795 ;
        RECT 75.440 125.735 75.760 125.995 ;
        RECT 79.670 125.980 79.810 126.135 ;
        RECT 80.055 126.090 80.345 126.135 ;
        RECT 81.880 126.075 82.200 126.335 ;
        RECT 94.760 126.075 95.080 126.335 ;
        RECT 95.235 126.275 95.525 126.320 ;
        RECT 97.980 126.275 98.300 126.335 ;
        RECT 95.235 126.135 98.300 126.275 ;
        RECT 95.235 126.090 95.525 126.135 ;
        RECT 97.980 126.075 98.300 126.135 ;
        RECT 98.440 126.275 98.760 126.335 ;
        RECT 100.295 126.275 100.585 126.320 ;
        RECT 98.440 126.135 100.585 126.275 ;
        RECT 98.440 126.075 98.760 126.135 ;
        RECT 100.295 126.090 100.585 126.135 ;
        RECT 79.595 125.935 79.885 125.980 ;
        RECT 85.160 125.935 85.450 125.980 ;
        RECT 79.485 125.795 79.885 125.935 ;
        RECT 79.595 125.750 79.885 125.795 ;
        RECT 82.915 125.795 85.450 125.935 ;
        RECT 56.110 125.595 56.400 125.640 ;
        RECT 52.850 125.455 56.400 125.595 ;
        RECT 52.850 125.410 53.140 125.455 ;
        RECT 54.280 125.395 54.600 125.455 ;
        RECT 56.110 125.410 56.400 125.455 ;
        RECT 57.030 125.595 57.320 125.640 ;
        RECT 58.890 125.595 59.180 125.640 ;
        RECT 57.030 125.455 59.180 125.595 ;
        RECT 57.030 125.410 57.320 125.455 ;
        RECT 58.890 125.410 59.180 125.455 ;
        RECT 69.935 125.595 70.225 125.640 ;
        RECT 71.760 125.595 72.080 125.655 ;
        RECT 82.915 125.640 83.130 125.795 ;
        RECT 85.160 125.750 85.450 125.795 ;
        RECT 86.020 125.935 86.340 125.995 ;
        RECT 92.000 125.935 92.320 125.995 ;
        RECT 92.475 125.935 92.765 125.980 ;
        RECT 86.020 125.795 92.765 125.935 ;
        RECT 94.850 125.935 94.990 126.075 ;
        RECT 98.530 125.935 98.670 126.075 ;
        RECT 94.850 125.795 98.670 125.935 ;
        RECT 100.830 125.935 100.970 126.475 ;
        RECT 108.070 126.475 113.000 126.615 ;
        RECT 108.070 126.430 108.360 126.475 ;
        RECT 110.850 126.430 111.140 126.475 ;
        RECT 112.710 126.430 113.000 126.475 ;
        RECT 109.480 126.275 109.800 126.335 ;
        RECT 111.335 126.275 111.625 126.320 ;
        RECT 109.480 126.135 111.625 126.275 ;
        RECT 109.480 126.075 109.800 126.135 ;
        RECT 111.335 126.090 111.625 126.135 ;
        RECT 113.160 126.275 113.480 126.335 ;
        RECT 114.080 126.275 114.400 126.335 ;
        RECT 113.160 126.135 114.400 126.275 ;
        RECT 113.160 126.075 113.480 126.135 ;
        RECT 114.080 126.075 114.400 126.135 ;
        RECT 101.215 125.935 101.505 125.980 ;
        RECT 100.830 125.795 101.505 125.935 ;
        RECT 86.020 125.735 86.340 125.795 ;
        RECT 92.000 125.735 92.320 125.795 ;
        RECT 92.475 125.750 92.765 125.795 ;
        RECT 101.215 125.750 101.505 125.795 ;
        RECT 101.660 125.935 101.980 125.995 ;
        RECT 104.205 125.935 104.495 125.980 ;
        RECT 101.660 125.795 104.495 125.935 ;
        RECT 101.660 125.735 101.980 125.795 ;
        RECT 104.205 125.750 104.495 125.795 ;
        RECT 108.070 125.935 108.360 125.980 ;
        RECT 108.070 125.795 110.605 125.935 ;
        RECT 108.070 125.750 108.360 125.795 ;
        RECT 69.935 125.455 72.080 125.595 ;
        RECT 69.935 125.410 70.225 125.455 ;
        RECT 71.760 125.395 72.080 125.455 ;
        RECT 80.980 125.595 81.270 125.640 ;
        RECT 82.840 125.595 83.130 125.640 ;
        RECT 80.980 125.455 83.130 125.595 ;
        RECT 80.980 125.410 81.270 125.455 ;
        RECT 82.840 125.410 83.130 125.455 ;
        RECT 83.760 125.595 84.050 125.640 ;
        RECT 87.020 125.595 87.310 125.640 ;
        RECT 91.540 125.595 91.860 125.655 ;
        RECT 95.220 125.595 95.540 125.655 ;
        RECT 95.695 125.595 95.985 125.640 ;
        RECT 83.760 125.455 91.860 125.595 ;
        RECT 83.760 125.410 84.050 125.455 ;
        RECT 87.020 125.410 87.310 125.455 ;
        RECT 91.540 125.395 91.860 125.455 ;
        RECT 92.550 125.455 95.985 125.595 ;
        RECT 17.480 125.055 17.800 125.315 ;
        RECT 18.860 125.255 19.180 125.315 ;
        RECT 21.635 125.255 21.925 125.300 ;
        RECT 18.860 125.115 21.925 125.255 ;
        RECT 18.860 125.055 19.180 125.115 ;
        RECT 21.635 125.070 21.925 125.115 ;
        RECT 27.140 125.055 27.460 125.315 ;
        RECT 33.580 125.255 33.900 125.315 ;
        RECT 34.515 125.255 34.805 125.300 ;
        RECT 33.580 125.115 34.805 125.255 ;
        RECT 33.580 125.055 33.900 125.115 ;
        RECT 34.515 125.070 34.805 125.115 ;
        RECT 36.815 125.255 37.105 125.300 ;
        RECT 37.720 125.255 38.040 125.315 ;
        RECT 36.815 125.115 38.040 125.255 ;
        RECT 36.815 125.070 37.105 125.115 ;
        RECT 37.720 125.055 38.040 125.115 ;
        RECT 44.160 125.055 44.480 125.315 ;
        RECT 47.840 125.255 48.160 125.315 ;
        RECT 54.740 125.255 55.060 125.315 ;
        RECT 47.840 125.115 55.060 125.255 ;
        RECT 47.840 125.055 48.160 125.115 ;
        RECT 54.740 125.055 55.060 125.115 ;
        RECT 70.380 125.055 70.700 125.315 ;
        RECT 72.235 125.255 72.525 125.300 ;
        RECT 76.360 125.255 76.680 125.315 ;
        RECT 72.235 125.115 76.680 125.255 ;
        RECT 72.235 125.070 72.525 125.115 ;
        RECT 76.360 125.055 76.680 125.115 ;
        RECT 88.320 125.255 88.640 125.315 ;
        RECT 92.550 125.255 92.690 125.455 ;
        RECT 95.220 125.395 95.540 125.455 ;
        RECT 95.695 125.410 95.985 125.455 ;
        RECT 106.210 125.595 106.500 125.640 ;
        RECT 107.180 125.595 107.500 125.655 ;
        RECT 110.390 125.640 110.605 125.795 ;
        RECT 109.470 125.595 109.760 125.640 ;
        RECT 106.210 125.455 109.760 125.595 ;
        RECT 106.210 125.410 106.500 125.455 ;
        RECT 107.180 125.395 107.500 125.455 ;
        RECT 109.470 125.410 109.760 125.455 ;
        RECT 110.390 125.595 110.680 125.640 ;
        RECT 112.250 125.595 112.540 125.640 ;
        RECT 110.390 125.455 112.540 125.595 ;
        RECT 110.390 125.410 110.680 125.455 ;
        RECT 112.250 125.410 112.540 125.455 ;
        RECT 88.320 125.115 92.690 125.255 ;
        RECT 92.935 125.255 93.225 125.300 ;
        RECT 93.840 125.255 94.160 125.315 ;
        RECT 92.935 125.115 94.160 125.255 ;
        RECT 88.320 125.055 88.640 125.115 ;
        RECT 92.935 125.070 93.225 125.115 ;
        RECT 93.840 125.055 94.160 125.115 ;
        RECT 97.060 125.255 97.380 125.315 ;
        RECT 97.535 125.255 97.825 125.300 ;
        RECT 97.060 125.115 97.825 125.255 ;
        RECT 97.060 125.055 97.380 125.115 ;
        RECT 97.535 125.070 97.825 125.115 ;
        RECT 10.510 124.435 115.850 124.915 ;
        RECT 18.400 124.235 18.720 124.295 ;
        RECT 23.920 124.235 24.240 124.295 ;
        RECT 18.400 124.095 24.240 124.235 ;
        RECT 18.400 124.035 18.720 124.095 ;
        RECT 23.920 124.035 24.240 124.095 ;
        RECT 48.300 124.235 48.620 124.295 ;
        RECT 55.675 124.235 55.965 124.280 ;
        RECT 66.025 124.235 66.315 124.280 ;
        RECT 70.380 124.235 70.700 124.295 ;
        RECT 48.300 124.095 55.965 124.235 ;
        RECT 48.300 124.035 48.620 124.095 ;
        RECT 55.675 124.050 55.965 124.095 ;
        RECT 56.210 124.095 60.030 124.235 ;
        RECT 33.070 123.895 33.360 123.940 ;
        RECT 34.040 123.895 34.360 123.955 ;
        RECT 36.330 123.895 36.620 123.940 ;
        RECT 33.070 123.755 36.620 123.895 ;
        RECT 33.070 123.710 33.360 123.755 ;
        RECT 34.040 123.695 34.360 123.755 ;
        RECT 36.330 123.710 36.620 123.755 ;
        RECT 37.250 123.895 37.540 123.940 ;
        RECT 39.110 123.895 39.400 123.940 ;
        RECT 37.250 123.755 39.400 123.895 ;
        RECT 37.250 123.710 37.540 123.755 ;
        RECT 39.110 123.710 39.400 123.755 ;
        RECT 42.730 123.895 43.020 123.940 ;
        RECT 44.160 123.895 44.480 123.955 ;
        RECT 45.990 123.895 46.280 123.940 ;
        RECT 42.730 123.755 46.280 123.895 ;
        RECT 42.730 123.710 43.020 123.755 ;
        RECT 14.260 123.355 14.580 123.615 ;
        RECT 15.655 123.555 15.945 123.600 ;
        RECT 17.480 123.555 17.800 123.615 ;
        RECT 15.655 123.415 17.800 123.555 ;
        RECT 15.655 123.370 15.945 123.415 ;
        RECT 17.480 123.355 17.800 123.415 ;
        RECT 24.840 123.355 25.160 123.615 ;
        RECT 26.680 123.555 27.000 123.615 ;
        RECT 28.520 123.555 28.840 123.615 ;
        RECT 26.680 123.415 28.840 123.555 ;
        RECT 26.680 123.355 27.000 123.415 ;
        RECT 28.520 123.355 28.840 123.415 ;
        RECT 31.065 123.555 31.355 123.600 ;
        RECT 33.580 123.555 33.900 123.615 ;
        RECT 31.065 123.415 33.900 123.555 ;
        RECT 31.065 123.370 31.355 123.415 ;
        RECT 33.580 123.355 33.900 123.415 ;
        RECT 34.930 123.555 35.220 123.600 ;
        RECT 37.250 123.555 37.465 123.710 ;
        RECT 44.160 123.695 44.480 123.755 ;
        RECT 45.990 123.710 46.280 123.755 ;
        RECT 46.910 123.895 47.200 123.940 ;
        RECT 48.770 123.895 49.060 123.940 ;
        RECT 46.910 123.755 49.060 123.895 ;
        RECT 46.910 123.710 47.200 123.755 ;
        RECT 48.770 123.710 49.060 123.755 ;
        RECT 51.980 123.895 52.300 123.955 ;
        RECT 56.210 123.940 56.350 124.095 ;
        RECT 56.135 123.895 56.425 123.940 ;
        RECT 51.980 123.755 56.425 123.895 ;
        RECT 34.930 123.415 37.465 123.555 ;
        RECT 40.035 123.555 40.325 123.600 ;
        RECT 43.240 123.555 43.560 123.615 ;
        RECT 40.035 123.415 43.560 123.555 ;
        RECT 34.930 123.370 35.220 123.415 ;
        RECT 40.035 123.370 40.325 123.415 ;
        RECT 43.240 123.355 43.560 123.415 ;
        RECT 44.590 123.555 44.880 123.600 ;
        RECT 46.910 123.555 47.125 123.710 ;
        RECT 51.980 123.695 52.300 123.755 ;
        RECT 56.135 123.710 56.425 123.755 ;
        RECT 56.580 123.895 56.900 123.955 ;
        RECT 59.355 123.895 59.645 123.940 ;
        RECT 56.580 123.755 59.645 123.895 ;
        RECT 56.580 123.695 56.900 123.755 ;
        RECT 59.355 123.710 59.645 123.755 ;
        RECT 59.890 123.615 60.030 124.095 ;
        RECT 66.025 124.095 70.700 124.235 ;
        RECT 66.025 124.050 66.315 124.095 ;
        RECT 70.380 124.035 70.700 124.095 ;
        RECT 78.660 124.035 78.980 124.295 ;
        RECT 91.540 124.035 91.860 124.295 ;
        RECT 104.880 124.235 105.200 124.295 ;
        RECT 104.880 124.095 114.310 124.235 ;
        RECT 104.880 124.035 105.200 124.095 ;
        RECT 68.030 123.895 68.320 123.940 ;
        RECT 69.000 123.895 69.320 123.955 ;
        RECT 71.290 123.895 71.580 123.940 ;
        RECT 68.030 123.755 71.580 123.895 ;
        RECT 68.030 123.710 68.320 123.755 ;
        RECT 69.000 123.695 69.320 123.755 ;
        RECT 71.290 123.710 71.580 123.755 ;
        RECT 72.210 123.895 72.500 123.940 ;
        RECT 74.070 123.895 74.360 123.940 ;
        RECT 78.750 123.895 78.890 124.035 ;
        RECT 72.210 123.755 74.360 123.895 ;
        RECT 72.210 123.710 72.500 123.755 ;
        RECT 74.070 123.710 74.360 123.755 ;
        RECT 75.070 123.755 78.890 123.895 ;
        RECT 86.020 123.895 86.340 123.955 ;
        RECT 93.395 123.895 93.685 123.940 ;
        RECT 86.020 123.755 93.685 123.895 ;
        RECT 44.590 123.415 47.125 123.555 ;
        RECT 47.855 123.555 48.145 123.600 ;
        RECT 49.220 123.555 49.540 123.615 ;
        RECT 47.855 123.415 49.540 123.555 ;
        RECT 44.590 123.370 44.880 123.415 ;
        RECT 47.855 123.370 48.145 123.415 ;
        RECT 49.220 123.355 49.540 123.415 ;
        RECT 51.535 123.555 51.825 123.600 ;
        RECT 51.535 123.415 54.050 123.555 ;
        RECT 51.535 123.370 51.825 123.415 ;
        RECT 20.240 123.215 20.560 123.275 ;
        RECT 26.220 123.215 26.540 123.275 ;
        RECT 27.155 123.215 27.445 123.260 ;
        RECT 20.240 123.075 27.445 123.215 ;
        RECT 20.240 123.015 20.560 123.075 ;
        RECT 26.220 123.015 26.540 123.075 ;
        RECT 27.155 123.030 27.445 123.075 ;
        RECT 28.060 123.015 28.380 123.275 ;
        RECT 38.180 123.015 38.500 123.275 ;
        RECT 43.330 123.215 43.470 123.355 ;
        RECT 48.300 123.215 48.620 123.275 ;
        RECT 49.695 123.215 49.985 123.260 ;
        RECT 43.330 123.075 49.985 123.215 ;
        RECT 48.300 123.015 48.620 123.075 ;
        RECT 49.695 123.030 49.985 123.075 ;
        RECT 13.815 122.875 14.105 122.920 ;
        RECT 17.020 122.875 17.340 122.935 ;
        RECT 53.910 122.920 54.050 123.415 ;
        RECT 59.800 123.355 60.120 123.615 ;
        RECT 69.890 123.555 70.180 123.600 ;
        RECT 72.210 123.555 72.425 123.710 ;
        RECT 75.070 123.600 75.210 123.755 ;
        RECT 86.020 123.695 86.340 123.755 ;
        RECT 93.395 123.710 93.685 123.755 ;
        RECT 105.750 123.895 106.040 123.940 ;
        RECT 106.720 123.895 107.040 123.955 ;
        RECT 109.010 123.895 109.300 123.940 ;
        RECT 105.750 123.755 109.300 123.895 ;
        RECT 105.750 123.710 106.040 123.755 ;
        RECT 106.720 123.695 107.040 123.755 ;
        RECT 109.010 123.710 109.300 123.755 ;
        RECT 109.930 123.895 110.220 123.940 ;
        RECT 111.790 123.895 112.080 123.940 ;
        RECT 109.930 123.755 112.080 123.895 ;
        RECT 109.930 123.710 110.220 123.755 ;
        RECT 111.790 123.710 112.080 123.755 ;
        RECT 69.890 123.415 72.425 123.555 ;
        RECT 69.890 123.370 70.180 123.415 ;
        RECT 74.995 123.370 75.285 123.600 ;
        RECT 76.360 123.355 76.680 123.615 ;
        RECT 83.260 123.555 83.580 123.615 ;
        RECT 86.480 123.555 86.800 123.615 ;
        RECT 88.795 123.555 89.085 123.600 ;
        RECT 83.260 123.415 89.085 123.555 ;
        RECT 83.260 123.355 83.580 123.415 ;
        RECT 86.480 123.355 86.800 123.415 ;
        RECT 88.795 123.370 89.085 123.415 ;
        RECT 92.000 123.355 92.320 123.615 ;
        RECT 107.610 123.555 107.900 123.600 ;
        RECT 109.930 123.555 110.145 123.710 ;
        RECT 107.610 123.415 110.145 123.555 ;
        RECT 112.715 123.555 113.005 123.600 ;
        RECT 113.160 123.555 113.480 123.615 ;
        RECT 114.170 123.600 114.310 124.095 ;
        RECT 112.715 123.415 113.480 123.555 ;
        RECT 107.610 123.370 107.900 123.415 ;
        RECT 112.715 123.370 113.005 123.415 ;
        RECT 113.160 123.355 113.480 123.415 ;
        RECT 114.095 123.370 114.385 123.600 ;
        RECT 54.740 123.215 55.060 123.275 ;
        RECT 57.055 123.215 57.345 123.260 ;
        RECT 58.435 123.215 58.725 123.260 ;
        RECT 54.740 123.075 58.725 123.215 ;
        RECT 54.740 123.015 55.060 123.075 ;
        RECT 57.055 123.030 57.345 123.075 ;
        RECT 58.435 123.030 58.725 123.075 ;
        RECT 73.155 123.215 73.445 123.260 ;
        RECT 73.155 123.075 75.670 123.215 ;
        RECT 73.155 123.030 73.445 123.075 ;
        RECT 75.530 122.920 75.670 123.075 ;
        RECT 87.875 123.030 88.165 123.260 ;
        RECT 13.815 122.735 17.340 122.875 ;
        RECT 13.815 122.690 14.105 122.735 ;
        RECT 17.020 122.675 17.340 122.735 ;
        RECT 34.930 122.875 35.220 122.920 ;
        RECT 37.710 122.875 38.000 122.920 ;
        RECT 39.570 122.875 39.860 122.920 ;
        RECT 34.930 122.735 39.860 122.875 ;
        RECT 34.930 122.690 35.220 122.735 ;
        RECT 37.710 122.690 38.000 122.735 ;
        RECT 39.570 122.690 39.860 122.735 ;
        RECT 44.590 122.875 44.880 122.920 ;
        RECT 47.370 122.875 47.660 122.920 ;
        RECT 49.230 122.875 49.520 122.920 ;
        RECT 44.590 122.735 49.520 122.875 ;
        RECT 44.590 122.690 44.880 122.735 ;
        RECT 47.370 122.690 47.660 122.735 ;
        RECT 49.230 122.690 49.520 122.735 ;
        RECT 53.835 122.690 54.125 122.920 ;
        RECT 69.890 122.875 70.180 122.920 ;
        RECT 72.670 122.875 72.960 122.920 ;
        RECT 74.530 122.875 74.820 122.920 ;
        RECT 69.890 122.735 74.820 122.875 ;
        RECT 69.890 122.690 70.180 122.735 ;
        RECT 72.670 122.690 72.960 122.735 ;
        RECT 74.530 122.690 74.820 122.735 ;
        RECT 75.455 122.690 75.745 122.920 ;
        RECT 87.950 122.875 88.090 123.030 ;
        RECT 88.320 123.015 88.640 123.275 ;
        RECT 110.875 123.215 111.165 123.260 ;
        RECT 110.875 123.075 113.390 123.215 ;
        RECT 110.875 123.030 111.165 123.075 ;
        RECT 98.440 122.875 98.760 122.935 ;
        RECT 113.250 122.920 113.390 123.075 ;
        RECT 87.950 122.735 98.760 122.875 ;
        RECT 98.440 122.675 98.760 122.735 ;
        RECT 107.610 122.875 107.900 122.920 ;
        RECT 110.390 122.875 110.680 122.920 ;
        RECT 112.250 122.875 112.540 122.920 ;
        RECT 107.610 122.735 112.540 122.875 ;
        RECT 107.610 122.690 107.900 122.735 ;
        RECT 110.390 122.690 110.680 122.735 ;
        RECT 112.250 122.690 112.540 122.735 ;
        RECT 113.175 122.690 113.465 122.920 ;
        RECT 14.735 122.535 15.025 122.580 ;
        RECT 15.180 122.535 15.500 122.595 ;
        RECT 14.735 122.395 15.500 122.535 ;
        RECT 14.735 122.350 15.025 122.395 ;
        RECT 15.180 122.335 15.500 122.395 ;
        RECT 30.360 122.335 30.680 122.595 ;
        RECT 40.020 122.535 40.340 122.595 ;
        RECT 40.725 122.535 41.015 122.580 ;
        RECT 40.020 122.395 41.015 122.535 ;
        RECT 40.020 122.335 40.340 122.395 ;
        RECT 40.725 122.350 41.015 122.395 ;
        RECT 52.455 122.535 52.745 122.580 ;
        RECT 55.200 122.535 55.520 122.595 ;
        RECT 52.455 122.395 55.520 122.535 ;
        RECT 52.455 122.350 52.745 122.395 ;
        RECT 55.200 122.335 55.520 122.395 ;
        RECT 61.655 122.535 61.945 122.580 ;
        RECT 65.320 122.535 65.640 122.595 ;
        RECT 61.655 122.395 65.640 122.535 ;
        RECT 61.655 122.350 61.945 122.395 ;
        RECT 65.320 122.335 65.640 122.395 ;
        RECT 89.700 122.535 90.020 122.595 ;
        RECT 90.635 122.535 90.925 122.580 ;
        RECT 89.700 122.395 90.925 122.535 ;
        RECT 89.700 122.335 90.020 122.395 ;
        RECT 90.635 122.350 90.925 122.395 ;
        RECT 99.360 122.535 99.680 122.595 ;
        RECT 99.835 122.535 100.125 122.580 ;
        RECT 99.360 122.395 100.125 122.535 ;
        RECT 99.360 122.335 99.680 122.395 ;
        RECT 99.835 122.350 100.125 122.395 ;
        RECT 100.280 122.535 100.600 122.595 ;
        RECT 103.745 122.535 104.035 122.580 ;
        RECT 100.280 122.395 104.035 122.535 ;
        RECT 100.280 122.335 100.600 122.395 ;
        RECT 103.745 122.350 104.035 122.395 ;
        RECT 10.510 121.715 115.850 122.195 ;
        RECT 23.000 121.315 23.320 121.575 ;
        RECT 28.060 121.560 28.380 121.575 ;
        RECT 27.845 121.330 28.380 121.560 ;
        RECT 32.660 121.515 32.980 121.575 ;
        RECT 28.060 121.315 28.380 121.330 ;
        RECT 28.610 121.375 32.980 121.515 ;
        RECT 13.820 121.175 14.110 121.220 ;
        RECT 15.680 121.175 15.970 121.220 ;
        RECT 18.460 121.175 18.750 121.220 ;
        RECT 13.820 121.035 18.750 121.175 ;
        RECT 13.820 120.990 14.110 121.035 ;
        RECT 15.680 120.990 15.970 121.035 ;
        RECT 18.460 120.990 18.750 121.035 ;
        RECT 19.320 121.175 19.640 121.235 ;
        RECT 22.325 121.175 22.615 121.220 ;
        RECT 28.610 121.175 28.750 121.375 ;
        RECT 32.660 121.315 32.980 121.375 ;
        RECT 52.440 121.515 52.760 121.575 ;
        RECT 54.525 121.515 54.815 121.560 ;
        RECT 56.580 121.515 56.900 121.575 ;
        RECT 52.440 121.375 56.900 121.515 ;
        RECT 52.440 121.315 52.760 121.375 ;
        RECT 54.525 121.330 54.815 121.375 ;
        RECT 56.580 121.315 56.900 121.375 ;
        RECT 69.000 121.315 69.320 121.575 ;
        RECT 88.320 121.515 88.640 121.575 ;
        RECT 90.405 121.515 90.695 121.560 ;
        RECT 88.320 121.375 90.695 121.515 ;
        RECT 88.320 121.315 88.640 121.375 ;
        RECT 90.405 121.330 90.695 121.375 ;
        RECT 19.320 121.035 28.750 121.175 ;
        RECT 31.710 121.175 32.000 121.220 ;
        RECT 34.490 121.175 34.780 121.220 ;
        RECT 36.350 121.175 36.640 121.220 ;
        RECT 31.710 121.035 36.640 121.175 ;
        RECT 19.320 120.975 19.640 121.035 ;
        RECT 22.325 120.990 22.615 121.035 ;
        RECT 15.180 120.635 15.500 120.895 ;
        RECT 25.390 120.880 25.530 121.035 ;
        RECT 31.710 120.990 32.000 121.035 ;
        RECT 34.490 120.990 34.780 121.035 ;
        RECT 36.350 120.990 36.640 121.035 ;
        RECT 58.390 121.175 58.680 121.220 ;
        RECT 61.170 121.175 61.460 121.220 ;
        RECT 63.030 121.175 63.320 121.220 ;
        RECT 58.390 121.035 63.320 121.175 ;
        RECT 58.390 120.990 58.680 121.035 ;
        RECT 61.170 120.990 61.460 121.035 ;
        RECT 63.030 120.990 63.320 121.035 ;
        RECT 84.150 121.175 84.440 121.220 ;
        RECT 86.930 121.175 87.220 121.220 ;
        RECT 88.790 121.175 89.080 121.220 ;
        RECT 84.150 121.035 89.080 121.175 ;
        RECT 84.150 120.990 84.440 121.035 ;
        RECT 86.930 120.990 87.220 121.035 ;
        RECT 88.790 120.990 89.080 121.035 ;
        RECT 94.270 121.175 94.560 121.220 ;
        RECT 97.050 121.175 97.340 121.220 ;
        RECT 98.910 121.175 99.200 121.220 ;
        RECT 94.270 121.035 99.200 121.175 ;
        RECT 94.270 120.990 94.560 121.035 ;
        RECT 97.050 120.990 97.340 121.035 ;
        RECT 98.910 120.990 99.200 121.035 ;
        RECT 103.930 121.175 104.220 121.220 ;
        RECT 106.710 121.175 107.000 121.220 ;
        RECT 108.570 121.175 108.860 121.220 ;
        RECT 103.930 121.035 108.860 121.175 ;
        RECT 103.930 120.990 104.220 121.035 ;
        RECT 106.710 120.990 107.000 121.035 ;
        RECT 108.570 120.990 108.860 121.035 ;
        RECT 25.315 120.650 25.605 120.880 ;
        RECT 26.220 120.835 26.540 120.895 ;
        RECT 32.660 120.835 32.980 120.895 ;
        RECT 26.220 120.695 32.980 120.835 ;
        RECT 26.220 120.635 26.540 120.695 ;
        RECT 32.660 120.635 32.980 120.695 ;
        RECT 63.480 120.635 63.800 120.895 ;
        RECT 70.855 120.835 71.145 120.880 ;
        RECT 76.820 120.835 77.140 120.895 ;
        RECT 70.855 120.695 77.140 120.835 ;
        RECT 70.855 120.650 71.145 120.695 ;
        RECT 76.820 120.635 77.140 120.695 ;
        RECT 78.660 120.835 78.980 120.895 ;
        RECT 78.660 120.695 87.170 120.835 ;
        RECT 78.660 120.635 78.980 120.695 ;
        RECT 87.030 120.555 87.170 120.695 ;
        RECT 87.400 120.635 87.720 120.895 ;
        RECT 109.020 120.835 109.340 120.895 ;
        RECT 113.160 120.835 113.480 120.895 ;
        RECT 109.020 120.695 113.480 120.835 ;
        RECT 109.020 120.635 109.340 120.695 ;
        RECT 113.160 120.635 113.480 120.695 ;
        RECT 13.355 120.495 13.645 120.540 ;
        RECT 18.460 120.495 18.750 120.540 ;
        RECT 13.355 120.355 14.030 120.495 ;
        RECT 13.355 120.310 13.645 120.355 ;
        RECT 13.890 119.815 14.030 120.355 ;
        RECT 16.215 120.355 18.750 120.495 ;
        RECT 16.215 120.200 16.430 120.355 ;
        RECT 18.460 120.310 18.750 120.355 ;
        RECT 31.710 120.495 32.000 120.540 ;
        RECT 34.500 120.495 34.820 120.555 ;
        RECT 34.975 120.495 35.265 120.540 ;
        RECT 31.710 120.355 34.245 120.495 ;
        RECT 31.710 120.310 32.000 120.355 ;
        RECT 14.280 120.155 14.570 120.200 ;
        RECT 16.140 120.155 16.430 120.200 ;
        RECT 14.280 120.015 16.430 120.155 ;
        RECT 14.280 119.970 14.570 120.015 ;
        RECT 16.140 119.970 16.430 120.015 ;
        RECT 17.020 120.200 17.340 120.215 ;
        RECT 17.020 120.155 17.350 120.200 ;
        RECT 20.320 120.155 20.610 120.200 ;
        RECT 17.020 120.015 20.610 120.155 ;
        RECT 17.020 119.970 17.350 120.015 ;
        RECT 20.320 119.970 20.610 120.015 ;
        RECT 27.140 120.155 27.460 120.215 ;
        RECT 34.030 120.200 34.245 120.355 ;
        RECT 34.500 120.355 35.265 120.495 ;
        RECT 34.500 120.295 34.820 120.355 ;
        RECT 34.975 120.310 35.265 120.355 ;
        RECT 36.815 120.495 37.105 120.540 ;
        RECT 37.260 120.495 37.580 120.555 ;
        RECT 36.815 120.355 37.580 120.495 ;
        RECT 36.815 120.310 37.105 120.355 ;
        RECT 37.260 120.295 37.580 120.355 ;
        RECT 40.020 120.295 40.340 120.555 ;
        RECT 48.300 120.495 48.620 120.555 ;
        RECT 51.535 120.495 51.825 120.540 ;
        RECT 48.300 120.355 51.825 120.495 ;
        RECT 48.300 120.295 48.620 120.355 ;
        RECT 51.535 120.310 51.825 120.355 ;
        RECT 52.915 120.495 53.205 120.540 ;
        RECT 53.820 120.495 54.140 120.555 ;
        RECT 52.915 120.355 54.140 120.495 ;
        RECT 52.915 120.310 53.205 120.355 ;
        RECT 29.850 120.155 30.140 120.200 ;
        RECT 33.110 120.155 33.400 120.200 ;
        RECT 27.140 120.015 33.400 120.155 ;
        RECT 17.020 119.955 17.340 119.970 ;
        RECT 27.140 119.955 27.460 120.015 ;
        RECT 29.850 119.970 30.140 120.015 ;
        RECT 33.110 119.970 33.400 120.015 ;
        RECT 34.030 120.155 34.320 120.200 ;
        RECT 35.890 120.155 36.180 120.200 ;
        RECT 40.480 120.155 40.800 120.215 ;
        RECT 34.030 120.015 36.180 120.155 ;
        RECT 34.030 119.970 34.320 120.015 ;
        RECT 35.890 119.970 36.180 120.015 ;
        RECT 36.430 120.015 40.800 120.155 ;
        RECT 18.400 119.815 18.720 119.875 ;
        RECT 13.890 119.675 18.720 119.815 ;
        RECT 18.400 119.615 18.720 119.675 ;
        RECT 24.840 119.815 25.160 119.875 ;
        RECT 36.430 119.815 36.570 120.015 ;
        RECT 40.480 119.955 40.800 120.015 ;
        RECT 24.840 119.675 36.570 119.815 ;
        RECT 38.180 119.815 38.500 119.875 ;
        RECT 39.115 119.815 39.405 119.860 ;
        RECT 38.180 119.675 39.405 119.815 ;
        RECT 51.610 119.815 51.750 120.310 ;
        RECT 53.820 120.295 54.140 120.355 ;
        RECT 58.390 120.495 58.680 120.540 ;
        RECT 61.655 120.495 61.945 120.540 ;
        RECT 58.390 120.355 60.925 120.495 ;
        RECT 58.390 120.310 58.680 120.355 ;
        RECT 60.710 120.200 60.925 120.355 ;
        RECT 61.655 120.355 64.630 120.495 ;
        RECT 61.655 120.310 61.945 120.355 ;
        RECT 53.375 120.155 53.665 120.200 ;
        RECT 56.530 120.155 56.820 120.200 ;
        RECT 59.790 120.155 60.080 120.200 ;
        RECT 53.375 120.015 60.080 120.155 ;
        RECT 53.375 119.970 53.665 120.015 ;
        RECT 56.530 119.970 56.820 120.015 ;
        RECT 59.790 119.970 60.080 120.015 ;
        RECT 60.710 120.155 61.000 120.200 ;
        RECT 62.570 120.155 62.860 120.200 ;
        RECT 60.710 120.015 62.860 120.155 ;
        RECT 60.710 119.970 61.000 120.015 ;
        RECT 62.570 119.970 62.860 120.015 ;
        RECT 59.340 119.815 59.660 119.875 ;
        RECT 63.480 119.815 63.800 119.875 ;
        RECT 64.490 119.860 64.630 120.355 ;
        RECT 65.320 120.295 65.640 120.555 ;
        RECT 68.555 120.310 68.845 120.540 ;
        RECT 71.315 120.495 71.605 120.540 ;
        RECT 72.220 120.495 72.540 120.555 ;
        RECT 77.755 120.495 78.045 120.540 ;
        RECT 83.260 120.495 83.580 120.555 ;
        RECT 71.315 120.355 78.045 120.495 ;
        RECT 71.315 120.310 71.605 120.355 ;
        RECT 68.630 120.155 68.770 120.310 ;
        RECT 72.220 120.295 72.540 120.355 ;
        RECT 77.755 120.310 78.045 120.355 ;
        RECT 81.970 120.355 83.580 120.495 ;
        RECT 75.440 120.155 75.760 120.215 ;
        RECT 68.630 120.015 75.760 120.155 ;
        RECT 75.440 119.955 75.760 120.015 ;
        RECT 77.295 120.155 77.585 120.200 ;
        RECT 80.285 120.155 80.575 120.200 ;
        RECT 81.970 120.155 82.110 120.355 ;
        RECT 83.260 120.295 83.580 120.355 ;
        RECT 84.150 120.495 84.440 120.540 ;
        RECT 86.940 120.495 87.260 120.555 ;
        RECT 89.255 120.495 89.545 120.540 ;
        RECT 84.150 120.355 86.685 120.495 ;
        RECT 84.150 120.310 84.440 120.355 ;
        RECT 82.340 120.200 82.660 120.215 ;
        RECT 86.470 120.200 86.685 120.355 ;
        RECT 86.940 120.355 89.545 120.495 ;
        RECT 86.940 120.295 87.260 120.355 ;
        RECT 89.255 120.310 89.545 120.355 ;
        RECT 94.270 120.495 94.560 120.540 ;
        RECT 94.270 120.355 96.805 120.495 ;
        RECT 94.270 120.310 94.560 120.355 ;
        RECT 77.295 120.015 82.110 120.155 ;
        RECT 82.290 120.155 82.660 120.200 ;
        RECT 85.550 120.155 85.840 120.200 ;
        RECT 82.290 120.015 85.840 120.155 ;
        RECT 77.295 119.970 77.585 120.015 ;
        RECT 80.285 119.970 80.575 120.015 ;
        RECT 82.290 119.970 82.660 120.015 ;
        RECT 85.550 119.970 85.840 120.015 ;
        RECT 86.470 120.155 86.760 120.200 ;
        RECT 88.330 120.155 88.620 120.200 ;
        RECT 86.470 120.015 88.620 120.155 ;
        RECT 86.470 119.970 86.760 120.015 ;
        RECT 88.330 119.970 88.620 120.015 ;
        RECT 92.410 120.155 92.700 120.200 ;
        RECT 93.840 120.155 94.160 120.215 ;
        RECT 96.590 120.200 96.805 120.355 ;
        RECT 97.520 120.295 97.840 120.555 ;
        RECT 99.360 120.295 99.680 120.555 ;
        RECT 103.930 120.495 104.220 120.540 ;
        RECT 103.930 120.355 106.465 120.495 ;
        RECT 103.930 120.310 104.220 120.355 ;
        RECT 95.670 120.155 95.960 120.200 ;
        RECT 92.410 120.015 95.960 120.155 ;
        RECT 92.410 119.970 92.700 120.015 ;
        RECT 82.340 119.955 82.660 119.970 ;
        RECT 93.840 119.955 94.160 120.015 ;
        RECT 95.670 119.970 95.960 120.015 ;
        RECT 96.590 120.155 96.880 120.200 ;
        RECT 98.450 120.155 98.740 120.200 ;
        RECT 96.590 120.015 98.740 120.155 ;
        RECT 96.590 119.970 96.880 120.015 ;
        RECT 98.450 119.970 98.740 120.015 ;
        RECT 98.900 120.155 99.220 120.215 ;
        RECT 106.250 120.200 106.465 120.355 ;
        RECT 107.180 120.295 107.500 120.555 ;
        RECT 102.070 120.155 102.360 120.200 ;
        RECT 105.330 120.155 105.620 120.200 ;
        RECT 98.900 120.015 105.620 120.155 ;
        RECT 98.900 119.955 99.220 120.015 ;
        RECT 102.070 119.970 102.360 120.015 ;
        RECT 105.330 119.970 105.620 120.015 ;
        RECT 106.250 120.155 106.540 120.200 ;
        RECT 108.110 120.155 108.400 120.200 ;
        RECT 106.250 120.015 108.400 120.155 ;
        RECT 106.250 119.970 106.540 120.015 ;
        RECT 108.110 119.970 108.400 120.015 ;
        RECT 51.610 119.675 63.800 119.815 ;
        RECT 24.840 119.615 25.160 119.675 ;
        RECT 38.180 119.615 38.500 119.675 ;
        RECT 39.115 119.630 39.405 119.675 ;
        RECT 59.340 119.615 59.660 119.675 ;
        RECT 63.480 119.615 63.800 119.675 ;
        RECT 64.415 119.630 64.705 119.860 ;
        RECT 71.760 119.615 72.080 119.875 ;
        RECT 73.615 119.815 73.905 119.860 ;
        RECT 74.060 119.815 74.380 119.875 ;
        RECT 73.615 119.675 74.380 119.815 ;
        RECT 73.615 119.630 73.905 119.675 ;
        RECT 74.060 119.615 74.380 119.675 ;
        RECT 79.595 119.815 79.885 119.860 ;
        RECT 87.860 119.815 88.180 119.875 ;
        RECT 79.595 119.675 88.180 119.815 ;
        RECT 79.595 119.630 79.885 119.675 ;
        RECT 87.860 119.615 88.180 119.675 ;
        RECT 97.980 119.815 98.300 119.875 ;
        RECT 100.065 119.815 100.355 119.860 ;
        RECT 97.980 119.675 100.355 119.815 ;
        RECT 97.980 119.615 98.300 119.675 ;
        RECT 100.065 119.630 100.355 119.675 ;
        RECT 10.510 118.995 115.850 119.475 ;
        RECT 18.860 118.795 19.180 118.855 ;
        RECT 14.350 118.655 19.180 118.795 ;
        RECT 14.350 118.115 14.490 118.655 ;
        RECT 18.860 118.595 19.180 118.655 ;
        RECT 22.785 118.795 23.075 118.840 ;
        RECT 24.840 118.795 25.160 118.855 ;
        RECT 22.785 118.655 25.160 118.795 ;
        RECT 22.785 118.610 23.075 118.655 ;
        RECT 24.840 118.595 25.160 118.655 ;
        RECT 26.005 118.795 26.295 118.840 ;
        RECT 28.520 118.795 28.840 118.855 ;
        RECT 26.005 118.655 28.840 118.795 ;
        RECT 26.005 118.610 26.295 118.655 ;
        RECT 28.520 118.595 28.840 118.655 ;
        RECT 34.500 118.795 34.820 118.855 ;
        RECT 35.435 118.795 35.725 118.840 ;
        RECT 34.500 118.655 35.725 118.795 ;
        RECT 34.500 118.595 34.820 118.655 ;
        RECT 35.435 118.610 35.725 118.655 ;
        RECT 39.115 118.795 39.405 118.840 ;
        RECT 40.480 118.795 40.800 118.855 ;
        RECT 39.115 118.655 40.800 118.795 ;
        RECT 39.115 118.610 39.405 118.655 ;
        RECT 40.480 118.595 40.800 118.655 ;
        RECT 41.415 118.610 41.705 118.840 ;
        RECT 14.740 118.455 15.030 118.500 ;
        RECT 16.600 118.455 16.890 118.500 ;
        RECT 14.740 118.315 16.890 118.455 ;
        RECT 14.740 118.270 15.030 118.315 ;
        RECT 16.600 118.270 16.890 118.315 ;
        RECT 17.520 118.455 17.810 118.500 ;
        RECT 19.320 118.455 19.640 118.515 ;
        RECT 20.780 118.455 21.070 118.500 ;
        RECT 17.520 118.315 21.070 118.455 ;
        RECT 17.520 118.270 17.810 118.315 ;
        RECT 15.655 118.115 15.945 118.160 ;
        RECT 14.350 117.975 15.945 118.115 ;
        RECT 16.675 118.115 16.890 118.270 ;
        RECT 19.320 118.255 19.640 118.315 ;
        RECT 20.780 118.270 21.070 118.315 ;
        RECT 28.010 118.455 28.300 118.500 ;
        RECT 29.440 118.455 29.760 118.515 ;
        RECT 31.270 118.455 31.560 118.500 ;
        RECT 28.010 118.315 31.560 118.455 ;
        RECT 28.010 118.270 28.300 118.315 ;
        RECT 29.440 118.255 29.760 118.315 ;
        RECT 31.270 118.270 31.560 118.315 ;
        RECT 32.190 118.455 32.480 118.500 ;
        RECT 34.050 118.455 34.340 118.500 ;
        RECT 32.190 118.315 34.340 118.455 ;
        RECT 32.190 118.270 32.480 118.315 ;
        RECT 34.050 118.270 34.340 118.315 ;
        RECT 18.920 118.115 19.210 118.160 ;
        RECT 16.675 117.975 19.210 118.115 ;
        RECT 15.655 117.930 15.945 117.975 ;
        RECT 18.920 117.930 19.210 117.975 ;
        RECT 29.870 118.115 30.160 118.160 ;
        RECT 32.190 118.115 32.405 118.270 ;
        RECT 29.870 117.975 32.405 118.115 ;
        RECT 29.870 117.930 30.160 117.975 ;
        RECT 33.120 117.915 33.440 118.175 ;
        RECT 36.355 118.115 36.645 118.160 ;
        RECT 37.720 118.115 38.040 118.175 ;
        RECT 36.355 117.975 38.040 118.115 ;
        RECT 36.355 117.930 36.645 117.975 ;
        RECT 37.720 117.915 38.040 117.975 ;
        RECT 39.560 117.915 39.880 118.175 ;
        RECT 41.490 118.115 41.630 118.610 ;
        RECT 48.300 118.595 48.620 118.855 ;
        RECT 49.220 118.795 49.540 118.855 ;
        RECT 51.535 118.795 51.825 118.840 ;
        RECT 49.220 118.655 51.825 118.795 ;
        RECT 49.220 118.595 49.540 118.655 ;
        RECT 51.535 118.610 51.825 118.655 ;
        RECT 59.800 118.795 60.120 118.855 ;
        RECT 62.345 118.795 62.635 118.840 ;
        RECT 59.800 118.655 62.635 118.795 ;
        RECT 59.800 118.595 60.120 118.655 ;
        RECT 62.345 118.610 62.635 118.655 ;
        RECT 66.025 118.795 66.315 118.840 ;
        RECT 71.760 118.795 72.080 118.855 ;
        RECT 66.025 118.655 72.080 118.795 ;
        RECT 66.025 118.610 66.315 118.655 ;
        RECT 71.760 118.595 72.080 118.655 ;
        RECT 87.400 118.795 87.720 118.855 ;
        RECT 88.795 118.795 89.085 118.840 ;
        RECT 87.400 118.655 89.085 118.795 ;
        RECT 87.400 118.595 87.720 118.655 ;
        RECT 88.795 118.610 89.085 118.655 ;
        RECT 97.075 118.795 97.365 118.840 ;
        RECT 97.520 118.795 97.840 118.855 ;
        RECT 97.075 118.655 97.840 118.795 ;
        RECT 97.075 118.610 97.365 118.655 ;
        RECT 97.520 118.595 97.840 118.655 ;
        RECT 97.980 118.795 98.300 118.855 ;
        RECT 100.295 118.795 100.585 118.840 ;
        RECT 97.980 118.655 100.585 118.795 ;
        RECT 97.980 118.595 98.300 118.655 ;
        RECT 100.295 118.610 100.585 118.655 ;
        RECT 106.720 118.595 107.040 118.855 ;
        RECT 41.860 118.255 42.180 118.515 ;
        RECT 48.390 118.455 48.530 118.595 ;
        RECT 57.040 118.500 57.360 118.515 ;
        RECT 54.300 118.455 54.590 118.500 ;
        RECT 56.160 118.455 56.450 118.500 ;
        RECT 48.390 118.315 53.590 118.455 ;
        RECT 53.450 118.160 53.590 118.315 ;
        RECT 54.300 118.315 56.450 118.455 ;
        RECT 54.300 118.270 54.590 118.315 ;
        RECT 56.160 118.270 56.450 118.315 ;
        RECT 52.455 118.115 52.745 118.160 ;
        RECT 41.490 117.975 52.745 118.115 ;
        RECT 52.455 117.930 52.745 117.975 ;
        RECT 53.375 117.930 53.665 118.160 ;
        RECT 55.200 117.915 55.520 118.175 ;
        RECT 56.235 118.115 56.450 118.270 ;
        RECT 57.040 118.455 57.370 118.500 ;
        RECT 60.340 118.455 60.630 118.500 ;
        RECT 57.040 118.315 60.630 118.455 ;
        RECT 57.040 118.270 57.370 118.315 ;
        RECT 60.340 118.270 60.630 118.315 ;
        RECT 68.030 118.455 68.320 118.500 ;
        RECT 69.460 118.455 69.780 118.515 ;
        RECT 71.290 118.455 71.580 118.500 ;
        RECT 68.030 118.315 71.580 118.455 ;
        RECT 68.030 118.270 68.320 118.315 ;
        RECT 57.040 118.255 57.360 118.270 ;
        RECT 69.460 118.255 69.780 118.315 ;
        RECT 71.290 118.270 71.580 118.315 ;
        RECT 72.210 118.455 72.500 118.500 ;
        RECT 74.070 118.455 74.360 118.500 ;
        RECT 72.210 118.315 74.360 118.455 ;
        RECT 72.210 118.270 72.500 118.315 ;
        RECT 74.070 118.270 74.360 118.315 ;
        RECT 75.915 118.455 76.205 118.500 ;
        RECT 79.530 118.455 79.820 118.500 ;
        RECT 82.790 118.455 83.080 118.500 ;
        RECT 75.915 118.315 83.080 118.455 ;
        RECT 75.915 118.270 76.205 118.315 ;
        RECT 79.530 118.270 79.820 118.315 ;
        RECT 82.790 118.270 83.080 118.315 ;
        RECT 83.710 118.455 84.000 118.500 ;
        RECT 85.570 118.455 85.860 118.500 ;
        RECT 83.710 118.315 85.860 118.455 ;
        RECT 83.710 118.270 84.000 118.315 ;
        RECT 85.570 118.270 85.860 118.315 ;
        RECT 95.235 118.455 95.525 118.500 ;
        RECT 98.900 118.455 99.220 118.515 ;
        RECT 95.235 118.315 99.220 118.455 ;
        RECT 95.235 118.270 95.525 118.315 ;
        RECT 58.480 118.115 58.770 118.160 ;
        RECT 56.235 117.975 58.770 118.115 ;
        RECT 58.480 117.930 58.770 117.975 ;
        RECT 69.890 118.115 70.180 118.160 ;
        RECT 72.210 118.115 72.425 118.270 ;
        RECT 69.890 117.975 72.425 118.115 ;
        RECT 69.890 117.930 70.180 117.975 ;
        RECT 75.440 117.915 75.760 118.175 ;
        RECT 81.390 118.115 81.680 118.160 ;
        RECT 83.710 118.115 83.925 118.270 ;
        RECT 98.900 118.255 99.220 118.315 ;
        RECT 99.360 118.455 99.680 118.515 ;
        RECT 103.975 118.455 104.265 118.500 ;
        RECT 109.020 118.455 109.340 118.515 ;
        RECT 99.360 118.315 109.340 118.455 ;
        RECT 99.360 118.255 99.680 118.315 ;
        RECT 103.975 118.270 104.265 118.315 ;
        RECT 109.020 118.255 109.340 118.315 ;
        RECT 81.390 117.975 83.925 118.115 ;
        RECT 86.495 118.115 86.785 118.160 ;
        RECT 86.940 118.115 87.260 118.175 ;
        RECT 86.495 117.975 87.260 118.115 ;
        RECT 81.390 117.930 81.680 117.975 ;
        RECT 86.495 117.930 86.785 117.975 ;
        RECT 86.940 117.915 87.260 117.975 ;
        RECT 87.860 117.915 88.180 118.175 ;
        RECT 89.700 117.915 90.020 118.175 ;
        RECT 94.775 117.930 95.065 118.160 ;
        RECT 96.155 118.115 96.445 118.160 ;
        RECT 97.060 118.115 97.380 118.175 ;
        RECT 96.155 117.975 97.380 118.115 ;
        RECT 96.155 117.930 96.445 117.975 ;
        RECT 13.815 117.775 14.105 117.820 ;
        RECT 18.400 117.775 18.720 117.835 ;
        RECT 24.380 117.775 24.700 117.835 ;
        RECT 34.975 117.775 35.265 117.820 ;
        RECT 37.260 117.775 37.580 117.835 ;
        RECT 13.815 117.635 37.580 117.775 ;
        RECT 13.815 117.590 14.105 117.635 ;
        RECT 18.400 117.575 18.720 117.635 ;
        RECT 24.380 117.575 24.700 117.635 ;
        RECT 34.975 117.590 35.265 117.635 ;
        RECT 37.260 117.575 37.580 117.635 ;
        RECT 38.195 117.590 38.485 117.820 ;
        RECT 14.280 117.435 14.570 117.480 ;
        RECT 16.140 117.435 16.430 117.480 ;
        RECT 18.920 117.435 19.210 117.480 ;
        RECT 14.280 117.295 19.210 117.435 ;
        RECT 14.280 117.250 14.570 117.295 ;
        RECT 16.140 117.250 16.430 117.295 ;
        RECT 18.920 117.250 19.210 117.295 ;
        RECT 29.870 117.435 30.160 117.480 ;
        RECT 32.650 117.435 32.940 117.480 ;
        RECT 34.510 117.435 34.800 117.480 ;
        RECT 38.270 117.435 38.410 117.590 ;
        RECT 73.140 117.575 73.460 117.835 ;
        RECT 73.600 117.775 73.920 117.835 ;
        RECT 74.995 117.775 75.285 117.820 ;
        RECT 78.660 117.775 78.980 117.835 ;
        RECT 73.600 117.635 78.980 117.775 ;
        RECT 73.600 117.575 73.920 117.635 ;
        RECT 74.995 117.590 75.285 117.635 ;
        RECT 78.660 117.575 78.980 117.635 ;
        RECT 84.655 117.775 84.945 117.820 ;
        RECT 84.655 117.635 87.170 117.775 ;
        RECT 84.655 117.590 84.945 117.635 ;
        RECT 87.030 117.480 87.170 117.635 ;
        RECT 29.870 117.295 34.800 117.435 ;
        RECT 29.870 117.250 30.160 117.295 ;
        RECT 32.650 117.250 32.940 117.295 ;
        RECT 34.510 117.250 34.800 117.295 ;
        RECT 35.050 117.295 38.410 117.435 ;
        RECT 53.840 117.435 54.130 117.480 ;
        RECT 55.700 117.435 55.990 117.480 ;
        RECT 58.480 117.435 58.770 117.480 ;
        RECT 53.840 117.295 58.770 117.435 ;
        RECT 35.050 117.155 35.190 117.295 ;
        RECT 53.840 117.250 54.130 117.295 ;
        RECT 55.700 117.250 55.990 117.295 ;
        RECT 58.480 117.250 58.770 117.295 ;
        RECT 69.890 117.435 70.180 117.480 ;
        RECT 72.670 117.435 72.960 117.480 ;
        RECT 74.530 117.435 74.820 117.480 ;
        RECT 69.890 117.295 74.820 117.435 ;
        RECT 69.890 117.250 70.180 117.295 ;
        RECT 72.670 117.250 72.960 117.295 ;
        RECT 74.530 117.250 74.820 117.295 ;
        RECT 81.390 117.435 81.680 117.480 ;
        RECT 84.170 117.435 84.460 117.480 ;
        RECT 86.030 117.435 86.320 117.480 ;
        RECT 81.390 117.295 86.320 117.435 ;
        RECT 81.390 117.250 81.680 117.295 ;
        RECT 84.170 117.250 84.460 117.295 ;
        RECT 86.030 117.250 86.320 117.295 ;
        RECT 86.955 117.250 87.245 117.480 ;
        RECT 94.850 117.435 94.990 117.930 ;
        RECT 97.060 117.915 97.380 117.975 ;
        RECT 99.835 118.115 100.125 118.160 ;
        RECT 100.280 118.115 100.600 118.175 ;
        RECT 99.835 117.975 100.600 118.115 ;
        RECT 99.835 117.930 100.125 117.975 ;
        RECT 100.280 117.915 100.600 117.975 ;
        RECT 106.260 117.915 106.580 118.175 ;
        RECT 98.440 117.775 98.760 117.835 ;
        RECT 98.915 117.775 99.205 117.820 ;
        RECT 98.440 117.635 99.205 117.775 ;
        RECT 98.440 117.575 98.760 117.635 ;
        RECT 98.915 117.590 99.205 117.635 ;
        RECT 106.350 117.435 106.490 117.915 ;
        RECT 94.850 117.295 106.490 117.435 ;
        RECT 34.960 116.895 35.280 117.155 ;
        RECT 72.220 117.095 72.540 117.155 ;
        RECT 77.525 117.095 77.815 117.140 ;
        RECT 72.220 116.955 77.815 117.095 ;
        RECT 72.220 116.895 72.540 116.955 ;
        RECT 77.525 116.910 77.815 116.955 ;
        RECT 102.120 116.895 102.440 117.155 ;
        RECT 10.510 116.275 115.850 116.755 ;
        RECT 17.955 116.075 18.245 116.120 ;
        RECT 19.320 116.075 19.640 116.135 ;
        RECT 17.955 115.935 19.640 116.075 ;
        RECT 17.955 115.890 18.245 115.935 ;
        RECT 19.320 115.875 19.640 115.935 ;
        RECT 29.440 115.875 29.760 116.135 ;
        RECT 33.120 115.875 33.440 116.135 ;
        RECT 37.735 116.075 38.025 116.120 ;
        RECT 40.020 116.075 40.340 116.135 ;
        RECT 37.735 115.935 40.340 116.075 ;
        RECT 37.735 115.890 38.025 115.935 ;
        RECT 40.020 115.875 40.340 115.935 ;
        RECT 57.040 116.075 57.360 116.135 ;
        RECT 57.515 116.075 57.805 116.120 ;
        RECT 57.040 115.935 57.805 116.075 ;
        RECT 57.040 115.875 57.360 115.935 ;
        RECT 57.515 115.890 57.805 115.935 ;
        RECT 69.460 115.875 69.780 116.135 ;
        RECT 72.695 116.075 72.985 116.120 ;
        RECT 73.140 116.075 73.460 116.135 ;
        RECT 72.695 115.935 73.460 116.075 ;
        RECT 72.695 115.890 72.985 115.935 ;
        RECT 73.140 115.875 73.460 115.935 ;
        RECT 81.895 116.075 82.185 116.120 ;
        RECT 82.340 116.075 82.660 116.135 ;
        RECT 81.895 115.935 82.660 116.075 ;
        RECT 81.895 115.890 82.185 115.935 ;
        RECT 82.340 115.875 82.660 115.935 ;
        RECT 102.135 116.075 102.425 116.120 ;
        RECT 107.180 116.075 107.500 116.135 ;
        RECT 102.135 115.935 107.500 116.075 ;
        RECT 102.135 115.890 102.425 115.935 ;
        RECT 107.180 115.875 107.500 115.935 ;
        RECT 34.040 115.735 34.360 115.795 ;
        RECT 41.875 115.735 42.165 115.780 ;
        RECT 34.040 115.595 42.165 115.735 ;
        RECT 34.040 115.535 34.360 115.595 ;
        RECT 41.875 115.550 42.165 115.595 ;
        RECT 105.340 115.735 105.660 115.795 ;
        RECT 110.415 115.735 110.705 115.780 ;
        RECT 105.340 115.595 110.705 115.735 ;
        RECT 105.340 115.535 105.660 115.595 ;
        RECT 110.415 115.550 110.705 115.595 ;
        RECT 32.660 115.395 32.980 115.455 ;
        RECT 34.515 115.395 34.805 115.440 ;
        RECT 34.960 115.395 35.280 115.455 ;
        RECT 32.660 115.255 35.280 115.395 ;
        RECT 32.660 115.195 32.980 115.255 ;
        RECT 34.515 115.210 34.805 115.255 ;
        RECT 34.960 115.195 35.280 115.255 ;
        RECT 35.435 115.395 35.725 115.440 ;
        RECT 39.560 115.395 39.880 115.455 ;
        RECT 75.440 115.395 75.760 115.455 ;
        RECT 35.435 115.255 39.880 115.395 ;
        RECT 35.435 115.210 35.725 115.255 ;
        RECT 39.560 115.195 39.880 115.255 ;
        RECT 69.090 115.255 75.760 115.395 ;
        RECT 18.415 115.055 18.705 115.100 ;
        RECT 23.920 115.055 24.240 115.115 ;
        RECT 28.995 115.055 29.285 115.100 ;
        RECT 18.415 114.915 29.285 115.055 ;
        RECT 18.415 114.870 18.705 114.915 ;
        RECT 23.920 114.855 24.240 114.915 ;
        RECT 28.995 114.870 29.285 114.915 ;
        RECT 30.360 115.055 30.680 115.115 ;
        RECT 32.215 115.055 32.505 115.100 ;
        RECT 30.360 114.915 32.505 115.055 ;
        RECT 29.070 114.715 29.210 114.870 ;
        RECT 30.360 114.855 30.680 114.915 ;
        RECT 32.215 114.870 32.505 114.915 ;
        RECT 33.580 115.055 33.900 115.115 ;
        RECT 35.895 115.055 36.185 115.100 ;
        RECT 33.580 114.915 36.185 115.055 ;
        RECT 33.580 114.855 33.900 114.915 ;
        RECT 35.895 114.870 36.185 114.915 ;
        RECT 42.335 115.055 42.625 115.100 ;
        RECT 43.700 115.055 44.020 115.115 ;
        RECT 46.015 115.055 46.305 115.100 ;
        RECT 42.335 114.915 46.305 115.055 ;
        RECT 42.335 114.870 42.625 114.915 ;
        RECT 42.410 114.715 42.550 114.870 ;
        RECT 43.700 114.855 44.020 114.915 ;
        RECT 46.015 114.870 46.305 114.915 ;
        RECT 47.395 115.055 47.685 115.100 ;
        RECT 53.820 115.055 54.140 115.115 ;
        RECT 69.090 115.100 69.230 115.255 ;
        RECT 75.440 115.195 75.760 115.255 ;
        RECT 57.055 115.055 57.345 115.100 ;
        RECT 47.395 114.915 57.345 115.055 ;
        RECT 47.395 114.870 47.685 114.915 ;
        RECT 53.820 114.855 54.140 114.915 ;
        RECT 57.055 114.870 57.345 114.915 ;
        RECT 69.015 114.870 69.305 115.100 ;
        RECT 73.615 115.055 73.905 115.100 ;
        RECT 74.060 115.055 74.380 115.115 ;
        RECT 73.615 114.915 74.380 115.055 ;
        RECT 75.530 115.055 75.670 115.195 ;
        RECT 81.435 115.055 81.725 115.100 ;
        RECT 75.530 114.915 81.725 115.055 ;
        RECT 73.615 114.870 73.905 114.915 ;
        RECT 74.060 114.855 74.380 114.915 ;
        RECT 81.435 114.870 81.725 114.915 ;
        RECT 101.215 115.055 101.505 115.100 ;
        RECT 102.120 115.055 102.440 115.115 ;
        RECT 101.215 114.915 102.440 115.055 ;
        RECT 101.215 114.870 101.505 114.915 ;
        RECT 102.120 114.855 102.440 114.915 ;
        RECT 107.640 114.855 107.960 115.115 ;
        RECT 108.100 114.855 108.420 115.115 ;
        RECT 111.335 115.055 111.625 115.100 ;
        RECT 112.240 115.055 112.560 115.115 ;
        RECT 111.335 114.915 112.560 115.055 ;
        RECT 111.335 114.870 111.625 114.915 ;
        RECT 112.240 114.855 112.560 114.915 ;
        RECT 29.070 114.575 42.550 114.715 ;
        RECT 105.800 114.375 106.120 114.435 ;
        RECT 106.735 114.375 107.025 114.420 ;
        RECT 105.800 114.235 107.025 114.375 ;
        RECT 105.800 114.175 106.120 114.235 ;
        RECT 106.735 114.190 107.025 114.235 ;
        RECT 108.560 114.175 108.880 114.435 ;
        RECT 10.510 113.555 115.850 114.035 ;
        RECT 67.620 113.355 67.940 113.415 ;
        RECT 67.620 113.215 85.330 113.355 ;
        RECT 67.620 113.155 67.940 113.215 ;
        RECT 53.820 113.015 54.140 113.075 ;
        RECT 52.990 112.875 54.140 113.015 ;
        RECT 23.460 112.475 23.780 112.735 ;
        RECT 31.740 112.475 32.060 112.735 ;
        RECT 32.200 112.675 32.520 112.735 ;
        RECT 38.195 112.675 38.485 112.720 ;
        RECT 32.200 112.535 38.485 112.675 ;
        RECT 32.200 112.475 32.520 112.535 ;
        RECT 38.195 112.490 38.485 112.535 ;
        RECT 47.380 112.675 47.700 112.735 ;
        RECT 52.990 112.720 53.130 112.875 ;
        RECT 53.820 112.815 54.140 112.875 ;
        RECT 59.200 112.875 71.530 113.015 ;
        RECT 49.695 112.675 49.985 112.720 ;
        RECT 47.380 112.535 49.985 112.675 ;
        RECT 47.380 112.475 47.700 112.535 ;
        RECT 49.695 112.490 49.985 112.535 ;
        RECT 52.915 112.675 53.205 112.720 ;
        RECT 59.200 112.675 59.340 112.875 ;
        RECT 52.915 112.535 59.340 112.675 ;
        RECT 52.915 112.490 53.205 112.535 ;
        RECT 68.540 112.475 68.860 112.735 ;
        RECT 71.390 112.720 71.530 112.875 ;
        RECT 85.190 112.720 85.330 113.215 ;
        RECT 105.340 112.815 105.660 113.075 ;
        RECT 107.635 113.015 108.285 113.060 ;
        RECT 108.560 113.015 108.880 113.075 ;
        RECT 111.235 113.015 111.525 113.060 ;
        RECT 107.635 112.875 111.525 113.015 ;
        RECT 107.635 112.830 108.285 112.875 ;
        RECT 108.560 112.815 108.880 112.875 ;
        RECT 110.935 112.830 111.525 112.875 ;
        RECT 69.935 112.490 70.225 112.720 ;
        RECT 71.315 112.490 71.605 112.720 ;
        RECT 85.115 112.490 85.405 112.720 ;
        RECT 51.980 112.335 52.300 112.395 ;
        RECT 53.835 112.335 54.125 112.380 ;
        RECT 51.980 112.195 54.125 112.335 ;
        RECT 51.980 112.135 52.300 112.195 ;
        RECT 53.835 112.150 54.125 112.195 ;
        RECT 68.080 112.335 68.400 112.395 ;
        RECT 70.010 112.335 70.150 112.490 ;
        RECT 90.160 112.475 90.480 112.735 ;
        RECT 94.300 112.675 94.620 112.735 ;
        RECT 95.695 112.675 95.985 112.720 ;
        RECT 94.300 112.535 95.985 112.675 ;
        RECT 94.300 112.475 94.620 112.535 ;
        RECT 95.695 112.490 95.985 112.535 ;
        RECT 99.820 112.475 100.140 112.735 ;
        RECT 101.215 112.675 101.505 112.720 ;
        RECT 102.580 112.675 102.900 112.735 ;
        RECT 101.215 112.535 102.900 112.675 ;
        RECT 101.215 112.490 101.505 112.535 ;
        RECT 102.580 112.475 102.900 112.535 ;
        RECT 104.440 112.675 104.730 112.720 ;
        RECT 106.275 112.675 106.565 112.720 ;
        RECT 109.855 112.675 110.145 112.720 ;
        RECT 104.440 112.535 110.145 112.675 ;
        RECT 104.440 112.490 104.730 112.535 ;
        RECT 106.275 112.490 106.565 112.535 ;
        RECT 109.855 112.490 110.145 112.535 ;
        RECT 110.935 112.515 111.225 112.830 ;
        RECT 68.080 112.195 70.150 112.335 ;
        RECT 68.080 112.135 68.400 112.195 ;
        RECT 72.680 112.135 73.000 112.395 ;
        RECT 103.960 112.335 104.280 112.395 ;
        RECT 109.020 112.335 109.340 112.395 ;
        RECT 103.960 112.195 109.340 112.335 ;
        RECT 103.960 112.135 104.280 112.195 ;
        RECT 109.020 112.135 109.340 112.195 ;
        RECT 114.095 112.335 114.385 112.380 ;
        RECT 115.460 112.335 115.780 112.395 ;
        RECT 114.095 112.195 115.780 112.335 ;
        RECT 114.095 112.150 114.385 112.195 ;
        RECT 115.460 112.135 115.780 112.195 ;
        RECT 69.475 111.995 69.765 112.040 ;
        RECT 72.220 111.995 72.540 112.055 ;
        RECT 69.475 111.855 72.540 111.995 ;
        RECT 69.475 111.810 69.765 111.855 ;
        RECT 72.220 111.795 72.540 111.855 ;
        RECT 104.845 111.995 105.135 112.040 ;
        RECT 106.735 111.995 107.025 112.040 ;
        RECT 109.855 111.995 110.145 112.040 ;
        RECT 104.845 111.855 110.145 111.995 ;
        RECT 104.845 111.810 105.135 111.855 ;
        RECT 106.735 111.810 107.025 111.855 ;
        RECT 109.855 111.810 110.145 111.855 ;
        RECT 22.080 111.655 22.400 111.715 ;
        RECT 22.555 111.655 22.845 111.700 ;
        RECT 22.080 111.515 22.845 111.655 ;
        RECT 22.080 111.455 22.400 111.515 ;
        RECT 22.555 111.470 22.845 111.515 ;
        RECT 32.675 111.655 32.965 111.700 ;
        RECT 34.500 111.655 34.820 111.715 ;
        RECT 32.675 111.515 34.820 111.655 ;
        RECT 32.675 111.470 32.965 111.515 ;
        RECT 34.500 111.455 34.820 111.515 ;
        RECT 36.340 111.655 36.660 111.715 ;
        RECT 37.275 111.655 37.565 111.700 ;
        RECT 36.340 111.515 37.565 111.655 ;
        RECT 36.340 111.455 36.660 111.515 ;
        RECT 37.275 111.470 37.565 111.515 ;
        RECT 50.615 111.655 50.905 111.700 ;
        RECT 54.740 111.655 55.060 111.715 ;
        RECT 50.615 111.515 55.060 111.655 ;
        RECT 50.615 111.470 50.905 111.515 ;
        RECT 54.740 111.455 55.060 111.515 ;
        RECT 70.855 111.655 71.145 111.700 ;
        RECT 71.760 111.655 72.080 111.715 ;
        RECT 70.855 111.515 72.080 111.655 ;
        RECT 70.855 111.470 71.145 111.515 ;
        RECT 71.760 111.455 72.080 111.515 ;
        RECT 86.020 111.455 86.340 111.715 ;
        RECT 91.080 111.455 91.400 111.715 ;
        RECT 96.600 111.455 96.920 111.715 ;
        RECT 100.755 111.655 101.045 111.700 ;
        RECT 101.200 111.655 101.520 111.715 ;
        RECT 100.755 111.515 101.520 111.655 ;
        RECT 100.755 111.470 101.045 111.515 ;
        RECT 101.200 111.455 101.520 111.515 ;
        RECT 102.135 111.655 102.425 111.700 ;
        RECT 103.500 111.655 103.820 111.715 ;
        RECT 102.135 111.515 103.820 111.655 ;
        RECT 102.135 111.470 102.425 111.515 ;
        RECT 103.500 111.455 103.820 111.515 ;
        RECT 10.510 110.835 115.850 111.315 ;
        RECT 32.660 110.635 32.980 110.695 ;
        RECT 41.415 110.635 41.705 110.680 ;
        RECT 32.660 110.495 41.705 110.635 ;
        RECT 32.660 110.435 32.980 110.495 ;
        RECT 41.415 110.450 41.705 110.495 ;
        RECT 61.640 110.635 61.960 110.695 ;
        RECT 66.715 110.635 67.005 110.680 ;
        RECT 61.640 110.495 67.005 110.635 ;
        RECT 61.640 110.435 61.960 110.495 ;
        RECT 66.715 110.450 67.005 110.495 ;
        RECT 86.940 110.635 87.260 110.695 ;
        RECT 86.940 110.495 89.010 110.635 ;
        RECT 86.940 110.435 87.260 110.495 ;
        RECT 18.515 110.295 18.805 110.340 ;
        RECT 21.635 110.295 21.925 110.340 ;
        RECT 23.525 110.295 23.815 110.340 ;
        RECT 18.515 110.155 23.815 110.295 ;
        RECT 18.515 110.110 18.805 110.155 ;
        RECT 21.635 110.110 21.925 110.155 ;
        RECT 23.525 110.110 23.815 110.155 ;
        RECT 31.855 110.295 32.145 110.340 ;
        RECT 34.975 110.295 35.265 110.340 ;
        RECT 36.865 110.295 37.155 110.340 ;
        RECT 31.855 110.155 37.155 110.295 ;
        RECT 31.855 110.110 32.145 110.155 ;
        RECT 34.975 110.110 35.265 110.155 ;
        RECT 36.865 110.110 37.155 110.155 ;
        RECT 50.255 110.295 50.545 110.340 ;
        RECT 53.375 110.295 53.665 110.340 ;
        RECT 55.265 110.295 55.555 110.340 ;
        RECT 50.255 110.155 55.555 110.295 ;
        RECT 50.255 110.110 50.545 110.155 ;
        RECT 53.375 110.110 53.665 110.155 ;
        RECT 55.265 110.110 55.555 110.155 ;
        RECT 65.795 110.110 66.085 110.340 ;
        RECT 68.505 110.295 68.795 110.340 ;
        RECT 70.395 110.295 70.685 110.340 ;
        RECT 73.515 110.295 73.805 110.340 ;
        RECT 68.505 110.155 73.805 110.295 ;
        RECT 68.505 110.110 68.795 110.155 ;
        RECT 70.395 110.110 70.685 110.155 ;
        RECT 73.515 110.110 73.805 110.155 ;
        RECT 83.375 110.295 83.665 110.340 ;
        RECT 86.495 110.295 86.785 110.340 ;
        RECT 88.385 110.295 88.675 110.340 ;
        RECT 83.375 110.155 88.675 110.295 ;
        RECT 83.375 110.110 83.665 110.155 ;
        RECT 86.495 110.110 86.785 110.155 ;
        RECT 88.385 110.110 88.675 110.155 ;
        RECT 24.380 109.755 24.700 110.015 ;
        RECT 31.280 109.955 31.600 110.015 ;
        RECT 25.850 109.815 31.600 109.955 ;
        RECT 14.275 109.615 14.565 109.660 ;
        RECT 15.640 109.615 15.960 109.675 ;
        RECT 25.850 109.660 25.990 109.815 ;
        RECT 31.280 109.755 31.600 109.815 ;
        RECT 36.340 109.755 36.660 110.015 ;
        RECT 37.720 109.755 38.040 110.015 ;
        RECT 46.015 109.955 46.305 110.000 ;
        RECT 48.760 109.955 49.080 110.015 ;
        RECT 46.015 109.815 49.080 109.955 ;
        RECT 46.015 109.770 46.305 109.815 ;
        RECT 48.760 109.755 49.080 109.815 ;
        RECT 54.740 109.755 55.060 110.015 ;
        RECT 56.135 109.955 56.425 110.000 ;
        RECT 59.340 109.955 59.660 110.015 ;
        RECT 56.135 109.815 59.660 109.955 ;
        RECT 65.870 109.955 66.010 110.110 ;
        RECT 69.015 109.955 69.305 110.000 ;
        RECT 65.870 109.815 69.305 109.955 ;
        RECT 56.135 109.770 56.425 109.815 ;
        RECT 59.340 109.755 59.660 109.815 ;
        RECT 69.015 109.770 69.305 109.815 ;
        RECT 71.300 109.955 71.620 110.015 ;
        RECT 77.755 109.955 78.045 110.000 ;
        RECT 71.300 109.815 78.045 109.955 ;
        RECT 71.300 109.755 71.620 109.815 ;
        RECT 77.755 109.770 78.045 109.815 ;
        RECT 79.135 109.955 79.425 110.000 ;
        RECT 81.880 109.955 82.200 110.015 ;
        RECT 79.135 109.815 82.200 109.955 ;
        RECT 79.135 109.770 79.425 109.815 ;
        RECT 81.880 109.755 82.200 109.815 ;
        RECT 86.020 109.955 86.340 110.015 ;
        RECT 87.875 109.955 88.165 110.000 ;
        RECT 86.020 109.815 88.165 109.955 ;
        RECT 88.870 109.955 89.010 110.495 ;
        RECT 94.415 110.295 94.705 110.340 ;
        RECT 97.535 110.295 97.825 110.340 ;
        RECT 99.425 110.295 99.715 110.340 ;
        RECT 94.415 110.155 99.715 110.295 ;
        RECT 94.415 110.110 94.705 110.155 ;
        RECT 97.535 110.110 97.825 110.155 ;
        RECT 99.425 110.110 99.715 110.155 ;
        RECT 104.845 110.295 105.135 110.340 ;
        RECT 106.735 110.295 107.025 110.340 ;
        RECT 109.855 110.295 110.145 110.340 ;
        RECT 104.845 110.155 110.145 110.295 ;
        RECT 104.845 110.110 105.135 110.155 ;
        RECT 106.735 110.110 107.025 110.155 ;
        RECT 109.855 110.110 110.145 110.155 ;
        RECT 89.255 109.955 89.545 110.000 ;
        RECT 88.870 109.815 89.545 109.955 ;
        RECT 86.020 109.755 86.340 109.815 ;
        RECT 87.875 109.770 88.165 109.815 ;
        RECT 89.255 109.770 89.545 109.815 ;
        RECT 90.175 109.955 90.465 110.000 ;
        RECT 92.920 109.955 93.240 110.015 ;
        RECT 90.175 109.815 93.240 109.955 ;
        RECT 90.175 109.770 90.465 109.815 ;
        RECT 92.920 109.755 93.240 109.815 ;
        RECT 96.600 109.955 96.920 110.015 ;
        RECT 98.915 109.955 99.205 110.000 ;
        RECT 96.600 109.815 99.205 109.955 ;
        RECT 96.600 109.755 96.920 109.815 ;
        RECT 98.915 109.770 99.205 109.815 ;
        RECT 105.355 109.955 105.645 110.000 ;
        RECT 105.800 109.955 106.120 110.015 ;
        RECT 105.355 109.815 106.120 109.955 ;
        RECT 105.355 109.770 105.645 109.815 ;
        RECT 105.800 109.755 106.120 109.815 ;
        RECT 14.275 109.475 15.960 109.615 ;
        RECT 14.275 109.430 14.565 109.475 ;
        RECT 15.640 109.415 15.960 109.475 ;
        RECT 13.800 109.275 14.120 109.335 ;
        RECT 17.435 109.320 17.725 109.635 ;
        RECT 18.515 109.615 18.805 109.660 ;
        RECT 22.095 109.615 22.385 109.660 ;
        RECT 23.930 109.615 24.220 109.660 ;
        RECT 18.515 109.475 24.220 109.615 ;
        RECT 18.515 109.430 18.805 109.475 ;
        RECT 22.095 109.430 22.385 109.475 ;
        RECT 23.930 109.430 24.220 109.475 ;
        RECT 25.775 109.430 26.065 109.660 ;
        RECT 27.155 109.615 27.445 109.660 ;
        RECT 29.900 109.615 30.220 109.675 ;
        RECT 27.155 109.475 30.220 109.615 ;
        RECT 27.155 109.430 27.445 109.475 ;
        RECT 29.900 109.415 30.220 109.475 ;
        RECT 17.135 109.275 17.725 109.320 ;
        RECT 20.375 109.275 21.025 109.320 ;
        RECT 13.800 109.135 21.025 109.275 ;
        RECT 13.800 109.075 14.120 109.135 ;
        RECT 17.135 109.090 17.425 109.135 ;
        RECT 20.375 109.090 21.025 109.135 ;
        RECT 23.015 109.090 23.305 109.320 ;
        RECT 23.460 109.275 23.780 109.335 ;
        RECT 23.460 109.135 26.450 109.275 ;
        RECT 23.090 108.935 23.230 109.090 ;
        RECT 23.460 109.075 23.780 109.135 ;
        RECT 26.310 108.980 26.450 109.135 ;
        RECT 27.615 109.090 27.905 109.320 ;
        RECT 28.980 109.275 29.300 109.335 ;
        RECT 30.775 109.320 31.065 109.635 ;
        RECT 31.855 109.615 32.145 109.660 ;
        RECT 35.435 109.615 35.725 109.660 ;
        RECT 37.270 109.615 37.560 109.660 ;
        RECT 31.855 109.475 37.560 109.615 ;
        RECT 31.855 109.430 32.145 109.475 ;
        RECT 35.435 109.430 35.725 109.475 ;
        RECT 37.270 109.430 37.560 109.475 ;
        RECT 40.495 109.430 40.785 109.660 ;
        RECT 40.940 109.615 41.260 109.675 ;
        RECT 42.335 109.615 42.625 109.660 ;
        RECT 40.940 109.475 42.625 109.615 ;
        RECT 30.475 109.275 31.065 109.320 ;
        RECT 33.715 109.275 34.365 109.320 ;
        RECT 28.980 109.135 34.365 109.275 ;
        RECT 40.570 109.275 40.710 109.430 ;
        RECT 40.940 109.415 41.260 109.475 ;
        RECT 42.335 109.430 42.625 109.475 ;
        RECT 44.620 109.415 44.940 109.675 ;
        RECT 49.220 109.635 49.540 109.675 ;
        RECT 49.175 109.415 49.540 109.635 ;
        RECT 50.255 109.615 50.545 109.660 ;
        RECT 53.835 109.615 54.125 109.660 ;
        RECT 55.670 109.615 55.960 109.660 ;
        RECT 50.255 109.475 55.960 109.615 ;
        RECT 50.255 109.430 50.545 109.475 ;
        RECT 53.835 109.430 54.125 109.475 ;
        RECT 55.670 109.430 55.960 109.475 ;
        RECT 56.580 109.615 56.900 109.675 ;
        RECT 57.055 109.615 57.345 109.660 ;
        RECT 58.435 109.615 58.725 109.660 ;
        RECT 56.580 109.475 57.345 109.615 ;
        RECT 56.580 109.415 56.900 109.475 ;
        RECT 57.055 109.430 57.345 109.475 ;
        RECT 57.590 109.475 58.725 109.615 ;
        RECT 46.000 109.275 46.320 109.335 ;
        RECT 49.175 109.320 49.465 109.415 ;
        RECT 40.570 109.135 46.320 109.275 ;
        RECT 24.855 108.935 25.145 108.980 ;
        RECT 23.090 108.795 25.145 108.935 ;
        RECT 24.855 108.750 25.145 108.795 ;
        RECT 26.235 108.750 26.525 108.980 ;
        RECT 27.690 108.935 27.830 109.090 ;
        RECT 28.980 109.075 29.300 109.135 ;
        RECT 30.475 109.090 30.765 109.135 ;
        RECT 33.715 109.090 34.365 109.135 ;
        RECT 46.000 109.075 46.320 109.135 ;
        RECT 48.875 109.275 49.465 109.320 ;
        RECT 52.115 109.275 52.765 109.320 ;
        RECT 48.875 109.135 52.765 109.275 ;
        RECT 48.875 109.090 49.165 109.135 ;
        RECT 52.115 109.090 52.765 109.135 ;
        RECT 32.200 108.935 32.520 108.995 ;
        RECT 27.690 108.795 32.520 108.935 ;
        RECT 32.200 108.735 32.520 108.795 ;
        RECT 40.020 108.735 40.340 108.995 ;
        RECT 45.555 108.935 45.845 108.980 ;
        RECT 47.840 108.935 48.160 108.995 ;
        RECT 45.555 108.795 48.160 108.935 ;
        RECT 45.555 108.750 45.845 108.795 ;
        RECT 47.840 108.735 48.160 108.795 ;
        RECT 51.520 108.935 51.840 108.995 ;
        RECT 57.590 108.935 57.730 109.475 ;
        RECT 58.435 109.430 58.725 109.475 ;
        RECT 60.260 109.615 60.580 109.675 ;
        RECT 61.195 109.615 61.485 109.660 ;
        RECT 60.260 109.475 61.485 109.615 ;
        RECT 60.260 109.415 60.580 109.475 ;
        RECT 61.195 109.430 61.485 109.475 ;
        RECT 63.940 109.615 64.260 109.675 ;
        RECT 64.875 109.615 65.165 109.660 ;
        RECT 63.940 109.475 65.165 109.615 ;
        RECT 63.940 109.415 64.260 109.475 ;
        RECT 64.875 109.430 65.165 109.475 ;
        RECT 67.160 109.415 67.480 109.675 ;
        RECT 67.635 109.430 67.925 109.660 ;
        RECT 68.100 109.615 68.390 109.660 ;
        RECT 69.935 109.615 70.225 109.660 ;
        RECT 73.515 109.615 73.805 109.660 ;
        RECT 68.100 109.475 73.805 109.615 ;
        RECT 68.100 109.430 68.390 109.475 ;
        RECT 69.935 109.430 70.225 109.475 ;
        RECT 73.515 109.430 73.805 109.475 ;
        RECT 74.520 109.635 74.840 109.675 ;
        RECT 51.520 108.795 57.730 108.935 ;
        RECT 51.520 108.735 51.840 108.795 ;
        RECT 57.960 108.735 58.280 108.995 ;
        RECT 58.880 108.735 59.200 108.995 ;
        RECT 62.100 108.735 62.420 108.995 ;
        RECT 67.710 108.935 67.850 109.430 ;
        RECT 74.520 109.415 74.885 109.635 ;
        RECT 74.595 109.320 74.885 109.415 ;
        RECT 82.295 109.320 82.585 109.635 ;
        RECT 83.375 109.615 83.665 109.660 ;
        RECT 86.955 109.615 87.245 109.660 ;
        RECT 88.790 109.615 89.080 109.660 ;
        RECT 83.375 109.475 89.080 109.615 ;
        RECT 83.375 109.430 83.665 109.475 ;
        RECT 86.955 109.430 87.245 109.475 ;
        RECT 88.790 109.430 89.080 109.475 ;
        RECT 71.295 109.275 71.945 109.320 ;
        RECT 74.595 109.275 75.185 109.320 ;
        RECT 71.295 109.135 75.185 109.275 ;
        RECT 71.295 109.090 71.945 109.135 ;
        RECT 74.895 109.090 75.185 109.135 ;
        RECT 81.995 109.275 82.585 109.320 ;
        RECT 84.180 109.275 84.500 109.335 ;
        RECT 93.335 109.320 93.625 109.635 ;
        RECT 94.415 109.615 94.705 109.660 ;
        RECT 97.995 109.615 98.285 109.660 ;
        RECT 99.830 109.615 100.120 109.660 ;
        RECT 94.415 109.475 100.120 109.615 ;
        RECT 94.415 109.430 94.705 109.475 ;
        RECT 97.995 109.430 98.285 109.475 ;
        RECT 99.830 109.430 100.120 109.475 ;
        RECT 100.295 109.615 100.585 109.660 ;
        RECT 100.740 109.615 101.060 109.675 ;
        RECT 101.660 109.615 101.980 109.675 ;
        RECT 103.960 109.615 104.280 109.675 ;
        RECT 100.295 109.475 104.280 109.615 ;
        RECT 100.295 109.430 100.585 109.475 ;
        RECT 100.740 109.415 101.060 109.475 ;
        RECT 101.660 109.415 101.980 109.475 ;
        RECT 103.960 109.415 104.280 109.475 ;
        RECT 104.440 109.615 104.730 109.660 ;
        RECT 106.275 109.615 106.565 109.660 ;
        RECT 109.855 109.615 110.145 109.660 ;
        RECT 104.440 109.475 110.145 109.615 ;
        RECT 104.440 109.430 104.730 109.475 ;
        RECT 106.275 109.430 106.565 109.475 ;
        RECT 109.855 109.430 110.145 109.475 ;
        RECT 85.235 109.275 85.885 109.320 ;
        RECT 81.995 109.135 85.885 109.275 ;
        RECT 81.995 109.090 82.285 109.135 ;
        RECT 84.180 109.075 84.500 109.135 ;
        RECT 85.235 109.090 85.885 109.135 ;
        RECT 93.035 109.275 93.625 109.320 ;
        RECT 96.275 109.275 96.925 109.320 ;
        RECT 98.900 109.275 99.220 109.335 ;
        RECT 93.035 109.135 99.220 109.275 ;
        RECT 93.035 109.090 93.325 109.135 ;
        RECT 96.275 109.090 96.925 109.135 ;
        RECT 98.900 109.075 99.220 109.135 ;
        RECT 107.635 109.275 108.285 109.320 ;
        RECT 108.560 109.275 108.880 109.335 ;
        RECT 110.935 109.320 111.225 109.635 ;
        RECT 110.935 109.275 111.525 109.320 ;
        RECT 107.635 109.135 111.525 109.275 ;
        RECT 107.635 109.090 108.285 109.135 ;
        RECT 108.560 109.075 108.880 109.135 ;
        RECT 111.235 109.090 111.525 109.135 ;
        RECT 114.095 109.090 114.385 109.320 ;
        RECT 73.600 108.935 73.920 108.995 ;
        RECT 67.710 108.795 73.920 108.935 ;
        RECT 73.600 108.735 73.920 108.795 ;
        RECT 109.480 108.935 109.800 108.995 ;
        RECT 114.170 108.935 114.310 109.090 ;
        RECT 109.480 108.795 114.310 108.935 ;
        RECT 109.480 108.735 109.800 108.795 ;
        RECT 10.510 108.115 115.850 108.595 ;
        RECT 13.800 107.715 14.120 107.975 ;
        RECT 17.110 107.775 26.910 107.915 ;
        RECT 12.895 107.235 13.185 107.280 ;
        RECT 13.355 107.235 13.645 107.280 ;
        RECT 17.110 107.235 17.250 107.775 ;
        RECT 21.160 107.620 21.480 107.635 ;
        RECT 17.595 107.575 17.885 107.620 ;
        RECT 20.835 107.575 21.485 107.620 ;
        RECT 17.595 107.435 21.485 107.575 ;
        RECT 17.595 107.390 18.185 107.435 ;
        RECT 20.835 107.390 21.485 107.435 ;
        RECT 12.895 107.095 17.250 107.235 ;
        RECT 12.895 107.050 13.185 107.095 ;
        RECT 13.355 107.050 13.645 107.095 ;
        RECT 17.895 107.075 18.185 107.390 ;
        RECT 21.160 107.375 21.480 107.390 ;
        RECT 23.460 107.375 23.780 107.635 ;
        RECT 26.770 107.280 26.910 107.775 ;
        RECT 28.980 107.715 29.300 107.975 ;
        RECT 46.000 107.915 46.320 107.975 ;
        RECT 59.340 107.915 59.660 107.975 ;
        RECT 29.530 107.775 46.320 107.915 ;
        RECT 18.975 107.235 19.265 107.280 ;
        RECT 22.555 107.235 22.845 107.280 ;
        RECT 24.390 107.235 24.680 107.280 ;
        RECT 18.975 107.095 24.680 107.235 ;
        RECT 18.975 107.050 19.265 107.095 ;
        RECT 22.555 107.050 22.845 107.095 ;
        RECT 24.390 107.050 24.680 107.095 ;
        RECT 26.695 107.235 26.985 107.280 ;
        RECT 27.155 107.235 27.445 107.280 ;
        RECT 28.535 107.235 28.825 107.280 ;
        RECT 29.530 107.235 29.670 107.775 ;
        RECT 46.000 107.715 46.320 107.775 ;
        RECT 50.690 107.775 62.330 107.915 ;
        RECT 31.295 107.575 31.585 107.620 ;
        RECT 32.660 107.575 32.980 107.635 ;
        RECT 31.295 107.435 32.980 107.575 ;
        RECT 31.295 107.390 31.585 107.435 ;
        RECT 32.660 107.375 32.980 107.435 ;
        RECT 33.575 107.575 34.225 107.620 ;
        RECT 37.175 107.575 37.465 107.620 ;
        RECT 40.020 107.575 40.340 107.635 ;
        RECT 33.575 107.435 40.340 107.575 ;
        RECT 33.575 107.390 34.225 107.435 ;
        RECT 36.875 107.390 37.465 107.435 ;
        RECT 26.695 107.095 29.670 107.235 ;
        RECT 30.380 107.235 30.670 107.280 ;
        RECT 32.215 107.235 32.505 107.280 ;
        RECT 35.795 107.235 36.085 107.280 ;
        RECT 30.380 107.095 36.085 107.235 ;
        RECT 26.695 107.050 26.985 107.095 ;
        RECT 27.155 107.050 27.445 107.095 ;
        RECT 28.535 107.050 28.825 107.095 ;
        RECT 30.380 107.050 30.670 107.095 ;
        RECT 32.215 107.050 32.505 107.095 ;
        RECT 35.795 107.050 36.085 107.095 ;
        RECT 36.875 107.075 37.165 107.390 ;
        RECT 40.020 107.375 40.340 107.435 ;
        RECT 43.355 107.575 43.645 107.620 ;
        RECT 44.160 107.575 44.480 107.635 ;
        RECT 46.595 107.575 47.245 107.620 ;
        RECT 43.355 107.435 47.245 107.575 ;
        RECT 43.355 107.390 43.945 107.435 ;
        RECT 43.655 107.075 43.945 107.390 ;
        RECT 44.160 107.375 44.480 107.435 ;
        RECT 46.595 107.390 47.245 107.435 ;
        RECT 47.840 107.575 48.160 107.635 ;
        RECT 49.235 107.575 49.525 107.620 ;
        RECT 47.840 107.435 49.525 107.575 ;
        RECT 47.840 107.375 48.160 107.435 ;
        RECT 49.235 107.390 49.525 107.435 ;
        RECT 50.690 107.280 50.830 107.775 ;
        RECT 59.340 107.715 59.660 107.775 ;
        RECT 52.440 107.575 52.760 107.635 ;
        RECT 54.855 107.575 55.145 107.620 ;
        RECT 58.095 107.575 58.745 107.620 ;
        RECT 52.440 107.435 58.745 107.575 ;
        RECT 52.440 107.375 52.760 107.435 ;
        RECT 54.855 107.390 55.445 107.435 ;
        RECT 58.095 107.390 58.745 107.435 ;
        RECT 44.735 107.235 45.025 107.280 ;
        RECT 48.315 107.235 48.605 107.280 ;
        RECT 50.150 107.235 50.440 107.280 ;
        RECT 44.735 107.095 50.440 107.235 ;
        RECT 44.735 107.050 45.025 107.095 ;
        RECT 48.315 107.050 48.605 107.095 ;
        RECT 50.150 107.050 50.440 107.095 ;
        RECT 50.615 107.050 50.905 107.280 ;
        RECT 55.155 107.075 55.445 107.390 ;
        RECT 62.190 107.280 62.330 107.775 ;
        RECT 74.520 107.715 74.840 107.975 ;
        RECT 98.900 107.715 99.220 107.975 ;
        RECT 100.740 107.715 101.060 107.975 ;
        RECT 63.495 107.575 63.785 107.620 ;
        RECT 64.400 107.575 64.720 107.635 ;
        RECT 69.920 107.620 70.240 107.635 ;
        RECT 63.495 107.435 64.720 107.575 ;
        RECT 63.495 107.390 63.785 107.435 ;
        RECT 64.400 107.375 64.720 107.435 ;
        RECT 66.355 107.575 66.645 107.620 ;
        RECT 69.595 107.575 70.245 107.620 ;
        RECT 66.355 107.435 70.245 107.575 ;
        RECT 66.355 107.390 66.945 107.435 ;
        RECT 69.595 107.390 70.245 107.435 ;
        RECT 56.235 107.235 56.525 107.280 ;
        RECT 59.815 107.235 60.105 107.280 ;
        RECT 61.650 107.235 61.940 107.280 ;
        RECT 56.235 107.095 61.940 107.235 ;
        RECT 56.235 107.050 56.525 107.095 ;
        RECT 59.815 107.050 60.105 107.095 ;
        RECT 61.650 107.050 61.940 107.095 ;
        RECT 62.115 107.235 62.405 107.280 ;
        RECT 62.115 107.095 63.710 107.235 ;
        RECT 62.115 107.050 62.405 107.095 ;
        RECT 63.570 106.955 63.710 107.095 ;
        RECT 66.655 107.075 66.945 107.390 ;
        RECT 69.920 107.375 70.240 107.390 ;
        RECT 72.220 107.375 72.540 107.635 ;
        RECT 72.680 107.575 73.000 107.635 ;
        RECT 75.915 107.575 76.205 107.620 ;
        RECT 80.155 107.575 80.445 107.620 ;
        RECT 83.395 107.575 84.045 107.620 ;
        RECT 72.680 107.435 75.210 107.575 ;
        RECT 72.680 107.375 73.000 107.435 ;
        RECT 67.735 107.235 68.025 107.280 ;
        RECT 71.315 107.235 71.605 107.280 ;
        RECT 73.150 107.235 73.440 107.280 ;
        RECT 67.735 107.095 73.440 107.235 ;
        RECT 67.735 107.050 68.025 107.095 ;
        RECT 71.315 107.050 71.605 107.095 ;
        RECT 73.150 107.050 73.440 107.095 ;
        RECT 73.600 107.035 73.920 107.295 ;
        RECT 75.070 107.280 75.210 107.435 ;
        RECT 75.915 107.435 84.045 107.575 ;
        RECT 75.915 107.390 76.205 107.435 ;
        RECT 80.155 107.390 80.745 107.435 ;
        RECT 83.395 107.390 84.045 107.435 ;
        RECT 88.780 107.575 89.100 107.635 ;
        RECT 90.735 107.575 91.025 107.620 ;
        RECT 93.975 107.575 94.625 107.620 ;
        RECT 100.830 107.575 100.970 107.715 ;
        RECT 88.780 107.435 94.625 107.575 ;
        RECT 74.995 107.235 75.285 107.280 ;
        RECT 75.440 107.235 75.760 107.295 ;
        RECT 74.995 107.095 75.760 107.235 ;
        RECT 74.995 107.050 75.285 107.095 ;
        RECT 75.440 107.035 75.760 107.095 ;
        RECT 80.455 107.075 80.745 107.390 ;
        RECT 88.780 107.375 89.100 107.435 ;
        RECT 90.735 107.390 91.325 107.435 ;
        RECT 93.975 107.390 94.625 107.435 ;
        RECT 98.070 107.435 100.970 107.575 ;
        RECT 101.675 107.575 101.965 107.620 ;
        RECT 105.915 107.575 106.205 107.620 ;
        RECT 109.155 107.575 109.805 107.620 ;
        RECT 101.675 107.435 109.805 107.575 ;
        RECT 81.535 107.235 81.825 107.280 ;
        RECT 85.115 107.235 85.405 107.280 ;
        RECT 86.950 107.235 87.240 107.280 ;
        RECT 81.535 107.095 87.240 107.235 ;
        RECT 81.535 107.050 81.825 107.095 ;
        RECT 85.115 107.050 85.405 107.095 ;
        RECT 86.950 107.050 87.240 107.095 ;
        RECT 87.400 107.035 87.720 107.295 ;
        RECT 91.035 107.075 91.325 107.390 ;
        RECT 98.070 107.280 98.210 107.435 ;
        RECT 101.675 107.390 101.965 107.435 ;
        RECT 105.915 107.390 106.505 107.435 ;
        RECT 109.155 107.390 109.805 107.435 ;
        RECT 92.115 107.235 92.405 107.280 ;
        RECT 95.695 107.235 95.985 107.280 ;
        RECT 97.530 107.235 97.820 107.280 ;
        RECT 92.115 107.095 97.820 107.235 ;
        RECT 92.115 107.050 92.405 107.095 ;
        RECT 95.695 107.050 95.985 107.095 ;
        RECT 97.530 107.050 97.820 107.095 ;
        RECT 97.995 107.050 98.285 107.280 ;
        RECT 98.440 107.235 98.760 107.295 ;
        RECT 99.375 107.235 99.665 107.280 ;
        RECT 100.755 107.235 101.045 107.280 ;
        RECT 101.215 107.235 101.505 107.280 ;
        RECT 98.440 107.095 105.110 107.235 ;
        RECT 98.440 107.035 98.760 107.095 ;
        RECT 99.375 107.050 99.665 107.095 ;
        RECT 100.755 107.050 101.045 107.095 ;
        RECT 101.215 107.050 101.505 107.095 ;
        RECT 12.435 106.895 12.725 106.940 ;
        RECT 13.800 106.895 14.120 106.955 ;
        RECT 12.435 106.755 14.120 106.895 ;
        RECT 12.435 106.710 12.725 106.755 ;
        RECT 13.800 106.695 14.120 106.755 ;
        RECT 14.735 106.895 15.025 106.940 ;
        RECT 23.000 106.895 23.320 106.955 ;
        RECT 14.735 106.755 23.320 106.895 ;
        RECT 14.735 106.710 15.025 106.755 ;
        RECT 23.000 106.695 23.320 106.755 ;
        RECT 24.840 106.695 25.160 106.955 ;
        RECT 27.600 106.695 27.920 106.955 ;
        RECT 29.915 106.895 30.205 106.940 ;
        RECT 36.340 106.895 36.660 106.955 ;
        RECT 29.915 106.755 36.660 106.895 ;
        RECT 29.915 106.710 30.205 106.755 ;
        RECT 36.340 106.695 36.660 106.755 ;
        RECT 38.180 106.895 38.500 106.955 ;
        RECT 40.035 106.895 40.325 106.940 ;
        RECT 38.180 106.755 40.325 106.895 ;
        RECT 38.180 106.695 38.500 106.755 ;
        RECT 40.035 106.710 40.325 106.755 ;
        RECT 40.495 106.895 40.785 106.940 ;
        RECT 43.240 106.895 43.560 106.955 ;
        RECT 40.495 106.755 43.560 106.895 ;
        RECT 40.495 106.710 40.785 106.755 ;
        RECT 43.240 106.695 43.560 106.755 ;
        RECT 51.995 106.895 52.285 106.940 ;
        RECT 54.740 106.895 55.060 106.955 ;
        RECT 51.995 106.755 55.060 106.895 ;
        RECT 51.995 106.710 52.285 106.755 ;
        RECT 54.740 106.695 55.060 106.755 ;
        RECT 57.960 106.895 58.280 106.955 ;
        RECT 60.735 106.895 61.025 106.940 ;
        RECT 57.960 106.755 61.025 106.895 ;
        RECT 57.960 106.695 58.280 106.755 ;
        RECT 60.735 106.710 61.025 106.755 ;
        RECT 63.480 106.695 63.800 106.955 ;
        RECT 76.820 106.895 77.140 106.955 ;
        RECT 77.295 106.895 77.585 106.940 ;
        RECT 76.820 106.755 77.585 106.895 ;
        RECT 76.820 106.695 77.140 106.755 ;
        RECT 77.295 106.710 77.585 106.755 ;
        RECT 87.860 106.695 88.180 106.955 ;
        RECT 100.280 106.695 100.600 106.955 ;
        RECT 103.055 106.895 103.345 106.940 ;
        RECT 104.420 106.895 104.740 106.955 ;
        RECT 103.055 106.755 104.740 106.895 ;
        RECT 104.970 106.895 105.110 107.095 ;
        RECT 106.215 107.075 106.505 107.390 ;
        RECT 107.295 107.235 107.585 107.280 ;
        RECT 110.875 107.235 111.165 107.280 ;
        RECT 112.710 107.235 113.000 107.280 ;
        RECT 107.295 107.095 113.000 107.235 ;
        RECT 107.295 107.050 107.585 107.095 ;
        RECT 110.875 107.050 111.165 107.095 ;
        RECT 112.710 107.050 113.000 107.095 ;
        RECT 108.100 106.895 108.420 106.955 ;
        RECT 104.970 106.755 108.420 106.895 ;
        RECT 103.055 106.710 103.345 106.755 ;
        RECT 104.420 106.695 104.740 106.755 ;
        RECT 108.100 106.695 108.420 106.755 ;
        RECT 109.020 106.895 109.340 106.955 ;
        RECT 113.175 106.895 113.465 106.940 ;
        RECT 109.020 106.755 113.465 106.895 ;
        RECT 109.020 106.695 109.340 106.755 ;
        RECT 113.175 106.710 113.465 106.755 ;
        RECT 135.660 106.690 136.800 133.400 ;
        RECT 133.100 106.600 136.850 106.690 ;
        RECT 18.975 106.555 19.265 106.600 ;
        RECT 22.095 106.555 22.385 106.600 ;
        RECT 23.985 106.555 24.275 106.600 ;
        RECT 18.975 106.415 24.275 106.555 ;
        RECT 18.975 106.370 19.265 106.415 ;
        RECT 22.095 106.370 22.385 106.415 ;
        RECT 23.985 106.370 24.275 106.415 ;
        RECT 30.785 106.555 31.075 106.600 ;
        RECT 32.675 106.555 32.965 106.600 ;
        RECT 35.795 106.555 36.085 106.600 ;
        RECT 30.785 106.415 36.085 106.555 ;
        RECT 30.785 106.370 31.075 106.415 ;
        RECT 32.675 106.370 32.965 106.415 ;
        RECT 35.795 106.370 36.085 106.415 ;
        RECT 44.735 106.555 45.025 106.600 ;
        RECT 47.855 106.555 48.145 106.600 ;
        RECT 49.745 106.555 50.035 106.600 ;
        RECT 44.735 106.415 50.035 106.555 ;
        RECT 44.735 106.370 45.025 106.415 ;
        RECT 47.855 106.370 48.145 106.415 ;
        RECT 49.745 106.370 50.035 106.415 ;
        RECT 56.235 106.555 56.525 106.600 ;
        RECT 59.355 106.555 59.645 106.600 ;
        RECT 61.245 106.555 61.535 106.600 ;
        RECT 56.235 106.415 61.535 106.555 ;
        RECT 56.235 106.370 56.525 106.415 ;
        RECT 59.355 106.370 59.645 106.415 ;
        RECT 61.245 106.370 61.535 106.415 ;
        RECT 67.735 106.555 68.025 106.600 ;
        RECT 70.855 106.555 71.145 106.600 ;
        RECT 72.745 106.555 73.035 106.600 ;
        RECT 67.735 106.415 73.035 106.555 ;
        RECT 67.735 106.370 68.025 106.415 ;
        RECT 70.855 106.370 71.145 106.415 ;
        RECT 72.745 106.370 73.035 106.415 ;
        RECT 81.535 106.555 81.825 106.600 ;
        RECT 84.655 106.555 84.945 106.600 ;
        RECT 86.545 106.555 86.835 106.600 ;
        RECT 81.535 106.415 86.835 106.555 ;
        RECT 81.535 106.370 81.825 106.415 ;
        RECT 84.655 106.370 84.945 106.415 ;
        RECT 86.545 106.370 86.835 106.415 ;
        RECT 92.115 106.555 92.405 106.600 ;
        RECT 95.235 106.555 95.525 106.600 ;
        RECT 97.125 106.555 97.415 106.600 ;
        RECT 92.115 106.415 97.415 106.555 ;
        RECT 92.115 106.370 92.405 106.415 ;
        RECT 95.235 106.370 95.525 106.415 ;
        RECT 97.125 106.370 97.415 106.415 ;
        RECT 107.295 106.555 107.585 106.600 ;
        RECT 110.415 106.555 110.705 106.600 ;
        RECT 112.305 106.555 112.595 106.600 ;
        RECT 107.295 106.415 112.595 106.555 ;
        RECT 107.295 106.370 107.585 106.415 ;
        RECT 110.415 106.370 110.705 106.415 ;
        RECT 112.305 106.370 112.595 106.415 ;
        RECT 21.160 106.215 21.480 106.275 ;
        RECT 26.235 106.215 26.525 106.260 ;
        RECT 21.160 106.075 26.525 106.215 ;
        RECT 21.160 106.015 21.480 106.075 ;
        RECT 26.235 106.030 26.525 106.075 ;
        RECT 71.760 106.215 72.080 106.275 ;
        RECT 86.100 106.215 86.390 106.260 ;
        RECT 71.760 106.075 86.390 106.215 ;
        RECT 71.760 106.015 72.080 106.075 ;
        RECT 86.100 106.030 86.390 106.075 ;
        RECT 91.080 106.215 91.400 106.275 ;
        RECT 96.680 106.215 96.970 106.260 ;
        RECT 91.080 106.075 96.970 106.215 ;
        RECT 91.080 106.015 91.400 106.075 ;
        RECT 96.680 106.030 96.970 106.075 ;
        RECT 103.500 106.215 103.820 106.275 ;
        RECT 111.860 106.215 112.150 106.260 ;
        RECT 103.500 106.075 112.150 106.215 ;
        RECT 103.500 106.015 103.820 106.075 ;
        RECT 111.860 106.030 112.150 106.075 ;
        RECT 10.510 105.395 115.850 105.875 ;
        RECT 129.700 105.630 136.850 106.600 ;
        RECT 133.100 105.500 136.850 105.630 ;
        RECT 44.160 105.195 44.480 105.255 ;
        RECT 45.555 105.195 45.845 105.240 ;
        RECT 44.160 105.055 45.845 105.195 ;
        RECT 44.160 104.995 44.480 105.055 ;
        RECT 45.555 105.010 45.845 105.055 ;
        RECT 49.220 105.195 49.540 105.255 ;
        RECT 50.155 105.195 50.445 105.240 ;
        RECT 49.220 105.055 50.445 105.195 ;
        RECT 49.220 104.995 49.540 105.055 ;
        RECT 50.155 105.010 50.445 105.055 ;
        RECT 52.440 104.995 52.760 105.255 ;
        RECT 69.920 105.195 70.240 105.255 ;
        RECT 70.395 105.195 70.685 105.240 ;
        RECT 69.920 105.055 70.685 105.195 ;
        RECT 69.920 104.995 70.240 105.055 ;
        RECT 70.395 105.010 70.685 105.055 ;
        RECT 84.180 104.995 84.500 105.255 ;
        RECT 88.780 104.995 89.100 105.255 ;
        RECT 98.440 105.195 98.760 105.255 ;
        RECT 91.630 105.055 98.760 105.195 ;
        RECT 17.135 104.855 17.425 104.900 ;
        RECT 20.255 104.855 20.545 104.900 ;
        RECT 22.145 104.855 22.435 104.900 ;
        RECT 17.135 104.715 22.435 104.855 ;
        RECT 17.135 104.670 17.425 104.715 ;
        RECT 20.255 104.670 20.545 104.715 ;
        RECT 22.145 104.670 22.435 104.715 ;
        RECT 30.015 104.855 30.305 104.900 ;
        RECT 33.135 104.855 33.425 104.900 ;
        RECT 35.025 104.855 35.315 104.900 ;
        RECT 30.015 104.715 35.315 104.855 ;
        RECT 30.015 104.670 30.305 104.715 ;
        RECT 33.135 104.670 33.425 104.715 ;
        RECT 35.025 104.670 35.315 104.715 ;
        RECT 57.615 104.855 57.905 104.900 ;
        RECT 60.735 104.855 61.025 104.900 ;
        RECT 62.625 104.855 62.915 104.900 ;
        RECT 57.615 104.715 62.915 104.855 ;
        RECT 57.615 104.670 57.905 104.715 ;
        RECT 60.735 104.670 61.025 104.715 ;
        RECT 62.625 104.670 62.915 104.715 ;
        RECT 23.015 104.515 23.305 104.560 ;
        RECT 24.380 104.515 24.700 104.575 ;
        RECT 23.015 104.375 24.700 104.515 ;
        RECT 23.015 104.330 23.305 104.375 ;
        RECT 24.380 104.315 24.700 104.375 ;
        RECT 34.500 104.315 34.820 104.575 ;
        RECT 35.895 104.515 36.185 104.560 ;
        RECT 36.340 104.515 36.660 104.575 ;
        RECT 35.895 104.375 36.660 104.515 ;
        RECT 35.895 104.330 36.185 104.375 ;
        RECT 36.340 104.315 36.660 104.375 ;
        RECT 53.375 104.515 53.665 104.560 ;
        RECT 60.260 104.515 60.580 104.575 ;
        RECT 53.375 104.375 60.580 104.515 ;
        RECT 53.375 104.330 53.665 104.375 ;
        RECT 60.260 104.315 60.580 104.375 ;
        RECT 62.100 104.315 62.420 104.575 ;
        RECT 63.480 104.315 63.800 104.575 ;
        RECT 10.580 103.835 10.900 103.895 ;
        RECT 12.895 103.835 13.185 103.880 ;
        RECT 10.580 103.695 13.185 103.835 ;
        RECT 10.580 103.635 10.900 103.695 ;
        RECT 12.895 103.650 13.185 103.695 ;
        RECT 13.800 103.835 14.120 103.895 ;
        RECT 16.055 103.880 16.345 104.195 ;
        RECT 17.135 104.175 17.425 104.220 ;
        RECT 20.715 104.175 21.005 104.220 ;
        RECT 22.550 104.175 22.840 104.220 ;
        RECT 17.135 104.035 22.840 104.175 ;
        RECT 17.135 103.990 17.425 104.035 ;
        RECT 20.715 103.990 21.005 104.035 ;
        RECT 22.550 103.990 22.840 104.035 ;
        RECT 15.755 103.835 16.345 103.880 ;
        RECT 18.995 103.835 19.645 103.880 ;
        RECT 13.800 103.695 19.645 103.835 ;
        RECT 13.800 103.635 14.120 103.695 ;
        RECT 15.755 103.650 16.045 103.695 ;
        RECT 18.995 103.650 19.645 103.695 ;
        RECT 21.635 103.835 21.925 103.880 ;
        RECT 22.080 103.835 22.400 103.895 ;
        RECT 21.635 103.695 22.400 103.835 ;
        RECT 21.635 103.650 21.925 103.695 ;
        RECT 22.080 103.635 22.400 103.695 ;
        RECT 25.775 103.835 26.065 103.880 ;
        RECT 27.140 103.835 27.460 103.895 ;
        RECT 25.775 103.695 27.460 103.835 ;
        RECT 25.775 103.650 26.065 103.695 ;
        RECT 27.140 103.635 27.460 103.695 ;
        RECT 27.600 103.835 27.920 103.895 ;
        RECT 28.935 103.880 29.225 104.195 ;
        RECT 30.015 104.175 30.305 104.220 ;
        RECT 33.595 104.175 33.885 104.220 ;
        RECT 35.430 104.175 35.720 104.220 ;
        RECT 30.015 104.035 35.720 104.175 ;
        RECT 30.015 103.990 30.305 104.035 ;
        RECT 33.595 103.990 33.885 104.035 ;
        RECT 35.430 103.990 35.720 104.035 ;
        RECT 46.000 104.175 46.320 104.235 ;
        RECT 49.695 104.175 49.985 104.220 ;
        RECT 51.980 104.175 52.300 104.235 ;
        RECT 46.000 104.035 52.300 104.175 ;
        RECT 46.000 103.975 46.320 104.035 ;
        RECT 49.695 103.990 49.985 104.035 ;
        RECT 51.980 103.975 52.300 104.035 ;
        RECT 56.535 103.880 56.825 104.195 ;
        RECT 57.615 104.175 57.905 104.220 ;
        RECT 61.195 104.175 61.485 104.220 ;
        RECT 63.030 104.175 63.320 104.220 ;
        RECT 57.615 104.035 63.320 104.175 ;
        RECT 57.615 103.990 57.905 104.035 ;
        RECT 61.195 103.990 61.485 104.035 ;
        RECT 63.030 103.990 63.320 104.035 ;
        RECT 70.855 104.175 71.145 104.220 ;
        RECT 75.440 104.175 75.760 104.235 ;
        RECT 84.655 104.175 84.945 104.220 ;
        RECT 88.335 104.175 88.625 104.220 ;
        RECT 91.630 104.175 91.770 105.055 ;
        RECT 98.440 104.995 98.760 105.055 ;
        RECT 108.560 104.995 108.880 105.255 ;
        RECT 96.255 104.855 96.545 104.900 ;
        RECT 99.375 104.855 99.665 104.900 ;
        RECT 101.265 104.855 101.555 104.900 ;
        RECT 96.255 104.715 101.555 104.855 ;
        RECT 96.255 104.670 96.545 104.715 ;
        RECT 99.375 104.670 99.665 104.715 ;
        RECT 101.265 104.670 101.555 104.715 ;
        RECT 92.015 104.515 92.305 104.560 ;
        RECT 98.900 104.515 99.220 104.575 ;
        RECT 92.015 104.375 99.220 104.515 ;
        RECT 92.015 104.330 92.305 104.375 ;
        RECT 98.900 104.315 99.220 104.375 ;
        RECT 100.740 104.315 101.060 104.575 ;
        RECT 102.120 104.315 102.440 104.575 ;
        RECT 70.855 104.035 91.770 104.175 ;
        RECT 70.855 103.990 71.145 104.035 ;
        RECT 75.440 103.975 75.760 104.035 ;
        RECT 84.655 103.990 84.945 104.035 ;
        RECT 88.335 103.990 88.625 104.035 ;
        RECT 28.635 103.835 29.225 103.880 ;
        RECT 31.875 103.835 32.525 103.880 ;
        RECT 27.600 103.695 32.525 103.835 ;
        RECT 27.600 103.635 27.920 103.695 ;
        RECT 28.635 103.650 28.925 103.695 ;
        RECT 31.875 103.650 32.525 103.695 ;
        RECT 56.235 103.835 56.825 103.880 ;
        RECT 58.880 103.835 59.200 103.895 ;
        RECT 95.175 103.880 95.465 104.195 ;
        RECT 96.255 104.175 96.545 104.220 ;
        RECT 99.835 104.175 100.125 104.220 ;
        RECT 101.670 104.175 101.960 104.220 ;
        RECT 96.255 104.035 101.960 104.175 ;
        RECT 96.255 103.990 96.545 104.035 ;
        RECT 99.835 103.990 100.125 104.035 ;
        RECT 101.670 103.990 101.960 104.035 ;
        RECT 108.100 103.975 108.420 104.235 ;
        RECT 114.095 104.175 114.385 104.220 ;
        RECT 119.140 104.175 119.460 104.235 ;
        RECT 114.095 104.035 119.460 104.175 ;
        RECT 114.095 103.990 114.385 104.035 ;
        RECT 119.140 103.975 119.460 104.035 ;
        RECT 59.475 103.835 60.125 103.880 ;
        RECT 56.235 103.695 60.125 103.835 ;
        RECT 56.235 103.650 56.525 103.695 ;
        RECT 58.880 103.635 59.200 103.695 ;
        RECT 59.475 103.650 60.125 103.695 ;
        RECT 94.875 103.835 95.465 103.880 ;
        RECT 98.115 103.835 98.765 103.880 ;
        RECT 100.280 103.835 100.600 103.895 ;
        RECT 94.875 103.695 100.600 103.835 ;
        RECT 94.875 103.650 95.165 103.695 ;
        RECT 98.115 103.650 98.765 103.695 ;
        RECT 100.280 103.635 100.600 103.695 ;
        RECT 113.160 103.295 113.480 103.555 ;
        RECT 10.510 102.675 115.850 103.155 ;
        RECT 67.160 102.475 67.480 102.535 ;
        RECT 113.160 102.475 113.480 102.535 ;
        RECT 67.160 102.335 113.480 102.475 ;
        RECT 67.160 102.275 67.480 102.335 ;
        RECT 113.160 102.275 113.480 102.335 ;
        RECT 133.330 76.630 136.060 77.830 ;
        RECT 137.920 77.810 143.450 77.960 ;
        RECT 21.115 74.380 23.065 74.390 ;
        RECT 19.415 73.240 23.065 74.380 ;
        RECT 19.415 73.230 21.125 73.240 ;
        RECT 28.135 73.230 30.305 74.410 ;
        RECT 32.315 74.390 34.265 74.400 ;
        RECT 30.615 73.250 34.265 74.390 ;
        RECT 30.615 73.240 32.325 73.250 ;
        RECT 39.425 73.200 41.595 74.380 ;
        RECT 43.535 74.360 45.485 74.370 ;
        RECT 41.835 73.220 45.485 74.360 ;
        RECT 54.785 74.340 56.735 74.350 ;
        RECT 41.835 73.210 43.545 73.220 ;
        RECT 3.910 73.080 6.100 73.190 ;
        RECT 50.005 73.140 52.175 74.320 ;
        RECT 53.085 73.200 56.735 74.340 ;
        RECT 53.085 73.190 54.795 73.200 ;
        RECT 61.425 73.170 63.595 74.350 ;
        RECT 66.005 74.330 67.955 74.340 ;
        RECT 64.305 73.190 67.955 74.330 ;
        RECT 64.305 73.180 66.015 73.190 ;
        RECT 72.535 73.180 74.705 74.360 ;
        RECT 77.245 74.320 79.195 74.330 ;
        RECT 75.545 73.180 79.195 74.320 ;
        RECT 75.545 73.170 77.255 73.180 ;
        RECT 83.805 73.170 85.975 74.350 ;
        RECT 88.495 74.330 90.445 74.340 ;
        RECT 86.795 73.190 90.445 74.330 ;
        RECT 99.775 74.320 101.725 74.330 ;
        RECT 86.795 73.180 88.505 73.190 ;
        RECT 94.995 73.110 97.165 74.290 ;
        RECT 98.075 73.180 101.725 74.320 ;
        RECT 98.075 73.170 99.785 73.180 ;
        RECT 106.405 73.160 108.575 74.340 ;
        RECT 111.045 74.320 112.995 74.330 ;
        RECT 109.345 73.180 112.995 74.320 ;
        RECT 109.345 73.170 111.055 73.180 ;
        RECT 117.605 73.160 119.775 74.340 ;
        RECT 122.295 74.320 124.245 74.330 ;
        RECT 120.595 73.180 124.245 74.320 ;
        RECT 129.455 73.240 131.625 74.420 ;
        RECT 120.595 73.170 122.305 73.180 ;
        RECT 3.910 72.820 12.240 73.080 ;
        RECT 29.635 72.840 43.235 72.850 ;
        RECT 18.435 72.820 43.235 72.840 ;
        RECT 3.910 72.800 54.455 72.820 ;
        RECT 3.910 72.790 65.705 72.800 ;
        RECT 133.960 72.790 135.640 76.630 ;
        RECT 137.190 76.610 143.450 77.810 ;
        RECT 137.920 75.460 143.450 76.610 ;
        RECT 3.910 72.780 76.925 72.790 ;
        RECT 85.815 72.780 99.415 72.790 ;
        RECT 132.085 72.780 140.600 72.790 ;
        RECT 3.910 71.700 140.600 72.780 ;
        RECT 3.910 71.690 32.035 71.700 ;
        RECT 3.910 71.670 19.135 71.690 ;
        RECT 40.855 71.670 140.600 71.700 ;
        RECT 3.910 71.500 12.240 71.670 ;
        RECT 52.105 71.650 140.600 71.670 ;
        RECT 63.325 71.640 140.600 71.650 ;
        RECT 74.565 71.630 88.165 71.640 ;
        RECT 97.095 71.630 133.215 71.640 ;
        RECT 3.910 71.370 6.100 71.500 ;
        RECT 10.800 71.180 11.950 71.500 ;
        RECT 10.800 69.480 11.915 71.180 ;
        RECT 29.635 71.170 43.285 71.180 ;
        RECT 15.510 71.155 17.040 71.160 ;
        RECT 18.435 71.155 43.285 71.170 ;
        RECT 12.285 71.150 43.285 71.155 ;
        RECT 12.285 71.130 54.505 71.150 ;
        RECT 141.810 71.140 143.230 75.460 ;
        RECT 12.285 71.120 65.755 71.130 ;
        RECT 12.285 71.110 76.975 71.120 ;
        RECT 85.815 71.110 99.465 71.120 ;
        RECT 140.220 71.110 143.240 71.140 ;
        RECT 12.285 70.030 143.240 71.110 ;
        RECT 12.285 70.020 32.085 70.030 ;
        RECT 12.285 70.005 19.375 70.020 ;
        RECT 10.800 13.800 11.950 69.480 ;
        RECT 12.320 15.450 13.470 70.005 ;
        RECT 15.510 68.660 17.040 70.005 ;
        RECT 40.855 70.000 143.240 70.030 ;
        RECT 52.105 69.980 143.240 70.000 ;
        RECT 63.325 69.970 143.240 69.980 ;
        RECT 74.565 69.960 88.215 69.970 ;
        RECT 97.095 69.960 143.240 69.970 ;
        RECT 140.220 69.910 143.240 69.960 ;
        RECT 29.645 69.670 43.315 69.680 ;
        RECT 18.445 69.650 43.315 69.670 ;
        RECT 18.445 69.630 54.535 69.650 ;
        RECT 18.445 69.620 65.785 69.630 ;
        RECT 139.590 69.620 150.610 69.640 ;
        RECT 18.445 69.610 77.005 69.620 ;
        RECT 85.825 69.610 99.495 69.620 ;
        RECT 132.155 69.610 150.610 69.620 ;
        RECT 18.445 69.570 150.610 69.610 ;
        RECT 18.445 68.530 150.740 69.570 ;
        RECT 18.445 68.520 32.115 68.530 ;
        RECT 40.865 68.500 150.740 68.530 ;
        RECT 52.115 68.490 143.320 68.500 ;
        RECT 52.115 68.480 140.670 68.490 ;
        RECT 63.335 68.470 140.670 68.480 ;
        RECT 74.575 68.460 88.245 68.470 ;
        RECT 97.105 68.460 133.295 68.470 ;
        RECT 141.080 68.450 142.300 68.490 ;
        RECT 149.360 68.470 150.740 68.500 ;
        RECT 29.655 68.100 43.325 68.110 ;
        RECT 13.950 68.080 43.325 68.100 ;
        RECT 13.950 68.060 54.545 68.080 ;
        RECT 13.950 68.050 65.795 68.060 ;
        RECT 13.950 68.040 77.015 68.050 ;
        RECT 85.835 68.040 99.505 68.050 ;
        RECT 139.530 68.040 143.320 68.060 ;
        RECT 13.950 66.960 152.870 68.040 ;
        RECT 13.950 66.950 32.125 66.960 ;
        RECT 13.950 18.530 15.100 66.950 ;
        RECT 40.875 66.930 152.870 66.960 ;
        RECT 52.125 66.910 152.870 66.930 ;
        RECT 63.345 66.900 152.870 66.910 ;
        RECT 74.585 66.890 88.255 66.900 ;
        RECT 97.115 66.890 143.320 66.900 ;
        RECT 141.030 66.770 142.490 66.890 ;
        RECT 21.405 65.510 26.555 65.790 ;
        RECT 27.815 65.490 28.965 65.800 ;
        RECT 32.605 65.520 37.755 65.800 ;
        RECT 39.015 65.500 40.165 65.810 ;
        RECT 43.825 65.490 48.975 65.770 ;
        RECT 50.235 65.470 51.385 65.780 ;
        RECT 149.460 65.760 150.600 65.780 ;
        RECT 55.075 65.470 60.225 65.750 ;
        RECT 61.485 65.450 62.635 65.760 ;
        RECT 66.295 65.460 71.445 65.740 ;
        RECT 72.705 65.440 73.855 65.750 ;
        RECT 77.535 65.450 82.685 65.730 ;
        RECT 83.945 65.430 85.095 65.740 ;
        RECT 88.785 65.460 93.935 65.740 ;
        RECT 95.195 65.440 96.345 65.750 ;
        RECT 100.065 65.450 105.215 65.730 ;
        RECT 106.475 65.430 107.625 65.740 ;
        RECT 111.335 65.450 116.485 65.730 ;
        RECT 117.745 65.430 118.895 65.740 ;
        RECT 122.585 65.450 127.735 65.730 ;
        RECT 128.995 65.430 130.145 65.740 ;
        RECT 133.315 65.430 138.455 65.690 ;
        RECT 21.205 65.140 21.435 65.320 ;
        RECT 26.495 65.190 26.725 65.320 ;
        RECT 21.125 55.220 21.485 65.140 ;
        RECT 26.435 55.240 26.805 65.190 ;
        RECT 27.635 65.150 27.865 65.320 ;
        RECT 27.565 55.200 27.935 65.150 ;
        RECT 28.925 65.140 29.155 65.320 ;
        RECT 32.405 65.150 32.635 65.330 ;
        RECT 37.695 65.200 37.925 65.330 ;
        RECT 28.835 55.250 29.255 65.140 ;
        RECT 32.325 55.230 32.685 65.150 ;
        RECT 37.635 55.250 38.005 65.200 ;
        RECT 38.835 65.160 39.065 65.330 ;
        RECT 38.765 55.210 39.135 65.160 ;
        RECT 40.125 65.150 40.355 65.330 ;
        RECT 40.035 55.260 40.455 65.150 ;
        RECT 43.625 65.120 43.855 65.300 ;
        RECT 48.915 65.170 49.145 65.300 ;
        RECT 43.545 55.200 43.905 65.120 ;
        RECT 48.855 55.220 49.225 65.170 ;
        RECT 50.055 65.130 50.285 65.300 ;
        RECT 49.985 55.180 50.355 65.130 ;
        RECT 51.345 65.120 51.575 65.300 ;
        RECT 51.255 55.230 51.675 65.120 ;
        RECT 54.875 65.100 55.105 65.280 ;
        RECT 60.165 65.150 60.395 65.280 ;
        RECT 54.795 55.180 55.155 65.100 ;
        RECT 60.105 55.200 60.475 65.150 ;
        RECT 61.305 65.110 61.535 65.280 ;
        RECT 61.235 55.160 61.605 65.110 ;
        RECT 62.595 65.100 62.825 65.280 ;
        RECT 62.505 55.210 62.925 65.100 ;
        RECT 66.095 65.090 66.325 65.270 ;
        RECT 71.385 65.140 71.615 65.270 ;
        RECT 66.015 55.170 66.375 65.090 ;
        RECT 71.325 55.190 71.695 65.140 ;
        RECT 72.525 65.100 72.755 65.270 ;
        RECT 72.455 55.150 72.825 65.100 ;
        RECT 73.815 65.090 74.045 65.270 ;
        RECT 73.725 55.200 74.145 65.090 ;
        RECT 77.335 65.080 77.565 65.260 ;
        RECT 82.625 65.130 82.855 65.260 ;
        RECT 77.255 55.160 77.615 65.080 ;
        RECT 82.565 55.180 82.935 65.130 ;
        RECT 83.765 65.090 83.995 65.260 ;
        RECT 83.695 55.140 84.065 65.090 ;
        RECT 85.055 65.080 85.285 65.260 ;
        RECT 88.585 65.090 88.815 65.270 ;
        RECT 93.875 65.140 94.105 65.270 ;
        RECT 84.965 55.190 85.385 65.080 ;
        RECT 88.505 55.170 88.865 65.090 ;
        RECT 93.815 55.190 94.185 65.140 ;
        RECT 95.015 65.100 95.245 65.270 ;
        RECT 94.945 55.150 95.315 65.100 ;
        RECT 96.305 65.090 96.535 65.270 ;
        RECT 96.215 55.200 96.635 65.090 ;
        RECT 99.865 65.080 100.095 65.260 ;
        RECT 105.155 65.130 105.385 65.260 ;
        RECT 99.785 55.160 100.145 65.080 ;
        RECT 105.095 55.180 105.465 65.130 ;
        RECT 106.295 65.090 106.525 65.260 ;
        RECT 106.225 55.140 106.595 65.090 ;
        RECT 107.585 65.080 107.815 65.260 ;
        RECT 111.135 65.080 111.365 65.260 ;
        RECT 116.425 65.130 116.655 65.260 ;
        RECT 107.495 55.190 107.915 65.080 ;
        RECT 111.055 55.160 111.415 65.080 ;
        RECT 116.365 55.180 116.735 65.130 ;
        RECT 117.565 65.090 117.795 65.260 ;
        RECT 117.495 55.140 117.865 65.090 ;
        RECT 118.855 65.080 119.085 65.260 ;
        RECT 122.385 65.080 122.615 65.260 ;
        RECT 127.675 65.130 127.905 65.260 ;
        RECT 118.765 55.190 119.185 65.080 ;
        RECT 122.305 55.160 122.665 65.080 ;
        RECT 127.615 55.180 127.985 65.130 ;
        RECT 128.815 65.090 129.045 65.260 ;
        RECT 128.745 55.140 129.115 65.090 ;
        RECT 130.105 65.080 130.335 65.260 ;
        RECT 133.135 65.130 133.365 65.230 ;
        RECT 130.015 55.190 130.435 65.080 ;
        RECT 133.005 55.240 133.405 65.130 ;
        RECT 138.425 65.100 138.655 65.230 ;
        RECT 133.135 55.230 133.365 55.240 ;
        RECT 138.345 55.130 138.725 65.100 ;
        RECT 149.340 64.660 150.720 65.760 ;
        RECT 20.815 54.230 25.555 54.530 ;
        RECT 32.015 54.240 36.755 54.540 ;
        RECT 43.235 54.210 47.975 54.510 ;
        RECT 54.485 54.190 59.225 54.490 ;
        RECT 65.705 54.180 70.445 54.480 ;
        RECT 76.945 54.170 81.685 54.470 ;
        RECT 88.195 54.180 92.935 54.480 ;
        RECT 99.475 54.170 104.215 54.470 ;
        RECT 110.745 54.170 115.485 54.470 ;
        RECT 121.995 54.170 126.735 54.470 ;
        RECT 21.655 52.320 22.115 52.550 ;
        RECT 25.625 52.280 26.255 52.560 ;
        RECT 25.735 52.240 26.195 52.280 ;
        RECT 27.665 52.240 28.125 52.470 ;
        RECT 32.855 52.330 33.315 52.560 ;
        RECT 36.825 52.290 37.455 52.570 ;
        RECT 36.935 52.250 37.395 52.290 ;
        RECT 38.865 52.250 39.325 52.480 ;
        RECT 44.075 52.300 44.535 52.530 ;
        RECT 48.045 52.260 48.675 52.540 ;
        RECT 48.155 52.220 48.615 52.260 ;
        RECT 50.085 52.220 50.545 52.450 ;
        RECT 55.325 52.280 55.785 52.510 ;
        RECT 59.295 52.240 59.925 52.520 ;
        RECT 59.405 52.200 59.865 52.240 ;
        RECT 61.335 52.200 61.795 52.430 ;
        RECT 66.545 52.270 67.005 52.500 ;
        RECT 70.515 52.230 71.145 52.510 ;
        RECT 70.625 52.190 71.085 52.230 ;
        RECT 72.555 52.190 73.015 52.420 ;
        RECT 77.785 52.260 78.245 52.490 ;
        RECT 81.755 52.220 82.385 52.500 ;
        RECT 81.865 52.180 82.325 52.220 ;
        RECT 83.795 52.180 84.255 52.410 ;
        RECT 89.035 52.270 89.495 52.500 ;
        RECT 93.005 52.230 93.635 52.510 ;
        RECT 93.115 52.190 93.575 52.230 ;
        RECT 95.045 52.190 95.505 52.420 ;
        RECT 100.315 52.260 100.775 52.490 ;
        RECT 104.285 52.220 104.915 52.500 ;
        RECT 104.395 52.180 104.855 52.220 ;
        RECT 106.325 52.180 106.785 52.410 ;
        RECT 111.585 52.260 112.045 52.490 ;
        RECT 115.555 52.220 116.185 52.500 ;
        RECT 115.665 52.180 116.125 52.220 ;
        RECT 117.595 52.180 118.055 52.410 ;
        RECT 122.835 52.260 123.295 52.490 ;
        RECT 126.805 52.220 127.435 52.500 ;
        RECT 126.915 52.180 127.375 52.220 ;
        RECT 128.845 52.180 129.305 52.410 ;
        RECT 21.375 52.010 21.605 52.115 ;
        RECT 21.245 50.290 21.615 52.010 ;
        RECT 22.165 51.890 22.395 52.115 ;
        RECT 25.455 51.980 25.685 52.035 ;
        RECT 21.375 50.115 21.605 50.290 ;
        RECT 22.155 50.210 22.525 51.890 ;
        RECT 22.165 50.115 22.395 50.210 ;
        RECT 21.525 49.670 22.245 49.930 ;
        RECT 19.295 46.650 20.065 47.720 ;
        RECT 21.385 47.490 22.105 47.750 ;
        RECT 21.225 47.200 21.455 47.340 ;
        RECT 21.085 46.430 21.475 47.200 ;
        RECT 22.015 47.190 22.245 47.340 ;
        RECT 22.005 46.450 22.375 47.190 ;
        RECT 25.305 47.010 25.735 51.980 ;
        RECT 26.245 51.970 26.475 52.035 ;
        RECT 27.385 51.970 27.615 52.035 ;
        RECT 26.185 46.970 26.585 51.970 ;
        RECT 27.265 46.970 27.665 51.970 ;
        RECT 28.175 51.940 28.405 52.035 ;
        RECT 32.575 52.020 32.805 52.125 ;
        RECT 28.115 46.970 28.545 51.940 ;
        RECT 32.445 50.300 32.815 52.020 ;
        RECT 33.365 51.900 33.595 52.125 ;
        RECT 36.655 51.990 36.885 52.045 ;
        RECT 32.575 50.125 32.805 50.300 ;
        RECT 33.355 50.220 33.725 51.900 ;
        RECT 33.365 50.125 33.595 50.220 ;
        RECT 32.725 49.680 33.445 49.940 ;
        RECT 25.735 46.600 26.195 46.830 ;
        RECT 27.665 46.710 28.125 46.830 ;
        RECT 27.515 46.600 28.125 46.710 ;
        RECT 30.495 46.660 31.265 47.730 ;
        RECT 32.585 47.500 33.305 47.760 ;
        RECT 32.425 47.210 32.655 47.350 ;
        RECT 21.225 46.340 21.455 46.430 ;
        RECT 22.015 46.340 22.245 46.450 ;
        RECT 27.515 46.430 28.095 46.600 ;
        RECT 32.285 46.440 32.675 47.210 ;
        RECT 33.215 47.200 33.445 47.350 ;
        RECT 33.205 46.460 33.575 47.200 ;
        RECT 36.505 47.020 36.935 51.990 ;
        RECT 37.445 51.980 37.675 52.045 ;
        RECT 38.585 51.980 38.815 52.045 ;
        RECT 37.385 46.980 37.785 51.980 ;
        RECT 38.465 46.980 38.865 51.980 ;
        RECT 39.375 51.950 39.605 52.045 ;
        RECT 43.795 51.990 44.025 52.095 ;
        RECT 39.315 46.980 39.745 51.950 ;
        RECT 43.665 50.270 44.035 51.990 ;
        RECT 44.585 51.870 44.815 52.095 ;
        RECT 47.875 51.960 48.105 52.015 ;
        RECT 43.795 50.095 44.025 50.270 ;
        RECT 44.575 50.190 44.945 51.870 ;
        RECT 44.585 50.095 44.815 50.190 ;
        RECT 43.945 49.650 44.665 49.910 ;
        RECT 36.935 46.610 37.395 46.840 ;
        RECT 38.865 46.720 39.325 46.840 ;
        RECT 38.715 46.610 39.325 46.720 ;
        RECT 41.715 46.630 42.485 47.700 ;
        RECT 43.805 47.470 44.525 47.730 ;
        RECT 43.645 47.180 43.875 47.320 ;
        RECT 32.425 46.350 32.655 46.440 ;
        RECT 33.215 46.350 33.445 46.460 ;
        RECT 38.715 46.440 39.295 46.610 ;
        RECT 43.505 46.410 43.895 47.180 ;
        RECT 44.435 47.170 44.665 47.320 ;
        RECT 44.425 46.430 44.795 47.170 ;
        RECT 47.725 46.990 48.155 51.960 ;
        RECT 48.665 51.950 48.895 52.015 ;
        RECT 49.805 51.950 50.035 52.015 ;
        RECT 48.605 46.950 49.005 51.950 ;
        RECT 49.685 46.950 50.085 51.950 ;
        RECT 50.595 51.920 50.825 52.015 ;
        RECT 55.045 51.970 55.275 52.075 ;
        RECT 50.535 46.950 50.965 51.920 ;
        RECT 54.915 50.250 55.285 51.970 ;
        RECT 55.835 51.850 56.065 52.075 ;
        RECT 59.125 51.940 59.355 51.995 ;
        RECT 55.045 50.075 55.275 50.250 ;
        RECT 55.825 50.170 56.195 51.850 ;
        RECT 55.835 50.075 56.065 50.170 ;
        RECT 55.195 49.630 55.915 49.890 ;
        RECT 48.155 46.580 48.615 46.810 ;
        RECT 50.085 46.690 50.545 46.810 ;
        RECT 49.935 46.580 50.545 46.690 ;
        RECT 52.965 46.610 53.735 47.680 ;
        RECT 55.055 47.450 55.775 47.710 ;
        RECT 54.895 47.160 55.125 47.300 ;
        RECT 43.645 46.320 43.875 46.410 ;
        RECT 44.435 46.320 44.665 46.430 ;
        RECT 49.935 46.410 50.515 46.580 ;
        RECT 54.755 46.390 55.145 47.160 ;
        RECT 55.685 47.150 55.915 47.300 ;
        RECT 55.675 46.410 56.045 47.150 ;
        RECT 58.975 46.970 59.405 51.940 ;
        RECT 59.915 51.930 60.145 51.995 ;
        RECT 61.055 51.930 61.285 51.995 ;
        RECT 59.855 46.930 60.255 51.930 ;
        RECT 60.935 46.930 61.335 51.930 ;
        RECT 61.845 51.900 62.075 51.995 ;
        RECT 66.265 51.960 66.495 52.065 ;
        RECT 61.785 46.930 62.215 51.900 ;
        RECT 66.135 50.240 66.505 51.960 ;
        RECT 67.055 51.840 67.285 52.065 ;
        RECT 70.345 51.930 70.575 51.985 ;
        RECT 66.265 50.065 66.495 50.240 ;
        RECT 67.045 50.160 67.415 51.840 ;
        RECT 67.055 50.065 67.285 50.160 ;
        RECT 66.415 49.620 67.135 49.880 ;
        RECT 59.405 46.560 59.865 46.790 ;
        RECT 61.335 46.670 61.795 46.790 ;
        RECT 61.185 46.560 61.795 46.670 ;
        RECT 64.185 46.600 64.955 47.670 ;
        RECT 66.275 47.440 66.995 47.700 ;
        RECT 66.115 47.150 66.345 47.290 ;
        RECT 54.895 46.300 55.125 46.390 ;
        RECT 55.685 46.300 55.915 46.410 ;
        RECT 61.185 46.390 61.765 46.560 ;
        RECT 65.975 46.380 66.365 47.150 ;
        RECT 66.905 47.140 67.135 47.290 ;
        RECT 66.895 46.400 67.265 47.140 ;
        RECT 70.195 46.960 70.625 51.930 ;
        RECT 71.135 51.920 71.365 51.985 ;
        RECT 72.275 51.920 72.505 51.985 ;
        RECT 71.075 46.920 71.475 51.920 ;
        RECT 72.155 46.920 72.555 51.920 ;
        RECT 73.065 51.890 73.295 51.985 ;
        RECT 77.505 51.950 77.735 52.055 ;
        RECT 73.005 46.920 73.435 51.890 ;
        RECT 77.375 50.230 77.745 51.950 ;
        RECT 78.295 51.830 78.525 52.055 ;
        RECT 81.585 51.920 81.815 51.975 ;
        RECT 77.505 50.055 77.735 50.230 ;
        RECT 78.285 50.150 78.655 51.830 ;
        RECT 78.295 50.055 78.525 50.150 ;
        RECT 77.655 49.610 78.375 49.870 ;
        RECT 70.625 46.550 71.085 46.780 ;
        RECT 72.555 46.660 73.015 46.780 ;
        RECT 72.405 46.550 73.015 46.660 ;
        RECT 75.425 46.590 76.195 47.660 ;
        RECT 77.515 47.430 78.235 47.690 ;
        RECT 77.355 47.140 77.585 47.280 ;
        RECT 66.115 46.290 66.345 46.380 ;
        RECT 66.905 46.290 67.135 46.400 ;
        RECT 72.405 46.380 72.985 46.550 ;
        RECT 77.215 46.370 77.605 47.140 ;
        RECT 78.145 47.130 78.375 47.280 ;
        RECT 78.135 46.390 78.505 47.130 ;
        RECT 81.435 46.950 81.865 51.920 ;
        RECT 82.375 51.910 82.605 51.975 ;
        RECT 83.515 51.910 83.745 51.975 ;
        RECT 82.315 46.910 82.715 51.910 ;
        RECT 83.395 46.910 83.795 51.910 ;
        RECT 84.305 51.880 84.535 51.975 ;
        RECT 88.755 51.960 88.985 52.065 ;
        RECT 84.245 46.910 84.675 51.880 ;
        RECT 88.625 50.240 88.995 51.960 ;
        RECT 89.545 51.840 89.775 52.065 ;
        RECT 92.835 51.930 93.065 51.985 ;
        RECT 88.755 50.065 88.985 50.240 ;
        RECT 89.535 50.160 89.905 51.840 ;
        RECT 89.545 50.065 89.775 50.160 ;
        RECT 88.905 49.620 89.625 49.880 ;
        RECT 81.865 46.540 82.325 46.770 ;
        RECT 83.795 46.650 84.255 46.770 ;
        RECT 83.645 46.540 84.255 46.650 ;
        RECT 86.675 46.600 87.445 47.670 ;
        RECT 88.765 47.440 89.485 47.700 ;
        RECT 88.605 47.150 88.835 47.290 ;
        RECT 77.355 46.280 77.585 46.370 ;
        RECT 78.145 46.280 78.375 46.390 ;
        RECT 83.645 46.370 84.225 46.540 ;
        RECT 88.465 46.380 88.855 47.150 ;
        RECT 89.395 47.140 89.625 47.290 ;
        RECT 89.385 46.400 89.755 47.140 ;
        RECT 92.685 46.960 93.115 51.930 ;
        RECT 93.625 51.920 93.855 51.985 ;
        RECT 94.765 51.920 94.995 51.985 ;
        RECT 93.565 46.920 93.965 51.920 ;
        RECT 94.645 46.920 95.045 51.920 ;
        RECT 95.555 51.890 95.785 51.985 ;
        RECT 100.035 51.950 100.265 52.055 ;
        RECT 95.495 46.920 95.925 51.890 ;
        RECT 99.905 50.230 100.275 51.950 ;
        RECT 100.825 51.830 101.055 52.055 ;
        RECT 104.115 51.920 104.345 51.975 ;
        RECT 100.035 50.055 100.265 50.230 ;
        RECT 100.815 50.150 101.185 51.830 ;
        RECT 100.825 50.055 101.055 50.150 ;
        RECT 100.185 49.610 100.905 49.870 ;
        RECT 93.115 46.550 93.575 46.780 ;
        RECT 95.045 46.660 95.505 46.780 ;
        RECT 94.895 46.550 95.505 46.660 ;
        RECT 97.955 46.590 98.725 47.660 ;
        RECT 100.045 47.430 100.765 47.690 ;
        RECT 99.885 47.140 100.115 47.280 ;
        RECT 88.605 46.290 88.835 46.380 ;
        RECT 89.395 46.290 89.625 46.400 ;
        RECT 94.895 46.380 95.475 46.550 ;
        RECT 99.745 46.370 100.135 47.140 ;
        RECT 100.675 47.130 100.905 47.280 ;
        RECT 100.665 46.390 101.035 47.130 ;
        RECT 103.965 46.950 104.395 51.920 ;
        RECT 104.905 51.910 105.135 51.975 ;
        RECT 106.045 51.910 106.275 51.975 ;
        RECT 104.845 46.910 105.245 51.910 ;
        RECT 105.925 46.910 106.325 51.910 ;
        RECT 106.835 51.880 107.065 51.975 ;
        RECT 111.305 51.950 111.535 52.055 ;
        RECT 106.775 46.910 107.205 51.880 ;
        RECT 111.175 50.230 111.545 51.950 ;
        RECT 112.095 51.830 112.325 52.055 ;
        RECT 115.385 51.920 115.615 51.975 ;
        RECT 111.305 50.055 111.535 50.230 ;
        RECT 112.085 50.150 112.455 51.830 ;
        RECT 112.095 50.055 112.325 50.150 ;
        RECT 111.455 49.610 112.175 49.870 ;
        RECT 104.395 46.540 104.855 46.770 ;
        RECT 106.325 46.650 106.785 46.770 ;
        RECT 106.175 46.540 106.785 46.650 ;
        RECT 109.225 46.590 109.995 47.660 ;
        RECT 111.315 47.430 112.035 47.690 ;
        RECT 111.155 47.140 111.385 47.280 ;
        RECT 99.885 46.280 100.115 46.370 ;
        RECT 100.675 46.280 100.905 46.390 ;
        RECT 106.175 46.370 106.755 46.540 ;
        RECT 111.015 46.370 111.405 47.140 ;
        RECT 111.945 47.130 112.175 47.280 ;
        RECT 111.935 46.390 112.305 47.130 ;
        RECT 115.235 46.950 115.665 51.920 ;
        RECT 116.175 51.910 116.405 51.975 ;
        RECT 117.315 51.910 117.545 51.975 ;
        RECT 116.115 46.910 116.515 51.910 ;
        RECT 117.195 46.910 117.595 51.910 ;
        RECT 118.105 51.880 118.335 51.975 ;
        RECT 122.555 51.950 122.785 52.055 ;
        RECT 118.045 46.910 118.475 51.880 ;
        RECT 122.425 50.230 122.795 51.950 ;
        RECT 123.345 51.830 123.575 52.055 ;
        RECT 126.635 51.920 126.865 51.975 ;
        RECT 122.555 50.055 122.785 50.230 ;
        RECT 123.335 50.150 123.705 51.830 ;
        RECT 123.345 50.055 123.575 50.150 ;
        RECT 122.705 49.610 123.425 49.870 ;
        RECT 115.665 46.540 116.125 46.770 ;
        RECT 117.595 46.650 118.055 46.770 ;
        RECT 117.445 46.540 118.055 46.650 ;
        RECT 120.475 46.590 121.245 47.660 ;
        RECT 122.565 47.430 123.285 47.690 ;
        RECT 122.405 47.140 122.635 47.280 ;
        RECT 111.155 46.280 111.385 46.370 ;
        RECT 111.945 46.280 112.175 46.390 ;
        RECT 117.445 46.370 118.025 46.540 ;
        RECT 122.265 46.370 122.655 47.140 ;
        RECT 123.195 47.130 123.425 47.280 ;
        RECT 123.185 46.390 123.555 47.130 ;
        RECT 126.485 46.950 126.915 51.920 ;
        RECT 127.425 51.910 127.655 51.975 ;
        RECT 128.565 51.910 128.795 51.975 ;
        RECT 127.365 46.910 127.765 51.910 ;
        RECT 128.445 46.910 128.845 51.910 ;
        RECT 129.355 51.880 129.585 51.975 ;
        RECT 129.295 46.910 129.725 51.880 ;
        RECT 126.915 46.540 127.375 46.770 ;
        RECT 128.845 46.650 129.305 46.770 ;
        RECT 128.695 46.540 129.305 46.650 ;
        RECT 122.405 46.280 122.635 46.370 ;
        RECT 123.195 46.280 123.425 46.390 ;
        RECT 128.695 46.370 129.275 46.540 ;
        RECT 21.505 45.950 21.965 46.180 ;
        RECT 32.705 45.960 33.165 46.190 ;
        RECT 43.925 45.930 44.385 46.160 ;
        RECT 55.175 45.910 55.635 46.140 ;
        RECT 66.395 45.900 66.855 46.130 ;
        RECT 77.635 45.890 78.095 46.120 ;
        RECT 88.885 45.900 89.345 46.130 ;
        RECT 100.165 45.890 100.625 46.120 ;
        RECT 111.435 45.890 111.895 46.120 ;
        RECT 122.685 45.890 123.145 46.120 ;
        RECT 29.055 45.020 41.225 45.030 ;
        RECT 17.855 45.005 41.225 45.020 ;
        RECT 15.900 45.000 41.225 45.005 ;
        RECT 15.900 44.980 52.445 45.000 ;
        RECT 15.900 44.970 63.695 44.980 ;
        RECT 15.900 44.960 74.915 44.970 ;
        RECT 85.235 44.960 97.405 44.970 ;
        RECT 15.900 43.880 131.205 44.960 ;
        RECT 15.900 43.870 30.025 43.880 ;
        RECT 15.900 43.855 18.690 43.870 ;
        RECT 15.900 41.620 17.050 43.855 ;
        RECT 40.275 43.850 131.205 43.880 ;
        RECT 51.525 43.830 131.205 43.850 ;
        RECT 62.745 43.820 131.205 43.830 ;
        RECT 73.985 43.810 86.155 43.820 ;
        RECT 96.515 43.810 131.205 43.820 ;
        RECT 29.015 43.330 41.185 43.340 ;
        RECT 17.815 43.310 41.185 43.330 ;
        RECT 142.830 43.320 144.150 43.340 ;
        RECT 17.815 43.290 52.405 43.310 ;
        RECT 140.750 43.300 144.150 43.320 ;
        RECT 17.815 43.280 63.655 43.290 ;
        RECT 119.895 43.280 144.150 43.300 ;
        RECT 17.815 43.270 74.875 43.280 ;
        RECT 85.195 43.270 97.365 43.280 ;
        RECT 108.685 43.270 144.150 43.280 ;
        RECT 17.815 42.180 144.150 43.270 ;
        RECT 18.755 42.150 144.150 42.180 ;
        RECT 18.755 42.120 131.165 42.150 ;
        RECT 18.755 42.090 109.655 42.120 ;
        RECT 18.755 42.080 98.445 42.090 ;
        RECT 41.325 42.070 98.445 42.080 ;
        RECT 142.830 42.070 144.150 42.150 ;
        RECT 41.325 42.060 87.205 42.070 ;
        RECT 75.035 42.050 87.205 42.060 ;
        RECT 15.900 41.540 19.685 41.620 ;
        RECT 142.070 41.610 146.210 41.640 ;
        RECT 119.855 41.590 146.210 41.610 ;
        RECT 108.645 41.550 146.210 41.590 ;
        RECT 15.900 41.520 42.165 41.540 ;
        RECT 97.445 41.530 146.210 41.550 ;
        RECT 15.900 41.510 75.875 41.520 ;
        RECT 86.235 41.510 146.210 41.530 ;
        RECT 15.900 40.500 146.210 41.510 ;
        RECT 15.900 40.480 142.320 40.500 ;
        RECT 15.900 40.470 140.920 40.480 ;
        RECT 18.715 40.460 140.920 40.470 ;
        RECT 142.070 40.460 142.250 40.480 ;
        RECT 18.715 40.440 120.815 40.460 ;
        RECT 18.715 40.400 109.615 40.440 ;
        RECT 18.715 40.390 98.405 40.400 ;
        RECT 41.285 40.380 98.405 40.390 ;
        RECT 41.285 40.370 87.165 40.380 ;
        RECT 74.995 40.360 87.165 40.370 ;
        RECT 26.775 39.230 27.235 39.460 ;
        RECT 38.055 39.230 38.515 39.460 ;
        RECT 49.345 39.210 49.805 39.440 ;
        RECT 60.565 39.210 61.025 39.440 ;
        RECT 71.765 39.210 72.225 39.440 ;
        RECT 83.055 39.200 83.515 39.430 ;
        RECT 94.295 39.220 94.755 39.450 ;
        RECT 105.505 39.240 105.965 39.470 ;
        RECT 116.705 39.280 117.165 39.510 ;
        RECT 127.915 39.300 128.375 39.530 ;
        RECT 20.645 38.810 21.225 38.980 ;
        RECT 26.495 38.960 26.725 39.070 ;
        RECT 27.285 38.980 27.515 39.070 ;
        RECT 20.615 38.700 21.225 38.810 ;
        RECT 20.615 38.580 21.075 38.700 ;
        RECT 22.545 38.580 23.005 38.810 ;
        RECT 20.195 33.470 20.625 38.440 ;
        RECT 20.335 33.375 20.565 33.470 ;
        RECT 21.075 33.440 21.475 38.440 ;
        RECT 22.155 33.440 22.555 38.440 ;
        RECT 21.125 33.375 21.355 33.440 ;
        RECT 22.265 33.375 22.495 33.440 ;
        RECT 23.005 33.430 23.435 38.400 ;
        RECT 26.365 38.220 26.735 38.960 ;
        RECT 26.495 38.070 26.725 38.220 ;
        RECT 27.265 38.210 27.655 38.980 ;
        RECT 31.925 38.810 32.505 38.980 ;
        RECT 37.775 38.960 38.005 39.070 ;
        RECT 38.565 38.980 38.795 39.070 ;
        RECT 27.285 38.070 27.515 38.210 ;
        RECT 26.635 37.660 27.355 37.920 ;
        RECT 28.675 37.690 29.445 38.760 ;
        RECT 31.895 38.700 32.505 38.810 ;
        RECT 31.895 38.580 32.355 38.700 ;
        RECT 33.825 38.580 34.285 38.810 ;
        RECT 26.495 35.480 27.215 35.740 ;
        RECT 26.345 35.200 26.575 35.295 ;
        RECT 26.215 33.520 26.585 35.200 ;
        RECT 27.135 35.120 27.365 35.295 ;
        RECT 23.055 33.375 23.285 33.430 ;
        RECT 26.345 33.295 26.575 33.520 ;
        RECT 27.125 33.400 27.495 35.120 ;
        RECT 31.475 33.470 31.905 38.440 ;
        RECT 27.135 33.295 27.365 33.400 ;
        RECT 31.615 33.375 31.845 33.470 ;
        RECT 32.355 33.440 32.755 38.440 ;
        RECT 33.435 33.440 33.835 38.440 ;
        RECT 32.405 33.375 32.635 33.440 ;
        RECT 33.545 33.375 33.775 33.440 ;
        RECT 34.285 33.430 34.715 38.400 ;
        RECT 37.645 38.220 38.015 38.960 ;
        RECT 37.775 38.070 38.005 38.220 ;
        RECT 38.545 38.210 38.935 38.980 ;
        RECT 43.215 38.790 43.795 38.960 ;
        RECT 49.065 38.940 49.295 39.050 ;
        RECT 49.855 38.960 50.085 39.050 ;
        RECT 38.565 38.070 38.795 38.210 ;
        RECT 37.915 37.660 38.635 37.920 ;
        RECT 39.955 37.690 40.725 38.760 ;
        RECT 43.185 38.680 43.795 38.790 ;
        RECT 43.185 38.560 43.645 38.680 ;
        RECT 45.115 38.560 45.575 38.790 ;
        RECT 37.775 35.480 38.495 35.740 ;
        RECT 37.625 35.200 37.855 35.295 ;
        RECT 37.495 33.520 37.865 35.200 ;
        RECT 38.415 35.120 38.645 35.295 ;
        RECT 34.335 33.375 34.565 33.430 ;
        RECT 37.625 33.295 37.855 33.520 ;
        RECT 38.405 33.400 38.775 35.120 ;
        RECT 42.765 33.450 43.195 38.420 ;
        RECT 38.415 33.295 38.645 33.400 ;
        RECT 42.905 33.355 43.135 33.450 ;
        RECT 43.645 33.420 44.045 38.420 ;
        RECT 44.725 33.420 45.125 38.420 ;
        RECT 43.695 33.355 43.925 33.420 ;
        RECT 44.835 33.355 45.065 33.420 ;
        RECT 45.575 33.410 46.005 38.380 ;
        RECT 48.935 38.200 49.305 38.940 ;
        RECT 49.065 38.050 49.295 38.200 ;
        RECT 49.835 38.190 50.225 38.960 ;
        RECT 54.435 38.790 55.015 38.960 ;
        RECT 60.285 38.940 60.515 39.050 ;
        RECT 61.075 38.960 61.305 39.050 ;
        RECT 49.855 38.050 50.085 38.190 ;
        RECT 49.205 37.640 49.925 37.900 ;
        RECT 51.245 37.670 52.015 38.740 ;
        RECT 54.405 38.680 55.015 38.790 ;
        RECT 54.405 38.560 54.865 38.680 ;
        RECT 56.335 38.560 56.795 38.790 ;
        RECT 49.065 35.460 49.785 35.720 ;
        RECT 48.915 35.180 49.145 35.275 ;
        RECT 48.785 33.500 49.155 35.180 ;
        RECT 49.705 35.100 49.935 35.275 ;
        RECT 45.625 33.355 45.855 33.410 ;
        RECT 48.915 33.275 49.145 33.500 ;
        RECT 49.695 33.380 50.065 35.100 ;
        RECT 53.985 33.450 54.415 38.420 ;
        RECT 49.705 33.275 49.935 33.380 ;
        RECT 54.125 33.355 54.355 33.450 ;
        RECT 54.865 33.420 55.265 38.420 ;
        RECT 55.945 33.420 56.345 38.420 ;
        RECT 54.915 33.355 55.145 33.420 ;
        RECT 56.055 33.355 56.285 33.420 ;
        RECT 56.795 33.410 57.225 38.380 ;
        RECT 60.155 38.200 60.525 38.940 ;
        RECT 60.285 38.050 60.515 38.200 ;
        RECT 61.055 38.190 61.445 38.960 ;
        RECT 65.635 38.790 66.215 38.960 ;
        RECT 71.485 38.940 71.715 39.050 ;
        RECT 72.275 38.960 72.505 39.050 ;
        RECT 61.075 38.050 61.305 38.190 ;
        RECT 60.425 37.640 61.145 37.900 ;
        RECT 62.465 37.670 63.235 38.740 ;
        RECT 65.605 38.680 66.215 38.790 ;
        RECT 65.605 38.560 66.065 38.680 ;
        RECT 67.535 38.560 67.995 38.790 ;
        RECT 60.285 35.460 61.005 35.720 ;
        RECT 60.135 35.180 60.365 35.275 ;
        RECT 60.005 33.500 60.375 35.180 ;
        RECT 60.925 35.100 61.155 35.275 ;
        RECT 56.845 33.355 57.075 33.410 ;
        RECT 60.135 33.275 60.365 33.500 ;
        RECT 60.915 33.380 61.285 35.100 ;
        RECT 65.185 33.450 65.615 38.420 ;
        RECT 60.925 33.275 61.155 33.380 ;
        RECT 65.325 33.355 65.555 33.450 ;
        RECT 66.065 33.420 66.465 38.420 ;
        RECT 67.145 33.420 67.545 38.420 ;
        RECT 66.115 33.355 66.345 33.420 ;
        RECT 67.255 33.355 67.485 33.420 ;
        RECT 67.995 33.410 68.425 38.380 ;
        RECT 71.355 38.200 71.725 38.940 ;
        RECT 71.485 38.050 71.715 38.200 ;
        RECT 72.255 38.190 72.645 38.960 ;
        RECT 76.925 38.780 77.505 38.950 ;
        RECT 82.775 38.930 83.005 39.040 ;
        RECT 83.565 38.950 83.795 39.040 ;
        RECT 72.275 38.050 72.505 38.190 ;
        RECT 71.625 37.640 72.345 37.900 ;
        RECT 73.665 37.670 74.435 38.740 ;
        RECT 76.895 38.670 77.505 38.780 ;
        RECT 76.895 38.550 77.355 38.670 ;
        RECT 78.825 38.550 79.285 38.780 ;
        RECT 71.485 35.460 72.205 35.720 ;
        RECT 71.335 35.180 71.565 35.275 ;
        RECT 71.205 33.500 71.575 35.180 ;
        RECT 72.125 35.100 72.355 35.275 ;
        RECT 68.045 33.355 68.275 33.410 ;
        RECT 71.335 33.275 71.565 33.500 ;
        RECT 72.115 33.380 72.485 35.100 ;
        RECT 76.475 33.440 76.905 38.410 ;
        RECT 72.125 33.275 72.355 33.380 ;
        RECT 76.615 33.345 76.845 33.440 ;
        RECT 77.355 33.410 77.755 38.410 ;
        RECT 78.435 33.410 78.835 38.410 ;
        RECT 77.405 33.345 77.635 33.410 ;
        RECT 78.545 33.345 78.775 33.410 ;
        RECT 79.285 33.400 79.715 38.370 ;
        RECT 82.645 38.190 83.015 38.930 ;
        RECT 82.775 38.040 83.005 38.190 ;
        RECT 83.545 38.180 83.935 38.950 ;
        RECT 88.165 38.800 88.745 38.970 ;
        RECT 94.015 38.950 94.245 39.060 ;
        RECT 94.805 38.970 95.035 39.060 ;
        RECT 83.565 38.040 83.795 38.180 ;
        RECT 82.915 37.630 83.635 37.890 ;
        RECT 84.955 37.660 85.725 38.730 ;
        RECT 88.135 38.690 88.745 38.800 ;
        RECT 88.135 38.570 88.595 38.690 ;
        RECT 90.065 38.570 90.525 38.800 ;
        RECT 82.775 35.450 83.495 35.710 ;
        RECT 82.625 35.170 82.855 35.265 ;
        RECT 82.495 33.490 82.865 35.170 ;
        RECT 83.415 35.090 83.645 35.265 ;
        RECT 79.335 33.345 79.565 33.400 ;
        RECT 82.625 33.265 82.855 33.490 ;
        RECT 83.405 33.370 83.775 35.090 ;
        RECT 87.715 33.460 88.145 38.430 ;
        RECT 83.415 33.265 83.645 33.370 ;
        RECT 87.855 33.365 88.085 33.460 ;
        RECT 88.595 33.430 88.995 38.430 ;
        RECT 89.675 33.430 90.075 38.430 ;
        RECT 88.645 33.365 88.875 33.430 ;
        RECT 89.785 33.365 90.015 33.430 ;
        RECT 90.525 33.420 90.955 38.390 ;
        RECT 93.885 38.210 94.255 38.950 ;
        RECT 94.015 38.060 94.245 38.210 ;
        RECT 94.785 38.200 95.175 38.970 ;
        RECT 99.375 38.820 99.955 38.990 ;
        RECT 105.225 38.970 105.455 39.080 ;
        RECT 106.015 38.990 106.245 39.080 ;
        RECT 94.805 38.060 95.035 38.200 ;
        RECT 94.155 37.650 94.875 37.910 ;
        RECT 96.195 37.680 96.965 38.750 ;
        RECT 99.345 38.710 99.955 38.820 ;
        RECT 99.345 38.590 99.805 38.710 ;
        RECT 101.275 38.590 101.735 38.820 ;
        RECT 94.015 35.470 94.735 35.730 ;
        RECT 93.865 35.190 94.095 35.285 ;
        RECT 93.735 33.510 94.105 35.190 ;
        RECT 94.655 35.110 94.885 35.285 ;
        RECT 90.575 33.365 90.805 33.420 ;
        RECT 93.865 33.285 94.095 33.510 ;
        RECT 94.645 33.390 95.015 35.110 ;
        RECT 98.925 33.480 99.355 38.450 ;
        RECT 94.655 33.285 94.885 33.390 ;
        RECT 99.065 33.385 99.295 33.480 ;
        RECT 99.805 33.450 100.205 38.450 ;
        RECT 100.885 33.450 101.285 38.450 ;
        RECT 99.855 33.385 100.085 33.450 ;
        RECT 100.995 33.385 101.225 33.450 ;
        RECT 101.735 33.440 102.165 38.410 ;
        RECT 105.095 38.230 105.465 38.970 ;
        RECT 105.225 38.080 105.455 38.230 ;
        RECT 105.995 38.220 106.385 38.990 ;
        RECT 110.575 38.860 111.155 39.030 ;
        RECT 116.425 39.010 116.655 39.120 ;
        RECT 117.215 39.030 117.445 39.120 ;
        RECT 106.015 38.080 106.245 38.220 ;
        RECT 105.365 37.670 106.085 37.930 ;
        RECT 107.405 37.700 108.175 38.770 ;
        RECT 110.545 38.750 111.155 38.860 ;
        RECT 110.545 38.630 111.005 38.750 ;
        RECT 112.475 38.630 112.935 38.860 ;
        RECT 105.225 35.490 105.945 35.750 ;
        RECT 105.075 35.210 105.305 35.305 ;
        RECT 104.945 33.530 105.315 35.210 ;
        RECT 105.865 35.130 106.095 35.305 ;
        RECT 101.785 33.385 102.015 33.440 ;
        RECT 105.075 33.305 105.305 33.530 ;
        RECT 105.855 33.410 106.225 35.130 ;
        RECT 110.125 33.520 110.555 38.490 ;
        RECT 110.265 33.425 110.495 33.520 ;
        RECT 111.005 33.490 111.405 38.490 ;
        RECT 112.085 33.490 112.485 38.490 ;
        RECT 111.055 33.425 111.285 33.490 ;
        RECT 112.195 33.425 112.425 33.490 ;
        RECT 112.935 33.480 113.365 38.450 ;
        RECT 116.295 38.270 116.665 39.010 ;
        RECT 116.425 38.120 116.655 38.270 ;
        RECT 117.195 38.260 117.585 39.030 ;
        RECT 121.785 38.880 122.365 39.050 ;
        RECT 127.635 39.030 127.865 39.140 ;
        RECT 128.425 39.050 128.655 39.140 ;
        RECT 117.215 38.120 117.445 38.260 ;
        RECT 116.565 37.710 117.285 37.970 ;
        RECT 118.605 37.740 119.375 38.810 ;
        RECT 121.755 38.770 122.365 38.880 ;
        RECT 121.755 38.650 122.215 38.770 ;
        RECT 123.685 38.650 124.145 38.880 ;
        RECT 116.425 35.530 117.145 35.790 ;
        RECT 116.275 35.250 116.505 35.345 ;
        RECT 116.145 33.570 116.515 35.250 ;
        RECT 117.065 35.170 117.295 35.345 ;
        RECT 112.985 33.425 113.215 33.480 ;
        RECT 105.865 33.305 106.095 33.410 ;
        RECT 116.275 33.345 116.505 33.570 ;
        RECT 117.055 33.450 117.425 35.170 ;
        RECT 121.335 33.540 121.765 38.510 ;
        RECT 117.065 33.345 117.295 33.450 ;
        RECT 121.475 33.445 121.705 33.540 ;
        RECT 122.215 33.510 122.615 38.510 ;
        RECT 123.295 33.510 123.695 38.510 ;
        RECT 122.265 33.445 122.495 33.510 ;
        RECT 123.405 33.445 123.635 33.510 ;
        RECT 124.145 33.500 124.575 38.470 ;
        RECT 127.505 38.290 127.875 39.030 ;
        RECT 127.635 38.140 127.865 38.290 ;
        RECT 128.405 38.280 128.795 39.050 ;
        RECT 128.425 38.140 128.655 38.280 ;
        RECT 127.775 37.730 128.495 37.990 ;
        RECT 129.815 37.760 130.585 38.830 ;
        RECT 142.850 37.630 144.170 38.900 ;
        RECT 127.635 35.550 128.355 35.810 ;
        RECT 127.485 35.270 127.715 35.365 ;
        RECT 127.355 33.590 127.725 35.270 ;
        RECT 128.275 35.190 128.505 35.365 ;
        RECT 124.195 33.445 124.425 33.500 ;
        RECT 127.485 33.365 127.715 33.590 ;
        RECT 128.265 33.470 128.635 35.190 ;
        RECT 128.275 33.365 128.505 33.470 ;
        RECT 20.615 32.940 21.075 33.170 ;
        RECT 22.545 33.130 23.005 33.170 ;
        RECT 22.485 32.850 23.115 33.130 ;
        RECT 26.625 32.860 27.085 33.090 ;
        RECT 31.895 32.940 32.355 33.170 ;
        RECT 33.825 33.130 34.285 33.170 ;
        RECT 33.765 32.850 34.395 33.130 ;
        RECT 37.905 32.860 38.365 33.090 ;
        RECT 43.185 32.920 43.645 33.150 ;
        RECT 45.115 33.110 45.575 33.150 ;
        RECT 45.055 32.830 45.685 33.110 ;
        RECT 49.195 32.840 49.655 33.070 ;
        RECT 54.405 32.920 54.865 33.150 ;
        RECT 56.335 33.110 56.795 33.150 ;
        RECT 56.275 32.830 56.905 33.110 ;
        RECT 60.415 32.840 60.875 33.070 ;
        RECT 65.605 32.920 66.065 33.150 ;
        RECT 67.535 33.110 67.995 33.150 ;
        RECT 67.475 32.830 68.105 33.110 ;
        RECT 71.615 32.840 72.075 33.070 ;
        RECT 76.895 32.910 77.355 33.140 ;
        RECT 78.825 33.100 79.285 33.140 ;
        RECT 78.765 32.820 79.395 33.100 ;
        RECT 82.905 32.830 83.365 33.060 ;
        RECT 88.135 32.930 88.595 33.160 ;
        RECT 90.065 33.120 90.525 33.160 ;
        RECT 90.005 32.840 90.635 33.120 ;
        RECT 94.145 32.850 94.605 33.080 ;
        RECT 99.345 32.950 99.805 33.180 ;
        RECT 101.275 33.140 101.735 33.180 ;
        RECT 101.215 32.860 101.845 33.140 ;
        RECT 105.355 32.870 105.815 33.100 ;
        RECT 110.545 32.990 111.005 33.220 ;
        RECT 112.475 33.180 112.935 33.220 ;
        RECT 112.415 32.900 113.045 33.180 ;
        RECT 116.555 32.910 117.015 33.140 ;
        RECT 121.755 33.010 122.215 33.240 ;
        RECT 123.685 33.200 124.145 33.240 ;
        RECT 123.625 32.920 124.255 33.200 ;
        RECT 127.765 32.930 128.225 33.160 ;
        RECT 23.185 30.880 27.925 31.180 ;
        RECT 34.465 30.880 39.205 31.180 ;
        RECT 45.755 30.860 50.495 31.160 ;
        RECT 56.975 30.860 61.715 31.160 ;
        RECT 68.175 30.860 72.915 31.160 ;
        RECT 79.465 30.850 84.205 31.150 ;
        RECT 90.705 30.870 95.445 31.170 ;
        RECT 101.915 30.890 106.655 31.190 ;
        RECT 113.115 30.930 117.855 31.230 ;
        RECT 124.325 30.950 129.065 31.250 ;
        RECT 19.485 20.270 19.905 30.160 ;
        RECT 19.585 20.090 19.815 20.270 ;
        RECT 20.805 20.260 21.175 30.210 ;
        RECT 20.875 20.090 21.105 20.260 ;
        RECT 21.935 20.220 22.305 30.170 ;
        RECT 27.255 20.270 27.615 30.190 ;
        RECT 30.765 20.270 31.185 30.160 ;
        RECT 22.015 20.090 22.245 20.220 ;
        RECT 27.305 20.090 27.535 20.270 ;
        RECT 30.865 20.090 31.095 20.270 ;
        RECT 32.085 20.260 32.455 30.210 ;
        RECT 32.155 20.090 32.385 20.260 ;
        RECT 33.215 20.220 33.585 30.170 ;
        RECT 38.535 20.270 38.895 30.190 ;
        RECT 33.295 20.090 33.525 20.220 ;
        RECT 38.585 20.090 38.815 20.270 ;
        RECT 42.055 20.250 42.475 30.140 ;
        RECT 42.155 20.070 42.385 20.250 ;
        RECT 43.375 20.240 43.745 30.190 ;
        RECT 43.445 20.070 43.675 20.240 ;
        RECT 44.505 20.200 44.875 30.150 ;
        RECT 49.825 20.250 50.185 30.170 ;
        RECT 53.275 20.250 53.695 30.140 ;
        RECT 44.585 20.070 44.815 20.200 ;
        RECT 49.875 20.070 50.105 20.250 ;
        RECT 53.375 20.070 53.605 20.250 ;
        RECT 54.595 20.240 54.965 30.190 ;
        RECT 54.665 20.070 54.895 20.240 ;
        RECT 55.725 20.200 56.095 30.150 ;
        RECT 61.045 20.250 61.405 30.170 ;
        RECT 64.475 20.250 64.895 30.140 ;
        RECT 55.805 20.070 56.035 20.200 ;
        RECT 61.095 20.070 61.325 20.250 ;
        RECT 64.575 20.070 64.805 20.250 ;
        RECT 65.795 20.240 66.165 30.190 ;
        RECT 65.865 20.070 66.095 20.240 ;
        RECT 66.925 20.200 67.295 30.150 ;
        RECT 72.245 20.250 72.605 30.170 ;
        RECT 67.005 20.070 67.235 20.200 ;
        RECT 72.295 20.070 72.525 20.250 ;
        RECT 75.765 20.240 76.185 30.130 ;
        RECT 75.865 20.060 76.095 20.240 ;
        RECT 77.085 20.230 77.455 30.180 ;
        RECT 77.155 20.060 77.385 20.230 ;
        RECT 78.215 20.190 78.585 30.140 ;
        RECT 83.535 20.240 83.895 30.160 ;
        RECT 87.005 20.260 87.425 30.150 ;
        RECT 78.295 20.060 78.525 20.190 ;
        RECT 83.585 20.060 83.815 20.240 ;
        RECT 87.105 20.080 87.335 20.260 ;
        RECT 88.325 20.250 88.695 30.200 ;
        RECT 88.395 20.080 88.625 20.250 ;
        RECT 89.455 20.210 89.825 30.160 ;
        RECT 94.775 20.260 95.135 30.180 ;
        RECT 98.215 20.280 98.635 30.170 ;
        RECT 89.535 20.080 89.765 20.210 ;
        RECT 94.825 20.080 95.055 20.260 ;
        RECT 98.315 20.100 98.545 20.280 ;
        RECT 99.535 20.270 99.905 30.220 ;
        RECT 99.605 20.100 99.835 20.270 ;
        RECT 100.665 20.230 101.035 30.180 ;
        RECT 105.985 20.280 106.345 30.200 ;
        RECT 109.415 20.320 109.835 30.210 ;
        RECT 100.745 20.100 100.975 20.230 ;
        RECT 106.035 20.100 106.265 20.280 ;
        RECT 109.515 20.140 109.745 20.320 ;
        RECT 110.735 20.310 111.105 30.260 ;
        RECT 110.805 20.140 111.035 20.310 ;
        RECT 111.865 20.270 112.235 30.220 ;
        RECT 117.185 20.320 117.545 30.240 ;
        RECT 120.625 20.340 121.045 30.230 ;
        RECT 111.945 20.140 112.175 20.270 ;
        RECT 117.235 20.140 117.465 20.320 ;
        RECT 120.725 20.160 120.955 20.340 ;
        RECT 121.945 20.330 122.315 30.280 ;
        RECT 122.015 20.160 122.245 20.330 ;
        RECT 123.075 20.290 123.445 30.240 ;
        RECT 128.395 20.340 128.755 30.260 ;
        RECT 123.155 20.160 123.385 20.290 ;
        RECT 128.445 20.160 128.675 20.340 ;
        RECT 132.345 20.170 132.755 30.180 ;
        RECT 137.735 30.120 137.965 30.130 ;
        RECT 132.445 20.130 132.675 20.170 ;
        RECT 137.665 20.080 138.055 30.120 ;
        RECT 19.775 19.610 20.925 19.920 ;
        RECT 22.185 19.620 27.335 19.900 ;
        RECT 31.055 19.610 32.205 19.920 ;
        RECT 33.465 19.620 38.615 19.900 ;
        RECT 42.345 19.590 43.495 19.900 ;
        RECT 44.755 19.600 49.905 19.880 ;
        RECT 53.565 19.590 54.715 19.900 ;
        RECT 55.975 19.600 61.125 19.880 ;
        RECT 64.765 19.590 65.915 19.900 ;
        RECT 67.175 19.600 72.325 19.880 ;
        RECT 76.055 19.580 77.205 19.890 ;
        RECT 78.465 19.590 83.615 19.870 ;
        RECT 87.295 19.600 88.445 19.910 ;
        RECT 89.705 19.610 94.855 19.890 ;
        RECT 98.505 19.620 99.655 19.930 ;
        RECT 100.915 19.630 106.065 19.910 ;
        RECT 109.705 19.660 110.855 19.970 ;
        RECT 112.115 19.670 117.265 19.950 ;
        RECT 120.915 19.680 122.065 19.990 ;
        RECT 123.325 19.690 128.475 19.970 ;
        RECT 132.635 19.640 138.025 19.930 ;
        RECT 142.940 19.110 144.080 37.630 ;
        RECT 13.940 18.460 17.635 18.530 ;
        RECT 117.755 18.510 131.425 18.530 ;
        RECT 106.545 18.470 131.425 18.510 ;
        RECT 13.940 18.440 41.565 18.460 ;
        RECT 95.345 18.450 131.425 18.470 ;
        RECT 13.940 18.430 75.275 18.440 ;
        RECT 84.135 18.430 131.425 18.450 ;
        RECT 13.940 17.380 131.425 18.430 ;
        RECT 142.890 17.990 144.140 19.110 ;
        RECT 145.070 18.880 146.210 40.500 ;
        RECT 145.030 17.960 146.250 18.880 ;
        RECT 13.950 17.370 15.100 17.380 ;
        RECT 16.615 17.360 120.215 17.380 ;
        RECT 16.615 17.320 109.015 17.360 ;
        RECT 16.615 17.310 97.805 17.320 ;
        RECT 39.185 17.300 97.805 17.310 ;
        RECT 39.185 17.290 86.565 17.300 ;
        RECT 72.895 17.280 86.565 17.290 ;
        RECT 117.765 16.950 140.620 16.960 ;
        RECT 142.040 16.950 148.010 16.980 ;
        RECT 117.765 16.940 148.010 16.950 ;
        RECT 106.555 16.900 148.010 16.940 ;
        RECT 16.625 16.870 41.575 16.890 ;
        RECT 95.355 16.880 148.010 16.900 ;
        RECT 16.625 16.860 75.285 16.870 ;
        RECT 84.145 16.860 148.010 16.880 ;
        RECT 16.625 15.840 148.010 16.860 ;
        RECT 16.625 15.820 142.660 15.840 ;
        RECT 16.625 15.810 140.620 15.820 ;
        RECT 142.040 15.810 142.660 15.820 ;
        RECT 16.625 15.790 120.225 15.810 ;
        RECT 16.625 15.750 109.025 15.790 ;
        RECT 16.625 15.740 97.815 15.750 ;
        RECT 39.195 15.730 97.815 15.740 ;
        RECT 39.195 15.720 86.575 15.730 ;
        RECT 72.905 15.710 86.575 15.720 ;
        RECT 131.215 15.460 132.585 15.470 ;
        RECT 12.290 15.390 17.625 15.450 ;
        RECT 117.795 15.440 132.785 15.460 ;
        RECT 106.585 15.400 132.785 15.440 ;
        RECT 12.290 15.370 41.585 15.390 ;
        RECT 95.385 15.380 132.785 15.400 ;
        RECT 12.290 15.360 75.295 15.370 ;
        RECT 84.175 15.360 132.785 15.380 ;
        RECT 12.290 14.320 132.785 15.360 ;
        RECT 142.905 15.040 144.045 15.050 ;
        RECT 12.290 14.310 131.445 14.320 ;
        RECT 12.290 14.300 120.235 14.310 ;
        RECT 12.320 14.280 13.470 14.300 ;
        RECT 16.655 14.290 120.235 14.300 ;
        RECT 16.655 14.250 109.035 14.290 ;
        RECT 16.655 14.240 97.825 14.250 ;
        RECT 39.225 14.230 97.825 14.240 ;
        RECT 39.225 14.220 86.585 14.230 ;
        RECT 72.935 14.210 86.585 14.220 ;
        RECT 142.850 13.920 144.100 15.040 ;
        RECT 145.020 14.870 146.160 14.980 ;
        RECT 144.980 13.950 146.200 14.870 ;
        RECT 16.965 13.800 17.435 13.810 ;
        RECT 10.800 13.780 17.435 13.800 ;
        RECT 10.800 13.720 17.555 13.780 ;
        RECT 117.845 13.770 131.445 13.790 ;
        RECT 106.635 13.730 131.445 13.770 ;
        RECT 10.800 13.700 41.585 13.720 ;
        RECT 95.435 13.710 131.445 13.730 ;
        RECT 10.800 13.690 75.295 13.700 ;
        RECT 84.225 13.690 131.445 13.710 ;
        RECT 10.800 12.650 131.445 13.690 ;
        RECT 16.705 12.640 131.445 12.650 ;
        RECT 16.705 12.620 120.235 12.640 ;
        RECT 16.705 12.580 109.035 12.620 ;
        RECT 16.705 12.570 97.825 12.580 ;
        RECT 39.275 12.560 97.825 12.570 ;
        RECT 39.275 12.550 86.585 12.560 ;
        RECT 72.985 12.540 86.585 12.550 ;
        RECT 128.755 12.240 130.465 12.250 ;
        RECT 117.545 12.220 119.255 12.230 ;
        RECT 106.345 12.180 108.055 12.190 ;
        RECT 27.615 12.170 29.325 12.180 ;
        RECT 38.895 12.170 40.605 12.180 ;
        RECT 25.675 11.030 29.325 12.170 ;
        RECT 36.955 11.030 40.605 12.170 ;
        RECT 95.135 12.160 96.845 12.170 ;
        RECT 50.185 12.150 51.895 12.160 ;
        RECT 61.405 12.150 63.115 12.160 ;
        RECT 72.605 12.150 74.315 12.160 ;
        RECT 25.675 11.020 27.625 11.030 ;
        RECT 36.955 11.020 38.905 11.030 ;
        RECT 48.245 11.010 51.895 12.150 ;
        RECT 59.465 11.010 63.115 12.150 ;
        RECT 70.665 11.010 74.315 12.150 ;
        RECT 83.895 12.140 85.605 12.150 ;
        RECT 48.245 11.000 50.195 11.010 ;
        RECT 59.465 11.000 61.415 11.010 ;
        RECT 70.665 11.000 72.615 11.010 ;
        RECT 81.955 11.000 85.605 12.140 ;
        RECT 93.195 11.020 96.845 12.160 ;
        RECT 104.405 11.040 108.055 12.180 ;
        RECT 115.605 11.080 119.255 12.220 ;
        RECT 126.815 11.100 130.465 12.240 ;
        RECT 126.815 11.090 128.765 11.100 ;
        RECT 115.605 11.070 117.555 11.080 ;
        RECT 104.405 11.030 106.355 11.040 ;
        RECT 93.195 11.010 95.145 11.020 ;
        RECT 81.955 10.990 83.905 11.000 ;
        RECT 142.905 8.580 144.045 13.920 ;
        RECT 74.420 7.440 144.045 8.580 ;
        RECT 74.420 1.410 75.560 7.440 ;
        RECT 145.020 6.630 146.160 13.950 ;
        RECT 93.650 5.490 146.160 6.630 ;
        RECT 93.650 1.480 94.790 5.490 ;
        RECT 146.870 4.560 148.010 15.840 ;
        RECT 113.130 3.420 148.010 4.560 ;
        RECT 113.130 1.610 114.270 3.420 ;
        RECT 149.460 2.770 150.600 64.660 ;
        RECT 131.940 1.880 150.600 2.770 ;
        RECT 131.800 1.630 150.600 1.880 ;
        RECT 74.290 0.160 75.680 1.410 ;
        RECT 93.500 0.230 94.890 1.480 ;
        RECT 112.900 0.360 114.290 1.610 ;
        RECT 131.800 1.380 133.490 1.630 ;
        RECT 151.730 1.420 152.870 66.900 ;
        RECT 131.800 0.430 133.540 1.380 ;
        RECT 113.130 0.330 114.270 0.360 ;
        RECT 151.600 0.300 152.970 1.420 ;
        RECT 93.650 0.150 94.790 0.230 ;
      LAYER met2 ;
        RECT 135.390 223.830 136.740 225.230 ;
        RECT 138.180 223.760 139.530 225.160 ;
        RECT 143.230 223.790 144.580 225.190 ;
        RECT 34.910 206.090 36.790 206.460 ;
        RECT 64.910 206.090 66.790 206.460 ;
        RECT 94.910 206.090 96.790 206.460 ;
        RECT 59.370 204.925 59.630 205.245 ;
        RECT 19.910 203.370 21.790 203.740 ;
        RECT 49.910 203.370 51.790 203.740 ;
        RECT 59.430 202.185 59.570 204.925 ;
        RECT 66.730 203.905 66.990 204.225 ;
        RECT 60.750 202.885 61.010 203.205 ;
        RECT 59.370 201.865 59.630 202.185 ;
        RECT 56.610 201.185 56.870 201.505 ;
        RECT 34.910 200.650 36.790 201.020 ;
        RECT 56.670 200.145 56.810 201.185 ;
        RECT 58.910 200.165 59.170 200.485 ;
        RECT 56.610 199.825 56.870 200.145 ;
        RECT 52.930 199.145 53.190 199.465 ;
        RECT 19.910 197.930 21.790 198.300 ;
        RECT 49.910 197.930 51.790 198.300 ;
        RECT 52.990 197.765 53.130 199.145 ;
        RECT 52.930 197.445 53.190 197.765 ;
        RECT 34.910 195.210 36.790 195.580 ;
        RECT 42.350 194.045 42.610 194.365 ;
        RECT 19.910 192.490 21.790 192.860 ;
        RECT 29.470 191.325 29.730 191.645 ;
        RECT 24.410 190.645 24.670 190.965 ;
        RECT 24.470 189.605 24.610 190.645 ;
        RECT 28.090 190.305 28.350 190.625 ;
        RECT 24.410 189.285 24.670 189.605 ;
        RECT 23.950 188.605 24.210 188.925 ;
        RECT 19.910 187.050 21.790 187.420 ;
        RECT 22.110 184.865 22.370 185.185 ;
        RECT 19.350 183.165 19.610 183.485 ;
        RECT 19.410 178.045 19.550 183.165 ;
        RECT 19.910 181.610 21.790 181.980 ;
        RECT 22.170 180.425 22.310 184.865 ;
        RECT 24.010 183.485 24.150 188.605 ;
        RECT 28.150 188.585 28.290 190.305 ;
        RECT 28.550 188.605 28.810 188.925 ;
        RECT 26.710 188.265 26.970 188.585 ;
        RECT 28.090 188.265 28.350 188.585 ;
        RECT 24.870 185.205 25.130 185.525 ;
        RECT 24.930 184.165 25.070 185.205 ;
        RECT 24.870 183.845 25.130 184.165 ;
        RECT 23.950 183.165 24.210 183.485 ;
        RECT 26.770 182.885 26.910 188.265 ;
        RECT 27.170 185.205 27.430 185.525 ;
        RECT 27.230 183.825 27.370 185.205 ;
        RECT 27.170 183.505 27.430 183.825 ;
        RECT 26.770 182.805 27.370 182.885 ;
        RECT 27.630 182.825 27.890 183.145 ;
        RECT 26.770 182.745 27.430 182.805 ;
        RECT 27.170 182.485 27.430 182.745 ;
        RECT 27.230 180.765 27.370 182.485 ;
        RECT 27.170 180.445 27.430 180.765 ;
        RECT 22.110 180.105 22.370 180.425 ;
        RECT 19.350 177.725 19.610 178.045 ;
        RECT 15.210 177.385 15.470 177.705 ;
        RECT 15.270 174.305 15.410 177.385 ;
        RECT 15.210 173.985 15.470 174.305 ;
        RECT 15.270 171.585 15.410 173.985 ;
        RECT 19.410 172.605 19.550 177.725 ;
        RECT 19.910 176.170 21.790 176.540 ;
        RECT 20.270 174.325 20.530 174.645 ;
        RECT 20.330 173.285 20.470 174.325 ;
        RECT 20.270 172.965 20.530 173.285 ;
        RECT 19.350 172.285 19.610 172.605 ;
        RECT 15.210 171.265 15.470 171.585 ;
        RECT 19.910 170.730 21.790 171.100 ;
        RECT 22.170 170.225 22.310 180.105 ;
        RECT 27.230 178.725 27.370 180.445 ;
        RECT 27.170 178.405 27.430 178.725 ;
        RECT 23.030 178.125 23.290 178.385 ;
        RECT 23.030 178.065 23.690 178.125 ;
        RECT 23.090 177.985 23.690 178.065 ;
        RECT 27.690 178.045 27.830 182.825 ;
        RECT 28.610 179.745 28.750 188.605 ;
        RECT 29.530 184.165 29.670 191.325 ;
        RECT 29.930 190.985 30.190 191.305 ;
        RECT 40.970 190.985 41.230 191.305 ;
        RECT 29.990 186.205 30.130 190.985 ;
        RECT 40.050 190.305 40.310 190.625 ;
        RECT 34.910 189.770 36.790 190.140 ;
        RECT 34.070 188.945 34.330 189.265 ;
        RECT 31.310 187.925 31.570 188.245 ;
        RECT 30.390 187.585 30.650 187.905 ;
        RECT 30.850 187.585 31.110 187.905 ;
        RECT 29.930 185.885 30.190 186.205 ;
        RECT 29.470 183.845 29.730 184.165 ;
        RECT 29.470 180.785 29.730 181.105 ;
        RECT 28.550 179.425 28.810 179.745 ;
        RECT 29.010 179.425 29.270 179.745 ;
        RECT 29.070 178.385 29.210 179.425 ;
        RECT 29.010 178.065 29.270 178.385 ;
        RECT 29.530 178.045 29.670 180.785 ;
        RECT 22.570 177.385 22.830 177.705 ;
        RECT 23.550 177.615 23.690 177.985 ;
        RECT 26.710 177.725 26.970 178.045 ;
        RECT 27.630 177.725 27.890 178.045 ;
        RECT 28.090 177.955 28.350 178.045 ;
        RECT 28.090 177.815 28.750 177.955 ;
        RECT 28.090 177.725 28.350 177.815 ;
        RECT 23.950 177.615 24.210 177.705 ;
        RECT 23.550 177.475 24.210 177.615 ;
        RECT 22.630 177.025 22.770 177.385 ;
        RECT 22.570 176.705 22.830 177.025 ;
        RECT 22.570 174.325 22.830 174.645 ;
        RECT 22.630 173.285 22.770 174.325 ;
        RECT 22.570 172.965 22.830 173.285 ;
        RECT 23.550 172.945 23.690 177.475 ;
        RECT 23.950 177.385 24.210 177.475 ;
        RECT 26.770 177.365 26.910 177.725 ;
        RECT 25.330 177.045 25.590 177.365 ;
        RECT 26.710 177.045 26.970 177.365 ;
        RECT 24.870 175.005 25.130 175.325 ;
        RECT 24.410 173.985 24.670 174.305 ;
        RECT 23.490 172.625 23.750 172.945 ;
        RECT 24.470 172.605 24.610 173.985 ;
        RECT 22.570 172.285 22.830 172.605 ;
        RECT 24.410 172.285 24.670 172.605 ;
        RECT 22.110 169.905 22.370 170.225 ;
        RECT 22.630 169.205 22.770 172.285 ;
        RECT 24.930 170.565 25.070 175.005 ;
        RECT 25.390 174.645 25.530 177.045 ;
        RECT 28.090 176.705 28.350 177.025 ;
        RECT 25.330 174.325 25.590 174.645 ;
        RECT 28.150 173.285 28.290 176.705 ;
        RECT 28.090 172.965 28.350 173.285 ;
        RECT 28.610 172.515 28.750 177.815 ;
        RECT 29.470 177.725 29.730 178.045 ;
        RECT 29.470 177.045 29.730 177.365 ;
        RECT 29.530 173.285 29.670 177.045 ;
        RECT 29.990 175.325 30.130 185.885 ;
        RECT 30.450 183.485 30.590 187.585 ;
        RECT 30.910 185.865 31.050 187.585 ;
        RECT 30.850 185.545 31.110 185.865 ;
        RECT 31.370 183.825 31.510 187.925 ;
        RECT 32.690 187.585 32.950 187.905 ;
        RECT 31.310 183.505 31.570 183.825 ;
        RECT 32.750 183.485 32.890 187.585 ;
        RECT 34.130 186.885 34.270 188.945 ;
        RECT 38.210 188.605 38.470 188.925 ;
        RECT 34.070 186.565 34.330 186.885 ;
        RECT 30.390 183.165 30.650 183.485 ;
        RECT 30.850 183.165 31.110 183.485 ;
        RECT 32.690 183.165 32.950 183.485 ;
        RECT 30.910 181.445 31.050 183.165 ;
        RECT 30.850 181.125 31.110 181.445 ;
        RECT 31.310 180.785 31.570 181.105 ;
        RECT 30.390 180.105 30.650 180.425 ;
        RECT 30.450 178.725 30.590 180.105 ;
        RECT 30.390 178.405 30.650 178.725 ;
        RECT 30.850 176.705 31.110 177.025 ;
        RECT 29.930 175.005 30.190 175.325 ;
        RECT 29.990 174.725 30.130 175.005 ;
        RECT 29.990 174.645 30.590 174.725 ;
        RECT 29.990 174.585 30.650 174.645 ;
        RECT 30.390 174.325 30.650 174.585 ;
        RECT 29.470 172.965 29.730 173.285 ;
        RECT 30.390 172.515 30.650 172.605 ;
        RECT 28.610 172.375 30.650 172.515 ;
        RECT 30.390 172.285 30.650 172.375 ;
        RECT 30.380 171.750 30.660 172.120 ;
        RECT 24.870 170.245 25.130 170.565 ;
        RECT 24.930 169.965 25.070 170.245 ;
        RECT 24.930 169.825 25.530 169.965 ;
        RECT 22.570 168.885 22.830 169.205 ;
        RECT 22.630 167.165 22.770 168.885 ;
        RECT 23.490 167.185 23.750 167.505 ;
        RECT 22.110 166.845 22.370 167.165 ;
        RECT 22.570 166.845 22.830 167.165 ;
        RECT 23.030 166.845 23.290 167.165 ;
        RECT 18.890 165.825 19.150 166.145 ;
        RECT 18.950 163.765 19.090 165.825 ;
        RECT 19.910 165.290 21.790 165.660 ;
        RECT 18.890 163.445 19.150 163.765 ;
        RECT 17.570 162.345 18.630 162.485 ;
        RECT 22.170 162.405 22.310 166.845 ;
        RECT 15.670 160.385 15.930 160.705 ;
        RECT 15.730 158.325 15.870 160.385 ;
        RECT 15.670 158.005 15.930 158.325 ;
        RECT 17.570 156.625 17.710 162.345 ;
        RECT 18.490 161.725 18.630 162.345 ;
        RECT 22.110 162.085 22.370 162.405 ;
        RECT 17.970 161.405 18.230 161.725 ;
        RECT 18.430 161.405 18.690 161.725 ;
        RECT 22.570 161.405 22.830 161.725 ;
        RECT 17.510 156.305 17.770 156.625 ;
        RECT 15.210 155.965 15.470 156.285 ;
        RECT 15.270 151.525 15.410 155.965 ;
        RECT 15.670 154.945 15.930 155.265 ;
        RECT 15.730 152.885 15.870 154.945 ;
        RECT 17.570 154.245 17.710 156.305 ;
        RECT 18.030 156.285 18.170 161.405 ;
        RECT 19.910 159.850 21.790 160.220 ;
        RECT 22.630 159.345 22.770 161.405 ;
        RECT 22.570 159.025 22.830 159.345 ;
        RECT 22.110 158.685 22.370 159.005 ;
        RECT 17.970 155.965 18.230 156.285 ;
        RECT 18.430 155.965 18.690 156.285 ;
        RECT 17.510 153.925 17.770 154.245 ;
        RECT 15.670 152.565 15.930 152.885 ;
        RECT 15.210 151.205 15.470 151.525 ;
        RECT 15.270 148.035 15.410 151.205 ;
        RECT 17.970 150.865 18.230 151.185 ;
        RECT 14.810 147.895 15.410 148.035 ;
        RECT 14.810 145.405 14.950 147.895 ;
        RECT 15.210 147.125 15.470 147.445 ;
        RECT 15.270 146.085 15.410 147.125 ;
        RECT 18.030 147.105 18.170 150.865 ;
        RECT 18.490 150.845 18.630 155.965 ;
        RECT 19.910 154.410 21.790 154.780 ;
        RECT 22.170 153.225 22.310 158.685 ;
        RECT 23.090 156.965 23.230 166.845 ;
        RECT 23.550 162.065 23.690 167.185 ;
        RECT 23.950 165.825 24.210 166.145 ;
        RECT 24.010 164.445 24.150 165.825 ;
        RECT 25.390 164.445 25.530 169.825 ;
        RECT 30.450 169.545 30.590 171.750 ;
        RECT 30.390 169.225 30.650 169.545 ;
        RECT 27.630 166.505 27.890 166.825 ;
        RECT 27.170 165.825 27.430 166.145 ;
        RECT 23.950 164.125 24.210 164.445 ;
        RECT 25.330 164.125 25.590 164.445 ;
        RECT 23.490 161.745 23.750 162.065 ;
        RECT 25.390 161.725 25.530 164.125 ;
        RECT 27.230 162.065 27.370 165.825 ;
        RECT 27.690 165.125 27.830 166.505 ;
        RECT 27.630 164.805 27.890 165.125 ;
        RECT 29.010 164.125 29.270 164.445 ;
        RECT 27.170 161.745 27.430 162.065 ;
        RECT 25.330 161.405 25.590 161.725 ;
        RECT 24.870 161.065 25.130 161.385 ;
        RECT 23.490 160.385 23.750 160.705 ;
        RECT 23.550 158.665 23.690 160.385 ;
        RECT 24.930 159.685 25.070 161.065 ;
        RECT 24.870 159.365 25.130 159.685 ;
        RECT 25.390 159.005 25.530 161.405 ;
        RECT 29.070 160.705 29.210 164.125 ;
        RECT 30.390 162.315 30.650 162.405 ;
        RECT 29.990 162.175 30.650 162.315 ;
        RECT 29.010 160.385 29.270 160.705 ;
        RECT 29.070 159.005 29.210 160.385 ;
        RECT 25.330 158.685 25.590 159.005 ;
        RECT 29.010 158.685 29.270 159.005 ;
        RECT 23.490 158.345 23.750 158.665 ;
        RECT 23.950 158.005 24.210 158.325 ;
        RECT 23.030 156.645 23.290 156.965 ;
        RECT 24.010 156.625 24.150 158.005 ;
        RECT 24.870 157.665 25.130 157.985 ;
        RECT 23.950 156.305 24.210 156.625 ;
        RECT 24.930 156.285 25.070 157.665 ;
        RECT 29.070 156.965 29.210 158.685 ;
        RECT 29.990 157.985 30.130 162.175 ;
        RECT 30.390 162.085 30.650 162.175 ;
        RECT 30.910 161.805 31.050 176.705 ;
        RECT 31.370 172.605 31.510 180.785 ;
        RECT 34.130 180.765 34.270 186.565 ;
        RECT 34.530 184.865 34.790 185.185 ;
        RECT 37.290 184.865 37.550 185.185 ;
        RECT 34.590 184.165 34.730 184.865 ;
        RECT 34.910 184.330 36.790 184.700 ;
        RECT 34.530 183.845 34.790 184.165 ;
        RECT 37.350 183.485 37.490 184.865 ;
        RECT 38.270 183.825 38.410 188.605 ;
        RECT 39.130 188.265 39.390 188.585 ;
        RECT 38.210 183.505 38.470 183.825 ;
        RECT 37.290 183.395 37.550 183.485 ;
        RECT 37.290 183.255 37.950 183.395 ;
        RECT 37.290 183.165 37.550 183.255 ;
        RECT 34.070 180.445 34.330 180.765 ;
        RECT 33.610 179.765 33.870 180.085 ;
        RECT 31.770 179.425 32.030 179.745 ;
        RECT 31.830 175.325 31.970 179.425 ;
        RECT 31.770 175.005 32.030 175.325 ;
        RECT 31.310 172.285 31.570 172.605 ;
        RECT 33.670 172.265 33.810 179.765 ;
        RECT 34.130 178.725 34.270 180.445 ;
        RECT 34.530 180.105 34.790 180.425 ;
        RECT 34.070 178.405 34.330 178.725 ;
        RECT 34.590 178.045 34.730 180.105 ;
        RECT 37.290 179.425 37.550 179.745 ;
        RECT 34.910 178.890 36.790 179.260 ;
        RECT 34.530 177.725 34.790 178.045 ;
        RECT 35.910 177.045 36.170 177.365 ;
        RECT 35.970 174.985 36.110 177.045 ;
        RECT 35.910 174.665 36.170 174.985 ;
        RECT 34.530 173.985 34.790 174.305 ;
        RECT 34.590 172.685 34.730 173.985 ;
        RECT 34.910 173.450 36.790 173.820 ;
        RECT 35.910 172.965 36.170 173.285 ;
        RECT 34.590 172.605 35.190 172.685 ;
        RECT 35.970 172.605 36.110 172.965 ;
        RECT 34.590 172.545 35.250 172.605 ;
        RECT 34.990 172.285 35.250 172.545 ;
        RECT 35.910 172.285 36.170 172.605 ;
        RECT 33.610 171.945 33.870 172.265 ;
        RECT 31.770 171.265 32.030 171.585 ;
        RECT 32.690 171.265 32.950 171.585 ;
        RECT 34.070 171.265 34.330 171.585 ;
        RECT 31.310 168.885 31.570 169.205 ;
        RECT 31.370 163.765 31.510 168.885 ;
        RECT 31.310 163.445 31.570 163.765 ;
        RECT 31.830 163.165 31.970 171.265 ;
        RECT 32.230 166.165 32.490 166.485 ;
        RECT 30.450 161.665 31.050 161.805 ;
        RECT 31.370 163.025 31.970 163.165 ;
        RECT 29.930 157.665 30.190 157.985 ;
        RECT 29.010 156.645 29.270 156.965 ;
        RECT 29.990 156.480 30.130 157.665 ;
        RECT 24.870 155.965 25.130 156.285 ;
        RECT 29.920 156.110 30.200 156.480 ;
        RECT 29.930 155.965 30.190 156.110 ;
        RECT 26.250 155.285 26.510 155.605 ;
        RECT 29.930 155.285 30.190 155.605 ;
        RECT 23.490 154.945 23.750 155.265 ;
        RECT 23.550 153.225 23.690 154.945 ;
        RECT 26.310 154.245 26.450 155.285 ;
        RECT 29.470 154.945 29.730 155.265 ;
        RECT 26.250 153.925 26.510 154.245 ;
        RECT 22.110 152.905 22.370 153.225 ;
        RECT 23.490 152.905 23.750 153.225 ;
        RECT 18.430 150.525 18.690 150.845 ;
        RECT 18.490 150.245 18.630 150.525 ;
        RECT 22.170 150.505 22.310 152.905 ;
        RECT 25.790 152.565 26.050 152.885 ;
        RECT 22.570 151.205 22.830 151.525 ;
        RECT 18.490 150.105 19.090 150.245 ;
        RECT 22.110 150.185 22.370 150.505 ;
        RECT 18.430 149.505 18.690 149.825 ;
        RECT 17.970 146.785 18.230 147.105 ;
        RECT 15.210 145.765 15.470 146.085 ;
        RECT 14.750 145.085 15.010 145.405 ;
        RECT 18.030 145.065 18.170 146.785 ;
        RECT 17.970 144.745 18.230 145.065 ;
        RECT 18.490 142.345 18.630 149.505 ;
        RECT 18.950 148.805 19.090 150.105 ;
        RECT 19.910 148.970 21.790 149.340 ;
        RECT 18.890 148.485 19.150 148.805 ;
        RECT 22.170 148.125 22.310 150.185 ;
        RECT 22.630 148.125 22.770 151.205 ;
        RECT 25.850 150.845 25.990 152.565 ;
        RECT 23.030 150.525 23.290 150.845 ;
        RECT 25.790 150.525 26.050 150.845 ;
        RECT 18.890 147.805 19.150 148.125 ;
        RECT 22.110 147.805 22.370 148.125 ;
        RECT 22.570 147.805 22.830 148.125 ;
        RECT 18.950 143.365 19.090 147.805 ;
        RECT 19.350 145.425 19.610 145.745 ;
        RECT 18.890 143.045 19.150 143.365 ;
        RECT 19.410 143.025 19.550 145.425 ;
        RECT 19.910 143.530 21.790 143.900 ;
        RECT 19.350 142.705 19.610 143.025 ;
        RECT 22.630 142.345 22.770 147.805 ;
        RECT 23.090 146.085 23.230 150.525 ;
        RECT 25.850 147.785 25.990 150.525 ;
        RECT 26.310 150.165 26.450 153.925 ;
        RECT 29.010 152.225 29.270 152.545 ;
        RECT 26.250 149.845 26.510 150.165 ;
        RECT 26.310 148.465 26.450 149.845 ;
        RECT 28.550 148.485 28.810 148.805 ;
        RECT 26.250 148.145 26.510 148.465 ;
        RECT 25.790 147.465 26.050 147.785 ;
        RECT 28.610 147.105 28.750 148.485 ;
        RECT 29.070 147.785 29.210 152.225 ;
        RECT 29.010 147.465 29.270 147.785 ;
        RECT 26.710 146.785 26.970 147.105 ;
        RECT 28.550 146.785 28.810 147.105 ;
        RECT 23.030 145.765 23.290 146.085 ;
        RECT 26.770 145.405 26.910 146.785 ;
        RECT 25.790 145.085 26.050 145.405 ;
        RECT 26.710 145.085 26.970 145.405 ;
        RECT 23.950 144.745 24.210 145.065 ;
        RECT 18.430 142.025 18.690 142.345 ;
        RECT 22.570 142.025 22.830 142.345 ;
        RECT 14.290 139.645 14.550 139.965 ;
        RECT 13.830 136.925 14.090 137.245 ;
        RECT 13.890 135.205 14.030 136.925 ;
        RECT 13.830 134.885 14.090 135.205 ;
        RECT 14.350 134.525 14.490 139.645 ;
        RECT 16.590 138.625 16.850 138.945 ;
        RECT 23.490 138.625 23.750 138.945 ;
        RECT 16.650 136.565 16.790 138.625 ;
        RECT 19.910 138.090 21.790 138.460 ;
        RECT 16.590 136.245 16.850 136.565 ;
        RECT 22.570 135.905 22.830 136.225 ;
        RECT 23.030 135.905 23.290 136.225 ;
        RECT 12.910 134.205 13.170 134.525 ;
        RECT 14.290 134.205 14.550 134.525 ;
        RECT 12.970 132.485 13.110 134.205 ;
        RECT 12.910 132.165 13.170 132.485 ;
        RECT 14.350 126.025 14.490 134.205 ;
        RECT 19.350 133.185 19.610 133.505 ;
        RECT 18.890 131.825 19.150 132.145 ;
        RECT 17.970 131.145 18.230 131.465 ;
        RECT 18.030 130.785 18.170 131.145 ;
        RECT 17.050 130.465 17.310 130.785 ;
        RECT 17.970 130.465 18.230 130.785 ;
        RECT 16.590 129.105 16.850 129.425 ;
        RECT 14.750 128.765 15.010 129.085 ;
        RECT 14.810 126.705 14.950 128.765 ;
        RECT 16.650 127.045 16.790 129.105 ;
        RECT 16.590 126.725 16.850 127.045 ;
        RECT 14.750 126.385 15.010 126.705 ;
        RECT 17.110 126.025 17.250 130.465 ;
        RECT 18.950 126.365 19.090 131.825 ;
        RECT 19.410 131.805 19.550 133.185 ;
        RECT 19.910 132.650 21.790 133.020 ;
        RECT 22.110 131.825 22.370 132.145 ;
        RECT 19.350 131.485 19.610 131.805 ;
        RECT 22.170 131.125 22.310 131.825 ;
        RECT 22.110 130.805 22.370 131.125 ;
        RECT 22.170 129.765 22.310 130.805 ;
        RECT 22.630 130.785 22.770 135.905 ;
        RECT 23.090 134.525 23.230 135.905 ;
        RECT 23.030 134.205 23.290 134.525 ;
        RECT 22.570 130.465 22.830 130.785 ;
        RECT 22.110 129.445 22.370 129.765 ;
        RECT 19.910 127.210 21.790 127.580 ;
        RECT 18.890 126.045 19.150 126.365 ;
        RECT 20.270 126.045 20.530 126.365 ;
        RECT 14.290 125.705 14.550 126.025 ;
        RECT 17.050 125.705 17.310 126.025 ;
        RECT 14.350 123.645 14.490 125.705 ;
        RECT 19.350 125.365 19.610 125.685 ;
        RECT 17.510 125.025 17.770 125.345 ;
        RECT 18.890 125.025 19.150 125.345 ;
        RECT 17.570 123.645 17.710 125.025 ;
        RECT 18.430 124.005 18.690 124.325 ;
        RECT 14.290 123.325 14.550 123.645 ;
        RECT 17.510 123.325 17.770 123.645 ;
        RECT 17.050 122.645 17.310 122.965 ;
        RECT 15.210 122.305 15.470 122.625 ;
        RECT 15.270 120.925 15.410 122.305 ;
        RECT 15.210 120.605 15.470 120.925 ;
        RECT 17.110 120.245 17.250 122.645 ;
        RECT 17.050 119.925 17.310 120.245 ;
        RECT 18.490 119.905 18.630 124.005 ;
        RECT 18.430 119.585 18.690 119.905 ;
        RECT 18.490 117.865 18.630 119.585 ;
        RECT 18.950 118.885 19.090 125.025 ;
        RECT 19.410 121.265 19.550 125.365 ;
        RECT 20.330 123.305 20.470 126.045 ;
        RECT 22.170 126.025 22.310 129.445 ;
        RECT 22.110 125.705 22.370 126.025 ;
        RECT 23.030 125.705 23.290 126.025 ;
        RECT 20.270 122.985 20.530 123.305 ;
        RECT 19.910 121.770 21.790 122.140 ;
        RECT 23.090 121.605 23.230 125.705 ;
        RECT 23.030 121.285 23.290 121.605 ;
        RECT 19.350 120.945 19.610 121.265 ;
        RECT 18.890 118.565 19.150 118.885 ;
        RECT 19.350 118.225 19.610 118.545 ;
        RECT 18.430 117.545 18.690 117.865 ;
        RECT 19.410 116.165 19.550 118.225 ;
        RECT 19.910 116.330 21.790 116.700 ;
        RECT 19.350 115.845 19.610 116.165 ;
        RECT 23.550 112.765 23.690 138.625 ;
        RECT 24.010 137.245 24.150 144.745 ;
        RECT 25.850 144.725 25.990 145.085 ;
        RECT 25.790 144.405 26.050 144.725 ;
        RECT 29.530 139.965 29.670 154.945 ;
        RECT 29.990 153.225 30.130 155.285 ;
        RECT 29.930 152.905 30.190 153.225 ;
        RECT 30.450 139.965 30.590 161.665 ;
        RECT 30.850 159.365 31.110 159.685 ;
        RECT 30.910 154.245 31.050 159.365 ;
        RECT 30.850 153.925 31.110 154.245 ;
        RECT 30.850 152.565 31.110 152.885 ;
        RECT 30.910 151.525 31.050 152.565 ;
        RECT 30.850 151.205 31.110 151.525 ;
        RECT 30.840 150.670 31.120 151.040 ;
        RECT 30.910 145.405 31.050 150.670 ;
        RECT 30.850 145.085 31.110 145.405 ;
        RECT 30.850 144.065 31.110 144.385 ;
        RECT 29.470 139.645 29.730 139.965 ;
        RECT 30.390 139.645 30.650 139.965 ;
        RECT 29.470 138.625 29.730 138.945 ;
        RECT 29.530 137.925 29.670 138.625 ;
        RECT 29.470 137.605 29.730 137.925 ;
        RECT 30.390 137.605 30.650 137.925 ;
        RECT 23.950 136.925 24.210 137.245 ;
        RECT 24.410 136.925 24.670 137.245 ;
        RECT 24.010 134.185 24.150 136.925 ;
        RECT 24.470 134.525 24.610 136.925 ;
        RECT 26.250 136.585 26.510 136.905 ;
        RECT 28.550 136.585 28.810 136.905 ;
        RECT 26.310 135.205 26.450 136.585 ;
        RECT 26.250 134.885 26.510 135.205 ;
        RECT 24.410 134.205 24.670 134.525 ;
        RECT 23.950 133.865 24.210 134.185 ;
        RECT 27.170 133.865 27.430 134.185 ;
        RECT 24.010 129.085 24.150 133.865 ;
        RECT 27.230 132.485 27.370 133.865 ;
        RECT 27.170 132.165 27.430 132.485 ;
        RECT 28.610 131.805 28.750 136.585 ;
        RECT 29.930 135.905 30.190 136.225 ;
        RECT 28.550 131.485 28.810 131.805 ;
        RECT 26.710 131.205 26.970 131.465 ;
        RECT 26.710 131.145 28.750 131.205 ;
        RECT 26.770 131.125 28.750 131.145 ;
        RECT 26.770 131.065 28.810 131.125 ;
        RECT 23.950 128.765 24.210 129.085 ;
        RECT 24.010 124.325 24.150 128.765 ;
        RECT 24.410 125.705 24.670 126.025 ;
        RECT 23.950 124.005 24.210 124.325 ;
        RECT 24.470 123.725 24.610 125.705 ;
        RECT 24.010 123.585 24.610 123.725 ;
        RECT 26.770 123.645 26.910 131.065 ;
        RECT 28.550 130.805 28.810 131.065 ;
        RECT 29.470 129.165 29.730 129.425 ;
        RECT 29.070 129.105 29.730 129.165 ;
        RECT 29.070 129.025 29.670 129.105 ;
        RECT 29.070 127.045 29.210 129.025 ;
        RECT 29.470 128.425 29.730 128.745 ;
        RECT 29.530 127.045 29.670 128.425 ;
        RECT 29.010 126.725 29.270 127.045 ;
        RECT 29.470 126.725 29.730 127.045 ;
        RECT 28.550 126.045 28.810 126.365 ;
        RECT 28.610 125.765 28.750 126.045 ;
        RECT 28.150 125.625 28.750 125.765 ;
        RECT 27.170 125.025 27.430 125.345 ;
        RECT 24.010 115.145 24.150 123.585 ;
        RECT 24.870 123.325 25.130 123.645 ;
        RECT 26.710 123.325 26.970 123.645 ;
        RECT 24.930 121.120 25.070 123.325 ;
        RECT 26.250 122.985 26.510 123.305 ;
        RECT 24.860 120.750 25.140 121.120 ;
        RECT 26.310 120.925 26.450 122.985 ;
        RECT 26.250 120.605 26.510 120.925 ;
        RECT 27.230 120.245 27.370 125.025 ;
        RECT 28.150 123.305 28.290 125.625 ;
        RECT 28.550 123.325 28.810 123.645 ;
        RECT 28.090 122.985 28.350 123.305 ;
        RECT 28.150 121.605 28.290 122.985 ;
        RECT 28.090 121.285 28.350 121.605 ;
        RECT 27.170 119.925 27.430 120.245 ;
        RECT 24.870 119.585 25.130 119.905 ;
        RECT 24.930 118.885 25.070 119.585 ;
        RECT 28.610 118.885 28.750 123.325 ;
        RECT 24.870 118.565 25.130 118.885 ;
        RECT 28.550 118.565 28.810 118.885 ;
        RECT 29.470 118.225 29.730 118.545 ;
        RECT 24.410 117.545 24.670 117.865 ;
        RECT 23.950 114.825 24.210 115.145 ;
        RECT 23.490 112.445 23.750 112.765 ;
        RECT 22.110 111.425 22.370 111.745 ;
        RECT 19.910 110.890 21.790 111.260 ;
        RECT 15.670 109.385 15.930 109.705 ;
        RECT 13.830 109.045 14.090 109.365 ;
        RECT 13.890 108.005 14.030 109.045 ;
        RECT 13.830 107.685 14.090 108.005 ;
        RECT 13.830 106.665 14.090 106.985 ;
        RECT 13.890 103.925 14.030 106.665 ;
        RECT 10.610 103.605 10.870 103.925 ;
        RECT 13.830 103.605 14.090 103.925 ;
        RECT 10.670 92.050 10.810 103.605 ;
        RECT 15.730 103.325 15.870 109.385 ;
        RECT 21.190 107.345 21.450 107.665 ;
        RECT 21.250 106.305 21.390 107.345 ;
        RECT 21.190 105.985 21.450 106.305 ;
        RECT 19.910 105.450 21.790 105.820 ;
        RECT 22.170 103.925 22.310 111.425 ;
        RECT 24.470 110.045 24.610 117.545 ;
        RECT 29.530 116.165 29.670 118.225 ;
        RECT 29.470 115.845 29.730 116.165 ;
        RECT 24.410 109.725 24.670 110.045 ;
        RECT 23.490 109.045 23.750 109.365 ;
        RECT 23.550 107.665 23.690 109.045 ;
        RECT 23.490 107.345 23.750 107.665 ;
        RECT 23.030 106.665 23.290 106.985 ;
        RECT 24.470 106.825 24.610 109.725 ;
        RECT 29.990 109.705 30.130 135.905 ;
        RECT 30.450 132.485 30.590 137.605 ;
        RECT 30.910 136.905 31.050 144.065 ;
        RECT 31.370 137.245 31.510 163.025 ;
        RECT 32.290 162.065 32.430 166.165 ;
        RECT 32.230 161.745 32.490 162.065 ;
        RECT 31.770 159.025 32.030 159.345 ;
        RECT 31.830 156.285 31.970 159.025 ;
        RECT 31.770 155.965 32.030 156.285 ;
        RECT 32.230 155.965 32.490 156.285 ;
        RECT 31.770 155.285 32.030 155.605 ;
        RECT 31.830 154.245 31.970 155.285 ;
        RECT 31.770 153.925 32.030 154.245 ;
        RECT 31.830 147.785 31.970 153.925 ;
        RECT 32.290 148.465 32.430 155.965 ;
        RECT 32.230 148.145 32.490 148.465 ;
        RECT 31.770 147.465 32.030 147.785 ;
        RECT 32.750 147.525 32.890 171.265 ;
        RECT 33.610 165.825 33.870 166.145 ;
        RECT 33.670 161.385 33.810 165.825 ;
        RECT 33.610 161.065 33.870 161.385 ;
        RECT 33.150 156.305 33.410 156.625 ;
        RECT 33.210 151.720 33.350 156.305 ;
        RECT 34.130 155.125 34.270 171.265 ;
        RECT 35.970 170.565 36.110 172.285 ;
        RECT 34.530 170.245 34.790 170.565 ;
        RECT 35.910 170.245 36.170 170.565 ;
        RECT 34.590 167.245 34.730 170.245 ;
        RECT 34.910 168.010 36.790 168.380 ;
        RECT 34.590 167.105 35.190 167.245 ;
        RECT 34.530 166.505 34.790 166.825 ;
        RECT 34.590 161.045 34.730 166.505 ;
        RECT 35.050 163.960 35.190 167.105 ;
        RECT 34.980 163.590 35.260 163.960 ;
        RECT 34.910 162.570 36.790 162.940 ;
        RECT 34.530 160.725 34.790 161.045 ;
        RECT 36.370 160.725 36.630 161.045 ;
        RECT 36.430 159.685 36.570 160.725 ;
        RECT 36.370 159.365 36.630 159.685 ;
        RECT 35.510 158.945 37.030 159.085 ;
        RECT 35.510 158.665 35.650 158.945 ;
        RECT 36.890 158.665 37.030 158.945 ;
        RECT 35.450 158.345 35.710 158.665 ;
        RECT 35.910 158.520 36.170 158.665 ;
        RECT 35.900 158.150 36.180 158.520 ;
        RECT 36.830 158.345 37.090 158.665 ;
        RECT 34.530 157.665 34.790 157.985 ;
        RECT 33.670 154.985 34.270 155.125 ;
        RECT 33.140 151.350 33.420 151.720 ;
        RECT 33.150 150.525 33.410 150.845 ;
        RECT 33.210 148.805 33.350 150.525 ;
        RECT 33.150 148.485 33.410 148.805 ;
        RECT 31.830 145.405 31.970 147.465 ;
        RECT 32.750 147.385 33.350 147.525 ;
        RECT 32.690 146.785 32.950 147.105 ;
        RECT 31.770 145.085 32.030 145.405 ;
        RECT 32.230 138.625 32.490 138.945 ;
        RECT 31.310 136.925 31.570 137.245 ;
        RECT 30.850 136.585 31.110 136.905 ;
        RECT 31.310 135.905 31.570 136.225 ;
        RECT 30.390 132.165 30.650 132.485 ;
        RECT 30.850 132.165 31.110 132.485 ;
        RECT 30.390 131.715 30.650 131.805 ;
        RECT 30.910 131.715 31.050 132.165 ;
        RECT 30.390 131.575 31.050 131.715 ;
        RECT 30.390 131.485 30.650 131.575 ;
        RECT 30.390 130.465 30.650 130.785 ;
        RECT 30.450 126.025 30.590 130.465 ;
        RECT 30.390 125.705 30.650 126.025 ;
        RECT 30.910 125.685 31.050 131.575 ;
        RECT 30.850 125.365 31.110 125.685 ;
        RECT 30.390 122.305 30.650 122.625 ;
        RECT 30.450 115.145 30.590 122.305 ;
        RECT 30.390 114.825 30.650 115.145 ;
        RECT 31.370 110.045 31.510 135.905 ;
        RECT 31.770 134.885 32.030 135.205 ;
        RECT 31.830 112.765 31.970 134.885 ;
        RECT 32.290 112.765 32.430 138.625 ;
        RECT 32.750 134.525 32.890 146.785 ;
        RECT 33.210 134.525 33.350 147.385 ;
        RECT 33.670 137.245 33.810 154.985 ;
        RECT 34.070 149.505 34.330 149.825 ;
        RECT 34.130 139.965 34.270 149.505 ;
        RECT 34.590 140.045 34.730 157.665 ;
        RECT 34.910 157.130 36.790 157.500 ;
        RECT 35.440 156.110 35.720 156.480 ;
        RECT 35.450 155.965 35.710 156.110 ;
        RECT 34.910 151.690 36.790 152.060 ;
        RECT 36.820 150.670 37.100 151.040 ;
        RECT 36.830 150.525 37.090 150.670 ;
        RECT 36.370 147.695 36.630 147.785 ;
        RECT 36.890 147.695 37.030 150.525 ;
        RECT 36.370 147.555 37.030 147.695 ;
        RECT 36.370 147.465 36.630 147.555 ;
        RECT 34.910 146.250 36.790 146.620 ;
        RECT 35.910 144.745 36.170 145.065 ;
        RECT 35.970 143.365 36.110 144.745 ;
        RECT 35.910 143.045 36.170 143.365 ;
        RECT 34.910 140.810 36.790 141.180 ;
        RECT 34.070 139.645 34.330 139.965 ;
        RECT 34.590 139.905 35.190 140.045 ;
        RECT 34.530 137.605 34.790 137.925 ;
        RECT 33.610 136.925 33.870 137.245 ;
        RECT 34.590 135.205 34.730 137.605 ;
        RECT 35.050 137.245 35.190 139.905 ;
        RECT 36.830 139.535 37.090 139.625 ;
        RECT 37.350 139.535 37.490 179.425 ;
        RECT 37.810 178.725 37.950 183.255 ;
        RECT 39.190 183.145 39.330 188.265 ;
        RECT 40.110 185.525 40.250 190.305 ;
        RECT 41.030 188.325 41.170 190.985 ;
        RECT 42.410 190.965 42.550 194.045 ;
        RECT 42.810 193.025 43.070 193.345 ;
        RECT 42.350 190.645 42.610 190.965 ;
        RECT 42.870 189.265 43.010 193.025 ;
        RECT 49.910 192.490 51.790 192.860 ;
        RECT 46.030 190.985 46.290 191.305 ;
        RECT 44.650 190.645 44.910 190.965 ;
        RECT 43.730 190.305 43.990 190.625 ;
        RECT 42.810 188.945 43.070 189.265 ;
        RECT 40.570 188.185 41.170 188.325 ;
        RECT 40.570 187.905 40.710 188.185 ;
        RECT 40.510 187.585 40.770 187.905 ;
        RECT 40.050 185.205 40.310 185.525 ;
        RECT 39.130 182.825 39.390 183.145 ;
        RECT 39.590 180.445 39.850 180.765 ;
        RECT 37.750 178.405 38.010 178.725 ;
        RECT 39.130 176.880 39.390 177.025 ;
        RECT 39.120 176.510 39.400 176.880 ;
        RECT 39.130 175.345 39.390 175.665 ;
        RECT 39.190 174.985 39.330 175.345 ;
        RECT 39.650 175.325 39.790 180.445 ;
        RECT 40.570 178.045 40.710 187.585 ;
        RECT 43.270 184.865 43.530 185.185 ;
        RECT 43.330 178.045 43.470 184.865 ;
        RECT 43.790 183.145 43.930 190.305 ;
        RECT 44.710 185.435 44.850 190.645 ;
        RECT 45.110 185.435 45.370 185.525 ;
        RECT 44.250 185.295 45.370 185.435 ;
        RECT 43.730 182.825 43.990 183.145 ;
        RECT 44.250 180.425 44.390 185.295 ;
        RECT 45.110 185.205 45.370 185.295 ;
        RECT 46.090 184.165 46.230 190.985 ;
        RECT 46.490 190.305 46.750 190.625 ;
        RECT 46.550 186.205 46.690 190.305 ;
        RECT 49.710 188.605 49.970 188.925 ;
        RECT 49.770 188.325 49.910 188.605 ;
        RECT 52.990 188.585 53.130 197.445 ;
        RECT 54.770 196.085 55.030 196.405 ;
        RECT 54.830 195.045 54.970 196.085 ;
        RECT 58.450 195.745 58.710 196.065 ;
        RECT 54.770 194.725 55.030 195.045 ;
        RECT 58.510 194.025 58.650 195.745 ;
        RECT 58.450 193.705 58.710 194.025 ;
        RECT 58.970 191.305 59.110 200.165 ;
        RECT 59.430 194.365 59.570 201.865 ;
        RECT 60.290 201.185 60.550 201.505 ;
        RECT 60.350 200.145 60.490 201.185 ;
        RECT 60.290 199.825 60.550 200.145 ;
        RECT 60.810 199.205 60.950 202.885 ;
        RECT 63.970 202.205 64.230 202.525 ;
        RECT 63.510 201.525 63.770 201.845 ;
        RECT 63.570 200.485 63.710 201.525 ;
        RECT 63.510 200.165 63.770 200.485 ;
        RECT 64.030 200.145 64.170 202.205 ;
        RECT 66.790 201.845 66.930 203.905 ;
        RECT 79.910 203.370 81.790 203.740 ;
        RECT 109.910 203.370 111.790 203.740 ;
        RECT 76.390 201.865 76.650 202.185 ;
        RECT 66.730 201.525 66.990 201.845 ;
        RECT 71.330 201.525 71.590 201.845 ;
        RECT 73.630 201.525 73.890 201.845 ;
        RECT 64.430 201.185 64.690 201.505 ;
        RECT 63.970 199.825 64.230 200.145 ;
        RECT 60.350 199.065 60.950 199.205 ;
        RECT 63.970 199.145 64.230 199.465 ;
        RECT 60.350 197.085 60.490 199.065 ;
        RECT 63.050 198.465 63.310 198.785 ;
        RECT 60.290 196.765 60.550 197.085 ;
        RECT 59.370 194.045 59.630 194.365 ;
        RECT 58.910 190.985 59.170 191.305 ;
        RECT 54.770 188.605 55.030 188.925 ;
        RECT 49.310 188.185 49.910 188.325 ;
        RECT 52.930 188.265 53.190 188.585 ;
        RECT 46.490 185.885 46.750 186.205 ;
        RECT 46.030 183.845 46.290 184.165 ;
        RECT 49.310 183.825 49.450 188.185 ;
        RECT 49.910 187.050 51.790 187.420 ;
        RECT 52.990 186.285 53.130 188.265 ;
        RECT 52.990 186.205 53.590 186.285 ;
        RECT 52.990 186.145 53.650 186.205 ;
        RECT 53.390 185.885 53.650 186.145 ;
        RECT 50.630 185.775 50.890 185.865 ;
        RECT 50.630 185.635 52.670 185.775 ;
        RECT 50.630 185.545 50.890 185.635 ;
        RECT 49.250 183.505 49.510 183.825 ;
        RECT 44.650 183.165 44.910 183.485 ;
        RECT 46.490 183.165 46.750 183.485 ;
        RECT 52.010 183.165 52.270 183.485 ;
        RECT 44.710 181.445 44.850 183.165 ;
        RECT 44.650 181.125 44.910 181.445 ;
        RECT 45.110 180.445 45.370 180.765 ;
        RECT 44.190 180.105 44.450 180.425 ;
        RECT 45.170 178.725 45.310 180.445 ;
        RECT 45.110 178.405 45.370 178.725 ;
        RECT 44.190 178.065 44.450 178.385 ;
        RECT 40.050 177.725 40.310 178.045 ;
        RECT 40.510 177.725 40.770 178.045 ;
        RECT 40.970 177.725 41.230 178.045 ;
        RECT 43.270 177.725 43.530 178.045 ;
        RECT 40.110 177.365 40.250 177.725 ;
        RECT 40.050 177.045 40.310 177.365 ;
        RECT 39.590 175.005 39.850 175.325 ;
        RECT 39.130 174.665 39.390 174.985 ;
        RECT 38.670 174.325 38.930 174.645 ;
        RECT 37.750 173.985 38.010 174.305 ;
        RECT 37.810 150.245 37.950 173.985 ;
        RECT 38.730 172.605 38.870 174.325 ;
        RECT 39.190 174.305 39.330 174.665 ;
        RECT 40.110 174.305 40.250 177.045 ;
        RECT 41.030 175.665 41.170 177.725 ;
        RECT 41.430 176.705 41.690 177.025 ;
        RECT 40.970 175.345 41.230 175.665 ;
        RECT 39.130 173.985 39.390 174.305 ;
        RECT 40.050 173.985 40.310 174.305 ;
        RECT 41.030 173.365 41.170 175.345 ;
        RECT 39.650 173.225 41.170 173.365 ;
        RECT 39.650 172.605 39.790 173.225 ;
        RECT 38.670 172.285 38.930 172.605 ;
        RECT 39.590 172.285 39.850 172.605 ;
        RECT 40.050 172.285 40.310 172.605 ;
        RECT 40.110 170.225 40.250 172.285 ;
        RECT 40.050 169.905 40.310 170.225 ;
        RECT 38.210 169.225 38.470 169.545 ;
        RECT 38.270 167.845 38.410 169.225 ;
        RECT 38.670 168.885 38.930 169.205 ;
        RECT 38.210 167.525 38.470 167.845 ;
        RECT 38.730 167.505 38.870 168.885 ;
        RECT 38.670 167.185 38.930 167.505 ;
        RECT 38.210 166.165 38.470 166.485 ;
        RECT 38.270 163.845 38.410 166.165 ;
        RECT 39.590 165.825 39.850 166.145 ;
        RECT 39.130 164.125 39.390 164.445 ;
        RECT 38.270 163.705 38.870 163.845 ;
        RECT 38.210 163.105 38.470 163.425 ;
        RECT 38.270 162.065 38.410 163.105 ;
        RECT 38.730 162.065 38.870 163.705 ;
        RECT 38.210 161.745 38.470 162.065 ;
        RECT 38.670 161.745 38.930 162.065 ;
        RECT 39.190 161.385 39.330 164.125 ;
        RECT 39.650 164.105 39.790 165.825 ;
        RECT 40.970 164.805 41.230 165.125 ;
        RECT 39.590 163.785 39.850 164.105 ;
        RECT 39.590 162.085 39.850 162.405 ;
        RECT 38.200 160.870 38.480 161.240 ;
        RECT 39.130 161.065 39.390 161.385 ;
        RECT 38.270 158.665 38.410 160.870 ;
        RECT 38.210 158.345 38.470 158.665 ;
        RECT 38.670 158.005 38.930 158.325 ;
        RECT 38.730 156.965 38.870 158.005 ;
        RECT 38.670 156.645 38.930 156.965 ;
        RECT 38.730 156.285 38.870 156.645 ;
        RECT 38.210 155.965 38.470 156.285 ;
        RECT 38.670 155.965 38.930 156.285 ;
        RECT 39.120 156.110 39.400 156.480 ;
        RECT 39.130 155.965 39.390 156.110 ;
        RECT 38.270 155.800 38.410 155.965 ;
        RECT 38.200 155.430 38.480 155.800 ;
        RECT 38.210 154.945 38.470 155.265 ;
        RECT 39.130 154.945 39.390 155.265 ;
        RECT 38.270 151.185 38.410 154.945 ;
        RECT 38.210 150.865 38.470 151.185 ;
        RECT 38.210 150.245 38.470 150.505 ;
        RECT 37.810 150.185 38.470 150.245 ;
        RECT 37.810 150.105 38.410 150.185 ;
        RECT 38.210 148.145 38.470 148.465 ;
        RECT 37.750 146.785 38.010 147.105 ;
        RECT 37.810 145.745 37.950 146.785 ;
        RECT 37.750 145.425 38.010 145.745 ;
        RECT 38.270 145.065 38.410 148.145 ;
        RECT 38.210 144.745 38.470 145.065 ;
        RECT 37.750 141.345 38.010 141.665 ;
        RECT 37.810 140.305 37.950 141.345 ;
        RECT 38.660 140.470 38.940 140.840 ;
        RECT 37.750 139.985 38.010 140.305 ;
        RECT 38.730 139.965 38.870 140.470 ;
        RECT 39.190 139.965 39.330 154.945 ;
        RECT 39.650 154.245 39.790 162.085 ;
        RECT 40.050 161.405 40.310 161.725 ;
        RECT 40.110 159.200 40.250 161.405 ;
        RECT 40.040 158.830 40.320 159.200 ;
        RECT 40.110 158.665 40.250 158.830 ;
        RECT 41.030 158.665 41.170 164.805 ;
        RECT 40.050 158.345 40.310 158.665 ;
        RECT 40.970 158.345 41.230 158.665 ;
        RECT 40.110 155.945 40.250 158.345 ;
        RECT 40.050 155.625 40.310 155.945 ;
        RECT 39.590 153.925 39.850 154.245 ;
        RECT 39.650 150.165 39.790 153.925 ;
        RECT 40.110 150.845 40.250 155.625 ;
        RECT 40.050 150.525 40.310 150.845 ;
        RECT 39.590 149.845 39.850 150.165 ;
        RECT 40.970 149.505 41.230 149.825 ;
        RECT 38.670 139.645 38.930 139.965 ;
        RECT 39.130 139.645 39.390 139.965 ;
        RECT 36.830 139.395 37.490 139.535 ;
        RECT 36.830 139.305 37.090 139.395 ;
        RECT 41.030 139.365 41.170 149.505 ;
        RECT 41.490 139.965 41.630 176.705 ;
        RECT 43.330 176.005 43.470 177.725 ;
        RECT 43.270 175.685 43.530 176.005 ;
        RECT 44.250 174.985 44.390 178.065 ;
        RECT 46.550 177.025 46.690 183.165 ;
        RECT 47.870 182.825 48.130 183.145 ;
        RECT 47.930 182.465 48.070 182.825 ;
        RECT 47.870 182.145 48.130 182.465 ;
        RECT 47.930 177.705 48.070 182.145 ;
        RECT 49.910 181.610 51.790 181.980 ;
        RECT 52.070 178.725 52.210 183.165 ;
        RECT 52.530 180.165 52.670 185.635 ;
        RECT 52.930 182.145 53.190 182.465 ;
        RECT 52.990 180.765 53.130 182.145 ;
        RECT 52.930 180.445 53.190 180.765 ;
        RECT 52.530 180.025 53.130 180.165 ;
        RECT 53.450 180.085 53.590 185.885 ;
        RECT 54.830 184.165 54.970 188.605 ;
        RECT 58.450 188.265 58.710 188.585 ;
        RECT 57.070 187.585 57.330 187.905 ;
        RECT 57.130 186.205 57.270 187.585 ;
        RECT 58.510 186.205 58.650 188.265 ;
        RECT 58.970 186.205 59.110 190.985 ;
        RECT 57.070 185.885 57.330 186.205 ;
        RECT 58.450 185.885 58.710 186.205 ;
        RECT 58.910 185.885 59.170 186.205 ;
        RECT 58.970 184.165 59.110 185.885 ;
        RECT 54.770 183.845 55.030 184.165 ;
        RECT 58.910 183.845 59.170 184.165 ;
        RECT 57.990 183.505 58.250 183.825 ;
        RECT 53.850 181.125 54.110 181.445 ;
        RECT 52.010 178.405 52.270 178.725 ;
        RECT 48.790 177.725 49.050 178.045 ;
        RECT 47.870 177.385 48.130 177.705 ;
        RECT 46.490 176.705 46.750 177.025 ;
        RECT 44.190 174.665 44.450 174.985 ;
        RECT 46.550 174.645 46.690 176.705 ;
        RECT 48.850 174.985 48.990 177.725 ;
        RECT 52.470 177.385 52.730 177.705 ;
        RECT 49.910 176.170 51.790 176.540 ;
        RECT 52.530 175.665 52.670 177.385 ;
        RECT 52.470 175.345 52.730 175.665 ;
        RECT 52.990 175.325 53.130 180.025 ;
        RECT 53.390 179.765 53.650 180.085 ;
        RECT 53.450 175.405 53.590 179.765 ;
        RECT 53.910 178.725 54.050 181.125 ;
        RECT 53.850 178.405 54.110 178.725 ;
        RECT 58.050 178.045 58.190 183.505 ;
        RECT 58.450 183.395 58.710 183.485 ;
        RECT 58.970 183.395 59.110 183.845 ;
        RECT 58.450 183.255 59.110 183.395 ;
        RECT 58.450 183.165 58.710 183.255 ;
        RECT 58.450 182.145 58.710 182.465 ;
        RECT 58.510 178.045 58.650 182.145 ;
        RECT 58.970 180.765 59.110 183.255 ;
        RECT 58.910 180.445 59.170 180.765 ;
        RECT 57.990 177.725 58.250 178.045 ;
        RECT 58.450 177.725 58.710 178.045 ;
        RECT 52.930 175.005 53.190 175.325 ;
        RECT 53.450 175.265 54.050 175.405 ;
        RECT 46.950 174.665 47.210 174.985 ;
        RECT 48.790 174.665 49.050 174.985 ;
        RECT 46.490 174.325 46.750 174.645 ;
        RECT 42.350 173.985 42.610 174.305 ;
        RECT 44.650 173.985 44.910 174.305 ;
        RECT 41.890 158.520 42.150 158.665 ;
        RECT 41.880 158.150 42.160 158.520 ;
        RECT 41.950 156.285 42.090 158.150 ;
        RECT 41.890 155.965 42.150 156.285 ;
        RECT 41.890 149.505 42.150 149.825 ;
        RECT 41.430 139.645 41.690 139.965 ;
        RECT 41.950 139.365 42.090 149.505 ;
        RECT 42.410 148.805 42.550 173.985 ;
        RECT 43.730 168.545 43.990 168.865 ;
        RECT 43.790 164.105 43.930 168.545 ;
        RECT 43.730 163.785 43.990 164.105 ;
        RECT 43.270 161.065 43.530 161.385 ;
        RECT 42.810 158.685 43.070 159.005 ;
        RECT 42.350 148.485 42.610 148.805 ;
        RECT 42.870 147.785 43.010 158.685 ;
        RECT 43.330 158.665 43.470 161.065 ;
        RECT 44.190 160.385 44.450 160.705 ;
        RECT 43.270 158.345 43.530 158.665 ;
        RECT 43.730 157.665 43.990 157.985 ;
        RECT 43.270 148.485 43.530 148.805 ;
        RECT 42.810 147.465 43.070 147.785 ;
        RECT 42.810 144.065 43.070 144.385 ;
        RECT 42.870 142.345 43.010 144.065 ;
        RECT 42.810 142.025 43.070 142.345 ;
        RECT 41.030 139.225 41.630 139.365 ;
        RECT 41.950 139.225 42.550 139.365 ;
        RECT 37.290 138.625 37.550 138.945 ;
        RECT 38.210 138.625 38.470 138.945 ;
        RECT 40.970 138.625 41.230 138.945 ;
        RECT 34.990 136.925 35.250 137.245 ;
        RECT 34.910 135.370 36.790 135.740 ;
        RECT 34.530 134.885 34.790 135.205 ;
        RECT 32.690 134.205 32.950 134.525 ;
        RECT 33.150 134.205 33.410 134.525 ;
        RECT 33.610 133.865 33.870 134.185 ;
        RECT 34.530 133.865 34.790 134.185 ;
        RECT 35.910 133.865 36.170 134.185 ;
        RECT 33.150 133.525 33.410 133.845 ;
        RECT 32.690 128.085 32.950 128.405 ;
        RECT 32.750 121.605 32.890 128.085 ;
        RECT 33.210 127.045 33.350 133.525 ;
        RECT 33.670 131.805 33.810 133.865 ;
        RECT 33.610 131.715 33.870 131.805 ;
        RECT 33.610 131.575 34.270 131.715 ;
        RECT 33.610 131.485 33.870 131.575 ;
        RECT 34.130 129.425 34.270 131.575 ;
        RECT 34.590 130.785 34.730 133.865 ;
        RECT 35.970 132.485 36.110 133.865 ;
        RECT 35.910 132.165 36.170 132.485 ;
        RECT 34.530 130.465 34.790 130.785 ;
        RECT 34.590 129.765 34.730 130.465 ;
        RECT 34.910 129.930 36.790 130.300 ;
        RECT 37.350 129.765 37.490 138.625 ;
        RECT 38.270 129.765 38.410 138.625 ;
        RECT 40.510 133.865 40.770 134.185 ;
        RECT 40.570 131.465 40.710 133.865 ;
        RECT 40.510 131.145 40.770 131.465 ;
        RECT 34.530 129.445 34.790 129.765 ;
        RECT 37.290 129.445 37.550 129.765 ;
        RECT 38.210 129.445 38.470 129.765 ;
        RECT 34.070 129.105 34.330 129.425 ;
        RECT 33.610 128.425 33.870 128.745 ;
        RECT 33.150 126.725 33.410 127.045 ;
        RECT 33.670 125.345 33.810 128.425 ;
        RECT 34.130 126.365 34.270 129.105 ;
        RECT 40.050 128.425 40.310 128.745 ;
        RECT 34.070 126.045 34.330 126.365 ;
        RECT 33.610 125.025 33.870 125.345 ;
        RECT 37.750 125.025 38.010 125.345 ;
        RECT 33.670 123.645 33.810 125.025 ;
        RECT 34.910 124.490 36.790 124.860 ;
        RECT 34.070 123.665 34.330 123.985 ;
        RECT 33.610 123.325 33.870 123.645 ;
        RECT 32.690 121.285 32.950 121.605 ;
        RECT 32.690 120.605 32.950 120.925 ;
        RECT 32.750 115.485 32.890 120.605 ;
        RECT 33.150 117.885 33.410 118.205 ;
        RECT 33.210 116.165 33.350 117.885 ;
        RECT 33.150 115.845 33.410 116.165 ;
        RECT 32.690 115.165 32.950 115.485 ;
        RECT 33.670 115.145 33.810 123.325 ;
        RECT 34.130 115.825 34.270 123.665 ;
        RECT 34.530 120.265 34.790 120.585 ;
        RECT 37.290 120.265 37.550 120.585 ;
        RECT 34.590 118.885 34.730 120.265 ;
        RECT 34.910 119.050 36.790 119.420 ;
        RECT 34.530 118.565 34.790 118.885 ;
        RECT 37.350 117.865 37.490 120.265 ;
        RECT 37.810 118.205 37.950 125.025 ;
        RECT 38.210 122.985 38.470 123.305 ;
        RECT 38.270 119.905 38.410 122.985 ;
        RECT 40.110 122.625 40.250 128.425 ;
        RECT 40.510 125.705 40.770 126.025 ;
        RECT 40.050 122.365 40.310 122.625 ;
        RECT 39.650 122.305 40.310 122.365 ;
        RECT 39.650 122.225 40.250 122.305 ;
        RECT 38.210 119.585 38.470 119.905 ;
        RECT 39.650 118.205 39.790 122.225 ;
        RECT 40.050 120.265 40.310 120.585 ;
        RECT 37.750 117.885 38.010 118.205 ;
        RECT 39.590 117.885 39.850 118.205 ;
        RECT 37.290 117.545 37.550 117.865 ;
        RECT 34.990 116.865 35.250 117.185 ;
        RECT 34.070 115.505 34.330 115.825 ;
        RECT 35.050 115.485 35.190 116.865 ;
        RECT 34.990 115.165 35.250 115.485 ;
        RECT 33.610 114.825 33.870 115.145 ;
        RECT 34.910 113.610 36.790 113.980 ;
        RECT 31.770 112.445 32.030 112.765 ;
        RECT 32.230 112.445 32.490 112.765 ;
        RECT 34.530 111.425 34.790 111.745 ;
        RECT 36.370 111.425 36.630 111.745 ;
        RECT 32.690 110.405 32.950 110.725 ;
        RECT 31.310 109.725 31.570 110.045 ;
        RECT 29.930 109.385 30.190 109.705 ;
        RECT 29.010 109.045 29.270 109.365 ;
        RECT 29.070 108.005 29.210 109.045 ;
        RECT 32.230 108.705 32.490 109.025 ;
        RECT 29.010 107.685 29.270 108.005 ;
        RECT 24.870 106.825 25.130 106.985 ;
        RECT 24.470 106.685 25.130 106.825 ;
        RECT 22.110 103.605 22.370 103.925 ;
        RECT 15.730 103.185 16.330 103.325 ;
        RECT 16.190 92.050 16.330 103.185 ;
        RECT 21.710 92.305 22.310 92.445 ;
        RECT 21.710 92.050 21.850 92.305 ;
        RECT 10.600 90.050 10.880 92.050 ;
        RECT 16.120 90.050 16.400 92.050 ;
        RECT 21.640 90.050 21.920 92.050 ;
        RECT 22.170 91.765 22.310 92.305 ;
        RECT 23.090 91.765 23.230 106.665 ;
        RECT 24.470 104.605 24.610 106.685 ;
        RECT 24.870 106.665 25.130 106.685 ;
        RECT 27.630 106.665 27.890 106.985 ;
        RECT 32.290 106.725 32.430 108.705 ;
        RECT 32.750 107.665 32.890 110.405 ;
        RECT 32.690 107.345 32.950 107.665 ;
        RECT 24.410 104.285 24.670 104.605 ;
        RECT 27.690 103.925 27.830 106.665 ;
        RECT 32.290 106.585 32.890 106.725 ;
        RECT 27.170 103.605 27.430 103.925 ;
        RECT 27.630 103.605 27.890 103.925 ;
        RECT 27.230 92.050 27.370 103.605 ;
        RECT 32.750 92.050 32.890 106.585 ;
        RECT 34.590 104.605 34.730 111.425 ;
        RECT 36.430 110.045 36.570 111.425 ;
        RECT 36.370 109.725 36.630 110.045 ;
        RECT 37.350 109.955 37.490 117.545 ;
        RECT 39.650 115.485 39.790 117.885 ;
        RECT 40.110 116.165 40.250 120.265 ;
        RECT 40.570 120.245 40.710 125.705 ;
        RECT 40.510 119.925 40.770 120.245 ;
        RECT 40.570 118.885 40.710 119.925 ;
        RECT 40.510 118.565 40.770 118.885 ;
        RECT 40.050 115.845 40.310 116.165 ;
        RECT 39.590 115.165 39.850 115.485 ;
        RECT 37.750 109.955 38.010 110.045 ;
        RECT 37.350 109.815 38.010 109.955 ;
        RECT 34.910 108.170 36.790 108.540 ;
        RECT 36.370 106.825 36.630 106.985 ;
        RECT 37.350 106.825 37.490 109.815 ;
        RECT 37.750 109.725 38.010 109.815 ;
        RECT 41.030 109.705 41.170 138.625 ;
        RECT 41.490 129.765 41.630 139.225 ;
        RECT 41.890 138.625 42.150 138.945 ;
        RECT 41.950 135.205 42.090 138.625 ;
        RECT 41.890 134.885 42.150 135.205 ;
        RECT 41.890 133.865 42.150 134.185 ;
        RECT 41.950 130.785 42.090 133.865 ;
        RECT 41.890 130.465 42.150 130.785 ;
        RECT 41.430 129.445 41.690 129.765 ;
        RECT 41.950 129.085 42.090 130.465 ;
        RECT 41.890 128.765 42.150 129.085 ;
        RECT 41.950 126.025 42.090 128.765 ;
        RECT 42.410 127.045 42.550 139.225 ;
        RECT 42.810 136.245 43.070 136.565 ;
        RECT 42.870 135.205 43.010 136.245 ;
        RECT 42.810 134.885 43.070 135.205 ;
        RECT 43.330 132.485 43.470 148.485 ;
        RECT 43.790 139.965 43.930 157.665 ;
        RECT 44.250 150.845 44.390 160.385 ;
        RECT 44.710 150.845 44.850 173.985 ;
        RECT 47.010 173.285 47.150 174.665 ;
        RECT 52.010 173.985 52.270 174.305 ;
        RECT 52.470 173.985 52.730 174.305 ;
        RECT 52.070 173.285 52.210 173.985 ;
        RECT 46.950 172.965 47.210 173.285 ;
        RECT 52.010 172.965 52.270 173.285 ;
        RECT 50.170 172.285 50.430 172.605 ;
        RECT 50.230 172.120 50.370 172.285 ;
        RECT 52.530 172.265 52.670 173.985 ;
        RECT 53.910 172.265 54.050 175.265 ;
        RECT 56.150 174.725 56.410 174.985 ;
        RECT 56.150 174.665 56.810 174.725 ;
        RECT 56.210 174.585 56.810 174.665 ;
        RECT 55.690 173.985 55.950 174.305 ;
        RECT 55.750 172.945 55.890 173.985 ;
        RECT 55.690 172.625 55.950 172.945 ;
        RECT 50.160 171.750 50.440 172.120 ;
        RECT 52.470 171.945 52.730 172.265 ;
        RECT 53.850 171.945 54.110 172.265 ;
        RECT 56.150 171.945 56.410 172.265 ;
        RECT 46.490 171.265 46.750 171.585 ;
        RECT 55.230 171.265 55.490 171.585 ;
        RECT 46.550 168.865 46.690 171.265 ;
        RECT 49.910 170.730 51.790 171.100 ;
        RECT 47.410 169.565 47.670 169.885 ;
        RECT 46.490 168.545 46.750 168.865 ;
        RECT 46.550 167.165 46.690 168.545 ;
        RECT 46.490 166.845 46.750 167.165 ;
        RECT 45.110 166.505 45.370 166.825 ;
        RECT 45.170 162.405 45.310 166.505 ;
        RECT 46.030 163.105 46.290 163.425 ;
        RECT 45.110 162.085 45.370 162.405 ;
        RECT 46.090 161.725 46.230 163.105 ;
        RECT 45.110 161.405 45.370 161.725 ;
        RECT 46.030 161.405 46.290 161.725 ;
        RECT 45.170 160.705 45.310 161.405 ;
        RECT 45.110 160.385 45.370 160.705 ;
        RECT 45.170 159.345 45.310 160.385 ;
        RECT 45.110 159.025 45.370 159.345 ;
        RECT 45.170 158.665 45.310 159.025 ;
        RECT 46.940 158.830 47.220 159.200 ;
        RECT 47.470 159.005 47.610 169.565 ;
        RECT 55.290 169.205 55.430 171.265 ;
        RECT 56.210 169.885 56.350 171.945 ;
        RECT 56.150 169.565 56.410 169.885 ;
        RECT 49.710 168.885 49.970 169.205 ;
        RECT 54.770 168.885 55.030 169.205 ;
        RECT 55.230 168.885 55.490 169.205 ;
        RECT 49.770 167.845 49.910 168.885 ;
        RECT 49.710 167.525 49.970 167.845 ;
        RECT 47.870 165.825 48.130 166.145 ;
        RECT 47.930 164.105 48.070 165.825 ;
        RECT 49.910 165.290 51.790 165.660 ;
        RECT 54.830 165.125 54.970 168.885 ;
        RECT 56.210 168.865 56.350 169.565 ;
        RECT 56.150 168.545 56.410 168.865 ;
        RECT 55.690 166.845 55.950 167.165 ;
        RECT 54.770 164.805 55.030 165.125 ;
        RECT 55.750 164.105 55.890 166.845 ;
        RECT 47.870 163.785 48.130 164.105 ;
        RECT 55.690 163.785 55.950 164.105 ;
        RECT 47.870 161.405 48.130 161.725 ;
        RECT 47.010 158.665 47.150 158.830 ;
        RECT 47.410 158.685 47.670 159.005 ;
        RECT 45.110 158.345 45.370 158.665 ;
        RECT 46.950 158.345 47.210 158.665 ;
        RECT 46.490 157.665 46.750 157.985 ;
        RECT 46.550 153.565 46.690 157.665 ;
        RECT 46.490 153.245 46.750 153.565 ;
        RECT 44.190 150.525 44.450 150.845 ;
        RECT 44.650 150.525 44.910 150.845 ;
        RECT 45.110 150.185 45.370 150.505 ;
        RECT 45.570 150.185 45.830 150.505 ;
        RECT 44.650 149.505 44.910 149.825 ;
        RECT 44.190 141.345 44.450 141.665 ;
        RECT 44.250 140.305 44.390 141.345 ;
        RECT 44.190 139.985 44.450 140.305 ;
        RECT 43.730 139.645 43.990 139.965 ;
        RECT 43.270 132.165 43.530 132.485 ;
        RECT 43.270 131.145 43.530 131.465 ;
        RECT 42.350 126.725 42.610 127.045 ;
        RECT 41.890 125.705 42.150 126.025 ;
        RECT 43.330 123.645 43.470 131.145 ;
        RECT 43.730 125.705 43.990 126.025 ;
        RECT 43.270 123.325 43.530 123.645 ;
        RECT 41.880 120.070 42.160 120.440 ;
        RECT 41.950 118.545 42.090 120.070 ;
        RECT 41.890 118.225 42.150 118.545 ;
        RECT 43.790 115.145 43.930 125.705 ;
        RECT 44.190 125.025 44.450 125.345 ;
        RECT 44.250 123.985 44.390 125.025 ;
        RECT 44.190 123.665 44.450 123.985 ;
        RECT 43.730 114.825 43.990 115.145 ;
        RECT 44.710 109.705 44.850 149.505 ;
        RECT 45.170 148.465 45.310 150.185 ;
        RECT 45.110 148.145 45.370 148.465 ;
        RECT 45.630 147.785 45.770 150.185 ;
        RECT 46.550 147.785 46.690 153.245 ;
        RECT 47.410 151.205 47.670 151.525 ;
        RECT 45.570 147.465 45.830 147.785 ;
        RECT 46.490 147.465 46.750 147.785 ;
        RECT 46.550 146.085 46.690 147.465 ;
        RECT 46.490 145.765 46.750 146.085 ;
        RECT 46.030 144.745 46.290 145.065 ;
        RECT 46.090 142.345 46.230 144.745 ;
        RECT 45.110 142.025 45.370 142.345 ;
        RECT 46.030 142.025 46.290 142.345 ;
        RECT 46.490 142.025 46.750 142.345 ;
        RECT 45.170 139.965 45.310 142.025 ;
        RECT 45.110 139.645 45.370 139.965 ;
        RECT 45.570 139.645 45.830 139.965 ;
        RECT 45.630 136.565 45.770 139.645 ;
        RECT 46.090 136.905 46.230 142.025 ;
        RECT 46.550 139.965 46.690 142.025 ;
        RECT 46.490 139.645 46.750 139.965 ;
        RECT 46.030 136.585 46.290 136.905 ;
        RECT 45.570 136.245 45.830 136.565 ;
        RECT 45.110 135.905 45.370 136.225 ;
        RECT 45.170 131.805 45.310 135.905 ;
        RECT 46.950 134.205 47.210 134.525 ;
        RECT 47.010 133.505 47.150 134.205 ;
        RECT 46.950 133.185 47.210 133.505 ;
        RECT 45.110 131.485 45.370 131.805 ;
        RECT 46.950 130.805 47.210 131.125 ;
        RECT 47.010 129.765 47.150 130.805 ;
        RECT 46.950 129.445 47.210 129.765 ;
        RECT 47.470 112.765 47.610 151.205 ;
        RECT 47.930 148.465 48.070 161.405 ;
        RECT 52.010 160.385 52.270 160.705 ;
        RECT 52.470 160.385 52.730 160.705 ;
        RECT 49.910 159.850 51.790 160.220 ;
        RECT 52.070 158.325 52.210 160.385 ;
        RECT 52.530 159.685 52.670 160.385 ;
        RECT 52.470 159.365 52.730 159.685 ;
        RECT 56.210 158.665 56.350 168.545 ;
        RECT 56.670 164.445 56.810 174.585 ;
        RECT 57.530 173.985 57.790 174.305 ;
        RECT 57.590 172.945 57.730 173.985 ;
        RECT 57.530 172.625 57.790 172.945 ;
        RECT 58.050 170.645 58.190 177.725 ;
        RECT 59.430 177.705 59.570 194.045 ;
        RECT 60.350 192.325 60.490 196.765 ;
        RECT 63.110 196.745 63.250 198.465 ;
        RECT 61.210 196.425 61.470 196.745 ;
        RECT 63.050 196.425 63.310 196.745 ;
        RECT 63.510 196.600 63.770 196.745 ;
        RECT 60.750 196.085 61.010 196.405 ;
        RECT 60.810 194.365 60.950 196.085 ;
        RECT 61.270 195.045 61.410 196.425 ;
        RECT 63.500 196.230 63.780 196.600 ;
        RECT 61.210 194.725 61.470 195.045 ;
        RECT 63.570 194.365 63.710 196.230 ;
        RECT 64.030 195.045 64.170 199.145 ;
        RECT 64.490 197.765 64.630 201.185 ;
        RECT 64.910 200.650 66.790 201.020 ;
        RECT 65.350 200.165 65.610 200.485 ;
        RECT 64.890 199.485 65.150 199.805 ;
        RECT 64.430 197.445 64.690 197.765 ;
        RECT 64.950 197.165 65.090 199.485 ;
        RECT 64.490 197.025 65.090 197.165 ;
        RECT 63.970 194.725 64.230 195.045 ;
        RECT 64.490 194.365 64.630 197.025 ;
        RECT 65.410 196.065 65.550 200.165 ;
        RECT 68.110 199.145 68.370 199.465 ;
        RECT 67.190 198.465 67.450 198.785 ;
        RECT 65.810 196.765 66.070 197.085 ;
        RECT 65.870 196.405 66.010 196.765 ;
        RECT 66.270 196.600 66.530 196.745 ;
        RECT 65.810 196.085 66.070 196.405 ;
        RECT 66.260 196.230 66.540 196.600 ;
        RECT 65.350 195.745 65.610 196.065 ;
        RECT 64.910 195.210 66.790 195.580 ;
        RECT 67.250 194.705 67.390 198.465 ;
        RECT 68.170 196.745 68.310 199.145 ;
        RECT 69.490 198.805 69.750 199.125 ;
        RECT 69.550 196.745 69.690 198.805 ;
        RECT 71.390 197.765 71.530 201.525 ;
        RECT 71.330 197.445 71.590 197.765 ;
        RECT 71.330 196.765 71.590 197.085 ;
        RECT 68.110 196.425 68.370 196.745 ;
        RECT 69.490 196.425 69.750 196.745 ;
        RECT 67.650 195.745 67.910 196.065 ;
        RECT 67.710 195.045 67.850 195.745 ;
        RECT 67.650 194.725 67.910 195.045 ;
        RECT 67.190 194.385 67.450 194.705 ;
        RECT 60.750 194.045 61.010 194.365 ;
        RECT 61.670 194.045 61.930 194.365 ;
        RECT 63.510 194.045 63.770 194.365 ;
        RECT 63.970 194.045 64.230 194.365 ;
        RECT 64.430 194.045 64.690 194.365 ;
        RECT 60.290 192.005 60.550 192.325 ;
        RECT 60.290 190.645 60.550 190.965 ;
        RECT 59.830 186.225 60.090 186.545 ;
        RECT 59.890 183.485 60.030 186.225 ;
        RECT 60.350 185.865 60.490 190.645 ;
        RECT 60.810 190.625 60.950 194.045 ;
        RECT 61.730 191.305 61.870 194.045 ;
        RECT 62.590 193.365 62.850 193.685 ;
        RECT 61.670 190.985 61.930 191.305 ;
        RECT 60.750 190.305 61.010 190.625 ;
        RECT 61.210 190.305 61.470 190.625 ;
        RECT 60.810 186.545 60.950 190.305 ;
        RECT 60.750 186.225 61.010 186.545 ;
        RECT 60.290 185.545 60.550 185.865 ;
        RECT 59.830 183.165 60.090 183.485 ;
        RECT 59.890 181.445 60.030 183.165 ;
        RECT 60.350 182.805 60.490 185.545 ;
        RECT 60.750 185.205 61.010 185.525 ;
        RECT 60.290 182.485 60.550 182.805 ;
        RECT 59.830 181.125 60.090 181.445 ;
        RECT 60.350 181.105 60.490 182.485 ;
        RECT 60.290 180.785 60.550 181.105 ;
        RECT 59.370 177.385 59.630 177.705 ;
        RECT 58.050 170.505 58.650 170.645 ;
        RECT 57.530 168.885 57.790 169.205 ;
        RECT 56.610 164.125 56.870 164.445 ;
        RECT 54.770 158.345 55.030 158.665 ;
        RECT 56.150 158.345 56.410 158.665 ;
        RECT 52.010 158.005 52.270 158.325 ;
        RECT 54.830 156.965 54.970 158.345 ;
        RECT 54.770 156.645 55.030 156.965 ;
        RECT 55.230 156.645 55.490 156.965 ;
        RECT 52.470 156.305 52.730 156.625 ;
        RECT 48.790 155.965 49.050 156.285 ;
        RECT 48.850 154.245 48.990 155.965 ;
        RECT 52.010 154.945 52.270 155.265 ;
        RECT 49.910 154.410 51.790 154.780 ;
        RECT 48.790 153.925 49.050 154.245 ;
        RECT 51.550 153.245 51.810 153.565 ;
        RECT 48.790 152.225 49.050 152.545 ;
        RECT 48.850 150.845 48.990 152.225 ;
        RECT 51.610 151.185 51.750 153.245 ;
        RECT 52.070 152.545 52.210 154.945 ;
        RECT 52.010 152.225 52.270 152.545 ;
        RECT 52.530 151.525 52.670 156.305 ;
        RECT 54.310 155.625 54.570 155.945 ;
        RECT 52.930 152.225 53.190 152.545 ;
        RECT 52.470 151.205 52.730 151.525 ;
        RECT 49.250 150.865 49.510 151.185 ;
        RECT 51.550 150.865 51.810 151.185 ;
        RECT 48.330 150.525 48.590 150.845 ;
        RECT 48.790 150.525 49.050 150.845 ;
        RECT 47.870 148.145 48.130 148.465 ;
        RECT 48.390 148.125 48.530 150.525 ;
        RECT 48.790 149.845 49.050 150.165 ;
        RECT 48.330 147.805 48.590 148.125 ;
        RECT 48.850 145.745 48.990 149.845 ;
        RECT 48.790 145.425 49.050 145.745 ;
        RECT 47.870 144.745 48.130 145.065 ;
        RECT 47.930 139.625 48.070 144.745 ;
        RECT 48.850 142.345 48.990 145.425 ;
        RECT 49.310 145.405 49.450 150.865 ;
        RECT 52.990 150.845 53.130 152.225 ;
        RECT 54.370 151.525 54.510 155.625 ;
        RECT 55.290 154.325 55.430 156.645 ;
        RECT 54.830 154.185 55.430 154.325 ;
        RECT 54.310 151.205 54.570 151.525 ;
        RECT 52.470 150.525 52.730 150.845 ;
        RECT 52.930 150.525 53.190 150.845 ;
        RECT 52.010 149.845 52.270 150.165 ;
        RECT 49.910 148.970 51.790 149.340 ;
        RECT 52.070 147.785 52.210 149.845 ;
        RECT 52.530 148.465 52.670 150.525 ;
        RECT 52.470 148.145 52.730 148.465 ;
        RECT 50.170 147.465 50.430 147.785 ;
        RECT 50.630 147.640 50.890 147.785 ;
        RECT 50.230 145.745 50.370 147.465 ;
        RECT 50.620 147.270 50.900 147.640 ;
        RECT 52.010 147.465 52.270 147.785 ;
        RECT 50.170 145.425 50.430 145.745 ;
        RECT 49.250 145.085 49.510 145.405 ;
        RECT 50.690 144.295 50.830 147.270 ;
        RECT 49.310 144.155 50.830 144.295 ;
        RECT 48.790 142.025 49.050 142.345 ;
        RECT 48.850 140.305 48.990 142.025 ;
        RECT 49.310 142.005 49.450 144.155 ;
        RECT 49.910 143.530 51.790 143.900 ;
        RECT 52.070 142.345 52.210 147.465 ;
        RECT 52.530 145.405 52.670 148.145 ;
        RECT 53.850 147.125 54.110 147.445 ;
        RECT 53.910 146.085 54.050 147.125 ;
        RECT 53.850 145.765 54.110 146.085 ;
        RECT 52.470 145.085 52.730 145.405 ;
        RECT 52.530 142.345 52.670 145.085 ;
        RECT 54.830 144.385 54.970 154.185 ;
        RECT 55.230 153.585 55.490 153.905 ;
        RECT 54.770 144.065 55.030 144.385 ;
        RECT 52.010 142.025 52.270 142.345 ;
        RECT 52.470 142.025 52.730 142.345 ;
        RECT 54.830 142.085 54.970 144.065 ;
        RECT 49.250 141.685 49.510 142.005 ;
        RECT 54.370 141.945 54.970 142.085 ;
        RECT 48.790 139.985 49.050 140.305 ;
        RECT 49.310 139.965 49.450 141.685 ;
        RECT 49.250 139.645 49.510 139.965 ;
        RECT 47.870 139.305 48.130 139.625 ;
        RECT 47.930 137.245 48.070 139.305 ;
        RECT 53.390 138.965 53.650 139.285 ;
        RECT 49.910 138.090 51.790 138.460 ;
        RECT 53.450 137.925 53.590 138.965 ;
        RECT 53.390 137.605 53.650 137.925 ;
        RECT 47.870 136.925 48.130 137.245 ;
        RECT 47.930 128.745 48.070 136.925 ;
        RECT 54.370 136.905 54.510 141.945 ;
        RECT 54.770 141.345 55.030 141.665 ;
        RECT 54.830 139.965 54.970 141.345 ;
        RECT 54.770 139.645 55.030 139.965 ;
        RECT 55.290 137.925 55.430 153.585 ;
        RECT 56.150 152.225 56.410 152.545 ;
        RECT 56.210 148.125 56.350 152.225 ;
        RECT 57.070 149.680 57.330 149.825 ;
        RECT 57.060 149.310 57.340 149.680 ;
        RECT 56.150 147.805 56.410 148.125 ;
        RECT 56.210 146.085 56.350 147.805 ;
        RECT 57.070 146.785 57.330 147.105 ;
        RECT 56.150 145.765 56.410 146.085 ;
        RECT 56.610 145.085 56.870 145.405 ;
        RECT 56.670 140.645 56.810 145.085 ;
        RECT 56.610 140.325 56.870 140.645 ;
        RECT 55.690 139.645 55.950 139.965 ;
        RECT 55.230 137.605 55.490 137.925 ;
        RECT 54.770 137.265 55.030 137.585 ;
        RECT 54.830 136.905 54.970 137.265 ;
        RECT 55.290 136.905 55.430 137.605 ;
        RECT 55.750 136.905 55.890 139.645 ;
        RECT 51.550 136.760 51.810 136.905 ;
        RECT 48.790 136.245 49.050 136.565 ;
        RECT 49.240 136.390 49.520 136.760 ;
        RECT 51.540 136.390 51.820 136.760 ;
        RECT 52.470 136.585 52.730 136.905 ;
        RECT 54.310 136.585 54.570 136.905 ;
        RECT 54.770 136.585 55.030 136.905 ;
        RECT 55.230 136.760 55.490 136.905 ;
        RECT 48.330 133.865 48.590 134.185 ;
        RECT 48.390 128.745 48.530 133.865 ;
        RECT 48.850 132.485 48.990 136.245 ;
        RECT 49.310 134.525 49.450 136.390 ;
        RECT 51.090 135.905 51.350 136.225 ;
        RECT 51.150 135.205 51.290 135.905 ;
        RECT 51.090 134.885 51.350 135.205 ;
        RECT 52.010 134.545 52.270 134.865 ;
        RECT 49.250 134.205 49.510 134.525 ;
        RECT 49.910 132.650 51.790 133.020 ;
        RECT 48.790 132.165 49.050 132.485 ;
        RECT 48.850 129.765 48.990 132.165 ;
        RECT 48.790 129.445 49.050 129.765 ;
        RECT 47.870 128.425 48.130 128.745 ;
        RECT 48.330 128.425 48.590 128.745 ;
        RECT 47.930 125.345 48.070 128.425 ;
        RECT 48.390 127.045 48.530 128.425 ;
        RECT 49.910 127.210 51.790 127.580 ;
        RECT 48.330 126.725 48.590 127.045 ;
        RECT 47.870 125.025 48.130 125.345 ;
        RECT 48.390 124.325 48.530 126.725 ;
        RECT 48.330 124.005 48.590 124.325 ;
        RECT 52.070 123.985 52.210 134.545 ;
        RECT 52.010 123.665 52.270 123.985 ;
        RECT 49.250 123.325 49.510 123.645 ;
        RECT 48.330 122.985 48.590 123.305 ;
        RECT 48.390 120.585 48.530 122.985 ;
        RECT 48.330 120.265 48.590 120.585 ;
        RECT 48.390 118.885 48.530 120.265 ;
        RECT 49.310 118.885 49.450 123.325 ;
        RECT 49.910 121.770 51.790 122.140 ;
        RECT 52.530 121.605 52.670 136.585 ;
        RECT 55.220 136.390 55.500 136.760 ;
        RECT 55.690 136.585 55.950 136.905 ;
        RECT 52.930 135.905 53.190 136.225 ;
        RECT 52.990 134.525 53.130 135.905 ;
        RECT 55.750 134.865 55.890 136.585 ;
        RECT 56.610 135.905 56.870 136.225 ;
        RECT 56.670 135.205 56.810 135.905 ;
        RECT 56.610 134.885 56.870 135.205 ;
        RECT 55.690 134.545 55.950 134.865 ;
        RECT 52.930 134.205 53.190 134.525 ;
        RECT 53.850 129.445 54.110 129.765 ;
        RECT 53.910 129.085 54.050 129.445 ;
        RECT 53.850 128.765 54.110 129.085 ;
        RECT 52.470 121.285 52.730 121.605 ;
        RECT 53.910 120.585 54.050 128.765 ;
        RECT 54.310 127.745 54.570 128.065 ;
        RECT 54.370 125.685 54.510 127.745 ;
        RECT 54.310 125.365 54.570 125.685 ;
        RECT 54.770 125.025 55.030 125.345 ;
        RECT 54.830 123.305 54.970 125.025 ;
        RECT 56.610 123.665 56.870 123.985 ;
        RECT 54.770 122.985 55.030 123.305 ;
        RECT 55.230 122.305 55.490 122.625 ;
        RECT 53.850 120.265 54.110 120.585 ;
        RECT 48.330 118.565 48.590 118.885 ;
        RECT 49.250 118.565 49.510 118.885 ;
        RECT 49.910 116.330 51.790 116.700 ;
        RECT 53.910 115.145 54.050 120.265 ;
        RECT 55.290 118.205 55.430 122.305 ;
        RECT 56.670 121.605 56.810 123.665 ;
        RECT 56.610 121.285 56.870 121.605 ;
        RECT 57.130 121.005 57.270 146.785 ;
        RECT 57.590 136.905 57.730 168.885 ;
        RECT 58.510 163.425 58.650 170.505 ;
        RECT 60.810 167.165 60.950 185.205 ;
        RECT 60.750 166.845 61.010 167.165 ;
        RECT 59.370 163.785 59.630 164.105 ;
        RECT 58.450 163.105 58.710 163.425 ;
        RECT 57.990 161.405 58.250 161.725 ;
        RECT 58.050 159.005 58.190 161.405 ;
        RECT 57.990 158.685 58.250 159.005 ;
        RECT 57.990 152.905 58.250 153.225 ;
        RECT 58.050 146.085 58.190 152.905 ;
        RECT 57.990 145.765 58.250 146.085 ;
        RECT 58.510 136.905 58.650 163.105 ;
        RECT 59.430 159.685 59.570 163.785 ;
        RECT 60.290 161.635 60.550 161.725 ;
        RECT 60.810 161.635 60.950 166.845 ;
        RECT 61.270 163.335 61.410 190.305 ;
        RECT 61.730 185.525 61.870 190.985 ;
        RECT 61.670 185.205 61.930 185.525 ;
        RECT 61.730 183.145 61.870 185.205 ;
        RECT 61.670 182.825 61.930 183.145 ;
        RECT 62.130 183.000 62.390 183.145 ;
        RECT 61.730 180.765 61.870 182.825 ;
        RECT 62.120 182.630 62.400 183.000 ;
        RECT 62.130 181.125 62.390 181.445 ;
        RECT 62.190 180.765 62.330 181.125 ;
        RECT 61.670 180.445 61.930 180.765 ;
        RECT 62.130 180.445 62.390 180.765 ;
        RECT 61.670 179.765 61.930 180.085 ;
        RECT 61.730 178.725 61.870 179.765 ;
        RECT 61.670 178.405 61.930 178.725 ;
        RECT 61.670 176.705 61.930 177.025 ;
        RECT 61.730 174.985 61.870 176.705 ;
        RECT 61.670 174.665 61.930 174.985 ;
        RECT 62.650 174.725 62.790 193.365 ;
        RECT 63.050 193.025 63.310 193.345 ;
        RECT 63.110 183.485 63.250 193.025 ;
        RECT 64.030 192.325 64.170 194.045 ;
        RECT 66.270 193.365 66.530 193.685 ;
        RECT 63.970 192.005 64.230 192.325 ;
        RECT 66.330 191.305 66.470 193.365 ;
        RECT 67.250 191.645 67.390 194.385 ;
        RECT 67.650 193.935 67.910 194.025 ;
        RECT 68.170 193.935 68.310 196.425 ;
        RECT 69.030 196.085 69.290 196.405 ;
        RECT 69.090 194.705 69.230 196.085 ;
        RECT 69.030 194.385 69.290 194.705 ;
        RECT 67.650 193.795 68.310 193.935 ;
        RECT 67.650 193.705 67.910 193.795 ;
        RECT 67.190 191.325 67.450 191.645 ;
        RECT 66.270 190.985 66.530 191.305 ;
        RECT 64.910 189.770 66.790 190.140 ;
        RECT 67.250 189.265 67.390 191.325 ;
        RECT 67.710 190.965 67.850 193.705 ;
        RECT 69.550 191.985 69.690 196.425 ;
        RECT 71.390 194.705 71.530 196.765 ;
        RECT 71.790 195.745 72.050 196.065 ;
        RECT 71.330 194.385 71.590 194.705 ;
        RECT 69.950 194.045 70.210 194.365 ;
        RECT 69.490 191.665 69.750 191.985 ;
        RECT 67.650 190.645 67.910 190.965 ;
        RECT 69.030 190.645 69.290 190.965 ;
        RECT 67.190 188.945 67.450 189.265 ;
        RECT 67.190 187.585 67.450 187.905 ;
        RECT 64.910 184.330 66.790 184.700 ;
        RECT 63.970 183.505 64.230 183.825 ;
        RECT 63.050 183.165 63.310 183.485 ;
        RECT 63.110 181.105 63.250 183.165 ;
        RECT 63.050 180.785 63.310 181.105 ;
        RECT 63.510 180.445 63.770 180.765 ;
        RECT 63.050 178.065 63.310 178.385 ;
        RECT 62.190 174.585 62.790 174.725 ;
        RECT 61.670 173.985 61.930 174.305 ;
        RECT 61.730 172.945 61.870 173.985 ;
        RECT 61.670 172.625 61.930 172.945 ;
        RECT 61.670 167.185 61.930 167.505 ;
        RECT 61.730 164.105 61.870 167.185 ;
        RECT 62.190 166.485 62.330 174.585 ;
        RECT 62.590 173.985 62.850 174.305 ;
        RECT 62.650 173.285 62.790 173.985 ;
        RECT 62.590 172.965 62.850 173.285 ;
        RECT 63.110 166.825 63.250 178.065 ;
        RECT 63.570 177.705 63.710 180.445 ;
        RECT 63.510 177.385 63.770 177.705 ;
        RECT 63.570 177.025 63.710 177.385 ;
        RECT 63.510 176.705 63.770 177.025 ;
        RECT 63.510 174.665 63.770 174.985 ;
        RECT 63.570 169.545 63.710 174.665 ;
        RECT 63.510 169.225 63.770 169.545 ;
        RECT 63.050 166.505 63.310 166.825 ;
        RECT 62.130 166.165 62.390 166.485 ;
        RECT 61.670 163.785 61.930 164.105 ;
        RECT 61.270 163.195 61.870 163.335 ;
        RECT 61.210 161.635 61.470 161.725 ;
        RECT 60.290 161.495 61.470 161.635 ;
        RECT 60.290 161.405 60.550 161.495 ;
        RECT 61.210 161.405 61.470 161.495 ;
        RECT 60.290 160.725 60.550 161.045 ;
        RECT 59.370 159.365 59.630 159.685 ;
        RECT 59.430 158.665 59.570 159.365 ;
        RECT 59.370 158.345 59.630 158.665 ;
        RECT 58.910 152.225 59.170 152.545 ;
        RECT 59.830 152.225 60.090 152.545 ;
        RECT 58.970 148.125 59.110 152.225 ;
        RECT 59.890 150.165 60.030 152.225 ;
        RECT 60.350 151.040 60.490 160.725 ;
        RECT 61.210 158.005 61.470 158.325 ;
        RECT 61.270 155.945 61.410 158.005 ;
        RECT 61.210 155.625 61.470 155.945 ;
        RECT 60.280 150.670 60.560 151.040 ;
        RECT 59.830 149.845 60.090 150.165 ;
        RECT 59.890 148.805 60.030 149.845 ;
        RECT 59.830 148.485 60.090 148.805 ;
        RECT 61.270 148.125 61.410 155.625 ;
        RECT 61.730 154.325 61.870 163.195 ;
        RECT 62.190 161.725 62.330 166.165 ;
        RECT 62.130 161.405 62.390 161.725 ;
        RECT 62.120 158.830 62.400 159.200 ;
        RECT 62.190 156.965 62.330 158.830 ;
        RECT 62.590 158.345 62.850 158.665 ;
        RECT 62.130 156.645 62.390 156.965 ;
        RECT 62.650 156.285 62.790 158.345 ;
        RECT 62.590 155.965 62.850 156.285 ;
        RECT 61.730 154.185 62.330 154.325 ;
        RECT 62.190 153.905 62.330 154.185 ;
        RECT 62.130 153.585 62.390 153.905 ;
        RECT 58.910 147.805 59.170 148.125 ;
        RECT 61.210 147.805 61.470 148.125 ;
        RECT 62.190 145.405 62.330 153.585 ;
        RECT 62.650 152.545 62.790 155.965 ;
        RECT 63.110 152.545 63.250 166.505 ;
        RECT 63.570 166.145 63.710 169.225 ;
        RECT 63.510 165.825 63.770 166.145 ;
        RECT 63.570 158.665 63.710 165.825 ;
        RECT 63.510 158.345 63.770 158.665 ;
        RECT 63.510 157.665 63.770 157.985 ;
        RECT 63.570 156.625 63.710 157.665 ;
        RECT 63.510 156.305 63.770 156.625 ;
        RECT 64.030 156.285 64.170 183.505 ;
        RECT 67.250 183.485 67.390 187.585 ;
        RECT 69.090 183.825 69.230 190.645 ;
        RECT 70.010 187.905 70.150 194.045 ;
        RECT 70.870 193.705 71.130 194.025 ;
        RECT 70.410 190.305 70.670 190.625 ;
        RECT 70.470 189.265 70.610 190.305 ;
        RECT 70.930 189.605 71.070 193.705 ;
        RECT 71.850 191.645 71.990 195.745 ;
        RECT 73.690 195.045 73.830 201.525 ;
        RECT 75.010 201.185 75.270 201.505 ;
        RECT 75.070 200.145 75.210 201.185 ;
        RECT 75.010 199.825 75.270 200.145 ;
        RECT 76.450 199.805 76.590 201.865 ;
        RECT 94.910 200.650 96.790 201.020 ;
        RECT 76.390 199.485 76.650 199.805 ;
        RECT 78.230 199.485 78.490 199.805 ;
        RECT 76.450 197.085 76.590 199.485 ;
        RECT 76.390 196.765 76.650 197.085 ;
        RECT 74.090 196.085 74.350 196.405 ;
        RECT 74.150 195.045 74.290 196.085 ;
        RECT 73.630 194.725 73.890 195.045 ;
        RECT 74.090 194.725 74.350 195.045 ;
        RECT 74.090 194.045 74.350 194.365 ;
        RECT 74.150 192.325 74.290 194.045 ;
        RECT 74.090 192.005 74.350 192.325 ;
        RECT 74.150 191.645 74.290 192.005 ;
        RECT 78.290 191.645 78.430 199.485 ;
        RECT 79.910 197.930 81.790 198.300 ;
        RECT 109.910 197.930 111.790 198.300 ;
        RECT 80.530 196.765 80.790 197.085 ;
        RECT 79.150 196.085 79.410 196.405 ;
        RECT 79.210 195.045 79.350 196.085 ;
        RECT 79.150 194.725 79.410 195.045 ;
        RECT 80.590 194.365 80.730 196.765 ;
        RECT 94.910 195.210 96.790 195.580 ;
        RECT 89.270 194.385 89.530 194.705 ;
        RECT 80.530 194.045 80.790 194.365 ;
        RECT 86.510 194.045 86.770 194.365 ;
        RECT 79.910 192.490 81.790 192.860 ;
        RECT 71.790 191.325 72.050 191.645 ;
        RECT 74.090 191.325 74.350 191.645 ;
        RECT 78.230 191.325 78.490 191.645 ;
        RECT 81.450 191.215 81.710 191.305 ;
        RECT 81.450 191.075 82.110 191.215 ;
        RECT 81.450 190.985 81.710 191.075 ;
        RECT 76.390 190.645 76.650 190.965 ;
        RECT 76.450 189.605 76.590 190.645 ;
        RECT 80.990 190.305 81.250 190.625 ;
        RECT 70.870 189.285 71.130 189.605 ;
        RECT 76.390 189.285 76.650 189.605 ;
        RECT 70.410 188.945 70.670 189.265 ;
        RECT 69.950 187.585 70.210 187.905 ;
        RECT 69.030 183.505 69.290 183.825 ;
        RECT 64.890 183.165 65.150 183.485 ;
        RECT 67.190 183.165 67.450 183.485 ;
        RECT 67.650 183.165 67.910 183.485 ;
        RECT 64.950 182.805 65.090 183.165 ;
        RECT 64.890 182.485 65.150 182.805 ;
        RECT 67.710 181.445 67.850 183.165 ;
        RECT 70.930 182.805 71.070 189.285 ;
        RECT 81.050 189.265 81.190 190.305 ;
        RECT 73.630 188.945 73.890 189.265 ;
        RECT 80.990 188.945 81.250 189.265 ;
        RECT 73.170 188.265 73.430 188.585 ;
        RECT 73.230 183.145 73.370 188.265 ;
        RECT 73.690 185.185 73.830 188.945 ;
        RECT 78.230 188.605 78.490 188.925 ;
        RECT 78.290 187.905 78.430 188.605 ;
        RECT 75.930 187.585 76.190 187.905 ;
        RECT 78.230 187.585 78.490 187.905 ;
        RECT 73.630 184.865 73.890 185.185 ;
        RECT 73.690 184.165 73.830 184.865 ;
        RECT 73.630 183.845 73.890 184.165 ;
        RECT 73.170 182.825 73.430 183.145 ;
        RECT 70.870 182.485 71.130 182.805 ;
        RECT 73.170 182.145 73.430 182.465 ;
        RECT 67.650 181.125 67.910 181.445 ;
        RECT 69.950 179.765 70.210 180.085 ;
        RECT 64.430 179.425 64.690 179.745 ;
        RECT 67.190 179.425 67.450 179.745 ;
        RECT 69.490 179.425 69.750 179.745 ;
        RECT 64.490 174.985 64.630 179.425 ;
        RECT 64.910 178.890 66.790 179.260 ;
        RECT 67.250 178.725 67.390 179.425 ;
        RECT 64.890 178.405 65.150 178.725 ;
        RECT 67.190 178.405 67.450 178.725 ;
        RECT 64.950 175.665 65.090 178.405 ;
        RECT 69.550 178.045 69.690 179.425 ;
        RECT 69.490 177.725 69.750 178.045 ;
        RECT 70.010 177.365 70.150 179.765 ;
        RECT 72.250 179.425 72.510 179.745 ;
        RECT 69.950 177.045 70.210 177.365 ;
        RECT 68.110 176.705 68.370 177.025 ;
        RECT 68.170 176.005 68.310 176.705 ;
        RECT 68.110 175.685 68.370 176.005 ;
        RECT 71.790 175.685 72.050 176.005 ;
        RECT 64.890 175.345 65.150 175.665 ;
        RECT 68.170 174.985 68.310 175.685 ;
        RECT 68.560 175.150 68.840 175.520 ;
        RECT 71.330 175.345 71.590 175.665 ;
        RECT 68.630 174.985 68.770 175.150 ;
        RECT 71.390 174.985 71.530 175.345 ;
        RECT 71.850 174.985 71.990 175.685 ;
        RECT 72.310 174.985 72.450 179.425 ;
        RECT 73.230 178.045 73.370 182.145 ;
        RECT 73.170 177.725 73.430 178.045 ;
        RECT 72.700 175.150 72.980 175.520 ;
        RECT 72.710 175.005 72.970 175.150 ;
        RECT 64.430 174.665 64.690 174.985 ;
        RECT 68.110 174.665 68.370 174.985 ;
        RECT 68.570 174.665 68.830 174.985 ;
        RECT 71.330 174.665 71.590 174.985 ;
        RECT 71.790 174.665 72.050 174.985 ;
        RECT 72.250 174.665 72.510 174.985 ;
        RECT 64.430 173.985 64.690 174.305 ;
        RECT 69.490 173.985 69.750 174.305 ;
        RECT 63.970 155.965 64.230 156.285 ;
        RECT 64.030 155.125 64.170 155.965 ;
        RECT 63.570 154.985 64.170 155.125 ;
        RECT 63.570 153.565 63.710 154.985 ;
        RECT 63.510 153.245 63.770 153.565 ;
        RECT 62.590 152.225 62.850 152.545 ;
        RECT 63.050 152.225 63.310 152.545 ;
        RECT 62.130 145.085 62.390 145.405 ;
        RECT 62.590 141.685 62.850 142.005 ;
        RECT 62.650 140.645 62.790 141.685 ;
        RECT 62.590 140.325 62.850 140.645 ;
        RECT 60.750 139.305 61.010 139.625 ;
        RECT 60.290 138.625 60.550 138.945 ;
        RECT 57.530 136.815 57.790 136.905 ;
        RECT 57.530 136.675 58.190 136.815 ;
        RECT 57.530 136.585 57.790 136.675 ;
        RECT 58.050 135.205 58.190 136.675 ;
        RECT 58.450 136.585 58.710 136.905 ;
        RECT 57.990 134.885 58.250 135.205 ;
        RECT 58.510 129.765 58.650 136.585 ;
        RECT 59.370 135.905 59.630 136.225 ;
        RECT 59.430 134.865 59.570 135.905 ;
        RECT 59.370 134.545 59.630 134.865 ;
        RECT 58.450 129.445 58.710 129.765 ;
        RECT 57.990 127.745 58.250 128.065 ;
        RECT 58.050 126.365 58.190 127.745 ;
        RECT 57.990 126.045 58.250 126.365 ;
        RECT 59.830 123.325 60.090 123.645 ;
        RECT 56.670 120.865 57.270 121.005 ;
        RECT 55.230 117.885 55.490 118.205 ;
        RECT 53.850 114.825 54.110 115.145 ;
        RECT 53.910 113.105 54.050 114.825 ;
        RECT 53.850 112.785 54.110 113.105 ;
        RECT 47.410 112.445 47.670 112.765 ;
        RECT 52.010 112.105 52.270 112.425 ;
        RECT 49.910 110.890 51.790 111.260 ;
        RECT 48.790 109.725 49.050 110.045 ;
        RECT 40.970 109.385 41.230 109.705 ;
        RECT 44.650 109.385 44.910 109.705 ;
        RECT 46.030 109.045 46.290 109.365 ;
        RECT 40.050 108.705 40.310 109.025 ;
        RECT 40.110 107.665 40.250 108.705 ;
        RECT 46.090 108.005 46.230 109.045 ;
        RECT 47.870 108.705 48.130 109.025 ;
        RECT 46.030 107.685 46.290 108.005 ;
        RECT 40.050 107.345 40.310 107.665 ;
        RECT 44.190 107.345 44.450 107.665 ;
        RECT 36.370 106.685 37.490 106.825 ;
        RECT 36.370 106.665 36.630 106.685 ;
        RECT 38.210 106.665 38.470 106.985 ;
        RECT 43.270 106.825 43.530 106.985 ;
        RECT 43.270 106.685 43.930 106.825 ;
        RECT 43.270 106.665 43.530 106.685 ;
        RECT 36.430 104.605 36.570 106.665 ;
        RECT 34.530 104.285 34.790 104.605 ;
        RECT 36.370 104.285 36.630 104.605 ;
        RECT 34.910 102.730 36.790 103.100 ;
        RECT 38.270 92.050 38.410 106.665 ;
        RECT 43.790 92.050 43.930 106.685 ;
        RECT 44.250 105.285 44.390 107.345 ;
        RECT 44.190 104.965 44.450 105.285 ;
        RECT 46.090 104.265 46.230 107.685 ;
        RECT 47.930 107.665 48.070 108.705 ;
        RECT 47.870 107.345 48.130 107.665 ;
        RECT 48.850 104.515 48.990 109.725 ;
        RECT 49.250 109.385 49.510 109.705 ;
        RECT 49.310 105.285 49.450 109.385 ;
        RECT 51.550 108.765 51.810 109.025 ;
        RECT 52.070 108.765 52.210 112.105 ;
        RECT 54.770 111.425 55.030 111.745 ;
        RECT 54.830 110.045 54.970 111.425 ;
        RECT 54.770 109.725 55.030 110.045 ;
        RECT 56.670 109.705 56.810 120.865 ;
        RECT 59.370 119.585 59.630 119.905 ;
        RECT 57.070 118.225 57.330 118.545 ;
        RECT 57.130 116.165 57.270 118.225 ;
        RECT 57.070 115.845 57.330 116.165 ;
        RECT 59.430 110.045 59.570 119.585 ;
        RECT 59.890 118.885 60.030 123.325 ;
        RECT 59.830 118.565 60.090 118.885 ;
        RECT 59.370 109.725 59.630 110.045 ;
        RECT 56.610 109.385 56.870 109.705 ;
        RECT 51.550 108.705 52.210 108.765 ;
        RECT 57.990 108.705 58.250 109.025 ;
        RECT 58.910 108.705 59.170 109.025 ;
        RECT 51.610 108.625 52.210 108.705 ;
        RECT 49.910 105.450 51.790 105.820 ;
        RECT 49.250 104.965 49.510 105.285 ;
        RECT 48.850 104.375 49.450 104.515 ;
        RECT 46.030 103.945 46.290 104.265 ;
        RECT 49.310 92.050 49.450 104.375 ;
        RECT 52.070 104.265 52.210 108.625 ;
        RECT 52.470 107.345 52.730 107.665 ;
        RECT 52.530 105.285 52.670 107.345 ;
        RECT 58.050 106.985 58.190 108.705 ;
        RECT 54.770 106.665 55.030 106.985 ;
        RECT 57.990 106.665 58.250 106.985 ;
        RECT 52.470 104.965 52.730 105.285 ;
        RECT 52.010 103.945 52.270 104.265 ;
        RECT 54.830 92.050 54.970 106.665 ;
        RECT 58.970 103.925 59.110 108.705 ;
        RECT 59.430 108.005 59.570 109.725 ;
        RECT 60.350 109.705 60.490 138.625 ;
        RECT 60.810 136.905 60.950 139.305 ;
        RECT 63.110 136.905 63.250 152.225 ;
        RECT 63.510 150.525 63.770 150.845 ;
        RECT 63.570 150.360 63.710 150.525 ;
        RECT 63.500 149.990 63.780 150.360 ;
        RECT 64.490 148.125 64.630 173.985 ;
        RECT 64.910 173.450 66.790 173.820 ;
        RECT 67.650 169.565 67.910 169.885 ;
        RECT 64.910 168.010 66.790 168.380 ;
        RECT 67.710 167.845 67.850 169.565 ;
        RECT 67.650 167.525 67.910 167.845 ;
        RECT 64.910 162.570 66.790 162.940 ;
        RECT 67.190 157.665 67.450 157.985 ;
        RECT 64.910 157.130 66.790 157.500 ;
        RECT 65.810 153.585 66.070 153.905 ;
        RECT 66.270 153.585 66.530 153.905 ;
        RECT 65.870 153.225 66.010 153.585 ;
        RECT 65.810 152.905 66.070 153.225 ;
        RECT 66.330 152.545 66.470 153.585 ;
        RECT 66.270 152.225 66.530 152.545 ;
        RECT 64.910 151.690 66.790 152.060 ;
        RECT 67.250 150.925 67.390 157.665 ;
        RECT 67.710 156.965 67.850 167.525 ;
        RECT 69.030 161.065 69.290 161.385 ;
        RECT 69.090 158.665 69.230 161.065 ;
        RECT 69.030 158.345 69.290 158.665 ;
        RECT 68.570 157.665 68.830 157.985 ;
        RECT 67.650 156.645 67.910 156.965 ;
        RECT 68.630 156.625 68.770 157.665 ;
        RECT 68.570 156.305 68.830 156.625 ;
        RECT 69.090 156.285 69.230 158.345 ;
        RECT 69.030 155.965 69.290 156.285 ;
        RECT 68.110 154.945 68.370 155.265 ;
        RECT 69.030 154.945 69.290 155.265 ;
        RECT 67.650 152.565 67.910 152.885 ;
        RECT 66.790 150.785 67.390 150.925 ;
        RECT 66.790 148.125 66.930 150.785 ;
        RECT 67.190 148.485 67.450 148.805 ;
        RECT 64.430 147.805 64.690 148.125 ;
        RECT 66.730 147.805 66.990 148.125 ;
        RECT 63.970 146.785 64.230 147.105 ;
        RECT 63.510 142.025 63.770 142.345 ;
        RECT 60.750 136.585 61.010 136.905 ;
        RECT 63.050 136.585 63.310 136.905 ;
        RECT 61.670 136.245 61.930 136.565 ;
        RECT 61.730 131.805 61.870 136.245 ;
        RECT 63.570 134.185 63.710 142.025 ;
        RECT 63.510 133.865 63.770 134.185 ;
        RECT 61.670 131.485 61.930 131.805 ;
        RECT 61.730 110.725 61.870 131.485 ;
        RECT 63.050 130.465 63.310 130.785 ;
        RECT 63.110 129.425 63.250 130.465 ;
        RECT 63.050 129.105 63.310 129.425 ;
        RECT 63.570 126.365 63.710 133.865 ;
        RECT 63.510 126.045 63.770 126.365 ;
        RECT 63.570 120.925 63.710 126.045 ;
        RECT 63.510 120.605 63.770 120.925 ;
        RECT 63.570 119.905 63.710 120.605 ;
        RECT 63.510 119.585 63.770 119.905 ;
        RECT 61.670 110.405 61.930 110.725 ;
        RECT 64.030 109.705 64.170 146.785 ;
        RECT 64.910 146.250 66.790 146.620 ;
        RECT 64.910 140.810 66.790 141.180 ;
        RECT 64.430 135.905 64.690 136.225 ;
        RECT 64.490 134.525 64.630 135.905 ;
        RECT 64.910 135.370 66.790 135.740 ;
        RECT 64.430 134.205 64.690 134.525 ;
        RECT 67.250 132.485 67.390 148.485 ;
        RECT 67.710 139.965 67.850 152.565 ;
        RECT 68.170 142.345 68.310 154.945 ;
        RECT 68.570 152.225 68.830 152.545 ;
        RECT 68.630 151.185 68.770 152.225 ;
        RECT 68.570 150.865 68.830 151.185 ;
        RECT 69.090 150.845 69.230 154.945 ;
        RECT 69.030 150.525 69.290 150.845 ;
        RECT 68.570 149.680 68.830 149.825 ;
        RECT 68.560 149.310 68.840 149.680 ;
        RECT 68.570 147.640 68.830 147.785 ;
        RECT 68.560 147.270 68.840 147.640 ;
        RECT 68.630 147.105 68.770 147.270 ;
        RECT 68.570 146.785 68.830 147.105 ;
        RECT 69.030 144.065 69.290 144.385 ;
        RECT 68.570 143.045 68.830 143.365 ;
        RECT 68.110 142.025 68.370 142.345 ;
        RECT 68.110 141.345 68.370 141.665 ;
        RECT 67.650 139.645 67.910 139.965 ;
        RECT 67.650 138.625 67.910 138.945 ;
        RECT 67.190 132.165 67.450 132.485 ;
        RECT 64.880 131.630 65.160 132.000 ;
        RECT 64.950 131.465 65.090 131.630 ;
        RECT 64.890 131.145 65.150 131.465 ;
        RECT 64.910 129.930 66.790 130.300 ;
        RECT 64.910 124.490 66.790 124.860 ;
        RECT 65.350 122.305 65.610 122.625 ;
        RECT 65.410 120.585 65.550 122.305 ;
        RECT 65.350 120.265 65.610 120.585 ;
        RECT 64.910 119.050 66.790 119.420 ;
        RECT 64.910 113.610 66.790 113.980 ;
        RECT 67.710 113.445 67.850 138.625 ;
        RECT 67.650 113.125 67.910 113.445 ;
        RECT 68.170 112.425 68.310 141.345 ;
        RECT 68.630 132.485 68.770 143.045 ;
        RECT 69.090 139.285 69.230 144.065 ;
        RECT 69.550 142.685 69.690 173.985 ;
        RECT 71.390 172.605 71.530 174.665 ;
        RECT 71.850 172.945 71.990 174.665 ;
        RECT 72.250 173.985 72.510 174.305 ;
        RECT 71.790 172.625 72.050 172.945 ;
        RECT 71.330 172.285 71.590 172.605 ;
        RECT 71.330 171.265 71.590 171.585 ;
        RECT 69.950 166.845 70.210 167.165 ;
        RECT 70.010 164.445 70.150 166.845 ;
        RECT 69.950 164.125 70.210 164.445 ;
        RECT 70.010 158.665 70.150 164.125 ;
        RECT 70.870 162.085 71.130 162.405 ;
        RECT 70.930 160.705 71.070 162.085 ;
        RECT 70.410 160.385 70.670 160.705 ;
        RECT 70.870 160.385 71.130 160.705 ;
        RECT 70.470 159.005 70.610 160.385 ;
        RECT 70.410 158.685 70.670 159.005 ;
        RECT 69.950 158.345 70.210 158.665 ;
        RECT 70.470 156.285 70.610 158.685 ;
        RECT 69.950 155.965 70.210 156.285 ;
        RECT 70.410 156.195 70.670 156.285 ;
        RECT 70.410 156.055 71.070 156.195 ;
        RECT 70.410 155.965 70.670 156.055 ;
        RECT 70.010 153.225 70.150 155.965 ;
        RECT 70.410 153.925 70.670 154.245 ;
        RECT 69.950 152.905 70.210 153.225 ;
        RECT 70.470 152.455 70.610 153.925 ;
        RECT 70.930 153.225 71.070 156.055 ;
        RECT 70.870 152.905 71.130 153.225 ;
        RECT 70.470 152.315 71.070 152.455 ;
        RECT 70.410 150.525 70.670 150.845 ;
        RECT 69.950 149.505 70.210 149.825 ;
        RECT 69.490 142.365 69.750 142.685 ;
        RECT 69.030 138.965 69.290 139.285 ;
        RECT 69.090 137.585 69.230 138.965 ;
        RECT 69.030 137.265 69.290 137.585 ;
        RECT 70.010 134.185 70.150 149.505 ;
        RECT 70.470 148.805 70.610 150.525 ;
        RECT 70.410 148.485 70.670 148.805 ;
        RECT 70.410 147.695 70.670 147.785 ;
        RECT 70.930 147.695 71.070 152.315 ;
        RECT 70.410 147.555 71.070 147.695 ;
        RECT 70.410 147.465 70.670 147.555 ;
        RECT 70.470 145.745 70.610 147.465 ;
        RECT 70.410 145.425 70.670 145.745 ;
        RECT 70.470 142.345 70.610 145.425 ;
        RECT 70.410 142.025 70.670 142.345 ;
        RECT 70.470 139.965 70.610 142.025 ;
        RECT 70.870 141.685 71.130 142.005 ;
        RECT 70.930 139.965 71.070 141.685 ;
        RECT 70.410 139.645 70.670 139.965 ;
        RECT 70.870 139.645 71.130 139.965 ;
        RECT 71.390 139.285 71.530 171.265 ;
        RECT 71.790 163.445 72.050 163.765 ;
        RECT 71.850 162.405 71.990 163.445 ;
        RECT 71.790 162.085 72.050 162.405 ;
        RECT 71.790 159.200 72.050 159.345 ;
        RECT 71.780 158.830 72.060 159.200 ;
        RECT 71.790 158.005 72.050 158.325 ;
        RECT 71.850 156.285 71.990 158.005 ;
        RECT 71.790 155.965 72.050 156.285 ;
        RECT 71.850 153.225 71.990 155.965 ;
        RECT 71.790 152.905 72.050 153.225 ;
        RECT 72.310 150.505 72.450 173.985 ;
        RECT 73.230 172.605 73.370 177.725 ;
        RECT 73.690 175.325 73.830 183.845 ;
        RECT 74.090 183.165 74.350 183.485 ;
        RECT 74.150 178.725 74.290 183.165 ;
        RECT 75.010 182.825 75.270 183.145 ;
        RECT 75.070 180.425 75.210 182.825 ;
        RECT 75.010 180.105 75.270 180.425 ;
        RECT 74.090 178.405 74.350 178.725 ;
        RECT 75.070 177.705 75.210 180.105 ;
        RECT 75.010 177.385 75.270 177.705 ;
        RECT 73.630 175.005 73.890 175.325 ;
        RECT 75.990 174.985 76.130 187.585 ;
        RECT 79.910 187.050 81.790 187.420 ;
        RECT 81.450 186.115 81.710 186.205 ;
        RECT 81.970 186.115 82.110 191.075 ;
        RECT 84.670 190.305 84.930 190.625 ;
        RECT 84.730 188.925 84.870 190.305 ;
        RECT 86.570 188.925 86.710 194.045 ;
        RECT 89.330 192.325 89.470 194.385 ;
        RECT 102.610 194.045 102.870 194.365 ;
        RECT 103.530 194.045 103.790 194.365 ;
        RECT 92.490 193.705 92.750 194.025 ;
        RECT 89.270 192.005 89.530 192.325 ;
        RECT 90.650 190.305 90.910 190.625 ;
        RECT 90.710 189.265 90.850 190.305 ;
        RECT 92.550 189.605 92.690 193.705 ;
        RECT 97.550 193.025 97.810 193.345 ;
        RECT 102.150 193.025 102.410 193.345 ;
        RECT 97.610 191.305 97.750 193.025 ;
        RECT 98.470 191.325 98.730 191.645 ;
        RECT 97.550 190.985 97.810 191.305 ;
        RECT 94.910 189.770 96.790 190.140 ;
        RECT 92.490 189.285 92.750 189.605 ;
        RECT 90.650 188.945 90.910 189.265 ;
        RECT 84.670 188.605 84.930 188.925 ;
        RECT 86.510 188.605 86.770 188.925 ;
        RECT 86.570 186.205 86.710 188.605 ;
        RECT 92.490 187.585 92.750 187.905 ;
        RECT 81.450 185.975 82.110 186.115 ;
        RECT 81.450 185.885 81.710 185.975 ;
        RECT 80.530 185.545 80.790 185.865 ;
        RECT 80.590 184.165 80.730 185.545 ;
        RECT 80.530 183.845 80.790 184.165 ;
        RECT 81.970 183.145 82.110 185.975 ;
        RECT 83.290 185.885 83.550 186.205 ;
        RECT 86.510 185.885 86.770 186.205 ;
        RECT 83.350 183.825 83.490 185.885 ;
        RECT 83.290 183.505 83.550 183.825 ;
        RECT 81.910 182.825 82.170 183.145 ;
        RECT 79.910 181.610 81.790 181.980 ;
        RECT 79.150 180.445 79.410 180.765 ;
        RECT 79.210 175.325 79.350 180.445 ;
        RECT 81.450 179.765 81.710 180.085 ;
        RECT 81.510 178.725 81.650 179.765 ;
        RECT 81.450 178.405 81.710 178.725 ;
        RECT 81.970 178.045 82.110 182.825 ;
        RECT 83.350 180.765 83.490 183.505 ;
        RECT 86.050 183.165 86.310 183.485 ;
        RECT 85.590 182.145 85.850 182.465 ;
        RECT 83.290 180.445 83.550 180.765 ;
        RECT 81.910 177.725 82.170 178.045 ;
        RECT 79.910 176.170 81.790 176.540 ;
        RECT 79.150 175.005 79.410 175.325 ;
        RECT 75.930 174.665 76.190 174.985 ;
        RECT 74.090 174.325 74.350 174.645 ;
        RECT 78.230 174.325 78.490 174.645 ;
        RECT 81.450 174.325 81.710 174.645 ;
        RECT 74.150 172.605 74.290 174.325 ;
        RECT 78.290 172.800 78.430 174.325 ;
        RECT 81.510 173.285 81.650 174.325 ;
        RECT 81.450 172.965 81.710 173.285 ;
        RECT 73.170 172.285 73.430 172.605 ;
        RECT 74.090 172.285 74.350 172.605 ;
        RECT 78.220 172.430 78.500 172.800 ;
        RECT 81.970 172.605 82.110 177.725 ;
        RECT 83.350 176.005 83.490 180.445 ;
        RECT 84.670 180.105 84.930 180.425 ;
        RECT 84.730 178.385 84.870 180.105 ;
        RECT 85.650 178.385 85.790 182.145 ;
        RECT 86.110 181.525 86.250 183.165 ;
        RECT 86.570 183.145 86.710 185.885 ;
        RECT 91.110 185.205 91.370 185.525 ;
        RECT 91.570 185.205 91.830 185.525 ;
        RECT 86.510 182.825 86.770 183.145 ;
        RECT 89.270 182.145 89.530 182.465 ;
        RECT 86.110 181.445 86.710 181.525 ;
        RECT 86.110 181.385 86.770 181.445 ;
        RECT 86.510 181.125 86.770 181.385 ;
        RECT 86.050 179.425 86.310 179.745 ;
        RECT 86.110 178.725 86.250 179.425 ;
        RECT 86.050 178.405 86.310 178.725 ;
        RECT 84.670 178.065 84.930 178.385 ;
        RECT 85.590 178.065 85.850 178.385 ;
        RECT 86.510 176.705 86.770 177.025 ;
        RECT 83.290 175.685 83.550 176.005 ;
        RECT 83.350 172.685 83.490 175.685 ;
        RECT 83.750 175.345 84.010 175.665 ;
        RECT 82.890 172.605 83.490 172.685 ;
        RECT 81.910 172.285 82.170 172.605 ;
        RECT 82.830 172.545 83.490 172.605 ;
        RECT 82.830 172.285 83.090 172.545 ;
        RECT 79.910 170.730 81.790 171.100 ;
        RECT 83.350 169.885 83.490 172.545 ;
        RECT 83.810 170.565 83.950 175.345 ;
        RECT 86.570 174.985 86.710 176.705 ;
        RECT 89.330 176.005 89.470 182.145 ;
        RECT 91.170 180.425 91.310 185.205 ;
        RECT 91.630 181.445 91.770 185.205 ;
        RECT 92.550 182.465 92.690 187.585 ;
        RECT 93.410 184.865 93.670 185.185 ;
        RECT 93.470 184.165 93.610 184.865 ;
        RECT 94.910 184.330 96.790 184.700 ;
        RECT 93.410 183.845 93.670 184.165 ;
        RECT 92.490 182.145 92.750 182.465 ;
        RECT 91.570 181.125 91.830 181.445 ;
        RECT 91.110 180.105 91.370 180.425 ;
        RECT 91.170 178.385 91.310 180.105 ;
        RECT 91.110 178.065 91.370 178.385 ;
        RECT 89.270 175.685 89.530 176.005 ;
        RECT 86.510 174.665 86.770 174.985 ;
        RECT 90.650 173.985 90.910 174.305 ;
        RECT 84.210 171.945 84.470 172.265 ;
        RECT 84.270 170.565 84.410 171.945 ;
        RECT 84.670 171.265 84.930 171.585 ;
        RECT 83.750 170.245 84.010 170.565 ;
        RECT 84.210 170.245 84.470 170.565 ;
        RECT 84.730 169.885 84.870 171.265 ;
        RECT 83.290 169.565 83.550 169.885 ;
        RECT 84.210 169.565 84.470 169.885 ;
        RECT 84.670 169.565 84.930 169.885 ;
        RECT 78.230 169.225 78.490 169.545 ;
        RECT 75.470 168.885 75.730 169.205 ;
        RECT 75.530 167.845 75.670 168.885 ;
        RECT 78.290 167.845 78.430 169.225 ;
        RECT 75.470 167.525 75.730 167.845 ;
        RECT 78.230 167.525 78.490 167.845 ;
        RECT 72.710 166.845 72.970 167.165 ;
        RECT 75.930 166.845 76.190 167.165 ;
        RECT 72.770 161.725 72.910 166.845 ;
        RECT 73.170 166.505 73.430 166.825 ;
        RECT 73.230 165.125 73.370 166.505 ;
        RECT 73.170 164.805 73.430 165.125 ;
        RECT 72.710 161.405 72.970 161.725 ;
        RECT 72.770 157.985 72.910 161.405 ;
        RECT 73.230 161.385 73.370 164.805 ;
        RECT 75.470 163.105 75.730 163.425 ;
        RECT 74.550 161.405 74.810 161.725 ;
        RECT 73.170 161.065 73.430 161.385 ;
        RECT 72.710 157.665 72.970 157.985 ;
        RECT 72.710 155.285 72.970 155.605 ;
        RECT 72.250 150.185 72.510 150.505 ;
        RECT 71.790 148.145 72.050 148.465 ;
        RECT 71.850 147.445 71.990 148.145 ;
        RECT 72.770 147.785 72.910 155.285 ;
        RECT 74.610 153.565 74.750 161.405 ;
        RECT 75.010 160.385 75.270 160.705 ;
        RECT 75.070 155.945 75.210 160.385 ;
        RECT 75.010 155.625 75.270 155.945 ;
        RECT 74.550 153.245 74.810 153.565 ;
        RECT 73.630 149.505 73.890 149.825 ;
        RECT 72.710 147.465 72.970 147.785 ;
        RECT 73.170 147.465 73.430 147.785 ;
        RECT 71.790 147.125 72.050 147.445 ;
        RECT 71.850 143.025 71.990 147.125 ;
        RECT 72.770 147.105 72.910 147.465 ;
        RECT 72.710 146.785 72.970 147.105 ;
        RECT 71.790 142.705 72.050 143.025 ;
        RECT 71.850 139.965 71.990 142.705 ;
        RECT 72.770 141.665 72.910 146.785 ;
        RECT 73.230 146.085 73.370 147.465 ;
        RECT 73.170 145.765 73.430 146.085 ;
        RECT 73.690 145.065 73.830 149.505 ;
        RECT 75.010 147.465 75.270 147.785 ;
        RECT 75.070 146.085 75.210 147.465 ;
        RECT 75.010 145.765 75.270 146.085 ;
        RECT 74.090 145.085 74.350 145.405 ;
        RECT 73.630 144.745 73.890 145.065 ;
        RECT 72.710 141.345 72.970 141.665 ;
        RECT 71.790 139.645 72.050 139.965 ;
        RECT 73.690 139.625 73.830 144.745 ;
        RECT 74.150 142.005 74.290 145.085 ;
        RECT 74.090 141.685 74.350 142.005 ;
        RECT 74.150 140.645 74.290 141.685 ;
        RECT 74.090 140.325 74.350 140.645 ;
        RECT 73.630 139.305 73.890 139.625 ;
        RECT 71.330 138.965 71.590 139.285 ;
        RECT 70.410 138.625 70.670 138.945 ;
        RECT 70.470 135.205 70.610 138.625 ;
        RECT 70.410 134.885 70.670 135.205 ;
        RECT 69.950 133.865 70.210 134.185 ;
        RECT 70.870 133.865 71.130 134.185 ;
        RECT 72.250 133.865 72.510 134.185 ;
        RECT 68.570 132.165 68.830 132.485 ;
        RECT 70.930 131.465 71.070 133.865 ;
        RECT 71.790 131.485 72.050 131.805 ;
        RECT 70.870 131.145 71.130 131.465 ;
        RECT 71.330 131.145 71.590 131.465 ;
        RECT 70.410 130.805 70.670 131.125 ;
        RECT 70.470 125.345 70.610 130.805 ;
        RECT 71.390 129.765 71.530 131.145 ;
        RECT 71.330 129.445 71.590 129.765 ;
        RECT 71.390 126.365 71.530 129.445 ;
        RECT 71.330 126.045 71.590 126.365 ;
        RECT 71.850 125.685 71.990 131.485 ;
        RECT 71.790 125.365 72.050 125.685 ;
        RECT 70.410 125.025 70.670 125.345 ;
        RECT 70.470 124.325 70.610 125.025 ;
        RECT 70.410 124.005 70.670 124.325 ;
        RECT 69.030 123.665 69.290 123.985 ;
        RECT 69.090 121.605 69.230 123.665 ;
        RECT 69.030 121.285 69.290 121.605 ;
        RECT 71.850 119.905 71.990 125.365 ;
        RECT 72.310 120.585 72.450 133.865 ;
        RECT 73.630 133.525 73.890 133.845 ;
        RECT 73.690 131.125 73.830 133.525 ;
        RECT 73.630 130.805 73.890 131.125 ;
        RECT 72.710 129.105 72.970 129.425 ;
        RECT 72.770 127.045 72.910 129.105 ;
        RECT 73.690 128.745 73.830 130.805 ;
        RECT 73.630 128.425 73.890 128.745 ;
        RECT 72.710 126.725 72.970 127.045 ;
        RECT 75.530 126.025 75.670 163.105 ;
        RECT 75.990 162.405 76.130 166.845 ;
        RECT 78.690 165.825 78.950 166.145 ;
        RECT 78.750 164.105 78.890 165.825 ;
        RECT 79.910 165.290 81.790 165.660 ;
        RECT 83.350 164.445 83.490 169.565 ;
        RECT 84.270 165.125 84.410 169.565 ;
        RECT 86.970 168.545 87.230 168.865 ;
        RECT 84.210 164.805 84.470 165.125 ;
        RECT 83.290 164.125 83.550 164.445 ;
        RECT 78.690 163.785 78.950 164.105 ;
        RECT 79.610 163.105 79.870 163.425 ;
        RECT 75.930 162.085 76.190 162.405 ;
        RECT 75.990 161.725 76.130 162.085 ;
        RECT 79.670 162.065 79.810 163.105 ;
        RECT 79.610 161.745 79.870 162.065 ;
        RECT 75.930 161.405 76.190 161.725 ;
        RECT 78.690 161.405 78.950 161.725 ;
        RECT 78.230 160.385 78.490 160.705 ;
        RECT 78.290 158.325 78.430 160.385 ;
        RECT 78.750 159.005 78.890 161.405 ;
        RECT 83.350 161.385 83.490 164.125 ;
        RECT 85.130 161.745 85.390 162.065 ;
        RECT 83.290 161.065 83.550 161.385 ;
        RECT 81.910 160.385 82.170 160.705 ;
        RECT 79.910 159.850 81.790 160.220 ;
        RECT 81.970 159.005 82.110 160.385 ;
        RECT 83.350 159.005 83.490 161.065 ;
        RECT 85.190 159.685 85.330 161.745 ;
        RECT 86.510 161.065 86.770 161.385 ;
        RECT 85.130 159.365 85.390 159.685 ;
        RECT 85.590 159.025 85.850 159.345 ;
        RECT 78.690 158.685 78.950 159.005 ;
        RECT 81.910 158.685 82.170 159.005 ;
        RECT 83.290 158.685 83.550 159.005 ;
        RECT 78.230 158.005 78.490 158.325 ;
        RECT 85.650 157.985 85.790 159.025 ;
        RECT 86.050 158.345 86.310 158.665 ;
        RECT 85.590 157.665 85.850 157.985 ;
        RECT 86.110 156.625 86.250 158.345 ;
        RECT 86.050 156.305 86.310 156.625 ;
        RECT 79.910 154.410 81.790 154.780 ;
        RECT 82.830 152.905 83.090 153.225 ;
        RECT 81.910 152.225 82.170 152.545 ;
        RECT 81.970 151.185 82.110 152.225 ;
        RECT 81.910 150.865 82.170 151.185 ;
        RECT 79.150 149.505 79.410 149.825 ;
        RECT 79.210 148.125 79.350 149.505 ;
        RECT 79.910 148.970 81.790 149.340 ;
        RECT 79.150 147.805 79.410 148.125 ;
        RECT 75.930 147.465 76.190 147.785 ;
        RECT 75.990 142.685 76.130 147.465 ;
        RECT 79.210 146.085 79.350 147.805 ;
        RECT 82.370 147.125 82.630 147.445 ;
        RECT 80.070 146.785 80.330 147.105 ;
        RECT 80.130 146.085 80.270 146.785 ;
        RECT 82.430 146.085 82.570 147.125 ;
        RECT 79.150 145.765 79.410 146.085 ;
        RECT 80.070 145.765 80.330 146.085 ;
        RECT 82.370 145.765 82.630 146.085 ;
        RECT 82.890 144.725 83.030 152.905 ;
        RECT 83.290 152.565 83.550 152.885 ;
        RECT 83.350 145.405 83.490 152.565 ;
        RECT 84.670 152.225 84.930 152.545 ;
        RECT 84.730 150.845 84.870 152.225 ;
        RECT 86.570 150.845 86.710 161.065 ;
        RECT 87.030 158.665 87.170 168.545 ;
        RECT 87.430 166.845 87.690 167.165 ;
        RECT 86.970 158.345 87.230 158.665 ;
        RECT 86.970 157.725 87.230 157.985 ;
        RECT 87.490 157.725 87.630 166.845 ;
        RECT 89.730 163.445 89.990 163.765 ;
        RECT 89.790 160.705 89.930 163.445 ;
        RECT 90.190 161.405 90.450 161.725 ;
        RECT 87.890 160.385 88.150 160.705 ;
        RECT 89.730 160.385 89.990 160.705 ;
        RECT 87.950 158.665 88.090 160.385 ;
        RECT 87.890 158.345 88.150 158.665 ;
        RECT 86.970 157.665 87.630 157.725 ;
        RECT 87.030 157.585 87.630 157.665 ;
        RECT 87.030 155.605 87.170 157.585 ;
        RECT 87.950 156.965 88.090 158.345 ;
        RECT 88.350 158.005 88.610 158.325 ;
        RECT 87.890 156.645 88.150 156.965 ;
        RECT 87.950 156.285 88.090 156.645 ;
        RECT 87.890 155.965 88.150 156.285 ;
        RECT 88.410 155.945 88.550 158.005 ;
        RECT 89.790 156.285 89.930 160.385 ;
        RECT 90.250 159.685 90.390 161.405 ;
        RECT 90.190 159.365 90.450 159.685 ;
        RECT 89.730 155.965 89.990 156.285 ;
        RECT 88.350 155.625 88.610 155.945 ;
        RECT 86.970 155.285 87.230 155.605 ;
        RECT 87.030 153.225 87.170 155.285 ;
        RECT 87.890 154.945 88.150 155.265 ;
        RECT 86.970 152.905 87.230 153.225 ;
        RECT 84.670 150.525 84.930 150.845 ;
        RECT 86.510 150.525 86.770 150.845 ;
        RECT 86.970 149.505 87.230 149.825 ;
        RECT 87.030 148.465 87.170 149.505 ;
        RECT 86.970 148.375 87.230 148.465 ;
        RECT 86.570 148.235 87.230 148.375 ;
        RECT 84.210 147.805 84.470 148.125 ;
        RECT 83.290 145.085 83.550 145.405 ;
        RECT 82.830 144.405 83.090 144.725 ;
        RECT 79.910 143.530 81.790 143.900 ;
        RECT 75.930 142.365 76.190 142.685 ;
        RECT 78.690 142.365 78.950 142.685 ;
        RECT 80.990 142.365 81.250 142.685 ;
        RECT 78.220 139.110 78.500 139.480 ;
        RECT 78.290 137.925 78.430 139.110 ;
        RECT 78.230 137.605 78.490 137.925 ;
        RECT 78.750 137.245 78.890 142.365 ;
        RECT 81.050 142.085 81.190 142.365 ;
        RECT 79.150 141.685 79.410 142.005 ;
        RECT 79.670 141.945 81.190 142.085 ;
        RECT 79.210 140.645 79.350 141.685 ;
        RECT 79.150 140.325 79.410 140.645 ;
        RECT 79.670 139.285 79.810 141.945 ;
        RECT 83.350 139.965 83.490 145.085 ;
        RECT 83.750 144.975 84.010 145.065 ;
        RECT 84.270 144.975 84.410 147.805 ;
        RECT 86.570 145.405 86.710 148.235 ;
        RECT 86.970 148.145 87.230 148.235 ;
        RECT 86.970 146.785 87.230 147.105 ;
        RECT 87.030 146.085 87.170 146.785 ;
        RECT 86.970 145.765 87.230 146.085 ;
        RECT 86.510 145.085 86.770 145.405 ;
        RECT 83.750 144.835 84.410 144.975 ;
        RECT 83.750 144.745 84.010 144.835 ;
        RECT 83.290 139.645 83.550 139.965 ;
        RECT 79.610 138.965 79.870 139.285 ;
        RECT 79.910 138.090 81.790 138.460 ;
        RECT 78.690 136.925 78.950 137.245 ;
        RECT 83.350 137.155 83.490 139.645 ;
        RECT 84.270 139.625 84.410 144.835 ;
        RECT 84.210 139.305 84.470 139.625 ;
        RECT 84.670 139.305 84.930 139.625 ;
        RECT 87.430 139.305 87.690 139.625 ;
        RECT 84.730 137.925 84.870 139.305 ;
        RECT 84.670 137.605 84.930 137.925 ;
        RECT 83.350 137.015 83.950 137.155 ;
        RECT 78.230 130.465 78.490 130.785 ;
        RECT 78.290 129.085 78.430 130.465 ;
        RECT 78.230 128.765 78.490 129.085 ;
        RECT 78.750 128.745 78.890 136.925 ;
        RECT 83.290 136.245 83.550 136.565 ;
        RECT 83.350 135.205 83.490 136.245 ;
        RECT 83.290 134.885 83.550 135.205 ;
        RECT 83.810 134.525 83.950 137.015 ;
        RECT 87.490 134.865 87.630 139.305 ;
        RECT 87.950 134.865 88.090 154.945 ;
        RECT 88.810 152.225 89.070 152.545 ;
        RECT 88.870 150.845 89.010 152.225 ;
        RECT 88.810 150.525 89.070 150.845 ;
        RECT 89.730 139.985 89.990 140.305 ;
        RECT 89.270 138.625 89.530 138.945 ;
        RECT 89.330 136.905 89.470 138.625 ;
        RECT 89.790 137.925 89.930 139.985 ;
        RECT 89.730 137.605 89.990 137.925 ;
        RECT 89.270 136.585 89.530 136.905 ;
        RECT 90.190 134.885 90.450 135.205 ;
        RECT 87.430 134.545 87.690 134.865 ;
        RECT 87.890 134.545 88.150 134.865 ;
        RECT 83.750 134.205 84.010 134.525 ;
        RECT 86.050 133.525 86.310 133.845 ;
        RECT 79.910 132.650 81.790 133.020 ;
        RECT 82.370 130.805 82.630 131.125 ;
        RECT 82.430 129.765 82.570 130.805 ;
        RECT 86.110 130.785 86.250 133.525 ;
        RECT 88.810 133.185 89.070 133.505 ;
        RECT 87.890 131.825 88.150 132.145 ;
        RECT 86.050 130.465 86.310 130.785 ;
        RECT 82.370 129.445 82.630 129.765 ;
        RECT 84.210 129.105 84.470 129.425 ;
        RECT 78.690 128.425 78.950 128.745 ;
        RECT 76.850 128.085 77.110 128.405 ;
        RECT 76.910 126.365 77.050 128.085 ;
        RECT 78.750 126.365 78.890 128.425 ;
        RECT 81.910 127.745 82.170 128.065 ;
        RECT 79.910 127.210 81.790 127.580 ;
        RECT 81.970 126.365 82.110 127.745 ;
        RECT 84.270 127.045 84.410 129.105 ;
        RECT 84.210 126.725 84.470 127.045 ;
        RECT 76.850 126.045 77.110 126.365 ;
        RECT 78.690 126.045 78.950 126.365 ;
        RECT 81.910 126.045 82.170 126.365 ;
        RECT 75.470 125.705 75.730 126.025 ;
        RECT 72.250 120.265 72.510 120.585 ;
        RECT 71.790 119.585 72.050 119.905 ;
        RECT 71.850 118.885 71.990 119.585 ;
        RECT 71.790 118.565 72.050 118.885 ;
        RECT 69.490 118.225 69.750 118.545 ;
        RECT 69.550 116.165 69.690 118.225 ;
        RECT 72.310 117.185 72.450 120.265 ;
        RECT 75.530 120.245 75.670 125.705 ;
        RECT 76.390 125.025 76.650 125.345 ;
        RECT 76.450 123.645 76.590 125.025 ;
        RECT 76.390 123.325 76.650 123.645 ;
        RECT 76.910 120.925 77.050 126.045 ;
        RECT 78.750 124.325 78.890 126.045 ;
        RECT 86.110 126.025 86.250 130.465 ;
        RECT 87.950 129.085 88.090 131.825 ;
        RECT 88.870 129.765 89.010 133.185 ;
        RECT 88.810 129.445 89.070 129.765 ;
        RECT 87.890 128.765 88.150 129.085 ;
        RECT 86.510 128.085 86.770 128.405 ;
        RECT 86.050 125.705 86.310 126.025 ;
        RECT 78.690 124.005 78.950 124.325 ;
        RECT 78.750 120.925 78.890 124.005 ;
        RECT 86.050 123.665 86.310 123.985 ;
        RECT 83.290 123.325 83.550 123.645 ;
        RECT 79.910 121.770 81.790 122.140 ;
        RECT 76.850 120.605 77.110 120.925 ;
        RECT 78.690 120.605 78.950 120.925 ;
        RECT 75.470 119.925 75.730 120.245 ;
        RECT 74.090 119.585 74.350 119.905 ;
        RECT 73.170 117.545 73.430 117.865 ;
        RECT 73.630 117.545 73.890 117.865 ;
        RECT 72.250 116.865 72.510 117.185 ;
        RECT 73.230 116.165 73.370 117.545 ;
        RECT 69.490 115.845 69.750 116.165 ;
        RECT 73.170 115.845 73.430 116.165 ;
        RECT 68.560 113.270 68.840 113.640 ;
        RECT 68.630 112.765 68.770 113.270 ;
        RECT 68.570 112.445 68.830 112.765 ;
        RECT 68.110 112.105 68.370 112.425 ;
        RECT 72.710 112.105 72.970 112.425 ;
        RECT 72.250 111.765 72.510 112.085 ;
        RECT 71.790 111.425 72.050 111.745 ;
        RECT 71.330 109.725 71.590 110.045 ;
        RECT 60.290 109.385 60.550 109.705 ;
        RECT 63.970 109.385 64.230 109.705 ;
        RECT 67.190 109.385 67.450 109.705 ;
        RECT 62.130 108.705 62.390 109.025 ;
        RECT 59.370 107.685 59.630 108.005 ;
        RECT 62.190 104.605 62.330 108.705 ;
        RECT 64.910 108.170 66.790 108.540 ;
        RECT 64.430 107.345 64.690 107.665 ;
        RECT 63.510 106.665 63.770 106.985 ;
        RECT 63.570 104.605 63.710 106.665 ;
        RECT 60.290 104.285 60.550 104.605 ;
        RECT 62.130 104.285 62.390 104.605 ;
        RECT 63.510 104.285 63.770 104.605 ;
        RECT 58.910 103.605 59.170 103.925 ;
        RECT 60.350 92.050 60.490 104.285 ;
        RECT 22.170 91.625 23.230 91.765 ;
        RECT 27.160 90.050 27.440 92.050 ;
        RECT 32.680 90.050 32.960 92.050 ;
        RECT 38.200 90.050 38.480 92.050 ;
        RECT 43.720 90.050 44.000 92.050 ;
        RECT 49.240 90.050 49.520 92.050 ;
        RECT 54.760 90.050 55.040 92.050 ;
        RECT 60.280 90.050 60.560 92.050 ;
        RECT 64.490 91.765 64.630 107.345 ;
        RECT 64.910 102.730 66.790 103.100 ;
        RECT 67.250 102.565 67.390 109.385 ;
        RECT 69.950 107.345 70.210 107.665 ;
        RECT 70.010 105.285 70.150 107.345 ;
        RECT 69.950 104.965 70.210 105.285 ;
        RECT 67.190 102.245 67.450 102.565 ;
        RECT 65.410 92.305 66.010 92.445 ;
        RECT 65.410 91.765 65.550 92.305 ;
        RECT 65.870 92.050 66.010 92.305 ;
        RECT 71.390 92.050 71.530 109.725 ;
        RECT 71.850 106.305 71.990 111.425 ;
        RECT 72.310 107.665 72.450 111.765 ;
        RECT 72.770 107.665 72.910 112.105 ;
        RECT 73.690 109.025 73.830 117.545 ;
        RECT 74.150 115.145 74.290 119.585 ;
        RECT 75.530 118.205 75.670 119.925 ;
        RECT 75.470 117.885 75.730 118.205 ;
        RECT 75.530 115.485 75.670 117.885 ;
        RECT 78.750 117.865 78.890 120.605 ;
        RECT 83.350 120.585 83.490 123.325 ;
        RECT 86.110 123.160 86.250 123.665 ;
        RECT 86.570 123.645 86.710 128.085 ;
        RECT 88.350 125.025 88.610 125.345 ;
        RECT 86.510 123.325 86.770 123.645 ;
        RECT 88.410 123.305 88.550 125.025 ;
        RECT 86.040 122.790 86.320 123.160 ;
        RECT 88.350 122.985 88.610 123.305 ;
        RECT 88.410 121.605 88.550 122.985 ;
        RECT 89.730 122.305 89.990 122.625 ;
        RECT 88.350 121.285 88.610 121.605 ;
        RECT 87.430 120.605 87.690 120.925 ;
        RECT 83.290 120.265 83.550 120.585 ;
        RECT 86.970 120.265 87.230 120.585 ;
        RECT 82.370 119.925 82.630 120.245 ;
        RECT 78.690 117.545 78.950 117.865 ;
        RECT 79.910 116.330 81.790 116.700 ;
        RECT 82.430 116.165 82.570 119.925 ;
        RECT 87.030 118.205 87.170 120.265 ;
        RECT 87.490 118.885 87.630 120.605 ;
        RECT 87.890 119.585 88.150 119.905 ;
        RECT 87.430 118.565 87.690 118.885 ;
        RECT 87.950 118.205 88.090 119.585 ;
        RECT 89.790 118.205 89.930 122.305 ;
        RECT 86.970 117.885 87.230 118.205 ;
        RECT 87.890 117.885 88.150 118.205 ;
        RECT 89.730 117.885 89.990 118.205 ;
        RECT 82.370 115.845 82.630 116.165 ;
        RECT 75.470 115.165 75.730 115.485 ;
        RECT 74.090 114.825 74.350 115.145 ;
        RECT 86.050 111.425 86.310 111.745 ;
        RECT 79.910 110.890 81.790 111.260 ;
        RECT 86.110 110.045 86.250 111.425 ;
        RECT 87.030 110.725 87.170 117.885 ;
        RECT 90.250 112.765 90.390 134.885 ;
        RECT 90.710 134.185 90.850 173.985 ;
        RECT 91.170 169.885 91.310 178.065 ;
        RECT 92.550 178.045 92.690 182.145 ;
        RECT 93.470 180.765 93.610 183.845 ;
        RECT 94.330 183.505 94.590 183.825 ;
        RECT 93.410 180.445 93.670 180.765 ;
        RECT 92.490 177.725 92.750 178.045 ;
        RECT 92.950 174.895 93.210 174.985 ;
        RECT 93.470 174.895 93.610 180.445 ;
        RECT 94.390 178.725 94.530 183.505 ;
        RECT 96.170 182.145 96.430 182.465 ;
        RECT 96.230 180.765 96.370 182.145 ;
        RECT 96.170 180.445 96.430 180.765 ;
        RECT 97.090 179.425 97.350 179.745 ;
        RECT 94.910 178.890 96.790 179.260 ;
        RECT 94.330 178.405 94.590 178.725 ;
        RECT 97.150 178.045 97.290 179.425 ;
        RECT 97.610 178.385 97.750 190.985 ;
        RECT 97.550 178.065 97.810 178.385 ;
        RECT 93.870 177.725 94.130 178.045 ;
        RECT 96.630 177.955 96.890 178.045 ;
        RECT 96.230 177.815 96.890 177.955 ;
        RECT 93.930 175.325 94.070 177.725 ;
        RECT 93.870 175.005 94.130 175.325 ;
        RECT 92.950 174.755 93.610 174.895 ;
        RECT 92.950 174.665 93.210 174.755 ;
        RECT 93.930 174.305 94.070 175.005 ;
        RECT 96.230 174.985 96.370 177.815 ;
        RECT 96.630 177.725 96.890 177.815 ;
        RECT 97.090 177.725 97.350 178.045 ;
        RECT 98.010 177.725 98.270 178.045 ;
        RECT 97.550 176.705 97.810 177.025 ;
        RECT 96.170 174.665 96.430 174.985 ;
        RECT 93.870 173.985 94.130 174.305 ;
        RECT 94.910 173.450 96.790 173.820 ;
        RECT 97.090 171.945 97.350 172.265 ;
        RECT 91.110 169.565 91.370 169.885 ;
        RECT 93.410 168.885 93.670 169.205 ;
        RECT 93.470 167.505 93.610 168.885 ;
        RECT 94.910 168.010 96.790 168.380 ;
        RECT 97.150 167.925 97.290 171.945 ;
        RECT 97.610 168.605 97.750 176.705 ;
        RECT 98.070 175.665 98.210 177.725 ;
        RECT 98.530 176.005 98.670 191.325 ;
        RECT 102.210 190.965 102.350 193.025 ;
        RECT 102.670 192.325 102.810 194.045 ;
        RECT 102.610 192.005 102.870 192.325 ;
        RECT 102.150 190.645 102.410 190.965 ;
        RECT 99.390 190.305 99.650 190.625 ;
        RECT 99.450 188.495 99.590 190.305 ;
        RECT 102.670 188.925 102.810 192.005 ;
        RECT 103.590 189.605 103.730 194.045 ;
        RECT 105.830 193.025 106.090 193.345 ;
        RECT 105.890 191.645 106.030 193.025 ;
        RECT 109.910 192.490 111.790 192.860 ;
        RECT 105.830 191.325 106.090 191.645 ;
        RECT 107.670 190.985 107.930 191.305 ;
        RECT 106.290 190.645 106.550 190.965 ;
        RECT 103.530 189.285 103.790 189.605 ;
        RECT 100.770 188.605 101.030 188.925 ;
        RECT 102.610 188.605 102.870 188.925 ;
        RECT 104.910 188.605 105.170 188.925 ;
        RECT 99.850 188.495 100.110 188.585 ;
        RECT 99.450 188.355 100.110 188.495 ;
        RECT 99.850 188.265 100.110 188.355 ;
        RECT 99.910 185.525 100.050 188.265 ;
        RECT 100.310 187.585 100.570 187.905 ;
        RECT 99.850 185.205 100.110 185.525 ;
        RECT 100.370 184.165 100.510 187.585 ;
        RECT 100.310 183.845 100.570 184.165 ;
        RECT 100.830 182.465 100.970 188.605 ;
        RECT 104.450 187.925 104.710 188.245 ;
        RECT 104.510 186.205 104.650 187.925 ;
        RECT 104.450 185.885 104.710 186.205 ;
        RECT 101.230 185.545 101.490 185.865 ;
        RECT 101.290 184.165 101.430 185.545 ;
        RECT 102.610 184.865 102.870 185.185 ;
        RECT 101.230 183.845 101.490 184.165 ;
        RECT 100.770 182.145 101.030 182.465 ;
        RECT 100.830 178.725 100.970 182.145 ;
        RECT 102.670 180.765 102.810 184.865 ;
        RECT 103.530 182.825 103.790 183.145 ;
        RECT 102.610 180.445 102.870 180.765 ;
        RECT 103.590 180.085 103.730 182.825 ;
        RECT 104.510 182.805 104.650 185.885 ;
        RECT 104.970 183.485 105.110 188.605 ;
        RECT 106.350 186.885 106.490 190.645 ;
        RECT 106.290 186.565 106.550 186.885 ;
        RECT 105.830 184.865 106.090 185.185 ;
        RECT 104.910 183.165 105.170 183.485 ;
        RECT 104.450 182.485 104.710 182.805 ;
        RECT 103.530 179.765 103.790 180.085 ;
        RECT 100.310 178.405 100.570 178.725 ;
        RECT 100.770 178.405 101.030 178.725 ;
        RECT 100.370 178.045 100.510 178.405 ;
        RECT 99.850 177.725 100.110 178.045 ;
        RECT 100.310 177.725 100.570 178.045 ;
        RECT 98.930 176.705 99.190 177.025 ;
        RECT 98.470 175.685 98.730 176.005 ;
        RECT 98.010 175.345 98.270 175.665 ;
        RECT 98.000 172.430 98.280 172.800 ;
        RECT 98.070 169.545 98.210 172.430 ;
        RECT 98.470 171.945 98.730 172.265 ;
        RECT 98.010 169.225 98.270 169.545 ;
        RECT 97.610 168.465 98.210 168.605 ;
        RECT 97.150 167.785 97.750 167.925 ;
        RECT 93.410 167.185 93.670 167.505 ;
        RECT 93.870 166.165 94.130 166.485 ;
        RECT 92.950 165.825 93.210 166.145 ;
        RECT 93.010 164.105 93.150 165.825 ;
        RECT 92.950 163.785 93.210 164.105 ;
        RECT 93.410 163.785 93.670 164.105 ;
        RECT 91.110 163.105 91.370 163.425 ;
        RECT 91.170 158.665 91.310 163.105 ;
        RECT 93.470 159.685 93.610 163.785 ;
        RECT 93.930 162.065 94.070 166.165 ;
        RECT 94.330 163.105 94.590 163.425 ;
        RECT 97.090 163.105 97.350 163.425 ;
        RECT 93.870 161.745 94.130 162.065 ;
        RECT 93.410 159.365 93.670 159.685 ;
        RECT 94.390 158.665 94.530 163.105 ;
        RECT 94.910 162.570 96.790 162.940 ;
        RECT 97.150 162.405 97.290 163.105 ;
        RECT 95.250 162.085 95.510 162.405 ;
        RECT 97.090 162.085 97.350 162.405 ;
        RECT 95.310 159.005 95.450 162.085 ;
        RECT 96.170 161.065 96.430 161.385 ;
        RECT 96.230 159.345 96.370 161.065 ;
        RECT 97.610 159.345 97.750 167.785 ;
        RECT 96.170 159.025 96.430 159.345 ;
        RECT 97.550 159.025 97.810 159.345 ;
        RECT 95.250 158.685 95.510 159.005 ;
        RECT 91.110 158.345 91.370 158.665 ;
        RECT 94.330 158.345 94.590 158.665 ;
        RECT 97.090 158.345 97.350 158.665 ;
        RECT 93.870 158.005 94.130 158.325 ;
        RECT 93.930 156.625 94.070 158.005 ;
        RECT 94.910 157.130 96.790 157.500 ;
        RECT 93.870 156.305 94.130 156.625 ;
        RECT 97.150 156.285 97.290 158.345 ;
        RECT 97.550 157.665 97.810 157.985 ;
        RECT 95.250 155.965 95.510 156.285 ;
        RECT 97.090 156.195 97.350 156.285 ;
        RECT 96.690 156.055 97.350 156.195 ;
        RECT 93.870 154.945 94.130 155.265 ;
        RECT 92.950 150.865 93.210 151.185 ;
        RECT 93.010 148.805 93.150 150.865 ;
        RECT 92.950 148.485 93.210 148.805 ;
        RECT 92.950 147.805 93.210 148.125 ;
        RECT 92.490 140.325 92.750 140.645 ;
        RECT 92.550 139.965 92.690 140.325 ;
        RECT 91.110 139.645 91.370 139.965 ;
        RECT 92.490 139.645 92.750 139.965 ;
        RECT 91.170 139.480 91.310 139.645 ;
        RECT 91.100 139.110 91.380 139.480 ;
        RECT 91.570 136.245 91.830 136.565 ;
        RECT 91.630 135.205 91.770 136.245 ;
        RECT 91.570 134.885 91.830 135.205 ;
        RECT 92.550 134.865 92.690 139.645 ;
        RECT 93.010 139.625 93.150 147.805 ;
        RECT 93.930 144.805 94.070 154.945 ;
        RECT 95.310 154.245 95.450 155.965 ;
        RECT 95.250 153.925 95.510 154.245 ;
        RECT 95.310 153.225 95.450 153.925 ;
        RECT 95.250 152.905 95.510 153.225 ;
        RECT 96.690 152.885 96.830 156.055 ;
        RECT 97.090 155.965 97.350 156.055 ;
        RECT 97.090 154.945 97.350 155.265 ;
        RECT 96.630 152.565 96.890 152.885 ;
        RECT 94.330 152.225 94.590 152.545 ;
        RECT 94.390 147.785 94.530 152.225 ;
        RECT 94.910 151.690 96.790 152.060 ;
        RECT 97.150 150.845 97.290 154.945 ;
        RECT 97.090 150.525 97.350 150.845 ;
        RECT 96.630 149.845 96.890 150.165 ;
        RECT 96.690 148.125 96.830 149.845 ;
        RECT 97.090 148.485 97.350 148.805 ;
        RECT 96.630 147.805 96.890 148.125 ;
        RECT 94.330 147.465 94.590 147.785 ;
        RECT 94.910 146.250 96.790 146.620 ;
        RECT 93.930 144.665 94.530 144.805 ;
        RECT 92.950 139.305 93.210 139.625 ;
        RECT 92.490 134.545 92.750 134.865 ;
        RECT 94.390 134.525 94.530 144.665 ;
        RECT 94.910 140.810 96.790 141.180 ;
        RECT 94.910 135.370 96.790 135.740 ;
        RECT 94.790 134.885 95.050 135.205 ;
        RECT 94.330 134.205 94.590 134.525 ;
        RECT 90.650 133.865 90.910 134.185 ;
        RECT 94.850 133.925 94.990 134.885 ;
        RECT 94.390 133.785 94.990 133.925 ;
        RECT 93.410 133.185 93.670 133.505 ;
        RECT 93.470 129.765 93.610 133.185 ;
        RECT 93.410 129.445 93.670 129.765 ;
        RECT 92.030 125.705 92.290 126.025 ;
        RECT 91.570 125.365 91.830 125.685 ;
        RECT 91.630 124.325 91.770 125.365 ;
        RECT 91.570 124.005 91.830 124.325 ;
        RECT 92.090 123.645 92.230 125.705 ;
        RECT 93.870 125.025 94.130 125.345 ;
        RECT 92.030 123.325 92.290 123.645 ;
        RECT 93.930 120.245 94.070 125.025 ;
        RECT 93.870 119.925 94.130 120.245 ;
        RECT 94.390 112.765 94.530 133.785 ;
        RECT 94.910 129.930 96.790 130.300 ;
        RECT 97.150 129.765 97.290 148.485 ;
        RECT 97.610 145.405 97.750 157.665 ;
        RECT 98.070 150.245 98.210 168.465 ;
        RECT 98.530 164.445 98.670 171.945 ;
        RECT 98.470 164.125 98.730 164.445 ;
        RECT 98.470 163.105 98.730 163.425 ;
        RECT 98.530 160.705 98.670 163.105 ;
        RECT 98.470 160.385 98.730 160.705 ;
        RECT 98.470 159.025 98.730 159.345 ;
        RECT 98.530 153.225 98.670 159.025 ;
        RECT 98.470 152.905 98.730 153.225 ;
        RECT 98.070 150.105 98.670 150.245 ;
        RECT 98.990 150.165 99.130 176.705 ;
        RECT 99.910 174.985 100.050 177.725 ;
        RECT 100.370 177.025 100.510 177.725 ;
        RECT 100.310 176.705 100.570 177.025 ;
        RECT 100.830 175.325 100.970 178.405 ;
        RECT 104.510 177.705 104.650 182.485 ;
        RECT 104.970 180.085 105.110 183.165 ;
        RECT 104.910 179.765 105.170 180.085 ;
        RECT 105.890 178.725 106.030 184.865 ;
        RECT 107.210 183.165 107.470 183.485 ;
        RECT 107.270 181.445 107.410 183.165 ;
        RECT 107.730 183.145 107.870 190.985 ;
        RECT 112.270 190.305 112.530 190.625 ;
        RECT 112.330 189.265 112.470 190.305 ;
        RECT 112.270 188.945 112.530 189.265 ;
        RECT 114.110 188.265 114.370 188.585 ;
        RECT 109.510 187.585 109.770 187.905 ;
        RECT 109.570 186.205 109.710 187.585 ;
        RECT 109.910 187.050 111.790 187.420 ;
        RECT 109.510 185.885 109.770 186.205 ;
        RECT 107.670 182.825 107.930 183.145 ;
        RECT 107.210 181.125 107.470 181.445 ;
        RECT 107.730 180.425 107.870 182.825 ;
        RECT 107.670 180.105 107.930 180.425 ;
        RECT 105.830 178.405 106.090 178.725 ;
        RECT 104.450 177.385 104.710 177.705 ;
        RECT 106.750 176.705 107.010 177.025 ;
        RECT 105.370 175.345 105.630 175.665 ;
        RECT 100.770 175.005 101.030 175.325 ;
        RECT 99.850 174.840 100.110 174.985 ;
        RECT 103.990 174.895 104.250 174.985 ;
        RECT 99.840 174.470 100.120 174.840 ;
        RECT 103.990 174.755 104.650 174.895 ;
        RECT 103.990 174.665 104.250 174.755 ;
        RECT 100.770 174.325 101.030 174.645 ;
        RECT 100.830 169.545 100.970 174.325 ;
        RECT 103.070 172.285 103.330 172.605 ;
        RECT 103.130 172.005 103.270 172.285 ;
        RECT 103.130 171.865 103.730 172.005 ;
        RECT 103.590 169.885 103.730 171.865 ;
        RECT 104.510 171.585 104.650 174.755 ;
        RECT 104.910 173.985 105.170 174.305 ;
        RECT 104.450 171.265 104.710 171.585 ;
        RECT 103.530 169.565 103.790 169.885 ;
        RECT 100.770 169.225 101.030 169.545 ;
        RECT 100.310 168.885 100.570 169.205 ;
        RECT 99.850 168.545 100.110 168.865 ;
        RECT 99.910 167.845 100.050 168.545 ;
        RECT 99.850 167.525 100.110 167.845 ;
        RECT 99.390 166.505 99.650 166.825 ;
        RECT 99.850 166.505 100.110 166.825 ;
        RECT 99.450 163.335 99.590 166.505 ;
        RECT 99.910 165.125 100.050 166.505 ;
        RECT 99.850 164.805 100.110 165.125 ;
        RECT 99.850 163.335 100.110 163.425 ;
        RECT 99.450 163.195 100.110 163.335 ;
        RECT 99.850 163.105 100.110 163.195 ;
        RECT 99.390 158.345 99.650 158.665 ;
        RECT 99.450 156.285 99.590 158.345 ;
        RECT 99.910 156.625 100.050 163.105 ;
        RECT 100.370 161.725 100.510 168.885 ;
        RECT 101.230 168.545 101.490 168.865 ;
        RECT 101.290 166.825 101.430 168.545 ;
        RECT 102.150 167.185 102.410 167.505 ;
        RECT 101.230 166.735 101.490 166.825 ;
        RECT 100.830 166.595 101.490 166.735 ;
        RECT 100.310 161.405 100.570 161.725 ;
        RECT 100.370 158.665 100.510 161.405 ;
        RECT 100.830 161.385 100.970 166.595 ;
        RECT 101.230 166.505 101.490 166.595 ;
        RECT 102.210 165.125 102.350 167.185 ;
        RECT 103.590 167.165 103.730 169.565 ;
        RECT 103.530 166.845 103.790 167.165 ;
        RECT 102.150 164.805 102.410 165.125 ;
        RECT 103.590 164.105 103.730 166.845 ;
        RECT 103.990 165.825 104.250 166.145 ;
        RECT 103.530 163.785 103.790 164.105 ;
        RECT 104.050 163.765 104.190 165.825 ;
        RECT 103.990 163.445 104.250 163.765 ;
        RECT 101.690 163.105 101.950 163.425 ;
        RECT 103.530 163.105 103.790 163.425 ;
        RECT 100.770 161.065 101.030 161.385 ;
        RECT 100.310 158.345 100.570 158.665 ;
        RECT 100.310 157.665 100.570 157.985 ;
        RECT 100.370 156.965 100.510 157.665 ;
        RECT 100.310 156.645 100.570 156.965 ;
        RECT 99.850 156.305 100.110 156.625 ;
        RECT 99.390 155.965 99.650 156.285 ;
        RECT 99.450 154.245 99.590 155.965 ;
        RECT 100.370 155.125 100.510 156.645 ;
        RECT 99.910 154.985 100.510 155.125 ;
        RECT 99.390 153.925 99.650 154.245 ;
        RECT 99.910 153.565 100.050 154.985 ;
        RECT 99.850 153.245 100.110 153.565 ;
        RECT 100.310 152.905 100.570 153.225 ;
        RECT 99.850 152.225 100.110 152.545 ;
        RECT 99.910 151.525 100.050 152.225 ;
        RECT 100.370 151.525 100.510 152.905 ;
        RECT 100.830 152.545 100.970 161.065 ;
        RECT 101.750 161.045 101.890 163.105 ;
        RECT 103.590 161.725 103.730 163.105 ;
        RECT 102.150 161.405 102.410 161.725 ;
        RECT 103.530 161.405 103.790 161.725 ;
        RECT 101.690 160.725 101.950 161.045 ;
        RECT 101.750 159.345 101.890 160.725 ;
        RECT 102.210 159.685 102.350 161.405 ;
        RECT 103.070 161.065 103.330 161.385 ;
        RECT 102.150 159.365 102.410 159.685 ;
        RECT 101.690 159.025 101.950 159.345 ;
        RECT 101.690 157.665 101.950 157.985 ;
        RECT 100.770 152.455 101.030 152.545 ;
        RECT 100.770 152.315 101.430 152.455 ;
        RECT 100.770 152.225 101.030 152.315 ;
        RECT 99.850 151.205 100.110 151.525 ;
        RECT 100.310 151.205 100.570 151.525 ;
        RECT 99.850 150.755 100.110 150.845 ;
        RECT 99.850 150.615 100.510 150.755 ;
        RECT 99.850 150.525 100.110 150.615 ;
        RECT 98.010 149.505 98.270 149.825 ;
        RECT 98.070 148.805 98.210 149.505 ;
        RECT 98.010 148.485 98.270 148.805 ;
        RECT 98.010 147.640 98.270 147.785 ;
        RECT 98.000 147.270 98.280 147.640 ;
        RECT 97.550 145.085 97.810 145.405 ;
        RECT 98.530 144.805 98.670 150.105 ;
        RECT 98.930 149.845 99.190 150.165 ;
        RECT 99.390 149.565 99.650 149.825 ;
        RECT 98.990 149.505 99.650 149.565 ;
        RECT 98.990 149.425 99.590 149.505 ;
        RECT 98.990 147.695 99.130 149.425 ;
        RECT 98.990 147.555 99.590 147.695 ;
        RECT 97.610 144.665 98.670 144.805 ;
        RECT 98.930 144.745 99.190 145.065 ;
        RECT 97.610 133.845 97.750 144.665 ;
        RECT 98.470 144.065 98.730 144.385 ;
        RECT 98.010 139.645 98.270 139.965 ;
        RECT 98.070 137.925 98.210 139.645 ;
        RECT 98.010 137.605 98.270 137.925 ;
        RECT 98.070 134.525 98.210 137.605 ;
        RECT 98.010 134.205 98.270 134.525 ;
        RECT 97.550 133.525 97.810 133.845 ;
        RECT 97.550 131.145 97.810 131.465 ;
        RECT 97.090 129.445 97.350 129.765 ;
        RECT 95.250 128.425 95.510 128.745 ;
        RECT 94.790 127.745 95.050 128.065 ;
        RECT 94.850 126.365 94.990 127.745 ;
        RECT 94.790 126.045 95.050 126.365 ;
        RECT 95.310 125.685 95.450 128.425 ;
        RECT 97.610 126.275 97.750 131.145 ;
        RECT 98.530 129.765 98.670 144.065 ;
        RECT 98.990 139.965 99.130 144.745 ;
        RECT 98.930 139.645 99.190 139.965 ;
        RECT 98.990 134.525 99.130 139.645 ;
        RECT 98.930 134.205 99.190 134.525 ;
        RECT 98.930 133.185 99.190 133.505 ;
        RECT 98.990 132.485 99.130 133.185 ;
        RECT 99.450 132.485 99.590 147.555 ;
        RECT 99.850 147.465 100.110 147.785 ;
        RECT 100.370 147.640 100.510 150.615 ;
        RECT 101.290 150.165 101.430 152.315 ;
        RECT 100.770 149.845 101.030 150.165 ;
        RECT 101.230 149.845 101.490 150.165 ;
        RECT 99.910 145.065 100.050 147.465 ;
        RECT 100.300 147.270 100.580 147.640 ;
        RECT 100.830 147.445 100.970 149.845 ;
        RECT 100.370 145.405 100.510 147.270 ;
        RECT 100.770 147.125 101.030 147.445 ;
        RECT 100.830 145.405 100.970 147.125 ;
        RECT 100.310 145.085 100.570 145.405 ;
        RECT 100.770 145.085 101.030 145.405 ;
        RECT 99.850 144.745 100.110 145.065 ;
        RECT 100.370 139.875 100.510 145.085 ;
        RECT 100.830 140.840 100.970 145.085 ;
        RECT 101.750 141.575 101.890 157.665 ;
        RECT 103.130 155.605 103.270 161.065 ;
        RECT 103.590 159.005 103.730 161.405 ;
        RECT 103.530 158.685 103.790 159.005 ;
        RECT 104.510 156.625 104.650 171.265 ;
        RECT 104.450 156.305 104.710 156.625 ;
        RECT 103.070 155.285 103.330 155.605 ;
        RECT 102.610 152.225 102.870 152.545 ;
        RECT 102.150 150.525 102.410 150.845 ;
        RECT 102.210 145.405 102.350 150.525 ;
        RECT 102.670 147.445 102.810 152.225 ;
        RECT 103.130 150.845 103.270 155.285 ;
        RECT 104.450 153.245 104.710 153.565 ;
        RECT 103.070 150.525 103.330 150.845 ;
        RECT 102.610 147.125 102.870 147.445 ;
        RECT 103.130 145.405 103.270 150.525 ;
        RECT 104.510 148.035 104.650 153.245 ;
        RECT 104.970 149.825 105.110 173.985 ;
        RECT 105.430 173.285 105.570 175.345 ;
        RECT 106.810 174.985 106.950 176.705 ;
        RECT 107.210 175.685 107.470 176.005 ;
        RECT 105.830 174.840 106.090 174.985 ;
        RECT 105.820 174.470 106.100 174.840 ;
        RECT 106.750 174.665 107.010 174.985 ;
        RECT 107.270 174.970 107.410 175.685 ;
        RECT 107.210 174.650 107.470 174.970 ;
        RECT 105.370 172.965 105.630 173.285 ;
        RECT 105.430 158.665 105.570 172.965 ;
        RECT 105.830 169.225 106.090 169.545 ;
        RECT 105.370 158.345 105.630 158.665 ;
        RECT 105.370 152.225 105.630 152.545 ;
        RECT 104.910 149.505 105.170 149.825 ;
        RECT 105.430 148.465 105.570 152.225 ;
        RECT 105.370 148.145 105.630 148.465 ;
        RECT 104.910 148.035 105.170 148.125 ;
        RECT 104.510 147.895 105.170 148.035 ;
        RECT 104.910 147.805 105.170 147.895 ;
        RECT 102.150 145.085 102.410 145.405 ;
        RECT 103.070 145.085 103.330 145.405 ;
        RECT 102.610 144.405 102.870 144.725 ;
        RECT 101.290 141.435 101.890 141.575 ;
        RECT 100.760 140.470 101.040 140.840 ;
        RECT 100.770 139.875 101.030 139.965 ;
        RECT 100.370 139.735 101.030 139.875 ;
        RECT 100.370 139.285 100.510 139.735 ;
        RECT 100.770 139.645 101.030 139.735 ;
        RECT 100.310 138.965 100.570 139.285 ;
        RECT 100.370 135.205 100.510 138.965 ;
        RECT 100.770 138.625 101.030 138.945 ;
        RECT 100.830 136.905 100.970 138.625 ;
        RECT 100.770 136.585 101.030 136.905 ;
        RECT 99.850 134.885 100.110 135.205 ;
        RECT 100.310 134.885 100.570 135.205 ;
        RECT 98.930 132.165 99.190 132.485 ;
        RECT 99.390 132.165 99.650 132.485 ;
        RECT 98.470 129.445 98.730 129.765 ;
        RECT 98.010 128.425 98.270 128.745 ;
        RECT 98.470 128.425 98.730 128.745 ;
        RECT 98.070 127.045 98.210 128.425 ;
        RECT 98.010 126.725 98.270 127.045 ;
        RECT 98.530 126.365 98.670 128.425 ;
        RECT 98.010 126.275 98.270 126.365 ;
        RECT 97.610 126.135 98.270 126.275 ;
        RECT 98.010 126.045 98.270 126.135 ;
        RECT 98.470 126.045 98.730 126.365 ;
        RECT 95.250 125.365 95.510 125.685 ;
        RECT 97.090 125.025 97.350 125.345 ;
        RECT 94.910 124.490 96.790 124.860 ;
        RECT 94.910 119.050 96.790 119.420 ;
        RECT 97.150 118.205 97.290 125.025 ;
        RECT 97.550 120.265 97.810 120.585 ;
        RECT 97.610 118.885 97.750 120.265 ;
        RECT 98.070 119.905 98.210 126.045 ;
        RECT 98.530 122.965 98.670 126.045 ;
        RECT 98.470 122.645 98.730 122.965 ;
        RECT 98.010 119.585 98.270 119.905 ;
        RECT 98.070 118.885 98.210 119.585 ;
        RECT 97.550 118.565 97.810 118.885 ;
        RECT 98.010 118.565 98.270 118.885 ;
        RECT 97.090 117.885 97.350 118.205 ;
        RECT 98.530 117.865 98.670 122.645 ;
        RECT 99.390 122.305 99.650 122.625 ;
        RECT 99.450 120.585 99.590 122.305 ;
        RECT 99.390 120.265 99.650 120.585 ;
        RECT 98.930 119.925 99.190 120.245 ;
        RECT 98.990 118.545 99.130 119.925 ;
        RECT 99.450 118.545 99.590 120.265 ;
        RECT 98.930 118.225 99.190 118.545 ;
        RECT 99.390 118.225 99.650 118.545 ;
        RECT 98.470 117.545 98.730 117.865 ;
        RECT 94.910 113.610 96.790 113.980 ;
        RECT 99.910 112.765 100.050 134.885 ;
        RECT 101.290 134.865 101.430 141.435 ;
        RECT 101.690 140.160 101.950 140.305 ;
        RECT 101.680 139.790 101.960 140.160 ;
        RECT 101.230 134.545 101.490 134.865 ;
        RECT 100.770 134.095 101.030 134.185 ;
        RECT 101.750 134.095 101.890 139.790 ;
        RECT 102.150 138.625 102.410 138.945 ;
        RECT 102.210 134.865 102.350 138.625 ;
        RECT 102.150 134.545 102.410 134.865 ;
        RECT 100.770 133.955 101.890 134.095 ;
        RECT 100.770 133.865 101.030 133.955 ;
        RECT 101.690 131.145 101.950 131.465 ;
        RECT 100.310 128.765 100.570 129.085 ;
        RECT 100.370 122.625 100.510 128.765 ;
        RECT 101.750 128.745 101.890 131.145 ;
        RECT 101.690 128.425 101.950 128.745 ;
        RECT 101.750 126.025 101.890 128.425 ;
        RECT 101.690 125.705 101.950 126.025 ;
        RECT 100.310 122.305 100.570 122.625 ;
        RECT 100.370 118.205 100.510 122.305 ;
        RECT 100.310 117.885 100.570 118.205 ;
        RECT 102.150 116.865 102.410 117.185 ;
        RECT 102.210 115.145 102.350 116.865 ;
        RECT 102.150 114.825 102.410 115.145 ;
        RECT 102.670 112.765 102.810 144.405 ;
        RECT 103.130 139.965 103.270 145.085 ;
        RECT 104.970 142.595 105.110 147.805 ;
        RECT 105.370 142.595 105.630 142.685 ;
        RECT 104.970 142.455 105.630 142.595 ;
        RECT 105.370 142.365 105.630 142.455 ;
        RECT 104.910 141.345 105.170 141.665 ;
        RECT 103.070 139.645 103.330 139.965 ;
        RECT 104.970 139.625 105.110 141.345 ;
        RECT 105.430 140.645 105.570 142.365 ;
        RECT 105.370 140.325 105.630 140.645 ;
        RECT 104.910 139.305 105.170 139.625 ;
        RECT 104.450 138.625 104.710 138.945 ;
        RECT 103.990 137.605 104.250 137.925 ;
        RECT 104.050 135.205 104.190 137.605 ;
        RECT 104.510 136.565 104.650 138.625 ;
        RECT 104.450 136.245 104.710 136.565 ;
        RECT 104.970 135.205 105.110 139.305 ;
        RECT 103.990 134.885 104.250 135.205 ;
        RECT 104.910 134.885 105.170 135.205 ;
        RECT 105.430 134.185 105.570 140.325 ;
        RECT 105.370 133.865 105.630 134.185 ;
        RECT 105.890 133.845 106.030 169.225 ;
        RECT 107.730 169.205 107.870 180.105 ;
        RECT 108.130 178.065 108.390 178.385 ;
        RECT 108.190 176.005 108.330 178.065 ;
        RECT 109.050 176.705 109.310 177.025 ;
        RECT 108.130 175.685 108.390 176.005 ;
        RECT 108.590 175.405 108.850 175.665 ;
        RECT 108.190 175.345 108.850 175.405 ;
        RECT 108.190 175.265 108.790 175.345 ;
        RECT 109.110 175.325 109.250 176.705 ;
        RECT 107.670 168.885 107.930 169.205 ;
        RECT 107.210 155.625 107.470 155.945 ;
        RECT 106.290 155.285 106.550 155.605 ;
        RECT 106.350 152.885 106.490 155.285 ;
        RECT 107.270 154.245 107.410 155.625 ;
        RECT 107.210 153.925 107.470 154.245 ;
        RECT 106.290 152.565 106.550 152.885 ;
        RECT 107.670 148.485 107.930 148.805 ;
        RECT 106.290 147.125 106.550 147.445 ;
        RECT 106.350 145.745 106.490 147.125 ;
        RECT 106.290 145.425 106.550 145.745 ;
        RECT 106.350 142.345 106.490 145.425 ;
        RECT 107.210 145.085 107.470 145.405 ;
        RECT 107.270 142.345 107.410 145.085 ;
        RECT 106.290 142.025 106.550 142.345 ;
        RECT 107.210 142.025 107.470 142.345 ;
        RECT 105.830 133.525 106.090 133.845 ;
        RECT 106.750 130.465 107.010 130.785 ;
        RECT 106.810 129.085 106.950 130.465 ;
        RECT 106.750 128.765 107.010 129.085 ;
        RECT 103.530 128.425 103.790 128.745 ;
        RECT 103.590 127.045 103.730 128.425 ;
        RECT 104.910 127.745 105.170 128.065 ;
        RECT 103.530 126.725 103.790 127.045 ;
        RECT 104.970 124.325 105.110 127.745 ;
        RECT 106.810 124.405 106.950 128.765 ;
        RECT 107.210 127.745 107.470 128.065 ;
        RECT 107.270 125.685 107.410 127.745 ;
        RECT 107.210 125.365 107.470 125.685 ;
        RECT 104.910 124.005 105.170 124.325 ;
        RECT 106.350 124.265 106.950 124.405 ;
        RECT 106.350 118.205 106.490 124.265 ;
        RECT 106.750 123.665 107.010 123.985 ;
        RECT 106.810 118.885 106.950 123.665 ;
        RECT 107.210 120.265 107.470 120.585 ;
        RECT 106.750 118.565 107.010 118.885 ;
        RECT 106.290 117.885 106.550 118.205 ;
        RECT 107.270 116.165 107.410 120.265 ;
        RECT 107.210 115.845 107.470 116.165 ;
        RECT 105.370 115.505 105.630 115.825 ;
        RECT 105.430 113.105 105.570 115.505 ;
        RECT 107.730 115.145 107.870 148.485 ;
        RECT 108.190 146.085 108.330 175.265 ;
        RECT 109.050 175.005 109.310 175.325 ;
        RECT 109.570 174.985 109.710 185.885 ;
        RECT 114.170 183.145 114.310 188.265 ;
        RECT 114.110 182.825 114.370 183.145 ;
        RECT 112.730 182.145 112.990 182.465 ;
        RECT 109.910 181.610 111.790 181.980 ;
        RECT 112.790 181.445 112.930 182.145 ;
        RECT 112.730 181.125 112.990 181.445 ;
        RECT 110.430 180.105 110.690 180.425 ;
        RECT 110.490 178.725 110.630 180.105 ;
        RECT 110.430 178.405 110.690 178.725 ;
        RECT 109.910 176.170 111.790 176.540 ;
        RECT 109.510 174.665 109.770 174.985 ;
        RECT 110.430 174.840 110.690 174.985 ;
        RECT 110.420 174.470 110.700 174.840 ;
        RECT 111.810 174.665 112.070 174.985 ;
        RECT 111.870 172.265 112.010 174.665 ;
        RECT 112.270 173.985 112.530 174.305 ;
        RECT 112.330 172.945 112.470 173.985 ;
        RECT 135.630 173.380 136.780 174.600 ;
        RECT 112.270 172.625 112.530 172.945 ;
        RECT 111.810 171.945 112.070 172.265 ;
        RECT 113.650 171.945 113.910 172.265 ;
        RECT 109.910 170.730 111.790 171.100 ;
        RECT 108.590 169.225 108.850 169.545 ;
        RECT 108.650 159.685 108.790 169.225 ;
        RECT 109.510 168.885 109.770 169.205 ;
        RECT 109.570 166.825 109.710 168.885 ;
        RECT 112.270 167.185 112.530 167.505 ;
        RECT 109.510 166.505 109.770 166.825 ;
        RECT 109.570 164.355 109.710 166.505 ;
        RECT 109.910 165.290 111.790 165.660 ;
        RECT 109.970 164.355 110.230 164.445 ;
        RECT 109.570 164.215 110.230 164.355 ;
        RECT 109.970 164.125 110.230 164.215 ;
        RECT 109.910 159.850 111.790 160.220 ;
        RECT 112.330 159.685 112.470 167.185 ;
        RECT 113.710 166.825 113.850 171.945 ;
        RECT 133.750 170.070 134.880 172.730 ;
        RECT 115.950 169.400 116.210 169.545 ;
        RECT 115.940 169.030 116.220 169.400 ;
        RECT 113.650 166.505 113.910 166.825 ;
        RECT 135.630 166.640 136.740 173.380 ;
        RECT 135.630 165.420 136.780 166.640 ;
        RECT 113.190 163.785 113.450 164.105 ;
        RECT 113.250 162.405 113.390 163.785 ;
        RECT 113.190 162.085 113.450 162.405 ;
        RECT 108.590 159.365 108.850 159.685 ;
        RECT 112.270 159.365 112.530 159.685 ;
        RECT 108.650 156.285 108.790 159.365 ;
        RECT 108.590 155.965 108.850 156.285 ;
        RECT 109.510 154.945 109.770 155.265 ;
        RECT 109.570 153.225 109.710 154.945 ;
        RECT 109.910 154.410 111.790 154.780 ;
        RECT 109.510 152.905 109.770 153.225 ;
        RECT 112.270 152.225 112.530 152.545 ;
        RECT 112.330 151.185 112.470 152.225 ;
        RECT 112.270 150.865 112.530 151.185 ;
        RECT 109.910 148.970 111.790 149.340 ;
        RECT 112.730 147.805 112.990 148.125 ;
        RECT 112.270 147.465 112.530 147.785 ;
        RECT 108.590 147.125 108.850 147.445 ;
        RECT 108.650 146.085 108.790 147.125 ;
        RECT 109.970 146.785 110.230 147.105 ;
        RECT 108.130 145.765 108.390 146.085 ;
        RECT 108.590 145.765 108.850 146.085 ;
        RECT 110.030 145.405 110.170 146.785 ;
        RECT 112.330 146.085 112.470 147.465 ;
        RECT 112.270 145.765 112.530 146.085 ;
        RECT 109.970 145.085 110.230 145.405 ;
        RECT 109.910 143.530 111.790 143.900 ;
        RECT 109.050 141.345 109.310 141.665 ;
        RECT 109.510 141.345 109.770 141.665 ;
        RECT 109.110 136.225 109.250 141.345 ;
        RECT 109.570 140.305 109.710 141.345 ;
        RECT 109.510 139.985 109.770 140.305 ;
        RECT 112.270 139.305 112.530 139.625 ;
        RECT 109.910 138.090 111.790 138.460 ;
        RECT 112.330 137.925 112.470 139.305 ;
        RECT 112.270 137.605 112.530 137.925 ;
        RECT 109.510 136.925 109.770 137.245 ;
        RECT 109.050 135.905 109.310 136.225 ;
        RECT 109.570 135.205 109.710 136.925 ;
        RECT 109.510 134.885 109.770 135.205 ;
        RECT 112.790 134.425 112.930 147.805 ;
        RECT 114.110 147.465 114.370 147.785 ;
        RECT 114.170 139.625 114.310 147.465 ;
        RECT 135.630 141.200 136.780 141.270 ;
        RECT 135.630 140.180 136.800 141.200 ;
        RECT 114.110 139.305 114.370 139.625 ;
        RECT 114.170 137.245 114.310 139.305 ;
        RECT 132.560 138.140 135.160 140.060 ;
        RECT 114.110 136.925 114.370 137.245 ;
        RECT 112.330 134.285 112.930 134.425 ;
        RECT 109.910 132.650 111.790 133.020 ;
        RECT 109.510 127.745 109.770 128.065 ;
        RECT 109.570 126.365 109.710 127.745 ;
        RECT 109.910 127.210 111.790 127.580 ;
        RECT 109.510 126.045 109.770 126.365 ;
        RECT 109.910 121.770 111.790 122.140 ;
        RECT 109.050 120.605 109.310 120.925 ;
        RECT 109.110 118.545 109.250 120.605 ;
        RECT 109.050 118.225 109.310 118.545 ;
        RECT 107.670 114.825 107.930 115.145 ;
        RECT 108.130 114.825 108.390 115.145 ;
        RECT 105.830 114.145 106.090 114.465 ;
        RECT 105.370 112.785 105.630 113.105 ;
        RECT 90.190 112.445 90.450 112.765 ;
        RECT 94.330 112.445 94.590 112.765 ;
        RECT 99.850 112.445 100.110 112.765 ;
        RECT 102.610 112.445 102.870 112.765 ;
        RECT 103.990 112.105 104.250 112.425 ;
        RECT 91.110 111.425 91.370 111.745 ;
        RECT 96.630 111.425 96.890 111.745 ;
        RECT 101.230 111.425 101.490 111.745 ;
        RECT 103.530 111.425 103.790 111.745 ;
        RECT 86.970 110.405 87.230 110.725 ;
        RECT 87.030 110.125 87.170 110.405 ;
        RECT 81.910 109.725 82.170 110.045 ;
        RECT 86.050 109.725 86.310 110.045 ;
        RECT 87.030 109.985 87.630 110.125 ;
        RECT 74.550 109.385 74.810 109.705 ;
        RECT 73.630 108.705 73.890 109.025 ;
        RECT 72.250 107.345 72.510 107.665 ;
        RECT 72.710 107.345 72.970 107.665 ;
        RECT 73.690 107.325 73.830 108.705 ;
        RECT 74.610 108.005 74.750 109.385 ;
        RECT 74.550 107.685 74.810 108.005 ;
        RECT 73.630 107.005 73.890 107.325 ;
        RECT 75.470 107.005 75.730 107.325 ;
        RECT 71.790 105.985 72.050 106.305 ;
        RECT 75.530 104.265 75.670 107.005 ;
        RECT 76.850 106.665 77.110 106.985 ;
        RECT 81.970 106.825 82.110 109.725 ;
        RECT 84.210 109.045 84.470 109.365 ;
        RECT 81.970 106.685 82.570 106.825 ;
        RECT 75.470 103.945 75.730 104.265 ;
        RECT 76.910 92.050 77.050 106.665 ;
        RECT 79.910 105.450 81.790 105.820 ;
        RECT 82.430 92.050 82.570 106.685 ;
        RECT 84.270 105.285 84.410 109.045 ;
        RECT 87.490 107.325 87.630 109.985 ;
        RECT 88.810 107.345 89.070 107.665 ;
        RECT 87.430 107.005 87.690 107.325 ;
        RECT 87.890 106.665 88.150 106.985 ;
        RECT 84.210 104.965 84.470 105.285 ;
        RECT 87.950 92.050 88.090 106.665 ;
        RECT 88.870 105.285 89.010 107.345 ;
        RECT 91.170 106.305 91.310 111.425 ;
        RECT 96.690 110.045 96.830 111.425 ;
        RECT 92.950 109.725 93.210 110.045 ;
        RECT 96.630 109.725 96.890 110.045 ;
        RECT 93.010 109.445 93.150 109.725 ;
        RECT 93.010 109.305 93.610 109.445 ;
        RECT 100.770 109.385 101.030 109.705 ;
        RECT 91.110 105.985 91.370 106.305 ;
        RECT 88.810 104.965 89.070 105.285 ;
        RECT 93.470 92.050 93.610 109.305 ;
        RECT 98.930 109.045 99.190 109.365 ;
        RECT 94.910 108.170 96.790 108.540 ;
        RECT 98.990 108.005 99.130 109.045 ;
        RECT 100.830 108.005 100.970 109.385 ;
        RECT 98.930 107.685 99.190 108.005 ;
        RECT 100.770 107.685 101.030 108.005 ;
        RECT 101.290 107.405 101.430 111.425 ;
        RECT 101.690 109.385 101.950 109.705 ;
        RECT 98.470 107.005 98.730 107.325 ;
        RECT 100.830 107.265 101.430 107.405 ;
        RECT 98.530 105.285 98.670 107.005 ;
        RECT 100.310 106.665 100.570 106.985 ;
        RECT 98.470 104.965 98.730 105.285 ;
        RECT 98.930 104.285 99.190 104.605 ;
        RECT 94.910 102.730 96.790 103.100 ;
        RECT 98.990 92.050 99.130 104.285 ;
        RECT 100.370 103.925 100.510 106.665 ;
        RECT 100.830 104.605 100.970 107.265 ;
        RECT 101.750 106.725 101.890 109.385 ;
        RECT 101.750 106.585 102.350 106.725 ;
        RECT 102.210 104.605 102.350 106.585 ;
        RECT 103.590 106.305 103.730 111.425 ;
        RECT 104.050 109.705 104.190 112.105 ;
        RECT 105.890 110.045 106.030 114.145 ;
        RECT 105.830 109.725 106.090 110.045 ;
        RECT 103.990 109.385 104.250 109.705 ;
        RECT 108.190 106.985 108.330 114.825 ;
        RECT 108.590 114.145 108.850 114.465 ;
        RECT 108.650 113.105 108.790 114.145 ;
        RECT 108.590 112.785 108.850 113.105 ;
        RECT 109.110 112.425 109.250 118.225 ;
        RECT 109.910 116.330 111.790 116.700 ;
        RECT 112.330 115.145 112.470 134.285 ;
        RECT 114.170 126.365 114.310 136.925 ;
        RECT 135.640 133.320 136.800 140.180 ;
        RECT 113.190 126.045 113.450 126.365 ;
        RECT 114.110 126.045 114.370 126.365 ;
        RECT 113.250 123.645 113.390 126.045 ;
        RECT 113.190 123.325 113.450 123.645 ;
        RECT 113.250 120.925 113.390 123.325 ;
        RECT 113.190 120.605 113.450 120.925 ;
        RECT 112.270 114.825 112.530 115.145 ;
        RECT 109.050 112.105 109.310 112.425 ;
        RECT 115.490 112.105 115.750 112.425 ;
        RECT 108.590 109.045 108.850 109.365 ;
        RECT 104.450 106.665 104.710 106.985 ;
        RECT 108.130 106.665 108.390 106.985 ;
        RECT 103.530 105.985 103.790 106.305 ;
        RECT 100.770 104.285 101.030 104.605 ;
        RECT 102.150 104.285 102.410 104.605 ;
        RECT 100.310 103.605 100.570 103.925 ;
        RECT 104.510 92.050 104.650 106.665 ;
        RECT 108.190 104.265 108.330 106.665 ;
        RECT 108.650 105.285 108.790 109.045 ;
        RECT 109.110 106.985 109.250 112.105 ;
        RECT 109.910 110.890 111.790 111.260 ;
        RECT 109.510 108.705 109.770 109.025 ;
        RECT 109.050 106.665 109.310 106.985 ;
        RECT 108.590 104.965 108.850 105.285 ;
        RECT 109.570 104.685 109.710 108.705 ;
        RECT 109.910 105.450 111.790 105.820 ;
        RECT 109.570 104.545 110.170 104.685 ;
        RECT 108.130 103.945 108.390 104.265 ;
        RECT 110.030 92.050 110.170 104.545 ;
        RECT 113.190 103.265 113.450 103.585 ;
        RECT 113.250 102.565 113.390 103.265 ;
        RECT 113.190 102.245 113.450 102.565 ;
        RECT 115.550 92.050 115.690 112.105 ;
        RECT 119.160 106.470 119.440 106.840 ;
        RECT 119.230 104.265 119.370 106.470 ;
        RECT 129.750 105.580 133.160 106.650 ;
        RECT 119.170 103.945 119.430 104.265 ;
        RECT 64.490 91.625 65.550 91.765 ;
        RECT 65.800 90.050 66.080 92.050 ;
        RECT 71.320 90.050 71.600 92.050 ;
        RECT 76.840 90.050 77.120 92.050 ;
        RECT 82.360 90.050 82.640 92.050 ;
        RECT 87.880 90.050 88.160 92.050 ;
        RECT 93.400 90.050 93.680 92.050 ;
        RECT 98.920 90.050 99.200 92.050 ;
        RECT 104.440 90.050 104.720 92.050 ;
        RECT 109.960 90.050 110.240 92.050 ;
        RECT 115.480 90.050 115.760 92.050 ;
        RECT 13.920 85.550 15.140 89.420 ;
        RECT 19.910 85.980 21.130 89.850 ;
        RECT 67.730 89.640 68.670 89.840 ;
        RECT 25.730 85.120 26.950 88.990 ;
        RECT 31.780 85.510 33.000 89.380 ;
        RECT 37.750 88.780 38.970 89.290 ;
        RECT 37.680 88.620 38.970 88.780 ;
        RECT 43.810 88.630 45.030 89.530 ;
        RECT 49.740 88.640 50.960 89.040 ;
        RECT 37.680 86.810 39.070 88.620 ;
        RECT 37.750 85.420 38.970 86.810 ;
        RECT 43.810 86.720 45.140 88.630 ;
        RECT 49.740 86.920 51.010 88.640 ;
        RECT 43.810 85.660 45.030 86.720 ;
        RECT 49.740 85.170 50.960 86.920 ;
        RECT 55.530 85.320 56.750 89.190 ;
        RECT 61.720 88.640 62.940 88.870 ;
        RECT 61.720 86.600 63.130 88.640 ;
        RECT 61.720 85.000 62.940 86.600 ;
        RECT 67.580 85.770 68.800 89.640 ;
        RECT 73.850 84.290 75.070 88.160 ;
        RECT 79.730 84.310 80.950 88.180 ;
        RECT 74.090 80.440 74.370 84.290 ;
        RECT 20.140 80.160 74.370 80.440 ;
        RECT 20.140 75.650 20.420 80.160 ;
        RECT 80.070 79.800 80.350 84.310 ;
        RECT 85.470 84.100 86.690 87.970 ;
        RECT 91.460 84.500 92.680 88.320 ;
        RECT 97.600 84.630 98.820 88.240 ;
        RECT 103.650 84.740 104.870 88.610 ;
        RECT 109.620 85.420 110.840 89.290 ;
        RECT 115.740 85.700 116.960 89.570 ;
        RECT 121.520 85.700 122.740 89.570 ;
        RECT 31.380 79.520 80.350 79.800 ;
        RECT 31.380 75.850 31.660 79.520 ;
        RECT 86.050 79.170 86.330 84.100 ;
        RECT 42.510 78.890 86.330 79.170 ;
        RECT 3.960 71.320 6.050 73.240 ;
        RECT 19.330 73.120 21.890 75.650 ;
        RECT 28.185 73.180 30.255 74.460 ;
        RECT 30.670 73.320 33.230 75.850 ;
        RECT 42.510 75.750 42.790 78.890 ;
        RECT 92.030 78.570 92.310 84.500 ;
        RECT 53.830 78.290 92.310 78.570 ;
        RECT 53.830 75.820 54.110 78.290 ;
        RECT 98.010 77.990 98.290 84.630 ;
        RECT 64.900 77.710 98.290 77.990 ;
        RECT 19.005 71.800 19.865 72.640 ;
        RECT 15.560 68.610 16.990 71.210 ;
        RECT 19.305 68.570 19.845 71.800 ;
        RECT 20.145 70.600 20.555 73.120 ;
        RECT 30.205 71.810 31.065 72.650 ;
        RECT 19.325 47.770 19.825 68.570 ;
        RECT 20.165 49.090 20.555 70.600 ;
        RECT 20.955 70.010 21.845 70.740 ;
        RECT 21.055 65.190 21.315 70.010 ;
        RECT 22.695 68.620 25.405 69.470 ;
        RECT 22.895 65.840 24.825 68.620 ;
        RECT 30.505 68.580 31.045 71.810 ;
        RECT 31.345 70.610 31.755 73.320 ;
        RECT 39.475 73.150 41.545 74.430 ;
        RECT 41.910 73.220 44.470 75.750 ;
        RECT 41.425 71.780 42.285 72.620 ;
        RECT 27.795 67.130 28.915 67.810 ;
        RECT 28.075 65.850 28.745 67.130 ;
        RECT 21.455 65.460 26.505 65.840 ;
        RECT 27.865 65.440 28.915 65.850 ;
        RECT 21.055 63.640 21.435 65.190 ;
        RECT 21.175 55.800 21.435 63.640 ;
        RECT 26.485 63.200 26.755 65.240 ;
        RECT 27.615 63.200 27.885 65.200 ;
        RECT 26.485 56.510 27.885 63.200 ;
        RECT 21.085 55.290 21.445 55.800 ;
        RECT 21.065 54.860 21.445 55.290 ;
        RECT 26.485 55.190 26.755 56.510 ;
        RECT 27.615 55.150 27.885 56.510 ;
        RECT 28.885 55.260 29.205 65.190 ;
        RECT 28.885 55.200 29.215 55.260 ;
        RECT 21.065 54.580 21.315 54.860 ;
        RECT 20.865 54.180 25.505 54.580 ;
        RECT 26.405 54.290 27.535 54.300 ;
        RECT 28.895 54.290 29.215 55.200 ;
        RECT 21.065 52.060 21.315 54.180 ;
        RECT 25.765 53.490 26.125 54.110 ;
        RECT 25.845 52.610 26.105 53.490 ;
        RECT 26.385 53.240 29.215 54.290 ;
        RECT 25.675 52.230 26.205 52.610 ;
        RECT 21.065 51.970 21.565 52.060 ;
        RECT 21.055 51.240 21.565 51.970 ;
        RECT 21.295 50.240 21.565 51.240 ;
        RECT 22.205 50.990 22.475 51.940 ;
        RECT 22.205 50.840 22.675 50.990 ;
        RECT 22.205 50.160 22.765 50.840 ;
        RECT 22.285 50.150 22.765 50.160 ;
        RECT 21.575 49.620 22.195 49.980 ;
        RECT 21.615 49.090 22.045 49.620 ;
        RECT 20.165 48.670 22.045 49.090 ;
        RECT 22.535 48.960 22.765 50.150 ;
        RECT 21.615 47.800 22.045 48.670 ;
        RECT 22.455 48.360 22.835 48.960 ;
        RECT 19.325 47.060 20.015 47.770 ;
        RECT 21.435 47.440 22.055 47.800 ;
        RECT 21.135 47.060 21.425 47.250 ;
        RECT 19.325 46.620 21.425 47.060 ;
        RECT 19.325 46.600 20.015 46.620 ;
        RECT 21.135 46.380 21.425 46.620 ;
        RECT 22.055 46.990 22.325 47.240 ;
        RECT 22.535 46.990 22.765 48.360 ;
        RECT 25.355 47.010 25.685 52.030 ;
        RECT 26.405 52.020 27.535 53.240 ;
        RECT 28.895 53.220 29.215 53.240 ;
        RECT 22.055 46.880 22.765 46.990 ;
        RECT 25.345 46.960 25.685 47.010 ;
        RECT 26.235 47.780 27.615 52.020 ;
        RECT 22.055 46.570 22.715 46.880 ;
        RECT 22.055 46.400 22.325 46.570 ;
        RECT 25.345 45.000 25.625 46.960 ;
        RECT 26.235 46.920 26.535 47.780 ;
        RECT 27.315 46.920 27.615 47.780 ;
        RECT 28.165 46.920 28.495 51.990 ;
        RECT 27.565 46.380 28.045 46.760 ;
        RECT 27.665 45.760 27.915 46.380 ;
        RECT 27.565 45.160 27.945 45.760 ;
        RECT 24.825 44.230 25.925 45.000 ;
        RECT 28.215 44.930 28.495 46.920 ;
        RECT 30.525 47.780 31.025 68.580 ;
        RECT 31.365 49.100 31.755 70.610 ;
        RECT 32.155 70.020 33.045 70.750 ;
        RECT 32.255 65.200 32.515 70.020 ;
        RECT 33.895 68.630 36.605 69.480 ;
        RECT 34.095 65.850 36.025 68.630 ;
        RECT 41.725 68.550 42.265 71.780 ;
        RECT 42.565 70.580 42.975 73.220 ;
        RECT 50.055 73.090 52.125 74.370 ;
        RECT 53.150 73.290 55.710 75.820 ;
        RECT 64.900 75.810 65.180 77.710 ;
        RECT 103.990 77.230 104.270 84.740 ;
        RECT 76.140 76.950 104.270 77.230 ;
        RECT 52.675 71.760 53.535 72.600 ;
        RECT 38.995 67.140 40.115 67.820 ;
        RECT 39.275 65.860 39.945 67.140 ;
        RECT 32.655 65.470 37.705 65.850 ;
        RECT 39.065 65.450 40.115 65.860 ;
        RECT 32.255 63.650 32.635 65.200 ;
        RECT 32.375 55.810 32.635 63.650 ;
        RECT 37.685 63.210 37.955 65.250 ;
        RECT 38.815 63.210 39.085 65.210 ;
        RECT 37.685 56.520 39.085 63.210 ;
        RECT 32.285 55.300 32.645 55.810 ;
        RECT 32.265 54.870 32.645 55.300 ;
        RECT 37.685 55.200 37.955 56.520 ;
        RECT 38.815 55.160 39.085 56.520 ;
        RECT 40.085 55.270 40.405 65.200 ;
        RECT 40.085 55.210 40.415 55.270 ;
        RECT 32.265 54.590 32.515 54.870 ;
        RECT 32.065 54.190 36.705 54.590 ;
        RECT 37.605 54.300 38.735 54.310 ;
        RECT 40.095 54.300 40.415 55.210 ;
        RECT 32.265 52.070 32.515 54.190 ;
        RECT 36.965 53.500 37.325 54.120 ;
        RECT 37.045 52.620 37.305 53.500 ;
        RECT 37.585 53.250 40.415 54.300 ;
        RECT 36.875 52.240 37.405 52.620 ;
        RECT 32.265 51.980 32.765 52.070 ;
        RECT 32.255 51.250 32.765 51.980 ;
        RECT 32.495 50.250 32.765 51.250 ;
        RECT 33.405 51.000 33.675 51.950 ;
        RECT 33.405 50.850 33.875 51.000 ;
        RECT 33.405 50.170 33.965 50.850 ;
        RECT 33.485 50.160 33.965 50.170 ;
        RECT 32.775 49.630 33.395 49.990 ;
        RECT 32.815 49.100 33.245 49.630 ;
        RECT 31.365 48.680 33.245 49.100 ;
        RECT 33.735 48.970 33.965 50.160 ;
        RECT 32.815 47.810 33.245 48.680 ;
        RECT 33.655 48.370 34.035 48.970 ;
        RECT 30.525 47.070 31.215 47.780 ;
        RECT 32.635 47.450 33.255 47.810 ;
        RECT 32.335 47.070 32.625 47.260 ;
        RECT 30.525 46.630 32.625 47.070 ;
        RECT 30.525 46.610 31.215 46.630 ;
        RECT 32.335 46.390 32.625 46.630 ;
        RECT 33.255 47.000 33.525 47.250 ;
        RECT 33.735 47.000 33.965 48.370 ;
        RECT 36.555 47.020 36.885 52.040 ;
        RECT 37.605 52.030 38.735 53.250 ;
        RECT 40.095 53.230 40.415 53.250 ;
        RECT 33.255 46.890 33.965 47.000 ;
        RECT 36.545 46.970 36.885 47.020 ;
        RECT 37.435 47.790 38.815 52.030 ;
        RECT 33.255 46.580 33.915 46.890 ;
        RECT 33.255 46.410 33.525 46.580 ;
        RECT 36.545 45.010 36.825 46.970 ;
        RECT 37.435 46.930 37.735 47.790 ;
        RECT 38.515 46.930 38.815 47.790 ;
        RECT 39.365 46.930 39.695 52.000 ;
        RECT 38.765 46.390 39.245 46.770 ;
        RECT 38.865 45.770 39.115 46.390 ;
        RECT 38.765 45.170 39.145 45.770 ;
        RECT 28.215 43.200 28.515 44.930 ;
        RECT 36.025 44.240 37.125 45.010 ;
        RECT 39.415 44.940 39.695 46.930 ;
        RECT 41.745 47.750 42.245 68.550 ;
        RECT 42.585 49.070 42.975 70.580 ;
        RECT 43.375 69.990 44.265 70.720 ;
        RECT 43.475 65.170 43.735 69.990 ;
        RECT 45.115 68.600 47.825 69.450 ;
        RECT 45.315 65.820 47.245 68.600 ;
        RECT 52.975 68.530 53.515 71.760 ;
        RECT 53.815 70.560 54.225 73.290 ;
        RECT 61.475 73.120 63.545 74.400 ;
        RECT 64.400 73.280 66.960 75.810 ;
        RECT 76.140 75.740 76.420 76.950 ;
        RECT 109.970 76.610 110.250 85.420 ;
        RECT 87.580 76.330 110.250 76.610 ;
        RECT 87.580 75.760 87.860 76.330 ;
        RECT 115.950 76.030 116.230 85.700 ;
        RECT 98.850 75.840 116.230 76.030 ;
        RECT 63.895 71.750 64.755 72.590 ;
        RECT 50.215 67.110 51.335 67.790 ;
        RECT 50.495 65.830 51.165 67.110 ;
        RECT 43.875 65.440 48.925 65.820 ;
        RECT 50.285 65.420 51.335 65.830 ;
        RECT 43.475 63.620 43.855 65.170 ;
        RECT 43.595 55.780 43.855 63.620 ;
        RECT 48.905 63.180 49.175 65.220 ;
        RECT 50.035 63.180 50.305 65.180 ;
        RECT 48.905 56.490 50.305 63.180 ;
        RECT 43.505 55.270 43.865 55.780 ;
        RECT 43.485 54.840 43.865 55.270 ;
        RECT 48.905 55.170 49.175 56.490 ;
        RECT 50.035 55.130 50.305 56.490 ;
        RECT 51.305 55.240 51.625 65.170 ;
        RECT 51.305 55.180 51.635 55.240 ;
        RECT 43.485 54.560 43.735 54.840 ;
        RECT 43.285 54.160 47.925 54.560 ;
        RECT 48.825 54.270 49.955 54.280 ;
        RECT 51.315 54.270 51.635 55.180 ;
        RECT 43.485 52.040 43.735 54.160 ;
        RECT 48.185 53.470 48.545 54.090 ;
        RECT 48.265 52.590 48.525 53.470 ;
        RECT 48.805 53.220 51.635 54.270 ;
        RECT 48.095 52.210 48.625 52.590 ;
        RECT 43.485 51.950 43.985 52.040 ;
        RECT 43.475 51.220 43.985 51.950 ;
        RECT 43.715 50.220 43.985 51.220 ;
        RECT 44.625 50.970 44.895 51.920 ;
        RECT 44.625 50.820 45.095 50.970 ;
        RECT 44.625 50.140 45.185 50.820 ;
        RECT 44.705 50.130 45.185 50.140 ;
        RECT 43.995 49.600 44.615 49.960 ;
        RECT 44.035 49.070 44.465 49.600 ;
        RECT 42.585 48.650 44.465 49.070 ;
        RECT 44.955 48.940 45.185 50.130 ;
        RECT 44.035 47.780 44.465 48.650 ;
        RECT 44.875 48.340 45.255 48.940 ;
        RECT 41.745 47.040 42.435 47.750 ;
        RECT 43.855 47.420 44.475 47.780 ;
        RECT 43.555 47.040 43.845 47.230 ;
        RECT 41.745 46.600 43.845 47.040 ;
        RECT 41.745 46.580 42.435 46.600 ;
        RECT 43.555 46.360 43.845 46.600 ;
        RECT 44.475 46.970 44.745 47.220 ;
        RECT 44.955 46.970 45.185 48.340 ;
        RECT 47.775 46.990 48.105 52.010 ;
        RECT 48.825 52.000 49.955 53.220 ;
        RECT 51.315 53.200 51.635 53.220 ;
        RECT 44.475 46.860 45.185 46.970 ;
        RECT 47.765 46.940 48.105 46.990 ;
        RECT 48.655 47.760 50.035 52.000 ;
        RECT 44.475 46.550 45.135 46.860 ;
        RECT 44.475 46.380 44.745 46.550 ;
        RECT 47.765 44.980 48.045 46.940 ;
        RECT 48.655 46.900 48.955 47.760 ;
        RECT 49.735 46.900 50.035 47.760 ;
        RECT 50.585 46.900 50.915 51.970 ;
        RECT 49.985 46.360 50.465 46.740 ;
        RECT 50.085 45.740 50.335 46.360 ;
        RECT 49.985 45.140 50.365 45.740 ;
        RECT 39.415 43.210 39.715 44.940 ;
        RECT 47.245 44.210 48.345 44.980 ;
        RECT 50.635 44.910 50.915 46.900 ;
        RECT 52.995 47.730 53.495 68.530 ;
        RECT 53.835 49.050 54.225 70.560 ;
        RECT 54.625 69.970 55.515 70.700 ;
        RECT 54.725 65.150 54.985 69.970 ;
        RECT 56.365 68.580 59.075 69.430 ;
        RECT 56.565 65.800 58.495 68.580 ;
        RECT 64.195 68.520 64.735 71.750 ;
        RECT 65.035 70.550 65.445 73.280 ;
        RECT 72.585 73.130 74.655 74.410 ;
        RECT 75.550 73.210 78.110 75.740 ;
        RECT 75.135 71.740 75.995 72.580 ;
        RECT 61.465 67.090 62.585 67.770 ;
        RECT 61.745 65.810 62.415 67.090 ;
        RECT 55.125 65.420 60.175 65.800 ;
        RECT 61.535 65.400 62.585 65.810 ;
        RECT 54.725 63.600 55.105 65.150 ;
        RECT 54.845 55.760 55.105 63.600 ;
        RECT 60.155 63.160 60.425 65.200 ;
        RECT 61.285 63.160 61.555 65.160 ;
        RECT 60.155 56.470 61.555 63.160 ;
        RECT 54.755 55.250 55.115 55.760 ;
        RECT 54.735 54.820 55.115 55.250 ;
        RECT 60.155 55.150 60.425 56.470 ;
        RECT 61.285 55.110 61.555 56.470 ;
        RECT 62.555 55.220 62.875 65.150 ;
        RECT 62.555 55.160 62.885 55.220 ;
        RECT 54.735 54.540 54.985 54.820 ;
        RECT 54.535 54.140 59.175 54.540 ;
        RECT 60.075 54.250 61.205 54.260 ;
        RECT 62.565 54.250 62.885 55.160 ;
        RECT 54.735 52.020 54.985 54.140 ;
        RECT 59.435 53.450 59.795 54.070 ;
        RECT 59.515 52.570 59.775 53.450 ;
        RECT 60.055 53.200 62.885 54.250 ;
        RECT 59.345 52.190 59.875 52.570 ;
        RECT 54.735 51.930 55.235 52.020 ;
        RECT 54.725 51.200 55.235 51.930 ;
        RECT 54.965 50.200 55.235 51.200 ;
        RECT 55.875 50.950 56.145 51.900 ;
        RECT 55.875 50.800 56.345 50.950 ;
        RECT 55.875 50.120 56.435 50.800 ;
        RECT 55.955 50.110 56.435 50.120 ;
        RECT 55.245 49.580 55.865 49.940 ;
        RECT 55.285 49.050 55.715 49.580 ;
        RECT 53.835 48.630 55.715 49.050 ;
        RECT 56.205 48.920 56.435 50.110 ;
        RECT 55.285 47.760 55.715 48.630 ;
        RECT 56.125 48.320 56.505 48.920 ;
        RECT 52.995 47.020 53.685 47.730 ;
        RECT 55.105 47.400 55.725 47.760 ;
        RECT 54.805 47.020 55.095 47.210 ;
        RECT 52.995 46.580 55.095 47.020 ;
        RECT 52.995 46.560 53.685 46.580 ;
        RECT 54.805 46.340 55.095 46.580 ;
        RECT 55.725 46.950 55.995 47.200 ;
        RECT 56.205 46.950 56.435 48.320 ;
        RECT 59.025 46.970 59.355 51.990 ;
        RECT 60.075 51.980 61.205 53.200 ;
        RECT 62.565 53.180 62.885 53.200 ;
        RECT 55.725 46.840 56.435 46.950 ;
        RECT 59.015 46.920 59.355 46.970 ;
        RECT 59.905 47.740 61.285 51.980 ;
        RECT 55.725 46.530 56.385 46.840 ;
        RECT 55.725 46.360 55.995 46.530 ;
        RECT 59.015 44.960 59.295 46.920 ;
        RECT 59.905 46.880 60.205 47.740 ;
        RECT 60.985 46.880 61.285 47.740 ;
        RECT 61.835 46.880 62.165 51.950 ;
        RECT 61.235 46.340 61.715 46.720 ;
        RECT 61.335 45.720 61.585 46.340 ;
        RECT 61.235 45.120 61.615 45.720 ;
        RECT 19.865 42.210 21.245 42.780 ;
        RECT 27.495 42.630 28.875 43.200 ;
        RECT 31.145 42.210 32.525 42.780 ;
        RECT 38.695 42.640 40.075 43.210 ;
        RECT 50.635 43.180 50.935 44.910 ;
        RECT 58.495 44.190 59.595 44.960 ;
        RECT 61.885 44.890 62.165 46.880 ;
        RECT 64.215 47.720 64.715 68.520 ;
        RECT 65.055 49.040 65.445 70.550 ;
        RECT 65.845 69.960 66.735 70.690 ;
        RECT 65.945 65.140 66.205 69.960 ;
        RECT 67.585 68.570 70.295 69.420 ;
        RECT 67.785 65.790 69.715 68.570 ;
        RECT 75.435 68.510 75.975 71.740 ;
        RECT 76.275 70.540 76.685 73.210 ;
        RECT 83.855 73.120 85.925 74.400 ;
        RECT 86.850 73.230 89.410 75.760 ;
        RECT 98.150 75.750 116.230 75.840 ;
        RECT 86.385 71.750 87.245 72.590 ;
        RECT 72.685 67.080 73.805 67.760 ;
        RECT 72.965 65.800 73.635 67.080 ;
        RECT 66.345 65.410 71.395 65.790 ;
        RECT 72.755 65.390 73.805 65.800 ;
        RECT 65.945 63.590 66.325 65.140 ;
        RECT 66.065 55.750 66.325 63.590 ;
        RECT 71.375 63.150 71.645 65.190 ;
        RECT 72.505 63.150 72.775 65.150 ;
        RECT 71.375 56.460 72.775 63.150 ;
        RECT 65.975 55.240 66.335 55.750 ;
        RECT 65.955 54.810 66.335 55.240 ;
        RECT 71.375 55.140 71.645 56.460 ;
        RECT 72.505 55.100 72.775 56.460 ;
        RECT 73.775 55.210 74.095 65.140 ;
        RECT 73.775 55.150 74.105 55.210 ;
        RECT 65.955 54.530 66.205 54.810 ;
        RECT 65.755 54.130 70.395 54.530 ;
        RECT 71.295 54.240 72.425 54.250 ;
        RECT 73.785 54.240 74.105 55.150 ;
        RECT 65.955 52.010 66.205 54.130 ;
        RECT 70.655 53.440 71.015 54.060 ;
        RECT 70.735 52.560 70.995 53.440 ;
        RECT 71.275 53.190 74.105 54.240 ;
        RECT 70.565 52.180 71.095 52.560 ;
        RECT 65.955 51.920 66.455 52.010 ;
        RECT 65.945 51.190 66.455 51.920 ;
        RECT 66.185 50.190 66.455 51.190 ;
        RECT 67.095 50.940 67.365 51.890 ;
        RECT 67.095 50.790 67.565 50.940 ;
        RECT 67.095 50.110 67.655 50.790 ;
        RECT 67.175 50.100 67.655 50.110 ;
        RECT 66.465 49.570 67.085 49.930 ;
        RECT 66.505 49.040 66.935 49.570 ;
        RECT 65.055 48.620 66.935 49.040 ;
        RECT 67.425 48.910 67.655 50.100 ;
        RECT 66.505 47.750 66.935 48.620 ;
        RECT 67.345 48.310 67.725 48.910 ;
        RECT 64.215 47.010 64.905 47.720 ;
        RECT 66.325 47.390 66.945 47.750 ;
        RECT 66.025 47.010 66.315 47.200 ;
        RECT 64.215 46.570 66.315 47.010 ;
        RECT 64.215 46.550 64.905 46.570 ;
        RECT 66.025 46.330 66.315 46.570 ;
        RECT 66.945 46.940 67.215 47.190 ;
        RECT 67.425 46.940 67.655 48.310 ;
        RECT 70.245 46.960 70.575 51.980 ;
        RECT 71.295 51.970 72.425 53.190 ;
        RECT 73.785 53.170 74.105 53.190 ;
        RECT 66.945 46.830 67.655 46.940 ;
        RECT 70.235 46.910 70.575 46.960 ;
        RECT 71.125 47.730 72.505 51.970 ;
        RECT 66.945 46.520 67.605 46.830 ;
        RECT 66.945 46.350 67.215 46.520 ;
        RECT 70.235 44.950 70.515 46.910 ;
        RECT 71.125 46.870 71.425 47.730 ;
        RECT 72.205 46.870 72.505 47.730 ;
        RECT 73.055 46.870 73.385 51.940 ;
        RECT 72.455 46.330 72.935 46.710 ;
        RECT 72.555 45.710 72.805 46.330 ;
        RECT 72.455 45.110 72.835 45.710 ;
        RECT 20.225 40.480 20.525 42.210 ;
        RECT 20.245 38.490 20.525 40.480 ;
        RECT 22.815 40.410 23.915 41.180 ;
        RECT 31.505 40.480 31.805 42.210 ;
        RECT 42.435 42.190 43.815 42.760 ;
        RECT 49.915 42.610 51.295 43.180 ;
        RECT 61.885 43.160 62.185 44.890 ;
        RECT 69.715 44.180 70.815 44.950 ;
        RECT 73.105 44.880 73.385 46.870 ;
        RECT 75.455 47.710 75.955 68.510 ;
        RECT 76.295 49.030 76.685 70.540 ;
        RECT 77.085 69.950 77.975 70.680 ;
        RECT 77.185 65.130 77.445 69.950 ;
        RECT 78.825 68.560 81.535 69.410 ;
        RECT 79.025 65.780 80.955 68.560 ;
        RECT 86.685 68.520 87.225 71.750 ;
        RECT 87.525 70.550 87.935 73.230 ;
        RECT 95.045 73.060 97.115 74.340 ;
        RECT 98.150 73.310 100.710 75.750 ;
        RECT 109.390 75.480 111.950 75.560 ;
        RECT 121.930 75.480 122.210 85.700 ;
        RECT 127.550 85.510 128.770 89.380 ;
        RECT 127.910 76.040 128.190 85.510 ;
        RECT 133.380 76.580 136.010 77.880 ;
        RECT 137.240 76.560 139.870 77.860 ;
        RECT 109.390 75.200 122.210 75.480 ;
        RECT 97.665 71.740 98.525 72.580 ;
        RECT 83.925 67.070 85.045 67.750 ;
        RECT 84.205 65.790 84.875 67.070 ;
        RECT 77.585 65.400 82.635 65.780 ;
        RECT 83.995 65.380 85.045 65.790 ;
        RECT 77.185 63.580 77.565 65.130 ;
        RECT 77.305 55.740 77.565 63.580 ;
        RECT 82.615 63.140 82.885 65.180 ;
        RECT 83.745 63.140 84.015 65.140 ;
        RECT 82.615 56.450 84.015 63.140 ;
        RECT 77.215 55.230 77.575 55.740 ;
        RECT 77.195 54.800 77.575 55.230 ;
        RECT 82.615 55.130 82.885 56.450 ;
        RECT 83.745 55.090 84.015 56.450 ;
        RECT 85.015 55.200 85.335 65.130 ;
        RECT 85.015 55.140 85.345 55.200 ;
        RECT 77.195 54.520 77.445 54.800 ;
        RECT 76.995 54.120 81.635 54.520 ;
        RECT 82.535 54.230 83.665 54.240 ;
        RECT 85.025 54.230 85.345 55.140 ;
        RECT 77.195 52.000 77.445 54.120 ;
        RECT 81.895 53.430 82.255 54.050 ;
        RECT 81.975 52.550 82.235 53.430 ;
        RECT 82.515 53.180 85.345 54.230 ;
        RECT 81.805 52.170 82.335 52.550 ;
        RECT 77.195 51.910 77.695 52.000 ;
        RECT 77.185 51.180 77.695 51.910 ;
        RECT 77.425 50.180 77.695 51.180 ;
        RECT 78.335 50.930 78.605 51.880 ;
        RECT 78.335 50.780 78.805 50.930 ;
        RECT 78.335 50.100 78.895 50.780 ;
        RECT 78.415 50.090 78.895 50.100 ;
        RECT 77.705 49.560 78.325 49.920 ;
        RECT 77.745 49.030 78.175 49.560 ;
        RECT 76.295 48.610 78.175 49.030 ;
        RECT 78.665 48.900 78.895 50.090 ;
        RECT 77.745 47.740 78.175 48.610 ;
        RECT 78.585 48.300 78.965 48.900 ;
        RECT 75.455 47.000 76.145 47.710 ;
        RECT 77.565 47.380 78.185 47.740 ;
        RECT 77.265 47.000 77.555 47.190 ;
        RECT 75.455 46.560 77.555 47.000 ;
        RECT 75.455 46.540 76.145 46.560 ;
        RECT 77.265 46.320 77.555 46.560 ;
        RECT 78.185 46.930 78.455 47.180 ;
        RECT 78.665 46.930 78.895 48.300 ;
        RECT 81.485 46.950 81.815 51.970 ;
        RECT 82.535 51.960 83.665 53.180 ;
        RECT 85.025 53.160 85.345 53.180 ;
        RECT 78.185 46.820 78.895 46.930 ;
        RECT 81.475 46.900 81.815 46.950 ;
        RECT 82.365 47.720 83.745 51.960 ;
        RECT 78.185 46.510 78.845 46.820 ;
        RECT 78.185 46.340 78.455 46.510 ;
        RECT 81.475 44.940 81.755 46.900 ;
        RECT 82.365 46.860 82.665 47.720 ;
        RECT 83.445 46.860 83.745 47.720 ;
        RECT 84.295 46.860 84.625 51.930 ;
        RECT 83.695 46.320 84.175 46.700 ;
        RECT 83.795 45.700 84.045 46.320 ;
        RECT 83.695 45.100 84.075 45.700 ;
        RECT 53.655 42.190 55.035 42.760 ;
        RECT 61.165 42.590 62.545 43.160 ;
        RECT 73.105 43.150 73.405 44.880 ;
        RECT 80.955 44.170 82.055 44.940 ;
        RECT 84.345 44.870 84.625 46.860 ;
        RECT 86.705 47.720 87.205 68.520 ;
        RECT 87.545 49.040 87.935 70.550 ;
        RECT 88.335 69.960 89.225 70.690 ;
        RECT 88.435 65.140 88.695 69.960 ;
        RECT 90.075 68.570 92.785 69.420 ;
        RECT 90.275 65.790 92.205 68.570 ;
        RECT 97.965 68.510 98.505 71.740 ;
        RECT 98.805 70.540 99.215 73.310 ;
        RECT 106.455 73.110 108.525 74.390 ;
        RECT 109.390 73.030 111.950 75.200 ;
        RECT 125.760 74.810 128.190 76.040 ;
        RECT 121.290 74.790 128.190 74.810 ;
        RECT 120.600 74.530 128.190 74.790 ;
        RECT 117.655 73.110 119.725 74.390 ;
        RECT 120.600 73.180 128.160 74.530 ;
        RECT 129.505 73.190 131.575 74.470 ;
        RECT 120.600 73.110 126.160 73.180 ;
        RECT 108.935 71.740 109.795 72.580 ;
        RECT 95.175 67.080 96.295 67.760 ;
        RECT 95.455 65.800 96.125 67.080 ;
        RECT 88.835 65.410 93.885 65.790 ;
        RECT 95.245 65.390 96.295 65.800 ;
        RECT 88.435 63.590 88.815 65.140 ;
        RECT 88.555 55.750 88.815 63.590 ;
        RECT 93.865 63.150 94.135 65.190 ;
        RECT 94.995 63.150 95.265 65.150 ;
        RECT 93.865 56.460 95.265 63.150 ;
        RECT 88.465 55.240 88.825 55.750 ;
        RECT 88.445 54.810 88.825 55.240 ;
        RECT 93.865 55.140 94.135 56.460 ;
        RECT 94.995 55.100 95.265 56.460 ;
        RECT 96.265 55.210 96.585 65.140 ;
        RECT 96.265 55.150 96.595 55.210 ;
        RECT 88.445 54.530 88.695 54.810 ;
        RECT 88.245 54.130 92.885 54.530 ;
        RECT 93.785 54.240 94.915 54.250 ;
        RECT 96.275 54.240 96.595 55.150 ;
        RECT 88.445 52.010 88.695 54.130 ;
        RECT 93.145 53.440 93.505 54.060 ;
        RECT 93.225 52.560 93.485 53.440 ;
        RECT 93.765 53.190 96.595 54.240 ;
        RECT 93.055 52.180 93.585 52.560 ;
        RECT 88.445 51.920 88.945 52.010 ;
        RECT 88.435 51.190 88.945 51.920 ;
        RECT 88.675 50.190 88.945 51.190 ;
        RECT 89.585 50.940 89.855 51.890 ;
        RECT 89.585 50.790 90.055 50.940 ;
        RECT 89.585 50.110 90.145 50.790 ;
        RECT 89.665 50.100 90.145 50.110 ;
        RECT 88.955 49.570 89.575 49.930 ;
        RECT 88.995 49.040 89.425 49.570 ;
        RECT 87.545 48.620 89.425 49.040 ;
        RECT 89.915 48.910 90.145 50.100 ;
        RECT 88.995 47.750 89.425 48.620 ;
        RECT 89.835 48.310 90.215 48.910 ;
        RECT 86.705 47.010 87.395 47.720 ;
        RECT 88.815 47.390 89.435 47.750 ;
        RECT 88.515 47.010 88.805 47.200 ;
        RECT 86.705 46.570 88.805 47.010 ;
        RECT 86.705 46.550 87.395 46.570 ;
        RECT 88.515 46.330 88.805 46.570 ;
        RECT 89.435 46.940 89.705 47.190 ;
        RECT 89.915 46.940 90.145 48.310 ;
        RECT 92.735 46.960 93.065 51.980 ;
        RECT 93.785 51.970 94.915 53.190 ;
        RECT 96.275 53.170 96.595 53.190 ;
        RECT 89.435 46.830 90.145 46.940 ;
        RECT 92.725 46.910 93.065 46.960 ;
        RECT 93.615 47.730 94.995 51.970 ;
        RECT 89.435 46.520 90.095 46.830 ;
        RECT 89.435 46.350 89.705 46.520 ;
        RECT 92.725 44.950 93.005 46.910 ;
        RECT 93.615 46.870 93.915 47.730 ;
        RECT 94.695 46.870 94.995 47.730 ;
        RECT 95.545 46.870 95.875 51.940 ;
        RECT 94.945 46.330 95.425 46.710 ;
        RECT 95.045 45.710 95.295 46.330 ;
        RECT 94.945 45.110 95.325 45.710 ;
        RECT 64.855 42.190 66.235 42.760 ;
        RECT 72.385 42.580 73.765 43.150 ;
        RECT 84.345 43.140 84.645 44.870 ;
        RECT 92.205 44.180 93.305 44.950 ;
        RECT 95.595 44.880 95.875 46.870 ;
        RECT 97.985 47.710 98.485 68.510 ;
        RECT 98.825 49.030 99.215 70.540 ;
        RECT 99.615 69.950 100.505 70.680 ;
        RECT 99.715 65.130 99.975 69.950 ;
        RECT 101.355 68.560 104.065 69.410 ;
        RECT 101.555 65.780 103.485 68.560 ;
        RECT 109.235 68.510 109.775 71.740 ;
        RECT 110.075 70.540 110.485 73.030 ;
        RECT 120.185 71.740 121.045 72.580 ;
        RECT 106.455 67.070 107.575 67.750 ;
        RECT 106.735 65.790 107.405 67.070 ;
        RECT 100.115 65.400 105.165 65.780 ;
        RECT 106.525 65.380 107.575 65.790 ;
        RECT 99.715 63.580 100.095 65.130 ;
        RECT 99.835 55.740 100.095 63.580 ;
        RECT 105.145 63.140 105.415 65.180 ;
        RECT 106.275 63.140 106.545 65.140 ;
        RECT 105.145 56.450 106.545 63.140 ;
        RECT 99.745 55.230 100.105 55.740 ;
        RECT 99.725 54.800 100.105 55.230 ;
        RECT 105.145 55.130 105.415 56.450 ;
        RECT 106.275 55.090 106.545 56.450 ;
        RECT 107.545 55.200 107.865 65.130 ;
        RECT 107.545 55.140 107.875 55.200 ;
        RECT 99.725 54.520 99.975 54.800 ;
        RECT 99.525 54.120 104.165 54.520 ;
        RECT 105.065 54.230 106.195 54.240 ;
        RECT 107.555 54.230 107.875 55.140 ;
        RECT 99.725 52.000 99.975 54.120 ;
        RECT 104.425 53.430 104.785 54.050 ;
        RECT 104.505 52.550 104.765 53.430 ;
        RECT 105.045 53.180 107.875 54.230 ;
        RECT 104.335 52.170 104.865 52.550 ;
        RECT 99.725 51.910 100.225 52.000 ;
        RECT 99.715 51.180 100.225 51.910 ;
        RECT 99.955 50.180 100.225 51.180 ;
        RECT 100.865 50.930 101.135 51.880 ;
        RECT 100.865 50.780 101.335 50.930 ;
        RECT 100.865 50.100 101.425 50.780 ;
        RECT 100.945 50.090 101.425 50.100 ;
        RECT 100.235 49.560 100.855 49.920 ;
        RECT 100.275 49.030 100.705 49.560 ;
        RECT 98.825 48.610 100.705 49.030 ;
        RECT 101.195 48.900 101.425 50.090 ;
        RECT 100.275 47.740 100.705 48.610 ;
        RECT 101.115 48.300 101.495 48.900 ;
        RECT 97.985 47.000 98.675 47.710 ;
        RECT 100.095 47.380 100.715 47.740 ;
        RECT 99.795 47.000 100.085 47.190 ;
        RECT 97.985 46.560 100.085 47.000 ;
        RECT 97.985 46.540 98.675 46.560 ;
        RECT 99.795 46.320 100.085 46.560 ;
        RECT 100.715 46.930 100.985 47.180 ;
        RECT 101.195 46.930 101.425 48.300 ;
        RECT 104.015 46.950 104.345 51.970 ;
        RECT 105.065 51.960 106.195 53.180 ;
        RECT 107.555 53.160 107.875 53.180 ;
        RECT 100.715 46.820 101.425 46.930 ;
        RECT 104.005 46.900 104.345 46.950 ;
        RECT 104.895 47.720 106.275 51.960 ;
        RECT 100.715 46.510 101.375 46.820 ;
        RECT 100.715 46.340 100.985 46.510 ;
        RECT 104.005 44.940 104.285 46.900 ;
        RECT 104.895 46.860 105.195 47.720 ;
        RECT 105.975 46.860 106.275 47.720 ;
        RECT 106.825 46.860 107.155 51.930 ;
        RECT 106.225 46.320 106.705 46.700 ;
        RECT 106.325 45.700 106.575 46.320 ;
        RECT 106.225 45.100 106.605 45.700 ;
        RECT 95.595 43.150 95.895 44.880 ;
        RECT 103.485 44.170 104.585 44.940 ;
        RECT 106.875 44.870 107.155 46.860 ;
        RECT 109.255 47.710 109.755 68.510 ;
        RECT 110.095 49.030 110.485 70.540 ;
        RECT 110.885 69.950 111.775 70.680 ;
        RECT 110.985 65.130 111.245 69.950 ;
        RECT 112.625 68.560 115.335 69.410 ;
        RECT 112.825 65.780 114.755 68.560 ;
        RECT 120.485 68.510 121.025 71.740 ;
        RECT 121.325 70.540 121.735 73.110 ;
        RECT 132.925 70.810 133.225 70.900 ;
        RECT 117.725 67.070 118.845 67.750 ;
        RECT 118.005 65.790 118.675 67.070 ;
        RECT 111.385 65.400 116.435 65.780 ;
        RECT 117.795 65.380 118.845 65.790 ;
        RECT 110.985 63.580 111.365 65.130 ;
        RECT 111.105 55.740 111.365 63.580 ;
        RECT 116.415 63.140 116.685 65.180 ;
        RECT 117.545 63.140 117.815 65.140 ;
        RECT 116.415 56.450 117.815 63.140 ;
        RECT 111.015 55.230 111.375 55.740 ;
        RECT 110.995 54.800 111.375 55.230 ;
        RECT 116.415 55.130 116.685 56.450 ;
        RECT 117.545 55.090 117.815 56.450 ;
        RECT 118.815 55.200 119.135 65.130 ;
        RECT 118.815 55.140 119.145 55.200 ;
        RECT 110.995 54.520 111.245 54.800 ;
        RECT 110.795 54.120 115.435 54.520 ;
        RECT 116.335 54.230 117.465 54.240 ;
        RECT 118.825 54.230 119.145 55.140 ;
        RECT 110.995 52.000 111.245 54.120 ;
        RECT 115.695 53.430 116.055 54.050 ;
        RECT 115.775 52.550 116.035 53.430 ;
        RECT 116.315 53.180 119.145 54.230 ;
        RECT 115.605 52.170 116.135 52.550 ;
        RECT 110.995 51.910 111.495 52.000 ;
        RECT 110.985 51.180 111.495 51.910 ;
        RECT 111.225 50.180 111.495 51.180 ;
        RECT 112.135 50.930 112.405 51.880 ;
        RECT 112.135 50.780 112.605 50.930 ;
        RECT 112.135 50.100 112.695 50.780 ;
        RECT 112.215 50.090 112.695 50.100 ;
        RECT 111.505 49.560 112.125 49.920 ;
        RECT 111.545 49.030 111.975 49.560 ;
        RECT 110.095 48.610 111.975 49.030 ;
        RECT 112.465 48.900 112.695 50.090 ;
        RECT 111.545 47.740 111.975 48.610 ;
        RECT 112.385 48.300 112.765 48.900 ;
        RECT 109.255 47.000 109.945 47.710 ;
        RECT 111.365 47.380 111.985 47.740 ;
        RECT 111.065 47.000 111.355 47.190 ;
        RECT 109.255 46.560 111.355 47.000 ;
        RECT 109.255 46.540 109.945 46.560 ;
        RECT 111.065 46.320 111.355 46.560 ;
        RECT 111.985 46.930 112.255 47.180 ;
        RECT 112.465 46.930 112.695 48.300 ;
        RECT 115.285 46.950 115.615 51.970 ;
        RECT 116.335 51.960 117.465 53.180 ;
        RECT 118.825 53.160 119.145 53.180 ;
        RECT 111.985 46.820 112.695 46.930 ;
        RECT 115.275 46.900 115.615 46.950 ;
        RECT 116.165 47.720 117.545 51.960 ;
        RECT 111.985 46.510 112.645 46.820 ;
        RECT 111.985 46.340 112.255 46.510 ;
        RECT 115.275 44.940 115.555 46.900 ;
        RECT 116.165 46.860 116.465 47.720 ;
        RECT 117.245 46.860 117.545 47.720 ;
        RECT 118.095 46.860 118.425 51.930 ;
        RECT 117.495 46.320 117.975 46.700 ;
        RECT 117.595 45.700 117.845 46.320 ;
        RECT 117.495 45.100 117.875 45.700 ;
        RECT 20.795 39.650 21.175 40.250 ;
        RECT 20.825 39.030 21.075 39.650 ;
        RECT 20.695 38.650 21.175 39.030 ;
        RECT 20.245 33.420 20.575 38.490 ;
        RECT 21.125 37.630 21.425 38.490 ;
        RECT 22.205 37.630 22.505 38.490 ;
        RECT 23.115 38.450 23.395 40.410 ;
        RECT 26.415 38.840 26.685 39.010 ;
        RECT 26.025 38.530 26.685 38.840 ;
        RECT 21.125 33.390 22.505 37.630 ;
        RECT 23.055 38.400 23.395 38.450 ;
        RECT 25.975 38.420 26.685 38.530 ;
        RECT 19.525 32.170 19.845 32.190 ;
        RECT 21.205 32.170 22.335 33.390 ;
        RECT 23.055 33.380 23.385 38.400 ;
        RECT 25.975 37.050 26.205 38.420 ;
        RECT 26.415 38.170 26.685 38.420 ;
        RECT 27.315 38.790 27.605 39.030 ;
        RECT 28.725 38.790 29.415 38.810 ;
        RECT 27.315 38.350 29.415 38.790 ;
        RECT 27.315 38.160 27.605 38.350 ;
        RECT 26.685 37.610 27.305 37.970 ;
        RECT 28.725 37.640 29.415 38.350 ;
        RECT 25.905 36.450 26.285 37.050 ;
        RECT 26.695 36.740 27.125 37.610 ;
        RECT 25.975 35.260 26.205 36.450 ;
        RECT 26.695 36.320 28.575 36.740 ;
        RECT 26.695 35.790 27.125 36.320 ;
        RECT 26.545 35.430 27.165 35.790 ;
        RECT 25.975 35.250 26.455 35.260 ;
        RECT 25.975 34.570 26.535 35.250 ;
        RECT 26.065 34.420 26.535 34.570 ;
        RECT 26.265 33.470 26.535 34.420 ;
        RECT 27.175 34.170 27.445 35.170 ;
        RECT 27.175 33.440 27.685 34.170 ;
        RECT 27.175 33.350 27.675 33.440 ;
        RECT 22.535 32.800 23.065 33.180 ;
        RECT 19.525 31.120 22.355 32.170 ;
        RECT 22.635 31.920 22.895 32.800 ;
        RECT 22.615 31.300 22.975 31.920 ;
        RECT 27.425 31.230 27.675 33.350 ;
        RECT 19.525 30.210 19.845 31.120 ;
        RECT 21.205 31.110 22.335 31.120 ;
        RECT 23.235 30.830 27.875 31.230 ;
        RECT 27.425 30.550 27.675 30.830 ;
        RECT 19.525 30.150 19.855 30.210 ;
        RECT 19.535 20.220 19.855 30.150 ;
        RECT 20.855 28.900 21.125 30.260 ;
        RECT 21.985 28.900 22.255 30.220 ;
        RECT 27.295 30.120 27.675 30.550 ;
        RECT 27.295 29.610 27.655 30.120 ;
        RECT 20.855 22.210 22.255 28.900 ;
        RECT 20.855 20.210 21.125 22.210 ;
        RECT 21.985 20.170 22.255 22.210 ;
        RECT 27.305 21.770 27.565 29.610 ;
        RECT 27.305 20.220 27.685 21.770 ;
        RECT 19.825 19.560 20.875 19.970 ;
        RECT 22.235 19.570 27.285 19.950 ;
        RECT 19.995 18.280 20.665 19.560 ;
        RECT 19.825 17.600 20.945 18.280 ;
        RECT 23.915 16.790 25.845 19.570 ;
        RECT 23.335 15.940 26.045 16.790 ;
        RECT 27.425 15.400 27.685 20.220 ;
        RECT 26.895 14.670 27.785 15.400 ;
        RECT 28.185 14.810 28.575 36.320 ;
        RECT 28.915 16.840 29.415 37.640 ;
        RECT 31.525 38.490 31.805 40.480 ;
        RECT 34.095 40.410 35.195 41.180 ;
        RECT 42.795 40.460 43.095 42.190 ;
        RECT 32.075 39.650 32.455 40.250 ;
        RECT 32.105 39.030 32.355 39.650 ;
        RECT 31.975 38.650 32.455 39.030 ;
        RECT 31.525 33.420 31.855 38.490 ;
        RECT 32.405 37.630 32.705 38.490 ;
        RECT 33.485 37.630 33.785 38.490 ;
        RECT 34.395 38.450 34.675 40.410 ;
        RECT 37.695 38.840 37.965 39.010 ;
        RECT 37.305 38.530 37.965 38.840 ;
        RECT 32.405 33.390 33.785 37.630 ;
        RECT 34.335 38.400 34.675 38.450 ;
        RECT 37.255 38.420 37.965 38.530 ;
        RECT 30.805 32.170 31.125 32.190 ;
        RECT 32.485 32.170 33.615 33.390 ;
        RECT 34.335 33.380 34.665 38.400 ;
        RECT 37.255 37.050 37.485 38.420 ;
        RECT 37.695 38.170 37.965 38.420 ;
        RECT 38.595 38.790 38.885 39.030 ;
        RECT 40.005 38.790 40.695 38.810 ;
        RECT 38.595 38.350 40.695 38.790 ;
        RECT 38.595 38.160 38.885 38.350 ;
        RECT 37.965 37.610 38.585 37.970 ;
        RECT 40.005 37.640 40.695 38.350 ;
        RECT 37.185 36.450 37.565 37.050 ;
        RECT 37.975 36.740 38.405 37.610 ;
        RECT 37.255 35.260 37.485 36.450 ;
        RECT 37.975 36.320 39.855 36.740 ;
        RECT 37.975 35.790 38.405 36.320 ;
        RECT 37.825 35.430 38.445 35.790 ;
        RECT 37.255 35.250 37.735 35.260 ;
        RECT 37.255 34.570 37.815 35.250 ;
        RECT 37.345 34.420 37.815 34.570 ;
        RECT 37.545 33.470 37.815 34.420 ;
        RECT 38.455 34.170 38.725 35.170 ;
        RECT 38.455 33.440 38.965 34.170 ;
        RECT 38.455 33.350 38.955 33.440 ;
        RECT 33.815 32.800 34.345 33.180 ;
        RECT 30.805 31.120 33.635 32.170 ;
        RECT 33.915 31.920 34.175 32.800 ;
        RECT 33.895 31.300 34.255 31.920 ;
        RECT 38.705 31.230 38.955 33.350 ;
        RECT 30.805 30.210 31.125 31.120 ;
        RECT 32.485 31.110 33.615 31.120 ;
        RECT 34.515 30.830 39.155 31.230 ;
        RECT 38.705 30.550 38.955 30.830 ;
        RECT 30.805 30.150 31.135 30.210 ;
        RECT 30.815 20.220 31.135 30.150 ;
        RECT 32.135 28.900 32.405 30.260 ;
        RECT 33.265 28.900 33.535 30.220 ;
        RECT 38.575 30.120 38.955 30.550 ;
        RECT 38.575 29.610 38.935 30.120 ;
        RECT 32.135 22.210 33.535 28.900 ;
        RECT 32.135 20.210 32.405 22.210 ;
        RECT 33.265 20.170 33.535 22.210 ;
        RECT 38.585 21.770 38.845 29.610 ;
        RECT 38.585 20.220 38.965 21.770 ;
        RECT 31.105 19.560 32.155 19.970 ;
        RECT 33.515 19.570 38.565 19.950 ;
        RECT 31.275 18.280 31.945 19.560 ;
        RECT 31.105 17.600 32.225 18.280 ;
        RECT 28.185 12.290 28.595 14.810 ;
        RECT 28.895 13.610 29.435 16.840 ;
        RECT 35.195 16.790 37.125 19.570 ;
        RECT 34.615 15.940 37.325 16.790 ;
        RECT 38.705 15.400 38.965 20.220 ;
        RECT 38.175 14.670 39.065 15.400 ;
        RECT 39.465 14.810 39.855 36.320 ;
        RECT 40.195 16.840 40.695 37.640 ;
        RECT 42.815 38.470 43.095 40.460 ;
        RECT 45.385 40.390 46.485 41.160 ;
        RECT 54.015 40.460 54.315 42.190 ;
        RECT 43.365 39.630 43.745 40.230 ;
        RECT 43.395 39.010 43.645 39.630 ;
        RECT 43.265 38.630 43.745 39.010 ;
        RECT 42.815 33.400 43.145 38.470 ;
        RECT 43.695 37.610 43.995 38.470 ;
        RECT 44.775 37.610 45.075 38.470 ;
        RECT 45.685 38.430 45.965 40.390 ;
        RECT 48.985 38.820 49.255 38.990 ;
        RECT 48.595 38.510 49.255 38.820 ;
        RECT 43.695 33.370 45.075 37.610 ;
        RECT 45.625 38.380 45.965 38.430 ;
        RECT 48.545 38.400 49.255 38.510 ;
        RECT 42.095 32.150 42.415 32.170 ;
        RECT 43.775 32.150 44.905 33.370 ;
        RECT 45.625 33.360 45.955 38.380 ;
        RECT 48.545 37.030 48.775 38.400 ;
        RECT 48.985 38.150 49.255 38.400 ;
        RECT 49.885 38.770 50.175 39.010 ;
        RECT 51.295 38.770 51.985 38.790 ;
        RECT 49.885 38.330 51.985 38.770 ;
        RECT 49.885 38.140 50.175 38.330 ;
        RECT 49.255 37.590 49.875 37.950 ;
        RECT 51.295 37.620 51.985 38.330 ;
        RECT 48.475 36.430 48.855 37.030 ;
        RECT 49.265 36.720 49.695 37.590 ;
        RECT 48.545 35.240 48.775 36.430 ;
        RECT 49.265 36.300 51.145 36.720 ;
        RECT 49.265 35.770 49.695 36.300 ;
        RECT 49.115 35.410 49.735 35.770 ;
        RECT 48.545 35.230 49.025 35.240 ;
        RECT 48.545 34.550 49.105 35.230 ;
        RECT 48.635 34.400 49.105 34.550 ;
        RECT 48.835 33.450 49.105 34.400 ;
        RECT 49.745 34.150 50.015 35.150 ;
        RECT 49.745 33.420 50.255 34.150 ;
        RECT 49.745 33.330 50.245 33.420 ;
        RECT 45.105 32.780 45.635 33.160 ;
        RECT 42.095 31.100 44.925 32.150 ;
        RECT 45.205 31.900 45.465 32.780 ;
        RECT 45.185 31.280 45.545 31.900 ;
        RECT 49.995 31.210 50.245 33.330 ;
        RECT 42.095 30.190 42.415 31.100 ;
        RECT 43.775 31.090 44.905 31.100 ;
        RECT 45.805 30.810 50.445 31.210 ;
        RECT 49.995 30.530 50.245 30.810 ;
        RECT 42.095 30.130 42.425 30.190 ;
        RECT 42.105 20.200 42.425 30.130 ;
        RECT 43.425 28.880 43.695 30.240 ;
        RECT 44.555 28.880 44.825 30.200 ;
        RECT 49.865 30.100 50.245 30.530 ;
        RECT 49.865 29.590 50.225 30.100 ;
        RECT 43.425 22.190 44.825 28.880 ;
        RECT 43.425 20.190 43.695 22.190 ;
        RECT 44.555 20.150 44.825 22.190 ;
        RECT 49.875 21.750 50.135 29.590 ;
        RECT 49.875 20.200 50.255 21.750 ;
        RECT 42.395 19.540 43.445 19.950 ;
        RECT 44.805 19.550 49.855 19.930 ;
        RECT 42.565 18.260 43.235 19.540 ;
        RECT 42.395 17.580 43.515 18.260 ;
        RECT 28.875 12.770 29.735 13.610 ;
        RECT 28.185 11.950 30.415 12.290 ;
        RECT 39.465 11.990 39.875 14.810 ;
        RECT 40.175 13.610 40.715 16.840 ;
        RECT 46.485 16.770 48.415 19.550 ;
        RECT 45.905 15.920 48.615 16.770 ;
        RECT 49.995 15.380 50.255 20.200 ;
        RECT 49.465 14.650 50.355 15.380 ;
        RECT 50.755 14.790 51.145 36.300 ;
        RECT 51.485 16.820 51.985 37.620 ;
        RECT 54.035 38.470 54.315 40.460 ;
        RECT 56.605 40.390 57.705 41.160 ;
        RECT 65.215 40.460 65.515 42.190 ;
        RECT 76.145 42.180 77.525 42.750 ;
        RECT 83.625 42.570 85.005 43.140 ;
        RECT 87.385 42.200 88.765 42.770 ;
        RECT 94.875 42.580 96.255 43.150 ;
        RECT 106.875 43.140 107.175 44.870 ;
        RECT 114.755 44.170 115.855 44.940 ;
        RECT 118.145 44.870 118.425 46.860 ;
        RECT 120.505 47.710 121.005 68.510 ;
        RECT 121.345 49.030 121.735 70.540 ;
        RECT 122.135 69.950 123.025 70.680 ;
        RECT 132.615 70.040 134.265 70.810 ;
        RECT 122.235 65.130 122.495 69.950 ;
        RECT 123.875 68.560 126.585 69.410 ;
        RECT 124.075 65.780 126.005 68.560 ;
        RECT 128.975 67.070 130.095 67.750 ;
        RECT 129.255 65.790 129.925 67.070 ;
        RECT 122.635 65.400 127.685 65.780 ;
        RECT 129.045 65.380 130.095 65.790 ;
        RECT 132.925 65.180 133.225 70.040 ;
        RECT 137.675 68.690 139.075 69.460 ;
        RECT 138.385 65.740 138.645 68.690 ;
        RECT 149.410 68.420 150.690 69.620 ;
        RECT 149.480 65.810 150.640 68.420 ;
        RECT 133.365 65.380 138.645 65.740 ;
        RECT 122.235 63.580 122.615 65.130 ;
        RECT 122.355 55.740 122.615 63.580 ;
        RECT 127.665 63.140 127.935 65.180 ;
        RECT 128.795 63.140 129.065 65.140 ;
        RECT 127.665 56.450 129.065 63.140 ;
        RECT 122.265 55.230 122.625 55.740 ;
        RECT 122.245 54.800 122.625 55.230 ;
        RECT 127.665 55.130 127.935 56.450 ;
        RECT 128.795 55.090 129.065 56.450 ;
        RECT 130.065 55.200 130.385 65.130 ;
        RECT 132.925 61.010 133.355 65.180 ;
        RECT 138.385 65.150 138.645 65.380 ;
        RECT 138.385 64.770 138.675 65.150 ;
        RECT 130.065 55.140 130.395 55.200 ;
        RECT 133.055 55.190 133.355 61.010 ;
        RECT 122.245 54.520 122.495 54.800 ;
        RECT 122.045 54.120 126.685 54.520 ;
        RECT 127.585 54.230 128.715 54.240 ;
        RECT 130.075 54.230 130.395 55.140 ;
        RECT 138.395 55.080 138.675 64.770 ;
        RECT 149.390 64.610 150.670 65.810 ;
        RECT 122.245 52.000 122.495 54.120 ;
        RECT 126.945 53.430 127.305 54.050 ;
        RECT 127.025 52.550 127.285 53.430 ;
        RECT 127.565 53.180 130.395 54.230 ;
        RECT 126.855 52.170 127.385 52.550 ;
        RECT 122.245 51.910 122.745 52.000 ;
        RECT 122.235 51.180 122.745 51.910 ;
        RECT 122.475 50.180 122.745 51.180 ;
        RECT 123.385 50.930 123.655 51.880 ;
        RECT 123.385 50.780 123.855 50.930 ;
        RECT 123.385 50.100 123.945 50.780 ;
        RECT 123.465 50.090 123.945 50.100 ;
        RECT 122.755 49.560 123.375 49.920 ;
        RECT 122.795 49.030 123.225 49.560 ;
        RECT 121.345 48.610 123.225 49.030 ;
        RECT 123.715 48.900 123.945 50.090 ;
        RECT 122.795 47.740 123.225 48.610 ;
        RECT 123.635 48.300 124.015 48.900 ;
        RECT 120.505 47.000 121.195 47.710 ;
        RECT 122.615 47.380 123.235 47.740 ;
        RECT 122.315 47.000 122.605 47.190 ;
        RECT 120.505 46.560 122.605 47.000 ;
        RECT 120.505 46.540 121.195 46.560 ;
        RECT 122.315 46.320 122.605 46.560 ;
        RECT 123.235 46.930 123.505 47.180 ;
        RECT 123.715 46.930 123.945 48.300 ;
        RECT 126.535 46.950 126.865 51.970 ;
        RECT 127.585 51.960 128.715 53.180 ;
        RECT 130.075 53.160 130.395 53.180 ;
        RECT 123.235 46.820 123.945 46.930 ;
        RECT 126.525 46.900 126.865 46.950 ;
        RECT 127.415 47.720 128.795 51.960 ;
        RECT 123.235 46.510 123.895 46.820 ;
        RECT 123.235 46.340 123.505 46.510 ;
        RECT 126.525 44.940 126.805 46.900 ;
        RECT 127.415 46.860 127.715 47.720 ;
        RECT 128.495 46.860 128.795 47.720 ;
        RECT 129.345 46.860 129.675 51.930 ;
        RECT 128.745 46.320 129.225 46.700 ;
        RECT 128.845 45.700 129.095 46.320 ;
        RECT 128.745 45.100 129.125 45.700 ;
        RECT 118.145 43.140 118.445 44.870 ;
        RECT 126.005 44.170 127.105 44.940 ;
        RECT 129.395 44.870 129.675 46.860 ;
        RECT 129.395 43.140 129.695 44.870 ;
        RECT 98.595 42.220 99.975 42.790 ;
        RECT 106.155 42.570 107.535 43.140 ;
        RECT 109.795 42.260 111.175 42.830 ;
        RECT 117.425 42.570 118.805 43.140 ;
        RECT 121.005 42.280 122.385 42.850 ;
        RECT 128.675 42.570 130.055 43.140 ;
        RECT 54.585 39.630 54.965 40.230 ;
        RECT 54.615 39.010 54.865 39.630 ;
        RECT 54.485 38.630 54.965 39.010 ;
        RECT 54.035 33.400 54.365 38.470 ;
        RECT 54.915 37.610 55.215 38.470 ;
        RECT 55.995 37.610 56.295 38.470 ;
        RECT 56.905 38.430 57.185 40.390 ;
        RECT 60.205 38.820 60.475 38.990 ;
        RECT 59.815 38.510 60.475 38.820 ;
        RECT 54.915 33.370 56.295 37.610 ;
        RECT 56.845 38.380 57.185 38.430 ;
        RECT 59.765 38.400 60.475 38.510 ;
        RECT 53.315 32.150 53.635 32.170 ;
        RECT 54.995 32.150 56.125 33.370 ;
        RECT 56.845 33.360 57.175 38.380 ;
        RECT 59.765 37.030 59.995 38.400 ;
        RECT 60.205 38.150 60.475 38.400 ;
        RECT 61.105 38.770 61.395 39.010 ;
        RECT 62.515 38.770 63.205 38.790 ;
        RECT 61.105 38.330 63.205 38.770 ;
        RECT 61.105 38.140 61.395 38.330 ;
        RECT 60.475 37.590 61.095 37.950 ;
        RECT 62.515 37.620 63.205 38.330 ;
        RECT 59.695 36.430 60.075 37.030 ;
        RECT 60.485 36.720 60.915 37.590 ;
        RECT 59.765 35.240 59.995 36.430 ;
        RECT 60.485 36.300 62.365 36.720 ;
        RECT 60.485 35.770 60.915 36.300 ;
        RECT 60.335 35.410 60.955 35.770 ;
        RECT 59.765 35.230 60.245 35.240 ;
        RECT 59.765 34.550 60.325 35.230 ;
        RECT 59.855 34.400 60.325 34.550 ;
        RECT 60.055 33.450 60.325 34.400 ;
        RECT 60.965 34.150 61.235 35.150 ;
        RECT 60.965 33.420 61.475 34.150 ;
        RECT 60.965 33.330 61.465 33.420 ;
        RECT 56.325 32.780 56.855 33.160 ;
        RECT 53.315 31.100 56.145 32.150 ;
        RECT 56.425 31.900 56.685 32.780 ;
        RECT 56.405 31.280 56.765 31.900 ;
        RECT 61.215 31.210 61.465 33.330 ;
        RECT 53.315 30.190 53.635 31.100 ;
        RECT 54.995 31.090 56.125 31.100 ;
        RECT 57.025 30.810 61.665 31.210 ;
        RECT 61.215 30.530 61.465 30.810 ;
        RECT 53.315 30.130 53.645 30.190 ;
        RECT 53.325 20.200 53.645 30.130 ;
        RECT 54.645 28.880 54.915 30.240 ;
        RECT 55.775 28.880 56.045 30.200 ;
        RECT 61.085 30.100 61.465 30.530 ;
        RECT 61.085 29.590 61.445 30.100 ;
        RECT 54.645 22.190 56.045 28.880 ;
        RECT 54.645 20.190 54.915 22.190 ;
        RECT 55.775 20.150 56.045 22.190 ;
        RECT 61.095 21.750 61.355 29.590 ;
        RECT 61.095 20.200 61.475 21.750 ;
        RECT 53.615 19.540 54.665 19.950 ;
        RECT 56.025 19.550 61.075 19.930 ;
        RECT 53.785 18.260 54.455 19.540 ;
        RECT 53.615 17.580 54.735 18.260 ;
        RECT 40.155 12.770 41.015 13.610 ;
        RECT 50.755 12.170 51.165 14.790 ;
        RECT 51.465 13.590 52.005 16.820 ;
        RECT 57.705 16.770 59.635 19.550 ;
        RECT 57.125 15.920 59.835 16.770 ;
        RECT 61.215 15.380 61.475 20.200 ;
        RECT 60.685 14.650 61.575 15.380 ;
        RECT 61.975 14.790 62.365 36.300 ;
        RECT 62.705 16.820 63.205 37.620 ;
        RECT 65.235 38.470 65.515 40.460 ;
        RECT 67.805 40.390 68.905 41.160 ;
        RECT 76.505 40.450 76.805 42.180 ;
        RECT 65.785 39.630 66.165 40.230 ;
        RECT 65.815 39.010 66.065 39.630 ;
        RECT 65.685 38.630 66.165 39.010 ;
        RECT 65.235 33.400 65.565 38.470 ;
        RECT 66.115 37.610 66.415 38.470 ;
        RECT 67.195 37.610 67.495 38.470 ;
        RECT 68.105 38.430 68.385 40.390 ;
        RECT 71.405 38.820 71.675 38.990 ;
        RECT 71.015 38.510 71.675 38.820 ;
        RECT 66.115 33.370 67.495 37.610 ;
        RECT 68.045 38.380 68.385 38.430 ;
        RECT 70.965 38.400 71.675 38.510 ;
        RECT 64.515 32.150 64.835 32.170 ;
        RECT 66.195 32.150 67.325 33.370 ;
        RECT 68.045 33.360 68.375 38.380 ;
        RECT 70.965 37.030 71.195 38.400 ;
        RECT 71.405 38.150 71.675 38.400 ;
        RECT 72.305 38.770 72.595 39.010 ;
        RECT 73.715 38.770 74.405 38.790 ;
        RECT 72.305 38.330 74.405 38.770 ;
        RECT 72.305 38.140 72.595 38.330 ;
        RECT 71.675 37.590 72.295 37.950 ;
        RECT 73.715 37.620 74.405 38.330 ;
        RECT 70.895 36.430 71.275 37.030 ;
        RECT 71.685 36.720 72.115 37.590 ;
        RECT 70.965 35.240 71.195 36.430 ;
        RECT 71.685 36.300 73.565 36.720 ;
        RECT 71.685 35.770 72.115 36.300 ;
        RECT 71.535 35.410 72.155 35.770 ;
        RECT 70.965 35.230 71.445 35.240 ;
        RECT 70.965 34.550 71.525 35.230 ;
        RECT 71.055 34.400 71.525 34.550 ;
        RECT 71.255 33.450 71.525 34.400 ;
        RECT 72.165 34.150 72.435 35.150 ;
        RECT 72.165 33.420 72.675 34.150 ;
        RECT 72.165 33.330 72.665 33.420 ;
        RECT 67.525 32.780 68.055 33.160 ;
        RECT 64.515 31.100 67.345 32.150 ;
        RECT 67.625 31.900 67.885 32.780 ;
        RECT 67.605 31.280 67.965 31.900 ;
        RECT 72.415 31.210 72.665 33.330 ;
        RECT 64.515 30.190 64.835 31.100 ;
        RECT 66.195 31.090 67.325 31.100 ;
        RECT 68.225 30.810 72.865 31.210 ;
        RECT 72.415 30.530 72.665 30.810 ;
        RECT 64.515 30.130 64.845 30.190 ;
        RECT 64.525 20.200 64.845 30.130 ;
        RECT 65.845 28.880 66.115 30.240 ;
        RECT 66.975 28.880 67.245 30.200 ;
        RECT 72.285 30.100 72.665 30.530 ;
        RECT 72.285 29.590 72.645 30.100 ;
        RECT 65.845 22.190 67.245 28.880 ;
        RECT 65.845 20.190 66.115 22.190 ;
        RECT 66.975 20.150 67.245 22.190 ;
        RECT 72.295 21.750 72.555 29.590 ;
        RECT 72.295 20.200 72.675 21.750 ;
        RECT 64.815 19.540 65.865 19.950 ;
        RECT 67.225 19.550 72.275 19.930 ;
        RECT 64.985 18.260 65.655 19.540 ;
        RECT 64.815 17.580 65.935 18.260 ;
        RECT 51.445 12.750 52.305 13.590 ;
        RECT 27.865 11.130 30.415 11.950 ;
        RECT 28.395 11.090 30.415 11.130 ;
        RECT 39.115 10.980 41.565 11.990 ;
        RECT 50.335 10.970 52.355 12.170 ;
        RECT 61.975 12.160 62.385 14.790 ;
        RECT 62.685 13.590 63.225 16.820 ;
        RECT 68.905 16.770 70.835 19.550 ;
        RECT 68.325 15.920 71.035 16.770 ;
        RECT 72.415 15.380 72.675 20.200 ;
        RECT 71.885 14.650 72.775 15.380 ;
        RECT 73.175 14.790 73.565 36.300 ;
        RECT 73.905 16.820 74.405 37.620 ;
        RECT 76.525 38.460 76.805 40.450 ;
        RECT 79.095 40.380 80.195 41.150 ;
        RECT 87.745 40.470 88.045 42.200 ;
        RECT 77.075 39.620 77.455 40.220 ;
        RECT 77.105 39.000 77.355 39.620 ;
        RECT 76.975 38.620 77.455 39.000 ;
        RECT 76.525 33.390 76.855 38.460 ;
        RECT 77.405 37.600 77.705 38.460 ;
        RECT 78.485 37.600 78.785 38.460 ;
        RECT 79.395 38.420 79.675 40.380 ;
        RECT 82.695 38.810 82.965 38.980 ;
        RECT 82.305 38.500 82.965 38.810 ;
        RECT 77.405 33.360 78.785 37.600 ;
        RECT 79.335 38.370 79.675 38.420 ;
        RECT 82.255 38.390 82.965 38.500 ;
        RECT 75.805 32.140 76.125 32.160 ;
        RECT 77.485 32.140 78.615 33.360 ;
        RECT 79.335 33.350 79.665 38.370 ;
        RECT 82.255 37.020 82.485 38.390 ;
        RECT 82.695 38.140 82.965 38.390 ;
        RECT 83.595 38.760 83.885 39.000 ;
        RECT 85.005 38.760 85.695 38.780 ;
        RECT 83.595 38.320 85.695 38.760 ;
        RECT 83.595 38.130 83.885 38.320 ;
        RECT 82.965 37.580 83.585 37.940 ;
        RECT 85.005 37.610 85.695 38.320 ;
        RECT 82.185 36.420 82.565 37.020 ;
        RECT 82.975 36.710 83.405 37.580 ;
        RECT 82.255 35.230 82.485 36.420 ;
        RECT 82.975 36.290 84.855 36.710 ;
        RECT 82.975 35.760 83.405 36.290 ;
        RECT 82.825 35.400 83.445 35.760 ;
        RECT 82.255 35.220 82.735 35.230 ;
        RECT 82.255 34.540 82.815 35.220 ;
        RECT 82.345 34.390 82.815 34.540 ;
        RECT 82.545 33.440 82.815 34.390 ;
        RECT 83.455 34.140 83.725 35.140 ;
        RECT 83.455 33.410 83.965 34.140 ;
        RECT 83.455 33.320 83.955 33.410 ;
        RECT 78.815 32.770 79.345 33.150 ;
        RECT 75.805 31.090 78.635 32.140 ;
        RECT 78.915 31.890 79.175 32.770 ;
        RECT 78.895 31.270 79.255 31.890 ;
        RECT 83.705 31.200 83.955 33.320 ;
        RECT 75.805 30.180 76.125 31.090 ;
        RECT 77.485 31.080 78.615 31.090 ;
        RECT 79.515 30.800 84.155 31.200 ;
        RECT 83.705 30.520 83.955 30.800 ;
        RECT 75.805 30.120 76.135 30.180 ;
        RECT 75.815 20.190 76.135 30.120 ;
        RECT 77.135 28.870 77.405 30.230 ;
        RECT 78.265 28.870 78.535 30.190 ;
        RECT 83.575 30.090 83.955 30.520 ;
        RECT 83.575 29.580 83.935 30.090 ;
        RECT 77.135 22.180 78.535 28.870 ;
        RECT 77.135 20.180 77.405 22.180 ;
        RECT 78.265 20.140 78.535 22.180 ;
        RECT 83.585 21.740 83.845 29.580 ;
        RECT 83.585 20.190 83.965 21.740 ;
        RECT 76.105 19.530 77.155 19.940 ;
        RECT 78.515 19.540 83.565 19.920 ;
        RECT 76.275 18.250 76.945 19.530 ;
        RECT 76.105 17.570 77.225 18.250 ;
        RECT 62.665 12.750 63.525 13.590 ;
        RECT 73.175 12.190 73.585 14.790 ;
        RECT 73.885 13.590 74.425 16.820 ;
        RECT 80.195 16.760 82.125 19.540 ;
        RECT 79.615 15.910 82.325 16.760 ;
        RECT 83.705 15.370 83.965 20.190 ;
        RECT 83.175 14.640 84.065 15.370 ;
        RECT 84.465 14.780 84.855 36.290 ;
        RECT 85.195 16.810 85.695 37.610 ;
        RECT 87.765 38.480 88.045 40.470 ;
        RECT 90.335 40.400 91.435 41.170 ;
        RECT 98.955 40.490 99.255 42.220 ;
        RECT 88.315 39.640 88.695 40.240 ;
        RECT 88.345 39.020 88.595 39.640 ;
        RECT 88.215 38.640 88.695 39.020 ;
        RECT 87.765 33.410 88.095 38.480 ;
        RECT 88.645 37.620 88.945 38.480 ;
        RECT 89.725 37.620 90.025 38.480 ;
        RECT 90.635 38.440 90.915 40.400 ;
        RECT 93.935 38.830 94.205 39.000 ;
        RECT 93.545 38.520 94.205 38.830 ;
        RECT 88.645 33.380 90.025 37.620 ;
        RECT 90.575 38.390 90.915 38.440 ;
        RECT 93.495 38.410 94.205 38.520 ;
        RECT 87.045 32.160 87.365 32.180 ;
        RECT 88.725 32.160 89.855 33.380 ;
        RECT 90.575 33.370 90.905 38.390 ;
        RECT 93.495 37.040 93.725 38.410 ;
        RECT 93.935 38.160 94.205 38.410 ;
        RECT 94.835 38.780 95.125 39.020 ;
        RECT 96.245 38.780 96.935 38.800 ;
        RECT 94.835 38.340 96.935 38.780 ;
        RECT 94.835 38.150 95.125 38.340 ;
        RECT 94.205 37.600 94.825 37.960 ;
        RECT 96.245 37.630 96.935 38.340 ;
        RECT 93.425 36.440 93.805 37.040 ;
        RECT 94.215 36.730 94.645 37.600 ;
        RECT 93.495 35.250 93.725 36.440 ;
        RECT 94.215 36.310 96.095 36.730 ;
        RECT 94.215 35.780 94.645 36.310 ;
        RECT 94.065 35.420 94.685 35.780 ;
        RECT 93.495 35.240 93.975 35.250 ;
        RECT 93.495 34.560 94.055 35.240 ;
        RECT 93.585 34.410 94.055 34.560 ;
        RECT 93.785 33.460 94.055 34.410 ;
        RECT 94.695 34.160 94.965 35.160 ;
        RECT 94.695 33.430 95.205 34.160 ;
        RECT 94.695 33.340 95.195 33.430 ;
        RECT 90.055 32.790 90.585 33.170 ;
        RECT 87.045 31.110 89.875 32.160 ;
        RECT 90.155 31.910 90.415 32.790 ;
        RECT 90.135 31.290 90.495 31.910 ;
        RECT 94.945 31.220 95.195 33.340 ;
        RECT 87.045 30.200 87.365 31.110 ;
        RECT 88.725 31.100 89.855 31.110 ;
        RECT 90.755 30.820 95.395 31.220 ;
        RECT 94.945 30.540 95.195 30.820 ;
        RECT 87.045 30.140 87.375 30.200 ;
        RECT 87.055 20.210 87.375 30.140 ;
        RECT 88.375 28.890 88.645 30.250 ;
        RECT 89.505 28.890 89.775 30.210 ;
        RECT 94.815 30.110 95.195 30.540 ;
        RECT 94.815 29.600 95.175 30.110 ;
        RECT 88.375 22.200 89.775 28.890 ;
        RECT 88.375 20.200 88.645 22.200 ;
        RECT 89.505 20.160 89.775 22.200 ;
        RECT 94.825 21.760 95.085 29.600 ;
        RECT 94.825 20.210 95.205 21.760 ;
        RECT 87.345 19.550 88.395 19.960 ;
        RECT 89.755 19.560 94.805 19.940 ;
        RECT 87.515 18.270 88.185 19.550 ;
        RECT 87.345 17.590 88.465 18.270 ;
        RECT 73.865 12.750 74.725 13.590 ;
        RECT 61.415 10.960 63.435 12.160 ;
        RECT 72.725 10.990 74.745 12.190 ;
        RECT 84.465 12.180 84.875 14.780 ;
        RECT 85.175 13.580 85.715 16.810 ;
        RECT 91.435 16.780 93.365 19.560 ;
        RECT 90.855 15.930 93.565 16.780 ;
        RECT 94.945 15.390 95.205 20.210 ;
        RECT 94.415 14.660 95.305 15.390 ;
        RECT 95.705 14.800 96.095 36.310 ;
        RECT 96.435 16.830 96.935 37.630 ;
        RECT 98.975 38.500 99.255 40.490 ;
        RECT 101.545 40.420 102.645 41.190 ;
        RECT 110.155 40.530 110.455 42.260 ;
        RECT 99.525 39.660 99.905 40.260 ;
        RECT 99.555 39.040 99.805 39.660 ;
        RECT 99.425 38.660 99.905 39.040 ;
        RECT 98.975 33.430 99.305 38.500 ;
        RECT 99.855 37.640 100.155 38.500 ;
        RECT 100.935 37.640 101.235 38.500 ;
        RECT 101.845 38.460 102.125 40.420 ;
        RECT 105.145 38.850 105.415 39.020 ;
        RECT 104.755 38.540 105.415 38.850 ;
        RECT 99.855 33.400 101.235 37.640 ;
        RECT 101.785 38.410 102.125 38.460 ;
        RECT 104.705 38.430 105.415 38.540 ;
        RECT 98.255 32.180 98.575 32.200 ;
        RECT 99.935 32.180 101.065 33.400 ;
        RECT 101.785 33.390 102.115 38.410 ;
        RECT 104.705 37.060 104.935 38.430 ;
        RECT 105.145 38.180 105.415 38.430 ;
        RECT 106.045 38.800 106.335 39.040 ;
        RECT 107.455 38.800 108.145 38.820 ;
        RECT 106.045 38.360 108.145 38.800 ;
        RECT 106.045 38.170 106.335 38.360 ;
        RECT 105.415 37.620 106.035 37.980 ;
        RECT 107.455 37.650 108.145 38.360 ;
        RECT 104.635 36.460 105.015 37.060 ;
        RECT 105.425 36.750 105.855 37.620 ;
        RECT 104.705 35.270 104.935 36.460 ;
        RECT 105.425 36.330 107.305 36.750 ;
        RECT 105.425 35.800 105.855 36.330 ;
        RECT 105.275 35.440 105.895 35.800 ;
        RECT 104.705 35.260 105.185 35.270 ;
        RECT 104.705 34.580 105.265 35.260 ;
        RECT 104.795 34.430 105.265 34.580 ;
        RECT 104.995 33.480 105.265 34.430 ;
        RECT 105.905 34.180 106.175 35.180 ;
        RECT 105.905 33.450 106.415 34.180 ;
        RECT 105.905 33.360 106.405 33.450 ;
        RECT 101.265 32.810 101.795 33.190 ;
        RECT 98.255 31.130 101.085 32.180 ;
        RECT 101.365 31.930 101.625 32.810 ;
        RECT 101.345 31.310 101.705 31.930 ;
        RECT 106.155 31.240 106.405 33.360 ;
        RECT 98.255 30.220 98.575 31.130 ;
        RECT 99.935 31.120 101.065 31.130 ;
        RECT 101.965 30.840 106.605 31.240 ;
        RECT 106.155 30.560 106.405 30.840 ;
        RECT 98.255 30.160 98.585 30.220 ;
        RECT 98.265 20.230 98.585 30.160 ;
        RECT 99.585 28.910 99.855 30.270 ;
        RECT 100.715 28.910 100.985 30.230 ;
        RECT 106.025 30.130 106.405 30.560 ;
        RECT 106.025 29.620 106.385 30.130 ;
        RECT 99.585 22.220 100.985 28.910 ;
        RECT 99.585 20.220 99.855 22.220 ;
        RECT 100.715 20.180 100.985 22.220 ;
        RECT 106.035 21.780 106.295 29.620 ;
        RECT 106.035 20.230 106.415 21.780 ;
        RECT 98.555 19.570 99.605 19.980 ;
        RECT 100.965 19.580 106.015 19.960 ;
        RECT 98.725 18.290 99.395 19.570 ;
        RECT 98.555 17.610 99.675 18.290 ;
        RECT 85.155 12.740 86.015 13.580 ;
        RECT 95.705 12.180 96.115 14.800 ;
        RECT 96.415 13.600 96.955 16.830 ;
        RECT 102.645 16.800 104.575 19.580 ;
        RECT 102.065 15.950 104.775 16.800 ;
        RECT 106.155 15.410 106.415 20.230 ;
        RECT 105.625 14.680 106.515 15.410 ;
        RECT 106.915 14.820 107.305 36.330 ;
        RECT 107.645 16.850 108.145 37.650 ;
        RECT 110.175 38.540 110.455 40.530 ;
        RECT 112.745 40.460 113.845 41.230 ;
        RECT 121.365 40.550 121.665 42.280 ;
        RECT 142.880 42.020 144.100 43.390 ;
        RECT 110.725 39.700 111.105 40.300 ;
        RECT 110.755 39.080 111.005 39.700 ;
        RECT 110.625 38.700 111.105 39.080 ;
        RECT 110.175 33.470 110.505 38.540 ;
        RECT 111.055 37.680 111.355 38.540 ;
        RECT 112.135 37.680 112.435 38.540 ;
        RECT 113.045 38.500 113.325 40.460 ;
        RECT 116.345 38.890 116.615 39.060 ;
        RECT 115.955 38.580 116.615 38.890 ;
        RECT 111.055 33.440 112.435 37.680 ;
        RECT 112.985 38.450 113.325 38.500 ;
        RECT 115.905 38.470 116.615 38.580 ;
        RECT 109.455 32.220 109.775 32.240 ;
        RECT 111.135 32.220 112.265 33.440 ;
        RECT 112.985 33.430 113.315 38.450 ;
        RECT 115.905 37.100 116.135 38.470 ;
        RECT 116.345 38.220 116.615 38.470 ;
        RECT 117.245 38.840 117.535 39.080 ;
        RECT 118.655 38.840 119.345 38.860 ;
        RECT 117.245 38.400 119.345 38.840 ;
        RECT 117.245 38.210 117.535 38.400 ;
        RECT 116.615 37.660 117.235 38.020 ;
        RECT 118.655 37.690 119.345 38.400 ;
        RECT 115.835 36.500 116.215 37.100 ;
        RECT 116.625 36.790 117.055 37.660 ;
        RECT 115.905 35.310 116.135 36.500 ;
        RECT 116.625 36.370 118.505 36.790 ;
        RECT 116.625 35.840 117.055 36.370 ;
        RECT 116.475 35.480 117.095 35.840 ;
        RECT 115.905 35.300 116.385 35.310 ;
        RECT 115.905 34.620 116.465 35.300 ;
        RECT 115.995 34.470 116.465 34.620 ;
        RECT 116.195 33.520 116.465 34.470 ;
        RECT 117.105 34.220 117.375 35.220 ;
        RECT 117.105 33.490 117.615 34.220 ;
        RECT 117.105 33.400 117.605 33.490 ;
        RECT 112.465 32.850 112.995 33.230 ;
        RECT 109.455 31.170 112.285 32.220 ;
        RECT 112.565 31.970 112.825 32.850 ;
        RECT 112.545 31.350 112.905 31.970 ;
        RECT 117.355 31.280 117.605 33.400 ;
        RECT 109.455 30.260 109.775 31.170 ;
        RECT 111.135 31.160 112.265 31.170 ;
        RECT 113.165 30.880 117.805 31.280 ;
        RECT 117.355 30.600 117.605 30.880 ;
        RECT 109.455 30.200 109.785 30.260 ;
        RECT 109.465 20.270 109.785 30.200 ;
        RECT 110.785 28.950 111.055 30.310 ;
        RECT 111.915 28.950 112.185 30.270 ;
        RECT 117.225 30.170 117.605 30.600 ;
        RECT 117.225 29.660 117.585 30.170 ;
        RECT 110.785 22.260 112.185 28.950 ;
        RECT 110.785 20.260 111.055 22.260 ;
        RECT 111.915 20.220 112.185 22.260 ;
        RECT 117.235 21.820 117.495 29.660 ;
        RECT 117.235 20.270 117.615 21.820 ;
        RECT 109.755 19.610 110.805 20.020 ;
        RECT 112.165 19.620 117.215 20.000 ;
        RECT 109.925 18.330 110.595 19.610 ;
        RECT 109.755 17.650 110.875 18.330 ;
        RECT 96.395 12.760 97.255 13.600 ;
        RECT 106.915 12.230 107.325 14.820 ;
        RECT 107.625 13.620 108.165 16.850 ;
        RECT 113.845 16.840 115.775 19.620 ;
        RECT 113.265 15.990 115.975 16.840 ;
        RECT 117.355 15.450 117.615 20.270 ;
        RECT 116.825 14.720 117.715 15.450 ;
        RECT 118.115 14.860 118.505 36.370 ;
        RECT 118.845 16.890 119.345 37.690 ;
        RECT 121.385 38.560 121.665 40.550 ;
        RECT 123.955 40.480 125.055 41.250 ;
        RECT 121.935 39.720 122.315 40.320 ;
        RECT 121.965 39.100 122.215 39.720 ;
        RECT 121.835 38.720 122.315 39.100 ;
        RECT 121.385 33.490 121.715 38.560 ;
        RECT 122.265 37.700 122.565 38.560 ;
        RECT 123.345 37.700 123.645 38.560 ;
        RECT 124.255 38.520 124.535 40.480 ;
        RECT 127.555 38.910 127.825 39.080 ;
        RECT 127.165 38.600 127.825 38.910 ;
        RECT 122.265 33.460 123.645 37.700 ;
        RECT 124.195 38.470 124.535 38.520 ;
        RECT 127.115 38.490 127.825 38.600 ;
        RECT 120.665 32.240 120.985 32.260 ;
        RECT 122.345 32.240 123.475 33.460 ;
        RECT 124.195 33.450 124.525 38.470 ;
        RECT 127.115 37.120 127.345 38.490 ;
        RECT 127.555 38.240 127.825 38.490 ;
        RECT 128.455 38.860 128.745 39.100 ;
        RECT 142.940 38.950 144.100 42.020 ;
        RECT 129.865 38.860 130.555 38.880 ;
        RECT 128.455 38.420 130.555 38.860 ;
        RECT 128.455 38.230 128.745 38.420 ;
        RECT 127.825 37.680 128.445 38.040 ;
        RECT 129.865 37.710 130.555 38.420 ;
        RECT 127.045 36.520 127.425 37.120 ;
        RECT 127.835 36.810 128.265 37.680 ;
        RECT 127.115 35.330 127.345 36.520 ;
        RECT 127.835 36.390 129.715 36.810 ;
        RECT 127.835 35.860 128.265 36.390 ;
        RECT 127.685 35.500 128.305 35.860 ;
        RECT 127.115 35.320 127.595 35.330 ;
        RECT 127.115 34.640 127.675 35.320 ;
        RECT 127.205 34.490 127.675 34.640 ;
        RECT 127.405 33.540 127.675 34.490 ;
        RECT 128.315 34.240 128.585 35.240 ;
        RECT 128.315 33.510 128.825 34.240 ;
        RECT 128.315 33.420 128.815 33.510 ;
        RECT 123.675 32.870 124.205 33.250 ;
        RECT 120.665 31.190 123.495 32.240 ;
        RECT 123.775 31.990 124.035 32.870 ;
        RECT 123.755 31.370 124.115 31.990 ;
        RECT 128.565 31.300 128.815 33.420 ;
        RECT 120.665 30.280 120.985 31.190 ;
        RECT 122.345 31.180 123.475 31.190 ;
        RECT 124.375 30.900 129.015 31.300 ;
        RECT 128.565 30.620 128.815 30.900 ;
        RECT 120.665 30.220 120.995 30.280 ;
        RECT 120.675 20.290 120.995 30.220 ;
        RECT 121.995 28.970 122.265 30.330 ;
        RECT 123.125 28.970 123.395 30.290 ;
        RECT 128.435 30.190 128.815 30.620 ;
        RECT 128.435 29.680 128.795 30.190 ;
        RECT 121.995 22.280 123.395 28.970 ;
        RECT 121.995 20.280 122.265 22.280 ;
        RECT 123.125 20.240 123.395 22.280 ;
        RECT 128.445 21.840 128.705 29.680 ;
        RECT 128.445 20.290 128.825 21.840 ;
        RECT 120.965 19.630 122.015 20.040 ;
        RECT 123.375 19.640 128.425 20.020 ;
        RECT 121.135 18.350 121.805 19.630 ;
        RECT 120.965 17.670 122.085 18.350 ;
        RECT 107.605 12.780 108.465 13.620 ;
        RECT 118.115 12.230 118.525 14.860 ;
        RECT 118.825 13.660 119.365 16.890 ;
        RECT 125.055 16.860 126.985 19.640 ;
        RECT 124.475 16.010 127.185 16.860 ;
        RECT 128.565 15.470 128.825 20.290 ;
        RECT 128.035 14.740 128.925 15.470 ;
        RECT 129.325 14.880 129.715 36.390 ;
        RECT 130.055 16.910 130.555 37.710 ;
        RECT 142.900 37.580 144.120 38.950 ;
        RECT 132.395 24.340 132.705 30.230 ;
        RECT 132.195 20.120 132.705 24.340 ;
        RECT 118.805 12.820 119.665 13.660 ;
        RECT 129.325 12.260 129.735 14.880 ;
        RECT 130.035 13.680 130.575 16.910 ;
        RECT 132.195 15.510 132.505 20.120 ;
        RECT 137.715 19.980 138.005 30.170 ;
        RECT 132.685 19.590 138.005 19.980 ;
        RECT 137.715 16.940 138.005 19.590 ;
        RECT 142.940 17.940 144.090 19.160 ;
        RECT 145.080 18.760 146.200 18.930 ;
        RECT 137.395 15.890 138.295 16.940 ;
        RECT 137.715 15.720 138.005 15.890 ;
        RECT 131.975 14.270 132.735 15.510 ;
        RECT 142.940 15.090 144.050 17.940 ;
        RECT 142.900 13.870 144.050 15.090 ;
        RECT 145.070 14.920 146.200 18.760 ;
        RECT 145.030 13.970 146.200 14.920 ;
        RECT 145.030 13.900 146.150 13.970 ;
        RECT 130.015 12.840 130.875 13.680 ;
        RECT 83.845 10.980 85.865 12.180 ;
        RECT 95.145 10.980 97.165 12.180 ;
        RECT 106.335 11.030 108.355 12.230 ;
        RECT 117.565 11.030 119.585 12.230 ;
        RECT 128.865 11.060 130.885 12.260 ;
        RECT 74.340 0.110 75.630 1.460 ;
        RECT 93.550 0.180 94.840 1.530 ;
        RECT 112.950 0.310 114.240 1.660 ;
        RECT 131.850 0.380 133.490 1.930 ;
        RECT 151.650 0.250 152.920 1.470 ;
      LAYER met3 ;
        RECT 135.340 223.855 136.790 225.205 ;
        RECT 138.130 223.785 139.580 225.135 ;
        RECT 143.180 223.815 144.630 225.165 ;
        RECT 34.860 206.110 36.840 206.440 ;
        RECT 64.860 206.110 66.840 206.440 ;
        RECT 94.860 206.110 96.840 206.440 ;
        RECT 19.860 203.390 21.840 203.720 ;
        RECT 49.860 203.390 51.840 203.720 ;
        RECT 79.860 203.390 81.840 203.720 ;
        RECT 109.860 203.390 111.840 203.720 ;
        RECT 34.860 200.670 36.840 201.000 ;
        RECT 64.860 200.670 66.840 201.000 ;
        RECT 94.860 200.670 96.840 201.000 ;
        RECT 19.860 197.950 21.840 198.280 ;
        RECT 49.860 197.950 51.840 198.280 ;
        RECT 79.860 197.950 81.840 198.280 ;
        RECT 109.860 197.950 111.840 198.280 ;
        RECT 63.475 196.565 63.805 196.580 ;
        RECT 66.235 196.565 66.565 196.580 ;
        RECT 63.475 196.265 66.565 196.565 ;
        RECT 63.475 196.250 63.805 196.265 ;
        RECT 66.235 196.250 66.565 196.265 ;
        RECT 34.860 195.230 36.840 195.560 ;
        RECT 64.860 195.230 66.840 195.560 ;
        RECT 94.860 195.230 96.840 195.560 ;
        RECT 19.860 192.510 21.840 192.840 ;
        RECT 49.860 192.510 51.840 192.840 ;
        RECT 79.860 192.510 81.840 192.840 ;
        RECT 109.860 192.510 111.840 192.840 ;
        RECT 34.860 189.790 36.840 190.120 ;
        RECT 64.860 189.790 66.840 190.120 ;
        RECT 94.860 189.790 96.840 190.120 ;
        RECT 19.860 187.070 21.840 187.400 ;
        RECT 49.860 187.070 51.840 187.400 ;
        RECT 79.860 187.070 81.840 187.400 ;
        RECT 109.860 187.070 111.840 187.400 ;
        RECT 34.860 184.350 36.840 184.680 ;
        RECT 64.860 184.350 66.840 184.680 ;
        RECT 94.860 184.350 96.840 184.680 ;
        RECT 62.095 182.965 62.425 182.980 ;
        RECT 63.680 182.965 64.060 182.975 ;
        RECT 62.095 182.665 64.060 182.965 ;
        RECT 62.095 182.650 62.425 182.665 ;
        RECT 63.680 182.655 64.060 182.665 ;
        RECT 19.860 181.630 21.840 181.960 ;
        RECT 49.860 181.630 51.840 181.960 ;
        RECT 79.860 181.630 81.840 181.960 ;
        RECT 109.860 181.630 111.840 181.960 ;
        RECT 34.860 178.910 36.840 179.240 ;
        RECT 64.860 178.910 66.840 179.240 ;
        RECT 94.860 178.910 96.840 179.240 ;
        RECT 39.095 176.855 39.425 176.860 ;
        RECT 38.840 176.845 39.425 176.855 ;
        RECT 38.840 176.545 39.650 176.845 ;
        RECT 38.840 176.535 39.425 176.545 ;
        RECT 39.095 176.530 39.425 176.535 ;
        RECT 19.860 176.190 21.840 176.520 ;
        RECT 49.860 176.190 51.840 176.520 ;
        RECT 79.860 176.190 81.840 176.520 ;
        RECT 109.860 176.190 111.840 176.520 ;
        RECT 68.535 175.485 68.865 175.500 ;
        RECT 72.675 175.485 73.005 175.500 ;
        RECT 68.535 175.185 73.005 175.485 ;
        RECT 68.535 175.170 68.865 175.185 ;
        RECT 72.675 175.170 73.005 175.185 ;
        RECT 99.815 174.805 100.145 174.820 ;
        RECT 105.795 174.805 106.125 174.820 ;
        RECT 110.395 174.805 110.725 174.820 ;
        RECT 99.815 174.505 110.725 174.805 ;
        RECT 99.815 174.490 100.145 174.505 ;
        RECT 105.795 174.490 106.125 174.505 ;
        RECT 110.395 174.490 110.725 174.505 ;
        RECT 34.860 173.470 36.840 173.800 ;
        RECT 64.860 173.470 66.840 173.800 ;
        RECT 94.860 173.470 96.840 173.800 ;
        RECT 78.195 172.765 78.525 172.780 ;
        RECT 97.975 172.765 98.305 172.780 ;
        RECT 59.120 172.465 98.305 172.765 ;
        RECT 133.700 172.500 134.930 172.705 ;
        RECT 30.355 172.085 30.685 172.100 ;
        RECT 50.135 172.085 50.465 172.100 ;
        RECT 57.240 172.085 57.620 172.095 ;
        RECT 59.120 172.085 59.420 172.465 ;
        RECT 78.195 172.450 78.525 172.465 ;
        RECT 97.975 172.450 98.305 172.465 ;
        RECT 30.355 171.785 59.420 172.085 ;
        RECT 30.355 171.770 30.685 171.785 ;
        RECT 50.135 171.770 50.465 171.785 ;
        RECT 57.240 171.775 57.620 171.785 ;
        RECT 19.860 170.750 21.840 171.080 ;
        RECT 49.860 170.750 51.840 171.080 ;
        RECT 79.860 170.750 81.840 171.080 ;
        RECT 109.860 170.750 111.840 171.080 ;
        RECT 129.030 170.130 134.930 172.500 ;
        RECT 133.700 170.095 134.930 170.130 ;
        RECT 115.915 169.365 116.245 169.380 ;
        RECT 119.370 169.365 121.370 169.515 ;
        RECT 115.915 169.065 121.370 169.365 ;
        RECT 115.915 169.050 116.245 169.065 ;
        RECT 119.370 168.915 121.370 169.065 ;
        RECT 34.860 168.030 36.840 168.360 ;
        RECT 64.860 168.030 66.840 168.360 ;
        RECT 94.860 168.030 96.840 168.360 ;
        RECT 19.860 165.310 21.840 165.640 ;
        RECT 49.860 165.310 51.840 165.640 ;
        RECT 79.860 165.310 81.840 165.640 ;
        RECT 109.860 165.310 111.840 165.640 ;
        RECT 34.955 163.925 35.285 163.940 ;
        RECT 34.955 163.625 38.260 163.925 ;
        RECT 34.955 163.610 35.285 163.625 ;
        RECT 34.860 162.590 36.840 162.920 ;
        RECT 37.960 161.220 38.260 163.625 ;
        RECT 64.860 162.590 66.840 162.920 ;
        RECT 94.860 162.590 96.840 162.920 ;
        RECT 37.960 160.905 38.505 161.220 ;
        RECT 38.175 160.890 38.505 160.905 ;
        RECT 19.860 159.870 21.840 160.200 ;
        RECT 49.860 159.870 51.840 160.200 ;
        RECT 79.860 159.870 81.840 160.200 ;
        RECT 109.860 159.870 111.840 160.200 ;
        RECT 40.015 159.165 40.345 159.180 ;
        RECT 46.915 159.165 47.245 159.180 ;
        RECT 40.015 158.865 47.245 159.165 ;
        RECT 40.015 158.850 40.345 158.865 ;
        RECT 46.915 158.850 47.245 158.865 ;
        RECT 62.095 159.165 62.425 159.180 ;
        RECT 71.755 159.165 72.085 159.180 ;
        RECT 62.095 158.865 72.085 159.165 ;
        RECT 62.095 158.850 62.425 158.865 ;
        RECT 71.755 158.850 72.085 158.865 ;
        RECT 35.875 158.485 36.205 158.500 ;
        RECT 41.855 158.485 42.185 158.500 ;
        RECT 35.875 158.185 42.185 158.485 ;
        RECT 35.875 158.170 36.205 158.185 ;
        RECT 41.855 158.170 42.185 158.185 ;
        RECT 34.860 157.150 36.840 157.480 ;
        RECT 64.860 157.150 66.840 157.480 ;
        RECT 94.860 157.150 96.840 157.480 ;
        RECT 29.895 156.445 30.225 156.460 ;
        RECT 35.415 156.445 35.745 156.460 ;
        RECT 39.095 156.445 39.425 156.460 ;
        RECT 29.895 156.145 34.580 156.445 ;
        RECT 29.895 156.130 30.225 156.145 ;
        RECT 34.280 155.765 34.580 156.145 ;
        RECT 35.415 156.145 39.425 156.445 ;
        RECT 35.415 156.130 35.745 156.145 ;
        RECT 39.095 156.130 39.425 156.145 ;
        RECT 38.175 155.765 38.505 155.780 ;
        RECT 34.280 155.465 38.505 155.765 ;
        RECT 38.175 155.450 38.505 155.465 ;
        RECT 19.860 154.430 21.840 154.760 ;
        RECT 49.860 154.430 51.840 154.760 ;
        RECT 79.860 154.430 81.840 154.760 ;
        RECT 109.860 154.430 111.840 154.760 ;
        RECT 34.860 151.710 36.840 152.040 ;
        RECT 64.860 151.710 66.840 152.040 ;
        RECT 94.860 151.710 96.840 152.040 ;
        RECT 33.115 151.685 33.445 151.700 ;
        RECT 33.115 151.370 33.660 151.685 ;
        RECT 30.815 151.005 31.145 151.020 ;
        RECT 33.360 151.005 33.660 151.370 ;
        RECT 36.795 151.005 37.125 151.020 ;
        RECT 60.255 151.005 60.585 151.020 ;
        RECT 30.815 150.705 60.585 151.005 ;
        RECT 30.815 150.690 31.145 150.705 ;
        RECT 36.795 150.690 37.125 150.705 ;
        RECT 60.255 150.690 60.585 150.705 ;
        RECT 63.475 150.325 63.805 150.340 ;
        RECT 100.480 150.325 100.860 150.335 ;
        RECT 63.475 150.025 100.860 150.325 ;
        RECT 63.475 150.010 63.805 150.025 ;
        RECT 100.480 150.015 100.860 150.025 ;
        RECT 57.035 149.655 57.365 149.660 ;
        RECT 68.535 149.655 68.865 149.660 ;
        RECT 57.035 149.645 57.620 149.655 ;
        RECT 56.810 149.345 57.620 149.645 ;
        RECT 57.035 149.335 57.620 149.345 ;
        RECT 68.280 149.645 68.865 149.655 ;
        RECT 68.280 149.345 69.090 149.645 ;
        RECT 68.280 149.335 68.865 149.345 ;
        RECT 57.035 149.330 57.365 149.335 ;
        RECT 68.535 149.330 68.865 149.335 ;
        RECT 19.860 148.990 21.840 149.320 ;
        RECT 49.860 148.990 51.840 149.320 ;
        RECT 79.860 148.990 81.840 149.320 ;
        RECT 109.860 148.990 111.840 149.320 ;
        RECT 50.595 147.605 50.925 147.620 ;
        RECT 68.535 147.605 68.865 147.620 ;
        RECT 50.595 147.305 68.865 147.605 ;
        RECT 50.595 147.290 50.925 147.305 ;
        RECT 68.535 147.290 68.865 147.305 ;
        RECT 97.975 147.605 98.305 147.620 ;
        RECT 100.275 147.605 100.605 147.620 ;
        RECT 97.975 147.305 100.605 147.605 ;
        RECT 97.975 147.290 98.305 147.305 ;
        RECT 100.275 147.290 100.605 147.305 ;
        RECT 34.860 146.270 36.840 146.600 ;
        RECT 64.860 146.270 66.840 146.600 ;
        RECT 94.860 146.270 96.840 146.600 ;
        RECT 19.860 143.550 21.840 143.880 ;
        RECT 49.860 143.550 51.840 143.880 ;
        RECT 79.860 143.550 81.840 143.880 ;
        RECT 109.860 143.550 111.840 143.880 ;
        RECT 34.860 140.830 36.840 141.160 ;
        RECT 64.860 140.830 66.840 141.160 ;
        RECT 94.860 140.830 96.840 141.160 ;
        RECT 38.635 140.815 38.965 140.820 ;
        RECT 38.635 140.805 39.220 140.815 ;
        RECT 100.735 140.805 101.065 140.820 ;
        RECT 38.635 140.505 39.420 140.805 ;
        RECT 38.635 140.495 39.220 140.505 ;
        RECT 38.635 140.490 38.965 140.495 ;
        RECT 100.520 140.490 101.065 140.805 ;
        RECT 100.520 140.125 100.820 140.490 ;
        RECT 101.655 140.125 101.985 140.140 ;
        RECT 99.600 139.825 101.985 140.125 ;
        RECT 78.195 139.445 78.525 139.460 ;
        RECT 91.075 139.445 91.405 139.460 ;
        RECT 99.600 139.445 99.900 139.825 ;
        RECT 101.655 139.810 101.985 139.825 ;
        RECT 78.195 139.145 99.900 139.445 ;
        RECT 100.480 139.445 100.860 139.455 ;
        RECT 100.480 139.145 112.780 139.445 ;
        RECT 78.195 139.130 78.525 139.145 ;
        RECT 91.075 139.130 91.405 139.145 ;
        RECT 100.480 139.135 100.860 139.145 ;
        RECT 19.860 138.110 21.840 138.440 ;
        RECT 49.860 138.110 51.840 138.440 ;
        RECT 79.860 138.110 81.840 138.440 ;
        RECT 109.860 138.110 111.840 138.440 ;
        RECT 112.480 138.085 112.780 139.145 ;
        RECT 119.370 138.085 121.370 138.235 ;
        RECT 132.510 138.165 135.210 140.035 ;
        RECT 112.480 137.785 121.370 138.085 ;
        RECT 119.370 137.635 121.370 137.785 ;
        RECT 49.215 136.725 49.545 136.740 ;
        RECT 51.515 136.725 51.845 136.740 ;
        RECT 55.195 136.725 55.525 136.740 ;
        RECT 49.215 136.425 55.525 136.725 ;
        RECT 49.215 136.410 49.545 136.425 ;
        RECT 51.515 136.410 51.845 136.425 ;
        RECT 55.195 136.410 55.525 136.425 ;
        RECT 34.860 135.390 36.840 135.720 ;
        RECT 64.860 135.390 66.840 135.720 ;
        RECT 94.860 135.390 96.840 135.720 ;
        RECT 19.860 132.670 21.840 133.000 ;
        RECT 49.860 132.670 51.840 133.000 ;
        RECT 79.860 132.670 81.840 133.000 ;
        RECT 109.860 132.670 111.840 133.000 ;
        RECT 63.680 131.965 64.060 131.975 ;
        RECT 64.855 131.965 65.185 131.980 ;
        RECT 63.680 131.665 65.185 131.965 ;
        RECT 63.680 131.655 64.060 131.665 ;
        RECT 64.855 131.650 65.185 131.665 ;
        RECT 34.860 129.950 36.840 130.280 ;
        RECT 64.860 129.950 66.840 130.280 ;
        RECT 94.860 129.950 96.840 130.280 ;
        RECT 19.860 127.230 21.840 127.560 ;
        RECT 49.860 127.230 51.840 127.560 ;
        RECT 79.860 127.230 81.840 127.560 ;
        RECT 109.860 127.230 111.840 127.560 ;
        RECT 34.860 124.510 36.840 124.840 ;
        RECT 64.860 124.510 66.840 124.840 ;
        RECT 94.860 124.510 96.840 124.840 ;
        RECT 57.240 123.125 57.620 123.135 ;
        RECT 86.015 123.125 86.345 123.140 ;
        RECT 57.240 122.825 86.345 123.125 ;
        RECT 57.240 122.815 57.620 122.825 ;
        RECT 19.860 121.790 21.840 122.120 ;
        RECT 49.860 121.790 51.840 122.120 ;
        RECT 24.835 121.085 25.165 121.100 ;
        RECT 59.120 121.085 59.420 122.825 ;
        RECT 86.015 122.810 86.345 122.825 ;
        RECT 79.860 121.790 81.840 122.120 ;
        RECT 109.860 121.790 111.840 122.120 ;
        RECT 24.835 120.785 59.420 121.085 ;
        RECT 24.835 120.770 25.165 120.785 ;
        RECT 41.640 120.420 41.940 120.785 ;
        RECT 41.640 120.105 42.185 120.420 ;
        RECT 41.855 120.090 42.185 120.105 ;
        RECT 34.860 119.070 36.840 119.400 ;
        RECT 64.860 119.070 66.840 119.400 ;
        RECT 94.860 119.070 96.840 119.400 ;
        RECT 19.860 116.350 21.840 116.680 ;
        RECT 49.860 116.350 51.840 116.680 ;
        RECT 79.860 116.350 81.840 116.680 ;
        RECT 109.860 116.350 111.840 116.680 ;
        RECT 34.860 113.630 36.840 113.960 ;
        RECT 64.860 113.630 66.840 113.960 ;
        RECT 94.860 113.630 96.840 113.960 ;
        RECT 68.535 113.615 68.865 113.620 ;
        RECT 68.280 113.605 68.865 113.615 ;
        RECT 68.080 113.305 68.865 113.605 ;
        RECT 68.280 113.295 68.865 113.305 ;
        RECT 68.535 113.290 68.865 113.295 ;
        RECT 19.860 110.910 21.840 111.240 ;
        RECT 49.860 110.910 51.840 111.240 ;
        RECT 79.860 110.910 81.840 111.240 ;
        RECT 109.860 110.910 111.840 111.240 ;
        RECT 34.860 108.190 36.840 108.520 ;
        RECT 64.860 108.190 66.840 108.520 ;
        RECT 94.860 108.190 96.840 108.520 ;
        RECT 119.370 106.820 121.370 106.955 ;
        RECT 119.135 106.490 121.370 106.820 ;
        RECT 119.370 106.355 121.370 106.490 ;
        RECT 19.860 105.470 21.840 105.800 ;
        RECT 49.860 105.470 51.840 105.800 ;
        RECT 79.860 105.470 81.840 105.800 ;
        RECT 109.860 105.470 111.840 105.800 ;
        RECT 129.700 105.605 133.210 106.625 ;
        RECT 34.860 102.750 36.840 103.080 ;
        RECT 64.860 102.750 66.840 103.080 ;
        RECT 94.860 102.750 96.840 103.080 ;
        RECT 37.630 88.620 38.970 88.755 ;
        RECT 13.950 87.980 14.980 88.515 ;
        RECT 13.950 87.500 14.990 87.980 ;
        RECT 13.950 87.175 14.980 87.500 ;
        RECT 14.070 86.570 14.810 87.175 ;
        RECT 20.050 87.105 20.920 88.515 ;
        RECT 14.070 75.715 14.700 86.570 ;
        RECT 20.170 77.115 20.800 87.105 ;
        RECT 25.910 87.055 26.860 88.515 ;
        RECT 26.070 78.385 26.700 87.055 ;
        RECT 31.730 86.965 32.910 88.585 ;
        RECT 32.005 79.615 32.635 86.965 ;
        RECT 37.630 86.835 39.120 88.620 ;
        RECT 38.060 81.125 38.690 86.835 ;
        RECT 43.790 86.745 45.190 88.605 ;
        RECT 49.710 86.945 51.060 88.615 ;
        RECT 44.175 82.625 44.805 86.745 ;
        RECT 50.070 83.875 50.700 86.945 ;
        RECT 55.530 86.785 56.750 88.545 ;
        RECT 55.825 85.115 56.455 86.785 ;
        RECT 61.670 86.625 63.180 88.615 ;
        RECT 67.680 88.305 68.720 89.815 ;
        RECT 67.885 87.225 68.515 88.305 ;
        RECT 62.110 86.175 62.740 86.625 ;
        RECT 67.885 86.595 130.605 87.225 ;
        RECT 62.110 85.545 118.855 86.175 ;
        RECT 55.825 84.485 107.605 85.115 ;
        RECT 50.070 83.245 96.285 83.875 ;
        RECT 44.175 81.995 85.055 82.625 ;
        RECT 38.060 80.495 73.765 81.125 ;
        RECT 32.005 78.985 62.635 79.615 ;
        RECT 26.070 77.755 51.245 78.385 ;
        RECT 20.170 76.485 40.645 77.115 ;
        RECT 14.070 75.660 29.295 75.715 ;
        RECT 40.015 75.710 40.645 76.485 ;
        RECT 14.070 75.085 30.410 75.660 ;
        RECT 27.850 74.670 30.410 75.085 ;
        RECT 3.910 71.345 6.100 73.215 ;
        RECT 27.850 73.120 30.450 74.670 ;
        RECT 39.060 74.510 41.620 75.710 ;
        RECT 50.615 75.580 51.245 77.755 ;
        RECT 62.005 75.690 62.635 78.985 ;
        RECT 49.930 74.650 52.490 75.580 ;
        RECT 0.970 70.330 3.070 70.430 ;
        RECT 15.510 70.330 17.040 71.185 ;
        RECT 0.960 68.750 17.040 70.330 ;
        RECT 0.970 68.710 3.070 68.750 ;
        RECT 15.510 68.635 17.040 68.750 ;
        RECT 20.145 54.060 20.605 54.135 ;
        RECT 25.715 54.060 26.175 54.085 ;
        RECT 20.145 53.620 26.175 54.060 ;
        RECT 20.145 53.565 20.605 53.620 ;
        RECT 25.715 53.515 26.175 53.620 ;
        RECT 22.405 48.870 22.885 48.935 ;
        RECT 22.405 48.550 24.205 48.870 ;
        RECT 22.405 48.385 22.885 48.550 ;
        RECT 23.635 45.710 24.195 48.550 ;
        RECT 27.515 45.710 27.995 45.735 ;
        RECT 23.635 45.290 27.995 45.710 ;
        RECT 23.635 45.280 24.195 45.290 ;
        RECT 27.515 45.185 27.995 45.290 ;
        RECT 20.745 40.120 21.225 40.225 ;
        RECT 24.545 40.120 25.105 40.130 ;
        RECT 20.745 39.700 25.105 40.120 ;
        RECT 20.745 39.675 21.225 39.700 ;
        RECT 24.545 36.860 25.105 39.700 ;
        RECT 25.855 36.860 26.335 37.025 ;
        RECT 24.535 36.540 26.335 36.860 ;
        RECT 25.855 36.475 26.335 36.540 ;
        RECT 22.565 31.790 23.025 31.895 ;
        RECT 28.135 31.790 28.595 31.845 ;
        RECT 22.565 31.350 28.595 31.790 ;
        RECT 22.565 31.325 23.025 31.350 ;
        RECT 28.135 31.275 28.595 31.350 ;
        RECT 29.765 12.265 30.255 73.120 ;
        RECT 38.960 73.080 41.730 74.510 ;
        RECT 31.345 54.070 31.805 54.145 ;
        RECT 36.915 54.070 37.375 54.095 ;
        RECT 31.345 53.630 37.375 54.070 ;
        RECT 31.345 53.575 31.805 53.630 ;
        RECT 36.915 53.525 37.375 53.630 ;
        RECT 33.605 48.880 34.085 48.945 ;
        RECT 33.605 48.560 35.405 48.880 ;
        RECT 33.605 48.395 34.085 48.560 ;
        RECT 34.835 45.720 35.395 48.560 ;
        RECT 38.715 45.720 39.195 45.745 ;
        RECT 34.835 45.300 39.195 45.720 ;
        RECT 34.835 45.290 35.395 45.300 ;
        RECT 38.715 45.195 39.195 45.300 ;
        RECT 32.025 40.120 32.505 40.225 ;
        RECT 35.825 40.120 36.385 40.130 ;
        RECT 32.025 39.700 36.385 40.120 ;
        RECT 32.025 39.675 32.505 39.700 ;
        RECT 35.825 36.860 36.385 39.700 ;
        RECT 37.135 36.860 37.615 37.025 ;
        RECT 35.815 36.540 37.615 36.860 ;
        RECT 37.135 36.475 37.615 36.540 ;
        RECT 33.845 31.790 34.305 31.895 ;
        RECT 39.415 31.790 39.875 31.845 ;
        RECT 33.845 31.350 39.875 31.790 ;
        RECT 33.845 31.325 34.305 31.350 ;
        RECT 39.415 31.275 39.875 31.350 ;
        RECT 41.055 12.360 41.545 73.080 ;
        RECT 49.930 73.030 52.530 74.650 ;
        RECT 61.330 74.530 63.890 75.690 ;
        RECT 73.135 75.580 73.765 80.495 ;
        RECT 84.425 75.690 85.055 81.995 ;
        RECT 72.340 74.980 74.900 75.580 ;
        RECT 42.565 54.040 43.025 54.115 ;
        RECT 48.135 54.040 48.595 54.065 ;
        RECT 42.565 53.600 48.595 54.040 ;
        RECT 42.565 53.545 43.025 53.600 ;
        RECT 48.135 53.495 48.595 53.600 ;
        RECT 44.825 48.850 45.305 48.915 ;
        RECT 44.825 48.530 46.625 48.850 ;
        RECT 44.825 48.365 45.305 48.530 ;
        RECT 46.055 45.690 46.615 48.530 ;
        RECT 49.935 45.690 50.415 45.715 ;
        RECT 46.055 45.270 50.415 45.690 ;
        RECT 46.055 45.260 46.615 45.270 ;
        RECT 49.935 45.165 50.415 45.270 ;
        RECT 43.315 40.100 43.795 40.205 ;
        RECT 47.115 40.100 47.675 40.110 ;
        RECT 43.315 39.680 47.675 40.100 ;
        RECT 43.315 39.655 43.795 39.680 ;
        RECT 47.115 36.840 47.675 39.680 ;
        RECT 48.425 36.840 48.905 37.005 ;
        RECT 47.105 36.520 48.905 36.840 ;
        RECT 48.425 36.455 48.905 36.520 ;
        RECT 45.135 31.770 45.595 31.875 ;
        RECT 50.705 31.770 51.165 31.825 ;
        RECT 45.135 31.330 51.165 31.770 ;
        RECT 45.135 31.305 45.595 31.330 ;
        RECT 50.705 31.255 51.165 31.330 ;
        RECT 41.055 12.350 41.555 12.360 ;
        RECT 28.345 11.115 30.465 12.265 ;
        RECT 41.065 11.965 41.555 12.350 ;
        RECT 51.635 12.145 52.125 73.030 ;
        RECT 61.260 73.010 64.060 74.530 ;
        RECT 72.340 73.050 75.020 74.980 ;
        RECT 83.730 74.540 86.290 75.690 ;
        RECT 95.655 75.580 96.285 83.245 ;
        RECT 106.975 75.640 107.605 84.485 ;
        RECT 118.225 75.650 118.855 85.545 ;
        RECT 129.975 75.650 130.605 86.595 ;
        RECT 133.330 76.605 136.060 77.855 ;
        RECT 137.190 76.585 139.920 77.835 ;
        RECT 53.815 54.020 54.275 54.095 ;
        RECT 59.385 54.020 59.845 54.045 ;
        RECT 53.815 53.580 59.845 54.020 ;
        RECT 53.815 53.525 54.275 53.580 ;
        RECT 59.385 53.475 59.845 53.580 ;
        RECT 56.075 48.830 56.555 48.895 ;
        RECT 56.075 48.510 57.875 48.830 ;
        RECT 56.075 48.345 56.555 48.510 ;
        RECT 57.305 45.670 57.865 48.510 ;
        RECT 61.185 45.670 61.665 45.695 ;
        RECT 57.305 45.250 61.665 45.670 ;
        RECT 57.305 45.240 57.865 45.250 ;
        RECT 61.185 45.145 61.665 45.250 ;
        RECT 54.535 40.100 55.015 40.205 ;
        RECT 58.335 40.100 58.895 40.110 ;
        RECT 54.535 39.680 58.895 40.100 ;
        RECT 54.535 39.655 55.015 39.680 ;
        RECT 58.335 36.840 58.895 39.680 ;
        RECT 59.645 36.840 60.125 37.005 ;
        RECT 58.325 36.520 60.125 36.840 ;
        RECT 59.645 36.455 60.125 36.520 ;
        RECT 56.355 31.770 56.815 31.875 ;
        RECT 61.925 31.770 62.385 31.825 ;
        RECT 56.355 31.330 62.385 31.770 ;
        RECT 56.355 31.305 56.815 31.330 ;
        RECT 61.925 31.255 62.385 31.330 ;
        RECT 29.765 11.100 30.255 11.115 ;
        RECT 39.065 11.005 41.615 11.965 ;
        RECT 50.285 10.995 52.405 12.145 ;
        RECT 62.915 12.135 63.405 73.010 ;
        RECT 65.035 54.010 65.495 54.085 ;
        RECT 70.605 54.010 71.065 54.035 ;
        RECT 65.035 53.570 71.065 54.010 ;
        RECT 65.035 53.515 65.495 53.570 ;
        RECT 70.605 53.465 71.065 53.570 ;
        RECT 67.295 48.820 67.775 48.885 ;
        RECT 67.295 48.500 69.095 48.820 ;
        RECT 67.295 48.335 67.775 48.500 ;
        RECT 68.525 45.660 69.085 48.500 ;
        RECT 72.405 45.660 72.885 45.685 ;
        RECT 68.525 45.240 72.885 45.660 ;
        RECT 68.525 45.230 69.085 45.240 ;
        RECT 72.405 45.135 72.885 45.240 ;
        RECT 65.735 40.100 66.215 40.205 ;
        RECT 69.535 40.100 70.095 40.110 ;
        RECT 65.735 39.680 70.095 40.100 ;
        RECT 65.735 39.655 66.215 39.680 ;
        RECT 69.535 36.840 70.095 39.680 ;
        RECT 70.845 36.840 71.325 37.005 ;
        RECT 69.525 36.520 71.325 36.840 ;
        RECT 70.845 36.455 71.325 36.520 ;
        RECT 67.555 31.770 68.015 31.875 ;
        RECT 73.125 31.770 73.585 31.825 ;
        RECT 67.555 31.330 73.585 31.770 ;
        RECT 67.555 31.305 68.015 31.330 ;
        RECT 73.125 31.255 73.585 31.330 ;
        RECT 74.055 12.165 74.545 73.050 ;
        RECT 83.690 73.000 86.290 74.540 ;
        RECT 94.960 74.710 97.520 75.580 ;
        RECT 94.960 73.020 97.570 74.710 ;
        RECT 106.340 74.460 108.900 75.640 ;
        RECT 117.470 74.720 120.030 75.650 ;
        RECT 76.275 54.000 76.735 54.075 ;
        RECT 81.845 54.000 82.305 54.025 ;
        RECT 76.275 53.560 82.305 54.000 ;
        RECT 76.275 53.505 76.735 53.560 ;
        RECT 81.845 53.455 82.305 53.560 ;
        RECT 78.535 48.810 79.015 48.875 ;
        RECT 78.535 48.490 80.335 48.810 ;
        RECT 78.535 48.325 79.015 48.490 ;
        RECT 79.765 45.650 80.325 48.490 ;
        RECT 83.645 45.650 84.125 45.675 ;
        RECT 79.765 45.230 84.125 45.650 ;
        RECT 79.765 45.220 80.325 45.230 ;
        RECT 83.645 45.125 84.125 45.230 ;
        RECT 77.025 40.090 77.505 40.195 ;
        RECT 80.825 40.090 81.385 40.100 ;
        RECT 77.025 39.670 81.385 40.090 ;
        RECT 77.025 39.645 77.505 39.670 ;
        RECT 80.825 36.830 81.385 39.670 ;
        RECT 82.135 36.830 82.615 36.995 ;
        RECT 80.815 36.510 82.615 36.830 ;
        RECT 82.135 36.445 82.615 36.510 ;
        RECT 78.845 31.760 79.305 31.865 ;
        RECT 84.415 31.760 84.875 31.815 ;
        RECT 78.845 31.320 84.875 31.760 ;
        RECT 78.845 31.295 79.305 31.320 ;
        RECT 84.415 31.245 84.875 31.320 ;
        RECT 61.365 10.985 63.485 12.135 ;
        RECT 72.675 11.015 74.795 12.165 ;
        RECT 85.375 12.155 85.865 73.000 ;
        RECT 87.525 54.010 87.985 54.085 ;
        RECT 93.095 54.010 93.555 54.035 ;
        RECT 87.525 53.570 93.555 54.010 ;
        RECT 87.525 53.515 87.985 53.570 ;
        RECT 93.095 53.465 93.555 53.570 ;
        RECT 89.785 48.820 90.265 48.885 ;
        RECT 89.785 48.500 91.585 48.820 ;
        RECT 89.785 48.335 90.265 48.500 ;
        RECT 91.015 45.660 91.575 48.500 ;
        RECT 94.895 45.660 95.375 45.685 ;
        RECT 91.015 45.240 95.375 45.660 ;
        RECT 91.015 45.230 91.575 45.240 ;
        RECT 94.895 45.135 95.375 45.240 ;
        RECT 88.265 40.110 88.745 40.215 ;
        RECT 92.065 40.110 92.625 40.120 ;
        RECT 88.265 39.690 92.625 40.110 ;
        RECT 88.265 39.665 88.745 39.690 ;
        RECT 92.065 36.850 92.625 39.690 ;
        RECT 93.375 36.850 93.855 37.015 ;
        RECT 92.055 36.530 93.855 36.850 ;
        RECT 93.375 36.465 93.855 36.530 ;
        RECT 90.085 31.780 90.545 31.885 ;
        RECT 95.655 31.780 96.115 31.835 ;
        RECT 90.085 31.340 96.115 31.780 ;
        RECT 90.085 31.315 90.545 31.340 ;
        RECT 95.655 31.265 96.115 31.340 ;
        RECT 96.605 12.155 97.095 73.020 ;
        RECT 106.150 73.000 109.060 74.460 ;
        RECT 117.470 73.070 120.000 74.720 ;
        RECT 129.290 74.650 131.850 75.650 ;
        RECT 129.300 73.140 131.820 74.650 ;
        RECT 98.805 54.000 99.265 54.075 ;
        RECT 104.375 54.000 104.835 54.025 ;
        RECT 98.805 53.560 104.835 54.000 ;
        RECT 98.805 53.505 99.265 53.560 ;
        RECT 104.375 53.455 104.835 53.560 ;
        RECT 101.065 48.810 101.545 48.875 ;
        RECT 101.065 48.490 102.865 48.810 ;
        RECT 101.065 48.325 101.545 48.490 ;
        RECT 102.295 45.650 102.855 48.490 ;
        RECT 106.175 45.650 106.655 45.675 ;
        RECT 102.295 45.230 106.655 45.650 ;
        RECT 102.295 45.220 102.855 45.230 ;
        RECT 106.175 45.125 106.655 45.230 ;
        RECT 99.475 40.130 99.955 40.235 ;
        RECT 103.275 40.130 103.835 40.140 ;
        RECT 99.475 39.710 103.835 40.130 ;
        RECT 99.475 39.685 99.955 39.710 ;
        RECT 103.275 36.870 103.835 39.710 ;
        RECT 104.585 36.870 105.065 37.035 ;
        RECT 103.265 36.550 105.065 36.870 ;
        RECT 104.585 36.485 105.065 36.550 ;
        RECT 101.295 31.800 101.755 31.905 ;
        RECT 106.865 31.800 107.325 31.855 ;
        RECT 101.295 31.360 107.325 31.800 ;
        RECT 101.295 31.335 101.755 31.360 ;
        RECT 106.865 31.285 107.325 31.360 ;
        RECT 107.865 12.205 108.355 73.000 ;
        RECT 110.075 54.000 110.535 54.075 ;
        RECT 115.645 54.000 116.105 54.025 ;
        RECT 110.075 53.560 116.105 54.000 ;
        RECT 110.075 53.505 110.535 53.560 ;
        RECT 115.645 53.455 116.105 53.560 ;
        RECT 112.335 48.810 112.815 48.875 ;
        RECT 112.335 48.490 114.135 48.810 ;
        RECT 112.335 48.325 112.815 48.490 ;
        RECT 113.565 45.650 114.125 48.490 ;
        RECT 117.445 45.650 117.925 45.675 ;
        RECT 113.565 45.230 117.925 45.650 ;
        RECT 113.565 45.220 114.125 45.230 ;
        RECT 117.445 45.125 117.925 45.230 ;
        RECT 110.675 40.170 111.155 40.275 ;
        RECT 114.475 40.170 115.035 40.180 ;
        RECT 110.675 39.750 115.035 40.170 ;
        RECT 110.675 39.725 111.155 39.750 ;
        RECT 114.475 36.910 115.035 39.750 ;
        RECT 115.785 36.910 116.265 37.075 ;
        RECT 114.465 36.590 116.265 36.910 ;
        RECT 115.785 36.525 116.265 36.590 ;
        RECT 112.495 31.840 112.955 31.945 ;
        RECT 118.065 31.840 118.525 31.895 ;
        RECT 112.495 31.400 118.525 31.840 ;
        RECT 112.495 31.375 112.955 31.400 ;
        RECT 118.065 31.325 118.525 31.400 ;
        RECT 119.085 12.205 119.575 73.070 ;
        RECT 121.325 54.000 121.785 54.075 ;
        RECT 126.895 54.000 127.355 54.025 ;
        RECT 121.325 53.560 127.355 54.000 ;
        RECT 121.325 53.505 121.785 53.560 ;
        RECT 126.895 53.455 127.355 53.560 ;
        RECT 123.585 48.810 124.065 48.875 ;
        RECT 123.585 48.490 125.385 48.810 ;
        RECT 123.585 48.325 124.065 48.490 ;
        RECT 124.815 45.650 125.375 48.490 ;
        RECT 128.695 45.650 129.175 45.675 ;
        RECT 124.815 45.230 129.175 45.650 ;
        RECT 124.815 45.220 125.375 45.230 ;
        RECT 128.695 45.125 129.175 45.230 ;
        RECT 121.885 40.190 122.365 40.295 ;
        RECT 125.685 40.190 126.245 40.200 ;
        RECT 121.885 39.770 126.245 40.190 ;
        RECT 121.885 39.745 122.365 39.770 ;
        RECT 125.685 36.930 126.245 39.770 ;
        RECT 126.995 36.930 127.475 37.095 ;
        RECT 125.675 36.610 127.475 36.930 ;
        RECT 126.995 36.545 127.475 36.610 ;
        RECT 123.705 31.860 124.165 31.965 ;
        RECT 129.275 31.860 129.735 31.915 ;
        RECT 123.705 31.420 129.735 31.860 ;
        RECT 123.705 31.395 124.165 31.420 ;
        RECT 129.275 31.345 129.735 31.420 ;
        RECT 130.335 12.235 130.825 73.140 ;
        RECT 74.055 11.010 74.545 11.015 ;
        RECT 83.795 11.005 85.915 12.155 ;
        RECT 95.095 11.005 97.215 12.155 ;
        RECT 106.285 11.055 108.405 12.205 ;
        RECT 117.515 11.055 119.635 12.205 ;
        RECT 128.815 11.085 130.935 12.235 ;
        RECT 107.865 11.010 108.355 11.055 ;
        RECT 119.085 11.050 119.575 11.055 ;
        RECT 85.375 11.000 85.865 11.005 ;
        RECT 96.605 10.980 97.095 11.005 ;
        RECT 74.290 0.135 75.680 1.435 ;
        RECT 93.500 0.205 94.890 1.505 ;
        RECT 112.900 0.335 114.290 1.635 ;
        RECT 131.800 0.405 133.540 1.905 ;
        RECT 151.600 0.275 152.970 1.445 ;
      LAYER met4 ;
        RECT 30.420 225.130 30.670 225.140 ;
        RECT 30.300 224.760 30.670 225.130 ;
        RECT 30.970 224.760 33.430 225.140 ;
        RECT 33.730 224.760 36.190 225.140 ;
        RECT 36.490 224.760 38.950 225.140 ;
        RECT 39.250 224.760 41.710 225.140 ;
        RECT 42.010 224.760 44.470 225.140 ;
        RECT 44.770 224.760 47.230 225.140 ;
        RECT 47.530 224.760 49.990 225.140 ;
        RECT 50.290 224.760 52.750 225.140 ;
        RECT 53.050 224.760 55.510 225.140 ;
        RECT 55.810 224.760 58.270 225.140 ;
        RECT 58.570 224.760 61.030 225.140 ;
        RECT 61.330 224.760 63.790 225.140 ;
        RECT 64.090 224.760 66.550 225.140 ;
        RECT 66.850 224.760 69.310 225.140 ;
        RECT 69.610 224.760 72.070 225.140 ;
        RECT 72.370 224.760 74.830 225.140 ;
        RECT 75.130 224.760 77.590 225.140 ;
        RECT 77.890 224.760 80.350 225.140 ;
        RECT 80.650 224.760 83.110 225.140 ;
        RECT 83.410 224.760 85.870 225.140 ;
        RECT 86.170 224.760 88.630 225.140 ;
        RECT 88.930 224.760 91.390 225.140 ;
        RECT 91.690 224.760 94.150 225.140 ;
        RECT 94.450 224.760 96.910 225.140 ;
        RECT 97.210 224.760 99.670 225.140 ;
        RECT 99.970 224.760 102.430 225.140 ;
        RECT 102.730 224.760 105.190 225.140 ;
        RECT 105.490 224.760 107.950 225.140 ;
        RECT 108.250 224.760 110.710 225.140 ;
        RECT 111.010 224.760 113.470 225.140 ;
        RECT 113.770 224.760 116.230 225.140 ;
        RECT 116.530 224.760 118.990 225.140 ;
        RECT 119.290 224.760 121.750 225.140 ;
        RECT 122.050 224.760 124.510 225.140 ;
        RECT 124.810 224.760 127.270 225.140 ;
        RECT 127.570 224.760 130.030 225.140 ;
        RECT 130.330 224.760 132.790 225.140 ;
        RECT 133.090 224.760 133.520 225.140 ;
        RECT 30.300 224.240 133.520 224.760 ;
        RECT 135.385 224.760 135.550 225.185 ;
        RECT 135.850 224.760 136.745 225.185 ;
        RECT 30.300 219.100 31.660 224.240 ;
        RECT 135.385 223.875 136.745 224.760 ;
        RECT 138.175 224.760 138.310 225.115 ;
        RECT 138.610 224.760 139.535 225.115 ;
        RECT 138.175 223.805 139.535 224.760 ;
        RECT 143.225 224.760 143.830 225.145 ;
        RECT 144.130 224.760 144.585 225.145 ;
        RECT 143.225 223.835 144.585 224.760 ;
        RECT 6.000 218.040 31.660 219.100 ;
        RECT 30.300 217.960 31.660 218.040 ;
        RECT 19.850 102.675 21.850 206.515 ;
        RECT 34.850 102.675 36.850 206.515 ;
        RECT 38.865 176.530 39.195 176.860 ;
        RECT 38.880 140.820 39.180 176.530 ;
        RECT 38.865 140.490 39.195 140.820 ;
        RECT 49.850 102.675 51.850 206.515 ;
        RECT 63.705 182.650 64.035 182.980 ;
        RECT 57.265 171.770 57.595 172.100 ;
        RECT 57.280 149.660 57.580 171.770 ;
        RECT 57.265 149.330 57.595 149.660 ;
        RECT 57.280 123.140 57.580 149.330 ;
        RECT 63.720 131.980 64.020 182.650 ;
        RECT 63.705 131.650 64.035 131.980 ;
        RECT 57.265 122.810 57.595 123.140 ;
        RECT 64.850 102.675 66.850 206.515 ;
        RECT 68.305 149.330 68.635 149.660 ;
        RECT 68.320 113.620 68.620 149.330 ;
        RECT 68.305 113.290 68.635 113.620 ;
        RECT 79.850 102.675 81.850 206.515 ;
        RECT 94.850 102.675 96.850 206.515 ;
        RECT 100.505 150.010 100.835 150.340 ;
        RECT 100.520 139.460 100.820 150.010 ;
        RECT 100.505 139.130 100.835 139.460 ;
        RECT 109.850 102.675 111.850 206.515 ;
        RECT 118.110 97.700 120.130 99.670 ;
        RECT 121.810 97.750 123.830 99.720 ;
        RECT 118.130 93.980 120.130 97.700 ;
        RECT 121.820 96.830 123.820 97.750 ;
        RECT 121.820 94.830 139.410 96.830 ;
        RECT 118.130 91.980 135.580 93.980 ;
        RECT 133.580 77.835 135.580 91.980 ;
        RECT 133.375 76.625 136.015 77.835 ;
        RECT 137.410 77.815 139.410 94.830 ;
        RECT 137.235 76.605 139.875 77.815 ;
        RECT 3.955 71.365 4.000 73.195 ;
        RECT 6.000 71.365 6.055 73.195 ;
        RECT 3.000 68.705 3.025 70.435 ;
        RECT 15.555 68.655 16.995 71.165 ;
        RECT 74.335 1.000 75.635 1.415 ;
        RECT 74.335 0.155 74.530 1.000 ;
        RECT 75.430 0.155 75.635 1.000 ;
        RECT 93.545 1.000 94.845 1.485 ;
        RECT 93.545 0.225 93.850 1.000 ;
        RECT 94.750 0.225 94.845 1.000 ;
        RECT 112.945 1.000 114.245 1.615 ;
        RECT 112.945 0.355 113.170 1.000 ;
        RECT 114.070 0.355 114.245 1.000 ;
        RECT 131.845 1.000 133.495 1.885 ;
        RECT 131.845 0.425 132.490 1.000 ;
        RECT 133.390 0.425 133.495 1.000 ;
        RECT 151.645 1.000 152.925 1.425 ;
        RECT 151.645 0.295 151.810 1.000 ;
        RECT 152.710 0.295 152.925 1.000 ;
  END
END tt_um_08_sws
END LIBRARY

