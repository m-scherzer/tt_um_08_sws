VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_08_sws
  CLASS BLOCK ;
  FOREIGN tt_um_08_sws ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 200.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNAGATEAREA 932.310486 ;
    ANTENNADIFFAREA 1102.580322 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 14.805 211.185 14.975 211.375 ;
        RECT 18.485 211.185 18.655 211.375 ;
        RECT 24.005 211.185 24.175 211.375 ;
        RECT 25.845 211.185 26.015 211.375 ;
        RECT 31.365 211.185 31.535 211.375 ;
        RECT 36.885 211.185 37.055 211.375 ;
        RECT 38.725 211.185 38.895 211.375 ;
        RECT 44.245 211.185 44.415 211.375 ;
        RECT 49.765 211.185 49.935 211.375 ;
        RECT 51.605 211.185 51.775 211.375 ;
        RECT 57.125 211.185 57.295 211.375 ;
        RECT 62.645 211.185 62.815 211.375 ;
        RECT 64.485 211.185 64.655 211.375 ;
        RECT 70.005 211.185 70.175 211.375 ;
        RECT 75.525 211.185 75.695 211.375 ;
        RECT 77.365 211.185 77.535 211.375 ;
        RECT 82.885 211.185 83.055 211.375 ;
        RECT 88.405 211.185 88.575 211.375 ;
        RECT 90.245 211.185 90.415 211.375 ;
        RECT 95.765 211.185 95.935 211.375 ;
        RECT 101.285 211.185 101.455 211.375 ;
        RECT 103.125 211.185 103.295 211.375 ;
        RECT 108.645 211.185 108.815 211.375 ;
        RECT 114.165 211.185 114.335 211.375 ;
        RECT 115.140 211.235 115.260 211.345 ;
        RECT 120.605 211.185 120.775 211.375 ;
        RECT 126.125 211.185 126.295 211.375 ;
        RECT 127.505 211.185 127.675 211.375 ;
        RECT 14.665 210.375 16.035 211.185 ;
        RECT 16.045 210.375 18.795 211.185 ;
        RECT 18.805 210.375 24.315 211.185 ;
        RECT 24.335 210.315 24.765 211.100 ;
        RECT 24.785 210.375 26.155 211.185 ;
        RECT 26.165 210.375 31.675 211.185 ;
        RECT 31.685 210.375 37.195 211.185 ;
        RECT 37.215 210.315 37.645 211.100 ;
        RECT 37.665 210.375 39.035 211.185 ;
        RECT 39.045 210.375 44.555 211.185 ;
        RECT 44.565 210.375 50.075 211.185 ;
        RECT 50.095 210.315 50.525 211.100 ;
        RECT 50.545 210.375 51.915 211.185 ;
        RECT 51.925 210.375 57.435 211.185 ;
        RECT 57.445 210.375 62.955 211.185 ;
        RECT 62.975 210.315 63.405 211.100 ;
        RECT 63.425 210.375 64.795 211.185 ;
        RECT 64.805 210.375 70.315 211.185 ;
        RECT 70.325 210.375 75.835 211.185 ;
        RECT 75.855 210.315 76.285 211.100 ;
        RECT 76.305 210.375 77.675 211.185 ;
        RECT 77.685 210.375 83.195 211.185 ;
        RECT 83.205 210.375 88.715 211.185 ;
        RECT 88.735 210.315 89.165 211.100 ;
        RECT 89.185 210.375 90.555 211.185 ;
        RECT 90.565 210.375 96.075 211.185 ;
        RECT 96.085 210.375 101.595 211.185 ;
        RECT 101.615 210.315 102.045 211.100 ;
        RECT 102.065 210.375 103.435 211.185 ;
        RECT 103.445 210.375 108.955 211.185 ;
        RECT 108.965 210.375 114.475 211.185 ;
        RECT 114.495 210.315 114.925 211.100 ;
        RECT 115.405 210.375 120.915 211.185 ;
        RECT 120.925 210.375 126.435 211.185 ;
        RECT 126.445 210.375 127.815 211.185 ;
      LAYER nwell ;
        RECT 14.470 207.155 128.010 209.985 ;
      LAYER pwell ;
        RECT 14.665 205.955 16.035 206.765 ;
        RECT 16.045 205.955 18.795 206.765 ;
        RECT 18.805 205.955 24.315 206.765 ;
        RECT 24.335 206.040 24.765 206.825 ;
        RECT 25.245 205.955 27.995 206.765 ;
        RECT 28.005 205.955 33.515 206.765 ;
        RECT 33.525 205.955 39.035 206.765 ;
        RECT 39.045 205.955 44.555 206.765 ;
        RECT 44.565 205.955 50.075 206.765 ;
        RECT 50.095 206.040 50.525 206.825 ;
        RECT 51.005 205.955 53.755 206.765 ;
        RECT 53.765 205.955 59.275 206.765 ;
        RECT 59.285 205.955 64.795 206.765 ;
        RECT 64.805 205.955 70.315 206.765 ;
        RECT 70.325 205.955 75.835 206.765 ;
        RECT 75.855 206.040 76.285 206.825 ;
        RECT 76.765 205.955 79.515 206.765 ;
        RECT 79.525 205.955 85.035 206.765 ;
        RECT 85.045 205.955 90.555 206.765 ;
        RECT 90.565 205.955 96.075 206.765 ;
        RECT 96.085 205.955 101.595 206.765 ;
        RECT 101.615 206.040 102.045 206.825 ;
        RECT 102.525 205.955 104.355 206.765 ;
        RECT 104.365 205.955 109.875 206.765 ;
        RECT 109.885 205.955 115.395 206.765 ;
        RECT 115.405 205.955 120.915 206.765 ;
        RECT 120.925 205.955 126.435 206.765 ;
        RECT 126.445 205.955 127.815 206.765 ;
        RECT 14.805 205.745 14.975 205.955 ;
        RECT 16.645 205.790 16.805 205.900 ;
        RECT 18.485 205.765 18.655 205.955 ;
        RECT 20.325 205.745 20.495 205.935 ;
        RECT 24.005 205.765 24.175 205.955 ;
        RECT 24.980 205.795 25.100 205.905 ;
        RECT 25.845 205.745 26.015 205.935 ;
        RECT 27.685 205.765 27.855 205.955 ;
        RECT 31.365 205.745 31.535 205.935 ;
        RECT 33.205 205.765 33.375 205.955 ;
        RECT 36.885 205.745 37.055 205.935 ;
        RECT 37.860 205.795 37.980 205.905 ;
        RECT 38.725 205.765 38.895 205.955 ;
        RECT 40.565 205.745 40.735 205.935 ;
        RECT 44.245 205.765 44.415 205.955 ;
        RECT 46.085 205.745 46.255 205.935 ;
        RECT 49.765 205.765 49.935 205.955 ;
        RECT 50.740 205.795 50.860 205.905 ;
        RECT 51.605 205.745 51.775 205.935 ;
        RECT 53.445 205.765 53.615 205.955 ;
        RECT 57.125 205.745 57.295 205.935 ;
        RECT 58.965 205.765 59.135 205.955 ;
        RECT 62.645 205.745 62.815 205.935 ;
        RECT 63.620 205.795 63.740 205.905 ;
        RECT 64.485 205.765 64.655 205.955 ;
        RECT 66.325 205.745 66.495 205.935 ;
        RECT 70.005 205.765 70.175 205.955 ;
        RECT 71.845 205.745 72.015 205.935 ;
        RECT 75.525 205.765 75.695 205.955 ;
        RECT 76.500 205.795 76.620 205.905 ;
        RECT 77.365 205.745 77.535 205.935 ;
        RECT 79.205 205.765 79.375 205.955 ;
        RECT 82.885 205.745 83.055 205.935 ;
        RECT 84.725 205.765 84.895 205.955 ;
        RECT 88.405 205.745 88.575 205.935 ;
        RECT 89.380 205.795 89.500 205.905 ;
        RECT 90.245 205.765 90.415 205.955 ;
        RECT 92.085 205.745 92.255 205.935 ;
        RECT 95.765 205.765 95.935 205.955 ;
        RECT 97.605 205.745 97.775 205.935 ;
        RECT 101.285 205.765 101.455 205.955 ;
        RECT 102.260 205.795 102.380 205.905 ;
        RECT 103.125 205.745 103.295 205.935 ;
        RECT 104.045 205.765 104.215 205.955 ;
        RECT 108.645 205.745 108.815 205.935 ;
        RECT 109.565 205.765 109.735 205.955 ;
        RECT 114.165 205.745 114.335 205.935 ;
        RECT 115.085 205.905 115.255 205.955 ;
        RECT 115.085 205.795 115.260 205.905 ;
        RECT 115.085 205.765 115.255 205.795 ;
        RECT 120.605 205.745 120.775 205.955 ;
        RECT 126.125 205.745 126.295 205.955 ;
        RECT 127.505 205.745 127.675 205.955 ;
        RECT 14.665 204.935 16.035 205.745 ;
        RECT 16.965 204.935 20.635 205.745 ;
        RECT 20.645 204.935 26.155 205.745 ;
        RECT 26.165 204.935 31.675 205.745 ;
        RECT 31.685 204.935 37.195 205.745 ;
        RECT 37.215 204.875 37.645 205.660 ;
        RECT 38.125 204.935 40.875 205.745 ;
        RECT 40.885 204.935 46.395 205.745 ;
        RECT 46.405 204.935 51.915 205.745 ;
        RECT 51.925 204.935 57.435 205.745 ;
        RECT 57.445 204.935 62.955 205.745 ;
        RECT 62.975 204.875 63.405 205.660 ;
        RECT 63.885 204.935 66.635 205.745 ;
        RECT 66.645 204.935 72.155 205.745 ;
        RECT 72.165 204.935 77.675 205.745 ;
        RECT 77.685 204.935 83.195 205.745 ;
        RECT 83.205 204.935 88.715 205.745 ;
        RECT 88.735 204.875 89.165 205.660 ;
        RECT 89.645 204.935 92.395 205.745 ;
        RECT 92.405 204.935 97.915 205.745 ;
        RECT 97.925 204.935 103.435 205.745 ;
        RECT 103.445 204.935 108.955 205.745 ;
        RECT 108.965 204.935 114.475 205.745 ;
        RECT 114.495 204.875 114.925 205.660 ;
        RECT 115.405 204.935 120.915 205.745 ;
        RECT 120.925 204.935 126.435 205.745 ;
        RECT 126.445 204.935 127.815 205.745 ;
      LAYER nwell ;
        RECT 14.470 201.715 128.010 204.545 ;
      LAYER pwell ;
        RECT 14.665 200.515 16.035 201.325 ;
        RECT 16.045 200.515 18.795 201.325 ;
        RECT 18.805 200.515 24.315 201.325 ;
        RECT 24.335 200.600 24.765 201.385 ;
        RECT 25.245 200.515 27.995 201.325 ;
        RECT 28.005 200.515 33.515 201.325 ;
        RECT 33.525 200.515 39.035 201.325 ;
        RECT 39.045 200.515 44.555 201.325 ;
        RECT 44.565 200.515 50.075 201.325 ;
        RECT 50.095 200.600 50.525 201.385 ;
        RECT 51.005 200.515 52.835 201.325 ;
        RECT 52.845 200.515 58.355 201.325 ;
        RECT 58.405 201.195 59.745 201.425 ;
        RECT 62.575 201.195 63.505 201.415 ;
        RECT 58.405 200.515 68.015 201.195 ;
        RECT 68.485 200.515 70.315 201.325 ;
        RECT 70.325 200.515 75.835 201.325 ;
        RECT 75.855 200.600 76.285 201.385 ;
        RECT 76.765 200.515 79.515 201.325 ;
        RECT 79.525 200.515 85.035 201.325 ;
        RECT 85.045 200.515 90.555 201.325 ;
        RECT 90.565 200.515 96.075 201.325 ;
        RECT 96.085 200.515 101.595 201.325 ;
        RECT 101.615 200.600 102.045 201.385 ;
        RECT 102.525 200.515 104.355 201.325 ;
        RECT 104.365 200.515 109.875 201.325 ;
        RECT 109.885 200.515 115.395 201.325 ;
        RECT 115.405 200.515 120.915 201.325 ;
        RECT 120.925 200.515 126.435 201.325 ;
        RECT 126.445 200.515 127.815 201.325 ;
        RECT 14.805 200.305 14.975 200.515 ;
        RECT 16.645 200.350 16.805 200.460 ;
        RECT 18.485 200.325 18.655 200.515 ;
        RECT 20.325 200.305 20.495 200.495 ;
        RECT 24.005 200.325 24.175 200.515 ;
        RECT 24.980 200.355 25.100 200.465 ;
        RECT 25.845 200.305 26.015 200.495 ;
        RECT 27.685 200.325 27.855 200.515 ;
        RECT 31.365 200.305 31.535 200.495 ;
        RECT 33.205 200.325 33.375 200.515 ;
        RECT 36.885 200.305 37.055 200.495 ;
        RECT 38.725 200.325 38.895 200.515 ;
        RECT 39.185 200.305 39.355 200.495 ;
        RECT 44.245 200.325 44.415 200.515 ;
        RECT 44.705 200.305 44.875 200.495 ;
        RECT 49.765 200.325 49.935 200.515 ;
        RECT 50.225 200.305 50.395 200.495 ;
        RECT 50.740 200.355 50.860 200.465 ;
        RECT 52.525 200.325 52.695 200.515 ;
        RECT 55.745 200.305 55.915 200.495 ;
        RECT 58.045 200.325 58.215 200.515 ;
        RECT 61.265 200.305 61.435 200.495 ;
        RECT 62.645 200.305 62.815 200.495 ;
        RECT 64.485 200.305 64.655 200.495 ;
        RECT 67.245 200.305 67.415 200.495 ;
        RECT 67.705 200.325 67.875 200.515 ;
        RECT 68.220 200.355 68.340 200.465 ;
        RECT 68.625 200.305 68.795 200.495 ;
        RECT 69.140 200.355 69.260 200.465 ;
        RECT 70.005 200.325 70.175 200.515 ;
        RECT 71.385 200.305 71.555 200.495 ;
        RECT 71.900 200.355 72.020 200.465 ;
        RECT 74.605 200.305 74.775 200.495 ;
        RECT 75.525 200.325 75.695 200.515 ;
        RECT 76.500 200.355 76.620 200.465 ;
        RECT 79.205 200.325 79.375 200.515 ;
        RECT 83.805 200.305 83.975 200.495 ;
        RECT 84.725 200.325 84.895 200.515 ;
        RECT 88.405 200.305 88.575 200.495 ;
        RECT 90.245 200.325 90.415 200.515 ;
        RECT 92.545 200.305 92.715 200.495 ;
        RECT 95.765 200.325 95.935 200.515 ;
        RECT 98.065 200.305 98.235 200.495 ;
        RECT 101.285 200.325 101.455 200.515 ;
        RECT 102.260 200.355 102.380 200.465 ;
        RECT 103.585 200.305 103.755 200.495 ;
        RECT 104.045 200.325 104.215 200.515 ;
        RECT 109.105 200.305 109.275 200.495 ;
        RECT 109.565 200.325 109.735 200.515 ;
        RECT 110.485 200.305 110.655 200.495 ;
        RECT 111.000 200.355 111.120 200.465 ;
        RECT 112.785 200.305 112.955 200.495 ;
        RECT 113.245 200.305 113.415 200.495 ;
        RECT 115.085 200.465 115.255 200.515 ;
        RECT 115.085 200.355 115.260 200.465 ;
        RECT 115.085 200.325 115.255 200.355 ;
        RECT 120.605 200.305 120.775 200.515 ;
        RECT 126.125 200.305 126.295 200.515 ;
        RECT 127.505 200.305 127.675 200.515 ;
        RECT 14.665 199.495 16.035 200.305 ;
        RECT 16.965 199.495 20.635 200.305 ;
        RECT 20.645 199.495 26.155 200.305 ;
        RECT 26.165 199.495 31.675 200.305 ;
        RECT 31.685 199.495 37.195 200.305 ;
        RECT 37.215 199.435 37.645 200.220 ;
        RECT 37.665 199.495 39.495 200.305 ;
        RECT 39.505 199.495 45.015 200.305 ;
        RECT 45.025 199.495 50.535 200.305 ;
        RECT 50.545 199.495 56.055 200.305 ;
        RECT 56.065 199.495 61.575 200.305 ;
        RECT 61.595 199.395 62.945 200.305 ;
        RECT 62.975 199.435 63.405 200.220 ;
        RECT 63.435 199.395 64.785 200.305 ;
        RECT 64.805 199.495 67.555 200.305 ;
        RECT 67.565 199.525 68.935 200.305 ;
        RECT 69.405 199.625 71.695 200.305 ;
        RECT 69.405 199.395 70.325 199.625 ;
        RECT 72.165 199.495 74.915 200.305 ;
        RECT 74.925 199.625 84.115 200.305 ;
        RECT 74.925 199.395 75.845 199.625 ;
        RECT 78.675 199.405 79.605 199.625 ;
        RECT 85.045 199.495 88.715 200.305 ;
        RECT 88.735 199.435 89.165 200.220 ;
        RECT 89.185 199.495 92.855 200.305 ;
        RECT 92.865 199.495 98.375 200.305 ;
        RECT 98.385 199.495 103.895 200.305 ;
        RECT 103.905 199.495 109.415 200.305 ;
        RECT 109.435 199.395 110.785 200.305 ;
        RECT 111.265 199.495 113.095 200.305 ;
        RECT 113.115 199.395 114.465 200.305 ;
        RECT 114.495 199.435 114.925 200.220 ;
        RECT 115.405 199.495 120.915 200.305 ;
        RECT 120.925 199.495 126.435 200.305 ;
        RECT 126.445 199.495 127.815 200.305 ;
      LAYER nwell ;
        RECT 14.470 196.275 128.010 199.105 ;
      LAYER pwell ;
        RECT 14.665 195.075 16.035 195.885 ;
        RECT 16.045 195.075 18.795 195.885 ;
        RECT 18.805 195.075 24.315 195.885 ;
        RECT 24.335 195.160 24.765 195.945 ;
        RECT 25.705 195.075 31.215 195.885 ;
        RECT 31.225 195.075 36.735 195.885 ;
        RECT 36.745 195.075 42.255 195.885 ;
        RECT 42.275 195.075 43.625 195.985 ;
        RECT 44.565 195.075 50.075 195.885 ;
        RECT 50.095 195.160 50.525 195.945 ;
        RECT 51.005 195.075 52.835 195.885 ;
        RECT 52.845 195.075 58.355 195.885 ;
        RECT 58.565 195.755 60.775 195.985 ;
        RECT 63.495 195.755 64.425 195.975 ;
        RECT 58.565 195.075 68.935 195.755 ;
        RECT 68.945 195.075 72.055 195.985 ;
        RECT 72.165 195.075 75.835 195.885 ;
        RECT 75.855 195.160 76.285 195.945 ;
        RECT 76.775 195.075 78.125 195.985 ;
        RECT 78.245 195.075 81.355 195.985 ;
        RECT 81.365 195.075 85.035 195.885 ;
        RECT 85.415 195.875 86.335 195.985 ;
        RECT 85.415 195.755 87.750 195.875 ;
        RECT 92.415 195.755 93.335 195.975 ;
        RECT 85.415 195.075 94.695 195.755 ;
        RECT 94.705 195.075 100.215 195.885 ;
        RECT 100.225 195.075 101.595 195.855 ;
        RECT 101.615 195.160 102.045 195.945 ;
        RECT 102.525 195.075 106.195 195.885 ;
        RECT 106.205 195.755 107.125 195.985 ;
        RECT 109.955 195.755 110.885 195.975 ;
        RECT 115.405 195.755 116.325 195.985 ;
        RECT 119.155 195.755 120.085 195.975 ;
        RECT 106.205 195.075 115.395 195.755 ;
        RECT 115.405 195.075 124.595 195.755 ;
        RECT 124.605 195.075 126.435 195.885 ;
        RECT 126.445 195.075 127.815 195.885 ;
        RECT 14.805 194.865 14.975 195.075 ;
        RECT 16.645 194.910 16.805 195.020 ;
        RECT 18.485 194.885 18.655 195.075 ;
        RECT 20.325 194.865 20.495 195.055 ;
        RECT 24.005 194.885 24.175 195.075 ;
        RECT 25.385 194.920 25.545 195.030 ;
        RECT 25.845 194.865 26.015 195.055 ;
        RECT 30.905 194.885 31.075 195.075 ;
        RECT 31.365 194.865 31.535 195.055 ;
        RECT 36.425 194.885 36.595 195.075 ;
        RECT 36.885 194.865 37.055 195.055 ;
        RECT 37.805 194.865 37.975 195.055 ;
        RECT 41.945 194.885 42.115 195.075 ;
        RECT 43.325 194.885 43.495 195.075 ;
        RECT 44.245 194.920 44.405 195.030 ;
        RECT 47.465 194.910 47.625 195.020 ;
        RECT 47.925 194.865 48.095 195.055 ;
        RECT 49.765 194.885 49.935 195.075 ;
        RECT 50.740 194.915 50.860 195.025 ;
        RECT 52.525 194.885 52.695 195.075 ;
        RECT 58.045 194.865 58.215 195.075 ;
        RECT 58.965 194.910 59.125 195.020 ;
        RECT 62.645 194.865 62.815 195.055 ;
        RECT 64.485 194.865 64.655 195.055 ;
        RECT 14.665 194.055 16.035 194.865 ;
        RECT 16.965 194.055 20.635 194.865 ;
        RECT 20.645 194.055 26.155 194.865 ;
        RECT 26.165 194.055 31.675 194.865 ;
        RECT 31.685 194.055 37.195 194.865 ;
        RECT 37.215 193.995 37.645 194.780 ;
        RECT 37.665 194.185 46.855 194.865 ;
        RECT 42.175 193.965 43.105 194.185 ;
        RECT 45.935 193.955 46.855 194.185 ;
        RECT 47.795 193.955 49.145 194.865 ;
        RECT 49.165 194.185 58.355 194.865 ;
        RECT 49.165 193.955 50.085 194.185 ;
        RECT 52.915 193.965 53.845 194.185 ;
        RECT 59.285 194.055 62.955 194.865 ;
        RECT 62.975 193.995 63.405 194.780 ;
        RECT 63.425 194.055 64.795 194.865 ;
        RECT 64.945 194.835 65.115 195.055 ;
        RECT 68.625 194.885 68.795 195.075 ;
        RECT 70.920 194.865 71.090 195.055 ;
        RECT 71.845 194.885 72.015 195.075 ;
        RECT 67.070 194.835 68.015 194.865 ;
        RECT 64.945 194.635 68.015 194.835 ;
        RECT 64.805 194.155 68.015 194.635 ;
        RECT 64.805 193.955 65.735 194.155 ;
        RECT 67.070 193.955 68.015 194.155 ;
        RECT 68.315 193.955 71.235 194.865 ;
        RECT 71.245 194.835 72.190 194.865 ;
        RECT 74.145 194.835 74.315 195.055 ;
        RECT 75.525 194.885 75.695 195.075 ;
        RECT 76.905 195.055 77.075 195.075 ;
        RECT 76.445 195.025 76.615 195.055 ;
        RECT 76.445 194.915 76.620 195.025 ;
        RECT 76.445 194.865 76.615 194.915 ;
        RECT 76.900 194.885 77.075 195.055 ;
        RECT 78.285 194.885 78.455 195.075 ;
        RECT 78.745 194.910 78.905 195.020 ;
        RECT 76.900 194.865 77.070 194.885 ;
        RECT 84.265 194.865 84.435 195.055 ;
        RECT 84.725 194.885 84.895 195.075 ;
        RECT 88.130 194.865 88.300 195.055 ;
        RECT 90.245 194.865 90.415 195.055 ;
        RECT 90.705 194.865 90.875 195.055 ;
        RECT 93.465 194.865 93.635 195.055 ;
        RECT 93.925 194.865 94.095 195.055 ;
        RECT 94.385 194.885 94.555 195.075 ;
        RECT 99.905 194.885 100.075 195.075 ;
        RECT 100.365 194.885 100.535 195.075 ;
        RECT 102.260 194.915 102.380 195.025 ;
        RECT 104.045 194.865 104.215 195.055 ;
        RECT 104.560 194.915 104.680 195.025 ;
        RECT 105.885 194.885 106.055 195.075 ;
        RECT 106.345 194.865 106.515 195.055 ;
        RECT 110.210 194.865 110.380 195.055 ;
        RECT 111.000 194.915 111.120 195.025 ;
        RECT 111.405 194.865 111.575 195.055 ;
        RECT 114.165 194.865 114.335 195.055 ;
        RECT 115.085 195.025 115.255 195.075 ;
        RECT 115.085 194.915 115.260 195.025 ;
        RECT 115.085 194.885 115.255 194.915 ;
        RECT 115.545 194.865 115.715 195.055 ;
        RECT 116.980 194.915 117.100 195.025 ;
        RECT 120.605 194.865 120.775 195.055 ;
        RECT 124.285 194.885 124.455 195.075 ;
        RECT 126.125 194.865 126.295 195.075 ;
        RECT 127.505 194.865 127.675 195.075 ;
        RECT 71.245 194.635 74.315 194.835 ;
        RECT 71.245 194.155 74.455 194.635 ;
        RECT 71.245 193.955 72.190 194.155 ;
        RECT 73.525 193.955 74.455 194.155 ;
        RECT 74.465 194.185 76.755 194.865 ;
        RECT 74.465 193.955 75.385 194.185 ;
        RECT 76.785 193.955 78.135 194.865 ;
        RECT 79.065 194.055 84.575 194.865 ;
        RECT 84.815 194.185 88.715 194.865 ;
        RECT 87.785 193.955 88.715 194.185 ;
        RECT 88.735 193.995 89.165 194.780 ;
        RECT 89.185 194.055 90.555 194.865 ;
        RECT 90.565 194.085 91.935 194.865 ;
        RECT 91.945 194.055 93.775 194.865 ;
        RECT 93.795 193.955 95.145 194.865 ;
        RECT 95.165 194.185 104.355 194.865 ;
        RECT 95.165 193.955 96.085 194.185 ;
        RECT 98.915 193.965 99.845 194.185 ;
        RECT 104.825 194.055 106.655 194.865 ;
        RECT 106.895 194.185 110.795 194.865 ;
        RECT 109.865 193.955 110.795 194.185 ;
        RECT 111.265 194.085 112.635 194.865 ;
        RECT 112.645 194.055 114.475 194.865 ;
        RECT 114.495 193.995 114.925 194.780 ;
        RECT 115.405 194.085 116.775 194.865 ;
        RECT 117.245 194.055 120.915 194.865 ;
        RECT 120.925 194.055 126.435 194.865 ;
        RECT 126.445 194.055 127.815 194.865 ;
      LAYER nwell ;
        RECT 14.470 190.835 128.010 193.665 ;
      LAYER pwell ;
        RECT 14.665 189.635 16.035 190.445 ;
        RECT 16.045 189.635 18.795 190.445 ;
        RECT 18.805 189.635 24.315 190.445 ;
        RECT 24.335 189.720 24.765 190.505 ;
        RECT 25.245 189.635 30.755 190.445 ;
        RECT 30.775 189.635 32.125 190.545 ;
        RECT 35.345 190.315 36.275 190.545 ;
        RECT 32.375 189.635 36.275 190.315 ;
        RECT 36.285 189.635 37.655 190.445 ;
        RECT 40.865 190.315 41.795 190.545 ;
        RECT 37.895 189.635 41.795 190.315 ;
        RECT 42.265 189.635 43.635 190.415 ;
        RECT 44.115 189.635 45.465 190.545 ;
        RECT 45.485 189.635 48.235 190.445 ;
        RECT 48.245 189.635 49.615 190.415 ;
        RECT 50.095 189.720 50.525 190.505 ;
        RECT 53.745 190.315 54.675 190.545 ;
        RECT 50.775 189.635 54.675 190.315 ;
        RECT 54.685 189.635 56.055 190.415 ;
        RECT 56.985 189.635 62.495 190.445 ;
        RECT 62.505 189.635 68.015 190.445 ;
        RECT 68.025 190.315 69.370 190.545 ;
        RECT 68.025 189.635 69.855 190.315 ;
        RECT 69.865 189.635 72.155 190.545 ;
        RECT 73.675 190.315 74.605 190.545 ;
        RECT 72.770 189.635 74.605 190.315 ;
        RECT 75.855 189.720 76.285 190.505 ;
        RECT 76.765 189.635 78.595 190.445 ;
        RECT 78.605 189.635 84.115 190.445 ;
        RECT 84.495 190.435 85.415 190.545 ;
        RECT 84.495 190.315 86.830 190.435 ;
        RECT 91.495 190.315 92.415 190.535 ;
        RECT 84.495 189.635 93.775 190.315 ;
        RECT 93.785 189.635 95.615 190.445 ;
        RECT 98.825 190.315 99.755 190.545 ;
        RECT 95.855 189.635 99.755 190.315 ;
        RECT 99.765 189.635 101.595 190.445 ;
        RECT 101.615 189.720 102.045 190.505 ;
        RECT 102.525 189.635 104.355 190.445 ;
        RECT 104.365 189.635 109.875 190.445 ;
        RECT 113.085 190.315 114.015 190.545 ;
        RECT 110.115 189.635 114.015 190.315 ;
        RECT 114.025 189.635 115.395 190.445 ;
        RECT 115.405 189.635 120.915 190.445 ;
        RECT 120.925 189.635 126.435 190.445 ;
        RECT 126.445 189.635 127.815 190.445 ;
        RECT 14.805 189.425 14.975 189.635 ;
        RECT 16.645 189.470 16.805 189.580 ;
        RECT 18.485 189.445 18.655 189.635 ;
        RECT 20.325 189.425 20.495 189.615 ;
        RECT 24.005 189.445 24.175 189.635 ;
        RECT 24.980 189.475 25.100 189.585 ;
        RECT 25.845 189.425 26.015 189.615 ;
        RECT 26.305 189.425 26.475 189.615 ;
        RECT 30.445 189.445 30.615 189.635 ;
        RECT 30.905 189.445 31.075 189.635 ;
        RECT 35.690 189.445 35.860 189.635 ;
        RECT 36.885 189.425 37.055 189.615 ;
        RECT 37.345 189.445 37.515 189.635 ;
        RECT 38.725 189.425 38.895 189.615 ;
        RECT 39.645 189.470 39.805 189.580 ;
        RECT 41.210 189.445 41.380 189.635 ;
        RECT 42.000 189.475 42.120 189.585 ;
        RECT 43.325 189.445 43.495 189.635 ;
        RECT 43.840 189.475 43.960 189.585 ;
        RECT 45.165 189.445 45.335 189.635 ;
        RECT 47.925 189.445 48.095 189.635 ;
        RECT 48.845 189.425 49.015 189.615 ;
        RECT 49.305 189.445 49.475 189.635 ;
        RECT 49.820 189.475 49.940 189.585 ;
        RECT 54.090 189.445 54.260 189.635 ;
        RECT 54.825 189.445 54.995 189.635 ;
        RECT 56.665 189.480 56.825 189.590 ;
        RECT 58.045 189.425 58.215 189.615 ;
        RECT 58.965 189.470 59.125 189.580 ;
        RECT 62.185 189.445 62.355 189.635 ;
        RECT 62.645 189.425 62.815 189.615 ;
        RECT 66.785 189.425 66.955 189.615 ;
        RECT 67.705 189.445 67.875 189.635 ;
        RECT 69.545 189.445 69.715 189.635 ;
        RECT 71.840 189.445 72.010 189.635 ;
        RECT 72.770 189.615 72.935 189.635 ;
        RECT 72.305 189.585 72.475 189.615 ;
        RECT 72.305 189.475 72.480 189.585 ;
        RECT 72.305 189.425 72.475 189.475 ;
        RECT 72.765 189.445 72.935 189.615 ;
        RECT 73.685 189.425 73.855 189.615 ;
        RECT 75.525 189.425 75.695 189.615 ;
        RECT 76.500 189.475 76.620 189.585 ;
        RECT 76.905 189.425 77.075 189.615 ;
        RECT 77.420 189.475 77.540 189.585 ;
        RECT 78.285 189.445 78.455 189.635 ;
        RECT 80.125 189.425 80.295 189.615 ;
        RECT 83.805 189.445 83.975 189.635 ;
        RECT 85.645 189.425 85.815 189.615 ;
        RECT 86.105 189.425 86.275 189.615 ;
        RECT 87.485 189.425 87.655 189.615 ;
        RECT 89.380 189.475 89.500 189.585 ;
        RECT 89.785 189.425 89.955 189.615 ;
        RECT 91.220 189.475 91.340 189.585 ;
        RECT 93.465 189.445 93.635 189.635 ;
        RECT 95.305 189.445 95.475 189.635 ;
        RECT 96.685 189.425 96.855 189.615 ;
        RECT 97.145 189.425 97.315 189.615 ;
        RECT 99.170 189.445 99.340 189.635 ;
        RECT 101.285 189.445 101.455 189.635 ;
        RECT 102.260 189.475 102.380 189.585 ;
        RECT 104.045 189.445 104.215 189.635 ;
        RECT 107.265 189.425 107.435 189.615 ;
        RECT 108.645 189.425 108.815 189.615 ;
        RECT 109.565 189.445 109.735 189.635 ;
        RECT 113.430 189.445 113.600 189.635 ;
        RECT 114.165 189.425 114.335 189.615 ;
        RECT 115.085 189.585 115.255 189.635 ;
        RECT 115.085 189.475 115.260 189.585 ;
        RECT 115.085 189.445 115.255 189.475 ;
        RECT 120.605 189.445 120.775 189.635 ;
        RECT 124.285 189.425 124.455 189.615 ;
        RECT 126.125 189.425 126.295 189.635 ;
        RECT 127.505 189.425 127.675 189.635 ;
        RECT 14.665 188.615 16.035 189.425 ;
        RECT 16.965 188.615 20.635 189.425 ;
        RECT 20.645 188.615 26.155 189.425 ;
        RECT 26.175 188.515 27.525 189.425 ;
        RECT 27.915 188.745 37.195 189.425 ;
        RECT 27.915 188.625 30.250 188.745 ;
        RECT 27.915 188.515 28.835 188.625 ;
        RECT 34.915 188.525 35.835 188.745 ;
        RECT 37.215 188.555 37.645 189.340 ;
        RECT 37.665 188.645 39.035 189.425 ;
        RECT 39.965 188.745 49.155 189.425 ;
        RECT 49.165 188.745 58.355 189.425 ;
        RECT 39.965 188.515 40.885 188.745 ;
        RECT 43.715 188.525 44.645 188.745 ;
        RECT 49.165 188.515 50.085 188.745 ;
        RECT 52.915 188.525 53.845 188.745 ;
        RECT 59.285 188.615 62.955 189.425 ;
        RECT 62.975 188.555 63.405 189.340 ;
        RECT 63.425 188.615 67.095 189.425 ;
        RECT 67.105 188.615 72.615 189.425 ;
        RECT 72.635 188.515 73.985 189.425 ;
        RECT 74.005 188.615 75.835 189.425 ;
        RECT 75.845 188.645 77.215 189.425 ;
        RECT 77.685 188.615 80.435 189.425 ;
        RECT 80.445 188.615 85.955 189.425 ;
        RECT 85.975 188.515 87.325 189.425 ;
        RECT 87.355 188.515 88.705 189.425 ;
        RECT 88.735 188.555 89.165 189.340 ;
        RECT 89.645 188.645 91.015 189.425 ;
        RECT 91.485 188.615 96.995 189.425 ;
        RECT 97.015 188.515 98.365 189.425 ;
        RECT 98.385 188.745 107.575 189.425 ;
        RECT 98.385 188.515 99.305 188.745 ;
        RECT 102.135 188.525 103.065 188.745 ;
        RECT 107.585 188.615 108.955 189.425 ;
        RECT 108.965 188.615 114.475 189.425 ;
        RECT 114.495 188.555 114.925 189.340 ;
        RECT 115.405 188.745 124.595 189.425 ;
        RECT 115.405 188.515 116.325 188.745 ;
        RECT 119.155 188.525 120.085 188.745 ;
        RECT 124.605 188.615 126.435 189.425 ;
        RECT 126.445 188.615 127.815 189.425 ;
      LAYER nwell ;
        RECT 14.470 185.395 128.010 188.225 ;
      LAYER pwell ;
        RECT 14.665 184.195 16.035 185.005 ;
        RECT 16.045 184.195 18.795 185.005 ;
        RECT 18.805 184.195 24.315 185.005 ;
        RECT 24.335 184.280 24.765 185.065 ;
        RECT 29.295 184.875 30.225 185.095 ;
        RECT 33.055 184.875 33.975 185.105 ;
        RECT 24.785 184.195 33.975 184.875 ;
        RECT 34.905 184.195 40.415 185.005 ;
        RECT 40.425 184.195 45.935 185.005 ;
        RECT 49.145 184.875 50.075 185.105 ;
        RECT 46.175 184.195 50.075 184.875 ;
        RECT 50.095 184.280 50.525 185.065 ;
        RECT 51.475 184.195 52.825 185.105 ;
        RECT 52.845 184.195 55.595 185.005 ;
        RECT 55.605 184.195 56.975 184.975 ;
        RECT 56.995 184.195 58.345 185.105 ;
        RECT 58.365 184.195 61.115 185.005 ;
        RECT 61.125 184.195 66.635 185.005 ;
        RECT 66.645 184.875 67.565 185.105 ;
        RECT 70.395 184.875 71.325 185.095 ;
        RECT 66.645 184.195 75.835 184.875 ;
        RECT 75.855 184.280 76.285 185.065 ;
        RECT 76.315 184.195 77.665 185.105 ;
        RECT 78.145 184.195 79.975 185.005 ;
        RECT 79.985 184.195 85.495 185.005 ;
        RECT 88.705 184.875 89.635 185.105 ;
        RECT 85.735 184.195 89.635 184.875 ;
        RECT 90.565 184.195 96.075 185.005 ;
        RECT 96.085 184.195 101.595 185.005 ;
        RECT 101.615 184.280 102.045 185.065 ;
        RECT 105.725 184.875 106.655 185.105 ;
        RECT 102.755 184.195 106.655 184.875 ;
        RECT 106.665 184.195 108.035 184.975 ;
        RECT 108.045 184.195 109.415 185.005 ;
        RECT 109.435 184.195 110.785 185.105 ;
        RECT 110.805 184.875 111.725 185.105 ;
        RECT 114.555 184.875 115.485 185.095 ;
        RECT 110.805 184.195 119.995 184.875 ;
        RECT 120.015 184.195 121.365 185.105 ;
        RECT 121.385 184.195 122.755 184.975 ;
        RECT 122.765 184.195 126.435 185.005 ;
        RECT 126.445 184.195 127.815 185.005 ;
        RECT 14.805 183.985 14.975 184.195 ;
        RECT 16.240 184.035 16.360 184.145 ;
        RECT 18.485 184.005 18.655 184.195 ;
        RECT 21.705 183.985 21.875 184.175 ;
        RECT 24.005 184.005 24.175 184.195 ;
        RECT 24.925 184.005 25.095 184.195 ;
        RECT 27.225 183.985 27.395 184.175 ;
        RECT 28.605 183.985 28.775 184.175 ;
        RECT 29.340 183.985 29.510 184.175 ;
        RECT 33.260 184.035 33.380 184.145 ;
        RECT 34.585 184.040 34.745 184.150 ;
        RECT 36.885 183.985 37.055 184.175 ;
        RECT 37.860 184.035 37.980 184.145 ;
        RECT 40.105 184.005 40.275 184.195 ;
        RECT 41.485 183.985 41.655 184.175 ;
        RECT 45.350 183.985 45.520 184.175 ;
        RECT 45.625 184.005 45.795 184.195 ;
        RECT 46.090 183.985 46.260 184.175 ;
        RECT 49.490 184.005 49.660 184.195 ;
        RECT 51.145 184.040 51.305 184.150 ;
        RECT 51.605 184.005 51.775 184.195 ;
        RECT 53.170 183.985 53.340 184.175 ;
        RECT 55.285 184.005 55.455 184.195 ;
        RECT 55.745 184.005 55.915 184.195 ;
        RECT 58.045 184.005 58.215 184.195 ;
        RECT 60.805 184.005 60.975 184.195 ;
        RECT 62.645 183.985 62.815 184.175 ;
        RECT 63.565 183.985 63.735 184.175 ;
        RECT 65.405 183.985 65.575 184.175 ;
        RECT 66.325 184.005 66.495 184.195 ;
        RECT 75.525 184.005 75.695 184.195 ;
        RECT 77.365 184.005 77.535 184.195 ;
        RECT 77.880 184.035 78.000 184.145 ;
        RECT 78.745 183.985 78.915 184.175 ;
        RECT 79.665 184.005 79.835 184.195 ;
        RECT 84.265 183.985 84.435 184.175 ;
        RECT 85.185 184.005 85.355 184.195 ;
        RECT 88.130 183.985 88.300 184.175 ;
        RECT 89.050 184.005 89.220 184.195 ;
        RECT 90.245 183.985 90.415 184.175 ;
        RECT 90.705 183.985 90.875 184.175 ;
        RECT 93.005 183.985 93.175 184.175 ;
        RECT 95.765 184.005 95.935 184.195 ;
        RECT 101.285 184.005 101.455 184.195 ;
        RECT 102.205 184.145 102.375 184.175 ;
        RECT 102.205 184.035 102.380 184.145 ;
        RECT 102.720 184.035 102.840 184.145 ;
        RECT 102.205 183.985 102.375 184.035 ;
        RECT 104.505 183.985 104.675 184.175 ;
        RECT 106.070 184.005 106.240 184.195 ;
        RECT 107.725 184.005 107.895 184.195 ;
        RECT 109.105 184.005 109.275 184.195 ;
        RECT 109.565 184.005 109.735 184.195 ;
        RECT 110.025 183.985 110.195 184.175 ;
        RECT 113.890 183.985 114.060 184.175 ;
        RECT 115.545 184.030 115.705 184.140 ;
        RECT 116.005 183.985 116.175 184.175 ;
        RECT 119.685 184.005 119.855 184.195 ;
        RECT 120.145 184.005 120.315 184.195 ;
        RECT 120.605 183.985 120.775 184.175 ;
        RECT 121.525 184.005 121.695 184.195 ;
        RECT 126.125 183.985 126.295 184.195 ;
        RECT 127.505 183.985 127.675 184.195 ;
        RECT 14.665 183.175 16.035 183.985 ;
        RECT 16.505 183.175 22.015 183.985 ;
        RECT 22.025 183.175 27.535 183.985 ;
        RECT 27.545 183.205 28.915 183.985 ;
        RECT 28.925 183.305 32.825 183.985 ;
        RECT 28.925 183.075 29.855 183.305 ;
        RECT 33.525 183.175 37.195 183.985 ;
        RECT 37.215 183.115 37.645 183.900 ;
        RECT 38.125 183.175 41.795 183.985 ;
        RECT 42.035 183.305 45.935 183.985 ;
        RECT 45.005 183.075 45.935 183.305 ;
        RECT 45.945 183.075 49.420 183.985 ;
        RECT 49.855 183.305 53.755 183.985 ;
        RECT 52.825 183.075 53.755 183.305 ;
        RECT 53.765 183.305 62.955 183.985 ;
        RECT 53.765 183.075 54.685 183.305 ;
        RECT 57.515 183.085 58.445 183.305 ;
        RECT 62.975 183.115 63.405 183.900 ;
        RECT 63.425 183.305 65.255 183.985 ;
        RECT 65.265 183.755 66.835 183.985 ;
        RECT 68.925 183.945 69.845 183.985 ;
        RECT 68.925 183.755 69.855 183.945 ;
        RECT 65.265 183.395 69.855 183.755 ;
        RECT 65.265 183.305 69.845 183.395 ;
        RECT 66.845 183.075 69.845 183.305 ;
        RECT 69.865 183.305 79.055 183.985 ;
        RECT 69.865 183.075 70.785 183.305 ;
        RECT 73.615 183.085 74.545 183.305 ;
        RECT 79.065 183.175 84.575 183.985 ;
        RECT 84.815 183.305 88.715 183.985 ;
        RECT 87.785 183.075 88.715 183.305 ;
        RECT 88.735 183.115 89.165 183.900 ;
        RECT 89.185 183.175 90.555 183.985 ;
        RECT 90.565 183.205 91.935 183.985 ;
        RECT 91.945 183.175 93.315 183.985 ;
        RECT 93.325 183.305 102.515 183.985 ;
        RECT 93.325 183.075 94.245 183.305 ;
        RECT 97.075 183.085 98.005 183.305 ;
        RECT 102.985 183.175 104.815 183.985 ;
        RECT 104.825 183.175 110.335 183.985 ;
        RECT 110.575 183.305 114.475 183.985 ;
        RECT 113.545 183.075 114.475 183.305 ;
        RECT 114.495 183.115 114.925 183.900 ;
        RECT 115.865 183.205 117.235 183.985 ;
        RECT 117.245 183.175 120.915 183.985 ;
        RECT 120.925 183.175 126.435 183.985 ;
        RECT 126.445 183.175 127.815 183.985 ;
      LAYER nwell ;
        RECT 14.470 179.955 128.010 182.785 ;
      LAYER pwell ;
        RECT 14.665 178.755 16.035 179.565 ;
        RECT 16.045 178.755 18.795 179.565 ;
        RECT 18.805 178.755 24.315 179.565 ;
        RECT 24.335 178.840 24.765 179.625 ;
        RECT 25.245 178.755 30.755 179.565 ;
        RECT 30.765 178.755 36.275 179.565 ;
        RECT 36.295 178.755 37.645 179.665 ;
        RECT 37.665 179.435 38.585 179.665 ;
        RECT 41.415 179.435 42.345 179.655 ;
        RECT 37.665 178.755 46.855 179.435 ;
        RECT 46.865 178.755 48.235 179.535 ;
        RECT 48.245 178.755 50.075 179.565 ;
        RECT 50.095 178.840 50.525 179.625 ;
        RECT 51.005 178.755 53.755 179.565 ;
        RECT 56.965 179.435 57.895 179.665 ;
        RECT 53.995 178.755 57.895 179.435 ;
        RECT 58.825 178.755 60.195 179.535 ;
        RECT 60.205 178.755 62.035 179.565 ;
        RECT 62.045 178.755 67.555 179.565 ;
        RECT 67.565 179.435 68.910 179.665 ;
        RECT 69.405 179.435 70.335 179.665 ;
        RECT 67.565 178.755 69.395 179.435 ;
        RECT 69.405 178.755 73.075 179.435 ;
        RECT 73.085 178.755 74.455 179.565 ;
        RECT 74.475 178.755 75.825 179.665 ;
        RECT 75.855 178.840 76.285 179.625 ;
        RECT 77.225 178.755 80.895 179.565 ;
        RECT 80.905 178.755 83.515 179.665 ;
        RECT 84.585 179.435 85.505 179.665 ;
        RECT 88.335 179.435 89.265 179.655 ;
        RECT 84.585 178.755 93.775 179.435 ;
        RECT 94.715 178.755 96.065 179.665 ;
        RECT 99.285 179.435 100.215 179.665 ;
        RECT 96.315 178.755 100.215 179.435 ;
        RECT 100.225 178.755 101.595 179.535 ;
        RECT 101.615 178.840 102.045 179.625 ;
        RECT 102.065 178.755 103.435 179.565 ;
        RECT 103.445 178.755 107.115 179.565 ;
        RECT 107.125 178.755 110.600 179.665 ;
        RECT 110.805 178.755 112.175 179.565 ;
        RECT 115.385 179.435 116.315 179.665 ;
        RECT 112.415 178.755 116.315 179.435 ;
        RECT 116.325 178.755 118.155 179.565 ;
        RECT 118.175 178.755 119.525 179.665 ;
        RECT 119.545 178.755 120.915 179.565 ;
        RECT 120.925 178.755 126.435 179.565 ;
        RECT 126.445 178.755 127.815 179.565 ;
        RECT 14.805 178.545 14.975 178.755 ;
        RECT 16.645 178.590 16.805 178.700 ;
        RECT 18.485 178.565 18.655 178.755 ;
        RECT 22.165 178.545 22.335 178.735 ;
        RECT 22.625 178.545 22.795 178.735 ;
        RECT 24.005 178.565 24.175 178.755 ;
        RECT 24.980 178.595 25.100 178.705 ;
        RECT 30.445 178.565 30.615 178.755 ;
        RECT 31.880 178.595 32.000 178.705 ;
        RECT 33.205 178.545 33.375 178.735 ;
        RECT 35.965 178.565 36.135 178.755 ;
        RECT 36.425 178.565 36.595 178.755 ;
        RECT 36.880 178.545 37.050 178.735 ;
        RECT 37.860 178.595 37.980 178.705 ;
        RECT 41.485 178.545 41.655 178.735 ;
        RECT 45.160 178.545 45.330 178.735 ;
        RECT 45.625 178.545 45.795 178.735 ;
        RECT 46.545 178.565 46.715 178.755 ;
        RECT 47.925 178.565 48.095 178.755 ;
        RECT 49.765 178.565 49.935 178.755 ;
        RECT 50.740 178.595 50.860 178.705 ;
        RECT 53.445 178.565 53.615 178.755 ;
        RECT 57.125 178.545 57.295 178.735 ;
        RECT 57.310 178.565 57.480 178.755 ;
        RECT 58.505 178.600 58.665 178.710 ;
        RECT 58.965 178.565 59.135 178.755 ;
        RECT 61.725 178.565 61.895 178.755 ;
        RECT 62.645 178.545 62.815 178.735 ;
        RECT 64.945 178.545 65.115 178.735 ;
        RECT 65.405 178.545 65.575 178.735 ;
        RECT 67.245 178.565 67.415 178.755 ;
        RECT 68.625 178.545 68.795 178.735 ;
        RECT 69.085 178.565 69.255 178.755 ;
        RECT 72.765 178.565 72.935 178.755 ;
        RECT 74.145 178.545 74.315 178.755 ;
        RECT 74.605 178.545 74.775 178.755 ;
        RECT 80.585 178.735 80.755 178.755 ;
        RECT 76.905 178.600 77.065 178.710 ;
        RECT 80.580 178.565 80.755 178.735 ;
        RECT 80.580 178.545 80.750 178.565 ;
        RECT 81.050 178.545 81.220 178.755 ;
        RECT 84.265 178.600 84.425 178.710 ;
        RECT 84.730 178.545 84.900 178.735 ;
        RECT 88.405 178.545 88.575 178.735 ;
        RECT 93.465 178.565 93.635 178.755 ;
        RECT 94.385 178.545 94.555 178.735 ;
        RECT 94.845 178.565 95.015 178.755 ;
        RECT 99.630 178.565 99.800 178.755 ;
        RECT 99.905 178.545 100.075 178.735 ;
        RECT 100.365 178.565 100.535 178.755 ;
        RECT 103.125 178.565 103.295 178.755 ;
        RECT 103.580 178.545 103.750 178.735 ;
        RECT 104.050 178.545 104.220 178.735 ;
        RECT 106.805 178.565 106.975 178.755 ;
        RECT 107.270 178.565 107.440 178.755 ;
        RECT 107.730 178.545 107.900 178.735 ;
        RECT 111.460 178.595 111.580 178.705 ;
        RECT 111.865 178.565 112.035 178.755 ;
        RECT 114.165 178.545 114.335 178.735 ;
        RECT 115.140 178.595 115.260 178.705 ;
        RECT 115.730 178.565 115.900 178.755 ;
        RECT 117.845 178.565 118.015 178.755 ;
        RECT 119.225 178.565 119.395 178.755 ;
        RECT 120.605 178.565 120.775 178.755 ;
        RECT 124.285 178.545 124.455 178.735 ;
        RECT 126.125 178.545 126.295 178.755 ;
        RECT 127.505 178.545 127.675 178.755 ;
        RECT 14.665 177.735 16.035 178.545 ;
        RECT 16.965 177.735 22.475 178.545 ;
        RECT 22.485 177.865 31.675 178.545 ;
        RECT 26.995 177.645 27.925 177.865 ;
        RECT 30.755 177.635 31.675 177.865 ;
        RECT 32.145 177.765 33.515 178.545 ;
        RECT 33.720 177.635 37.195 178.545 ;
        RECT 37.215 177.675 37.645 178.460 ;
        RECT 38.125 177.735 41.795 178.545 ;
        RECT 42.000 177.635 45.475 178.545 ;
        RECT 45.485 177.865 54.590 178.545 ;
        RECT 54.685 177.735 57.435 178.545 ;
        RECT 57.445 177.735 62.955 178.545 ;
        RECT 62.975 177.675 63.405 178.460 ;
        RECT 63.425 177.865 65.255 178.545 ;
        RECT 65.265 177.865 67.095 178.545 ;
        RECT 63.425 177.635 64.770 177.865 ;
        RECT 65.750 177.635 67.095 177.865 ;
        RECT 67.105 177.735 68.935 178.545 ;
        RECT 68.945 177.735 74.455 178.545 ;
        RECT 74.465 177.865 77.205 178.545 ;
        RECT 77.420 177.635 80.895 178.545 ;
        RECT 80.905 177.635 84.380 178.545 ;
        RECT 84.585 177.635 87.195 178.545 ;
        RECT 87.355 177.635 88.705 178.545 ;
        RECT 88.735 177.675 89.165 178.460 ;
        RECT 89.185 177.735 94.695 178.545 ;
        RECT 94.705 177.735 100.215 178.545 ;
        RECT 100.420 177.635 103.895 178.545 ;
        RECT 103.905 177.635 107.380 178.545 ;
        RECT 107.585 177.635 111.060 178.545 ;
        RECT 111.725 177.735 114.475 178.545 ;
        RECT 114.495 177.675 114.925 178.460 ;
        RECT 115.405 177.865 124.595 178.545 ;
        RECT 115.405 177.635 116.325 177.865 ;
        RECT 119.155 177.645 120.085 177.865 ;
        RECT 124.605 177.735 126.435 178.545 ;
        RECT 126.445 177.735 127.815 178.545 ;
      LAYER nwell ;
        RECT 14.470 174.515 128.010 177.345 ;
      LAYER pwell ;
        RECT 14.665 173.315 16.035 174.125 ;
        RECT 16.045 173.315 21.555 174.125 ;
        RECT 21.575 173.315 22.925 174.225 ;
        RECT 22.955 173.315 24.305 174.225 ;
        RECT 24.335 173.400 24.765 174.185 ;
        RECT 25.705 173.315 27.075 174.095 ;
        RECT 31.595 173.995 32.525 174.215 ;
        RECT 35.355 173.995 36.275 174.225 ;
        RECT 27.085 173.315 36.275 173.995 ;
        RECT 36.285 173.995 37.215 174.225 ;
        RECT 36.285 173.315 40.185 173.995 ;
        RECT 40.885 173.315 42.715 174.125 ;
        RECT 42.725 173.315 46.200 174.225 ;
        RECT 46.600 173.315 50.075 174.225 ;
        RECT 50.095 173.400 50.525 174.185 ;
        RECT 51.465 173.315 54.940 174.225 ;
        RECT 55.145 173.315 56.515 174.125 ;
        RECT 56.535 173.315 59.275 173.995 ;
        RECT 59.285 173.315 62.035 174.125 ;
        RECT 62.045 173.995 63.390 174.225 ;
        RECT 62.045 173.315 63.875 173.995 ;
        RECT 64.125 173.545 66.880 174.225 ;
        RECT 67.345 173.545 70.100 174.225 ;
        RECT 70.565 173.545 73.320 174.225 ;
        RECT 64.125 173.315 66.395 173.545 ;
        RECT 67.345 173.315 69.615 173.545 ;
        RECT 70.565 173.315 72.835 173.545 ;
        RECT 74.005 173.315 75.835 174.125 ;
        RECT 75.855 173.400 76.285 174.185 ;
        RECT 77.420 173.315 80.895 174.225 ;
        RECT 81.365 173.315 84.115 174.125 ;
        RECT 84.210 173.315 93.315 173.995 ;
        RECT 94.245 173.315 97.915 174.125 ;
        RECT 97.925 173.315 101.400 174.225 ;
        RECT 101.615 173.400 102.045 174.185 ;
        RECT 102.525 173.315 104.355 174.125 ;
        RECT 104.375 173.315 107.115 173.995 ;
        RECT 107.125 173.315 110.600 174.225 ;
        RECT 110.805 173.315 112.635 174.125 ;
        RECT 112.645 173.315 118.155 174.125 ;
        RECT 118.175 173.315 119.525 174.225 ;
        RECT 120.005 173.315 121.375 174.095 ;
        RECT 121.385 173.315 122.755 174.125 ;
        RECT 122.765 173.315 126.435 174.125 ;
        RECT 126.445 173.315 127.815 174.125 ;
        RECT 14.805 173.105 14.975 173.315 ;
        RECT 17.105 173.105 17.275 173.295 ;
        RECT 20.785 173.105 20.955 173.295 ;
        RECT 21.245 173.125 21.415 173.315 ;
        RECT 22.625 173.125 22.795 173.315 ;
        RECT 23.085 173.125 23.255 173.315 ;
        RECT 25.385 173.160 25.545 173.270 ;
        RECT 26.765 173.125 26.935 173.315 ;
        RECT 27.225 173.125 27.395 173.315 ;
        RECT 31.820 173.105 31.990 173.295 ;
        RECT 32.560 173.105 32.730 173.295 ;
        RECT 36.700 173.125 36.870 173.315 ;
        RECT 36.885 173.150 37.045 173.260 ;
        RECT 37.810 173.105 37.980 173.295 ;
        RECT 40.620 173.155 40.740 173.265 ;
        RECT 41.540 173.155 41.660 173.265 ;
        RECT 41.950 173.105 42.120 173.295 ;
        RECT 42.405 173.125 42.575 173.315 ;
        RECT 42.870 173.125 43.040 173.315 ;
        RECT 45.630 173.105 45.800 173.295 ;
        RECT 49.760 173.125 49.930 173.315 ;
        RECT 51.145 173.160 51.305 173.270 ;
        RECT 51.610 173.125 51.780 173.315 ;
        RECT 52.525 173.105 52.695 173.295 ;
        RECT 54.365 173.125 54.535 173.295 ;
        RECT 56.205 173.125 56.375 173.315 ;
        RECT 57.125 173.105 57.295 173.295 ;
        RECT 58.965 173.125 59.135 173.315 ;
        RECT 61.725 173.125 61.895 173.315 ;
        RECT 62.645 173.105 62.815 173.295 ;
        RECT 63.565 173.125 63.735 173.315 ;
        RECT 64.125 173.295 64.195 173.315 ;
        RECT 67.345 173.295 67.415 173.315 ;
        RECT 70.565 173.295 70.635 173.315 ;
        RECT 64.025 173.125 64.195 173.295 ;
        RECT 65.865 173.105 66.035 173.295 ;
        RECT 67.245 173.125 67.415 173.295 ;
        RECT 70.465 173.105 70.635 173.295 ;
        RECT 73.740 173.155 73.860 173.265 ;
        RECT 75.065 173.105 75.235 173.295 ;
        RECT 75.525 173.105 75.695 173.315 ;
        RECT 76.905 173.160 77.065 173.270 ;
        RECT 77.825 173.150 77.985 173.260 ;
        RECT 80.580 173.125 80.750 173.315 ;
        RECT 81.100 173.155 81.220 173.265 ;
        RECT 81.505 173.105 81.675 173.295 ;
        RECT 81.970 173.105 82.140 173.295 ;
        RECT 83.805 173.125 83.975 173.315 ;
        RECT 85.700 173.155 85.820 173.265 ;
        RECT 88.405 173.105 88.575 173.295 ;
        RECT 89.380 173.155 89.500 173.265 ;
        RECT 91.165 173.105 91.335 173.295 ;
        RECT 93.005 173.125 93.175 173.315 ;
        RECT 93.925 173.160 94.085 173.270 ;
        RECT 95.765 173.105 95.935 173.295 ;
        RECT 96.225 173.105 96.395 173.295 ;
        RECT 97.605 173.265 97.775 173.315 ;
        RECT 97.605 173.155 97.780 173.265 ;
        RECT 97.605 173.125 97.775 173.155 ;
        RECT 98.070 173.125 98.240 173.315 ;
        RECT 100.365 173.105 100.535 173.295 ;
        RECT 102.260 173.155 102.380 173.265 ;
        RECT 104.045 173.125 104.215 173.315 ;
        RECT 106.805 173.125 106.975 173.315 ;
        RECT 107.270 173.125 107.440 173.315 ;
        RECT 109.565 173.105 109.735 173.295 ;
        RECT 110.080 173.155 110.200 173.265 ;
        RECT 112.325 173.125 112.495 173.315 ;
        RECT 113.890 173.105 114.060 173.295 ;
        RECT 115.545 173.150 115.705 173.260 ;
        RECT 117.845 173.125 118.015 173.315 ;
        RECT 118.305 173.125 118.475 173.315 ;
        RECT 119.740 173.155 119.860 173.265 ;
        RECT 120.145 173.125 120.315 173.315 ;
        RECT 122.445 173.125 122.615 173.315 ;
        RECT 124.745 173.105 124.915 173.295 ;
        RECT 126.125 173.105 126.295 173.315 ;
        RECT 127.505 173.105 127.675 173.315 ;
        RECT 14.665 172.295 16.035 173.105 ;
        RECT 16.045 172.295 17.415 173.105 ;
        RECT 17.425 172.295 21.095 173.105 ;
        RECT 21.125 172.195 32.135 173.105 ;
        RECT 32.145 172.425 36.045 173.105 ;
        RECT 32.145 172.195 33.075 172.425 ;
        RECT 37.215 172.235 37.645 173.020 ;
        RECT 37.665 172.195 41.140 173.105 ;
        RECT 41.805 172.195 45.280 173.105 ;
        RECT 45.485 172.195 48.960 173.105 ;
        RECT 49.165 172.295 52.835 173.105 ;
        RECT 52.845 172.425 54.210 173.105 ;
        RECT 54.685 172.295 57.435 173.105 ;
        RECT 57.445 172.295 62.955 173.105 ;
        RECT 62.975 172.235 63.405 173.020 ;
        RECT 64.345 172.425 66.175 173.105 ;
        RECT 64.345 172.195 65.690 172.425 ;
        RECT 66.225 172.195 70.775 173.105 ;
        RECT 70.795 173.065 71.715 173.105 ;
        RECT 70.785 172.875 71.715 173.065 ;
        RECT 73.805 172.875 75.375 173.105 ;
        RECT 70.785 172.515 75.375 172.875 ;
        RECT 70.795 172.425 75.375 172.515 ;
        RECT 75.385 172.425 77.215 173.105 ;
        RECT 70.795 172.195 73.795 172.425 ;
        RECT 75.870 172.195 77.215 172.425 ;
        RECT 78.145 172.295 81.815 173.105 ;
        RECT 81.825 172.195 85.300 173.105 ;
        RECT 85.965 172.295 88.715 173.105 ;
        RECT 88.735 172.235 89.165 173.020 ;
        RECT 89.645 172.295 91.475 173.105 ;
        RECT 91.485 172.425 92.850 173.105 ;
        RECT 93.325 172.295 96.075 173.105 ;
        RECT 96.085 172.325 97.455 173.105 ;
        RECT 97.925 172.295 100.675 173.105 ;
        RECT 100.770 172.425 109.875 173.105 ;
        RECT 110.575 172.425 114.475 173.105 ;
        RECT 113.545 172.195 114.475 172.425 ;
        RECT 114.495 172.235 114.925 173.020 ;
        RECT 115.865 172.425 125.055 173.105 ;
        RECT 115.865 172.195 116.785 172.425 ;
        RECT 119.615 172.205 120.545 172.425 ;
        RECT 125.065 172.295 126.435 173.105 ;
        RECT 126.445 172.295 127.815 173.105 ;
      LAYER nwell ;
        RECT 14.470 169.075 128.010 171.905 ;
      LAYER pwell ;
        RECT 14.665 167.875 16.035 168.685 ;
        RECT 16.045 167.875 18.795 168.685 ;
        RECT 18.805 167.875 24.315 168.685 ;
        RECT 24.335 167.960 24.765 168.745 ;
        RECT 24.870 167.875 33.975 168.555 ;
        RECT 34.180 167.875 37.655 168.785 ;
        RECT 37.665 167.875 39.035 168.685 ;
        RECT 39.045 167.875 44.555 168.685 ;
        RECT 44.565 167.875 50.075 168.685 ;
        RECT 50.095 167.960 50.525 168.745 ;
        RECT 51.465 167.875 55.135 168.685 ;
        RECT 55.155 167.875 56.505 168.785 ;
        RECT 57.445 167.875 58.815 168.655 ;
        RECT 58.965 167.875 61.575 168.785 ;
        RECT 61.585 167.875 62.955 168.685 ;
        RECT 62.965 167.875 68.475 168.685 ;
        RECT 68.495 167.875 69.845 168.785 ;
        RECT 70.105 168.105 72.860 168.785 ;
        RECT 70.105 167.875 72.375 168.105 ;
        RECT 73.085 167.875 75.835 168.685 ;
        RECT 75.855 167.960 76.285 168.745 ;
        RECT 76.765 167.875 82.275 168.685 ;
        RECT 85.485 168.555 86.415 168.785 ;
        RECT 82.515 167.875 86.415 168.555 ;
        RECT 86.435 167.875 87.785 168.785 ;
        RECT 88.265 167.875 90.095 168.685 ;
        RECT 90.115 167.875 91.465 168.785 ;
        RECT 91.485 168.555 92.405 168.785 ;
        RECT 95.235 168.555 96.165 168.775 ;
        RECT 91.485 167.875 100.675 168.555 ;
        RECT 101.615 167.960 102.045 168.745 ;
        RECT 102.535 167.875 103.885 168.785 ;
        RECT 103.905 168.555 104.825 168.785 ;
        RECT 107.655 168.555 108.585 168.775 ;
        RECT 103.905 167.875 113.095 168.555 ;
        RECT 113.105 167.875 114.935 168.685 ;
        RECT 114.945 167.875 120.455 168.685 ;
        RECT 120.465 167.875 121.835 168.655 ;
        RECT 121.845 167.875 123.675 168.555 ;
        RECT 123.685 167.875 126.435 168.685 ;
        RECT 126.445 167.875 127.815 168.685 ;
        RECT 14.805 167.665 14.975 167.875 ;
        RECT 18.485 167.685 18.655 167.875 ;
        RECT 24.005 167.685 24.175 167.875 ;
        RECT 25.385 167.665 25.555 167.855 ;
        RECT 25.900 167.715 26.020 167.825 ;
        RECT 31.365 167.665 31.535 167.855 ;
        RECT 33.665 167.685 33.835 167.875 ;
        RECT 36.885 167.665 37.055 167.855 ;
        RECT 37.340 167.685 37.510 167.875 ;
        RECT 37.860 167.715 37.980 167.825 ;
        RECT 38.725 167.685 38.895 167.875 ;
        RECT 40.565 167.665 40.735 167.855 ;
        RECT 44.245 167.685 44.415 167.875 ;
        RECT 46.085 167.665 46.255 167.855 ;
        RECT 49.765 167.685 49.935 167.875 ;
        RECT 51.145 167.720 51.305 167.830 ;
        RECT 51.605 167.665 51.775 167.855 ;
        RECT 54.825 167.685 54.995 167.875 ;
        RECT 56.205 167.685 56.375 167.875 ;
        RECT 57.125 167.720 57.285 167.830 ;
        RECT 57.585 167.685 57.755 167.875 ;
        RECT 60.805 167.665 60.975 167.855 ;
        RECT 61.260 167.685 61.430 167.875 ;
        RECT 62.645 167.665 62.815 167.875 ;
        RECT 64.485 167.665 64.655 167.855 ;
        RECT 68.165 167.685 68.335 167.875 ;
        RECT 68.625 167.685 68.795 167.875 ;
        RECT 70.105 167.855 70.175 167.875 ;
        RECT 70.005 167.665 70.175 167.855 ;
        RECT 71.845 167.665 72.015 167.855 ;
        RECT 73.225 167.665 73.395 167.855 ;
        RECT 75.525 167.685 75.695 167.875 ;
        RECT 76.500 167.715 76.620 167.825 ;
        RECT 78.745 167.665 78.915 167.855 ;
        RECT 79.205 167.665 79.375 167.855 ;
        RECT 81.965 167.685 82.135 167.875 ;
        RECT 85.830 167.685 86.000 167.875 ;
        RECT 87.485 167.685 87.655 167.875 ;
        RECT 88.000 167.715 88.120 167.825 ;
        RECT 89.785 167.685 89.955 167.875 ;
        RECT 90.245 167.665 90.415 167.875 ;
        RECT 91.165 167.710 91.325 167.820 ;
        RECT 95.030 167.665 95.200 167.855 ;
        RECT 96.685 167.665 96.855 167.855 ;
        RECT 100.365 167.685 100.535 167.875 ;
        RECT 101.285 167.720 101.445 167.830 ;
        RECT 102.205 167.825 102.375 167.855 ;
        RECT 102.205 167.715 102.380 167.825 ;
        RECT 102.205 167.665 102.375 167.715 ;
        RECT 102.665 167.685 102.835 167.875 ;
        RECT 106.070 167.665 106.240 167.855 ;
        RECT 106.860 167.715 106.980 167.825 ;
        RECT 110.670 167.665 110.840 167.855 ;
        RECT 112.325 167.665 112.495 167.855 ;
        RECT 112.785 167.685 112.955 167.875 ;
        RECT 114.165 167.665 114.335 167.855 ;
        RECT 114.625 167.685 114.795 167.875 ;
        RECT 118.490 167.665 118.660 167.855 ;
        RECT 119.225 167.665 119.395 167.855 ;
        RECT 120.145 167.685 120.315 167.875 ;
        RECT 120.605 167.825 120.775 167.875 ;
        RECT 120.605 167.715 120.780 167.825 ;
        RECT 120.605 167.685 120.775 167.715 ;
        RECT 121.065 167.665 121.235 167.855 ;
        RECT 122.500 167.715 122.620 167.825 ;
        RECT 123.365 167.685 123.535 167.875 ;
        RECT 126.125 167.665 126.295 167.875 ;
        RECT 127.505 167.665 127.675 167.875 ;
        RECT 14.665 166.855 16.035 167.665 ;
        RECT 16.415 166.985 25.695 167.665 ;
        RECT 16.415 166.865 18.750 166.985 ;
        RECT 16.415 166.755 17.335 166.865 ;
        RECT 23.415 166.765 24.335 166.985 ;
        RECT 26.165 166.855 31.675 167.665 ;
        RECT 31.685 166.855 37.195 167.665 ;
        RECT 37.215 166.795 37.645 167.580 ;
        RECT 38.125 166.855 40.875 167.665 ;
        RECT 40.885 166.855 46.395 167.665 ;
        RECT 46.405 166.855 51.915 167.665 ;
        RECT 51.925 166.985 61.115 167.665 ;
        RECT 51.925 166.755 52.845 166.985 ;
        RECT 55.675 166.765 56.605 166.985 ;
        RECT 61.125 166.855 62.955 167.665 ;
        RECT 62.975 166.795 63.405 167.580 ;
        RECT 63.425 166.855 64.795 167.665 ;
        RECT 64.805 166.855 70.315 167.665 ;
        RECT 70.325 166.985 72.155 167.665 ;
        RECT 70.325 166.755 71.670 166.985 ;
        RECT 72.165 166.855 73.535 167.665 ;
        RECT 73.545 166.855 79.055 167.665 ;
        RECT 79.065 166.985 88.345 167.665 ;
        RECT 80.425 166.765 81.345 166.985 ;
        RECT 86.010 166.865 88.345 166.985 ;
        RECT 87.425 166.755 88.345 166.865 ;
        RECT 88.735 166.795 89.165 167.580 ;
        RECT 89.185 166.885 90.555 167.665 ;
        RECT 91.715 166.985 95.615 167.665 ;
        RECT 94.685 166.755 95.615 166.985 ;
        RECT 95.625 166.855 96.995 167.665 ;
        RECT 97.005 166.855 102.515 167.665 ;
        RECT 102.755 166.985 106.655 167.665 ;
        RECT 107.355 166.985 111.255 167.665 ;
        RECT 105.725 166.755 106.655 166.985 ;
        RECT 110.325 166.755 111.255 166.985 ;
        RECT 111.265 166.885 112.635 167.665 ;
        RECT 112.645 166.855 114.475 167.665 ;
        RECT 114.495 166.795 114.925 167.580 ;
        RECT 115.175 166.985 119.075 167.665 ;
        RECT 118.145 166.755 119.075 166.985 ;
        RECT 119.095 166.755 120.445 167.665 ;
        RECT 120.925 166.885 122.295 167.665 ;
        RECT 122.765 166.855 126.435 167.665 ;
        RECT 126.445 166.855 127.815 167.665 ;
      LAYER nwell ;
        RECT 14.470 163.635 128.010 166.465 ;
      LAYER pwell ;
        RECT 14.665 162.435 16.035 163.245 ;
        RECT 16.045 162.435 18.795 163.245 ;
        RECT 18.815 162.435 20.165 163.345 ;
        RECT 23.385 163.115 24.315 163.345 ;
        RECT 20.415 162.435 24.315 163.115 ;
        RECT 24.335 162.520 24.765 163.305 ;
        RECT 25.245 162.435 26.615 163.215 ;
        RECT 26.625 162.435 28.455 163.245 ;
        RECT 28.475 162.435 29.825 163.345 ;
        RECT 29.845 163.115 30.765 163.345 ;
        RECT 33.595 163.115 34.525 163.335 ;
        RECT 39.045 163.115 39.975 163.345 ;
        RECT 29.845 162.435 39.035 163.115 ;
        RECT 39.045 162.435 42.945 163.115 ;
        RECT 43.195 162.435 44.545 163.345 ;
        RECT 44.565 162.435 45.935 163.245 ;
        RECT 49.145 163.115 50.075 163.345 ;
        RECT 46.175 162.435 50.075 163.115 ;
        RECT 50.095 162.520 50.525 163.305 ;
        RECT 50.545 162.435 52.375 163.245 ;
        RECT 52.395 162.435 53.745 163.345 ;
        RECT 53.765 163.115 54.685 163.345 ;
        RECT 57.515 163.115 58.445 163.335 ;
        RECT 53.765 162.435 62.955 163.115 ;
        RECT 62.965 162.435 64.335 163.245 ;
        RECT 64.485 162.435 67.095 163.345 ;
        RECT 67.245 162.435 69.855 163.345 ;
        RECT 70.325 162.435 73.045 163.345 ;
        RECT 73.085 162.435 75.825 163.115 ;
        RECT 75.855 162.520 76.285 163.305 ;
        RECT 77.135 163.235 78.055 163.345 ;
        RECT 77.135 163.115 79.470 163.235 ;
        RECT 84.135 163.115 85.055 163.335 ;
        RECT 77.135 162.435 86.415 163.115 ;
        RECT 86.425 162.435 87.795 163.215 ;
        RECT 87.815 162.435 89.165 163.345 ;
        RECT 89.645 162.435 95.155 163.245 ;
        RECT 98.365 163.115 99.295 163.345 ;
        RECT 95.395 162.435 99.295 163.115 ;
        RECT 100.235 162.435 101.585 163.345 ;
        RECT 101.615 162.520 102.045 163.305 ;
        RECT 102.435 163.235 103.355 163.345 ;
        RECT 102.435 163.115 104.770 163.235 ;
        RECT 109.435 163.115 110.355 163.335 ;
        RECT 115.385 163.115 116.315 163.345 ;
        RECT 102.435 162.435 111.715 163.115 ;
        RECT 112.415 162.435 116.315 163.115 ;
        RECT 116.325 163.115 117.245 163.345 ;
        RECT 120.075 163.115 121.005 163.335 ;
        RECT 116.325 162.435 125.515 163.115 ;
        RECT 126.445 162.435 127.815 163.245 ;
        RECT 14.805 162.225 14.975 162.435 ;
        RECT 16.240 162.275 16.360 162.385 ;
        RECT 17.565 162.225 17.735 162.415 ;
        RECT 18.485 162.245 18.655 162.435 ;
        RECT 18.945 162.245 19.115 162.435 ;
        RECT 23.730 162.245 23.900 162.435 ;
        RECT 24.980 162.275 25.100 162.385 ;
        RECT 25.385 162.245 25.555 162.435 ;
        RECT 27.225 162.225 27.395 162.415 ;
        RECT 27.685 162.225 27.855 162.415 ;
        RECT 28.145 162.245 28.315 162.435 ;
        RECT 28.605 162.245 28.775 162.435 ;
        RECT 38.725 162.225 38.895 162.435 ;
        RECT 39.460 162.245 39.630 162.435 ;
        RECT 40.105 162.225 40.275 162.415 ;
        RECT 44.245 162.245 44.415 162.435 ;
        RECT 45.625 162.245 45.795 162.435 ;
        RECT 49.305 162.225 49.475 162.415 ;
        RECT 49.490 162.245 49.660 162.435 ;
        RECT 50.685 162.225 50.855 162.415 ;
        RECT 51.605 162.270 51.765 162.380 ;
        RECT 52.065 162.225 52.235 162.435 ;
        RECT 52.525 162.245 52.695 162.435 ;
        RECT 62.645 162.415 62.815 162.435 ;
        RECT 56.850 162.225 57.020 162.415 ;
        RECT 58.505 162.225 58.675 162.415 ;
        RECT 58.965 162.225 59.135 162.415 ;
        RECT 62.640 162.245 62.815 162.415 ;
        RECT 63.620 162.275 63.740 162.385 ;
        RECT 64.025 162.245 64.195 162.435 ;
        RECT 62.640 162.225 62.810 162.245 ;
        RECT 65.405 162.225 65.575 162.415 ;
        RECT 66.780 162.245 66.950 162.435 ;
        RECT 69.540 162.415 69.710 162.435 ;
        RECT 68.165 162.225 68.335 162.415 ;
        RECT 69.540 162.245 69.715 162.415 ;
        RECT 70.060 162.275 70.180 162.385 ;
        RECT 70.465 162.245 70.635 162.435 ;
        RECT 69.545 162.225 69.715 162.245 ;
        RECT 71.385 162.225 71.555 162.415 ;
        RECT 71.900 162.275 72.020 162.385 ;
        RECT 73.225 162.245 73.395 162.435 ;
        RECT 73.685 162.225 73.855 162.415 ;
        RECT 76.500 162.275 76.620 162.385 ;
        RECT 79.205 162.225 79.375 162.415 ;
        RECT 83.070 162.225 83.240 162.415 ;
        RECT 84.265 162.270 84.425 162.380 ;
        RECT 85.645 162.225 85.815 162.415 ;
        RECT 86.105 162.245 86.275 162.435 ;
        RECT 86.565 162.270 86.725 162.380 ;
        RECT 87.025 162.225 87.195 162.415 ;
        RECT 87.485 162.245 87.655 162.435 ;
        RECT 88.460 162.275 88.580 162.385 ;
        RECT 88.865 162.245 89.035 162.435 ;
        RECT 89.380 162.275 89.500 162.385 ;
        RECT 90.245 162.225 90.415 162.415 ;
        RECT 94.845 162.245 95.015 162.435 ;
        RECT 98.710 162.245 98.880 162.435 ;
        RECT 99.905 162.225 100.075 162.415 ;
        RECT 100.365 162.245 100.535 162.435 ;
        RECT 101.285 162.225 101.455 162.415 ;
        RECT 102.205 162.270 102.365 162.380 ;
        RECT 105.885 162.225 106.055 162.415 ;
        RECT 106.345 162.225 106.515 162.415 ;
        RECT 108.645 162.225 108.815 162.415 ;
        RECT 111.405 162.245 111.575 162.435 ;
        RECT 111.920 162.275 112.040 162.385 ;
        RECT 114.165 162.225 114.335 162.415 ;
        RECT 115.140 162.275 115.260 162.385 ;
        RECT 115.730 162.245 115.900 162.435 ;
        RECT 116.925 162.225 117.095 162.415 ;
        RECT 119.680 162.225 119.850 162.415 ;
        RECT 120.605 162.270 120.765 162.380 ;
        RECT 125.205 162.245 125.375 162.435 ;
        RECT 126.125 162.225 126.295 162.415 ;
        RECT 127.505 162.225 127.675 162.435 ;
        RECT 14.665 161.415 16.035 162.225 ;
        RECT 16.515 161.315 17.865 162.225 ;
        RECT 18.255 161.545 27.535 162.225 ;
        RECT 27.545 161.545 36.825 162.225 ;
        RECT 18.255 161.425 20.590 161.545 ;
        RECT 18.255 161.315 19.175 161.425 ;
        RECT 25.255 161.325 26.175 161.545 ;
        RECT 28.905 161.325 29.825 161.545 ;
        RECT 34.490 161.425 36.825 161.545 ;
        RECT 35.905 161.315 36.825 161.425 ;
        RECT 37.215 161.355 37.645 162.140 ;
        RECT 37.665 161.445 39.035 162.225 ;
        RECT 39.045 161.445 40.415 162.225 ;
        RECT 40.425 161.545 49.615 162.225 ;
        RECT 40.425 161.315 41.345 161.545 ;
        RECT 44.175 161.325 45.105 161.545 ;
        RECT 49.625 161.445 50.995 162.225 ;
        RECT 51.935 161.315 53.285 162.225 ;
        RECT 53.535 161.545 57.435 162.225 ;
        RECT 56.505 161.315 57.435 161.545 ;
        RECT 57.445 161.415 58.815 162.225 ;
        RECT 58.825 161.445 60.195 162.225 ;
        RECT 60.345 161.315 62.955 162.225 ;
        RECT 62.975 161.355 63.405 162.140 ;
        RECT 63.885 161.415 65.715 162.225 ;
        RECT 65.735 161.545 68.475 162.225 ;
        RECT 68.485 161.415 69.855 162.225 ;
        RECT 69.865 161.545 71.695 162.225 ;
        RECT 69.865 161.315 71.210 161.545 ;
        RECT 72.165 161.415 73.995 162.225 ;
        RECT 74.005 161.415 79.515 162.225 ;
        RECT 79.755 161.545 83.655 162.225 ;
        RECT 82.725 161.315 83.655 161.545 ;
        RECT 84.595 161.315 85.945 162.225 ;
        RECT 86.885 161.445 88.255 162.225 ;
        RECT 88.735 161.355 89.165 162.140 ;
        RECT 89.185 161.415 90.555 162.225 ;
        RECT 90.935 161.545 100.215 162.225 ;
        RECT 90.935 161.425 93.270 161.545 ;
        RECT 90.935 161.315 91.855 161.425 ;
        RECT 97.935 161.325 98.855 161.545 ;
        RECT 100.225 161.445 101.595 162.225 ;
        RECT 102.525 161.415 106.195 162.225 ;
        RECT 106.205 161.445 107.575 162.225 ;
        RECT 107.585 161.415 108.955 162.225 ;
        RECT 108.965 161.415 114.475 162.225 ;
        RECT 114.495 161.355 114.925 162.140 ;
        RECT 115.405 161.415 117.235 162.225 ;
        RECT 117.385 161.315 119.995 162.225 ;
        RECT 120.925 161.415 126.435 162.225 ;
        RECT 126.445 161.415 127.815 162.225 ;
      LAYER nwell ;
        RECT 14.470 158.195 128.010 161.025 ;
      LAYER pwell ;
        RECT 14.665 156.995 16.035 157.805 ;
        RECT 16.045 156.995 18.795 157.805 ;
        RECT 18.805 156.995 20.175 157.775 ;
        RECT 20.185 157.675 21.115 157.905 ;
        RECT 20.185 156.995 24.085 157.675 ;
        RECT 24.335 157.080 24.765 157.865 ;
        RECT 24.785 156.995 26.155 157.805 ;
        RECT 26.165 156.995 31.675 157.805 ;
        RECT 31.695 156.995 33.045 157.905 ;
        RECT 36.265 157.675 37.195 157.905 ;
        RECT 33.295 156.995 37.195 157.675 ;
        RECT 37.205 156.995 39.955 157.805 ;
        RECT 39.965 156.995 43.440 157.905 ;
        RECT 44.105 156.995 45.935 157.805 ;
        RECT 49.145 157.675 50.075 157.905 ;
        RECT 46.175 156.995 50.075 157.675 ;
        RECT 50.095 157.080 50.525 157.865 ;
        RECT 50.545 156.995 51.915 157.805 ;
        RECT 51.925 157.675 52.845 157.905 ;
        RECT 55.675 157.675 56.605 157.895 ;
        RECT 51.925 156.995 61.115 157.675 ;
        RECT 61.585 156.995 64.335 157.805 ;
        RECT 64.345 157.675 65.690 157.905 ;
        RECT 66.185 157.675 67.530 157.905 ;
        RECT 68.510 157.675 69.855 157.905 ;
        RECT 70.350 157.675 71.695 157.905 ;
        RECT 64.345 156.995 66.175 157.675 ;
        RECT 66.185 156.995 68.015 157.675 ;
        RECT 68.025 156.995 69.855 157.675 ;
        RECT 69.865 156.995 71.695 157.675 ;
        RECT 72.165 156.995 75.835 157.805 ;
        RECT 75.855 157.080 76.285 157.865 ;
        RECT 77.225 156.995 80.895 157.805 ;
        RECT 81.275 157.795 82.195 157.905 ;
        RECT 81.275 157.675 83.610 157.795 ;
        RECT 88.275 157.675 89.195 157.895 ;
        RECT 81.275 156.995 90.555 157.675 ;
        RECT 90.565 156.995 94.235 157.805 ;
        RECT 94.255 156.995 95.605 157.905 ;
        RECT 96.085 156.995 101.595 157.805 ;
        RECT 101.615 157.080 102.045 157.865 ;
        RECT 102.525 156.995 104.355 157.805 ;
        RECT 104.365 156.995 107.840 157.905 ;
        RECT 108.505 156.995 110.335 157.805 ;
        RECT 110.345 156.995 115.855 157.805 ;
        RECT 115.865 156.995 118.475 157.905 ;
        RECT 119.085 156.995 120.915 157.805 ;
        RECT 120.925 156.995 126.435 157.805 ;
        RECT 126.445 156.995 127.815 157.805 ;
        RECT 14.805 156.785 14.975 156.995 ;
        RECT 16.645 156.830 16.805 156.940 ;
        RECT 18.485 156.805 18.655 156.995 ;
        RECT 18.945 156.805 19.115 156.995 ;
        RECT 20.600 156.805 20.770 156.995 ;
        RECT 25.845 156.805 26.015 156.995 ;
        RECT 26.305 156.785 26.475 156.975 ;
        RECT 27.685 156.785 27.855 156.975 ;
        RECT 31.365 156.785 31.535 156.995 ;
        RECT 31.825 156.805 31.995 156.995 ;
        RECT 36.610 156.805 36.780 156.995 ;
        RECT 36.885 156.785 37.055 156.975 ;
        RECT 37.860 156.835 37.980 156.945 ;
        RECT 39.645 156.785 39.815 156.995 ;
        RECT 40.110 156.805 40.280 156.995 ;
        RECT 43.840 156.835 43.960 156.945 ;
        RECT 45.165 156.785 45.335 156.975 ;
        RECT 45.625 156.805 45.795 156.995 ;
        RECT 49.490 156.805 49.660 156.995 ;
        RECT 50.685 156.785 50.855 156.975 ;
        RECT 51.605 156.805 51.775 156.995 ;
        RECT 54.550 156.785 54.720 156.975 ;
        RECT 56.205 156.785 56.375 156.975 ;
        RECT 56.665 156.785 56.835 156.975 ;
        RECT 58.965 156.785 59.135 156.975 ;
        RECT 60.805 156.805 60.975 156.995 ;
        RECT 61.320 156.835 61.440 156.945 ;
        RECT 62.645 156.785 62.815 156.975 ;
        RECT 64.025 156.805 64.195 156.995 ;
        RECT 65.865 156.785 66.035 156.995 ;
        RECT 67.705 156.785 67.875 156.995 ;
        RECT 68.165 156.785 68.335 156.995 ;
        RECT 70.005 156.785 70.175 156.995 ;
        RECT 71.900 156.835 72.020 156.945 ;
        RECT 73.225 156.785 73.395 156.975 ;
        RECT 74.605 156.785 74.775 156.975 ;
        RECT 75.525 156.805 75.695 156.995 ;
        RECT 76.905 156.840 77.065 156.950 ;
        RECT 78.285 156.785 78.455 156.975 ;
        RECT 78.750 156.785 78.920 156.975 ;
        RECT 80.585 156.805 80.755 156.995 ;
        RECT 82.480 156.835 82.600 156.945 ;
        RECT 86.290 156.785 86.460 156.975 ;
        RECT 88.405 156.785 88.575 156.975 ;
        RECT 89.380 156.835 89.500 156.945 ;
        RECT 90.245 156.805 90.415 156.995 ;
        RECT 92.085 156.785 92.255 156.975 ;
        RECT 93.925 156.805 94.095 156.995 ;
        RECT 95.305 156.805 95.475 156.995 ;
        RECT 95.820 156.835 95.940 156.945 ;
        RECT 97.605 156.785 97.775 156.975 ;
        RECT 98.070 156.785 98.240 156.975 ;
        RECT 101.285 156.805 101.455 156.995 ;
        RECT 102.260 156.835 102.380 156.945 ;
        RECT 103.125 156.785 103.295 156.975 ;
        RECT 103.590 156.785 103.760 156.975 ;
        RECT 104.045 156.805 104.215 156.995 ;
        RECT 104.510 156.805 104.680 156.995 ;
        RECT 107.270 156.785 107.440 156.975 ;
        RECT 108.240 156.835 108.360 156.945 ;
        RECT 110.025 156.805 110.195 156.995 ;
        RECT 110.950 156.785 111.120 156.975 ;
        RECT 115.085 156.785 115.255 156.975 ;
        RECT 115.545 156.805 115.715 156.995 ;
        RECT 116.010 156.805 116.180 156.995 ;
        RECT 118.820 156.835 118.940 156.945 ;
        RECT 120.605 156.805 120.775 156.995 ;
        RECT 125.205 156.785 125.375 156.975 ;
        RECT 126.125 156.805 126.295 156.995 ;
        RECT 127.505 156.785 127.675 156.995 ;
        RECT 14.665 155.975 16.035 156.785 ;
        RECT 17.335 156.105 26.615 156.785 ;
        RECT 17.335 155.985 19.670 156.105 ;
        RECT 17.335 155.875 18.255 155.985 ;
        RECT 24.335 155.885 25.255 156.105 ;
        RECT 26.625 155.975 27.995 156.785 ;
        RECT 28.005 155.975 31.675 156.785 ;
        RECT 31.685 155.975 37.195 156.785 ;
        RECT 37.215 155.915 37.645 156.700 ;
        RECT 38.125 155.975 39.955 156.785 ;
        RECT 39.965 155.975 45.475 156.785 ;
        RECT 45.485 155.975 50.995 156.785 ;
        RECT 51.235 156.105 55.135 156.785 ;
        RECT 54.205 155.875 55.135 156.105 ;
        RECT 55.145 155.975 56.515 156.785 ;
        RECT 56.525 156.005 57.895 156.785 ;
        RECT 57.905 155.975 59.275 156.785 ;
        RECT 59.285 155.975 62.955 156.785 ;
        RECT 62.975 155.915 63.405 156.700 ;
        RECT 63.425 155.975 66.175 156.785 ;
        RECT 66.185 156.105 68.015 156.785 ;
        RECT 68.025 156.105 69.855 156.785 ;
        RECT 69.865 156.105 71.695 156.785 ;
        RECT 66.185 155.875 67.530 156.105 ;
        RECT 68.510 155.875 69.855 156.105 ;
        RECT 70.350 155.875 71.695 156.105 ;
        RECT 71.705 156.105 73.535 156.785 ;
        RECT 71.705 155.875 73.050 156.105 ;
        RECT 73.545 155.975 74.915 156.785 ;
        RECT 74.925 155.975 78.595 156.785 ;
        RECT 78.605 155.875 82.080 156.785 ;
        RECT 82.975 156.105 86.875 156.785 ;
        RECT 85.945 155.875 86.875 156.105 ;
        RECT 86.885 155.975 88.715 156.785 ;
        RECT 88.735 155.915 89.165 156.700 ;
        RECT 89.645 155.975 92.395 156.785 ;
        RECT 92.405 155.975 97.915 156.785 ;
        RECT 97.925 155.875 101.400 156.785 ;
        RECT 101.605 155.975 103.435 156.785 ;
        RECT 103.445 155.875 106.920 156.785 ;
        RECT 107.125 155.875 110.600 156.785 ;
        RECT 110.805 155.875 114.280 156.785 ;
        RECT 114.495 155.915 114.925 156.700 ;
        RECT 114.955 155.875 116.305 156.785 ;
        RECT 116.325 156.105 125.515 156.785 ;
        RECT 116.325 155.875 117.245 156.105 ;
        RECT 120.075 155.885 121.005 156.105 ;
        RECT 126.445 155.975 127.815 156.785 ;
      LAYER nwell ;
        RECT 14.470 152.755 128.010 155.585 ;
      LAYER pwell ;
        RECT 14.665 151.555 16.035 152.365 ;
        RECT 16.505 151.555 20.175 152.365 ;
        RECT 23.385 152.235 24.315 152.465 ;
        RECT 20.415 151.555 24.315 152.235 ;
        RECT 24.335 151.640 24.765 152.425 ;
        RECT 24.785 151.555 26.615 152.365 ;
        RECT 29.825 152.235 30.755 152.465 ;
        RECT 26.855 151.555 30.755 152.235 ;
        RECT 31.420 151.555 34.895 152.465 ;
        RECT 34.905 151.555 38.380 152.465 ;
        RECT 39.045 151.555 42.715 152.365 ;
        RECT 42.920 151.555 46.395 152.465 ;
        RECT 46.600 151.555 50.075 152.465 ;
        RECT 50.095 151.640 50.525 152.425 ;
        RECT 50.545 151.555 54.020 152.465 ;
        RECT 54.685 151.555 56.515 152.365 ;
        RECT 56.525 151.555 62.035 152.365 ;
        RECT 62.055 151.555 63.405 152.465 ;
        RECT 63.425 152.235 64.770 152.465 ;
        RECT 63.425 151.555 65.255 152.235 ;
        RECT 65.265 151.555 68.740 152.465 ;
        RECT 69.875 151.555 72.615 152.235 ;
        RECT 72.625 151.555 75.345 152.465 ;
        RECT 75.855 151.640 76.285 152.425 ;
        RECT 76.305 151.555 77.675 152.365 ;
        RECT 77.685 151.555 81.160 152.465 ;
        RECT 81.365 151.555 84.840 152.465 ;
        RECT 85.965 151.555 89.635 152.365 ;
        RECT 89.645 151.555 95.155 152.365 ;
        RECT 95.175 151.555 96.525 152.465 ;
        RECT 97.465 151.555 98.835 152.335 ;
        RECT 98.845 151.555 101.595 152.365 ;
        RECT 101.615 151.640 102.045 152.425 ;
        RECT 102.065 151.555 107.575 152.365 ;
        RECT 107.585 151.555 111.060 152.465 ;
        RECT 111.265 151.555 114.935 152.365 ;
        RECT 118.145 152.235 119.075 152.465 ;
        RECT 115.175 151.555 119.075 152.235 ;
        RECT 119.555 151.555 120.905 152.465 ;
        RECT 121.385 151.555 122.755 152.335 ;
        RECT 122.765 151.555 124.135 152.335 ;
        RECT 124.605 151.555 126.435 152.365 ;
        RECT 126.445 151.555 127.815 152.365 ;
        RECT 14.805 151.345 14.975 151.555 ;
        RECT 16.240 151.395 16.360 151.505 ;
        RECT 16.645 151.390 16.805 151.500 ;
        RECT 18.025 151.345 18.195 151.535 ;
        RECT 18.485 151.345 18.655 151.535 ;
        RECT 19.865 151.365 20.035 151.555 ;
        RECT 23.730 151.365 23.900 151.555 ;
        RECT 26.305 151.365 26.475 151.555 ;
        RECT 29.065 151.345 29.235 151.535 ;
        RECT 30.170 151.365 30.340 151.555 ;
        RECT 30.445 151.345 30.615 151.535 ;
        RECT 30.960 151.395 31.080 151.505 ;
        RECT 33.205 151.345 33.375 151.535 ;
        RECT 34.580 151.365 34.750 151.555 ;
        RECT 35.050 151.365 35.220 151.555 ;
        RECT 42.405 151.535 42.575 151.555 ;
        RECT 36.880 151.345 37.050 151.535 ;
        RECT 38.265 151.390 38.425 151.500 ;
        RECT 38.730 151.345 38.900 151.535 ;
        RECT 42.405 151.365 42.580 151.535 ;
        RECT 46.080 151.365 46.250 151.555 ;
        RECT 42.410 151.345 42.580 151.365 ;
        RECT 48.385 151.345 48.555 151.535 ;
        RECT 48.850 151.345 49.020 151.535 ;
        RECT 49.760 151.365 49.930 151.555 ;
        RECT 50.690 151.365 50.860 151.555 ;
        RECT 53.445 151.345 53.615 151.535 ;
        RECT 54.420 151.395 54.540 151.505 ;
        RECT 56.205 151.365 56.375 151.555 ;
        RECT 58.965 151.345 59.135 151.535 ;
        RECT 59.430 151.345 59.600 151.535 ;
        RECT 61.725 151.365 61.895 151.555 ;
        RECT 62.185 151.365 62.355 151.555 ;
        RECT 64.945 151.365 65.115 151.555 ;
        RECT 65.410 151.365 65.580 151.555 ;
        RECT 69.545 151.400 69.705 151.510 ;
        RECT 72.305 151.345 72.475 151.555 ;
        RECT 72.765 151.345 72.935 151.555 ;
        RECT 74.605 151.345 74.775 151.535 ;
        RECT 75.580 151.395 75.700 151.505 ;
        RECT 76.445 151.345 76.615 151.535 ;
        RECT 77.365 151.365 77.535 151.555 ;
        RECT 77.830 151.365 78.000 151.555 ;
        RECT 79.260 151.395 79.380 151.505 ;
        RECT 79.670 151.345 79.840 151.535 ;
        RECT 81.510 151.365 81.680 151.555 ;
        RECT 85.645 151.400 85.805 151.510 ;
        RECT 88.405 151.345 88.575 151.535 ;
        RECT 89.325 151.505 89.495 151.555 ;
        RECT 89.325 151.395 89.500 151.505 ;
        RECT 89.325 151.365 89.495 151.395 ;
        RECT 90.705 151.345 90.875 151.535 ;
        RECT 91.165 151.345 91.335 151.535 ;
        RECT 94.845 151.365 95.015 151.555 ;
        RECT 96.225 151.365 96.395 151.555 ;
        RECT 97.145 151.400 97.305 151.510 ;
        RECT 97.605 151.365 97.775 151.555 ;
        RECT 101.285 151.345 101.455 151.555 ;
        RECT 103.125 151.345 103.295 151.535 ;
        RECT 14.665 150.535 16.035 151.345 ;
        RECT 16.975 150.435 18.325 151.345 ;
        RECT 18.355 150.435 19.705 151.345 ;
        RECT 20.095 150.665 29.375 151.345 ;
        RECT 20.095 150.545 22.430 150.665 ;
        RECT 20.095 150.435 21.015 150.545 ;
        RECT 27.095 150.445 28.015 150.665 ;
        RECT 29.385 150.565 30.755 151.345 ;
        RECT 30.765 150.535 33.515 151.345 ;
        RECT 33.720 150.435 37.195 151.345 ;
        RECT 37.215 150.475 37.645 151.260 ;
        RECT 38.585 150.435 42.060 151.345 ;
        RECT 42.265 150.435 45.740 151.345 ;
        RECT 45.945 150.535 48.695 151.345 ;
        RECT 48.705 150.435 52.180 151.345 ;
        RECT 52.385 150.535 53.755 151.345 ;
        RECT 53.765 150.535 59.275 151.345 ;
        RECT 59.285 150.435 62.760 151.345 ;
        RECT 62.975 150.475 63.405 151.260 ;
        RECT 63.510 150.665 72.615 151.345 ;
        RECT 72.625 150.665 74.455 151.345 ;
        RECT 74.465 150.665 76.295 151.345 ;
        RECT 76.305 150.665 79.045 151.345 ;
        RECT 73.110 150.435 74.455 150.665 ;
        RECT 74.950 150.435 76.295 150.665 ;
        RECT 79.525 150.435 83.000 151.345 ;
        RECT 83.205 150.535 88.715 151.345 ;
        RECT 88.735 150.475 89.165 151.260 ;
        RECT 89.655 150.435 91.005 151.345 ;
        RECT 91.025 150.565 92.395 151.345 ;
        RECT 92.405 150.665 101.595 151.345 ;
        RECT 92.405 150.435 93.325 150.665 ;
        RECT 96.155 150.445 97.085 150.665 ;
        RECT 101.605 150.535 103.435 151.345 ;
        RECT 103.445 151.315 104.390 151.345 ;
        RECT 105.880 151.315 106.050 151.535 ;
        RECT 106.350 151.315 106.520 151.535 ;
        RECT 107.265 151.365 107.435 151.555 ;
        RECT 107.730 151.365 107.900 151.555 ;
        RECT 109.110 151.345 109.280 151.535 ;
        RECT 114.165 151.345 114.335 151.535 ;
        RECT 114.625 151.365 114.795 151.555 ;
        RECT 116.005 151.345 116.175 151.535 ;
        RECT 118.490 151.365 118.660 151.555 ;
        RECT 119.280 151.395 119.400 151.505 ;
        RECT 119.685 151.365 119.855 151.555 ;
        RECT 121.120 151.395 121.240 151.505 ;
        RECT 121.525 151.365 121.695 151.555 ;
        RECT 122.905 151.365 123.075 151.555 ;
        RECT 124.340 151.395 124.460 151.505 ;
        RECT 125.665 151.345 125.835 151.535 ;
        RECT 126.125 151.505 126.295 151.555 ;
        RECT 126.125 151.395 126.300 151.505 ;
        RECT 126.125 151.365 126.295 151.395 ;
        RECT 127.505 151.345 127.675 151.555 ;
        RECT 108.010 151.315 108.955 151.345 ;
        RECT 103.445 150.635 106.195 151.315 ;
        RECT 106.205 150.635 108.955 151.315 ;
        RECT 103.445 150.435 104.390 150.635 ;
        RECT 108.010 150.435 108.955 150.635 ;
        RECT 108.965 150.435 112.440 151.345 ;
        RECT 112.645 150.535 114.475 151.345 ;
        RECT 114.495 150.475 114.925 151.260 ;
        RECT 114.945 150.535 116.315 151.345 ;
        RECT 116.695 150.665 125.975 151.345 ;
        RECT 116.695 150.545 119.030 150.665 ;
        RECT 116.695 150.435 117.615 150.545 ;
        RECT 123.695 150.445 124.615 150.665 ;
        RECT 126.445 150.535 127.815 151.345 ;
      LAYER nwell ;
        RECT 14.470 147.315 128.010 150.145 ;
      LAYER pwell ;
        RECT 14.665 146.115 16.035 146.925 ;
        RECT 16.045 146.115 17.415 146.925 ;
        RECT 17.425 146.115 22.935 146.925 ;
        RECT 22.945 146.115 24.315 146.895 ;
        RECT 24.335 146.200 24.765 146.985 ;
        RECT 25.245 146.115 27.995 146.925 ;
        RECT 28.005 146.115 33.515 146.925 ;
        RECT 33.525 146.825 34.470 147.025 ;
        RECT 33.525 146.145 36.275 146.825 ;
        RECT 33.525 146.115 34.470 146.145 ;
        RECT 14.805 145.905 14.975 146.115 ;
        RECT 17.105 145.925 17.275 146.115 ;
        RECT 22.625 145.925 22.795 146.115 ;
        RECT 23.085 145.925 23.255 146.115 ;
        RECT 24.980 145.955 25.100 146.065 ;
        RECT 25.385 145.905 25.555 146.095 ;
        RECT 27.225 145.905 27.395 146.095 ;
        RECT 27.685 145.925 27.855 146.115 ;
        RECT 32.745 145.905 32.915 146.095 ;
        RECT 33.205 145.925 33.375 146.115 ;
        RECT 14.665 145.095 16.035 145.905 ;
        RECT 16.415 145.225 25.695 145.905 ;
        RECT 16.415 145.105 18.750 145.225 ;
        RECT 16.415 144.995 17.335 145.105 ;
        RECT 23.415 145.005 24.335 145.225 ;
        RECT 25.705 145.095 27.535 145.905 ;
        RECT 27.545 145.095 33.055 145.905 ;
        RECT 33.065 145.875 34.010 145.905 ;
        RECT 35.500 145.875 35.670 146.095 ;
        RECT 35.960 145.925 36.130 146.145 ;
        RECT 36.285 146.115 38.115 146.925 ;
        RECT 38.125 146.825 39.070 147.025 ;
        RECT 38.125 146.145 40.875 146.825 ;
        RECT 38.125 146.115 39.070 146.145 ;
        RECT 36.885 145.905 37.055 146.095 ;
        RECT 37.805 145.925 37.975 146.115 ;
        RECT 38.725 145.905 38.895 146.095 ;
        RECT 40.560 145.925 40.730 146.145 ;
        RECT 40.885 146.115 44.555 146.925 ;
        RECT 44.565 146.115 50.075 146.925 ;
        RECT 50.095 146.200 50.525 146.985 ;
        RECT 50.545 146.115 53.295 146.925 ;
        RECT 53.315 146.115 54.665 147.025 ;
        RECT 55.605 146.115 59.275 146.925 ;
        RECT 59.655 146.915 60.575 147.025 ;
        RECT 59.655 146.795 61.990 146.915 ;
        RECT 66.655 146.795 67.575 147.015 ;
        RECT 59.655 146.115 68.935 146.795 ;
        RECT 68.945 146.115 72.155 147.025 ;
        RECT 72.165 146.115 75.835 146.925 ;
        RECT 75.855 146.200 76.285 146.985 ;
        RECT 76.765 146.115 80.435 146.925 ;
        RECT 80.445 146.115 85.955 146.925 ;
        RECT 86.335 146.915 87.255 147.025 ;
        RECT 86.335 146.795 88.670 146.915 ;
        RECT 93.335 146.795 94.255 147.015 ;
        RECT 86.335 146.115 95.615 146.795 ;
        RECT 96.085 146.115 101.595 146.925 ;
        RECT 101.615 146.200 102.045 146.985 ;
        RECT 102.525 146.825 103.470 147.025 ;
        RECT 102.525 146.145 105.275 146.825 ;
        RECT 102.525 146.115 103.470 146.145 ;
        RECT 44.245 145.905 44.415 146.115 ;
        RECT 33.065 145.195 35.815 145.875 ;
        RECT 33.065 144.995 34.010 145.195 ;
        RECT 35.825 145.095 37.195 145.905 ;
        RECT 37.215 145.035 37.645 145.820 ;
        RECT 37.665 145.095 39.035 145.905 ;
        RECT 39.045 145.095 44.555 145.905 ;
        RECT 44.710 145.875 44.880 146.095 ;
        RECT 47.470 145.905 47.640 146.095 ;
        RECT 49.765 145.925 49.935 146.115 ;
        RECT 52.985 145.925 53.155 146.115 ;
        RECT 53.445 145.925 53.615 146.115 ;
        RECT 55.285 145.960 55.445 146.070 ;
        RECT 58.965 145.925 59.135 146.115 ;
        RECT 59.885 145.905 60.055 146.095 ;
        RECT 61.265 145.905 61.435 146.095 ;
        RECT 62.645 145.905 62.815 146.095 ;
        RECT 63.620 145.955 63.740 146.065 ;
        RECT 64.030 145.905 64.200 146.095 ;
        RECT 68.165 145.950 68.325 146.060 ;
        RECT 68.625 145.925 68.795 146.115 ;
        RECT 71.845 145.925 72.015 146.115 ;
        RECT 72.030 145.905 72.200 146.095 ;
        RECT 73.225 145.950 73.385 146.060 ;
        RECT 73.685 145.905 73.855 146.095 ;
        RECT 75.120 145.955 75.240 146.065 ;
        RECT 75.525 145.925 75.695 146.115 ;
        RECT 76.500 145.955 76.620 146.065 ;
        RECT 77.825 145.905 77.995 146.095 ;
        RECT 80.125 145.925 80.295 146.115 ;
        RECT 46.370 145.875 47.315 145.905 ;
        RECT 44.565 145.195 47.315 145.875 ;
        RECT 46.370 144.995 47.315 145.195 ;
        RECT 47.325 144.995 50.800 145.905 ;
        RECT 51.005 145.225 60.195 145.905 ;
        RECT 51.005 144.995 51.925 145.225 ;
        RECT 54.755 145.005 55.685 145.225 ;
        RECT 60.205 145.125 61.575 145.905 ;
        RECT 61.585 145.095 62.955 145.905 ;
        RECT 62.975 145.035 63.405 145.820 ;
        RECT 63.885 144.995 67.360 145.905 ;
        RECT 68.715 145.225 72.615 145.905 ;
        RECT 71.685 144.995 72.615 145.225 ;
        RECT 73.545 145.125 74.915 145.905 ;
        RECT 75.385 145.095 78.135 145.905 ;
        RECT 78.145 145.875 79.090 145.905 ;
        RECT 80.580 145.875 80.750 146.095 ;
        RECT 81.050 145.905 81.220 146.095 ;
        RECT 85.645 145.925 85.815 146.115 ;
        RECT 88.130 145.905 88.300 146.095 ;
        RECT 92.545 145.905 92.715 146.095 ;
        RECT 95.305 145.925 95.475 146.115 ;
        RECT 95.820 145.955 95.940 146.065 ;
        RECT 96.410 145.905 96.580 146.095 ;
        RECT 97.200 145.955 97.320 146.065 ;
        RECT 101.285 145.925 101.455 146.115 ;
        RECT 102.260 145.955 102.380 146.065 ;
        RECT 102.665 145.905 102.835 146.095 ;
        RECT 104.960 145.925 105.130 146.145 ;
        RECT 105.285 146.115 108.760 147.025 ;
        RECT 108.965 146.115 112.440 147.025 ;
        RECT 112.645 146.115 116.315 146.925 ;
        RECT 119.525 146.795 120.455 147.025 ;
        RECT 116.555 146.115 120.455 146.795 ;
        RECT 120.925 146.115 126.435 146.925 ;
        RECT 126.445 146.115 127.815 146.925 ;
        RECT 105.430 145.925 105.600 146.115 ;
        RECT 108.185 145.905 108.355 146.095 ;
        RECT 108.650 145.905 108.820 146.095 ;
        RECT 109.110 145.925 109.280 146.115 ;
        RECT 112.380 145.955 112.500 146.065 ;
        RECT 114.165 145.905 114.335 146.095 ;
        RECT 115.140 145.955 115.260 146.065 ;
        RECT 116.005 145.925 116.175 146.115 ;
        RECT 119.870 145.925 120.040 146.115 ;
        RECT 120.605 146.065 120.775 146.095 ;
        RECT 120.605 145.955 120.780 146.065 ;
        RECT 120.605 145.905 120.775 145.955 ;
        RECT 126.125 145.905 126.295 146.115 ;
        RECT 127.505 145.905 127.675 146.115 ;
        RECT 78.145 145.195 80.895 145.875 ;
        RECT 78.145 144.995 79.090 145.195 ;
        RECT 80.905 144.995 84.380 145.905 ;
        RECT 84.815 145.225 88.715 145.905 ;
        RECT 87.785 144.995 88.715 145.225 ;
        RECT 88.735 145.035 89.165 145.820 ;
        RECT 89.185 145.095 92.855 145.905 ;
        RECT 93.095 145.225 96.995 145.905 ;
        RECT 96.065 144.995 96.995 145.225 ;
        RECT 97.465 145.095 102.975 145.905 ;
        RECT 102.985 145.095 108.495 145.905 ;
        RECT 108.505 144.995 111.980 145.905 ;
        RECT 112.645 145.095 114.475 145.905 ;
        RECT 114.495 145.035 114.925 145.820 ;
        RECT 115.405 145.095 120.915 145.905 ;
        RECT 120.925 145.095 126.435 145.905 ;
        RECT 126.445 145.095 127.815 145.905 ;
      LAYER nwell ;
        RECT 14.470 141.875 128.010 144.705 ;
      LAYER pwell ;
        RECT 14.665 140.675 16.035 141.485 ;
        RECT 16.045 140.675 18.795 141.485 ;
        RECT 18.805 140.675 24.315 141.485 ;
        RECT 24.335 140.760 24.765 141.545 ;
        RECT 33.285 141.495 34.235 141.585 ;
        RECT 24.785 140.675 26.615 141.485 ;
        RECT 26.625 140.675 32.135 141.485 ;
        RECT 32.305 140.675 34.235 141.495 ;
        RECT 34.445 141.385 35.390 141.585 ;
        RECT 34.445 140.705 37.195 141.385 ;
        RECT 34.445 140.675 35.390 140.705 ;
        RECT 14.805 140.465 14.975 140.675 ;
        RECT 16.240 140.515 16.360 140.625 ;
        RECT 18.485 140.485 18.655 140.675 ;
        RECT 24.005 140.485 24.175 140.675 ;
        RECT 25.845 140.465 26.015 140.655 ;
        RECT 26.305 140.625 26.475 140.675 ;
        RECT 26.305 140.515 26.480 140.625 ;
        RECT 26.305 140.485 26.475 140.515 ;
        RECT 29.985 140.465 30.155 140.655 ;
        RECT 30.445 140.485 30.615 140.655 ;
        RECT 31.825 140.485 31.995 140.675 ;
        RECT 32.305 140.655 32.455 140.675 ;
        RECT 32.285 140.485 32.455 140.655 ;
        RECT 32.745 140.485 32.915 140.655 ;
        RECT 35.045 140.485 35.215 140.655 ;
        RECT 36.880 140.485 37.050 140.705 ;
        RECT 37.205 140.675 39.035 141.485 ;
        RECT 39.045 140.675 44.555 141.485 ;
        RECT 44.565 140.675 50.075 141.485 ;
        RECT 50.095 140.760 50.525 141.545 ;
        RECT 51.005 140.675 56.515 141.485 ;
        RECT 59.725 141.355 60.655 141.585 ;
        RECT 56.755 140.675 60.655 141.355 ;
        RECT 60.665 140.675 62.495 141.485 ;
        RECT 62.505 140.675 65.980 141.585 ;
        RECT 66.555 141.475 67.475 141.585 ;
        RECT 66.555 141.355 68.890 141.475 ;
        RECT 73.555 141.355 74.475 141.575 ;
        RECT 66.555 140.675 75.835 141.355 ;
        RECT 75.855 140.760 76.285 141.545 ;
        RECT 76.305 140.675 77.675 141.485 ;
        RECT 79.490 141.385 80.435 141.585 ;
        RECT 77.685 140.705 80.435 141.385 ;
        RECT 37.860 140.515 37.980 140.625 ;
        RECT 38.725 140.485 38.895 140.675 ;
        RECT 30.465 140.465 30.615 140.485 ;
        RECT 32.765 140.465 32.915 140.485 ;
        RECT 35.065 140.465 35.215 140.485 ;
        RECT 39.645 140.465 39.815 140.655 ;
        RECT 44.245 140.485 44.415 140.675 ;
        RECT 45.165 140.465 45.335 140.655 ;
        RECT 45.625 140.485 45.795 140.655 ;
        RECT 45.645 140.465 45.795 140.485 ;
        RECT 48.845 140.465 49.015 140.655 ;
        RECT 14.665 139.655 16.035 140.465 ;
        RECT 16.875 139.785 26.155 140.465 ;
        RECT 16.875 139.665 19.210 139.785 ;
        RECT 16.875 139.555 17.795 139.665 ;
        RECT 23.875 139.565 24.795 139.785 ;
        RECT 26.625 139.655 30.295 140.465 ;
        RECT 30.465 139.645 32.395 140.465 ;
        RECT 32.765 139.645 34.695 140.465 ;
        RECT 35.065 139.645 36.995 140.465 ;
        RECT 31.445 139.555 32.395 139.645 ;
        RECT 33.745 139.555 34.695 139.645 ;
        RECT 36.045 139.555 36.995 139.645 ;
        RECT 37.215 139.595 37.645 140.380 ;
        RECT 38.125 139.655 39.955 140.465 ;
        RECT 39.965 139.655 45.475 140.465 ;
        RECT 45.645 139.645 47.575 140.465 ;
        RECT 47.785 139.655 49.155 140.465 ;
        RECT 49.310 140.435 49.480 140.655 ;
        RECT 49.765 140.485 49.935 140.675 ;
        RECT 50.740 140.515 50.860 140.625 ;
        RECT 52.070 140.465 52.240 140.655 ;
        RECT 55.800 140.515 55.920 140.625 ;
        RECT 56.205 140.485 56.375 140.675 ;
        RECT 59.610 140.465 59.780 140.655 ;
        RECT 60.070 140.485 60.240 140.675 ;
        RECT 60.345 140.465 60.515 140.655 ;
        RECT 62.185 140.485 62.355 140.675 ;
        RECT 62.650 140.655 62.820 140.675 ;
        RECT 62.645 140.485 62.820 140.655 ;
        RECT 63.620 140.515 63.740 140.625 ;
        RECT 62.645 140.465 62.815 140.485 ;
        RECT 66.325 140.465 66.495 140.655 ;
        RECT 71.845 140.465 72.015 140.655 ;
        RECT 73.225 140.465 73.395 140.655 ;
        RECT 75.525 140.485 75.695 140.675 ;
        RECT 77.365 140.485 77.535 140.675 ;
        RECT 77.830 140.485 78.000 140.705 ;
        RECT 79.490 140.675 80.435 140.705 ;
        RECT 80.445 140.675 83.920 141.585 ;
        RECT 87.785 141.355 88.715 141.585 ;
        RECT 84.815 140.675 88.715 141.355 ;
        RECT 88.735 140.675 90.085 141.585 ;
        RECT 90.565 140.675 96.075 141.485 ;
        RECT 96.085 140.675 101.595 141.485 ;
        RECT 101.615 140.760 102.045 141.545 ;
        RECT 102.065 140.675 103.435 141.485 ;
        RECT 103.445 141.385 104.390 141.585 ;
        RECT 103.445 140.705 106.195 141.385 ;
        RECT 103.445 140.675 104.390 140.705 ;
        RECT 78.745 140.465 78.915 140.655 ;
        RECT 80.590 140.485 80.760 140.675 ;
        RECT 84.320 140.515 84.440 140.625 ;
        RECT 88.130 140.485 88.300 140.675 ;
        RECT 88.405 140.465 88.575 140.655 ;
        RECT 89.785 140.485 89.955 140.675 ;
        RECT 90.245 140.625 90.415 140.655 ;
        RECT 90.245 140.515 90.420 140.625 ;
        RECT 90.760 140.515 90.880 140.625 ;
        RECT 90.245 140.465 90.415 140.515 ;
        RECT 95.765 140.485 95.935 140.675 ;
        RECT 96.225 140.465 96.395 140.655 ;
        RECT 50.970 140.435 51.915 140.465 ;
        RECT 49.165 139.755 51.915 140.435 ;
        RECT 46.625 139.555 47.575 139.645 ;
        RECT 50.970 139.555 51.915 139.755 ;
        RECT 51.925 139.555 55.400 140.465 ;
        RECT 56.295 139.785 60.195 140.465 ;
        RECT 59.265 139.555 60.195 139.785 ;
        RECT 60.205 139.685 61.575 140.465 ;
        RECT 61.585 139.655 62.955 140.465 ;
        RECT 62.975 139.595 63.405 140.380 ;
        RECT 63.885 139.655 66.635 140.465 ;
        RECT 66.645 139.655 72.155 140.465 ;
        RECT 72.175 139.555 73.525 140.465 ;
        RECT 73.545 139.655 79.055 140.465 ;
        RECT 79.435 139.785 88.715 140.465 ;
        RECT 79.435 139.665 81.770 139.785 ;
        RECT 79.435 139.555 80.355 139.665 ;
        RECT 86.435 139.565 87.355 139.785 ;
        RECT 88.735 139.595 89.165 140.380 ;
        RECT 89.185 139.685 90.555 140.465 ;
        RECT 91.025 139.655 96.535 140.465 ;
        RECT 96.690 140.435 96.860 140.655 ;
        RECT 99.450 140.465 99.620 140.655 ;
        RECT 101.285 140.485 101.455 140.675 ;
        RECT 103.125 140.625 103.295 140.675 ;
        RECT 103.125 140.515 103.300 140.625 ;
        RECT 103.125 140.485 103.295 140.515 ;
        RECT 98.350 140.435 99.295 140.465 ;
        RECT 96.545 139.755 99.295 140.435 ;
        RECT 98.350 139.555 99.295 139.755 ;
        RECT 99.305 139.555 102.780 140.465 ;
        RECT 103.445 140.435 104.390 140.465 ;
        RECT 105.880 140.435 106.050 140.705 ;
        RECT 106.205 140.675 109.680 141.585 ;
        RECT 110.345 140.675 112.175 141.485 ;
        RECT 115.385 141.355 116.315 141.585 ;
        RECT 112.415 140.675 116.315 141.355 ;
        RECT 116.325 141.355 117.255 141.585 ;
        RECT 116.325 140.675 120.225 141.355 ;
        RECT 120.475 140.675 121.825 141.585 ;
        RECT 122.765 140.675 126.435 141.485 ;
        RECT 126.445 140.675 127.815 141.485 ;
        RECT 106.350 140.485 106.520 140.675 ;
        RECT 107.265 140.465 107.435 140.655 ;
        RECT 110.080 140.515 110.200 140.625 ;
        RECT 111.130 140.465 111.300 140.655 ;
        RECT 111.865 140.485 112.035 140.675 ;
        RECT 112.785 140.465 112.955 140.655 ;
        RECT 113.245 140.465 113.415 140.655 ;
        RECT 115.085 140.465 115.255 140.655 ;
        RECT 115.730 140.485 115.900 140.675 ;
        RECT 116.740 140.485 116.910 140.675 ;
        RECT 120.605 140.485 120.775 140.675 ;
        RECT 122.445 140.520 122.605 140.630 ;
        RECT 125.665 140.465 125.835 140.655 ;
        RECT 126.125 140.625 126.295 140.675 ;
        RECT 126.125 140.515 126.300 140.625 ;
        RECT 126.125 140.485 126.295 140.515 ;
        RECT 127.505 140.465 127.675 140.675 ;
        RECT 103.445 139.755 106.195 140.435 ;
        RECT 103.445 139.555 104.390 139.755 ;
        RECT 106.205 139.655 107.575 140.465 ;
        RECT 107.815 139.785 111.715 140.465 ;
        RECT 110.785 139.555 111.715 139.785 ;
        RECT 111.725 139.655 113.095 140.465 ;
        RECT 113.105 139.685 114.475 140.465 ;
        RECT 114.495 139.595 114.925 140.380 ;
        RECT 114.955 139.555 116.305 140.465 ;
        RECT 116.695 139.785 125.975 140.465 ;
        RECT 116.695 139.665 119.030 139.785 ;
        RECT 116.695 139.555 117.615 139.665 ;
        RECT 123.695 139.565 124.615 139.785 ;
        RECT 126.445 139.655 127.815 140.465 ;
      LAYER nwell ;
        RECT 14.470 136.435 128.010 139.265 ;
      LAYER pwell ;
        RECT 14.665 135.235 16.035 136.045 ;
        RECT 16.045 135.235 17.415 136.045 ;
        RECT 17.435 135.235 18.785 136.145 ;
        RECT 18.815 135.235 20.165 136.145 ;
        RECT 23.385 135.915 24.315 136.145 ;
        RECT 20.415 135.235 24.315 135.915 ;
        RECT 24.335 135.320 24.765 136.105 ;
        RECT 24.785 135.235 26.155 136.015 ;
        RECT 26.635 135.235 27.985 136.145 ;
        RECT 31.205 135.915 32.135 136.145 ;
        RECT 28.235 135.235 32.135 135.915 ;
        RECT 32.515 136.035 33.435 136.145 ;
        RECT 32.515 135.915 34.850 136.035 ;
        RECT 39.515 135.915 40.435 136.135 ;
        RECT 45.925 135.915 46.855 136.145 ;
        RECT 32.515 135.235 41.795 135.915 ;
        RECT 42.955 135.235 46.855 135.915 ;
        RECT 47.065 136.055 48.015 136.145 ;
        RECT 47.065 135.235 48.995 136.055 ;
        RECT 50.095 135.320 50.525 136.105 ;
        RECT 50.545 135.235 54.215 136.045 ;
        RECT 54.595 136.035 55.515 136.145 ;
        RECT 54.595 135.915 56.930 136.035 ;
        RECT 61.595 135.915 62.515 136.135 ;
        RECT 54.595 135.235 63.875 135.915 ;
        RECT 64.805 135.235 70.315 136.045 ;
        RECT 70.325 135.235 75.835 136.045 ;
        RECT 75.855 135.320 76.285 136.105 ;
        RECT 76.305 135.235 81.815 136.045 ;
        RECT 81.825 135.235 85.300 136.145 ;
        RECT 85.505 135.235 91.015 136.045 ;
        RECT 91.025 135.235 96.535 136.045 ;
        RECT 99.745 135.915 100.675 136.145 ;
        RECT 96.775 135.235 100.675 135.915 ;
        RECT 101.615 135.320 102.045 136.105 ;
        RECT 102.065 135.235 104.815 136.045 ;
        RECT 105.195 136.035 106.115 136.145 ;
        RECT 105.195 135.915 107.530 136.035 ;
        RECT 112.195 135.915 113.115 136.135 ;
        RECT 105.195 135.235 114.475 135.915 ;
        RECT 114.485 135.235 115.855 136.045 ;
        RECT 116.235 136.035 117.155 136.145 ;
        RECT 116.235 135.915 118.570 136.035 ;
        RECT 123.235 135.915 124.155 136.135 ;
        RECT 116.235 135.235 125.515 135.915 ;
        RECT 126.445 135.235 127.815 136.045 ;
        RECT 14.805 135.025 14.975 135.235 ;
        RECT 16.240 135.075 16.360 135.185 ;
        RECT 17.105 135.045 17.275 135.235 ;
        RECT 17.565 135.045 17.735 135.235 ;
        RECT 18.025 135.025 18.195 135.215 ;
        RECT 18.485 135.025 18.655 135.215 ;
        RECT 18.945 135.045 19.115 135.235 ;
        RECT 20.140 135.025 20.310 135.215 ;
        RECT 23.730 135.045 23.900 135.235 ;
        RECT 25.845 135.045 26.015 135.235 ;
        RECT 26.360 135.075 26.480 135.185 ;
        RECT 26.765 135.045 26.935 135.235 ;
        RECT 31.550 135.045 31.720 135.235 ;
        RECT 33.205 135.025 33.375 135.215 ;
        RECT 35.045 135.025 35.215 135.215 ;
        RECT 35.505 135.025 35.675 135.215 ;
        RECT 36.940 135.075 37.060 135.185 ;
        RECT 37.860 135.075 37.980 135.185 ;
        RECT 38.265 135.025 38.435 135.215 ;
        RECT 41.485 135.045 41.655 135.235 ;
        RECT 42.405 135.080 42.565 135.190 ;
        RECT 46.270 135.045 46.440 135.235 ;
        RECT 48.845 135.215 48.995 135.235 ;
        RECT 48.845 135.025 49.015 135.215 ;
        RECT 49.765 135.080 49.925 135.190 ;
        RECT 51.605 135.025 51.775 135.215 ;
        RECT 53.905 135.045 54.075 135.235 ;
        RECT 57.125 135.025 57.295 135.215 ;
        RECT 57.585 135.025 57.755 135.215 ;
        RECT 59.020 135.075 59.140 135.185 ;
        RECT 62.645 135.025 62.815 135.215 ;
        RECT 63.565 135.045 63.735 135.235 ;
        RECT 64.485 135.080 64.645 135.190 ;
        RECT 65.865 135.025 66.035 135.215 ;
        RECT 67.705 135.025 67.875 135.215 ;
        RECT 70.005 135.045 70.175 135.235 ;
        RECT 71.570 135.025 71.740 135.215 ;
        RECT 72.305 135.025 72.475 135.215 ;
        RECT 74.200 135.075 74.320 135.185 ;
        RECT 75.525 135.045 75.695 135.235 ;
        RECT 77.825 135.025 77.995 135.215 ;
        RECT 14.665 134.215 16.035 135.025 ;
        RECT 16.505 134.215 18.335 135.025 ;
        RECT 18.345 134.245 19.715 135.025 ;
        RECT 19.725 134.345 23.625 135.025 ;
        RECT 24.235 134.345 33.515 135.025 ;
        RECT 19.725 134.115 20.655 134.345 ;
        RECT 24.235 134.225 26.570 134.345 ;
        RECT 24.235 134.115 25.155 134.225 ;
        RECT 31.235 134.125 32.155 134.345 ;
        RECT 33.525 134.215 35.355 135.025 ;
        RECT 35.375 134.115 36.725 135.025 ;
        RECT 37.215 134.155 37.645 134.940 ;
        RECT 38.125 134.245 39.495 135.025 ;
        RECT 39.875 134.345 49.155 135.025 ;
        RECT 39.875 134.225 42.210 134.345 ;
        RECT 39.875 134.115 40.795 134.225 ;
        RECT 46.875 134.125 47.795 134.345 ;
        RECT 49.165 134.215 51.915 135.025 ;
        RECT 51.925 134.215 57.435 135.025 ;
        RECT 57.455 134.115 58.805 135.025 ;
        RECT 59.285 134.215 62.955 135.025 ;
        RECT 62.975 134.155 63.405 134.940 ;
        RECT 63.425 134.215 66.175 135.025 ;
        RECT 66.185 134.345 68.015 135.025 ;
        RECT 68.255 134.345 72.155 135.025 ;
        RECT 72.165 134.345 73.995 135.025 ;
        RECT 71.225 134.115 72.155 134.345 ;
        RECT 74.465 134.215 78.135 135.025 ;
        RECT 78.145 134.995 79.090 135.025 ;
        RECT 80.580 134.995 80.750 135.215 ;
        RECT 81.050 135.025 81.220 135.215 ;
        RECT 81.505 135.045 81.675 135.235 ;
        RECT 81.970 135.045 82.140 135.235 ;
        RECT 88.130 135.025 88.300 135.215 ;
        RECT 90.245 135.025 90.415 135.215 ;
        RECT 90.705 135.025 90.875 135.235 ;
        RECT 92.140 135.075 92.260 135.185 ;
        RECT 96.225 135.045 96.395 135.235 ;
        RECT 100.090 135.045 100.260 135.235 ;
        RECT 101.285 135.080 101.445 135.190 ;
        RECT 101.745 135.025 101.915 135.215 ;
        RECT 103.125 135.025 103.295 135.215 ;
        RECT 104.505 135.025 104.675 135.235 ;
        RECT 108.185 135.025 108.355 135.215 ;
        RECT 109.565 135.025 109.735 135.215 ;
        RECT 110.945 135.025 111.115 135.215 ;
        RECT 111.405 135.025 111.575 135.215 ;
        RECT 114.165 135.025 114.335 135.235 ;
        RECT 115.140 135.075 115.260 135.185 ;
        RECT 115.545 135.045 115.715 135.235 ;
        RECT 120.605 135.025 120.775 135.215 ;
        RECT 121.065 135.025 121.235 135.215 ;
        RECT 122.500 135.075 122.620 135.185 ;
        RECT 125.205 135.045 125.375 135.235 ;
        RECT 126.125 135.025 126.295 135.215 ;
        RECT 127.505 135.025 127.675 135.235 ;
        RECT 78.145 134.315 80.895 134.995 ;
        RECT 78.145 134.115 79.090 134.315 ;
        RECT 80.905 134.115 84.380 135.025 ;
        RECT 84.815 134.345 88.715 135.025 ;
        RECT 87.785 134.115 88.715 134.345 ;
        RECT 88.735 134.155 89.165 134.940 ;
        RECT 89.195 134.115 90.545 135.025 ;
        RECT 90.565 134.245 91.935 135.025 ;
        RECT 92.775 134.345 102.055 135.025 ;
        RECT 92.775 134.225 95.110 134.345 ;
        RECT 92.775 134.115 93.695 134.225 ;
        RECT 99.775 134.125 100.695 134.345 ;
        RECT 102.065 134.245 103.435 135.025 ;
        RECT 103.445 134.215 104.815 135.025 ;
        RECT 104.825 134.215 108.495 135.025 ;
        RECT 108.515 134.115 109.865 135.025 ;
        RECT 109.885 134.215 111.255 135.025 ;
        RECT 111.265 134.245 112.635 135.025 ;
        RECT 112.645 134.215 114.475 135.025 ;
        RECT 114.495 134.155 114.925 134.940 ;
        RECT 115.405 134.215 120.915 135.025 ;
        RECT 120.925 134.245 122.295 135.025 ;
        RECT 122.765 134.215 126.435 135.025 ;
        RECT 126.445 134.215 127.815 135.025 ;
      LAYER nwell ;
        RECT 14.470 130.995 128.010 133.825 ;
      LAYER pwell ;
        RECT 14.665 129.795 16.035 130.605 ;
        RECT 16.045 129.795 18.795 130.605 ;
        RECT 18.805 129.795 24.315 130.605 ;
        RECT 24.335 129.880 24.765 130.665 ;
        RECT 25.245 129.795 30.755 130.605 ;
        RECT 30.765 129.795 32.135 130.575 ;
        RECT 32.145 129.795 34.895 130.605 ;
        RECT 38.105 130.475 39.035 130.705 ;
        RECT 35.135 129.795 39.035 130.475 ;
        RECT 39.045 129.795 42.715 130.605 ;
        RECT 42.735 129.795 44.085 130.705 ;
        RECT 44.105 129.795 45.475 130.605 ;
        RECT 45.485 129.795 46.855 130.575 ;
        RECT 47.325 129.795 50.075 130.605 ;
        RECT 50.095 129.880 50.525 130.665 ;
        RECT 50.545 129.795 51.915 130.605 ;
        RECT 51.925 129.795 55.595 130.605 ;
        RECT 55.615 129.795 56.965 130.705 ;
        RECT 60.185 130.475 61.115 130.705 ;
        RECT 57.215 129.795 61.115 130.475 ;
        RECT 61.125 129.795 62.495 130.605 ;
        RECT 62.505 129.795 66.175 130.605 ;
        RECT 66.555 130.595 67.475 130.705 ;
        RECT 66.555 130.475 68.890 130.595 ;
        RECT 73.555 130.475 74.475 130.695 ;
        RECT 66.555 129.795 75.835 130.475 ;
        RECT 75.855 129.880 76.285 130.665 ;
        RECT 76.305 129.795 77.675 130.575 ;
        RECT 77.685 129.795 79.515 130.605 ;
        RECT 81.330 130.505 82.275 130.705 ;
        RECT 79.525 129.825 82.275 130.505 ;
        RECT 14.805 129.585 14.975 129.795 ;
        RECT 18.485 129.605 18.655 129.795 ;
        RECT 24.005 129.605 24.175 129.795 ;
        RECT 24.980 129.635 25.100 129.745 ;
        RECT 25.385 129.585 25.555 129.775 ;
        RECT 25.900 129.635 26.020 129.745 ;
        RECT 30.445 129.605 30.615 129.795 ;
        RECT 31.365 129.585 31.535 129.775 ;
        RECT 31.825 129.605 31.995 129.795 ;
        RECT 34.585 129.605 34.755 129.795 ;
        RECT 36.885 129.585 37.055 129.775 ;
        RECT 38.265 129.630 38.425 129.740 ;
        RECT 38.450 129.605 38.620 129.795 ;
        RECT 42.405 129.605 42.575 129.795 ;
        RECT 42.865 129.605 43.035 129.795 ;
        RECT 43.785 129.585 43.955 129.775 ;
        RECT 45.165 129.605 45.335 129.795 ;
        RECT 45.625 129.605 45.795 129.795 ;
        RECT 49.765 129.775 49.935 129.795 ;
        RECT 46.545 129.585 46.715 129.775 ;
        RECT 14.665 128.775 16.035 129.585 ;
        RECT 16.415 128.905 25.695 129.585 ;
        RECT 16.415 128.785 18.750 128.905 ;
        RECT 16.415 128.675 17.335 128.785 ;
        RECT 23.415 128.685 24.335 128.905 ;
        RECT 26.165 128.775 31.675 129.585 ;
        RECT 31.685 128.775 37.195 129.585 ;
        RECT 37.215 128.715 37.645 129.500 ;
        RECT 38.585 128.775 44.095 129.585 ;
        RECT 44.115 128.905 46.855 129.585 ;
        RECT 47.010 129.555 47.180 129.775 ;
        RECT 49.765 129.605 49.940 129.775 ;
        RECT 51.605 129.605 51.775 129.795 ;
        RECT 55.285 129.605 55.455 129.795 ;
        RECT 55.745 129.605 55.915 129.795 ;
        RECT 60.530 129.605 60.700 129.795 ;
        RECT 62.185 129.605 62.355 129.795 ;
        RECT 49.770 129.585 49.940 129.605 ;
        RECT 62.645 129.585 62.815 129.775 ;
        RECT 64.485 129.585 64.655 129.775 ;
        RECT 65.000 129.635 65.120 129.745 ;
        RECT 65.865 129.605 66.035 129.795 ;
        RECT 67.705 129.585 67.875 129.775 ;
        RECT 68.165 129.585 68.335 129.775 ;
        RECT 69.545 129.605 69.715 129.775 ;
        RECT 69.565 129.585 69.715 129.605 ;
        RECT 71.845 129.585 72.015 129.775 ;
        RECT 75.525 129.585 75.695 129.795 ;
        RECT 77.365 129.605 77.535 129.795 ;
        RECT 79.205 129.585 79.375 129.795 ;
        RECT 79.670 129.605 79.840 129.825 ;
        RECT 81.330 129.795 82.275 129.825 ;
        RECT 82.285 129.795 85.035 130.605 ;
        RECT 85.415 130.595 86.335 130.705 ;
        RECT 85.415 130.475 87.750 130.595 ;
        RECT 92.415 130.475 93.335 130.695 ;
        RECT 85.415 129.795 94.695 130.475 ;
        RECT 95.635 129.795 96.985 130.705 ;
        RECT 97.665 130.615 98.615 130.705 ;
        RECT 97.665 129.795 99.595 130.615 ;
        RECT 99.765 129.795 101.595 130.605 ;
        RECT 101.615 129.880 102.045 130.665 ;
        RECT 104.585 130.615 105.535 130.705 ;
        RECT 102.065 129.795 103.435 130.605 ;
        RECT 103.605 129.795 105.535 130.615 ;
        RECT 107.785 130.615 108.735 130.705 ;
        RECT 105.745 129.795 107.575 130.605 ;
        RECT 107.785 129.795 109.715 130.615 ;
        RECT 109.885 129.795 115.395 130.605 ;
        RECT 115.405 129.795 120.915 130.605 ;
        RECT 120.925 129.795 126.435 130.605 ;
        RECT 126.445 129.795 127.815 130.605 ;
        RECT 81.505 129.605 81.675 129.775 ;
        RECT 83.805 129.605 83.975 129.775 ;
        RECT 84.725 129.605 84.895 129.795 ;
        RECT 81.505 129.585 81.655 129.605 ;
        RECT 83.805 129.585 83.955 129.605 ;
        RECT 88.405 129.585 88.575 129.775 ;
        RECT 90.245 129.585 90.415 129.775 ;
        RECT 93.925 129.585 94.095 129.775 ;
        RECT 94.385 129.605 94.555 129.795 ;
        RECT 95.305 129.640 95.465 129.750 ;
        RECT 95.765 129.605 95.935 129.795 ;
        RECT 99.445 129.775 99.595 129.795 ;
        RECT 97.200 129.635 97.320 129.745 ;
        RECT 99.445 129.585 99.615 129.775 ;
        RECT 101.285 129.605 101.455 129.795 ;
        RECT 103.125 129.605 103.295 129.795 ;
        RECT 103.605 129.775 103.755 129.795 ;
        RECT 103.585 129.605 103.755 129.775 ;
        RECT 104.965 129.585 105.135 129.775 ;
        RECT 107.265 129.605 107.435 129.795 ;
        RECT 109.565 129.775 109.715 129.795 ;
        RECT 109.565 129.605 109.735 129.775 ;
        RECT 111.865 129.605 112.035 129.775 ;
        RECT 112.380 129.635 112.500 129.745 ;
        RECT 107.265 129.585 107.415 129.605 ;
        RECT 109.565 129.585 109.715 129.605 ;
        RECT 111.865 129.585 112.015 129.605 ;
        RECT 114.165 129.585 114.335 129.775 ;
        RECT 115.085 129.605 115.255 129.795 ;
        RECT 118.490 129.585 118.660 129.775 ;
        RECT 120.605 129.585 120.775 129.795 ;
        RECT 126.125 129.585 126.295 129.795 ;
        RECT 127.505 129.585 127.675 129.795 ;
        RECT 48.670 129.555 49.615 129.585 ;
        RECT 46.865 128.875 49.615 129.555 ;
        RECT 48.670 128.675 49.615 128.875 ;
        RECT 49.625 128.675 53.100 129.585 ;
        RECT 53.675 128.905 62.955 129.585 ;
        RECT 53.675 128.785 56.010 128.905 ;
        RECT 53.675 128.675 54.595 128.785 ;
        RECT 60.675 128.685 61.595 128.905 ;
        RECT 62.975 128.715 63.405 129.500 ;
        RECT 63.425 128.805 64.795 129.585 ;
        RECT 65.265 128.775 68.015 129.585 ;
        RECT 68.035 128.675 69.385 129.585 ;
        RECT 69.565 128.765 71.495 129.585 ;
        RECT 71.705 128.905 74.445 129.585 ;
        RECT 74.465 128.775 75.835 129.585 ;
        RECT 75.845 128.775 79.515 129.585 ;
        RECT 70.545 128.675 71.495 128.765 ;
        RECT 79.725 128.765 81.655 129.585 ;
        RECT 82.025 128.765 83.955 129.585 ;
        RECT 85.045 128.775 88.715 129.585 ;
        RECT 79.725 128.675 80.675 128.765 ;
        RECT 82.025 128.675 82.975 128.765 ;
        RECT 88.735 128.715 89.165 129.500 ;
        RECT 89.185 128.775 90.555 129.585 ;
        RECT 90.565 128.775 94.235 129.585 ;
        RECT 94.245 128.775 99.755 129.585 ;
        RECT 99.765 128.775 105.275 129.585 ;
        RECT 105.485 128.765 107.415 129.585 ;
        RECT 107.785 128.765 109.715 129.585 ;
        RECT 110.085 128.765 112.015 129.585 ;
        RECT 112.645 128.775 114.475 129.585 ;
        RECT 105.485 128.675 106.435 128.765 ;
        RECT 107.785 128.675 108.735 128.765 ;
        RECT 110.085 128.675 111.035 128.765 ;
        RECT 114.495 128.715 114.925 129.500 ;
        RECT 115.175 128.905 119.075 129.585 ;
        RECT 118.145 128.675 119.075 128.905 ;
        RECT 119.085 128.775 120.915 129.585 ;
        RECT 120.925 128.775 126.435 129.585 ;
        RECT 126.445 128.775 127.815 129.585 ;
      LAYER nwell ;
        RECT 14.470 125.555 128.010 128.385 ;
      LAYER pwell ;
        RECT 14.665 124.355 16.035 125.165 ;
        RECT 16.045 124.355 18.795 125.165 ;
        RECT 18.805 124.355 24.315 125.165 ;
        RECT 24.335 124.440 24.765 125.225 ;
        RECT 25.705 124.355 29.375 125.165 ;
        RECT 29.385 124.355 30.755 125.135 ;
        RECT 30.775 124.355 33.515 125.035 ;
        RECT 34.445 124.355 38.115 125.165 ;
        RECT 38.125 125.065 39.070 125.265 ;
        RECT 40.885 125.065 41.830 125.265 ;
        RECT 45.450 125.065 46.395 125.265 ;
        RECT 38.125 124.385 40.875 125.065 ;
        RECT 40.885 124.385 43.635 125.065 ;
        RECT 43.645 124.385 46.395 125.065 ;
        RECT 38.125 124.355 39.070 124.385 ;
        RECT 14.805 124.145 14.975 124.355 ;
        RECT 16.240 124.195 16.360 124.305 ;
        RECT 18.485 124.165 18.655 124.355 ;
        RECT 21.705 124.145 21.875 124.335 ;
        RECT 22.165 124.145 22.335 124.335 ;
        RECT 24.005 124.165 24.175 124.355 ;
        RECT 25.385 124.200 25.545 124.310 ;
        RECT 29.065 124.165 29.235 124.355 ;
        RECT 29.525 124.165 29.695 124.355 ;
        RECT 32.745 124.145 32.915 124.335 ;
        RECT 33.205 124.165 33.375 124.355 ;
        RECT 33.480 124.145 33.650 124.335 ;
        RECT 34.125 124.200 34.285 124.310 ;
        RECT 37.805 124.165 37.975 124.355 ;
        RECT 40.105 124.165 40.275 124.335 ;
        RECT 40.560 124.165 40.730 124.385 ;
        RECT 40.885 124.355 41.830 124.385 ;
        RECT 42.405 124.165 42.575 124.335 ;
        RECT 43.320 124.165 43.490 124.385 ;
        RECT 43.790 124.165 43.960 124.385 ;
        RECT 45.450 124.355 46.395 124.385 ;
        RECT 46.405 124.355 49.880 125.265 ;
        RECT 50.095 124.440 50.525 125.225 ;
        RECT 50.545 124.355 54.020 125.265 ;
        RECT 57.425 125.035 58.355 125.265 ;
        RECT 54.455 124.355 58.355 125.035 ;
        RECT 58.735 125.155 59.655 125.265 ;
        RECT 58.735 125.035 61.070 125.155 ;
        RECT 65.735 125.035 66.655 125.255 ;
        RECT 58.735 124.355 68.015 125.035 ;
        RECT 68.485 124.355 70.315 125.165 ;
        RECT 70.325 124.355 75.835 125.165 ;
        RECT 75.855 124.440 76.285 125.225 ;
        RECT 78.365 125.175 79.315 125.265 ;
        RECT 77.385 124.355 79.315 125.175 ;
        RECT 79.525 124.355 81.355 125.165 ;
        RECT 84.565 125.035 85.495 125.265 ;
        RECT 81.595 124.355 85.495 125.035 ;
        RECT 85.705 125.175 86.655 125.265 ;
        RECT 85.705 124.355 87.635 125.175 ;
        RECT 88.265 124.355 91.935 125.165 ;
        RECT 91.945 124.355 97.455 125.165 ;
        RECT 100.665 125.035 101.595 125.265 ;
        RECT 97.695 124.355 101.595 125.035 ;
        RECT 101.615 124.440 102.045 125.225 ;
        RECT 102.065 124.355 103.895 125.165 ;
        RECT 103.915 124.355 105.265 125.265 ;
        RECT 108.485 125.035 109.415 125.265 ;
        RECT 105.515 124.355 109.415 125.035 ;
        RECT 109.885 124.355 112.635 125.165 ;
        RECT 112.655 124.355 114.005 125.265 ;
        RECT 114.395 125.155 115.315 125.265 ;
        RECT 114.395 125.035 116.730 125.155 ;
        RECT 121.395 125.035 122.315 125.255 ;
        RECT 114.395 124.355 123.675 125.035 ;
        RECT 123.685 124.355 126.435 125.165 ;
        RECT 126.445 124.355 127.815 125.165 ;
        RECT 44.705 124.165 44.875 124.335 ;
        RECT 46.550 124.165 46.720 124.355 ;
        RECT 47.060 124.195 47.180 124.305 ;
        RECT 50.690 124.165 50.860 124.355 ;
        RECT 37.825 124.145 37.975 124.165 ;
        RECT 40.125 124.145 40.275 124.165 ;
        RECT 42.425 124.145 42.575 124.165 ;
        RECT 44.725 124.145 44.875 124.165 ;
        RECT 56.205 124.145 56.375 124.335 ;
        RECT 57.125 124.190 57.285 124.300 ;
        RECT 57.770 124.165 57.940 124.355 ;
        RECT 60.805 124.145 60.975 124.335 ;
        RECT 61.265 124.145 61.435 124.335 ;
        RECT 62.700 124.195 62.820 124.305 ;
        RECT 63.620 124.195 63.740 124.305 ;
        RECT 64.025 124.145 64.195 124.335 ;
        RECT 65.460 124.195 65.580 124.305 ;
        RECT 67.245 124.145 67.415 124.335 ;
        RECT 67.705 124.165 67.875 124.355 ;
        RECT 68.220 124.195 68.340 124.305 ;
        RECT 70.005 124.165 70.175 124.355 ;
        RECT 72.765 124.145 72.935 124.335 ;
        RECT 74.145 124.145 74.315 124.335 ;
        RECT 75.065 124.190 75.225 124.300 ;
        RECT 75.525 124.165 75.695 124.355 ;
        RECT 77.385 124.335 77.535 124.355 ;
        RECT 76.905 124.200 77.065 124.310 ;
        RECT 77.365 124.165 77.535 124.335 ;
        RECT 78.930 124.145 79.100 124.335 ;
        RECT 81.045 124.165 81.215 124.355 ;
        RECT 84.910 124.165 85.080 124.355 ;
        RECT 87.485 124.335 87.635 124.355 ;
        RECT 87.485 124.165 87.655 124.335 ;
        RECT 88.000 124.195 88.120 124.305 ;
        RECT 88.405 124.145 88.575 124.335 ;
        RECT 90.705 124.145 90.875 124.335 ;
        RECT 91.165 124.145 91.335 124.335 ;
        RECT 91.625 124.165 91.795 124.355 ;
        RECT 97.145 124.165 97.315 124.355 ;
        RECT 101.010 124.165 101.180 124.355 ;
        RECT 101.745 124.145 101.915 124.335 ;
        RECT 103.585 124.165 103.755 124.355 ;
        RECT 104.045 124.165 104.215 124.355 ;
        RECT 108.830 124.165 109.000 124.355 ;
        RECT 109.620 124.195 109.740 124.305 ;
        RECT 111.405 124.145 111.575 124.335 ;
        RECT 112.325 124.165 112.495 124.355 ;
        RECT 112.785 124.145 112.955 124.355 ;
        RECT 113.245 124.145 113.415 124.335 ;
        RECT 115.545 124.190 115.705 124.300 ;
        RECT 123.365 124.165 123.535 124.355 ;
        RECT 125.205 124.145 125.375 124.335 ;
        RECT 126.125 124.165 126.295 124.355 ;
        RECT 127.505 124.145 127.675 124.355 ;
        RECT 14.665 123.335 16.035 124.145 ;
        RECT 16.505 123.335 22.015 124.145 ;
        RECT 22.025 123.365 23.395 124.145 ;
        RECT 23.775 123.465 33.055 124.145 ;
        RECT 33.065 123.465 36.965 124.145 ;
        RECT 23.775 123.345 26.110 123.465 ;
        RECT 23.775 123.235 24.695 123.345 ;
        RECT 30.775 123.245 31.695 123.465 ;
        RECT 33.065 123.235 33.995 123.465 ;
        RECT 37.215 123.275 37.645 124.060 ;
        RECT 37.825 123.325 39.755 124.145 ;
        RECT 40.125 123.325 42.055 124.145 ;
        RECT 42.425 123.325 44.355 124.145 ;
        RECT 44.725 123.325 46.655 124.145 ;
        RECT 47.410 123.465 56.515 124.145 ;
        RECT 57.445 123.335 61.115 124.145 ;
        RECT 38.805 123.235 39.755 123.325 ;
        RECT 41.105 123.235 42.055 123.325 ;
        RECT 43.405 123.235 44.355 123.325 ;
        RECT 45.705 123.235 46.655 123.325 ;
        RECT 61.135 123.235 62.485 124.145 ;
        RECT 62.975 123.275 63.405 124.060 ;
        RECT 63.885 123.365 65.255 124.145 ;
        RECT 65.725 123.335 67.555 124.145 ;
        RECT 67.565 123.335 73.075 124.145 ;
        RECT 73.095 123.235 74.445 124.145 ;
        RECT 75.615 123.465 79.515 124.145 ;
        RECT 79.610 123.465 88.715 124.145 ;
        RECT 78.585 123.235 79.515 123.465 ;
        RECT 88.735 123.275 89.165 124.060 ;
        RECT 89.185 123.335 91.015 124.145 ;
        RECT 91.035 123.235 92.385 124.145 ;
        RECT 92.775 123.465 102.055 124.145 ;
        RECT 102.435 123.465 111.715 124.145 ;
        RECT 92.775 123.345 95.110 123.465 ;
        RECT 92.775 123.235 93.695 123.345 ;
        RECT 99.775 123.245 100.695 123.465 ;
        RECT 102.435 123.345 104.770 123.465 ;
        RECT 102.435 123.235 103.355 123.345 ;
        RECT 109.435 123.245 110.355 123.465 ;
        RECT 111.725 123.335 113.095 124.145 ;
        RECT 113.115 123.235 114.465 124.145 ;
        RECT 114.495 123.275 114.925 124.060 ;
        RECT 116.235 123.465 125.515 124.145 ;
        RECT 116.235 123.345 118.570 123.465 ;
        RECT 116.235 123.235 117.155 123.345 ;
        RECT 123.235 123.245 124.155 123.465 ;
        RECT 126.445 123.335 127.815 124.145 ;
      LAYER nwell ;
        RECT 14.470 120.115 128.010 122.945 ;
      LAYER pwell ;
        RECT 14.665 118.915 16.035 119.725 ;
        RECT 16.055 118.915 17.405 119.825 ;
        RECT 17.435 118.915 18.785 119.825 ;
        RECT 18.815 118.915 20.165 119.825 ;
        RECT 23.385 119.595 24.315 119.825 ;
        RECT 20.415 118.915 24.315 119.595 ;
        RECT 24.335 119.000 24.765 119.785 ;
        RECT 24.785 119.595 25.715 119.825 ;
        RECT 29.295 119.715 30.215 119.825 ;
        RECT 29.295 119.595 31.630 119.715 ;
        RECT 36.295 119.595 37.215 119.815 ;
        RECT 24.785 118.915 28.685 119.595 ;
        RECT 29.295 118.915 38.575 119.595 ;
        RECT 38.585 118.915 41.335 119.725 ;
        RECT 44.545 119.595 45.475 119.825 ;
        RECT 41.575 118.915 45.475 119.595 ;
        RECT 45.485 118.915 48.235 119.725 ;
        RECT 48.245 118.915 49.610 119.595 ;
        RECT 50.095 119.000 50.525 119.785 ;
        RECT 50.545 118.915 54.020 119.825 ;
        RECT 54.235 118.915 55.585 119.825 ;
        RECT 58.805 119.595 59.735 119.825 ;
        RECT 55.835 118.915 59.735 119.595 ;
        RECT 60.665 118.915 66.175 119.725 ;
        RECT 67.545 119.595 68.465 119.815 ;
        RECT 74.545 119.715 75.465 119.825 ;
        RECT 73.130 119.595 75.465 119.715 ;
        RECT 66.185 118.915 75.465 119.595 ;
        RECT 75.855 119.000 76.285 119.785 ;
        RECT 76.675 119.715 77.595 119.825 ;
        RECT 76.675 119.595 79.010 119.715 ;
        RECT 83.675 119.595 84.595 119.815 ;
        RECT 88.175 119.715 89.095 119.825 ;
        RECT 76.675 118.915 85.955 119.595 ;
        RECT 85.965 118.915 87.335 119.695 ;
        RECT 88.175 119.595 90.510 119.715 ;
        RECT 95.175 119.595 96.095 119.815 ;
        RECT 88.175 118.915 97.455 119.595 ;
        RECT 97.475 118.915 98.825 119.825 ;
        RECT 98.845 118.915 100.215 119.695 ;
        RECT 100.225 118.915 101.595 119.695 ;
        RECT 101.615 119.000 102.045 119.785 ;
        RECT 102.065 118.915 111.170 119.595 ;
        RECT 111.275 118.915 114.015 119.595 ;
        RECT 114.025 118.915 115.395 119.725 ;
        RECT 118.605 119.595 119.535 119.825 ;
        RECT 115.635 118.915 119.535 119.595 ;
        RECT 119.545 118.915 120.915 119.695 ;
        RECT 120.925 118.915 122.295 119.695 ;
        RECT 122.765 118.915 126.435 119.725 ;
        RECT 126.445 118.915 127.815 119.725 ;
        RECT 14.805 118.705 14.975 118.915 ;
        RECT 17.105 118.725 17.275 118.915 ;
        RECT 17.565 118.705 17.735 118.915 ;
        RECT 18.945 118.725 19.115 118.915 ;
        RECT 23.730 118.725 23.900 118.915 ;
        RECT 25.200 118.725 25.370 118.915 ;
        RECT 27.225 118.705 27.395 118.895 ;
        RECT 36.425 118.705 36.595 118.895 ;
        RECT 36.940 118.755 37.060 118.865 ;
        RECT 38.265 118.725 38.435 118.915 ;
        RECT 41.025 118.725 41.195 118.915 ;
        RECT 44.890 118.725 45.060 118.915 ;
        RECT 47.005 118.705 47.175 118.895 ;
        RECT 47.925 118.725 48.095 118.915 ;
        RECT 49.760 118.725 49.935 118.895 ;
        RECT 50.690 118.725 50.860 118.915 ;
        RECT 49.760 118.705 49.930 118.725 ;
        RECT 51.145 118.705 51.315 118.895 ;
        RECT 54.365 118.725 54.535 118.915 ;
        RECT 59.150 118.725 59.320 118.915 ;
        RECT 60.345 118.760 60.505 118.870 ;
        RECT 60.805 118.705 60.975 118.895 ;
        RECT 62.185 118.705 62.355 118.895 ;
        RECT 62.700 118.755 62.820 118.865 ;
        RECT 63.620 118.755 63.740 118.865 ;
        RECT 65.405 118.705 65.575 118.895 ;
        RECT 65.865 118.725 66.035 118.915 ;
        RECT 66.325 118.725 66.495 118.915 ;
        RECT 69.270 118.705 69.440 118.895 ;
        RECT 70.060 118.755 70.180 118.865 ;
        RECT 70.465 118.705 70.635 118.895 ;
        RECT 72.305 118.750 72.465 118.860 ;
        RECT 75.985 118.705 76.155 118.895 ;
        RECT 76.445 118.705 76.615 118.895 ;
        RECT 78.745 118.705 78.915 118.895 ;
        RECT 79.205 118.705 79.375 118.895 ;
        RECT 85.645 118.725 85.815 118.915 ;
        RECT 87.025 118.725 87.195 118.915 ;
        RECT 87.540 118.755 87.660 118.865 ;
        RECT 90.245 118.705 90.415 118.895 ;
        RECT 91.165 118.750 91.325 118.860 ;
        RECT 95.030 118.705 95.200 118.895 ;
        RECT 95.820 118.755 95.940 118.865 ;
        RECT 97.145 118.725 97.315 118.915 ;
        RECT 97.605 118.705 97.775 118.915 ;
        RECT 99.905 118.725 100.075 118.915 ;
        RECT 101.285 118.725 101.455 118.915 ;
        RECT 102.205 118.725 102.375 118.915 ;
        RECT 103.125 118.705 103.295 118.895 ;
        RECT 103.585 118.705 103.755 118.895 ;
        RECT 108.370 118.705 108.540 118.895 ;
        RECT 109.105 118.705 109.275 118.895 ;
        RECT 113.705 118.725 113.875 118.915 ;
        RECT 113.890 118.705 114.060 118.895 ;
        RECT 115.085 118.725 115.255 118.915 ;
        RECT 116.005 118.705 116.175 118.895 ;
        RECT 117.385 118.705 117.555 118.895 ;
        RECT 118.305 118.750 118.465 118.860 ;
        RECT 118.765 118.705 118.935 118.895 ;
        RECT 118.950 118.725 119.120 118.915 ;
        RECT 119.685 118.725 119.855 118.915 ;
        RECT 120.605 118.750 120.765 118.860 ;
        RECT 121.065 118.725 121.235 118.915 ;
        RECT 122.500 118.755 122.620 118.865 ;
        RECT 126.125 118.705 126.295 118.915 ;
        RECT 127.505 118.705 127.675 118.915 ;
        RECT 14.665 117.895 16.035 118.705 ;
        RECT 16.045 117.895 17.875 118.705 ;
        RECT 18.255 118.025 27.535 118.705 ;
        RECT 27.630 118.025 36.735 118.705 ;
        RECT 18.255 117.905 20.590 118.025 ;
        RECT 18.255 117.795 19.175 117.905 ;
        RECT 25.255 117.805 26.175 118.025 ;
        RECT 37.215 117.835 37.645 118.620 ;
        RECT 38.035 118.025 47.315 118.705 ;
        RECT 38.035 117.905 40.370 118.025 ;
        RECT 38.035 117.795 38.955 117.905 ;
        RECT 45.035 117.805 45.955 118.025 ;
        RECT 47.465 117.795 50.075 118.705 ;
        RECT 50.085 117.895 51.455 118.705 ;
        RECT 51.835 118.025 61.115 118.705 ;
        RECT 51.835 117.905 54.170 118.025 ;
        RECT 51.835 117.795 52.755 117.905 ;
        RECT 58.835 117.805 59.755 118.025 ;
        RECT 61.125 117.925 62.495 118.705 ;
        RECT 62.975 117.835 63.405 118.620 ;
        RECT 63.885 117.895 65.715 118.705 ;
        RECT 65.955 118.025 69.855 118.705 ;
        RECT 68.925 117.795 69.855 118.025 ;
        RECT 70.325 117.925 71.695 118.705 ;
        RECT 72.625 117.895 76.295 118.705 ;
        RECT 76.315 117.795 77.665 118.705 ;
        RECT 77.685 117.925 79.055 118.705 ;
        RECT 79.065 118.025 88.345 118.705 ;
        RECT 80.425 117.805 81.345 118.025 ;
        RECT 86.010 117.905 88.345 118.025 ;
        RECT 87.425 117.795 88.345 117.905 ;
        RECT 88.735 117.835 89.165 118.620 ;
        RECT 89.195 117.795 90.545 118.705 ;
        RECT 91.715 118.025 95.615 118.705 ;
        RECT 94.685 117.795 95.615 118.025 ;
        RECT 96.085 117.895 97.915 118.705 ;
        RECT 97.925 117.895 103.435 118.705 ;
        RECT 103.455 117.795 104.805 118.705 ;
        RECT 105.055 118.025 108.955 118.705 ;
        RECT 108.025 117.795 108.955 118.025 ;
        RECT 108.965 117.925 110.335 118.705 ;
        RECT 110.575 118.025 114.475 118.705 ;
        RECT 113.545 117.795 114.475 118.025 ;
        RECT 114.495 117.835 114.925 118.620 ;
        RECT 114.945 117.895 116.315 118.705 ;
        RECT 116.335 117.795 117.685 118.705 ;
        RECT 118.625 117.925 119.995 118.705 ;
        RECT 120.925 117.895 126.435 118.705 ;
        RECT 126.445 117.895 127.815 118.705 ;
      LAYER nwell ;
        RECT 14.470 114.675 128.010 117.505 ;
      LAYER pwell ;
        RECT 14.665 113.475 16.035 114.285 ;
        RECT 16.045 113.475 17.415 114.285 ;
        RECT 17.425 113.475 22.935 114.285 ;
        RECT 22.945 113.475 24.315 114.255 ;
        RECT 24.335 113.560 24.765 114.345 ;
        RECT 25.245 113.475 27.995 114.285 ;
        RECT 28.015 113.475 29.365 114.385 ;
        RECT 29.385 114.155 30.315 114.385 ;
        RECT 29.385 113.475 33.285 114.155 ;
        RECT 34.445 113.475 35.815 114.255 ;
        RECT 35.835 113.475 37.185 114.385 ;
        RECT 37.205 113.475 39.035 114.285 ;
        RECT 39.045 113.475 44.555 114.285 ;
        RECT 44.565 113.475 45.935 114.255 ;
        RECT 46.405 113.475 50.075 114.285 ;
        RECT 50.095 113.560 50.525 114.345 ;
        RECT 50.545 113.475 51.915 114.285 ;
        RECT 51.925 113.475 55.595 114.285 ;
        RECT 58.805 114.155 59.735 114.385 ;
        RECT 55.835 113.475 59.735 114.155 ;
        RECT 59.745 113.475 65.255 114.285 ;
        RECT 65.635 114.275 66.555 114.385 ;
        RECT 65.635 114.155 67.970 114.275 ;
        RECT 72.635 114.155 73.555 114.375 ;
        RECT 65.635 113.475 74.915 114.155 ;
        RECT 75.855 113.560 76.285 114.345 ;
        RECT 76.765 113.475 79.515 114.285 ;
        RECT 79.525 113.475 85.035 114.285 ;
        RECT 88.245 114.155 89.175 114.385 ;
        RECT 85.275 113.475 89.175 114.155 ;
        RECT 89.185 113.475 90.555 114.255 ;
        RECT 90.565 113.475 96.075 114.285 ;
        RECT 96.085 113.475 101.595 114.285 ;
        RECT 101.615 113.560 102.045 114.345 ;
        RECT 102.895 114.275 103.815 114.385 ;
        RECT 102.895 114.155 105.230 114.275 ;
        RECT 109.895 114.155 110.815 114.375 ;
        RECT 113.015 114.275 113.935 114.385 ;
        RECT 113.015 114.155 115.350 114.275 ;
        RECT 120.015 114.155 120.935 114.375 ;
        RECT 102.895 113.475 112.175 114.155 ;
        RECT 113.015 113.475 122.295 114.155 ;
        RECT 122.765 113.475 126.435 114.285 ;
        RECT 126.445 113.475 127.815 114.285 ;
        RECT 14.805 113.265 14.975 113.475 ;
        RECT 16.645 113.310 16.805 113.420 ;
        RECT 17.105 113.285 17.275 113.475 ;
        RECT 20.325 113.265 20.495 113.455 ;
        RECT 22.625 113.285 22.795 113.475 ;
        RECT 23.085 113.285 23.255 113.475 ;
        RECT 24.980 113.315 25.100 113.425 ;
        RECT 27.685 113.285 27.855 113.475 ;
        RECT 28.145 113.285 28.315 113.475 ;
        RECT 29.525 113.265 29.695 113.455 ;
        RECT 29.800 113.285 29.970 113.475 ;
        RECT 31.365 113.265 31.535 113.455 ;
        RECT 34.125 113.320 34.285 113.430 ;
        RECT 34.585 113.285 34.755 113.475 ;
        RECT 35.965 113.285 36.135 113.475 ;
        RECT 36.885 113.265 37.055 113.455 ;
        RECT 37.860 113.315 37.980 113.425 ;
        RECT 38.725 113.285 38.895 113.475 ;
        RECT 41.485 113.265 41.655 113.455 ;
        RECT 41.945 113.265 42.115 113.455 ;
        RECT 43.380 113.315 43.500 113.425 ;
        RECT 44.245 113.285 44.415 113.475 ;
        RECT 44.705 113.285 44.875 113.475 ;
        RECT 46.140 113.315 46.260 113.425 ;
        RECT 47.005 113.265 47.175 113.455 ;
        RECT 49.765 113.285 49.935 113.475 ;
        RECT 51.605 113.285 51.775 113.475 ;
        RECT 52.525 113.265 52.695 113.455 ;
        RECT 55.285 113.285 55.455 113.475 ;
        RECT 59.150 113.285 59.320 113.475 ;
        RECT 62.185 113.265 62.355 113.455 ;
        RECT 62.700 113.315 62.820 113.425 ;
        RECT 64.945 113.285 65.115 113.475 ;
        RECT 68.625 113.265 68.795 113.455 ;
        RECT 70.005 113.265 70.175 113.455 ;
        RECT 71.845 113.265 72.015 113.455 ;
        RECT 74.605 113.285 74.775 113.475 ;
        RECT 75.525 113.320 75.685 113.430 ;
        RECT 76.500 113.315 76.620 113.425 ;
        RECT 77.365 113.265 77.535 113.455 ;
        RECT 79.205 113.285 79.375 113.475 ;
        RECT 82.885 113.265 83.055 113.455 ;
        RECT 84.725 113.285 84.895 113.475 ;
        RECT 88.405 113.265 88.575 113.455 ;
        RECT 88.590 113.285 88.760 113.475 ;
        RECT 89.380 113.315 89.500 113.425 ;
        RECT 90.245 113.285 90.415 113.475 ;
        RECT 93.005 113.265 93.175 113.455 ;
        RECT 95.765 113.285 95.935 113.475 ;
        RECT 98.525 113.265 98.695 113.455 ;
        RECT 98.985 113.265 99.155 113.455 ;
        RECT 101.285 113.285 101.455 113.475 ;
        RECT 102.260 113.315 102.380 113.425 ;
        RECT 102.665 113.265 102.835 113.455 ;
        RECT 108.185 113.265 108.355 113.455 ;
        RECT 108.645 113.265 108.815 113.455 ;
        RECT 110.485 113.310 110.645 113.420 ;
        RECT 111.865 113.285 112.035 113.475 ;
        RECT 112.380 113.315 112.500 113.425 ;
        RECT 114.165 113.265 114.335 113.455 ;
        RECT 115.140 113.315 115.260 113.425 ;
        RECT 120.605 113.265 120.775 113.455 ;
        RECT 121.065 113.265 121.235 113.455 ;
        RECT 121.985 113.285 122.155 113.475 ;
        RECT 122.500 113.315 122.620 113.425 ;
        RECT 123.365 113.265 123.535 113.455 ;
        RECT 126.125 113.265 126.295 113.475 ;
        RECT 127.505 113.265 127.675 113.475 ;
        RECT 14.665 112.455 16.035 113.265 ;
        RECT 16.965 112.455 20.635 113.265 ;
        RECT 20.645 112.585 29.835 113.265 ;
        RECT 20.645 112.355 21.565 112.585 ;
        RECT 24.395 112.365 25.325 112.585 ;
        RECT 29.845 112.455 31.675 113.265 ;
        RECT 31.685 112.455 37.195 113.265 ;
        RECT 37.215 112.395 37.645 113.180 ;
        RECT 38.125 112.455 41.795 113.265 ;
        RECT 41.805 112.485 43.175 113.265 ;
        RECT 43.645 112.455 47.315 113.265 ;
        RECT 47.325 112.455 52.835 113.265 ;
        RECT 53.215 112.585 62.495 113.265 ;
        RECT 53.215 112.465 55.550 112.585 ;
        RECT 53.215 112.355 54.135 112.465 ;
        RECT 60.215 112.365 61.135 112.585 ;
        RECT 62.975 112.395 63.405 113.180 ;
        RECT 63.425 112.455 68.935 113.265 ;
        RECT 68.955 112.355 70.305 113.265 ;
        RECT 70.325 112.455 72.155 113.265 ;
        RECT 72.165 112.455 77.675 113.265 ;
        RECT 77.685 112.455 83.195 113.265 ;
        RECT 83.205 112.455 88.715 113.265 ;
        RECT 88.735 112.395 89.165 113.180 ;
        RECT 89.645 112.455 93.315 113.265 ;
        RECT 93.325 112.455 98.835 113.265 ;
        RECT 98.845 112.485 100.215 113.265 ;
        RECT 100.225 112.455 102.975 113.265 ;
        RECT 102.985 112.455 108.495 113.265 ;
        RECT 108.505 112.485 109.875 113.265 ;
        RECT 110.805 112.455 114.475 113.265 ;
        RECT 114.495 112.395 114.925 113.180 ;
        RECT 115.405 112.455 120.915 113.265 ;
        RECT 120.925 112.485 122.295 113.265 ;
        RECT 122.305 112.485 123.675 113.265 ;
        RECT 123.685 112.455 126.435 113.265 ;
        RECT 126.445 112.455 127.815 113.265 ;
      LAYER nwell ;
        RECT 14.470 109.235 128.010 112.065 ;
      LAYER pwell ;
        RECT 14.665 108.035 16.035 108.845 ;
        RECT 16.045 108.035 17.415 108.845 ;
        RECT 17.425 108.035 22.935 108.845 ;
        RECT 22.955 108.035 24.305 108.945 ;
        RECT 24.335 108.120 24.765 108.905 ;
        RECT 25.255 108.035 26.605 108.945 ;
        RECT 26.625 108.035 27.995 108.815 ;
        RECT 28.005 108.035 29.835 108.845 ;
        RECT 29.855 108.035 31.205 108.945 ;
        RECT 31.225 108.035 32.595 108.815 ;
        RECT 32.605 108.035 33.975 108.815 ;
        RECT 33.985 108.035 35.355 108.815 ;
        RECT 35.365 108.715 36.285 108.945 ;
        RECT 39.115 108.715 40.045 108.935 ;
        RECT 35.365 108.035 44.555 108.715 ;
        RECT 45.025 108.035 46.395 108.815 ;
        RECT 47.465 108.035 50.075 108.945 ;
        RECT 50.095 108.120 50.525 108.905 ;
        RECT 50.545 108.035 56.055 108.845 ;
        RECT 56.075 108.035 57.425 108.945 ;
        RECT 57.445 108.035 59.275 108.845 ;
        RECT 59.285 108.035 60.655 108.815 ;
        RECT 60.665 108.035 62.035 108.845 ;
        RECT 62.045 108.035 67.555 108.845 ;
        RECT 67.565 108.035 68.935 108.815 ;
        RECT 68.945 108.035 74.455 108.845 ;
        RECT 74.475 108.035 75.825 108.945 ;
        RECT 75.855 108.120 76.285 108.905 ;
        RECT 76.305 108.035 78.135 108.845 ;
        RECT 78.155 108.035 79.505 108.945 ;
        RECT 79.525 108.035 80.895 108.815 ;
        RECT 80.905 108.035 83.515 108.945 ;
        RECT 84.125 108.035 86.875 108.845 ;
        RECT 86.895 108.035 88.245 108.945 ;
        RECT 88.265 108.035 89.635 108.845 ;
        RECT 89.655 108.035 91.005 108.945 ;
        RECT 91.025 108.035 92.395 108.815 ;
        RECT 92.405 108.715 93.325 108.945 ;
        RECT 96.155 108.715 97.085 108.935 ;
        RECT 92.405 108.035 101.595 108.715 ;
        RECT 101.615 108.120 102.045 108.905 ;
        RECT 102.535 108.035 103.885 108.945 ;
        RECT 104.365 108.035 105.735 108.815 ;
        RECT 105.745 108.035 107.115 108.845 ;
        RECT 107.135 108.035 108.485 108.945 ;
        RECT 108.505 108.035 110.335 108.845 ;
        RECT 110.345 108.035 115.855 108.845 ;
        RECT 115.875 108.035 117.225 108.945 ;
        RECT 117.245 108.715 118.165 108.945 ;
        RECT 120.995 108.715 121.925 108.935 ;
        RECT 117.245 108.035 126.435 108.715 ;
        RECT 126.445 108.035 127.815 108.845 ;
        RECT 14.805 107.825 14.975 108.035 ;
        RECT 17.105 107.825 17.275 108.035 ;
        RECT 18.485 107.825 18.655 108.015 ;
        RECT 22.625 107.845 22.795 108.035 ;
        RECT 23.085 107.845 23.255 108.035 ;
        RECT 24.980 107.875 25.100 107.985 ;
        RECT 26.305 107.845 26.475 108.035 ;
        RECT 26.765 107.845 26.935 108.035 ;
        RECT 27.685 107.825 27.855 108.015 ;
        RECT 29.525 107.845 29.695 108.035 ;
        RECT 29.985 107.845 30.155 108.035 ;
        RECT 32.285 107.845 32.455 108.035 ;
        RECT 33.665 107.845 33.835 108.035 ;
        RECT 34.125 107.845 34.295 108.035 ;
        RECT 36.885 107.825 37.055 108.015 ;
        RECT 37.860 107.875 37.980 107.985 ;
        RECT 38.265 107.825 38.435 108.015 ;
        RECT 44.245 107.845 44.415 108.035 ;
        RECT 44.760 107.875 44.880 107.985 ;
        RECT 45.165 107.845 45.335 108.035 ;
        RECT 49.760 108.015 49.930 108.035 ;
        RECT 47.005 107.880 47.165 107.990 ;
        RECT 48.385 107.825 48.555 108.015 ;
        RECT 49.760 107.845 49.935 108.015 ;
        RECT 49.765 107.825 49.935 107.845 ;
        RECT 51.145 107.825 51.315 108.015 ;
        RECT 51.605 107.825 51.775 108.015 ;
        RECT 53.445 107.870 53.605 107.980 ;
        RECT 54.825 107.825 54.995 108.015 ;
        RECT 55.340 107.875 55.460 107.985 ;
        RECT 55.745 107.825 55.915 108.035 ;
        RECT 56.205 107.845 56.375 108.035 ;
        RECT 57.585 107.870 57.745 107.980 ;
        RECT 58.965 107.845 59.135 108.035 ;
        RECT 59.425 107.845 59.595 108.035 ;
        RECT 61.265 107.825 61.435 108.015 ;
        RECT 61.725 107.825 61.895 108.035 ;
        RECT 67.245 107.845 67.415 108.035 ;
        RECT 67.705 107.845 67.875 108.035 ;
        RECT 72.305 107.825 72.475 108.015 ;
        RECT 73.225 107.870 73.385 107.980 ;
        RECT 74.145 107.845 74.315 108.035 ;
        RECT 75.525 107.845 75.695 108.035 ;
        RECT 77.825 107.845 77.995 108.035 ;
        RECT 79.205 107.845 79.375 108.035 ;
        RECT 79.665 107.845 79.835 108.035 ;
        RECT 81.050 107.845 81.220 108.035 ;
        RECT 82.425 107.825 82.595 108.015 ;
        RECT 82.885 107.825 83.055 108.015 ;
        RECT 83.860 107.875 83.980 107.985 ;
        RECT 85.185 107.825 85.355 108.015 ;
        RECT 86.105 107.870 86.265 107.980 ;
        RECT 86.565 107.825 86.735 108.035 ;
        RECT 87.025 107.845 87.195 108.035 ;
        RECT 88.405 107.870 88.565 107.980 ;
        RECT 89.325 107.845 89.495 108.035 ;
        RECT 89.785 107.845 89.955 108.035 ;
        RECT 91.165 107.845 91.335 108.035 ;
        RECT 98.065 107.825 98.235 108.015 ;
        RECT 99.445 107.825 99.615 108.015 ;
        RECT 101.285 107.845 101.455 108.035 ;
        RECT 102.260 107.875 102.380 107.985 ;
        RECT 103.585 107.845 103.755 108.035 ;
        RECT 104.100 107.875 104.220 107.985 ;
        RECT 104.505 107.845 104.675 108.035 ;
        RECT 106.805 107.845 106.975 108.035 ;
        RECT 108.185 107.845 108.355 108.035 ;
        RECT 108.645 107.825 108.815 108.015 ;
        RECT 109.105 107.825 109.275 108.015 ;
        RECT 110.025 107.845 110.195 108.035 ;
        RECT 111.405 107.825 111.575 108.015 ;
        RECT 111.865 107.825 112.035 108.015 ;
        RECT 113.245 107.825 113.415 108.015 ;
        RECT 115.085 107.825 115.255 108.015 ;
        RECT 115.545 107.845 115.715 108.035 ;
        RECT 116.005 107.845 116.175 108.035 ;
        RECT 116.925 107.870 117.085 107.980 ;
        RECT 117.385 107.825 117.555 108.015 ;
        RECT 126.125 107.845 126.295 108.035 ;
        RECT 127.505 107.825 127.675 108.035 ;
        RECT 14.665 107.015 16.035 107.825 ;
        RECT 16.045 107.015 17.415 107.825 ;
        RECT 17.435 106.915 18.785 107.825 ;
        RECT 18.805 107.145 27.995 107.825 ;
        RECT 28.005 107.145 37.195 107.825 ;
        RECT 18.805 106.915 19.725 107.145 ;
        RECT 22.555 106.925 23.485 107.145 ;
        RECT 28.005 106.915 28.925 107.145 ;
        RECT 31.755 106.925 32.685 107.145 ;
        RECT 37.215 106.955 37.645 107.740 ;
        RECT 38.135 106.915 39.485 107.825 ;
        RECT 39.505 107.145 48.695 107.825 ;
        RECT 39.505 106.915 40.425 107.145 ;
        RECT 43.255 106.925 44.185 107.145 ;
        RECT 48.705 107.045 50.075 107.825 ;
        RECT 50.085 107.015 51.455 107.825 ;
        RECT 51.465 107.045 52.835 107.825 ;
        RECT 53.765 107.045 55.135 107.825 ;
        RECT 55.615 106.915 56.965 107.825 ;
        RECT 57.905 107.015 61.575 107.825 ;
        RECT 61.595 106.915 62.945 107.825 ;
        RECT 62.975 106.955 63.405 107.740 ;
        RECT 63.425 107.145 72.615 107.825 ;
        RECT 73.545 107.145 82.735 107.825 ;
        RECT 63.425 106.915 64.345 107.145 ;
        RECT 67.175 106.925 68.105 107.145 ;
        RECT 73.545 106.915 74.465 107.145 ;
        RECT 77.295 106.925 78.225 107.145 ;
        RECT 82.745 107.045 84.115 107.825 ;
        RECT 84.135 106.915 85.485 107.825 ;
        RECT 86.425 107.045 87.795 107.825 ;
        RECT 88.735 106.955 89.165 107.740 ;
        RECT 89.185 107.145 98.375 107.825 ;
        RECT 89.185 106.915 90.105 107.145 ;
        RECT 92.935 106.925 93.865 107.145 ;
        RECT 98.395 106.915 99.745 107.825 ;
        RECT 99.765 107.145 108.955 107.825 ;
        RECT 99.765 106.915 100.685 107.145 ;
        RECT 103.515 106.925 104.445 107.145 ;
        RECT 108.965 107.045 110.335 107.825 ;
        RECT 110.345 107.015 111.715 107.825 ;
        RECT 111.735 106.915 113.085 107.825 ;
        RECT 113.105 107.045 114.475 107.825 ;
        RECT 114.495 106.955 114.925 107.740 ;
        RECT 114.955 106.915 116.305 107.825 ;
        RECT 117.245 107.145 126.435 107.825 ;
        RECT 121.755 106.925 122.685 107.145 ;
        RECT 125.515 106.915 126.435 107.145 ;
        RECT 126.445 107.015 127.815 107.825 ;
      LAYER nwell ;
        RECT 14.470 103.795 128.010 106.625 ;
      LAYER pwell ;
        RECT 14.665 102.595 16.035 103.405 ;
        RECT 16.045 102.595 18.795 103.405 ;
        RECT 18.805 102.595 24.315 103.405 ;
        RECT 24.335 102.680 24.765 103.465 ;
        RECT 24.785 103.275 25.705 103.505 ;
        RECT 28.535 103.275 29.465 103.495 ;
        RECT 24.785 102.595 33.975 103.275 ;
        RECT 34.445 102.595 38.115 103.405 ;
        RECT 38.135 102.595 39.485 103.505 ;
        RECT 39.505 102.595 40.875 103.405 ;
        RECT 45.395 103.275 46.325 103.495 ;
        RECT 49.155 103.275 50.075 103.505 ;
        RECT 40.885 102.595 50.075 103.275 ;
        RECT 50.095 102.680 50.525 103.465 ;
        RECT 55.515 103.275 56.445 103.495 ;
        RECT 59.275 103.275 60.195 103.505 ;
        RECT 51.005 102.595 60.195 103.275 ;
        RECT 60.205 103.275 61.125 103.505 ;
        RECT 63.955 103.275 64.885 103.495 ;
        RECT 60.205 102.595 69.395 103.275 ;
        RECT 70.325 102.595 75.835 103.405 ;
        RECT 75.855 102.680 76.285 103.465 ;
        RECT 76.305 103.275 77.225 103.505 ;
        RECT 80.055 103.275 80.985 103.495 ;
        RECT 85.505 103.275 86.425 103.505 ;
        RECT 89.255 103.275 90.185 103.495 ;
        RECT 76.305 102.595 85.495 103.275 ;
        RECT 85.505 102.595 94.695 103.275 ;
        RECT 94.705 102.595 96.075 103.405 ;
        RECT 96.085 102.595 101.595 103.405 ;
        RECT 101.615 102.680 102.045 103.465 ;
        RECT 102.525 102.595 104.355 103.405 ;
        RECT 104.365 103.275 105.285 103.505 ;
        RECT 108.115 103.275 109.045 103.495 ;
        RECT 113.565 103.275 114.485 103.505 ;
        RECT 117.315 103.275 118.245 103.495 ;
        RECT 104.365 102.595 113.555 103.275 ;
        RECT 113.565 102.595 122.755 103.275 ;
        RECT 123.225 102.595 125.055 103.405 ;
        RECT 125.065 102.595 126.435 103.375 ;
        RECT 126.445 102.595 127.815 103.405 ;
        RECT 14.805 102.385 14.975 102.595 ;
        RECT 18.485 102.385 18.655 102.595 ;
        RECT 24.005 102.385 24.175 102.595 ;
        RECT 25.845 102.385 26.015 102.575 ;
        RECT 31.365 102.385 31.535 102.575 ;
        RECT 33.665 102.405 33.835 102.595 ;
        RECT 34.180 102.435 34.300 102.545 ;
        RECT 36.885 102.385 37.055 102.575 ;
        RECT 37.805 102.405 37.975 102.595 ;
        RECT 39.185 102.405 39.355 102.595 ;
        RECT 40.565 102.405 40.735 102.595 ;
        RECT 41.025 102.385 41.195 102.595 ;
        RECT 46.545 102.385 46.715 102.575 ;
        RECT 47.925 102.385 48.095 102.575 ;
        RECT 49.765 102.385 49.935 102.575 ;
        RECT 50.740 102.435 50.860 102.545 ;
        RECT 51.145 102.405 51.315 102.595 ;
        RECT 51.605 102.385 51.775 102.575 ;
        RECT 57.125 102.385 57.295 102.575 ;
        RECT 62.645 102.385 62.815 102.575 ;
        RECT 64.025 102.430 64.185 102.540 ;
        RECT 64.485 102.385 64.655 102.575 ;
        RECT 66.325 102.430 66.485 102.540 ;
        RECT 69.085 102.405 69.255 102.595 ;
        RECT 70.005 102.385 70.175 102.575 ;
        RECT 75.525 102.385 75.695 102.595 ;
        RECT 77.365 102.385 77.535 102.575 ;
        RECT 82.885 102.385 83.055 102.575 ;
        RECT 85.185 102.405 85.355 102.595 ;
        RECT 88.405 102.385 88.575 102.575 ;
        RECT 90.245 102.385 90.415 102.575 ;
        RECT 94.385 102.405 94.555 102.595 ;
        RECT 95.765 102.385 95.935 102.595 ;
        RECT 101.285 102.385 101.455 102.595 ;
        RECT 102.260 102.435 102.380 102.545 ;
        RECT 103.125 102.385 103.295 102.575 ;
        RECT 104.045 102.405 104.215 102.595 ;
        RECT 108.645 102.385 108.815 102.575 ;
        RECT 113.245 102.405 113.415 102.595 ;
        RECT 114.165 102.385 114.335 102.575 ;
        RECT 115.140 102.435 115.260 102.545 ;
        RECT 120.605 102.385 120.775 102.575 ;
        RECT 122.445 102.405 122.615 102.595 ;
        RECT 122.960 102.435 123.080 102.545 ;
        RECT 124.745 102.405 124.915 102.595 ;
        RECT 126.115 102.575 126.285 102.595 ;
        RECT 126.115 102.405 126.295 102.575 ;
        RECT 126.125 102.385 126.295 102.405 ;
        RECT 127.505 102.385 127.675 102.595 ;
        RECT 14.665 101.575 16.035 102.385 ;
        RECT 16.045 101.575 18.795 102.385 ;
        RECT 18.805 101.575 24.315 102.385 ;
        RECT 24.335 101.515 24.765 102.300 ;
        RECT 24.785 101.575 26.155 102.385 ;
        RECT 26.165 101.575 31.675 102.385 ;
        RECT 31.685 101.575 37.195 102.385 ;
        RECT 37.215 101.515 37.645 102.300 ;
        RECT 37.665 101.575 41.335 102.385 ;
        RECT 41.345 101.575 46.855 102.385 ;
        RECT 46.875 101.475 48.225 102.385 ;
        RECT 48.245 101.575 50.075 102.385 ;
        RECT 50.095 101.515 50.525 102.300 ;
        RECT 50.545 101.575 51.915 102.385 ;
        RECT 51.925 101.575 57.435 102.385 ;
        RECT 57.445 101.575 62.955 102.385 ;
        RECT 62.975 101.515 63.405 102.300 ;
        RECT 64.355 101.475 65.705 102.385 ;
        RECT 66.645 101.575 70.315 102.385 ;
        RECT 70.325 101.575 75.835 102.385 ;
        RECT 75.855 101.515 76.285 102.300 ;
        RECT 76.305 101.575 77.675 102.385 ;
        RECT 77.685 101.575 83.195 102.385 ;
        RECT 83.205 101.575 88.715 102.385 ;
        RECT 88.735 101.515 89.165 102.300 ;
        RECT 89.185 101.575 90.555 102.385 ;
        RECT 90.565 101.575 96.075 102.385 ;
        RECT 96.085 101.575 101.595 102.385 ;
        RECT 101.615 101.515 102.045 102.300 ;
        RECT 102.065 101.575 103.435 102.385 ;
        RECT 103.445 101.575 108.955 102.385 ;
        RECT 108.965 101.575 114.475 102.385 ;
        RECT 114.495 101.515 114.925 102.300 ;
        RECT 115.405 101.575 120.915 102.385 ;
        RECT 120.925 101.575 126.435 102.385 ;
        RECT 126.445 101.575 127.815 102.385 ;
      LAYER nwell ;
        RECT 14.470 99.580 128.010 101.185 ;
        RECT 20.485 54.580 29.875 66.420 ;
        RECT 31.685 54.590 41.075 66.430 ;
        RECT 42.905 54.560 52.295 66.400 ;
        RECT 54.155 54.540 63.545 66.380 ;
        RECT 65.375 54.530 74.765 66.370 ;
        RECT 76.615 54.520 86.005 66.360 ;
        RECT 87.865 54.530 97.255 66.370 ;
        RECT 99.145 54.520 108.535 66.360 ;
        RECT 110.415 54.520 119.805 66.360 ;
        RECT 121.665 54.520 131.055 66.360 ;
        RECT 132.415 54.490 139.375 66.330 ;
        RECT 20.655 49.020 23.115 53.210 ;
      LAYER pwell ;
        RECT 20.555 45.340 22.915 48.340 ;
      LAYER nwell ;
        RECT 24.735 45.940 29.125 53.130 ;
        RECT 31.855 49.030 34.315 53.220 ;
      LAYER pwell ;
        RECT 31.755 45.350 34.115 48.350 ;
      LAYER nwell ;
        RECT 35.935 45.950 40.325 53.140 ;
        RECT 43.075 49.000 45.535 53.190 ;
      LAYER pwell ;
        RECT 42.975 45.320 45.335 48.320 ;
      LAYER nwell ;
        RECT 47.155 45.920 51.545 53.110 ;
        RECT 54.325 48.980 56.785 53.170 ;
      LAYER pwell ;
        RECT 54.225 45.300 56.585 48.300 ;
      LAYER nwell ;
        RECT 58.405 45.900 62.795 53.090 ;
        RECT 65.545 48.970 68.005 53.160 ;
      LAYER pwell ;
        RECT 65.445 45.290 67.805 48.290 ;
      LAYER nwell ;
        RECT 69.625 45.890 74.015 53.080 ;
        RECT 76.785 48.960 79.245 53.150 ;
      LAYER pwell ;
        RECT 76.685 45.280 79.045 48.280 ;
      LAYER nwell ;
        RECT 80.865 45.880 85.255 53.070 ;
        RECT 88.035 48.970 90.495 53.160 ;
      LAYER pwell ;
        RECT 87.935 45.290 90.295 48.290 ;
      LAYER nwell ;
        RECT 92.115 45.890 96.505 53.080 ;
        RECT 99.315 48.960 101.775 53.150 ;
      LAYER pwell ;
        RECT 99.215 45.280 101.575 48.280 ;
      LAYER nwell ;
        RECT 103.395 45.880 107.785 53.070 ;
        RECT 110.585 48.960 113.045 53.150 ;
      LAYER pwell ;
        RECT 110.485 45.280 112.845 48.280 ;
      LAYER nwell ;
        RECT 114.665 45.880 119.055 53.070 ;
        RECT 121.835 48.960 124.295 53.150 ;
      LAYER pwell ;
        RECT 121.735 45.280 124.095 48.280 ;
      LAYER nwell ;
        RECT 125.915 45.880 130.305 53.070 ;
        RECT 19.615 32.280 24.005 39.470 ;
      LAYER pwell ;
        RECT 25.825 37.070 28.185 40.070 ;
      LAYER nwell ;
        RECT 25.625 32.200 28.085 36.390 ;
        RECT 30.895 32.280 35.285 39.470 ;
      LAYER pwell ;
        RECT 37.105 37.070 39.465 40.070 ;
      LAYER nwell ;
        RECT 36.905 32.200 39.365 36.390 ;
        RECT 42.185 32.260 46.575 39.450 ;
      LAYER pwell ;
        RECT 48.395 37.050 50.755 40.050 ;
      LAYER nwell ;
        RECT 48.195 32.180 50.655 36.370 ;
        RECT 53.405 32.260 57.795 39.450 ;
      LAYER pwell ;
        RECT 59.615 37.050 61.975 40.050 ;
      LAYER nwell ;
        RECT 59.415 32.180 61.875 36.370 ;
        RECT 64.605 32.260 68.995 39.450 ;
      LAYER pwell ;
        RECT 70.815 37.050 73.175 40.050 ;
      LAYER nwell ;
        RECT 70.615 32.180 73.075 36.370 ;
        RECT 75.895 32.250 80.285 39.440 ;
      LAYER pwell ;
        RECT 82.105 37.040 84.465 40.040 ;
      LAYER nwell ;
        RECT 81.905 32.170 84.365 36.360 ;
        RECT 87.135 32.270 91.525 39.460 ;
      LAYER pwell ;
        RECT 93.345 37.060 95.705 40.060 ;
      LAYER nwell ;
        RECT 93.145 32.190 95.605 36.380 ;
        RECT 98.345 32.290 102.735 39.480 ;
      LAYER pwell ;
        RECT 104.555 37.080 106.915 40.080 ;
      LAYER nwell ;
        RECT 104.355 32.210 106.815 36.400 ;
        RECT 109.545 32.330 113.935 39.520 ;
      LAYER pwell ;
        RECT 115.755 37.120 118.115 40.120 ;
      LAYER nwell ;
        RECT 115.555 32.250 118.015 36.440 ;
        RECT 120.755 32.350 125.145 39.540 ;
      LAYER pwell ;
        RECT 126.965 37.140 129.325 40.140 ;
      LAYER nwell ;
        RECT 126.765 32.270 129.225 36.460 ;
        RECT 18.865 18.990 28.255 30.830 ;
        RECT 30.145 18.990 39.535 30.830 ;
        RECT 41.435 18.970 50.825 30.810 ;
        RECT 52.655 18.970 62.045 30.810 ;
        RECT 63.855 18.970 73.245 30.810 ;
        RECT 75.145 18.960 84.535 30.800 ;
        RECT 86.385 18.980 95.775 30.820 ;
        RECT 97.595 19.000 106.985 30.840 ;
        RECT 108.795 19.040 118.185 30.880 ;
        RECT 120.005 19.060 129.395 30.900 ;
        RECT 131.725 19.030 138.685 30.870 ;
      LAYER li1 ;
        RECT 14.660 211.205 127.820 211.375 ;
        RECT 14.745 210.455 15.955 211.205 ;
        RECT 14.745 209.915 15.265 210.455 ;
        RECT 16.125 210.435 18.715 211.205 ;
        RECT 18.890 210.660 24.235 211.205 ;
        RECT 15.435 209.745 15.955 210.285 ;
        RECT 14.745 208.655 15.955 209.745 ;
        RECT 16.125 209.745 17.335 210.265 ;
        RECT 17.505 209.915 18.715 210.435 ;
        RECT 16.125 208.655 18.715 209.745 ;
        RECT 20.480 209.090 20.830 210.340 ;
        RECT 22.310 209.830 22.650 210.660 ;
        RECT 24.405 210.480 24.695 211.205 ;
        RECT 24.865 210.455 26.075 211.205 ;
        RECT 26.250 210.660 31.595 211.205 ;
        RECT 31.770 210.660 37.115 211.205 ;
        RECT 18.890 208.655 24.235 209.090 ;
        RECT 24.405 208.655 24.695 209.820 ;
        RECT 24.865 209.745 25.385 210.285 ;
        RECT 25.555 209.915 26.075 210.455 ;
        RECT 24.865 208.655 26.075 209.745 ;
        RECT 27.840 209.090 28.190 210.340 ;
        RECT 29.670 209.830 30.010 210.660 ;
        RECT 33.360 209.090 33.710 210.340 ;
        RECT 35.190 209.830 35.530 210.660 ;
        RECT 37.285 210.480 37.575 211.205 ;
        RECT 37.745 210.455 38.955 211.205 ;
        RECT 39.130 210.660 44.475 211.205 ;
        RECT 44.650 210.660 49.995 211.205 ;
        RECT 26.250 208.655 31.595 209.090 ;
        RECT 31.770 208.655 37.115 209.090 ;
        RECT 37.285 208.655 37.575 209.820 ;
        RECT 37.745 209.745 38.265 210.285 ;
        RECT 38.435 209.915 38.955 210.455 ;
        RECT 37.745 208.655 38.955 209.745 ;
        RECT 40.720 209.090 41.070 210.340 ;
        RECT 42.550 209.830 42.890 210.660 ;
        RECT 46.240 209.090 46.590 210.340 ;
        RECT 48.070 209.830 48.410 210.660 ;
        RECT 50.165 210.480 50.455 211.205 ;
        RECT 50.625 210.455 51.835 211.205 ;
        RECT 52.010 210.660 57.355 211.205 ;
        RECT 57.530 210.660 62.875 211.205 ;
        RECT 39.130 208.655 44.475 209.090 ;
        RECT 44.650 208.655 49.995 209.090 ;
        RECT 50.165 208.655 50.455 209.820 ;
        RECT 50.625 209.745 51.145 210.285 ;
        RECT 51.315 209.915 51.835 210.455 ;
        RECT 50.625 208.655 51.835 209.745 ;
        RECT 53.600 209.090 53.950 210.340 ;
        RECT 55.430 209.830 55.770 210.660 ;
        RECT 59.120 209.090 59.470 210.340 ;
        RECT 60.950 209.830 61.290 210.660 ;
        RECT 63.045 210.480 63.335 211.205 ;
        RECT 63.505 210.455 64.715 211.205 ;
        RECT 64.890 210.660 70.235 211.205 ;
        RECT 70.410 210.660 75.755 211.205 ;
        RECT 52.010 208.655 57.355 209.090 ;
        RECT 57.530 208.655 62.875 209.090 ;
        RECT 63.045 208.655 63.335 209.820 ;
        RECT 63.505 209.745 64.025 210.285 ;
        RECT 64.195 209.915 64.715 210.455 ;
        RECT 63.505 208.655 64.715 209.745 ;
        RECT 66.480 209.090 66.830 210.340 ;
        RECT 68.310 209.830 68.650 210.660 ;
        RECT 72.000 209.090 72.350 210.340 ;
        RECT 73.830 209.830 74.170 210.660 ;
        RECT 75.925 210.480 76.215 211.205 ;
        RECT 76.385 210.455 77.595 211.205 ;
        RECT 77.770 210.660 83.115 211.205 ;
        RECT 83.290 210.660 88.635 211.205 ;
        RECT 64.890 208.655 70.235 209.090 ;
        RECT 70.410 208.655 75.755 209.090 ;
        RECT 75.925 208.655 76.215 209.820 ;
        RECT 76.385 209.745 76.905 210.285 ;
        RECT 77.075 209.915 77.595 210.455 ;
        RECT 76.385 208.655 77.595 209.745 ;
        RECT 79.360 209.090 79.710 210.340 ;
        RECT 81.190 209.830 81.530 210.660 ;
        RECT 84.880 209.090 85.230 210.340 ;
        RECT 86.710 209.830 87.050 210.660 ;
        RECT 88.805 210.480 89.095 211.205 ;
        RECT 89.265 210.455 90.475 211.205 ;
        RECT 90.650 210.660 95.995 211.205 ;
        RECT 96.170 210.660 101.515 211.205 ;
        RECT 77.770 208.655 83.115 209.090 ;
        RECT 83.290 208.655 88.635 209.090 ;
        RECT 88.805 208.655 89.095 209.820 ;
        RECT 89.265 209.745 89.785 210.285 ;
        RECT 89.955 209.915 90.475 210.455 ;
        RECT 89.265 208.655 90.475 209.745 ;
        RECT 92.240 209.090 92.590 210.340 ;
        RECT 94.070 209.830 94.410 210.660 ;
        RECT 97.760 209.090 98.110 210.340 ;
        RECT 99.590 209.830 99.930 210.660 ;
        RECT 101.685 210.480 101.975 211.205 ;
        RECT 102.145 210.455 103.355 211.205 ;
        RECT 103.530 210.660 108.875 211.205 ;
        RECT 109.050 210.660 114.395 211.205 ;
        RECT 90.650 208.655 95.995 209.090 ;
        RECT 96.170 208.655 101.515 209.090 ;
        RECT 101.685 208.655 101.975 209.820 ;
        RECT 102.145 209.745 102.665 210.285 ;
        RECT 102.835 209.915 103.355 210.455 ;
        RECT 102.145 208.655 103.355 209.745 ;
        RECT 105.120 209.090 105.470 210.340 ;
        RECT 106.950 209.830 107.290 210.660 ;
        RECT 110.640 209.090 110.990 210.340 ;
        RECT 112.470 209.830 112.810 210.660 ;
        RECT 114.565 210.480 114.855 211.205 ;
        RECT 115.490 210.660 120.835 211.205 ;
        RECT 121.010 210.660 126.355 211.205 ;
        RECT 103.530 208.655 108.875 209.090 ;
        RECT 109.050 208.655 114.395 209.090 ;
        RECT 114.565 208.655 114.855 209.820 ;
        RECT 117.080 209.090 117.430 210.340 ;
        RECT 118.910 209.830 119.250 210.660 ;
        RECT 122.600 209.090 122.950 210.340 ;
        RECT 124.430 209.830 124.770 210.660 ;
        RECT 126.525 210.455 127.735 211.205 ;
        RECT 126.525 209.745 127.045 210.285 ;
        RECT 127.215 209.915 127.735 210.455 ;
        RECT 115.490 208.655 120.835 209.090 ;
        RECT 121.010 208.655 126.355 209.090 ;
        RECT 126.525 208.655 127.735 209.745 ;
        RECT 14.660 208.485 127.820 208.655 ;
        RECT 14.745 207.395 15.955 208.485 ;
        RECT 14.745 206.685 15.265 207.225 ;
        RECT 15.435 206.855 15.955 207.395 ;
        RECT 16.125 207.395 18.715 208.485 ;
        RECT 18.890 208.050 24.235 208.485 ;
        RECT 16.125 206.875 17.335 207.395 ;
        RECT 17.505 206.705 18.715 207.225 ;
        RECT 20.480 206.800 20.830 208.050 ;
        RECT 24.405 207.320 24.695 208.485 ;
        RECT 25.325 207.395 27.915 208.485 ;
        RECT 28.090 208.050 33.435 208.485 ;
        RECT 33.610 208.050 38.955 208.485 ;
        RECT 39.130 208.050 44.475 208.485 ;
        RECT 44.650 208.050 49.995 208.485 ;
        RECT 14.745 205.935 15.955 206.685 ;
        RECT 16.125 205.935 18.715 206.705 ;
        RECT 22.310 206.480 22.650 207.310 ;
        RECT 25.325 206.875 26.535 207.395 ;
        RECT 26.705 206.705 27.915 207.225 ;
        RECT 29.680 206.800 30.030 208.050 ;
        RECT 18.890 205.935 24.235 206.480 ;
        RECT 24.405 205.935 24.695 206.660 ;
        RECT 25.325 205.935 27.915 206.705 ;
        RECT 31.510 206.480 31.850 207.310 ;
        RECT 35.200 206.800 35.550 208.050 ;
        RECT 37.030 206.480 37.370 207.310 ;
        RECT 40.720 206.800 41.070 208.050 ;
        RECT 42.550 206.480 42.890 207.310 ;
        RECT 46.240 206.800 46.590 208.050 ;
        RECT 50.165 207.320 50.455 208.485 ;
        RECT 51.085 207.395 53.675 208.485 ;
        RECT 53.850 208.050 59.195 208.485 ;
        RECT 59.370 208.050 64.715 208.485 ;
        RECT 64.890 208.050 70.235 208.485 ;
        RECT 70.410 208.050 75.755 208.485 ;
        RECT 48.070 206.480 48.410 207.310 ;
        RECT 51.085 206.875 52.295 207.395 ;
        RECT 52.465 206.705 53.675 207.225 ;
        RECT 55.440 206.800 55.790 208.050 ;
        RECT 28.090 205.935 33.435 206.480 ;
        RECT 33.610 205.935 38.955 206.480 ;
        RECT 39.130 205.935 44.475 206.480 ;
        RECT 44.650 205.935 49.995 206.480 ;
        RECT 50.165 205.935 50.455 206.660 ;
        RECT 51.085 205.935 53.675 206.705 ;
        RECT 57.270 206.480 57.610 207.310 ;
        RECT 60.960 206.800 61.310 208.050 ;
        RECT 62.790 206.480 63.130 207.310 ;
        RECT 66.480 206.800 66.830 208.050 ;
        RECT 68.310 206.480 68.650 207.310 ;
        RECT 72.000 206.800 72.350 208.050 ;
        RECT 75.925 207.320 76.215 208.485 ;
        RECT 76.845 207.395 79.435 208.485 ;
        RECT 79.610 208.050 84.955 208.485 ;
        RECT 85.130 208.050 90.475 208.485 ;
        RECT 90.650 208.050 95.995 208.485 ;
        RECT 96.170 208.050 101.515 208.485 ;
        RECT 73.830 206.480 74.170 207.310 ;
        RECT 76.845 206.875 78.055 207.395 ;
        RECT 78.225 206.705 79.435 207.225 ;
        RECT 81.200 206.800 81.550 208.050 ;
        RECT 53.850 205.935 59.195 206.480 ;
        RECT 59.370 205.935 64.715 206.480 ;
        RECT 64.890 205.935 70.235 206.480 ;
        RECT 70.410 205.935 75.755 206.480 ;
        RECT 75.925 205.935 76.215 206.660 ;
        RECT 76.845 205.935 79.435 206.705 ;
        RECT 83.030 206.480 83.370 207.310 ;
        RECT 86.720 206.800 87.070 208.050 ;
        RECT 88.550 206.480 88.890 207.310 ;
        RECT 92.240 206.800 92.590 208.050 ;
        RECT 94.070 206.480 94.410 207.310 ;
        RECT 97.760 206.800 98.110 208.050 ;
        RECT 101.685 207.320 101.975 208.485 ;
        RECT 102.605 207.395 104.275 208.485 ;
        RECT 104.450 208.050 109.795 208.485 ;
        RECT 109.970 208.050 115.315 208.485 ;
        RECT 115.490 208.050 120.835 208.485 ;
        RECT 121.010 208.050 126.355 208.485 ;
        RECT 99.590 206.480 99.930 207.310 ;
        RECT 102.605 206.875 103.355 207.395 ;
        RECT 103.525 206.705 104.275 207.225 ;
        RECT 106.040 206.800 106.390 208.050 ;
        RECT 79.610 205.935 84.955 206.480 ;
        RECT 85.130 205.935 90.475 206.480 ;
        RECT 90.650 205.935 95.995 206.480 ;
        RECT 96.170 205.935 101.515 206.480 ;
        RECT 101.685 205.935 101.975 206.660 ;
        RECT 102.605 205.935 104.275 206.705 ;
        RECT 107.870 206.480 108.210 207.310 ;
        RECT 111.560 206.800 111.910 208.050 ;
        RECT 113.390 206.480 113.730 207.310 ;
        RECT 117.080 206.800 117.430 208.050 ;
        RECT 118.910 206.480 119.250 207.310 ;
        RECT 122.600 206.800 122.950 208.050 ;
        RECT 126.525 207.395 127.735 208.485 ;
        RECT 124.430 206.480 124.770 207.310 ;
        RECT 126.525 206.855 127.045 207.395 ;
        RECT 127.215 206.685 127.735 207.225 ;
        RECT 104.450 205.935 109.795 206.480 ;
        RECT 109.970 205.935 115.315 206.480 ;
        RECT 115.490 205.935 120.835 206.480 ;
        RECT 121.010 205.935 126.355 206.480 ;
        RECT 126.525 205.935 127.735 206.685 ;
        RECT 14.660 205.765 127.820 205.935 ;
        RECT 14.745 205.015 15.955 205.765 ;
        RECT 14.745 204.475 15.265 205.015 ;
        RECT 17.045 204.995 20.555 205.765 ;
        RECT 20.730 205.220 26.075 205.765 ;
        RECT 26.250 205.220 31.595 205.765 ;
        RECT 31.770 205.220 37.115 205.765 ;
        RECT 15.435 204.305 15.955 204.845 ;
        RECT 14.745 203.215 15.955 204.305 ;
        RECT 17.045 204.305 18.735 204.825 ;
        RECT 18.905 204.475 20.555 204.995 ;
        RECT 17.045 203.215 20.555 204.305 ;
        RECT 22.320 203.650 22.670 204.900 ;
        RECT 24.150 204.390 24.490 205.220 ;
        RECT 27.840 203.650 28.190 204.900 ;
        RECT 29.670 204.390 30.010 205.220 ;
        RECT 33.360 203.650 33.710 204.900 ;
        RECT 35.190 204.390 35.530 205.220 ;
        RECT 37.285 205.040 37.575 205.765 ;
        RECT 38.205 204.995 40.795 205.765 ;
        RECT 40.970 205.220 46.315 205.765 ;
        RECT 46.490 205.220 51.835 205.765 ;
        RECT 52.010 205.220 57.355 205.765 ;
        RECT 57.530 205.220 62.875 205.765 ;
        RECT 20.730 203.215 26.075 203.650 ;
        RECT 26.250 203.215 31.595 203.650 ;
        RECT 31.770 203.215 37.115 203.650 ;
        RECT 37.285 203.215 37.575 204.380 ;
        RECT 38.205 204.305 39.415 204.825 ;
        RECT 39.585 204.475 40.795 204.995 ;
        RECT 38.205 203.215 40.795 204.305 ;
        RECT 42.560 203.650 42.910 204.900 ;
        RECT 44.390 204.390 44.730 205.220 ;
        RECT 48.080 203.650 48.430 204.900 ;
        RECT 49.910 204.390 50.250 205.220 ;
        RECT 53.600 203.650 53.950 204.900 ;
        RECT 55.430 204.390 55.770 205.220 ;
        RECT 59.120 203.650 59.470 204.900 ;
        RECT 60.950 204.390 61.290 205.220 ;
        RECT 63.045 205.040 63.335 205.765 ;
        RECT 63.965 204.995 66.555 205.765 ;
        RECT 66.730 205.220 72.075 205.765 ;
        RECT 72.250 205.220 77.595 205.765 ;
        RECT 77.770 205.220 83.115 205.765 ;
        RECT 83.290 205.220 88.635 205.765 ;
        RECT 40.970 203.215 46.315 203.650 ;
        RECT 46.490 203.215 51.835 203.650 ;
        RECT 52.010 203.215 57.355 203.650 ;
        RECT 57.530 203.215 62.875 203.650 ;
        RECT 63.045 203.215 63.335 204.380 ;
        RECT 63.965 204.305 65.175 204.825 ;
        RECT 65.345 204.475 66.555 204.995 ;
        RECT 63.965 203.215 66.555 204.305 ;
        RECT 68.320 203.650 68.670 204.900 ;
        RECT 70.150 204.390 70.490 205.220 ;
        RECT 73.840 203.650 74.190 204.900 ;
        RECT 75.670 204.390 76.010 205.220 ;
        RECT 79.360 203.650 79.710 204.900 ;
        RECT 81.190 204.390 81.530 205.220 ;
        RECT 84.880 203.650 85.230 204.900 ;
        RECT 86.710 204.390 87.050 205.220 ;
        RECT 88.805 205.040 89.095 205.765 ;
        RECT 89.725 204.995 92.315 205.765 ;
        RECT 92.490 205.220 97.835 205.765 ;
        RECT 98.010 205.220 103.355 205.765 ;
        RECT 103.530 205.220 108.875 205.765 ;
        RECT 109.050 205.220 114.395 205.765 ;
        RECT 66.730 203.215 72.075 203.650 ;
        RECT 72.250 203.215 77.595 203.650 ;
        RECT 77.770 203.215 83.115 203.650 ;
        RECT 83.290 203.215 88.635 203.650 ;
        RECT 88.805 203.215 89.095 204.380 ;
        RECT 89.725 204.305 90.935 204.825 ;
        RECT 91.105 204.475 92.315 204.995 ;
        RECT 89.725 203.215 92.315 204.305 ;
        RECT 94.080 203.650 94.430 204.900 ;
        RECT 95.910 204.390 96.250 205.220 ;
        RECT 99.600 203.650 99.950 204.900 ;
        RECT 101.430 204.390 101.770 205.220 ;
        RECT 105.120 203.650 105.470 204.900 ;
        RECT 106.950 204.390 107.290 205.220 ;
        RECT 110.640 203.650 110.990 204.900 ;
        RECT 112.470 204.390 112.810 205.220 ;
        RECT 114.565 205.040 114.855 205.765 ;
        RECT 115.490 205.220 120.835 205.765 ;
        RECT 121.010 205.220 126.355 205.765 ;
        RECT 92.490 203.215 97.835 203.650 ;
        RECT 98.010 203.215 103.355 203.650 ;
        RECT 103.530 203.215 108.875 203.650 ;
        RECT 109.050 203.215 114.395 203.650 ;
        RECT 114.565 203.215 114.855 204.380 ;
        RECT 117.080 203.650 117.430 204.900 ;
        RECT 118.910 204.390 119.250 205.220 ;
        RECT 122.600 203.650 122.950 204.900 ;
        RECT 124.430 204.390 124.770 205.220 ;
        RECT 126.525 205.015 127.735 205.765 ;
        RECT 126.525 204.305 127.045 204.845 ;
        RECT 127.215 204.475 127.735 205.015 ;
        RECT 115.490 203.215 120.835 203.650 ;
        RECT 121.010 203.215 126.355 203.650 ;
        RECT 126.525 203.215 127.735 204.305 ;
        RECT 14.660 203.045 127.820 203.215 ;
        RECT 14.745 201.955 15.955 203.045 ;
        RECT 14.745 201.245 15.265 201.785 ;
        RECT 15.435 201.415 15.955 201.955 ;
        RECT 16.125 201.955 18.715 203.045 ;
        RECT 18.890 202.610 24.235 203.045 ;
        RECT 16.125 201.435 17.335 201.955 ;
        RECT 17.505 201.265 18.715 201.785 ;
        RECT 20.480 201.360 20.830 202.610 ;
        RECT 24.405 201.880 24.695 203.045 ;
        RECT 25.325 201.955 27.915 203.045 ;
        RECT 28.090 202.610 33.435 203.045 ;
        RECT 33.610 202.610 38.955 203.045 ;
        RECT 39.130 202.610 44.475 203.045 ;
        RECT 44.650 202.610 49.995 203.045 ;
        RECT 14.745 200.495 15.955 201.245 ;
        RECT 16.125 200.495 18.715 201.265 ;
        RECT 22.310 201.040 22.650 201.870 ;
        RECT 25.325 201.435 26.535 201.955 ;
        RECT 26.705 201.265 27.915 201.785 ;
        RECT 29.680 201.360 30.030 202.610 ;
        RECT 18.890 200.495 24.235 201.040 ;
        RECT 24.405 200.495 24.695 201.220 ;
        RECT 25.325 200.495 27.915 201.265 ;
        RECT 31.510 201.040 31.850 201.870 ;
        RECT 35.200 201.360 35.550 202.610 ;
        RECT 37.030 201.040 37.370 201.870 ;
        RECT 40.720 201.360 41.070 202.610 ;
        RECT 42.550 201.040 42.890 201.870 ;
        RECT 46.240 201.360 46.590 202.610 ;
        RECT 50.165 201.880 50.455 203.045 ;
        RECT 51.085 201.955 52.755 203.045 ;
        RECT 52.930 202.610 58.275 203.045 ;
        RECT 48.070 201.040 48.410 201.870 ;
        RECT 51.085 201.435 51.835 201.955 ;
        RECT 52.005 201.265 52.755 201.785 ;
        RECT 54.520 201.360 54.870 202.610 ;
        RECT 58.495 201.905 58.745 203.045 ;
        RECT 28.090 200.495 33.435 201.040 ;
        RECT 33.610 200.495 38.955 201.040 ;
        RECT 39.130 200.495 44.475 201.040 ;
        RECT 44.650 200.495 49.995 201.040 ;
        RECT 50.165 200.495 50.455 201.220 ;
        RECT 51.085 200.495 52.755 201.265 ;
        RECT 56.350 201.040 56.690 201.870 ;
        RECT 58.915 201.855 59.165 202.735 ;
        RECT 59.335 201.905 59.640 203.045 ;
        RECT 59.980 202.665 60.310 203.045 ;
        RECT 60.490 202.495 60.660 202.785 ;
        RECT 60.830 202.585 61.080 203.045 ;
        RECT 59.860 202.325 60.660 202.495 ;
        RECT 61.250 202.535 62.120 202.875 ;
        RECT 52.930 200.495 58.275 201.040 ;
        RECT 58.495 200.495 58.745 201.250 ;
        RECT 58.915 201.205 59.120 201.855 ;
        RECT 59.860 201.735 60.030 202.325 ;
        RECT 61.250 202.155 61.420 202.535 ;
        RECT 62.355 202.415 62.525 202.875 ;
        RECT 62.695 202.585 63.065 203.045 ;
        RECT 63.360 202.445 63.530 202.785 ;
        RECT 63.700 202.615 64.030 203.045 ;
        RECT 64.265 202.445 64.435 202.785 ;
        RECT 60.200 201.985 61.420 202.155 ;
        RECT 61.590 202.075 62.050 202.365 ;
        RECT 62.355 202.245 62.915 202.415 ;
        RECT 63.360 202.275 64.435 202.445 ;
        RECT 64.605 202.545 65.285 202.875 ;
        RECT 65.500 202.545 65.750 202.875 ;
        RECT 65.920 202.585 66.170 203.045 ;
        RECT 62.745 202.105 62.915 202.245 ;
        RECT 61.590 202.065 62.555 202.075 ;
        RECT 61.250 201.895 61.420 201.985 ;
        RECT 61.880 201.905 62.555 202.065 ;
        RECT 59.290 201.705 60.030 201.735 ;
        RECT 59.290 201.405 60.205 201.705 ;
        RECT 59.880 201.230 60.205 201.405 ;
        RECT 58.915 200.675 59.165 201.205 ;
        RECT 59.335 200.495 59.640 200.955 ;
        RECT 59.885 200.875 60.205 201.230 ;
        RECT 60.375 201.445 60.915 201.815 ;
        RECT 61.250 201.725 61.655 201.895 ;
        RECT 60.375 201.045 60.615 201.445 ;
        RECT 61.095 201.275 61.315 201.555 ;
        RECT 60.785 201.105 61.315 201.275 ;
        RECT 60.785 200.875 60.955 201.105 ;
        RECT 61.485 200.945 61.655 201.725 ;
        RECT 61.825 201.115 62.175 201.735 ;
        RECT 62.345 201.115 62.555 201.905 ;
        RECT 62.745 201.935 64.245 202.105 ;
        RECT 62.745 201.245 62.915 201.935 ;
        RECT 64.605 201.765 64.775 202.545 ;
        RECT 65.580 202.415 65.750 202.545 ;
        RECT 63.085 201.595 64.775 201.765 ;
        RECT 64.945 201.985 65.410 202.375 ;
        RECT 65.580 202.245 65.975 202.415 ;
        RECT 63.085 201.415 63.255 201.595 ;
        RECT 59.885 200.705 60.955 200.875 ;
        RECT 61.125 200.495 61.315 200.935 ;
        RECT 61.485 200.665 62.435 200.945 ;
        RECT 62.745 200.855 63.005 201.245 ;
        RECT 63.425 201.175 64.215 201.425 ;
        RECT 62.655 200.685 63.005 200.855 ;
        RECT 63.215 200.495 63.545 200.955 ;
        RECT 64.420 200.885 64.590 201.595 ;
        RECT 64.945 201.395 65.115 201.985 ;
        RECT 64.760 201.175 65.115 201.395 ;
        RECT 65.285 201.175 65.635 201.795 ;
        RECT 65.805 200.885 65.975 202.245 ;
        RECT 66.340 202.075 66.665 202.860 ;
        RECT 66.145 201.025 66.605 202.075 ;
        RECT 64.420 200.715 65.275 200.885 ;
        RECT 65.480 200.715 65.975 200.885 ;
        RECT 66.145 200.495 66.475 200.855 ;
        RECT 66.835 200.755 67.005 202.875 ;
        RECT 67.175 202.545 67.505 203.045 ;
        RECT 67.675 202.375 67.930 202.875 ;
        RECT 67.180 202.205 67.930 202.375 ;
        RECT 67.180 201.215 67.410 202.205 ;
        RECT 67.580 201.385 67.930 202.035 ;
        RECT 68.565 201.955 70.235 203.045 ;
        RECT 70.410 202.610 75.755 203.045 ;
        RECT 68.565 201.435 69.315 201.955 ;
        RECT 69.485 201.265 70.235 201.785 ;
        RECT 72.000 201.360 72.350 202.610 ;
        RECT 75.925 201.880 76.215 203.045 ;
        RECT 76.845 201.955 79.435 203.045 ;
        RECT 79.610 202.610 84.955 203.045 ;
        RECT 85.130 202.610 90.475 203.045 ;
        RECT 90.650 202.610 95.995 203.045 ;
        RECT 96.170 202.610 101.515 203.045 ;
        RECT 67.180 201.045 67.930 201.215 ;
        RECT 67.175 200.495 67.505 200.875 ;
        RECT 67.675 200.755 67.930 201.045 ;
        RECT 68.565 200.495 70.235 201.265 ;
        RECT 73.830 201.040 74.170 201.870 ;
        RECT 76.845 201.435 78.055 201.955 ;
        RECT 78.225 201.265 79.435 201.785 ;
        RECT 81.200 201.360 81.550 202.610 ;
        RECT 70.410 200.495 75.755 201.040 ;
        RECT 75.925 200.495 76.215 201.220 ;
        RECT 76.845 200.495 79.435 201.265 ;
        RECT 83.030 201.040 83.370 201.870 ;
        RECT 86.720 201.360 87.070 202.610 ;
        RECT 88.550 201.040 88.890 201.870 ;
        RECT 92.240 201.360 92.590 202.610 ;
        RECT 94.070 201.040 94.410 201.870 ;
        RECT 97.760 201.360 98.110 202.610 ;
        RECT 101.685 201.880 101.975 203.045 ;
        RECT 102.605 201.955 104.275 203.045 ;
        RECT 104.450 202.610 109.795 203.045 ;
        RECT 109.970 202.610 115.315 203.045 ;
        RECT 115.490 202.610 120.835 203.045 ;
        RECT 121.010 202.610 126.355 203.045 ;
        RECT 99.590 201.040 99.930 201.870 ;
        RECT 102.605 201.435 103.355 201.955 ;
        RECT 103.525 201.265 104.275 201.785 ;
        RECT 106.040 201.360 106.390 202.610 ;
        RECT 79.610 200.495 84.955 201.040 ;
        RECT 85.130 200.495 90.475 201.040 ;
        RECT 90.650 200.495 95.995 201.040 ;
        RECT 96.170 200.495 101.515 201.040 ;
        RECT 101.685 200.495 101.975 201.220 ;
        RECT 102.605 200.495 104.275 201.265 ;
        RECT 107.870 201.040 108.210 201.870 ;
        RECT 111.560 201.360 111.910 202.610 ;
        RECT 113.390 201.040 113.730 201.870 ;
        RECT 117.080 201.360 117.430 202.610 ;
        RECT 118.910 201.040 119.250 201.870 ;
        RECT 122.600 201.360 122.950 202.610 ;
        RECT 126.525 201.955 127.735 203.045 ;
        RECT 124.430 201.040 124.770 201.870 ;
        RECT 126.525 201.415 127.045 201.955 ;
        RECT 127.215 201.245 127.735 201.785 ;
        RECT 104.450 200.495 109.795 201.040 ;
        RECT 109.970 200.495 115.315 201.040 ;
        RECT 115.490 200.495 120.835 201.040 ;
        RECT 121.010 200.495 126.355 201.040 ;
        RECT 126.525 200.495 127.735 201.245 ;
        RECT 14.660 200.325 127.820 200.495 ;
        RECT 14.745 199.575 15.955 200.325 ;
        RECT 14.745 199.035 15.265 199.575 ;
        RECT 17.045 199.555 20.555 200.325 ;
        RECT 20.730 199.780 26.075 200.325 ;
        RECT 26.250 199.780 31.595 200.325 ;
        RECT 31.770 199.780 37.115 200.325 ;
        RECT 15.435 198.865 15.955 199.405 ;
        RECT 14.745 197.775 15.955 198.865 ;
        RECT 17.045 198.865 18.735 199.385 ;
        RECT 18.905 199.035 20.555 199.555 ;
        RECT 17.045 197.775 20.555 198.865 ;
        RECT 22.320 198.210 22.670 199.460 ;
        RECT 24.150 198.950 24.490 199.780 ;
        RECT 27.840 198.210 28.190 199.460 ;
        RECT 29.670 198.950 30.010 199.780 ;
        RECT 33.360 198.210 33.710 199.460 ;
        RECT 35.190 198.950 35.530 199.780 ;
        RECT 37.285 199.600 37.575 200.325 ;
        RECT 37.745 199.555 39.415 200.325 ;
        RECT 39.590 199.780 44.935 200.325 ;
        RECT 45.110 199.780 50.455 200.325 ;
        RECT 50.630 199.780 55.975 200.325 ;
        RECT 56.150 199.780 61.495 200.325 ;
        RECT 20.730 197.775 26.075 198.210 ;
        RECT 26.250 197.775 31.595 198.210 ;
        RECT 31.770 197.775 37.115 198.210 ;
        RECT 37.285 197.775 37.575 198.940 ;
        RECT 37.745 198.865 38.495 199.385 ;
        RECT 38.665 199.035 39.415 199.555 ;
        RECT 37.745 197.775 39.415 198.865 ;
        RECT 41.180 198.210 41.530 199.460 ;
        RECT 43.010 198.950 43.350 199.780 ;
        RECT 46.700 198.210 47.050 199.460 ;
        RECT 48.530 198.950 48.870 199.780 ;
        RECT 52.220 198.210 52.570 199.460 ;
        RECT 54.050 198.950 54.390 199.780 ;
        RECT 57.740 198.210 58.090 199.460 ;
        RECT 59.570 198.950 59.910 199.780 ;
        RECT 61.725 199.505 61.935 200.325 ;
        RECT 62.105 199.525 62.435 200.155 ;
        RECT 62.105 198.925 62.355 199.525 ;
        RECT 62.605 199.505 62.835 200.325 ;
        RECT 63.045 199.600 63.335 200.325 ;
        RECT 63.565 199.505 63.775 200.325 ;
        RECT 63.945 199.525 64.275 200.155 ;
        RECT 62.525 199.085 62.855 199.335 ;
        RECT 39.590 197.775 44.935 198.210 ;
        RECT 45.110 197.775 50.455 198.210 ;
        RECT 50.630 197.775 55.975 198.210 ;
        RECT 56.150 197.775 61.495 198.210 ;
        RECT 61.725 197.775 61.935 198.915 ;
        RECT 62.105 197.945 62.435 198.925 ;
        RECT 62.605 197.775 62.835 198.915 ;
        RECT 63.045 197.775 63.335 198.940 ;
        RECT 63.945 198.925 64.195 199.525 ;
        RECT 64.445 199.505 64.675 200.325 ;
        RECT 64.885 199.555 67.475 200.325 ;
        RECT 64.365 199.085 64.695 199.335 ;
        RECT 63.565 197.775 63.775 198.915 ;
        RECT 63.945 197.945 64.275 198.925 ;
        RECT 64.445 197.775 64.675 198.915 ;
        RECT 64.885 198.865 66.095 199.385 ;
        RECT 66.265 199.035 67.475 199.555 ;
        RECT 67.645 199.650 67.905 200.155 ;
        RECT 68.085 199.945 68.415 200.325 ;
        RECT 68.595 199.775 68.765 200.155 ;
        RECT 64.885 197.775 67.475 198.865 ;
        RECT 67.645 198.850 67.815 199.650 ;
        RECT 68.100 199.605 68.765 199.775 ;
        RECT 69.485 199.675 69.745 200.155 ;
        RECT 69.915 199.785 70.165 200.325 ;
        RECT 68.100 199.350 68.270 199.605 ;
        RECT 67.985 199.020 68.270 199.350 ;
        RECT 68.505 199.055 68.835 199.425 ;
        RECT 68.100 198.875 68.270 199.020 ;
        RECT 67.645 197.945 67.915 198.850 ;
        RECT 68.100 198.705 68.765 198.875 ;
        RECT 68.085 197.775 68.415 198.535 ;
        RECT 68.595 197.945 68.765 198.705 ;
        RECT 69.485 198.645 69.655 199.675 ;
        RECT 70.335 199.620 70.555 200.105 ;
        RECT 69.825 199.025 70.055 199.420 ;
        RECT 70.225 199.195 70.555 199.620 ;
        RECT 70.725 199.945 71.615 200.115 ;
        RECT 70.725 199.220 70.895 199.945 ;
        RECT 71.065 199.390 71.615 199.775 ;
        RECT 72.245 199.555 74.835 200.325 ;
        RECT 70.725 199.150 71.615 199.220 ;
        RECT 70.720 199.125 71.615 199.150 ;
        RECT 70.710 199.110 71.615 199.125 ;
        RECT 70.705 199.095 71.615 199.110 ;
        RECT 70.695 199.090 71.615 199.095 ;
        RECT 70.690 199.080 71.615 199.090 ;
        RECT 70.685 199.070 71.615 199.080 ;
        RECT 70.675 199.065 71.615 199.070 ;
        RECT 70.665 199.055 71.615 199.065 ;
        RECT 70.655 199.050 71.615 199.055 ;
        RECT 70.655 199.045 70.990 199.050 ;
        RECT 70.640 199.040 70.990 199.045 ;
        RECT 70.625 199.030 70.990 199.040 ;
        RECT 70.600 199.025 70.990 199.030 ;
        RECT 69.825 199.020 70.990 199.025 ;
        RECT 69.825 198.985 70.960 199.020 ;
        RECT 69.825 198.960 70.925 198.985 ;
        RECT 69.825 198.930 70.895 198.960 ;
        RECT 69.825 198.900 70.875 198.930 ;
        RECT 69.825 198.870 70.855 198.900 ;
        RECT 69.825 198.860 70.785 198.870 ;
        RECT 69.825 198.850 70.760 198.860 ;
        RECT 69.825 198.835 70.740 198.850 ;
        RECT 69.825 198.820 70.720 198.835 ;
        RECT 69.930 198.810 70.715 198.820 ;
        RECT 69.930 198.775 70.700 198.810 ;
        RECT 69.485 197.945 69.760 198.645 ;
        RECT 69.930 198.525 70.685 198.775 ;
        RECT 70.855 198.455 71.185 198.700 ;
        RECT 71.355 198.600 71.615 199.050 ;
        RECT 72.245 198.865 73.455 199.385 ;
        RECT 73.625 199.035 74.835 199.555 ;
        RECT 75.010 199.615 75.265 200.145 ;
        RECT 75.435 199.865 75.740 200.325 ;
        RECT 75.985 199.945 77.055 200.115 ;
        RECT 75.010 198.965 75.220 199.615 ;
        RECT 75.985 199.590 76.305 199.945 ;
        RECT 75.980 199.415 76.305 199.590 ;
        RECT 75.390 199.115 76.305 199.415 ;
        RECT 76.475 199.375 76.715 199.775 ;
        RECT 76.885 199.715 77.055 199.945 ;
        RECT 77.225 199.885 77.415 200.325 ;
        RECT 77.585 199.875 78.535 200.155 ;
        RECT 78.755 199.965 79.105 200.135 ;
        RECT 76.885 199.545 77.415 199.715 ;
        RECT 75.390 199.085 76.130 199.115 ;
        RECT 71.000 198.430 71.185 198.455 ;
        RECT 71.000 198.330 71.615 198.430 ;
        RECT 69.930 197.775 70.185 198.320 ;
        RECT 70.355 197.945 70.835 198.285 ;
        RECT 71.010 197.775 71.615 198.330 ;
        RECT 72.245 197.775 74.835 198.865 ;
        RECT 75.010 198.085 75.265 198.965 ;
        RECT 75.435 197.775 75.740 198.915 ;
        RECT 75.960 198.495 76.130 199.085 ;
        RECT 76.475 199.005 77.015 199.375 ;
        RECT 77.195 199.265 77.415 199.545 ;
        RECT 77.585 199.095 77.755 199.875 ;
        RECT 77.350 198.925 77.755 199.095 ;
        RECT 77.925 199.085 78.275 199.705 ;
        RECT 77.350 198.835 77.520 198.925 ;
        RECT 78.445 198.915 78.655 199.705 ;
        RECT 76.300 198.665 77.520 198.835 ;
        RECT 77.980 198.755 78.655 198.915 ;
        RECT 75.960 198.325 76.760 198.495 ;
        RECT 76.080 197.775 76.410 198.155 ;
        RECT 76.590 198.035 76.760 198.325 ;
        RECT 77.350 198.285 77.520 198.665 ;
        RECT 77.690 198.745 78.655 198.755 ;
        RECT 78.845 199.575 79.105 199.965 ;
        RECT 79.315 199.865 79.645 200.325 ;
        RECT 80.520 199.935 81.375 200.105 ;
        RECT 81.580 199.935 82.075 200.105 ;
        RECT 82.245 199.965 82.575 200.325 ;
        RECT 78.845 198.885 79.015 199.575 ;
        RECT 79.185 199.225 79.355 199.405 ;
        RECT 79.525 199.395 80.315 199.645 ;
        RECT 80.520 199.225 80.690 199.935 ;
        RECT 80.860 199.425 81.215 199.645 ;
        RECT 79.185 199.055 80.875 199.225 ;
        RECT 77.690 198.455 78.150 198.745 ;
        RECT 78.845 198.715 80.345 198.885 ;
        RECT 78.845 198.575 79.015 198.715 ;
        RECT 78.455 198.405 79.015 198.575 ;
        RECT 76.930 197.775 77.180 198.235 ;
        RECT 77.350 197.945 78.220 198.285 ;
        RECT 78.455 197.945 78.625 198.405 ;
        RECT 79.460 198.375 80.535 198.545 ;
        RECT 78.795 197.775 79.165 198.235 ;
        RECT 79.460 198.035 79.630 198.375 ;
        RECT 79.800 197.775 80.130 198.205 ;
        RECT 80.365 198.035 80.535 198.375 ;
        RECT 80.705 198.275 80.875 199.055 ;
        RECT 81.045 198.835 81.215 199.425 ;
        RECT 81.385 199.025 81.735 199.645 ;
        RECT 81.045 198.445 81.510 198.835 ;
        RECT 81.905 198.575 82.075 199.935 ;
        RECT 82.245 198.745 82.705 199.795 ;
        RECT 81.680 198.405 82.075 198.575 ;
        RECT 81.680 198.275 81.850 198.405 ;
        RECT 80.705 197.945 81.385 198.275 ;
        RECT 81.600 197.945 81.850 198.275 ;
        RECT 82.020 197.775 82.270 198.235 ;
        RECT 82.440 197.960 82.765 198.745 ;
        RECT 82.935 197.945 83.105 200.065 ;
        RECT 83.275 199.945 83.605 200.325 ;
        RECT 83.775 199.775 84.030 200.065 ;
        RECT 83.280 199.605 84.030 199.775 ;
        RECT 83.280 198.615 83.510 199.605 ;
        RECT 85.125 199.555 88.635 200.325 ;
        RECT 88.805 199.600 89.095 200.325 ;
        RECT 89.265 199.555 92.775 200.325 ;
        RECT 92.950 199.780 98.295 200.325 ;
        RECT 98.470 199.780 103.815 200.325 ;
        RECT 103.990 199.780 109.335 200.325 ;
        RECT 83.680 198.785 84.030 199.435 ;
        RECT 85.125 198.865 86.815 199.385 ;
        RECT 86.985 199.035 88.635 199.555 ;
        RECT 83.280 198.445 84.030 198.615 ;
        RECT 83.275 197.775 83.605 198.275 ;
        RECT 83.775 197.945 84.030 198.445 ;
        RECT 85.125 197.775 88.635 198.865 ;
        RECT 88.805 197.775 89.095 198.940 ;
        RECT 89.265 198.865 90.955 199.385 ;
        RECT 91.125 199.035 92.775 199.555 ;
        RECT 89.265 197.775 92.775 198.865 ;
        RECT 94.540 198.210 94.890 199.460 ;
        RECT 96.370 198.950 96.710 199.780 ;
        RECT 100.060 198.210 100.410 199.460 ;
        RECT 101.890 198.950 102.230 199.780 ;
        RECT 105.580 198.210 105.930 199.460 ;
        RECT 107.410 198.950 107.750 199.780 ;
        RECT 109.565 199.505 109.775 200.325 ;
        RECT 109.945 199.525 110.275 200.155 ;
        RECT 109.945 198.925 110.195 199.525 ;
        RECT 110.445 199.505 110.675 200.325 ;
        RECT 111.345 199.555 113.015 200.325 ;
        RECT 110.365 199.085 110.695 199.335 ;
        RECT 92.950 197.775 98.295 198.210 ;
        RECT 98.470 197.775 103.815 198.210 ;
        RECT 103.990 197.775 109.335 198.210 ;
        RECT 109.565 197.775 109.775 198.915 ;
        RECT 109.945 197.945 110.275 198.925 ;
        RECT 110.445 197.775 110.675 198.915 ;
        RECT 111.345 198.865 112.095 199.385 ;
        RECT 112.265 199.035 113.015 199.555 ;
        RECT 113.225 199.505 113.455 200.325 ;
        RECT 113.625 199.525 113.955 200.155 ;
        RECT 113.205 199.085 113.535 199.335 ;
        RECT 113.705 198.925 113.955 199.525 ;
        RECT 114.125 199.505 114.335 200.325 ;
        RECT 114.565 199.600 114.855 200.325 ;
        RECT 115.490 199.780 120.835 200.325 ;
        RECT 121.010 199.780 126.355 200.325 ;
        RECT 111.345 197.775 113.015 198.865 ;
        RECT 113.225 197.775 113.455 198.915 ;
        RECT 113.625 197.945 113.955 198.925 ;
        RECT 114.125 197.775 114.335 198.915 ;
        RECT 114.565 197.775 114.855 198.940 ;
        RECT 117.080 198.210 117.430 199.460 ;
        RECT 118.910 198.950 119.250 199.780 ;
        RECT 122.600 198.210 122.950 199.460 ;
        RECT 124.430 198.950 124.770 199.780 ;
        RECT 126.525 199.575 127.735 200.325 ;
        RECT 126.525 198.865 127.045 199.405 ;
        RECT 127.215 199.035 127.735 199.575 ;
        RECT 115.490 197.775 120.835 198.210 ;
        RECT 121.010 197.775 126.355 198.210 ;
        RECT 126.525 197.775 127.735 198.865 ;
        RECT 14.660 197.605 127.820 197.775 ;
        RECT 14.745 196.515 15.955 197.605 ;
        RECT 14.745 195.805 15.265 196.345 ;
        RECT 15.435 195.975 15.955 196.515 ;
        RECT 16.125 196.515 18.715 197.605 ;
        RECT 18.890 197.170 24.235 197.605 ;
        RECT 16.125 195.995 17.335 196.515 ;
        RECT 17.505 195.825 18.715 196.345 ;
        RECT 20.480 195.920 20.830 197.170 ;
        RECT 24.405 196.440 24.695 197.605 ;
        RECT 25.790 197.170 31.135 197.605 ;
        RECT 31.310 197.170 36.655 197.605 ;
        RECT 36.830 197.170 42.175 197.605 ;
        RECT 14.745 195.055 15.955 195.805 ;
        RECT 16.125 195.055 18.715 195.825 ;
        RECT 22.310 195.600 22.650 196.430 ;
        RECT 27.380 195.920 27.730 197.170 ;
        RECT 18.890 195.055 24.235 195.600 ;
        RECT 24.405 195.055 24.695 195.780 ;
        RECT 29.210 195.600 29.550 196.430 ;
        RECT 32.900 195.920 33.250 197.170 ;
        RECT 34.730 195.600 35.070 196.430 ;
        RECT 38.420 195.920 38.770 197.170 ;
        RECT 42.405 196.465 42.615 197.605 ;
        RECT 42.785 196.455 43.115 197.435 ;
        RECT 43.285 196.465 43.515 197.605 ;
        RECT 44.650 197.170 49.995 197.605 ;
        RECT 40.250 195.600 40.590 196.430 ;
        RECT 25.790 195.055 31.135 195.600 ;
        RECT 31.310 195.055 36.655 195.600 ;
        RECT 36.830 195.055 42.175 195.600 ;
        RECT 42.405 195.055 42.615 195.875 ;
        RECT 42.785 195.855 43.035 196.455 ;
        RECT 43.205 196.045 43.535 196.295 ;
        RECT 46.240 195.920 46.590 197.170 ;
        RECT 50.165 196.440 50.455 197.605 ;
        RECT 51.085 196.515 52.755 197.605 ;
        RECT 52.930 197.170 58.275 197.605 ;
        RECT 42.785 195.225 43.115 195.855 ;
        RECT 43.285 195.055 43.515 195.875 ;
        RECT 48.070 195.600 48.410 196.430 ;
        RECT 51.085 195.995 51.835 196.515 ;
        RECT 52.005 195.825 52.755 196.345 ;
        RECT 54.520 195.920 54.870 197.170 ;
        RECT 58.755 196.765 58.925 197.605 ;
        RECT 59.135 196.595 59.385 197.435 ;
        RECT 59.595 196.765 59.765 197.605 ;
        RECT 59.935 196.595 60.225 197.435 ;
        RECT 44.650 195.055 49.995 195.600 ;
        RECT 50.165 195.055 50.455 195.780 ;
        RECT 51.085 195.055 52.755 195.825 ;
        RECT 56.350 195.600 56.690 196.430 ;
        RECT 58.500 196.425 60.225 196.595 ;
        RECT 60.435 196.545 60.605 197.605 ;
        RECT 60.900 197.225 61.230 197.605 ;
        RECT 61.410 197.055 61.580 197.345 ;
        RECT 61.750 197.145 62.000 197.605 ;
        RECT 60.780 196.885 61.580 197.055 ;
        RECT 62.170 197.095 63.040 197.435 ;
        RECT 58.500 195.875 58.910 196.425 ;
        RECT 60.780 196.265 60.950 196.885 ;
        RECT 62.170 196.715 62.340 197.095 ;
        RECT 63.275 196.975 63.445 197.435 ;
        RECT 63.615 197.145 63.985 197.605 ;
        RECT 64.280 197.005 64.450 197.345 ;
        RECT 64.620 197.175 64.950 197.605 ;
        RECT 65.185 197.005 65.355 197.345 ;
        RECT 61.120 196.545 62.340 196.715 ;
        RECT 62.510 196.635 62.970 196.925 ;
        RECT 63.275 196.805 63.835 196.975 ;
        RECT 64.280 196.835 65.355 197.005 ;
        RECT 65.525 197.105 66.205 197.435 ;
        RECT 66.420 197.105 66.670 197.435 ;
        RECT 66.840 197.145 67.090 197.605 ;
        RECT 63.665 196.665 63.835 196.805 ;
        RECT 62.510 196.625 63.475 196.635 ;
        RECT 62.170 196.455 62.340 196.545 ;
        RECT 62.800 196.465 63.475 196.625 ;
        RECT 60.780 196.255 61.125 196.265 ;
        RECT 59.095 196.045 61.125 196.255 ;
        RECT 58.500 195.705 60.265 195.875 ;
        RECT 52.930 195.055 58.275 195.600 ;
        RECT 58.755 195.055 58.925 195.525 ;
        RECT 59.095 195.225 59.425 195.705 ;
        RECT 59.595 195.055 59.765 195.525 ;
        RECT 59.935 195.225 60.265 195.705 ;
        RECT 60.435 195.055 60.605 195.865 ;
        RECT 60.800 195.790 61.125 196.045 ;
        RECT 60.805 195.435 61.125 195.790 ;
        RECT 61.295 196.005 61.835 196.375 ;
        RECT 62.170 196.285 62.575 196.455 ;
        RECT 61.295 195.605 61.535 196.005 ;
        RECT 62.015 195.835 62.235 196.115 ;
        RECT 61.705 195.665 62.235 195.835 ;
        RECT 61.705 195.435 61.875 195.665 ;
        RECT 62.405 195.505 62.575 196.285 ;
        RECT 62.745 195.675 63.095 196.295 ;
        RECT 63.265 195.675 63.475 196.465 ;
        RECT 63.665 196.495 65.165 196.665 ;
        RECT 63.665 195.805 63.835 196.495 ;
        RECT 65.525 196.325 65.695 197.105 ;
        RECT 66.500 196.975 66.670 197.105 ;
        RECT 64.005 196.155 65.695 196.325 ;
        RECT 65.865 196.545 66.330 196.935 ;
        RECT 66.500 196.805 66.895 196.975 ;
        RECT 64.005 195.975 64.175 196.155 ;
        RECT 60.805 195.265 61.875 195.435 ;
        RECT 62.045 195.055 62.235 195.495 ;
        RECT 62.405 195.225 63.355 195.505 ;
        RECT 63.665 195.415 63.925 195.805 ;
        RECT 64.345 195.735 65.135 195.985 ;
        RECT 63.575 195.245 63.925 195.415 ;
        RECT 64.135 195.055 64.465 195.515 ;
        RECT 65.340 195.445 65.510 196.155 ;
        RECT 65.865 195.955 66.035 196.545 ;
        RECT 65.680 195.735 66.035 195.955 ;
        RECT 66.205 195.735 66.555 196.355 ;
        RECT 66.725 195.445 66.895 196.805 ;
        RECT 67.260 196.635 67.585 197.420 ;
        RECT 67.065 195.585 67.525 196.635 ;
        RECT 65.340 195.275 66.195 195.445 ;
        RECT 66.400 195.275 66.895 195.445 ;
        RECT 67.065 195.055 67.395 195.415 ;
        RECT 67.755 195.315 67.925 197.435 ;
        RECT 68.095 197.105 68.425 197.605 ;
        RECT 68.595 196.935 68.850 197.435 ;
        RECT 69.045 197.095 69.345 197.605 ;
        RECT 69.515 197.095 69.895 197.265 ;
        RECT 70.475 197.095 71.105 197.605 ;
        RECT 68.100 196.765 68.850 196.935 ;
        RECT 69.515 196.925 69.685 197.095 ;
        RECT 71.275 196.925 71.605 197.435 ;
        RECT 71.775 197.095 72.075 197.605 ;
        RECT 68.100 195.775 68.330 196.765 ;
        RECT 69.025 196.725 69.685 196.925 ;
        RECT 69.855 196.755 72.075 196.925 ;
        RECT 68.500 195.945 68.850 196.595 ;
        RECT 69.025 195.795 69.195 196.725 ;
        RECT 69.855 196.555 70.025 196.755 ;
        RECT 69.365 196.385 70.025 196.555 ;
        RECT 70.195 196.415 71.735 196.585 ;
        RECT 69.365 195.965 69.535 196.385 ;
        RECT 70.195 196.215 70.365 196.415 ;
        RECT 69.765 196.045 70.365 196.215 ;
        RECT 70.535 196.045 71.230 196.245 ;
        RECT 71.490 195.965 71.735 196.415 ;
        RECT 69.855 195.795 70.765 195.875 ;
        RECT 68.100 195.605 68.850 195.775 ;
        RECT 68.095 195.055 68.425 195.435 ;
        RECT 68.595 195.315 68.850 195.605 ;
        RECT 69.025 195.315 69.345 195.795 ;
        RECT 69.515 195.705 70.765 195.795 ;
        RECT 69.515 195.625 70.025 195.705 ;
        RECT 69.515 195.225 69.745 195.625 ;
        RECT 69.915 195.055 70.265 195.445 ;
        RECT 70.435 195.225 70.765 195.705 ;
        RECT 70.935 195.055 71.105 195.875 ;
        RECT 71.905 195.795 72.075 196.755 ;
        RECT 72.245 196.515 75.755 197.605 ;
        RECT 72.245 195.995 73.935 196.515 ;
        RECT 75.925 196.440 76.215 197.605 ;
        RECT 76.885 196.465 77.115 197.605 ;
        RECT 77.285 196.455 77.615 197.435 ;
        RECT 77.785 196.465 77.995 197.605 ;
        RECT 78.225 197.095 78.525 197.605 ;
        RECT 78.695 196.925 79.025 197.435 ;
        RECT 79.195 197.095 79.825 197.605 ;
        RECT 80.405 197.095 80.785 197.265 ;
        RECT 80.955 197.095 81.255 197.605 ;
        RECT 80.615 196.925 80.785 197.095 ;
        RECT 78.225 196.755 80.445 196.925 ;
        RECT 74.105 195.825 75.755 196.345 ;
        RECT 76.865 196.045 77.195 196.295 ;
        RECT 71.610 195.250 72.075 195.795 ;
        RECT 72.245 195.055 75.755 195.825 ;
        RECT 75.925 195.055 76.215 195.780 ;
        RECT 76.885 195.055 77.115 195.875 ;
        RECT 77.365 195.855 77.615 196.455 ;
        RECT 77.285 195.225 77.615 195.855 ;
        RECT 77.785 195.055 77.995 195.875 ;
        RECT 78.225 195.795 78.395 196.755 ;
        RECT 78.565 196.415 80.105 196.585 ;
        RECT 78.565 195.965 78.810 196.415 ;
        RECT 79.070 196.045 79.765 196.245 ;
        RECT 79.935 196.215 80.105 196.415 ;
        RECT 80.275 196.555 80.445 196.755 ;
        RECT 80.615 196.725 81.275 196.925 ;
        RECT 80.275 196.385 80.935 196.555 ;
        RECT 79.935 196.045 80.535 196.215 ;
        RECT 80.765 195.965 80.935 196.385 ;
        RECT 78.225 195.250 78.690 195.795 ;
        RECT 79.195 195.055 79.365 195.875 ;
        RECT 79.535 195.795 80.445 195.875 ;
        RECT 81.105 195.795 81.275 196.725 ;
        RECT 81.445 196.515 84.955 197.605 ;
        RECT 85.500 196.625 85.755 197.295 ;
        RECT 85.935 196.805 86.220 197.605 ;
        RECT 86.400 196.885 86.730 197.395 ;
        RECT 81.445 195.995 83.135 196.515 ;
        RECT 83.305 195.825 84.955 196.345 ;
        RECT 79.535 195.705 80.785 195.795 ;
        RECT 79.535 195.225 79.865 195.705 ;
        RECT 80.275 195.625 80.785 195.705 ;
        RECT 80.035 195.055 80.385 195.445 ;
        RECT 80.555 195.225 80.785 195.625 ;
        RECT 80.955 195.315 81.275 195.795 ;
        RECT 81.445 195.055 84.955 195.825 ;
        RECT 85.500 195.765 85.680 196.625 ;
        RECT 86.400 196.295 86.650 196.885 ;
        RECT 87.000 196.735 87.170 197.345 ;
        RECT 87.340 196.915 87.670 197.605 ;
        RECT 87.900 197.055 88.140 197.345 ;
        RECT 88.340 197.225 88.760 197.605 ;
        RECT 88.940 197.135 89.570 197.385 ;
        RECT 90.040 197.225 90.370 197.605 ;
        RECT 88.940 197.055 89.110 197.135 ;
        RECT 90.540 197.055 90.710 197.345 ;
        RECT 90.890 197.225 91.270 197.605 ;
        RECT 91.510 197.220 92.340 197.390 ;
        RECT 87.900 196.885 89.110 197.055 ;
        RECT 85.850 195.965 86.650 196.295 ;
        RECT 85.500 195.565 85.755 195.765 ;
        RECT 85.415 195.395 85.755 195.565 ;
        RECT 85.500 195.235 85.755 195.395 ;
        RECT 85.935 195.055 86.220 195.515 ;
        RECT 86.400 195.315 86.650 195.965 ;
        RECT 86.850 196.715 87.170 196.735 ;
        RECT 86.850 196.545 88.770 196.715 ;
        RECT 86.850 195.650 87.040 196.545 ;
        RECT 88.940 196.375 89.110 196.885 ;
        RECT 89.280 196.625 89.800 196.935 ;
        RECT 87.210 196.205 89.110 196.375 ;
        RECT 87.210 196.145 87.540 196.205 ;
        RECT 87.690 195.975 88.020 196.035 ;
        RECT 87.360 195.705 88.020 195.975 ;
        RECT 86.850 195.320 87.170 195.650 ;
        RECT 87.350 195.055 88.010 195.535 ;
        RECT 88.210 195.445 88.380 196.205 ;
        RECT 89.280 196.035 89.460 196.445 ;
        RECT 88.550 195.865 88.880 195.985 ;
        RECT 89.630 195.865 89.800 196.625 ;
        RECT 88.550 195.695 89.800 195.865 ;
        RECT 89.970 196.805 91.340 197.055 ;
        RECT 89.970 196.035 90.160 196.805 ;
        RECT 91.090 196.545 91.340 196.805 ;
        RECT 90.330 196.375 90.580 196.535 ;
        RECT 91.510 196.375 91.680 197.220 ;
        RECT 92.575 196.935 92.745 197.435 ;
        RECT 92.915 197.105 93.245 197.605 ;
        RECT 91.850 196.545 92.350 196.925 ;
        RECT 92.575 196.765 93.270 196.935 ;
        RECT 90.330 196.205 91.680 196.375 ;
        RECT 91.260 196.165 91.680 196.205 ;
        RECT 89.970 195.695 90.390 196.035 ;
        RECT 90.680 195.705 91.090 196.035 ;
        RECT 88.210 195.275 89.060 195.445 ;
        RECT 89.620 195.055 89.940 195.515 ;
        RECT 90.140 195.265 90.390 195.695 ;
        RECT 90.680 195.055 91.090 195.495 ;
        RECT 91.260 195.435 91.430 196.165 ;
        RECT 91.600 195.615 91.950 195.985 ;
        RECT 92.130 195.675 92.350 196.545 ;
        RECT 92.520 195.975 92.930 196.595 ;
        RECT 93.100 195.795 93.270 196.765 ;
        RECT 92.575 195.605 93.270 195.795 ;
        RECT 91.260 195.235 92.275 195.435 ;
        RECT 92.575 195.275 92.745 195.605 ;
        RECT 92.915 195.055 93.245 195.435 ;
        RECT 93.460 195.315 93.685 197.435 ;
        RECT 93.855 197.105 94.185 197.605 ;
        RECT 94.355 196.935 94.525 197.435 ;
        RECT 94.790 197.170 100.135 197.605 ;
        RECT 93.860 196.765 94.525 196.935 ;
        RECT 93.860 195.775 94.090 196.765 ;
        RECT 94.260 195.945 94.610 196.595 ;
        RECT 96.380 195.920 96.730 197.170 ;
        RECT 100.395 196.675 100.565 197.435 ;
        RECT 100.745 196.845 101.075 197.605 ;
        RECT 100.395 196.505 101.060 196.675 ;
        RECT 101.245 196.530 101.515 197.435 ;
        RECT 93.860 195.605 94.525 195.775 ;
        RECT 93.855 195.055 94.185 195.435 ;
        RECT 94.355 195.315 94.525 195.605 ;
        RECT 98.210 195.600 98.550 196.430 ;
        RECT 100.890 196.360 101.060 196.505 ;
        RECT 100.325 195.955 100.655 196.325 ;
        RECT 100.890 196.030 101.175 196.360 ;
        RECT 100.890 195.775 101.060 196.030 ;
        RECT 100.395 195.605 101.060 195.775 ;
        RECT 101.345 195.730 101.515 196.530 ;
        RECT 101.685 196.440 101.975 197.605 ;
        RECT 102.605 196.515 106.115 197.605 ;
        RECT 102.605 195.995 104.295 196.515 ;
        RECT 106.290 196.415 106.545 197.295 ;
        RECT 106.715 196.465 107.020 197.605 ;
        RECT 107.360 197.225 107.690 197.605 ;
        RECT 107.870 197.055 108.040 197.345 ;
        RECT 108.210 197.145 108.460 197.605 ;
        RECT 107.240 196.885 108.040 197.055 ;
        RECT 108.630 197.095 109.500 197.435 ;
        RECT 104.465 195.825 106.115 196.345 ;
        RECT 94.790 195.055 100.135 195.600 ;
        RECT 100.395 195.225 100.565 195.605 ;
        RECT 100.745 195.055 101.075 195.435 ;
        RECT 101.255 195.225 101.515 195.730 ;
        RECT 101.685 195.055 101.975 195.780 ;
        RECT 102.605 195.055 106.115 195.825 ;
        RECT 106.290 195.765 106.500 196.415 ;
        RECT 107.240 196.295 107.410 196.885 ;
        RECT 108.630 196.715 108.800 197.095 ;
        RECT 109.735 196.975 109.905 197.435 ;
        RECT 110.075 197.145 110.445 197.605 ;
        RECT 110.740 197.005 110.910 197.345 ;
        RECT 111.080 197.175 111.410 197.605 ;
        RECT 111.645 197.005 111.815 197.345 ;
        RECT 107.580 196.545 108.800 196.715 ;
        RECT 108.970 196.635 109.430 196.925 ;
        RECT 109.735 196.805 110.295 196.975 ;
        RECT 110.740 196.835 111.815 197.005 ;
        RECT 111.985 197.105 112.665 197.435 ;
        RECT 112.880 197.105 113.130 197.435 ;
        RECT 113.300 197.145 113.550 197.605 ;
        RECT 110.125 196.665 110.295 196.805 ;
        RECT 108.970 196.625 109.935 196.635 ;
        RECT 108.630 196.455 108.800 196.545 ;
        RECT 109.260 196.465 109.935 196.625 ;
        RECT 106.670 196.265 107.410 196.295 ;
        RECT 106.670 195.965 107.585 196.265 ;
        RECT 107.260 195.790 107.585 195.965 ;
        RECT 106.290 195.235 106.545 195.765 ;
        RECT 106.715 195.055 107.020 195.515 ;
        RECT 107.265 195.435 107.585 195.790 ;
        RECT 107.755 196.005 108.295 196.375 ;
        RECT 108.630 196.285 109.035 196.455 ;
        RECT 107.755 195.605 107.995 196.005 ;
        RECT 108.475 195.835 108.695 196.115 ;
        RECT 108.165 195.665 108.695 195.835 ;
        RECT 108.165 195.435 108.335 195.665 ;
        RECT 108.865 195.505 109.035 196.285 ;
        RECT 109.205 195.675 109.555 196.295 ;
        RECT 109.725 195.675 109.935 196.465 ;
        RECT 110.125 196.495 111.625 196.665 ;
        RECT 110.125 195.805 110.295 196.495 ;
        RECT 111.985 196.325 112.155 197.105 ;
        RECT 112.960 196.975 113.130 197.105 ;
        RECT 110.465 196.155 112.155 196.325 ;
        RECT 112.325 196.545 112.790 196.935 ;
        RECT 112.960 196.805 113.355 196.975 ;
        RECT 110.465 195.975 110.635 196.155 ;
        RECT 107.265 195.265 108.335 195.435 ;
        RECT 108.505 195.055 108.695 195.495 ;
        RECT 108.865 195.225 109.815 195.505 ;
        RECT 110.125 195.415 110.385 195.805 ;
        RECT 110.805 195.735 111.595 195.985 ;
        RECT 110.035 195.245 110.385 195.415 ;
        RECT 110.595 195.055 110.925 195.515 ;
        RECT 111.800 195.445 111.970 196.155 ;
        RECT 112.325 195.955 112.495 196.545 ;
        RECT 112.140 195.735 112.495 195.955 ;
        RECT 112.665 195.735 113.015 196.355 ;
        RECT 113.185 195.445 113.355 196.805 ;
        RECT 113.720 196.635 114.045 197.420 ;
        RECT 113.525 195.585 113.985 196.635 ;
        RECT 111.800 195.275 112.655 195.445 ;
        RECT 112.860 195.275 113.355 195.445 ;
        RECT 113.525 195.055 113.855 195.415 ;
        RECT 114.215 195.315 114.385 197.435 ;
        RECT 114.555 197.105 114.885 197.605 ;
        RECT 115.055 196.935 115.310 197.435 ;
        RECT 114.560 196.765 115.310 196.935 ;
        RECT 114.560 195.775 114.790 196.765 ;
        RECT 114.960 195.945 115.310 196.595 ;
        RECT 115.490 196.415 115.745 197.295 ;
        RECT 115.915 196.465 116.220 197.605 ;
        RECT 116.560 197.225 116.890 197.605 ;
        RECT 117.070 197.055 117.240 197.345 ;
        RECT 117.410 197.145 117.660 197.605 ;
        RECT 116.440 196.885 117.240 197.055 ;
        RECT 117.830 197.095 118.700 197.435 ;
        RECT 114.560 195.605 115.310 195.775 ;
        RECT 114.555 195.055 114.885 195.435 ;
        RECT 115.055 195.315 115.310 195.605 ;
        RECT 115.490 195.765 115.700 196.415 ;
        RECT 116.440 196.295 116.610 196.885 ;
        RECT 117.830 196.715 118.000 197.095 ;
        RECT 118.935 196.975 119.105 197.435 ;
        RECT 119.275 197.145 119.645 197.605 ;
        RECT 119.940 197.005 120.110 197.345 ;
        RECT 120.280 197.175 120.610 197.605 ;
        RECT 120.845 197.005 121.015 197.345 ;
        RECT 116.780 196.545 118.000 196.715 ;
        RECT 118.170 196.635 118.630 196.925 ;
        RECT 118.935 196.805 119.495 196.975 ;
        RECT 119.940 196.835 121.015 197.005 ;
        RECT 121.185 197.105 121.865 197.435 ;
        RECT 122.080 197.105 122.330 197.435 ;
        RECT 122.500 197.145 122.750 197.605 ;
        RECT 119.325 196.665 119.495 196.805 ;
        RECT 118.170 196.625 119.135 196.635 ;
        RECT 117.830 196.455 118.000 196.545 ;
        RECT 118.460 196.465 119.135 196.625 ;
        RECT 115.870 196.265 116.610 196.295 ;
        RECT 115.870 195.965 116.785 196.265 ;
        RECT 116.460 195.790 116.785 195.965 ;
        RECT 115.490 195.235 115.745 195.765 ;
        RECT 115.915 195.055 116.220 195.515 ;
        RECT 116.465 195.435 116.785 195.790 ;
        RECT 116.955 196.005 117.495 196.375 ;
        RECT 117.830 196.285 118.235 196.455 ;
        RECT 116.955 195.605 117.195 196.005 ;
        RECT 117.675 195.835 117.895 196.115 ;
        RECT 117.365 195.665 117.895 195.835 ;
        RECT 117.365 195.435 117.535 195.665 ;
        RECT 118.065 195.505 118.235 196.285 ;
        RECT 118.405 195.675 118.755 196.295 ;
        RECT 118.925 195.675 119.135 196.465 ;
        RECT 119.325 196.495 120.825 196.665 ;
        RECT 119.325 195.805 119.495 196.495 ;
        RECT 121.185 196.325 121.355 197.105 ;
        RECT 122.160 196.975 122.330 197.105 ;
        RECT 119.665 196.155 121.355 196.325 ;
        RECT 121.525 196.545 121.990 196.935 ;
        RECT 122.160 196.805 122.555 196.975 ;
        RECT 119.665 195.975 119.835 196.155 ;
        RECT 116.465 195.265 117.535 195.435 ;
        RECT 117.705 195.055 117.895 195.495 ;
        RECT 118.065 195.225 119.015 195.505 ;
        RECT 119.325 195.415 119.585 195.805 ;
        RECT 120.005 195.735 120.795 195.985 ;
        RECT 119.235 195.245 119.585 195.415 ;
        RECT 119.795 195.055 120.125 195.515 ;
        RECT 121.000 195.445 121.170 196.155 ;
        RECT 121.525 195.955 121.695 196.545 ;
        RECT 121.340 195.735 121.695 195.955 ;
        RECT 121.865 195.735 122.215 196.355 ;
        RECT 122.385 195.445 122.555 196.805 ;
        RECT 122.920 196.635 123.245 197.420 ;
        RECT 122.725 195.585 123.185 196.635 ;
        RECT 121.000 195.275 121.855 195.445 ;
        RECT 122.060 195.275 122.555 195.445 ;
        RECT 122.725 195.055 123.055 195.415 ;
        RECT 123.415 195.315 123.585 197.435 ;
        RECT 123.755 197.105 124.085 197.605 ;
        RECT 124.255 196.935 124.510 197.435 ;
        RECT 123.760 196.765 124.510 196.935 ;
        RECT 123.760 195.775 123.990 196.765 ;
        RECT 124.160 195.945 124.510 196.595 ;
        RECT 124.685 196.515 126.355 197.605 ;
        RECT 126.525 196.515 127.735 197.605 ;
        RECT 124.685 195.995 125.435 196.515 ;
        RECT 125.605 195.825 126.355 196.345 ;
        RECT 126.525 195.975 127.045 196.515 ;
        RECT 123.760 195.605 124.510 195.775 ;
        RECT 123.755 195.055 124.085 195.435 ;
        RECT 124.255 195.315 124.510 195.605 ;
        RECT 124.685 195.055 126.355 195.825 ;
        RECT 127.215 195.805 127.735 196.345 ;
        RECT 126.525 195.055 127.735 195.805 ;
        RECT 14.660 194.885 127.820 195.055 ;
        RECT 14.745 194.135 15.955 194.885 ;
        RECT 14.745 193.595 15.265 194.135 ;
        RECT 17.045 194.115 20.555 194.885 ;
        RECT 20.730 194.340 26.075 194.885 ;
        RECT 26.250 194.340 31.595 194.885 ;
        RECT 31.770 194.340 37.115 194.885 ;
        RECT 15.435 193.425 15.955 193.965 ;
        RECT 14.745 192.335 15.955 193.425 ;
        RECT 17.045 193.425 18.735 193.945 ;
        RECT 18.905 193.595 20.555 194.115 ;
        RECT 17.045 192.335 20.555 193.425 ;
        RECT 22.320 192.770 22.670 194.020 ;
        RECT 24.150 193.510 24.490 194.340 ;
        RECT 27.840 192.770 28.190 194.020 ;
        RECT 29.670 193.510 30.010 194.340 ;
        RECT 33.360 192.770 33.710 194.020 ;
        RECT 35.190 193.510 35.530 194.340 ;
        RECT 37.285 194.160 37.575 194.885 ;
        RECT 37.750 194.335 38.005 194.625 ;
        RECT 38.175 194.505 38.505 194.885 ;
        RECT 37.750 194.165 38.500 194.335 ;
        RECT 20.730 192.335 26.075 192.770 ;
        RECT 26.250 192.335 31.595 192.770 ;
        RECT 31.770 192.335 37.115 192.770 ;
        RECT 37.285 192.335 37.575 193.500 ;
        RECT 37.750 193.345 38.100 193.995 ;
        RECT 38.270 193.175 38.500 194.165 ;
        RECT 37.750 193.005 38.500 193.175 ;
        RECT 37.750 192.505 38.005 193.005 ;
        RECT 38.175 192.335 38.505 192.835 ;
        RECT 38.675 192.505 38.845 194.625 ;
        RECT 39.205 194.525 39.535 194.885 ;
        RECT 39.705 194.495 40.200 194.665 ;
        RECT 40.405 194.495 41.260 194.665 ;
        RECT 39.075 193.305 39.535 194.355 ;
        RECT 39.015 192.520 39.340 193.305 ;
        RECT 39.705 193.135 39.875 194.495 ;
        RECT 40.045 193.585 40.395 194.205 ;
        RECT 40.565 193.985 40.920 194.205 ;
        RECT 40.565 193.395 40.735 193.985 ;
        RECT 41.090 193.785 41.260 194.495 ;
        RECT 42.135 194.425 42.465 194.885 ;
        RECT 42.675 194.525 43.025 194.695 ;
        RECT 41.465 193.955 42.255 194.205 ;
        RECT 42.675 194.135 42.935 194.525 ;
        RECT 43.245 194.435 44.195 194.715 ;
        RECT 44.365 194.445 44.555 194.885 ;
        RECT 44.725 194.505 45.795 194.675 ;
        RECT 42.425 193.785 42.595 193.965 ;
        RECT 39.705 192.965 40.100 193.135 ;
        RECT 40.270 193.005 40.735 193.395 ;
        RECT 40.905 193.615 42.595 193.785 ;
        RECT 39.930 192.835 40.100 192.965 ;
        RECT 40.905 192.835 41.075 193.615 ;
        RECT 42.765 193.445 42.935 194.135 ;
        RECT 41.435 193.275 42.935 193.445 ;
        RECT 43.125 193.475 43.335 194.265 ;
        RECT 43.505 193.645 43.855 194.265 ;
        RECT 44.025 193.655 44.195 194.435 ;
        RECT 44.725 194.275 44.895 194.505 ;
        RECT 44.365 194.105 44.895 194.275 ;
        RECT 44.365 193.825 44.585 194.105 ;
        RECT 45.065 193.935 45.305 194.335 ;
        RECT 44.025 193.485 44.430 193.655 ;
        RECT 44.765 193.565 45.305 193.935 ;
        RECT 45.475 194.150 45.795 194.505 ;
        RECT 46.040 194.425 46.345 194.885 ;
        RECT 46.515 194.175 46.770 194.705 ;
        RECT 45.475 193.975 45.800 194.150 ;
        RECT 45.475 193.675 46.390 193.975 ;
        RECT 45.650 193.645 46.390 193.675 ;
        RECT 43.125 193.315 43.800 193.475 ;
        RECT 44.260 193.395 44.430 193.485 ;
        RECT 43.125 193.305 44.090 193.315 ;
        RECT 42.765 193.135 42.935 193.275 ;
        RECT 39.510 192.335 39.760 192.795 ;
        RECT 39.930 192.505 40.180 192.835 ;
        RECT 40.395 192.505 41.075 192.835 ;
        RECT 41.245 192.935 42.320 193.105 ;
        RECT 42.765 192.965 43.325 193.135 ;
        RECT 43.630 193.015 44.090 193.305 ;
        RECT 44.260 193.225 45.480 193.395 ;
        RECT 41.245 192.595 41.415 192.935 ;
        RECT 41.650 192.335 41.980 192.765 ;
        RECT 42.150 192.595 42.320 192.935 ;
        RECT 42.615 192.335 42.985 192.795 ;
        RECT 43.155 192.505 43.325 192.965 ;
        RECT 44.260 192.845 44.430 193.225 ;
        RECT 45.650 193.055 45.820 193.645 ;
        RECT 46.560 193.525 46.770 194.175 ;
        RECT 47.905 194.065 48.135 194.885 ;
        RECT 48.305 194.085 48.635 194.715 ;
        RECT 47.885 193.645 48.215 193.895 ;
        RECT 43.560 192.505 44.430 192.845 ;
        RECT 45.020 192.885 45.820 193.055 ;
        RECT 44.600 192.335 44.850 192.795 ;
        RECT 45.020 192.595 45.190 192.885 ;
        RECT 45.370 192.335 45.700 192.715 ;
        RECT 46.040 192.335 46.345 193.475 ;
        RECT 46.515 192.645 46.770 193.525 ;
        RECT 48.385 193.485 48.635 194.085 ;
        RECT 48.805 194.065 49.015 194.885 ;
        RECT 49.250 194.175 49.505 194.705 ;
        RECT 49.675 194.425 49.980 194.885 ;
        RECT 50.225 194.505 51.295 194.675 ;
        RECT 47.905 192.335 48.135 193.475 ;
        RECT 48.305 192.505 48.635 193.485 ;
        RECT 49.250 193.525 49.460 194.175 ;
        RECT 50.225 194.150 50.545 194.505 ;
        RECT 50.220 193.975 50.545 194.150 ;
        RECT 49.630 193.675 50.545 193.975 ;
        RECT 50.715 193.935 50.955 194.335 ;
        RECT 51.125 194.275 51.295 194.505 ;
        RECT 51.465 194.445 51.655 194.885 ;
        RECT 51.825 194.435 52.775 194.715 ;
        RECT 52.995 194.525 53.345 194.695 ;
        RECT 51.125 194.105 51.655 194.275 ;
        RECT 49.630 193.645 50.370 193.675 ;
        RECT 48.805 192.335 49.015 193.475 ;
        RECT 49.250 192.645 49.505 193.525 ;
        RECT 49.675 192.335 49.980 193.475 ;
        RECT 50.200 193.055 50.370 193.645 ;
        RECT 50.715 193.565 51.255 193.935 ;
        RECT 51.435 193.825 51.655 194.105 ;
        RECT 51.825 193.655 51.995 194.435 ;
        RECT 51.590 193.485 51.995 193.655 ;
        RECT 52.165 193.645 52.515 194.265 ;
        RECT 51.590 193.395 51.760 193.485 ;
        RECT 52.685 193.475 52.895 194.265 ;
        RECT 50.540 193.225 51.760 193.395 ;
        RECT 52.220 193.315 52.895 193.475 ;
        RECT 50.200 192.885 51.000 193.055 ;
        RECT 50.320 192.335 50.650 192.715 ;
        RECT 50.830 192.595 51.000 192.885 ;
        RECT 51.590 192.845 51.760 193.225 ;
        RECT 51.930 193.305 52.895 193.315 ;
        RECT 53.085 194.135 53.345 194.525 ;
        RECT 53.555 194.425 53.885 194.885 ;
        RECT 54.760 194.495 55.615 194.665 ;
        RECT 55.820 194.495 56.315 194.665 ;
        RECT 56.485 194.525 56.815 194.885 ;
        RECT 53.085 193.445 53.255 194.135 ;
        RECT 53.425 193.785 53.595 193.965 ;
        RECT 53.765 193.955 54.555 194.205 ;
        RECT 54.760 193.785 54.930 194.495 ;
        RECT 55.100 193.985 55.455 194.205 ;
        RECT 53.425 193.615 55.115 193.785 ;
        RECT 51.930 193.015 52.390 193.305 ;
        RECT 53.085 193.275 54.585 193.445 ;
        RECT 53.085 193.135 53.255 193.275 ;
        RECT 52.695 192.965 53.255 193.135 ;
        RECT 51.170 192.335 51.420 192.795 ;
        RECT 51.590 192.505 52.460 192.845 ;
        RECT 52.695 192.505 52.865 192.965 ;
        RECT 53.700 192.935 54.775 193.105 ;
        RECT 53.035 192.335 53.405 192.795 ;
        RECT 53.700 192.595 53.870 192.935 ;
        RECT 54.040 192.335 54.370 192.765 ;
        RECT 54.605 192.595 54.775 192.935 ;
        RECT 54.945 192.835 55.115 193.615 ;
        RECT 55.285 193.395 55.455 193.985 ;
        RECT 55.625 193.585 55.975 194.205 ;
        RECT 55.285 193.005 55.750 193.395 ;
        RECT 56.145 193.135 56.315 194.495 ;
        RECT 56.485 193.305 56.945 194.355 ;
        RECT 55.920 192.965 56.315 193.135 ;
        RECT 55.920 192.835 56.090 192.965 ;
        RECT 54.945 192.505 55.625 192.835 ;
        RECT 55.840 192.505 56.090 192.835 ;
        RECT 56.260 192.335 56.510 192.795 ;
        RECT 56.680 192.520 57.005 193.305 ;
        RECT 57.175 192.505 57.345 194.625 ;
        RECT 57.515 194.505 57.845 194.885 ;
        RECT 58.015 194.335 58.270 194.625 ;
        RECT 57.520 194.165 58.270 194.335 ;
        RECT 57.520 193.175 57.750 194.165 ;
        RECT 59.365 194.115 62.875 194.885 ;
        RECT 63.045 194.160 63.335 194.885 ;
        RECT 63.505 194.135 64.715 194.885 ;
        RECT 57.920 193.345 58.270 193.995 ;
        RECT 59.365 193.425 61.055 193.945 ;
        RECT 61.225 193.595 62.875 194.115 ;
        RECT 57.520 193.005 58.270 193.175 ;
        RECT 57.515 192.335 57.845 192.835 ;
        RECT 58.015 192.505 58.270 193.005 ;
        RECT 59.365 192.335 62.875 193.425 ;
        RECT 63.045 192.335 63.335 193.500 ;
        RECT 63.505 193.425 64.025 193.965 ;
        RECT 64.195 193.595 64.715 194.135 ;
        RECT 64.885 194.065 65.145 194.885 ;
        RECT 65.315 194.065 65.645 194.485 ;
        RECT 65.825 194.315 66.085 194.715 ;
        RECT 66.255 194.485 66.585 194.885 ;
        RECT 66.755 194.315 66.925 194.665 ;
        RECT 67.095 194.485 67.470 194.885 ;
        RECT 65.825 194.145 67.490 194.315 ;
        RECT 67.660 194.210 67.935 194.555 ;
        RECT 68.435 194.485 68.765 194.885 ;
        RECT 68.935 194.315 69.265 194.655 ;
        RECT 70.315 194.485 70.645 194.885 ;
        RECT 65.395 193.975 65.645 194.065 ;
        RECT 67.320 193.975 67.490 194.145 ;
        RECT 64.890 193.645 65.225 193.895 ;
        RECT 65.395 193.645 66.110 193.975 ;
        RECT 66.325 193.645 67.150 193.975 ;
        RECT 67.320 193.645 67.595 193.975 ;
        RECT 63.505 192.335 64.715 193.425 ;
        RECT 64.885 192.335 65.145 193.475 ;
        RECT 65.395 193.085 65.565 193.645 ;
        RECT 65.825 193.185 66.155 193.475 ;
        RECT 66.325 193.355 66.570 193.645 ;
        RECT 67.320 193.475 67.490 193.645 ;
        RECT 67.765 193.475 67.935 194.210 ;
        RECT 66.830 193.305 67.490 193.475 ;
        RECT 66.830 193.185 67.000 193.305 ;
        RECT 65.825 193.015 67.000 193.185 ;
        RECT 65.385 192.515 67.000 192.845 ;
        RECT 67.170 192.335 67.450 193.135 ;
        RECT 67.660 192.505 67.935 193.475 ;
        RECT 68.280 194.145 70.645 194.315 ;
        RECT 70.815 194.160 71.145 194.670 ;
        RECT 68.280 193.145 68.450 194.145 ;
        RECT 70.475 193.975 70.645 194.145 ;
        RECT 68.620 193.315 68.865 193.975 ;
        RECT 69.080 193.315 69.345 193.975 ;
        RECT 69.540 193.315 69.825 193.975 ;
        RECT 70.000 193.645 70.305 193.975 ;
        RECT 70.475 193.645 70.785 193.975 ;
        RECT 70.000 193.315 70.215 193.645 ;
        RECT 68.280 192.975 68.735 193.145 ;
        RECT 68.405 192.545 68.735 192.975 ;
        RECT 68.915 192.975 70.205 193.145 ;
        RECT 68.915 192.555 69.165 192.975 ;
        RECT 69.395 192.335 69.725 192.805 ;
        RECT 69.955 192.555 70.205 192.975 ;
        RECT 70.395 192.335 70.645 193.475 ;
        RECT 70.955 193.395 71.145 194.160 ;
        RECT 70.815 192.545 71.145 193.395 ;
        RECT 71.325 194.210 71.600 194.555 ;
        RECT 71.790 194.485 72.165 194.885 ;
        RECT 72.335 194.315 72.505 194.665 ;
        RECT 72.675 194.485 73.005 194.885 ;
        RECT 73.175 194.315 73.435 194.715 ;
        RECT 71.325 193.475 71.495 194.210 ;
        RECT 71.770 194.145 73.435 194.315 ;
        RECT 71.770 193.975 71.940 194.145 ;
        RECT 73.615 194.065 73.945 194.485 ;
        RECT 74.115 194.065 74.375 194.885 ;
        RECT 74.545 194.235 74.805 194.715 ;
        RECT 74.975 194.345 75.225 194.885 ;
        RECT 73.615 193.975 73.865 194.065 ;
        RECT 71.665 193.645 71.940 193.975 ;
        RECT 72.110 193.645 72.935 193.975 ;
        RECT 73.150 193.645 73.865 193.975 ;
        RECT 74.035 193.645 74.370 193.895 ;
        RECT 71.770 193.475 71.940 193.645 ;
        RECT 71.325 192.505 71.600 193.475 ;
        RECT 71.770 193.305 72.430 193.475 ;
        RECT 72.690 193.355 72.935 193.645 ;
        RECT 72.260 193.185 72.430 193.305 ;
        RECT 73.105 193.185 73.435 193.475 ;
        RECT 71.810 192.335 72.090 193.135 ;
        RECT 72.260 193.015 73.435 193.185 ;
        RECT 73.695 193.085 73.865 193.645 ;
        RECT 72.260 192.515 73.875 192.845 ;
        RECT 74.115 192.335 74.375 193.475 ;
        RECT 74.545 193.205 74.715 194.235 ;
        RECT 75.395 194.205 75.615 194.665 ;
        RECT 75.365 194.180 75.615 194.205 ;
        RECT 74.885 193.585 75.115 193.980 ;
        RECT 75.285 193.755 75.615 194.180 ;
        RECT 75.785 194.505 76.675 194.675 ;
        RECT 75.785 193.780 75.955 194.505 ;
        RECT 76.125 193.950 76.675 194.335 ;
        RECT 76.845 194.085 77.155 194.885 ;
        RECT 77.360 194.085 78.055 194.715 ;
        RECT 79.150 194.340 84.495 194.885 ;
        RECT 75.785 193.710 76.675 193.780 ;
        RECT 75.780 193.685 76.675 193.710 ;
        RECT 75.770 193.670 76.675 193.685 ;
        RECT 75.765 193.655 76.675 193.670 ;
        RECT 75.755 193.650 76.675 193.655 ;
        RECT 75.750 193.640 76.675 193.650 ;
        RECT 76.855 193.645 77.190 193.915 ;
        RECT 75.745 193.630 76.675 193.640 ;
        RECT 75.735 193.625 76.675 193.630 ;
        RECT 75.725 193.615 76.675 193.625 ;
        RECT 75.715 193.610 76.675 193.615 ;
        RECT 75.715 193.605 76.050 193.610 ;
        RECT 75.700 193.600 76.050 193.605 ;
        RECT 75.685 193.590 76.050 193.600 ;
        RECT 75.660 193.585 76.050 193.590 ;
        RECT 74.885 193.580 76.050 193.585 ;
        RECT 74.885 193.545 76.020 193.580 ;
        RECT 74.885 193.520 75.985 193.545 ;
        RECT 74.885 193.490 75.955 193.520 ;
        RECT 74.885 193.460 75.935 193.490 ;
        RECT 74.885 193.430 75.915 193.460 ;
        RECT 74.885 193.420 75.845 193.430 ;
        RECT 74.885 193.410 75.820 193.420 ;
        RECT 74.885 193.395 75.800 193.410 ;
        RECT 74.885 193.380 75.780 193.395 ;
        RECT 74.990 193.370 75.775 193.380 ;
        RECT 74.990 193.335 75.760 193.370 ;
        RECT 74.545 192.505 74.820 193.205 ;
        RECT 74.990 193.085 75.745 193.335 ;
        RECT 75.915 193.015 76.245 193.260 ;
        RECT 76.415 193.160 76.675 193.610 ;
        RECT 77.360 193.485 77.530 194.085 ;
        RECT 77.700 193.645 78.035 193.895 ;
        RECT 76.060 192.990 76.245 193.015 ;
        RECT 76.060 192.890 76.675 192.990 ;
        RECT 74.990 192.335 75.245 192.880 ;
        RECT 75.415 192.505 75.895 192.845 ;
        RECT 76.070 192.335 76.675 192.890 ;
        RECT 76.845 192.335 77.125 193.475 ;
        RECT 77.295 192.505 77.625 193.485 ;
        RECT 77.795 192.335 78.055 193.475 ;
        RECT 80.740 192.770 81.090 194.020 ;
        RECT 82.570 193.510 82.910 194.340 ;
        RECT 84.940 194.075 85.185 194.680 ;
        RECT 85.405 194.350 85.915 194.885 ;
        RECT 84.665 193.905 85.895 194.075 ;
        RECT 84.665 193.095 85.005 193.905 ;
        RECT 85.175 193.340 85.925 193.530 ;
        RECT 79.150 192.335 84.495 192.770 ;
        RECT 84.665 192.685 85.180 193.095 ;
        RECT 85.415 192.335 85.585 193.095 ;
        RECT 85.755 192.675 85.925 193.340 ;
        RECT 86.095 193.355 86.285 194.715 ;
        RECT 86.455 194.205 86.730 194.715 ;
        RECT 86.920 194.350 87.450 194.715 ;
        RECT 87.875 194.485 88.205 194.885 ;
        RECT 87.275 194.315 87.450 194.350 ;
        RECT 86.455 194.035 86.735 194.205 ;
        RECT 86.455 193.555 86.730 194.035 ;
        RECT 86.935 193.355 87.105 194.155 ;
        RECT 86.095 193.185 87.105 193.355 ;
        RECT 87.275 194.145 88.205 194.315 ;
        RECT 88.375 194.145 88.630 194.715 ;
        RECT 88.805 194.160 89.095 194.885 ;
        RECT 87.275 193.015 87.445 194.145 ;
        RECT 88.035 193.975 88.205 194.145 ;
        RECT 86.320 192.845 87.445 193.015 ;
        RECT 87.615 193.645 87.810 193.975 ;
        RECT 88.035 193.645 88.290 193.975 ;
        RECT 87.615 192.675 87.785 193.645 ;
        RECT 88.460 193.475 88.630 194.145 ;
        RECT 89.265 194.135 90.475 194.885 ;
        RECT 90.735 194.335 90.905 194.715 ;
        RECT 91.085 194.505 91.415 194.885 ;
        RECT 90.735 194.165 91.400 194.335 ;
        RECT 91.595 194.210 91.855 194.715 ;
        RECT 85.755 192.505 87.785 192.675 ;
        RECT 87.955 192.335 88.125 193.475 ;
        RECT 88.295 192.505 88.630 193.475 ;
        RECT 88.805 192.335 89.095 193.500 ;
        RECT 89.265 193.425 89.785 193.965 ;
        RECT 89.955 193.595 90.475 194.135 ;
        RECT 90.665 193.615 90.995 193.985 ;
        RECT 91.230 193.910 91.400 194.165 ;
        RECT 91.230 193.580 91.515 193.910 ;
        RECT 91.230 193.435 91.400 193.580 ;
        RECT 89.265 192.335 90.475 193.425 ;
        RECT 90.735 193.265 91.400 193.435 ;
        RECT 91.685 193.410 91.855 194.210 ;
        RECT 92.025 194.115 93.695 194.885 ;
        RECT 90.735 192.505 90.905 193.265 ;
        RECT 91.085 192.335 91.415 193.095 ;
        RECT 91.585 192.505 91.855 193.410 ;
        RECT 92.025 193.425 92.775 193.945 ;
        RECT 92.945 193.595 93.695 194.115 ;
        RECT 93.905 194.065 94.135 194.885 ;
        RECT 94.305 194.085 94.635 194.715 ;
        RECT 93.885 193.645 94.215 193.895 ;
        RECT 94.385 193.485 94.635 194.085 ;
        RECT 94.805 194.065 95.015 194.885 ;
        RECT 95.250 194.175 95.505 194.705 ;
        RECT 95.675 194.425 95.980 194.885 ;
        RECT 96.225 194.505 97.295 194.675 ;
        RECT 92.025 192.335 93.695 193.425 ;
        RECT 93.905 192.335 94.135 193.475 ;
        RECT 94.305 192.505 94.635 193.485 ;
        RECT 95.250 193.525 95.460 194.175 ;
        RECT 96.225 194.150 96.545 194.505 ;
        RECT 96.220 193.975 96.545 194.150 ;
        RECT 95.630 193.675 96.545 193.975 ;
        RECT 96.715 193.935 96.955 194.335 ;
        RECT 97.125 194.275 97.295 194.505 ;
        RECT 97.465 194.445 97.655 194.885 ;
        RECT 97.825 194.435 98.775 194.715 ;
        RECT 98.995 194.525 99.345 194.695 ;
        RECT 97.125 194.105 97.655 194.275 ;
        RECT 95.630 193.645 96.370 193.675 ;
        RECT 94.805 192.335 95.015 193.475 ;
        RECT 95.250 192.645 95.505 193.525 ;
        RECT 95.675 192.335 95.980 193.475 ;
        RECT 96.200 193.055 96.370 193.645 ;
        RECT 96.715 193.565 97.255 193.935 ;
        RECT 97.435 193.825 97.655 194.105 ;
        RECT 97.825 193.655 97.995 194.435 ;
        RECT 97.590 193.485 97.995 193.655 ;
        RECT 98.165 193.645 98.515 194.265 ;
        RECT 97.590 193.395 97.760 193.485 ;
        RECT 98.685 193.475 98.895 194.265 ;
        RECT 96.540 193.225 97.760 193.395 ;
        RECT 98.220 193.315 98.895 193.475 ;
        RECT 96.200 192.885 97.000 193.055 ;
        RECT 96.320 192.335 96.650 192.715 ;
        RECT 96.830 192.595 97.000 192.885 ;
        RECT 97.590 192.845 97.760 193.225 ;
        RECT 97.930 193.305 98.895 193.315 ;
        RECT 99.085 194.135 99.345 194.525 ;
        RECT 99.555 194.425 99.885 194.885 ;
        RECT 100.760 194.495 101.615 194.665 ;
        RECT 101.820 194.495 102.315 194.665 ;
        RECT 102.485 194.525 102.815 194.885 ;
        RECT 99.085 193.445 99.255 194.135 ;
        RECT 99.425 193.785 99.595 193.965 ;
        RECT 99.765 193.955 100.555 194.205 ;
        RECT 100.760 193.785 100.930 194.495 ;
        RECT 101.100 193.985 101.455 194.205 ;
        RECT 99.425 193.615 101.115 193.785 ;
        RECT 97.930 193.015 98.390 193.305 ;
        RECT 99.085 193.275 100.585 193.445 ;
        RECT 99.085 193.135 99.255 193.275 ;
        RECT 98.695 192.965 99.255 193.135 ;
        RECT 97.170 192.335 97.420 192.795 ;
        RECT 97.590 192.505 98.460 192.845 ;
        RECT 98.695 192.505 98.865 192.965 ;
        RECT 99.700 192.935 100.775 193.105 ;
        RECT 99.035 192.335 99.405 192.795 ;
        RECT 99.700 192.595 99.870 192.935 ;
        RECT 100.040 192.335 100.370 192.765 ;
        RECT 100.605 192.595 100.775 192.935 ;
        RECT 100.945 192.835 101.115 193.615 ;
        RECT 101.285 193.395 101.455 193.985 ;
        RECT 101.625 193.585 101.975 194.205 ;
        RECT 101.285 193.005 101.750 193.395 ;
        RECT 102.145 193.135 102.315 194.495 ;
        RECT 102.485 193.305 102.945 194.355 ;
        RECT 101.920 192.965 102.315 193.135 ;
        RECT 101.920 192.835 102.090 192.965 ;
        RECT 100.945 192.505 101.625 192.835 ;
        RECT 101.840 192.505 102.090 192.835 ;
        RECT 102.260 192.335 102.510 192.795 ;
        RECT 102.680 192.520 103.005 193.305 ;
        RECT 103.175 192.505 103.345 194.625 ;
        RECT 103.515 194.505 103.845 194.885 ;
        RECT 104.015 194.335 104.270 194.625 ;
        RECT 103.520 194.165 104.270 194.335 ;
        RECT 103.520 193.175 103.750 194.165 ;
        RECT 104.905 194.115 106.575 194.885 ;
        RECT 103.920 193.345 104.270 193.995 ;
        RECT 104.905 193.425 105.655 193.945 ;
        RECT 105.825 193.595 106.575 194.115 ;
        RECT 107.020 194.075 107.265 194.680 ;
        RECT 107.485 194.350 107.995 194.885 ;
        RECT 106.745 193.905 107.975 194.075 ;
        RECT 103.520 193.005 104.270 193.175 ;
        RECT 103.515 192.335 103.845 192.835 ;
        RECT 104.015 192.505 104.270 193.005 ;
        RECT 104.905 192.335 106.575 193.425 ;
        RECT 106.745 193.095 107.085 193.905 ;
        RECT 107.255 193.340 108.005 193.530 ;
        RECT 106.745 192.685 107.260 193.095 ;
        RECT 107.495 192.335 107.665 193.095 ;
        RECT 107.835 192.675 108.005 193.340 ;
        RECT 108.175 193.355 108.365 194.715 ;
        RECT 108.535 194.205 108.810 194.715 ;
        RECT 109.000 194.350 109.530 194.715 ;
        RECT 109.955 194.485 110.285 194.885 ;
        RECT 109.355 194.315 109.530 194.350 ;
        RECT 108.535 194.035 108.815 194.205 ;
        RECT 108.535 193.555 108.810 194.035 ;
        RECT 109.015 193.355 109.185 194.155 ;
        RECT 108.175 193.185 109.185 193.355 ;
        RECT 109.355 194.145 110.285 194.315 ;
        RECT 110.455 194.145 110.710 194.715 ;
        RECT 111.435 194.335 111.605 194.715 ;
        RECT 111.785 194.505 112.115 194.885 ;
        RECT 111.435 194.165 112.100 194.335 ;
        RECT 112.295 194.210 112.555 194.715 ;
        RECT 109.355 193.015 109.525 194.145 ;
        RECT 110.115 193.975 110.285 194.145 ;
        RECT 108.400 192.845 109.525 193.015 ;
        RECT 109.695 193.645 109.890 193.975 ;
        RECT 110.115 193.645 110.370 193.975 ;
        RECT 109.695 192.675 109.865 193.645 ;
        RECT 110.540 193.475 110.710 194.145 ;
        RECT 111.365 193.615 111.695 193.985 ;
        RECT 111.930 193.910 112.100 194.165 ;
        RECT 107.835 192.505 109.865 192.675 ;
        RECT 110.035 192.335 110.205 193.475 ;
        RECT 110.375 192.505 110.710 193.475 ;
        RECT 111.930 193.580 112.215 193.910 ;
        RECT 111.930 193.435 112.100 193.580 ;
        RECT 111.435 193.265 112.100 193.435 ;
        RECT 112.385 193.410 112.555 194.210 ;
        RECT 112.725 194.115 114.395 194.885 ;
        RECT 114.565 194.160 114.855 194.885 ;
        RECT 115.575 194.335 115.745 194.715 ;
        RECT 115.925 194.505 116.255 194.885 ;
        RECT 115.575 194.165 116.240 194.335 ;
        RECT 116.435 194.210 116.695 194.715 ;
        RECT 111.435 192.505 111.605 193.265 ;
        RECT 111.785 192.335 112.115 193.095 ;
        RECT 112.285 192.505 112.555 193.410 ;
        RECT 112.725 193.425 113.475 193.945 ;
        RECT 113.645 193.595 114.395 194.115 ;
        RECT 115.505 193.615 115.835 193.985 ;
        RECT 116.070 193.910 116.240 194.165 ;
        RECT 116.070 193.580 116.355 193.910 ;
        RECT 112.725 192.335 114.395 193.425 ;
        RECT 114.565 192.335 114.855 193.500 ;
        RECT 116.070 193.435 116.240 193.580 ;
        RECT 115.575 193.265 116.240 193.435 ;
        RECT 116.525 193.410 116.695 194.210 ;
        RECT 117.325 194.115 120.835 194.885 ;
        RECT 121.010 194.340 126.355 194.885 ;
        RECT 115.575 192.505 115.745 193.265 ;
        RECT 115.925 192.335 116.255 193.095 ;
        RECT 116.425 192.505 116.695 193.410 ;
        RECT 117.325 193.425 119.015 193.945 ;
        RECT 119.185 193.595 120.835 194.115 ;
        RECT 117.325 192.335 120.835 193.425 ;
        RECT 122.600 192.770 122.950 194.020 ;
        RECT 124.430 193.510 124.770 194.340 ;
        RECT 126.525 194.135 127.735 194.885 ;
        RECT 126.525 193.425 127.045 193.965 ;
        RECT 127.215 193.595 127.735 194.135 ;
        RECT 121.010 192.335 126.355 192.770 ;
        RECT 126.525 192.335 127.735 193.425 ;
        RECT 14.660 192.165 127.820 192.335 ;
        RECT 14.745 191.075 15.955 192.165 ;
        RECT 14.745 190.365 15.265 190.905 ;
        RECT 15.435 190.535 15.955 191.075 ;
        RECT 16.125 191.075 18.715 192.165 ;
        RECT 18.890 191.730 24.235 192.165 ;
        RECT 16.125 190.555 17.335 191.075 ;
        RECT 17.505 190.385 18.715 190.905 ;
        RECT 20.480 190.480 20.830 191.730 ;
        RECT 24.405 191.000 24.695 192.165 ;
        RECT 25.330 191.730 30.675 192.165 ;
        RECT 14.745 189.615 15.955 190.365 ;
        RECT 16.125 189.615 18.715 190.385 ;
        RECT 22.310 190.160 22.650 190.990 ;
        RECT 26.920 190.480 27.270 191.730 ;
        RECT 30.885 191.025 31.115 192.165 ;
        RECT 31.285 191.015 31.615 191.995 ;
        RECT 31.785 191.025 31.995 192.165 ;
        RECT 32.225 191.405 32.740 191.815 ;
        RECT 32.975 191.405 33.145 192.165 ;
        RECT 33.315 191.825 35.345 191.995 ;
        RECT 18.890 189.615 24.235 190.160 ;
        RECT 24.405 189.615 24.695 190.340 ;
        RECT 28.750 190.160 29.090 190.990 ;
        RECT 30.865 190.605 31.195 190.855 ;
        RECT 25.330 189.615 30.675 190.160 ;
        RECT 30.885 189.615 31.115 190.435 ;
        RECT 31.365 190.415 31.615 191.015 ;
        RECT 32.225 190.595 32.565 191.405 ;
        RECT 33.315 191.160 33.485 191.825 ;
        RECT 33.880 191.485 35.005 191.655 ;
        RECT 32.735 190.970 33.485 191.160 ;
        RECT 33.655 191.145 34.665 191.315 ;
        RECT 31.285 189.785 31.615 190.415 ;
        RECT 31.785 189.615 31.995 190.435 ;
        RECT 32.225 190.425 33.455 190.595 ;
        RECT 32.500 189.820 32.745 190.425 ;
        RECT 32.965 189.615 33.475 190.150 ;
        RECT 33.655 189.785 33.845 191.145 ;
        RECT 34.015 190.125 34.290 190.945 ;
        RECT 34.495 190.345 34.665 191.145 ;
        RECT 34.835 190.355 35.005 191.485 ;
        RECT 35.175 190.855 35.345 191.825 ;
        RECT 35.515 191.025 35.685 192.165 ;
        RECT 35.855 191.025 36.190 191.995 ;
        RECT 35.175 190.525 35.370 190.855 ;
        RECT 35.595 190.525 35.850 190.855 ;
        RECT 35.595 190.355 35.765 190.525 ;
        RECT 36.020 190.355 36.190 191.025 ;
        RECT 36.365 191.075 37.575 192.165 ;
        RECT 37.745 191.405 38.260 191.815 ;
        RECT 38.495 191.405 38.665 192.165 ;
        RECT 38.835 191.825 40.865 191.995 ;
        RECT 36.365 190.535 36.885 191.075 ;
        RECT 37.055 190.365 37.575 190.905 ;
        RECT 37.745 190.595 38.085 191.405 ;
        RECT 38.835 191.160 39.005 191.825 ;
        RECT 39.400 191.485 40.525 191.655 ;
        RECT 38.255 190.970 39.005 191.160 ;
        RECT 39.175 191.145 40.185 191.315 ;
        RECT 37.745 190.425 38.975 190.595 ;
        RECT 34.835 190.185 35.765 190.355 ;
        RECT 34.835 190.150 35.010 190.185 ;
        RECT 34.015 189.955 34.295 190.125 ;
        RECT 34.015 189.785 34.290 189.955 ;
        RECT 34.480 189.785 35.010 190.150 ;
        RECT 35.435 189.615 35.765 190.015 ;
        RECT 35.935 189.785 36.190 190.355 ;
        RECT 36.365 189.615 37.575 190.365 ;
        RECT 38.020 189.820 38.265 190.425 ;
        RECT 38.485 189.615 38.995 190.150 ;
        RECT 39.175 189.785 39.365 191.145 ;
        RECT 39.535 190.465 39.810 190.945 ;
        RECT 39.535 190.295 39.815 190.465 ;
        RECT 40.015 190.345 40.185 191.145 ;
        RECT 40.355 190.355 40.525 191.485 ;
        RECT 40.695 190.855 40.865 191.825 ;
        RECT 41.035 191.025 41.205 192.165 ;
        RECT 41.375 191.025 41.710 191.995 ;
        RECT 40.695 190.525 40.890 190.855 ;
        RECT 41.115 190.525 41.370 190.855 ;
        RECT 41.115 190.355 41.285 190.525 ;
        RECT 41.540 190.355 41.710 191.025 ;
        RECT 39.535 189.785 39.810 190.295 ;
        RECT 40.355 190.185 41.285 190.355 ;
        RECT 40.355 190.150 40.530 190.185 ;
        RECT 40.000 189.785 40.530 190.150 ;
        RECT 40.955 189.615 41.285 190.015 ;
        RECT 41.455 189.785 41.710 190.355 ;
        RECT 42.345 191.090 42.615 191.995 ;
        RECT 42.785 191.405 43.115 192.165 ;
        RECT 43.295 191.235 43.465 191.995 ;
        RECT 42.345 190.290 42.515 191.090 ;
        RECT 42.800 191.065 43.465 191.235 ;
        RECT 42.800 190.920 42.970 191.065 ;
        RECT 44.245 191.025 44.455 192.165 ;
        RECT 42.685 190.590 42.970 190.920 ;
        RECT 44.625 191.015 44.955 191.995 ;
        RECT 45.125 191.025 45.355 192.165 ;
        RECT 45.565 191.075 48.155 192.165 ;
        RECT 48.325 191.090 48.595 191.995 ;
        RECT 48.765 191.405 49.095 192.165 ;
        RECT 49.275 191.235 49.445 191.995 ;
        RECT 42.800 190.335 42.970 190.590 ;
        RECT 43.205 190.515 43.535 190.885 ;
        RECT 42.345 189.785 42.605 190.290 ;
        RECT 42.800 190.165 43.465 190.335 ;
        RECT 42.785 189.615 43.115 189.995 ;
        RECT 43.295 189.785 43.465 190.165 ;
        RECT 44.245 189.615 44.455 190.435 ;
        RECT 44.625 190.415 44.875 191.015 ;
        RECT 45.045 190.605 45.375 190.855 ;
        RECT 45.565 190.555 46.775 191.075 ;
        RECT 44.625 189.785 44.955 190.415 ;
        RECT 45.125 189.615 45.355 190.435 ;
        RECT 46.945 190.385 48.155 190.905 ;
        RECT 45.565 189.615 48.155 190.385 ;
        RECT 48.325 190.290 48.495 191.090 ;
        RECT 48.780 191.065 49.445 191.235 ;
        RECT 48.780 190.920 48.950 191.065 ;
        RECT 50.165 191.000 50.455 192.165 ;
        RECT 50.625 191.405 51.140 191.815 ;
        RECT 51.375 191.405 51.545 192.165 ;
        RECT 51.715 191.825 53.745 191.995 ;
        RECT 48.665 190.590 48.950 190.920 ;
        RECT 48.780 190.335 48.950 190.590 ;
        RECT 49.185 190.515 49.515 190.885 ;
        RECT 50.625 190.595 50.965 191.405 ;
        RECT 51.715 191.160 51.885 191.825 ;
        RECT 52.280 191.485 53.405 191.655 ;
        RECT 51.135 190.970 51.885 191.160 ;
        RECT 52.055 191.145 53.065 191.315 ;
        RECT 50.625 190.425 51.855 190.595 ;
        RECT 48.325 189.785 48.585 190.290 ;
        RECT 48.780 190.165 49.445 190.335 ;
        RECT 48.765 189.615 49.095 189.995 ;
        RECT 49.275 189.785 49.445 190.165 ;
        RECT 50.165 189.615 50.455 190.340 ;
        RECT 50.900 189.820 51.145 190.425 ;
        RECT 51.365 189.615 51.875 190.150 ;
        RECT 52.055 189.785 52.245 191.145 ;
        RECT 52.415 190.465 52.690 190.945 ;
        RECT 52.415 190.295 52.695 190.465 ;
        RECT 52.895 190.345 53.065 191.145 ;
        RECT 53.235 190.355 53.405 191.485 ;
        RECT 53.575 190.855 53.745 191.825 ;
        RECT 53.915 191.025 54.085 192.165 ;
        RECT 54.255 191.025 54.590 191.995 ;
        RECT 54.855 191.235 55.025 191.995 ;
        RECT 55.205 191.405 55.535 192.165 ;
        RECT 54.855 191.065 55.520 191.235 ;
        RECT 55.705 191.090 55.975 191.995 ;
        RECT 57.070 191.730 62.415 192.165 ;
        RECT 62.590 191.730 67.935 192.165 ;
        RECT 53.575 190.525 53.770 190.855 ;
        RECT 53.995 190.525 54.250 190.855 ;
        RECT 53.995 190.355 54.165 190.525 ;
        RECT 54.420 190.355 54.590 191.025 ;
        RECT 55.350 190.920 55.520 191.065 ;
        RECT 54.785 190.515 55.115 190.885 ;
        RECT 55.350 190.590 55.635 190.920 ;
        RECT 52.415 189.785 52.690 190.295 ;
        RECT 53.235 190.185 54.165 190.355 ;
        RECT 53.235 190.150 53.410 190.185 ;
        RECT 52.880 189.785 53.410 190.150 ;
        RECT 53.835 189.615 54.165 190.015 ;
        RECT 54.335 189.785 54.590 190.355 ;
        RECT 55.350 190.335 55.520 190.590 ;
        RECT 54.855 190.165 55.520 190.335 ;
        RECT 55.805 190.290 55.975 191.090 ;
        RECT 58.660 190.480 59.010 191.730 ;
        RECT 54.855 189.785 55.025 190.165 ;
        RECT 55.205 189.615 55.535 189.995 ;
        RECT 55.715 189.785 55.975 190.290 ;
        RECT 60.490 190.160 60.830 190.990 ;
        RECT 64.180 190.480 64.530 191.730 ;
        RECT 68.110 191.015 68.370 192.165 ;
        RECT 68.545 191.090 68.800 191.995 ;
        RECT 68.970 191.405 69.300 192.165 ;
        RECT 69.515 191.235 69.685 191.995 ;
        RECT 69.965 191.365 70.245 192.165 ;
        RECT 66.010 190.160 66.350 190.990 ;
        RECT 57.070 189.615 62.415 190.160 ;
        RECT 62.590 189.615 67.935 190.160 ;
        RECT 68.110 189.615 68.370 190.455 ;
        RECT 68.545 190.360 68.715 191.090 ;
        RECT 68.970 191.065 69.685 191.235 ;
        RECT 70.445 191.195 70.775 191.995 ;
        RECT 70.975 191.365 71.145 192.165 ;
        RECT 71.315 191.195 71.645 191.995 ;
        RECT 68.970 190.855 69.140 191.065 ;
        RECT 68.885 190.525 69.140 190.855 ;
        RECT 68.545 189.785 68.800 190.360 ;
        RECT 68.970 190.335 69.140 190.525 ;
        RECT 69.420 190.515 69.775 190.885 ;
        RECT 69.945 190.525 70.185 191.195 ;
        RECT 70.365 191.025 71.645 191.195 ;
        RECT 71.815 191.025 72.075 192.165 ;
        RECT 72.890 191.195 73.280 191.370 ;
        RECT 73.765 191.365 74.095 192.165 ;
        RECT 74.265 191.375 74.800 191.995 ;
        RECT 72.890 191.025 74.315 191.195 ;
        RECT 70.365 190.355 70.535 191.025 ;
        RECT 70.705 190.525 71.015 190.855 ;
        RECT 71.185 190.525 71.565 190.855 ;
        RECT 71.765 190.525 72.050 190.855 ;
        RECT 70.810 190.355 71.015 190.525 ;
        RECT 68.970 190.165 69.685 190.335 ;
        RECT 68.970 189.615 69.300 189.995 ;
        RECT 69.515 189.785 69.685 190.165 ;
        RECT 69.945 189.785 70.640 190.355 ;
        RECT 70.810 189.830 71.160 190.355 ;
        RECT 71.350 189.830 71.565 190.525 ;
        RECT 71.735 189.615 72.070 190.355 ;
        RECT 72.765 190.295 73.120 190.855 ;
        RECT 73.290 190.125 73.460 191.025 ;
        RECT 73.630 190.295 73.895 190.855 ;
        RECT 74.145 190.525 74.315 191.025 ;
        RECT 74.485 190.355 74.800 191.375 ;
        RECT 75.925 191.000 76.215 192.165 ;
        RECT 76.845 191.075 78.515 192.165 ;
        RECT 78.690 191.730 84.035 192.165 ;
        RECT 76.845 190.555 77.595 191.075 ;
        RECT 77.765 190.385 78.515 190.905 ;
        RECT 80.280 190.480 80.630 191.730 ;
        RECT 84.580 191.185 84.835 191.855 ;
        RECT 85.015 191.365 85.300 192.165 ;
        RECT 85.480 191.445 85.810 191.955 ;
        RECT 72.870 189.615 73.110 190.125 ;
        RECT 73.290 189.795 73.570 190.125 ;
        RECT 73.800 189.615 74.015 190.125 ;
        RECT 74.185 189.785 74.800 190.355 ;
        RECT 75.925 189.615 76.215 190.340 ;
        RECT 76.845 189.615 78.515 190.385 ;
        RECT 82.110 190.160 82.450 190.990 ;
        RECT 84.580 190.325 84.760 191.185 ;
        RECT 85.480 190.855 85.730 191.445 ;
        RECT 86.080 191.295 86.250 191.905 ;
        RECT 86.420 191.475 86.750 192.165 ;
        RECT 86.980 191.615 87.220 191.905 ;
        RECT 87.420 191.785 87.840 192.165 ;
        RECT 88.020 191.695 88.650 191.945 ;
        RECT 89.120 191.785 89.450 192.165 ;
        RECT 88.020 191.615 88.190 191.695 ;
        RECT 89.620 191.615 89.790 191.905 ;
        RECT 89.970 191.785 90.350 192.165 ;
        RECT 90.590 191.780 91.420 191.950 ;
        RECT 86.980 191.445 88.190 191.615 ;
        RECT 84.930 190.525 85.730 190.855 ;
        RECT 78.690 189.615 84.035 190.160 ;
        RECT 84.580 190.125 84.835 190.325 ;
        RECT 84.495 189.955 84.835 190.125 ;
        RECT 84.580 189.795 84.835 189.955 ;
        RECT 85.015 189.615 85.300 190.075 ;
        RECT 85.480 189.875 85.730 190.525 ;
        RECT 85.930 191.275 86.250 191.295 ;
        RECT 85.930 191.105 87.850 191.275 ;
        RECT 85.930 190.210 86.120 191.105 ;
        RECT 88.020 190.935 88.190 191.445 ;
        RECT 88.360 191.185 88.880 191.495 ;
        RECT 86.290 190.765 88.190 190.935 ;
        RECT 86.290 190.705 86.620 190.765 ;
        RECT 86.770 190.535 87.100 190.595 ;
        RECT 86.440 190.265 87.100 190.535 ;
        RECT 85.930 189.880 86.250 190.210 ;
        RECT 86.430 189.615 87.090 190.095 ;
        RECT 87.290 190.005 87.460 190.765 ;
        RECT 88.360 190.595 88.540 191.005 ;
        RECT 87.630 190.425 87.960 190.545 ;
        RECT 88.710 190.425 88.880 191.185 ;
        RECT 87.630 190.255 88.880 190.425 ;
        RECT 89.050 191.365 90.420 191.615 ;
        RECT 89.050 190.595 89.240 191.365 ;
        RECT 90.170 191.105 90.420 191.365 ;
        RECT 89.410 190.935 89.660 191.095 ;
        RECT 90.590 190.935 90.760 191.780 ;
        RECT 91.655 191.495 91.825 191.995 ;
        RECT 91.995 191.665 92.325 192.165 ;
        RECT 90.930 191.105 91.430 191.485 ;
        RECT 91.655 191.325 92.350 191.495 ;
        RECT 89.410 190.765 90.760 190.935 ;
        RECT 90.340 190.725 90.760 190.765 ;
        RECT 89.050 190.255 89.470 190.595 ;
        RECT 89.760 190.265 90.170 190.595 ;
        RECT 87.290 189.835 88.140 190.005 ;
        RECT 88.700 189.615 89.020 190.075 ;
        RECT 89.220 189.825 89.470 190.255 ;
        RECT 89.760 189.615 90.170 190.055 ;
        RECT 90.340 189.995 90.510 190.725 ;
        RECT 90.680 190.175 91.030 190.545 ;
        RECT 91.210 190.235 91.430 191.105 ;
        RECT 91.600 190.535 92.010 191.155 ;
        RECT 92.180 190.355 92.350 191.325 ;
        RECT 91.655 190.165 92.350 190.355 ;
        RECT 90.340 189.795 91.355 189.995 ;
        RECT 91.655 189.835 91.825 190.165 ;
        RECT 91.995 189.615 92.325 189.995 ;
        RECT 92.540 189.875 92.765 191.995 ;
        RECT 92.935 191.665 93.265 192.165 ;
        RECT 93.435 191.495 93.605 191.995 ;
        RECT 92.940 191.325 93.605 191.495 ;
        RECT 92.940 190.335 93.170 191.325 ;
        RECT 93.340 190.505 93.690 191.155 ;
        RECT 93.865 191.075 95.535 192.165 ;
        RECT 95.705 191.405 96.220 191.815 ;
        RECT 96.455 191.405 96.625 192.165 ;
        RECT 96.795 191.825 98.825 191.995 ;
        RECT 93.865 190.555 94.615 191.075 ;
        RECT 94.785 190.385 95.535 190.905 ;
        RECT 95.705 190.595 96.045 191.405 ;
        RECT 96.795 191.160 96.965 191.825 ;
        RECT 97.360 191.485 98.485 191.655 ;
        RECT 96.215 190.970 96.965 191.160 ;
        RECT 97.135 191.145 98.145 191.315 ;
        RECT 95.705 190.425 96.935 190.595 ;
        RECT 92.940 190.165 93.605 190.335 ;
        RECT 92.935 189.615 93.265 189.995 ;
        RECT 93.435 189.875 93.605 190.165 ;
        RECT 93.865 189.615 95.535 190.385 ;
        RECT 95.980 189.820 96.225 190.425 ;
        RECT 96.445 189.615 96.955 190.150 ;
        RECT 97.135 189.785 97.325 191.145 ;
        RECT 97.495 190.805 97.770 190.945 ;
        RECT 97.495 190.635 97.775 190.805 ;
        RECT 97.495 189.785 97.770 190.635 ;
        RECT 97.975 190.345 98.145 191.145 ;
        RECT 98.315 190.355 98.485 191.485 ;
        RECT 98.655 190.855 98.825 191.825 ;
        RECT 98.995 191.025 99.165 192.165 ;
        RECT 99.335 191.025 99.670 191.995 ;
        RECT 98.655 190.525 98.850 190.855 ;
        RECT 99.075 190.525 99.330 190.855 ;
        RECT 99.075 190.355 99.245 190.525 ;
        RECT 99.500 190.355 99.670 191.025 ;
        RECT 99.845 191.075 101.515 192.165 ;
        RECT 99.845 190.555 100.595 191.075 ;
        RECT 101.685 191.000 101.975 192.165 ;
        RECT 102.605 191.075 104.275 192.165 ;
        RECT 104.450 191.730 109.795 192.165 ;
        RECT 100.765 190.385 101.515 190.905 ;
        RECT 102.605 190.555 103.355 191.075 ;
        RECT 103.525 190.385 104.275 190.905 ;
        RECT 106.040 190.480 106.390 191.730 ;
        RECT 109.965 191.405 110.480 191.815 ;
        RECT 110.715 191.405 110.885 192.165 ;
        RECT 111.055 191.825 113.085 191.995 ;
        RECT 98.315 190.185 99.245 190.355 ;
        RECT 98.315 190.150 98.490 190.185 ;
        RECT 97.960 189.785 98.490 190.150 ;
        RECT 98.915 189.615 99.245 190.015 ;
        RECT 99.415 189.785 99.670 190.355 ;
        RECT 99.845 189.615 101.515 190.385 ;
        RECT 101.685 189.615 101.975 190.340 ;
        RECT 102.605 189.615 104.275 190.385 ;
        RECT 107.870 190.160 108.210 190.990 ;
        RECT 109.965 190.595 110.305 191.405 ;
        RECT 111.055 191.160 111.225 191.825 ;
        RECT 111.620 191.485 112.745 191.655 ;
        RECT 110.475 190.970 111.225 191.160 ;
        RECT 111.395 191.145 112.405 191.315 ;
        RECT 109.965 190.425 111.195 190.595 ;
        RECT 104.450 189.615 109.795 190.160 ;
        RECT 110.240 189.820 110.485 190.425 ;
        RECT 110.705 189.615 111.215 190.150 ;
        RECT 111.395 189.785 111.585 191.145 ;
        RECT 111.755 190.125 112.030 190.945 ;
        RECT 112.235 190.345 112.405 191.145 ;
        RECT 112.575 190.355 112.745 191.485 ;
        RECT 112.915 190.855 113.085 191.825 ;
        RECT 113.255 191.025 113.425 192.165 ;
        RECT 113.595 191.025 113.930 191.995 ;
        RECT 112.915 190.525 113.110 190.855 ;
        RECT 113.335 190.525 113.590 190.855 ;
        RECT 113.335 190.355 113.505 190.525 ;
        RECT 113.760 190.355 113.930 191.025 ;
        RECT 114.105 191.075 115.315 192.165 ;
        RECT 115.490 191.730 120.835 192.165 ;
        RECT 121.010 191.730 126.355 192.165 ;
        RECT 114.105 190.535 114.625 191.075 ;
        RECT 114.795 190.365 115.315 190.905 ;
        RECT 117.080 190.480 117.430 191.730 ;
        RECT 112.575 190.185 113.505 190.355 ;
        RECT 112.575 190.150 112.750 190.185 ;
        RECT 111.755 189.955 112.035 190.125 ;
        RECT 111.755 189.785 112.030 189.955 ;
        RECT 112.220 189.785 112.750 190.150 ;
        RECT 113.175 189.615 113.505 190.015 ;
        RECT 113.675 189.785 113.930 190.355 ;
        RECT 114.105 189.615 115.315 190.365 ;
        RECT 118.910 190.160 119.250 190.990 ;
        RECT 122.600 190.480 122.950 191.730 ;
        RECT 126.525 191.075 127.735 192.165 ;
        RECT 124.430 190.160 124.770 190.990 ;
        RECT 126.525 190.535 127.045 191.075 ;
        RECT 127.215 190.365 127.735 190.905 ;
        RECT 115.490 189.615 120.835 190.160 ;
        RECT 121.010 189.615 126.355 190.160 ;
        RECT 126.525 189.615 127.735 190.365 ;
        RECT 14.660 189.445 127.820 189.615 ;
        RECT 14.745 188.695 15.955 189.445 ;
        RECT 14.745 188.155 15.265 188.695 ;
        RECT 17.045 188.675 20.555 189.445 ;
        RECT 20.730 188.900 26.075 189.445 ;
        RECT 15.435 187.985 15.955 188.525 ;
        RECT 14.745 186.895 15.955 187.985 ;
        RECT 17.045 187.985 18.735 188.505 ;
        RECT 18.905 188.155 20.555 188.675 ;
        RECT 17.045 186.895 20.555 187.985 ;
        RECT 22.320 187.330 22.670 188.580 ;
        RECT 24.150 188.070 24.490 188.900 ;
        RECT 26.285 188.625 26.515 189.445 ;
        RECT 26.685 188.645 27.015 189.275 ;
        RECT 26.265 188.205 26.595 188.455 ;
        RECT 26.765 188.045 27.015 188.645 ;
        RECT 27.185 188.625 27.395 189.445 ;
        RECT 28.000 189.105 28.255 189.265 ;
        RECT 27.915 188.935 28.255 189.105 ;
        RECT 28.435 188.985 28.720 189.445 ;
        RECT 28.000 188.735 28.255 188.935 ;
        RECT 20.730 186.895 26.075 187.330 ;
        RECT 26.285 186.895 26.515 188.035 ;
        RECT 26.685 187.065 27.015 188.045 ;
        RECT 27.185 186.895 27.395 188.035 ;
        RECT 28.000 187.875 28.180 188.735 ;
        RECT 28.900 188.535 29.150 189.185 ;
        RECT 28.350 188.205 29.150 188.535 ;
        RECT 28.000 187.205 28.255 187.875 ;
        RECT 28.435 186.895 28.720 187.695 ;
        RECT 28.900 187.615 29.150 188.205 ;
        RECT 29.350 188.850 29.670 189.180 ;
        RECT 29.850 188.965 30.510 189.445 ;
        RECT 30.710 189.055 31.560 189.225 ;
        RECT 29.350 187.955 29.540 188.850 ;
        RECT 29.860 188.525 30.520 188.795 ;
        RECT 30.190 188.465 30.520 188.525 ;
        RECT 29.710 188.295 30.040 188.355 ;
        RECT 30.710 188.295 30.880 189.055 ;
        RECT 32.120 188.985 32.440 189.445 ;
        RECT 32.640 188.805 32.890 189.235 ;
        RECT 33.180 189.005 33.590 189.445 ;
        RECT 33.760 189.065 34.775 189.265 ;
        RECT 31.050 188.635 32.300 188.805 ;
        RECT 31.050 188.515 31.380 188.635 ;
        RECT 29.710 188.125 31.610 188.295 ;
        RECT 29.350 187.785 31.270 187.955 ;
        RECT 29.350 187.765 29.670 187.785 ;
        RECT 28.900 187.105 29.230 187.615 ;
        RECT 29.500 187.155 29.670 187.765 ;
        RECT 31.440 187.615 31.610 188.125 ;
        RECT 31.780 188.055 31.960 188.465 ;
        RECT 32.130 187.875 32.300 188.635 ;
        RECT 29.840 186.895 30.170 187.585 ;
        RECT 30.400 187.445 31.610 187.615 ;
        RECT 31.780 187.565 32.300 187.875 ;
        RECT 32.470 188.465 32.890 188.805 ;
        RECT 33.180 188.465 33.590 188.795 ;
        RECT 32.470 187.695 32.660 188.465 ;
        RECT 33.760 188.335 33.930 189.065 ;
        RECT 35.075 188.895 35.245 189.225 ;
        RECT 35.415 189.065 35.745 189.445 ;
        RECT 34.100 188.515 34.450 188.885 ;
        RECT 33.760 188.295 34.180 188.335 ;
        RECT 32.830 188.125 34.180 188.295 ;
        RECT 32.830 187.965 33.080 188.125 ;
        RECT 33.590 187.695 33.840 187.955 ;
        RECT 32.470 187.445 33.840 187.695 ;
        RECT 30.400 187.155 30.640 187.445 ;
        RECT 31.440 187.365 31.610 187.445 ;
        RECT 30.840 186.895 31.260 187.275 ;
        RECT 31.440 187.115 32.070 187.365 ;
        RECT 32.540 186.895 32.870 187.275 ;
        RECT 33.040 187.155 33.210 187.445 ;
        RECT 34.010 187.280 34.180 188.125 ;
        RECT 34.630 187.955 34.850 188.825 ;
        RECT 35.075 188.705 35.770 188.895 ;
        RECT 34.350 187.575 34.850 187.955 ;
        RECT 35.020 187.905 35.430 188.525 ;
        RECT 35.600 187.735 35.770 188.705 ;
        RECT 35.075 187.565 35.770 187.735 ;
        RECT 33.390 186.895 33.770 187.275 ;
        RECT 34.010 187.110 34.840 187.280 ;
        RECT 35.075 187.065 35.245 187.565 ;
        RECT 35.415 186.895 35.745 187.395 ;
        RECT 35.960 187.065 36.185 189.185 ;
        RECT 36.355 189.065 36.685 189.445 ;
        RECT 36.855 188.895 37.025 189.185 ;
        RECT 36.360 188.725 37.025 188.895 ;
        RECT 36.360 187.735 36.590 188.725 ;
        RECT 37.285 188.720 37.575 189.445 ;
        RECT 37.745 188.770 38.005 189.275 ;
        RECT 38.185 189.065 38.515 189.445 ;
        RECT 38.695 188.895 38.865 189.275 ;
        RECT 36.760 187.905 37.110 188.555 ;
        RECT 36.360 187.565 37.025 187.735 ;
        RECT 36.355 186.895 36.685 187.395 ;
        RECT 36.855 187.065 37.025 187.565 ;
        RECT 37.285 186.895 37.575 188.060 ;
        RECT 37.745 187.970 37.915 188.770 ;
        RECT 38.200 188.725 38.865 188.895 ;
        RECT 40.050 188.735 40.305 189.265 ;
        RECT 40.475 188.985 40.780 189.445 ;
        RECT 41.025 189.065 42.095 189.235 ;
        RECT 38.200 188.470 38.370 188.725 ;
        RECT 38.085 188.140 38.370 188.470 ;
        RECT 38.605 188.175 38.935 188.545 ;
        RECT 38.200 187.995 38.370 188.140 ;
        RECT 40.050 188.085 40.260 188.735 ;
        RECT 41.025 188.710 41.345 189.065 ;
        RECT 41.020 188.535 41.345 188.710 ;
        RECT 40.430 188.235 41.345 188.535 ;
        RECT 41.515 188.495 41.755 188.895 ;
        RECT 41.925 188.835 42.095 189.065 ;
        RECT 42.265 189.005 42.455 189.445 ;
        RECT 42.625 188.995 43.575 189.275 ;
        RECT 43.795 189.085 44.145 189.255 ;
        RECT 41.925 188.665 42.455 188.835 ;
        RECT 40.430 188.205 41.170 188.235 ;
        RECT 37.745 187.065 38.015 187.970 ;
        RECT 38.200 187.825 38.865 187.995 ;
        RECT 38.185 186.895 38.515 187.655 ;
        RECT 38.695 187.065 38.865 187.825 ;
        RECT 40.050 187.205 40.305 188.085 ;
        RECT 40.475 186.895 40.780 188.035 ;
        RECT 41.000 187.615 41.170 188.205 ;
        RECT 41.515 188.125 42.055 188.495 ;
        RECT 42.235 188.385 42.455 188.665 ;
        RECT 42.625 188.215 42.795 188.995 ;
        RECT 42.390 188.045 42.795 188.215 ;
        RECT 42.965 188.205 43.315 188.825 ;
        RECT 42.390 187.955 42.560 188.045 ;
        RECT 43.485 188.035 43.695 188.825 ;
        RECT 41.340 187.785 42.560 187.955 ;
        RECT 43.020 187.875 43.695 188.035 ;
        RECT 41.000 187.445 41.800 187.615 ;
        RECT 41.120 186.895 41.450 187.275 ;
        RECT 41.630 187.155 41.800 187.445 ;
        RECT 42.390 187.405 42.560 187.785 ;
        RECT 42.730 187.865 43.695 187.875 ;
        RECT 43.885 188.695 44.145 189.085 ;
        RECT 44.355 188.985 44.685 189.445 ;
        RECT 45.560 189.055 46.415 189.225 ;
        RECT 46.620 189.055 47.115 189.225 ;
        RECT 47.285 189.085 47.615 189.445 ;
        RECT 43.885 188.005 44.055 188.695 ;
        RECT 44.225 188.345 44.395 188.525 ;
        RECT 44.565 188.515 45.355 188.765 ;
        RECT 45.560 188.345 45.730 189.055 ;
        RECT 45.900 188.545 46.255 188.765 ;
        RECT 44.225 188.175 45.915 188.345 ;
        RECT 42.730 187.575 43.190 187.865 ;
        RECT 43.885 187.835 45.385 188.005 ;
        RECT 43.885 187.695 44.055 187.835 ;
        RECT 43.495 187.525 44.055 187.695 ;
        RECT 41.970 186.895 42.220 187.355 ;
        RECT 42.390 187.065 43.260 187.405 ;
        RECT 43.495 187.065 43.665 187.525 ;
        RECT 44.500 187.495 45.575 187.665 ;
        RECT 43.835 186.895 44.205 187.355 ;
        RECT 44.500 187.155 44.670 187.495 ;
        RECT 44.840 186.895 45.170 187.325 ;
        RECT 45.405 187.155 45.575 187.495 ;
        RECT 45.745 187.395 45.915 188.175 ;
        RECT 46.085 187.955 46.255 188.545 ;
        RECT 46.425 188.145 46.775 188.765 ;
        RECT 46.085 187.565 46.550 187.955 ;
        RECT 46.945 187.695 47.115 189.055 ;
        RECT 47.285 187.865 47.745 188.915 ;
        RECT 46.720 187.525 47.115 187.695 ;
        RECT 46.720 187.395 46.890 187.525 ;
        RECT 45.745 187.065 46.425 187.395 ;
        RECT 46.640 187.065 46.890 187.395 ;
        RECT 47.060 186.895 47.310 187.355 ;
        RECT 47.480 187.080 47.805 187.865 ;
        RECT 47.975 187.065 48.145 189.185 ;
        RECT 48.315 189.065 48.645 189.445 ;
        RECT 48.815 188.895 49.070 189.185 ;
        RECT 48.320 188.725 49.070 188.895 ;
        RECT 49.250 188.735 49.505 189.265 ;
        RECT 49.675 188.985 49.980 189.445 ;
        RECT 50.225 189.065 51.295 189.235 ;
        RECT 48.320 187.735 48.550 188.725 ;
        RECT 48.720 187.905 49.070 188.555 ;
        RECT 49.250 188.085 49.460 188.735 ;
        RECT 50.225 188.710 50.545 189.065 ;
        RECT 50.220 188.535 50.545 188.710 ;
        RECT 49.630 188.235 50.545 188.535 ;
        RECT 50.715 188.495 50.955 188.895 ;
        RECT 51.125 188.835 51.295 189.065 ;
        RECT 51.465 189.005 51.655 189.445 ;
        RECT 51.825 188.995 52.775 189.275 ;
        RECT 52.995 189.085 53.345 189.255 ;
        RECT 51.125 188.665 51.655 188.835 ;
        RECT 49.630 188.205 50.370 188.235 ;
        RECT 48.320 187.565 49.070 187.735 ;
        RECT 48.315 186.895 48.645 187.395 ;
        RECT 48.815 187.065 49.070 187.565 ;
        RECT 49.250 187.205 49.505 188.085 ;
        RECT 49.675 186.895 49.980 188.035 ;
        RECT 50.200 187.615 50.370 188.205 ;
        RECT 50.715 188.125 51.255 188.495 ;
        RECT 51.435 188.385 51.655 188.665 ;
        RECT 51.825 188.215 51.995 188.995 ;
        RECT 51.590 188.045 51.995 188.215 ;
        RECT 52.165 188.205 52.515 188.825 ;
        RECT 51.590 187.955 51.760 188.045 ;
        RECT 52.685 188.035 52.895 188.825 ;
        RECT 50.540 187.785 51.760 187.955 ;
        RECT 52.220 187.875 52.895 188.035 ;
        RECT 50.200 187.445 51.000 187.615 ;
        RECT 50.320 186.895 50.650 187.275 ;
        RECT 50.830 187.155 51.000 187.445 ;
        RECT 51.590 187.405 51.760 187.785 ;
        RECT 51.930 187.865 52.895 187.875 ;
        RECT 53.085 188.695 53.345 189.085 ;
        RECT 53.555 188.985 53.885 189.445 ;
        RECT 54.760 189.055 55.615 189.225 ;
        RECT 55.820 189.055 56.315 189.225 ;
        RECT 56.485 189.085 56.815 189.445 ;
        RECT 53.085 188.005 53.255 188.695 ;
        RECT 53.425 188.345 53.595 188.525 ;
        RECT 53.765 188.515 54.555 188.765 ;
        RECT 54.760 188.345 54.930 189.055 ;
        RECT 55.100 188.545 55.455 188.765 ;
        RECT 53.425 188.175 55.115 188.345 ;
        RECT 51.930 187.575 52.390 187.865 ;
        RECT 53.085 187.835 54.585 188.005 ;
        RECT 53.085 187.695 53.255 187.835 ;
        RECT 52.695 187.525 53.255 187.695 ;
        RECT 51.170 186.895 51.420 187.355 ;
        RECT 51.590 187.065 52.460 187.405 ;
        RECT 52.695 187.065 52.865 187.525 ;
        RECT 53.700 187.495 54.775 187.665 ;
        RECT 53.035 186.895 53.405 187.355 ;
        RECT 53.700 187.155 53.870 187.495 ;
        RECT 54.040 186.895 54.370 187.325 ;
        RECT 54.605 187.155 54.775 187.495 ;
        RECT 54.945 187.395 55.115 188.175 ;
        RECT 55.285 187.955 55.455 188.545 ;
        RECT 55.625 188.145 55.975 188.765 ;
        RECT 55.285 187.565 55.750 187.955 ;
        RECT 56.145 187.695 56.315 189.055 ;
        RECT 56.485 187.865 56.945 188.915 ;
        RECT 55.920 187.525 56.315 187.695 ;
        RECT 55.920 187.395 56.090 187.525 ;
        RECT 54.945 187.065 55.625 187.395 ;
        RECT 55.840 187.065 56.090 187.395 ;
        RECT 56.260 186.895 56.510 187.355 ;
        RECT 56.680 187.080 57.005 187.865 ;
        RECT 57.175 187.065 57.345 189.185 ;
        RECT 57.515 189.065 57.845 189.445 ;
        RECT 58.015 188.895 58.270 189.185 ;
        RECT 57.520 188.725 58.270 188.895 ;
        RECT 57.520 187.735 57.750 188.725 ;
        RECT 59.365 188.675 62.875 189.445 ;
        RECT 63.045 188.720 63.335 189.445 ;
        RECT 63.505 188.675 67.015 189.445 ;
        RECT 67.190 188.900 72.535 189.445 ;
        RECT 57.920 187.905 58.270 188.555 ;
        RECT 59.365 187.985 61.055 188.505 ;
        RECT 61.225 188.155 62.875 188.675 ;
        RECT 57.520 187.565 58.270 187.735 ;
        RECT 57.515 186.895 57.845 187.395 ;
        RECT 58.015 187.065 58.270 187.565 ;
        RECT 59.365 186.895 62.875 187.985 ;
        RECT 63.045 186.895 63.335 188.060 ;
        RECT 63.505 187.985 65.195 188.505 ;
        RECT 65.365 188.155 67.015 188.675 ;
        RECT 63.505 186.895 67.015 187.985 ;
        RECT 68.780 187.330 69.130 188.580 ;
        RECT 70.610 188.070 70.950 188.900 ;
        RECT 72.765 188.625 72.975 189.445 ;
        RECT 73.145 188.645 73.475 189.275 ;
        RECT 73.145 188.045 73.395 188.645 ;
        RECT 73.645 188.625 73.875 189.445 ;
        RECT 74.085 188.675 75.755 189.445 ;
        RECT 73.565 188.205 73.895 188.455 ;
        RECT 67.190 186.895 72.535 187.330 ;
        RECT 72.765 186.895 72.975 188.035 ;
        RECT 73.145 187.065 73.475 188.045 ;
        RECT 73.645 186.895 73.875 188.035 ;
        RECT 74.085 187.985 74.835 188.505 ;
        RECT 75.005 188.155 75.755 188.675 ;
        RECT 75.925 188.770 76.185 189.275 ;
        RECT 76.365 189.065 76.695 189.445 ;
        RECT 76.875 188.895 77.045 189.275 ;
        RECT 74.085 186.895 75.755 187.985 ;
        RECT 75.925 187.970 76.095 188.770 ;
        RECT 76.380 188.725 77.045 188.895 ;
        RECT 76.380 188.470 76.550 188.725 ;
        RECT 77.765 188.675 80.355 189.445 ;
        RECT 80.530 188.900 85.875 189.445 ;
        RECT 76.265 188.140 76.550 188.470 ;
        RECT 76.785 188.175 77.115 188.545 ;
        RECT 76.380 187.995 76.550 188.140 ;
        RECT 75.925 187.065 76.195 187.970 ;
        RECT 76.380 187.825 77.045 187.995 ;
        RECT 76.365 186.895 76.695 187.655 ;
        RECT 76.875 187.065 77.045 187.825 ;
        RECT 77.765 187.985 78.975 188.505 ;
        RECT 79.145 188.155 80.355 188.675 ;
        RECT 77.765 186.895 80.355 187.985 ;
        RECT 82.120 187.330 82.470 188.580 ;
        RECT 83.950 188.070 84.290 188.900 ;
        RECT 86.085 188.625 86.315 189.445 ;
        RECT 86.485 188.645 86.815 189.275 ;
        RECT 86.065 188.205 86.395 188.455 ;
        RECT 86.565 188.045 86.815 188.645 ;
        RECT 86.985 188.625 87.195 189.445 ;
        RECT 87.465 188.625 87.695 189.445 ;
        RECT 87.865 188.645 88.195 189.275 ;
        RECT 87.445 188.205 87.775 188.455 ;
        RECT 87.945 188.045 88.195 188.645 ;
        RECT 88.365 188.625 88.575 189.445 ;
        RECT 88.805 188.720 89.095 189.445 ;
        RECT 89.815 188.895 89.985 189.275 ;
        RECT 90.165 189.065 90.495 189.445 ;
        RECT 89.815 188.725 90.480 188.895 ;
        RECT 90.675 188.770 90.935 189.275 ;
        RECT 91.570 188.900 96.915 189.445 ;
        RECT 89.745 188.175 90.075 188.545 ;
        RECT 90.310 188.470 90.480 188.725 ;
        RECT 90.310 188.140 90.595 188.470 ;
        RECT 80.530 186.895 85.875 187.330 ;
        RECT 86.085 186.895 86.315 188.035 ;
        RECT 86.485 187.065 86.815 188.045 ;
        RECT 86.985 186.895 87.195 188.035 ;
        RECT 87.465 186.895 87.695 188.035 ;
        RECT 87.865 187.065 88.195 188.045 ;
        RECT 88.365 186.895 88.575 188.035 ;
        RECT 88.805 186.895 89.095 188.060 ;
        RECT 90.310 187.995 90.480 188.140 ;
        RECT 89.815 187.825 90.480 187.995 ;
        RECT 90.765 187.970 90.935 188.770 ;
        RECT 89.815 187.065 89.985 187.825 ;
        RECT 90.165 186.895 90.495 187.655 ;
        RECT 90.665 187.065 90.935 187.970 ;
        RECT 93.160 187.330 93.510 188.580 ;
        RECT 94.990 188.070 95.330 188.900 ;
        RECT 97.125 188.625 97.355 189.445 ;
        RECT 97.525 188.645 97.855 189.275 ;
        RECT 97.105 188.205 97.435 188.455 ;
        RECT 97.605 188.045 97.855 188.645 ;
        RECT 98.025 188.625 98.235 189.445 ;
        RECT 98.470 188.735 98.725 189.265 ;
        RECT 98.895 188.985 99.200 189.445 ;
        RECT 99.445 189.065 100.515 189.235 ;
        RECT 91.570 186.895 96.915 187.330 ;
        RECT 97.125 186.895 97.355 188.035 ;
        RECT 97.525 187.065 97.855 188.045 ;
        RECT 98.470 188.085 98.680 188.735 ;
        RECT 99.445 188.710 99.765 189.065 ;
        RECT 99.440 188.535 99.765 188.710 ;
        RECT 98.850 188.235 99.765 188.535 ;
        RECT 99.935 188.495 100.175 188.895 ;
        RECT 100.345 188.835 100.515 189.065 ;
        RECT 100.685 189.005 100.875 189.445 ;
        RECT 101.045 188.995 101.995 189.275 ;
        RECT 102.215 189.085 102.565 189.255 ;
        RECT 100.345 188.665 100.875 188.835 ;
        RECT 98.850 188.205 99.590 188.235 ;
        RECT 98.025 186.895 98.235 188.035 ;
        RECT 98.470 187.205 98.725 188.085 ;
        RECT 98.895 186.895 99.200 188.035 ;
        RECT 99.420 187.615 99.590 188.205 ;
        RECT 99.935 188.125 100.475 188.495 ;
        RECT 100.655 188.385 100.875 188.665 ;
        RECT 101.045 188.215 101.215 188.995 ;
        RECT 100.810 188.045 101.215 188.215 ;
        RECT 101.385 188.205 101.735 188.825 ;
        RECT 100.810 187.955 100.980 188.045 ;
        RECT 101.905 188.035 102.115 188.825 ;
        RECT 99.760 187.785 100.980 187.955 ;
        RECT 101.440 187.875 102.115 188.035 ;
        RECT 99.420 187.445 100.220 187.615 ;
        RECT 99.540 186.895 99.870 187.275 ;
        RECT 100.050 187.155 100.220 187.445 ;
        RECT 100.810 187.405 100.980 187.785 ;
        RECT 101.150 187.865 102.115 187.875 ;
        RECT 102.305 188.695 102.565 189.085 ;
        RECT 102.775 188.985 103.105 189.445 ;
        RECT 103.980 189.055 104.835 189.225 ;
        RECT 105.040 189.055 105.535 189.225 ;
        RECT 105.705 189.085 106.035 189.445 ;
        RECT 102.305 188.005 102.475 188.695 ;
        RECT 102.645 188.345 102.815 188.525 ;
        RECT 102.985 188.515 103.775 188.765 ;
        RECT 103.980 188.345 104.150 189.055 ;
        RECT 104.320 188.545 104.675 188.765 ;
        RECT 102.645 188.175 104.335 188.345 ;
        RECT 101.150 187.575 101.610 187.865 ;
        RECT 102.305 187.835 103.805 188.005 ;
        RECT 102.305 187.695 102.475 187.835 ;
        RECT 101.915 187.525 102.475 187.695 ;
        RECT 100.390 186.895 100.640 187.355 ;
        RECT 100.810 187.065 101.680 187.405 ;
        RECT 101.915 187.065 102.085 187.525 ;
        RECT 102.920 187.495 103.995 187.665 ;
        RECT 102.255 186.895 102.625 187.355 ;
        RECT 102.920 187.155 103.090 187.495 ;
        RECT 103.260 186.895 103.590 187.325 ;
        RECT 103.825 187.155 103.995 187.495 ;
        RECT 104.165 187.395 104.335 188.175 ;
        RECT 104.505 187.955 104.675 188.545 ;
        RECT 104.845 188.145 105.195 188.765 ;
        RECT 104.505 187.565 104.970 187.955 ;
        RECT 105.365 187.695 105.535 189.055 ;
        RECT 105.705 187.865 106.165 188.915 ;
        RECT 105.140 187.525 105.535 187.695 ;
        RECT 105.140 187.395 105.310 187.525 ;
        RECT 104.165 187.065 104.845 187.395 ;
        RECT 105.060 187.065 105.310 187.395 ;
        RECT 105.480 186.895 105.730 187.355 ;
        RECT 105.900 187.080 106.225 187.865 ;
        RECT 106.395 187.065 106.565 189.185 ;
        RECT 106.735 189.065 107.065 189.445 ;
        RECT 107.235 188.895 107.490 189.185 ;
        RECT 106.740 188.725 107.490 188.895 ;
        RECT 106.740 187.735 106.970 188.725 ;
        RECT 107.665 188.695 108.875 189.445 ;
        RECT 109.050 188.900 114.395 189.445 ;
        RECT 107.140 187.905 107.490 188.555 ;
        RECT 107.665 187.985 108.185 188.525 ;
        RECT 108.355 188.155 108.875 188.695 ;
        RECT 106.740 187.565 107.490 187.735 ;
        RECT 106.735 186.895 107.065 187.395 ;
        RECT 107.235 187.065 107.490 187.565 ;
        RECT 107.665 186.895 108.875 187.985 ;
        RECT 110.640 187.330 110.990 188.580 ;
        RECT 112.470 188.070 112.810 188.900 ;
        RECT 114.565 188.720 114.855 189.445 ;
        RECT 115.490 188.735 115.745 189.265 ;
        RECT 115.915 188.985 116.220 189.445 ;
        RECT 116.465 189.065 117.535 189.235 ;
        RECT 115.490 188.085 115.700 188.735 ;
        RECT 116.465 188.710 116.785 189.065 ;
        RECT 116.460 188.535 116.785 188.710 ;
        RECT 115.870 188.235 116.785 188.535 ;
        RECT 116.955 188.495 117.195 188.895 ;
        RECT 117.365 188.835 117.535 189.065 ;
        RECT 117.705 189.005 117.895 189.445 ;
        RECT 118.065 188.995 119.015 189.275 ;
        RECT 119.235 189.085 119.585 189.255 ;
        RECT 117.365 188.665 117.895 188.835 ;
        RECT 115.870 188.205 116.610 188.235 ;
        RECT 109.050 186.895 114.395 187.330 ;
        RECT 114.565 186.895 114.855 188.060 ;
        RECT 115.490 187.205 115.745 188.085 ;
        RECT 115.915 186.895 116.220 188.035 ;
        RECT 116.440 187.615 116.610 188.205 ;
        RECT 116.955 188.125 117.495 188.495 ;
        RECT 117.675 188.385 117.895 188.665 ;
        RECT 118.065 188.215 118.235 188.995 ;
        RECT 117.830 188.045 118.235 188.215 ;
        RECT 118.405 188.205 118.755 188.825 ;
        RECT 117.830 187.955 118.000 188.045 ;
        RECT 118.925 188.035 119.135 188.825 ;
        RECT 116.780 187.785 118.000 187.955 ;
        RECT 118.460 187.875 119.135 188.035 ;
        RECT 116.440 187.445 117.240 187.615 ;
        RECT 116.560 186.895 116.890 187.275 ;
        RECT 117.070 187.155 117.240 187.445 ;
        RECT 117.830 187.405 118.000 187.785 ;
        RECT 118.170 187.865 119.135 187.875 ;
        RECT 119.325 188.695 119.585 189.085 ;
        RECT 119.795 188.985 120.125 189.445 ;
        RECT 121.000 189.055 121.855 189.225 ;
        RECT 122.060 189.055 122.555 189.225 ;
        RECT 122.725 189.085 123.055 189.445 ;
        RECT 119.325 188.005 119.495 188.695 ;
        RECT 119.665 188.345 119.835 188.525 ;
        RECT 120.005 188.515 120.795 188.765 ;
        RECT 121.000 188.345 121.170 189.055 ;
        RECT 121.340 188.545 121.695 188.765 ;
        RECT 119.665 188.175 121.355 188.345 ;
        RECT 118.170 187.575 118.630 187.865 ;
        RECT 119.325 187.835 120.825 188.005 ;
        RECT 119.325 187.695 119.495 187.835 ;
        RECT 118.935 187.525 119.495 187.695 ;
        RECT 117.410 186.895 117.660 187.355 ;
        RECT 117.830 187.065 118.700 187.405 ;
        RECT 118.935 187.065 119.105 187.525 ;
        RECT 119.940 187.495 121.015 187.665 ;
        RECT 119.275 186.895 119.645 187.355 ;
        RECT 119.940 187.155 120.110 187.495 ;
        RECT 120.280 186.895 120.610 187.325 ;
        RECT 120.845 187.155 121.015 187.495 ;
        RECT 121.185 187.395 121.355 188.175 ;
        RECT 121.525 187.955 121.695 188.545 ;
        RECT 121.865 188.145 122.215 188.765 ;
        RECT 121.525 187.565 121.990 187.955 ;
        RECT 122.385 187.695 122.555 189.055 ;
        RECT 122.725 187.865 123.185 188.915 ;
        RECT 122.160 187.525 122.555 187.695 ;
        RECT 122.160 187.395 122.330 187.525 ;
        RECT 121.185 187.065 121.865 187.395 ;
        RECT 122.080 187.065 122.330 187.395 ;
        RECT 122.500 186.895 122.750 187.355 ;
        RECT 122.920 187.080 123.245 187.865 ;
        RECT 123.415 187.065 123.585 189.185 ;
        RECT 123.755 189.065 124.085 189.445 ;
        RECT 124.255 188.895 124.510 189.185 ;
        RECT 123.760 188.725 124.510 188.895 ;
        RECT 123.760 187.735 123.990 188.725 ;
        RECT 124.685 188.675 126.355 189.445 ;
        RECT 126.525 188.695 127.735 189.445 ;
        RECT 124.160 187.905 124.510 188.555 ;
        RECT 124.685 187.985 125.435 188.505 ;
        RECT 125.605 188.155 126.355 188.675 ;
        RECT 126.525 187.985 127.045 188.525 ;
        RECT 127.215 188.155 127.735 188.695 ;
        RECT 123.760 187.565 124.510 187.735 ;
        RECT 123.755 186.895 124.085 187.395 ;
        RECT 124.255 187.065 124.510 187.565 ;
        RECT 124.685 186.895 126.355 187.985 ;
        RECT 126.525 186.895 127.735 187.985 ;
        RECT 14.660 186.725 127.820 186.895 ;
        RECT 14.745 185.635 15.955 186.725 ;
        RECT 14.745 184.925 15.265 185.465 ;
        RECT 15.435 185.095 15.955 185.635 ;
        RECT 16.125 185.635 18.715 186.725 ;
        RECT 18.890 186.290 24.235 186.725 ;
        RECT 16.125 185.115 17.335 185.635 ;
        RECT 17.505 184.945 18.715 185.465 ;
        RECT 20.480 185.040 20.830 186.290 ;
        RECT 24.405 185.560 24.695 186.725 ;
        RECT 24.870 186.055 25.125 186.555 ;
        RECT 25.295 186.225 25.625 186.725 ;
        RECT 24.870 185.885 25.620 186.055 ;
        RECT 14.745 184.175 15.955 184.925 ;
        RECT 16.125 184.175 18.715 184.945 ;
        RECT 22.310 184.720 22.650 185.550 ;
        RECT 24.870 185.065 25.220 185.715 ;
        RECT 18.890 184.175 24.235 184.720 ;
        RECT 24.405 184.175 24.695 184.900 ;
        RECT 25.390 184.895 25.620 185.885 ;
        RECT 24.870 184.725 25.620 184.895 ;
        RECT 24.870 184.435 25.125 184.725 ;
        RECT 25.295 184.175 25.625 184.555 ;
        RECT 25.795 184.435 25.965 186.555 ;
        RECT 26.135 185.755 26.460 186.540 ;
        RECT 26.630 186.265 26.880 186.725 ;
        RECT 27.050 186.225 27.300 186.555 ;
        RECT 27.515 186.225 28.195 186.555 ;
        RECT 27.050 186.095 27.220 186.225 ;
        RECT 26.825 185.925 27.220 186.095 ;
        RECT 26.195 184.705 26.655 185.755 ;
        RECT 26.825 184.565 26.995 185.925 ;
        RECT 27.390 185.665 27.855 186.055 ;
        RECT 27.165 184.855 27.515 185.475 ;
        RECT 27.685 185.075 27.855 185.665 ;
        RECT 28.025 185.445 28.195 186.225 ;
        RECT 28.365 186.125 28.535 186.465 ;
        RECT 28.770 186.295 29.100 186.725 ;
        RECT 29.270 186.125 29.440 186.465 ;
        RECT 29.735 186.265 30.105 186.725 ;
        RECT 28.365 185.955 29.440 186.125 ;
        RECT 30.275 186.095 30.445 186.555 ;
        RECT 30.680 186.215 31.550 186.555 ;
        RECT 31.720 186.265 31.970 186.725 ;
        RECT 29.885 185.925 30.445 186.095 ;
        RECT 29.885 185.785 30.055 185.925 ;
        RECT 28.555 185.615 30.055 185.785 ;
        RECT 30.750 185.755 31.210 186.045 ;
        RECT 28.025 185.275 29.715 185.445 ;
        RECT 27.685 184.855 28.040 185.075 ;
        RECT 28.210 184.565 28.380 185.275 ;
        RECT 28.585 184.855 29.375 185.105 ;
        RECT 29.545 185.095 29.715 185.275 ;
        RECT 29.885 184.925 30.055 185.615 ;
        RECT 26.325 184.175 26.655 184.535 ;
        RECT 26.825 184.395 27.320 184.565 ;
        RECT 27.525 184.395 28.380 184.565 ;
        RECT 29.255 184.175 29.585 184.635 ;
        RECT 29.795 184.535 30.055 184.925 ;
        RECT 30.245 185.745 31.210 185.755 ;
        RECT 31.380 185.835 31.550 186.215 ;
        RECT 32.140 186.175 32.310 186.465 ;
        RECT 32.490 186.345 32.820 186.725 ;
        RECT 32.140 186.005 32.940 186.175 ;
        RECT 30.245 185.585 30.920 185.745 ;
        RECT 31.380 185.665 32.600 185.835 ;
        RECT 30.245 184.795 30.455 185.585 ;
        RECT 31.380 185.575 31.550 185.665 ;
        RECT 30.625 184.795 30.975 185.415 ;
        RECT 31.145 185.405 31.550 185.575 ;
        RECT 31.145 184.625 31.315 185.405 ;
        RECT 31.485 184.955 31.705 185.235 ;
        RECT 31.885 185.125 32.425 185.495 ;
        RECT 32.770 185.415 32.940 186.005 ;
        RECT 33.160 185.585 33.465 186.725 ;
        RECT 33.635 185.535 33.890 186.415 ;
        RECT 34.990 186.290 40.335 186.725 ;
        RECT 40.510 186.290 45.855 186.725 ;
        RECT 32.770 185.385 33.510 185.415 ;
        RECT 31.485 184.785 32.015 184.955 ;
        RECT 29.795 184.365 30.145 184.535 ;
        RECT 30.365 184.345 31.315 184.625 ;
        RECT 31.485 184.175 31.675 184.615 ;
        RECT 31.845 184.555 32.015 184.785 ;
        RECT 32.185 184.725 32.425 185.125 ;
        RECT 32.595 185.085 33.510 185.385 ;
        RECT 32.595 184.910 32.920 185.085 ;
        RECT 32.595 184.555 32.915 184.910 ;
        RECT 33.680 184.885 33.890 185.535 ;
        RECT 36.580 185.040 36.930 186.290 ;
        RECT 31.845 184.385 32.915 184.555 ;
        RECT 33.160 184.175 33.465 184.635 ;
        RECT 33.635 184.355 33.890 184.885 ;
        RECT 38.410 184.720 38.750 185.550 ;
        RECT 42.100 185.040 42.450 186.290 ;
        RECT 46.025 185.965 46.540 186.375 ;
        RECT 46.775 185.965 46.945 186.725 ;
        RECT 47.115 186.385 49.145 186.555 ;
        RECT 43.930 184.720 44.270 185.550 ;
        RECT 46.025 185.155 46.365 185.965 ;
        RECT 47.115 185.720 47.285 186.385 ;
        RECT 47.680 186.045 48.805 186.215 ;
        RECT 46.535 185.530 47.285 185.720 ;
        RECT 47.455 185.705 48.465 185.875 ;
        RECT 46.025 184.985 47.255 185.155 ;
        RECT 34.990 184.175 40.335 184.720 ;
        RECT 40.510 184.175 45.855 184.720 ;
        RECT 46.300 184.380 46.545 184.985 ;
        RECT 46.765 184.175 47.275 184.710 ;
        RECT 47.455 184.345 47.645 185.705 ;
        RECT 47.815 185.365 48.090 185.505 ;
        RECT 47.815 185.195 48.095 185.365 ;
        RECT 47.815 184.345 48.090 185.195 ;
        RECT 48.295 184.905 48.465 185.705 ;
        RECT 48.635 184.915 48.805 186.045 ;
        RECT 48.975 185.415 49.145 186.385 ;
        RECT 49.315 185.585 49.485 186.725 ;
        RECT 49.655 185.585 49.990 186.555 ;
        RECT 48.975 185.085 49.170 185.415 ;
        RECT 49.395 185.085 49.650 185.415 ;
        RECT 49.395 184.915 49.565 185.085 ;
        RECT 49.820 184.915 49.990 185.585 ;
        RECT 50.165 185.560 50.455 186.725 ;
        RECT 51.585 185.585 51.815 186.725 ;
        RECT 51.985 185.575 52.315 186.555 ;
        RECT 52.485 185.585 52.695 186.725 ;
        RECT 52.925 185.635 55.515 186.725 ;
        RECT 55.775 185.795 55.945 186.555 ;
        RECT 56.125 185.965 56.455 186.725 ;
        RECT 51.565 185.165 51.895 185.415 ;
        RECT 48.635 184.745 49.565 184.915 ;
        RECT 48.635 184.710 48.810 184.745 ;
        RECT 48.280 184.345 48.810 184.710 ;
        RECT 49.235 184.175 49.565 184.575 ;
        RECT 49.735 184.345 49.990 184.915 ;
        RECT 50.165 184.175 50.455 184.900 ;
        RECT 51.585 184.175 51.815 184.995 ;
        RECT 52.065 184.975 52.315 185.575 ;
        RECT 52.925 185.115 54.135 185.635 ;
        RECT 55.775 185.625 56.440 185.795 ;
        RECT 56.625 185.650 56.895 186.555 ;
        RECT 56.270 185.480 56.440 185.625 ;
        RECT 51.985 184.345 52.315 184.975 ;
        RECT 52.485 184.175 52.695 184.995 ;
        RECT 54.305 184.945 55.515 185.465 ;
        RECT 55.705 185.075 56.035 185.445 ;
        RECT 56.270 185.150 56.555 185.480 ;
        RECT 52.925 184.175 55.515 184.945 ;
        RECT 56.270 184.895 56.440 185.150 ;
        RECT 55.775 184.725 56.440 184.895 ;
        RECT 56.725 184.850 56.895 185.650 ;
        RECT 57.125 185.585 57.335 186.725 ;
        RECT 57.505 185.575 57.835 186.555 ;
        RECT 58.005 185.585 58.235 186.725 ;
        RECT 58.445 185.635 61.035 186.725 ;
        RECT 61.210 186.290 66.555 186.725 ;
        RECT 55.775 184.345 55.945 184.725 ;
        RECT 56.125 184.175 56.455 184.555 ;
        RECT 56.635 184.345 56.895 184.850 ;
        RECT 57.125 184.175 57.335 184.995 ;
        RECT 57.505 184.975 57.755 185.575 ;
        RECT 57.925 185.165 58.255 185.415 ;
        RECT 58.445 185.115 59.655 185.635 ;
        RECT 57.505 184.345 57.835 184.975 ;
        RECT 58.005 184.175 58.235 184.995 ;
        RECT 59.825 184.945 61.035 185.465 ;
        RECT 62.800 185.040 63.150 186.290 ;
        RECT 58.445 184.175 61.035 184.945 ;
        RECT 64.630 184.720 64.970 185.550 ;
        RECT 66.730 185.535 66.985 186.415 ;
        RECT 67.155 185.585 67.460 186.725 ;
        RECT 67.800 186.345 68.130 186.725 ;
        RECT 68.310 186.175 68.480 186.465 ;
        RECT 68.650 186.265 68.900 186.725 ;
        RECT 67.680 186.005 68.480 186.175 ;
        RECT 69.070 186.215 69.940 186.555 ;
        RECT 66.730 184.885 66.940 185.535 ;
        RECT 67.680 185.415 67.850 186.005 ;
        RECT 69.070 185.835 69.240 186.215 ;
        RECT 70.175 186.095 70.345 186.555 ;
        RECT 70.515 186.265 70.885 186.725 ;
        RECT 71.180 186.125 71.350 186.465 ;
        RECT 71.520 186.295 71.850 186.725 ;
        RECT 72.085 186.125 72.255 186.465 ;
        RECT 68.020 185.665 69.240 185.835 ;
        RECT 69.410 185.755 69.870 186.045 ;
        RECT 70.175 185.925 70.735 186.095 ;
        RECT 71.180 185.955 72.255 186.125 ;
        RECT 72.425 186.225 73.105 186.555 ;
        RECT 73.320 186.225 73.570 186.555 ;
        RECT 73.740 186.265 73.990 186.725 ;
        RECT 70.565 185.785 70.735 185.925 ;
        RECT 69.410 185.745 70.375 185.755 ;
        RECT 69.070 185.575 69.240 185.665 ;
        RECT 69.700 185.585 70.375 185.745 ;
        RECT 67.110 185.385 67.850 185.415 ;
        RECT 67.110 185.085 68.025 185.385 ;
        RECT 67.700 184.910 68.025 185.085 ;
        RECT 61.210 184.175 66.555 184.720 ;
        RECT 66.730 184.355 66.985 184.885 ;
        RECT 67.155 184.175 67.460 184.635 ;
        RECT 67.705 184.555 68.025 184.910 ;
        RECT 68.195 185.125 68.735 185.495 ;
        RECT 69.070 185.405 69.475 185.575 ;
        RECT 68.195 184.725 68.435 185.125 ;
        RECT 68.915 184.955 69.135 185.235 ;
        RECT 68.605 184.785 69.135 184.955 ;
        RECT 68.605 184.555 68.775 184.785 ;
        RECT 69.305 184.625 69.475 185.405 ;
        RECT 69.645 184.795 69.995 185.415 ;
        RECT 70.165 184.795 70.375 185.585 ;
        RECT 70.565 185.615 72.065 185.785 ;
        RECT 70.565 184.925 70.735 185.615 ;
        RECT 72.425 185.445 72.595 186.225 ;
        RECT 73.400 186.095 73.570 186.225 ;
        RECT 70.905 185.275 72.595 185.445 ;
        RECT 72.765 185.665 73.230 186.055 ;
        RECT 73.400 185.925 73.795 186.095 ;
        RECT 70.905 185.095 71.075 185.275 ;
        RECT 67.705 184.385 68.775 184.555 ;
        RECT 68.945 184.175 69.135 184.615 ;
        RECT 69.305 184.345 70.255 184.625 ;
        RECT 70.565 184.535 70.825 184.925 ;
        RECT 71.245 184.855 72.035 185.105 ;
        RECT 70.475 184.365 70.825 184.535 ;
        RECT 71.035 184.175 71.365 184.635 ;
        RECT 72.240 184.565 72.410 185.275 ;
        RECT 72.765 185.075 72.935 185.665 ;
        RECT 72.580 184.855 72.935 185.075 ;
        RECT 73.105 184.855 73.455 185.475 ;
        RECT 73.625 184.565 73.795 185.925 ;
        RECT 74.160 185.755 74.485 186.540 ;
        RECT 73.965 184.705 74.425 185.755 ;
        RECT 72.240 184.395 73.095 184.565 ;
        RECT 73.300 184.395 73.795 184.565 ;
        RECT 73.965 184.175 74.295 184.535 ;
        RECT 74.655 184.435 74.825 186.555 ;
        RECT 74.995 186.225 75.325 186.725 ;
        RECT 75.495 186.055 75.750 186.555 ;
        RECT 75.000 185.885 75.750 186.055 ;
        RECT 75.000 184.895 75.230 185.885 ;
        RECT 75.400 185.065 75.750 185.715 ;
        RECT 75.925 185.560 76.215 186.725 ;
        RECT 76.445 185.585 76.655 186.725 ;
        RECT 76.825 185.575 77.155 186.555 ;
        RECT 77.325 185.585 77.555 186.725 ;
        RECT 78.225 185.635 79.895 186.725 ;
        RECT 80.070 186.290 85.415 186.725 ;
        RECT 75.000 184.725 75.750 184.895 ;
        RECT 74.995 184.175 75.325 184.555 ;
        RECT 75.495 184.435 75.750 184.725 ;
        RECT 75.925 184.175 76.215 184.900 ;
        RECT 76.445 184.175 76.655 184.995 ;
        RECT 76.825 184.975 77.075 185.575 ;
        RECT 77.245 185.165 77.575 185.415 ;
        RECT 78.225 185.115 78.975 185.635 ;
        RECT 76.825 184.345 77.155 184.975 ;
        RECT 77.325 184.175 77.555 184.995 ;
        RECT 79.145 184.945 79.895 185.465 ;
        RECT 81.660 185.040 82.010 186.290 ;
        RECT 85.585 185.965 86.100 186.375 ;
        RECT 86.335 185.965 86.505 186.725 ;
        RECT 86.675 186.385 88.705 186.555 ;
        RECT 78.225 184.175 79.895 184.945 ;
        RECT 83.490 184.720 83.830 185.550 ;
        RECT 85.585 185.155 85.925 185.965 ;
        RECT 86.675 185.720 86.845 186.385 ;
        RECT 87.240 186.045 88.365 186.215 ;
        RECT 86.095 185.530 86.845 185.720 ;
        RECT 87.015 185.705 88.025 185.875 ;
        RECT 85.585 184.985 86.815 185.155 ;
        RECT 80.070 184.175 85.415 184.720 ;
        RECT 85.860 184.380 86.105 184.985 ;
        RECT 86.325 184.175 86.835 184.710 ;
        RECT 87.015 184.345 87.205 185.705 ;
        RECT 87.375 185.025 87.650 185.505 ;
        RECT 87.375 184.855 87.655 185.025 ;
        RECT 87.855 184.905 88.025 185.705 ;
        RECT 88.195 184.915 88.365 186.045 ;
        RECT 88.535 185.415 88.705 186.385 ;
        RECT 88.875 185.585 89.045 186.725 ;
        RECT 89.215 185.585 89.550 186.555 ;
        RECT 90.650 186.290 95.995 186.725 ;
        RECT 96.170 186.290 101.515 186.725 ;
        RECT 88.535 185.085 88.730 185.415 ;
        RECT 88.955 185.085 89.210 185.415 ;
        RECT 88.955 184.915 89.125 185.085 ;
        RECT 89.380 184.915 89.550 185.585 ;
        RECT 92.240 185.040 92.590 186.290 ;
        RECT 87.375 184.345 87.650 184.855 ;
        RECT 88.195 184.745 89.125 184.915 ;
        RECT 88.195 184.710 88.370 184.745 ;
        RECT 87.840 184.345 88.370 184.710 ;
        RECT 88.795 184.175 89.125 184.575 ;
        RECT 89.295 184.345 89.550 184.915 ;
        RECT 94.070 184.720 94.410 185.550 ;
        RECT 97.760 185.040 98.110 186.290 ;
        RECT 101.685 185.560 101.975 186.725 ;
        RECT 102.605 185.965 103.120 186.375 ;
        RECT 103.355 185.965 103.525 186.725 ;
        RECT 103.695 186.385 105.725 186.555 ;
        RECT 99.590 184.720 99.930 185.550 ;
        RECT 102.605 185.155 102.945 185.965 ;
        RECT 103.695 185.720 103.865 186.385 ;
        RECT 104.260 186.045 105.385 186.215 ;
        RECT 103.115 185.530 103.865 185.720 ;
        RECT 104.035 185.705 105.045 185.875 ;
        RECT 102.605 184.985 103.835 185.155 ;
        RECT 90.650 184.175 95.995 184.720 ;
        RECT 96.170 184.175 101.515 184.720 ;
        RECT 101.685 184.175 101.975 184.900 ;
        RECT 102.880 184.380 103.125 184.985 ;
        RECT 103.345 184.175 103.855 184.710 ;
        RECT 104.035 184.345 104.225 185.705 ;
        RECT 104.395 184.685 104.670 185.505 ;
        RECT 104.875 184.905 105.045 185.705 ;
        RECT 105.215 184.915 105.385 186.045 ;
        RECT 105.555 185.415 105.725 186.385 ;
        RECT 105.895 185.585 106.065 186.725 ;
        RECT 106.235 185.585 106.570 186.555 ;
        RECT 105.555 185.085 105.750 185.415 ;
        RECT 105.975 185.085 106.230 185.415 ;
        RECT 105.975 184.915 106.145 185.085 ;
        RECT 106.400 184.915 106.570 185.585 ;
        RECT 105.215 184.745 106.145 184.915 ;
        RECT 105.215 184.710 105.390 184.745 ;
        RECT 104.395 184.515 104.675 184.685 ;
        RECT 104.395 184.345 104.670 184.515 ;
        RECT 104.860 184.345 105.390 184.710 ;
        RECT 105.815 184.175 106.145 184.575 ;
        RECT 106.315 184.345 106.570 184.915 ;
        RECT 106.745 185.650 107.015 186.555 ;
        RECT 107.185 185.965 107.515 186.725 ;
        RECT 107.695 185.795 107.865 186.555 ;
        RECT 106.745 184.850 106.915 185.650 ;
        RECT 107.200 185.625 107.865 185.795 ;
        RECT 108.125 185.635 109.335 186.725 ;
        RECT 107.200 185.480 107.370 185.625 ;
        RECT 107.085 185.150 107.370 185.480 ;
        RECT 107.200 184.895 107.370 185.150 ;
        RECT 107.605 185.075 107.935 185.445 ;
        RECT 108.125 185.095 108.645 185.635 ;
        RECT 109.545 185.585 109.775 186.725 ;
        RECT 109.945 185.575 110.275 186.555 ;
        RECT 110.445 185.585 110.655 186.725 ;
        RECT 108.815 184.925 109.335 185.465 ;
        RECT 109.525 185.165 109.855 185.415 ;
        RECT 106.745 184.345 107.005 184.850 ;
        RECT 107.200 184.725 107.865 184.895 ;
        RECT 107.185 184.175 107.515 184.555 ;
        RECT 107.695 184.345 107.865 184.725 ;
        RECT 108.125 184.175 109.335 184.925 ;
        RECT 109.545 184.175 109.775 184.995 ;
        RECT 110.025 184.975 110.275 185.575 ;
        RECT 110.890 185.535 111.145 186.415 ;
        RECT 111.315 185.585 111.620 186.725 ;
        RECT 111.960 186.345 112.290 186.725 ;
        RECT 112.470 186.175 112.640 186.465 ;
        RECT 112.810 186.265 113.060 186.725 ;
        RECT 111.840 186.005 112.640 186.175 ;
        RECT 113.230 186.215 114.100 186.555 ;
        RECT 109.945 184.345 110.275 184.975 ;
        RECT 110.445 184.175 110.655 184.995 ;
        RECT 110.890 184.885 111.100 185.535 ;
        RECT 111.840 185.415 112.010 186.005 ;
        RECT 113.230 185.835 113.400 186.215 ;
        RECT 114.335 186.095 114.505 186.555 ;
        RECT 114.675 186.265 115.045 186.725 ;
        RECT 115.340 186.125 115.510 186.465 ;
        RECT 115.680 186.295 116.010 186.725 ;
        RECT 116.245 186.125 116.415 186.465 ;
        RECT 112.180 185.665 113.400 185.835 ;
        RECT 113.570 185.755 114.030 186.045 ;
        RECT 114.335 185.925 114.895 186.095 ;
        RECT 115.340 185.955 116.415 186.125 ;
        RECT 116.585 186.225 117.265 186.555 ;
        RECT 117.480 186.225 117.730 186.555 ;
        RECT 117.900 186.265 118.150 186.725 ;
        RECT 114.725 185.785 114.895 185.925 ;
        RECT 113.570 185.745 114.535 185.755 ;
        RECT 113.230 185.575 113.400 185.665 ;
        RECT 113.860 185.585 114.535 185.745 ;
        RECT 111.270 185.385 112.010 185.415 ;
        RECT 111.270 185.085 112.185 185.385 ;
        RECT 111.860 184.910 112.185 185.085 ;
        RECT 110.890 184.355 111.145 184.885 ;
        RECT 111.315 184.175 111.620 184.635 ;
        RECT 111.865 184.555 112.185 184.910 ;
        RECT 112.355 185.125 112.895 185.495 ;
        RECT 113.230 185.405 113.635 185.575 ;
        RECT 112.355 184.725 112.595 185.125 ;
        RECT 113.075 184.955 113.295 185.235 ;
        RECT 112.765 184.785 113.295 184.955 ;
        RECT 112.765 184.555 112.935 184.785 ;
        RECT 113.465 184.625 113.635 185.405 ;
        RECT 113.805 184.795 114.155 185.415 ;
        RECT 114.325 184.795 114.535 185.585 ;
        RECT 114.725 185.615 116.225 185.785 ;
        RECT 114.725 184.925 114.895 185.615 ;
        RECT 116.585 185.445 116.755 186.225 ;
        RECT 117.560 186.095 117.730 186.225 ;
        RECT 115.065 185.275 116.755 185.445 ;
        RECT 116.925 185.665 117.390 186.055 ;
        RECT 117.560 185.925 117.955 186.095 ;
        RECT 115.065 185.095 115.235 185.275 ;
        RECT 111.865 184.385 112.935 184.555 ;
        RECT 113.105 184.175 113.295 184.615 ;
        RECT 113.465 184.345 114.415 184.625 ;
        RECT 114.725 184.535 114.985 184.925 ;
        RECT 115.405 184.855 116.195 185.105 ;
        RECT 114.635 184.365 114.985 184.535 ;
        RECT 115.195 184.175 115.525 184.635 ;
        RECT 116.400 184.565 116.570 185.275 ;
        RECT 116.925 185.075 117.095 185.665 ;
        RECT 116.740 184.855 117.095 185.075 ;
        RECT 117.265 184.855 117.615 185.475 ;
        RECT 117.785 184.565 117.955 185.925 ;
        RECT 118.320 185.755 118.645 186.540 ;
        RECT 118.125 184.705 118.585 185.755 ;
        RECT 116.400 184.395 117.255 184.565 ;
        RECT 117.460 184.395 117.955 184.565 ;
        RECT 118.125 184.175 118.455 184.535 ;
        RECT 118.815 184.435 118.985 186.555 ;
        RECT 119.155 186.225 119.485 186.725 ;
        RECT 119.655 186.055 119.910 186.555 ;
        RECT 119.160 185.885 119.910 186.055 ;
        RECT 119.160 184.895 119.390 185.885 ;
        RECT 119.560 185.065 119.910 185.715 ;
        RECT 120.125 185.585 120.355 186.725 ;
        RECT 120.525 185.575 120.855 186.555 ;
        RECT 121.025 185.585 121.235 186.725 ;
        RECT 121.555 185.795 121.725 186.555 ;
        RECT 121.905 185.965 122.235 186.725 ;
        RECT 121.555 185.625 122.220 185.795 ;
        RECT 122.405 185.650 122.675 186.555 ;
        RECT 120.105 185.165 120.435 185.415 ;
        RECT 119.160 184.725 119.910 184.895 ;
        RECT 119.155 184.175 119.485 184.555 ;
        RECT 119.655 184.435 119.910 184.725 ;
        RECT 120.125 184.175 120.355 184.995 ;
        RECT 120.605 184.975 120.855 185.575 ;
        RECT 122.050 185.480 122.220 185.625 ;
        RECT 121.485 185.075 121.815 185.445 ;
        RECT 122.050 185.150 122.335 185.480 ;
        RECT 120.525 184.345 120.855 184.975 ;
        RECT 121.025 184.175 121.235 184.995 ;
        RECT 122.050 184.895 122.220 185.150 ;
        RECT 121.555 184.725 122.220 184.895 ;
        RECT 122.505 184.850 122.675 185.650 ;
        RECT 122.845 185.635 126.355 186.725 ;
        RECT 126.525 185.635 127.735 186.725 ;
        RECT 122.845 185.115 124.535 185.635 ;
        RECT 124.705 184.945 126.355 185.465 ;
        RECT 126.525 185.095 127.045 185.635 ;
        RECT 121.555 184.345 121.725 184.725 ;
        RECT 121.905 184.175 122.235 184.555 ;
        RECT 122.415 184.345 122.675 184.850 ;
        RECT 122.845 184.175 126.355 184.945 ;
        RECT 127.215 184.925 127.735 185.465 ;
        RECT 126.525 184.175 127.735 184.925 ;
        RECT 14.660 184.005 127.820 184.175 ;
        RECT 14.745 183.255 15.955 184.005 ;
        RECT 16.590 183.460 21.935 184.005 ;
        RECT 22.110 183.460 27.455 184.005 ;
        RECT 14.745 182.715 15.265 183.255 ;
        RECT 15.435 182.545 15.955 183.085 ;
        RECT 14.745 181.455 15.955 182.545 ;
        RECT 18.180 181.890 18.530 183.140 ;
        RECT 20.010 182.630 20.350 183.460 ;
        RECT 23.700 181.890 24.050 183.140 ;
        RECT 25.530 182.630 25.870 183.460 ;
        RECT 27.625 183.330 27.885 183.835 ;
        RECT 28.065 183.625 28.395 184.005 ;
        RECT 28.575 183.455 28.745 183.835 ;
        RECT 27.625 182.530 27.795 183.330 ;
        RECT 28.080 183.285 28.745 183.455 ;
        RECT 28.080 183.030 28.250 183.285 ;
        RECT 29.010 183.265 29.265 183.835 ;
        RECT 29.435 183.605 29.765 184.005 ;
        RECT 30.190 183.470 30.720 183.835 ;
        RECT 30.190 183.435 30.365 183.470 ;
        RECT 29.435 183.265 30.365 183.435 ;
        RECT 27.965 182.700 28.250 183.030 ;
        RECT 28.485 182.735 28.815 183.105 ;
        RECT 28.080 182.555 28.250 182.700 ;
        RECT 29.010 182.595 29.180 183.265 ;
        RECT 29.435 183.095 29.605 183.265 ;
        RECT 29.350 182.765 29.605 183.095 ;
        RECT 29.830 182.765 30.025 183.095 ;
        RECT 16.590 181.455 21.935 181.890 ;
        RECT 22.110 181.455 27.455 181.890 ;
        RECT 27.625 181.625 27.895 182.530 ;
        RECT 28.080 182.385 28.745 182.555 ;
        RECT 28.065 181.455 28.395 182.215 ;
        RECT 28.575 181.625 28.745 182.385 ;
        RECT 29.010 181.625 29.345 182.595 ;
        RECT 29.515 181.455 29.685 182.595 ;
        RECT 29.855 181.795 30.025 182.765 ;
        RECT 30.195 182.135 30.365 183.265 ;
        RECT 30.535 182.475 30.705 183.275 ;
        RECT 30.910 182.985 31.185 183.835 ;
        RECT 30.905 182.815 31.185 182.985 ;
        RECT 30.910 182.675 31.185 182.815 ;
        RECT 31.355 182.475 31.545 183.835 ;
        RECT 31.725 183.470 32.235 184.005 ;
        RECT 32.455 183.195 32.700 183.800 ;
        RECT 33.605 183.235 37.115 184.005 ;
        RECT 37.285 183.280 37.575 184.005 ;
        RECT 38.205 183.235 41.715 184.005 ;
        RECT 31.745 183.025 32.975 183.195 ;
        RECT 30.535 182.305 31.545 182.475 ;
        RECT 31.715 182.460 32.465 182.650 ;
        RECT 30.195 181.965 31.320 182.135 ;
        RECT 31.715 181.795 31.885 182.460 ;
        RECT 32.635 182.215 32.975 183.025 ;
        RECT 29.855 181.625 31.885 181.795 ;
        RECT 32.055 181.455 32.225 182.215 ;
        RECT 32.460 181.805 32.975 182.215 ;
        RECT 33.605 182.545 35.295 183.065 ;
        RECT 35.465 182.715 37.115 183.235 ;
        RECT 33.605 181.455 37.115 182.545 ;
        RECT 37.285 181.455 37.575 182.620 ;
        RECT 38.205 182.545 39.895 183.065 ;
        RECT 40.065 182.715 41.715 183.235 ;
        RECT 42.160 183.195 42.405 183.800 ;
        RECT 42.625 183.470 43.135 184.005 ;
        RECT 41.885 183.025 43.115 183.195 ;
        RECT 38.205 181.455 41.715 182.545 ;
        RECT 41.885 182.215 42.225 183.025 ;
        RECT 42.395 182.460 43.145 182.650 ;
        RECT 41.885 181.805 42.400 182.215 ;
        RECT 42.635 181.455 42.805 182.215 ;
        RECT 42.975 181.795 43.145 182.460 ;
        RECT 43.315 182.475 43.505 183.835 ;
        RECT 43.675 183.325 43.950 183.835 ;
        RECT 44.140 183.470 44.670 183.835 ;
        RECT 45.095 183.605 45.425 184.005 ;
        RECT 44.495 183.435 44.670 183.470 ;
        RECT 43.675 183.155 43.955 183.325 ;
        RECT 43.675 182.675 43.950 183.155 ;
        RECT 44.155 182.475 44.325 183.275 ;
        RECT 43.315 182.305 44.325 182.475 ;
        RECT 44.495 183.265 45.425 183.435 ;
        RECT 45.595 183.265 45.850 183.835 ;
        RECT 44.495 182.135 44.665 183.265 ;
        RECT 45.255 183.095 45.425 183.265 ;
        RECT 43.540 181.965 44.665 182.135 ;
        RECT 44.835 182.765 45.030 183.095 ;
        RECT 45.255 182.765 45.510 183.095 ;
        RECT 44.835 181.795 45.005 182.765 ;
        RECT 45.680 182.595 45.850 183.265 ;
        RECT 42.975 181.625 45.005 181.795 ;
        RECT 45.175 181.455 45.345 182.595 ;
        RECT 45.515 181.625 45.850 182.595 ;
        RECT 46.025 183.205 46.365 183.835 ;
        RECT 46.535 183.205 46.785 184.005 ;
        RECT 46.975 183.355 47.305 183.835 ;
        RECT 47.475 183.545 47.700 184.005 ;
        RECT 47.870 183.355 48.200 183.835 ;
        RECT 46.025 182.595 46.200 183.205 ;
        RECT 46.975 183.185 48.200 183.355 ;
        RECT 48.830 183.225 49.330 183.835 ;
        RECT 46.370 182.845 47.065 183.015 ;
        RECT 46.895 182.595 47.065 182.845 ;
        RECT 47.240 182.815 47.660 183.015 ;
        RECT 47.830 182.815 48.160 183.015 ;
        RECT 48.330 182.815 48.660 183.015 ;
        RECT 48.830 182.595 49.000 183.225 ;
        RECT 49.980 183.195 50.225 183.800 ;
        RECT 50.445 183.470 50.955 184.005 ;
        RECT 49.705 183.025 50.935 183.195 ;
        RECT 49.185 182.765 49.535 183.015 ;
        RECT 46.025 181.625 46.365 182.595 ;
        RECT 46.535 181.455 46.705 182.595 ;
        RECT 46.895 182.425 49.330 182.595 ;
        RECT 46.975 181.455 47.225 182.255 ;
        RECT 47.870 181.625 48.200 182.425 ;
        RECT 48.500 181.455 48.830 182.255 ;
        RECT 49.000 181.625 49.330 182.425 ;
        RECT 49.705 182.215 50.045 183.025 ;
        RECT 50.215 182.460 50.965 182.650 ;
        RECT 49.705 181.805 50.220 182.215 ;
        RECT 50.455 181.455 50.625 182.215 ;
        RECT 50.795 181.795 50.965 182.460 ;
        RECT 51.135 182.475 51.325 183.835 ;
        RECT 51.495 182.985 51.770 183.835 ;
        RECT 51.960 183.470 52.490 183.835 ;
        RECT 52.915 183.605 53.245 184.005 ;
        RECT 52.315 183.435 52.490 183.470 ;
        RECT 51.495 182.815 51.775 182.985 ;
        RECT 51.495 182.675 51.770 182.815 ;
        RECT 51.975 182.475 52.145 183.275 ;
        RECT 51.135 182.305 52.145 182.475 ;
        RECT 52.315 183.265 53.245 183.435 ;
        RECT 53.415 183.265 53.670 183.835 ;
        RECT 52.315 182.135 52.485 183.265 ;
        RECT 53.075 183.095 53.245 183.265 ;
        RECT 51.360 181.965 52.485 182.135 ;
        RECT 52.655 182.765 52.850 183.095 ;
        RECT 53.075 182.765 53.330 183.095 ;
        RECT 52.655 181.795 52.825 182.765 ;
        RECT 53.500 182.595 53.670 183.265 ;
        RECT 50.795 181.625 52.825 181.795 ;
        RECT 52.995 181.455 53.165 182.595 ;
        RECT 53.335 181.625 53.670 182.595 ;
        RECT 53.850 183.295 54.105 183.825 ;
        RECT 54.275 183.545 54.580 184.005 ;
        RECT 54.825 183.625 55.895 183.795 ;
        RECT 53.850 182.645 54.060 183.295 ;
        RECT 54.825 183.270 55.145 183.625 ;
        RECT 54.820 183.095 55.145 183.270 ;
        RECT 54.230 182.795 55.145 183.095 ;
        RECT 55.315 183.055 55.555 183.455 ;
        RECT 55.725 183.395 55.895 183.625 ;
        RECT 56.065 183.565 56.255 184.005 ;
        RECT 56.425 183.555 57.375 183.835 ;
        RECT 57.595 183.645 57.945 183.815 ;
        RECT 55.725 183.225 56.255 183.395 ;
        RECT 54.230 182.765 54.970 182.795 ;
        RECT 53.850 181.765 54.105 182.645 ;
        RECT 54.275 181.455 54.580 182.595 ;
        RECT 54.800 182.175 54.970 182.765 ;
        RECT 55.315 182.685 55.855 183.055 ;
        RECT 56.035 182.945 56.255 183.225 ;
        RECT 56.425 182.775 56.595 183.555 ;
        RECT 56.190 182.605 56.595 182.775 ;
        RECT 56.765 182.765 57.115 183.385 ;
        RECT 56.190 182.515 56.360 182.605 ;
        RECT 57.285 182.595 57.495 183.385 ;
        RECT 55.140 182.345 56.360 182.515 ;
        RECT 56.820 182.435 57.495 182.595 ;
        RECT 54.800 182.005 55.600 182.175 ;
        RECT 54.920 181.455 55.250 181.835 ;
        RECT 55.430 181.715 55.600 182.005 ;
        RECT 56.190 181.965 56.360 182.345 ;
        RECT 56.530 182.425 57.495 182.435 ;
        RECT 57.685 183.255 57.945 183.645 ;
        RECT 58.155 183.545 58.485 184.005 ;
        RECT 59.360 183.615 60.215 183.785 ;
        RECT 60.420 183.615 60.915 183.785 ;
        RECT 61.085 183.645 61.415 184.005 ;
        RECT 57.685 182.565 57.855 183.255 ;
        RECT 58.025 182.905 58.195 183.085 ;
        RECT 58.365 183.075 59.155 183.325 ;
        RECT 59.360 182.905 59.530 183.615 ;
        RECT 59.700 183.105 60.055 183.325 ;
        RECT 58.025 182.735 59.715 182.905 ;
        RECT 56.530 182.135 56.990 182.425 ;
        RECT 57.685 182.395 59.185 182.565 ;
        RECT 57.685 182.255 57.855 182.395 ;
        RECT 57.295 182.085 57.855 182.255 ;
        RECT 55.770 181.455 56.020 181.915 ;
        RECT 56.190 181.625 57.060 181.965 ;
        RECT 57.295 181.625 57.465 182.085 ;
        RECT 58.300 182.055 59.375 182.225 ;
        RECT 57.635 181.455 58.005 181.915 ;
        RECT 58.300 181.715 58.470 182.055 ;
        RECT 58.640 181.455 58.970 181.885 ;
        RECT 59.205 181.715 59.375 182.055 ;
        RECT 59.545 181.955 59.715 182.735 ;
        RECT 59.885 182.515 60.055 183.105 ;
        RECT 60.225 182.705 60.575 183.325 ;
        RECT 59.885 182.125 60.350 182.515 ;
        RECT 60.745 182.255 60.915 183.615 ;
        RECT 61.085 182.425 61.545 183.475 ;
        RECT 60.520 182.085 60.915 182.255 ;
        RECT 60.520 181.955 60.690 182.085 ;
        RECT 59.545 181.625 60.225 181.955 ;
        RECT 60.440 181.625 60.690 181.955 ;
        RECT 60.860 181.455 61.110 181.915 ;
        RECT 61.280 181.640 61.605 182.425 ;
        RECT 61.775 181.625 61.945 183.745 ;
        RECT 62.115 183.625 62.445 184.005 ;
        RECT 62.615 183.455 62.870 183.745 ;
        RECT 62.120 183.285 62.870 183.455 ;
        RECT 62.120 182.295 62.350 183.285 ;
        RECT 63.045 183.280 63.335 184.005 ;
        RECT 63.505 183.505 63.765 183.835 ;
        RECT 63.975 183.525 64.250 184.005 ;
        RECT 62.520 182.465 62.870 183.115 ;
        RECT 62.120 182.125 62.870 182.295 ;
        RECT 62.115 181.455 62.445 181.955 ;
        RECT 62.615 181.625 62.870 182.125 ;
        RECT 63.045 181.455 63.335 182.620 ;
        RECT 63.505 182.595 63.675 183.505 ;
        RECT 64.460 183.435 64.665 183.835 ;
        RECT 64.835 183.605 65.170 184.005 ;
        RECT 65.345 183.505 65.605 183.835 ;
        RECT 65.915 183.625 66.245 184.005 ;
        RECT 66.425 183.665 67.905 183.835 ;
        RECT 63.845 182.765 64.205 183.345 ;
        RECT 64.460 183.265 65.145 183.435 ;
        RECT 64.385 182.595 64.635 183.095 ;
        RECT 63.505 182.425 64.635 182.595 ;
        RECT 63.505 181.655 63.775 182.425 ;
        RECT 64.805 182.235 65.145 183.265 ;
        RECT 63.945 181.455 64.275 182.235 ;
        RECT 64.480 182.060 65.145 182.235 ;
        RECT 65.345 182.805 65.515 183.505 ;
        RECT 66.425 183.335 66.825 183.665 ;
        RECT 65.865 183.145 66.075 183.325 ;
        RECT 65.865 182.975 66.485 183.145 ;
        RECT 66.655 182.855 66.825 183.335 ;
        RECT 67.015 183.165 67.565 183.495 ;
        RECT 65.345 182.635 66.475 182.805 ;
        RECT 66.655 182.685 67.225 182.855 ;
        RECT 64.480 181.655 64.665 182.060 ;
        RECT 65.345 181.955 65.515 182.635 ;
        RECT 66.305 182.515 66.475 182.635 ;
        RECT 65.685 182.135 66.035 182.465 ;
        RECT 66.305 182.345 66.885 182.515 ;
        RECT 67.055 182.175 67.225 182.685 ;
        RECT 66.485 182.005 67.225 182.175 ;
        RECT 67.395 182.175 67.565 183.165 ;
        RECT 67.735 182.765 67.905 183.665 ;
        RECT 68.155 183.095 68.340 183.675 ;
        RECT 68.610 183.095 68.805 183.670 ;
        RECT 69.015 183.625 69.345 184.005 ;
        RECT 68.155 182.765 68.385 183.095 ;
        RECT 68.610 182.765 68.865 183.095 ;
        RECT 68.155 182.455 68.340 182.765 ;
        RECT 68.610 182.455 68.805 182.765 ;
        RECT 69.175 182.175 69.345 183.095 ;
        RECT 67.395 182.005 69.345 182.175 ;
        RECT 64.835 181.455 65.170 181.880 ;
        RECT 65.345 181.625 65.605 181.955 ;
        RECT 65.915 181.455 66.245 181.835 ;
        RECT 66.485 181.625 66.675 182.005 ;
        RECT 66.925 181.455 67.255 181.835 ;
        RECT 67.465 181.625 67.635 182.005 ;
        RECT 67.830 181.455 68.160 181.835 ;
        RECT 68.420 181.625 68.590 182.005 ;
        RECT 69.015 181.455 69.345 181.835 ;
        RECT 69.515 181.625 69.775 183.835 ;
        RECT 69.950 183.295 70.205 183.825 ;
        RECT 70.375 183.545 70.680 184.005 ;
        RECT 70.925 183.625 71.995 183.795 ;
        RECT 69.950 182.645 70.160 183.295 ;
        RECT 70.925 183.270 71.245 183.625 ;
        RECT 70.920 183.095 71.245 183.270 ;
        RECT 70.330 182.795 71.245 183.095 ;
        RECT 71.415 183.055 71.655 183.455 ;
        RECT 71.825 183.395 71.995 183.625 ;
        RECT 72.165 183.565 72.355 184.005 ;
        RECT 72.525 183.555 73.475 183.835 ;
        RECT 73.695 183.645 74.045 183.815 ;
        RECT 71.825 183.225 72.355 183.395 ;
        RECT 70.330 182.765 71.070 182.795 ;
        RECT 69.950 181.765 70.205 182.645 ;
        RECT 70.375 181.455 70.680 182.595 ;
        RECT 70.900 182.175 71.070 182.765 ;
        RECT 71.415 182.685 71.955 183.055 ;
        RECT 72.135 182.945 72.355 183.225 ;
        RECT 72.525 182.775 72.695 183.555 ;
        RECT 72.290 182.605 72.695 182.775 ;
        RECT 72.865 182.765 73.215 183.385 ;
        RECT 72.290 182.515 72.460 182.605 ;
        RECT 73.385 182.595 73.595 183.385 ;
        RECT 71.240 182.345 72.460 182.515 ;
        RECT 72.920 182.435 73.595 182.595 ;
        RECT 70.900 182.005 71.700 182.175 ;
        RECT 71.020 181.455 71.350 181.835 ;
        RECT 71.530 181.715 71.700 182.005 ;
        RECT 72.290 181.965 72.460 182.345 ;
        RECT 72.630 182.425 73.595 182.435 ;
        RECT 73.785 183.255 74.045 183.645 ;
        RECT 74.255 183.545 74.585 184.005 ;
        RECT 75.460 183.615 76.315 183.785 ;
        RECT 76.520 183.615 77.015 183.785 ;
        RECT 77.185 183.645 77.515 184.005 ;
        RECT 73.785 182.565 73.955 183.255 ;
        RECT 74.125 182.905 74.295 183.085 ;
        RECT 74.465 183.075 75.255 183.325 ;
        RECT 75.460 182.905 75.630 183.615 ;
        RECT 75.800 183.105 76.155 183.325 ;
        RECT 74.125 182.735 75.815 182.905 ;
        RECT 72.630 182.135 73.090 182.425 ;
        RECT 73.785 182.395 75.285 182.565 ;
        RECT 73.785 182.255 73.955 182.395 ;
        RECT 73.395 182.085 73.955 182.255 ;
        RECT 71.870 181.455 72.120 181.915 ;
        RECT 72.290 181.625 73.160 181.965 ;
        RECT 73.395 181.625 73.565 182.085 ;
        RECT 74.400 182.055 75.475 182.225 ;
        RECT 73.735 181.455 74.105 181.915 ;
        RECT 74.400 181.715 74.570 182.055 ;
        RECT 74.740 181.455 75.070 181.885 ;
        RECT 75.305 181.715 75.475 182.055 ;
        RECT 75.645 181.955 75.815 182.735 ;
        RECT 75.985 182.515 76.155 183.105 ;
        RECT 76.325 182.705 76.675 183.325 ;
        RECT 75.985 182.125 76.450 182.515 ;
        RECT 76.845 182.255 77.015 183.615 ;
        RECT 77.185 182.425 77.645 183.475 ;
        RECT 76.620 182.085 77.015 182.255 ;
        RECT 76.620 181.955 76.790 182.085 ;
        RECT 75.645 181.625 76.325 181.955 ;
        RECT 76.540 181.625 76.790 181.955 ;
        RECT 76.960 181.455 77.210 181.915 ;
        RECT 77.380 181.640 77.705 182.425 ;
        RECT 77.875 181.625 78.045 183.745 ;
        RECT 78.215 183.625 78.545 184.005 ;
        RECT 78.715 183.455 78.970 183.745 ;
        RECT 79.150 183.460 84.495 184.005 ;
        RECT 78.220 183.285 78.970 183.455 ;
        RECT 78.220 182.295 78.450 183.285 ;
        RECT 78.620 182.465 78.970 183.115 ;
        RECT 78.220 182.125 78.970 182.295 ;
        RECT 78.215 181.455 78.545 181.955 ;
        RECT 78.715 181.625 78.970 182.125 ;
        RECT 80.740 181.890 81.090 183.140 ;
        RECT 82.570 182.630 82.910 183.460 ;
        RECT 84.940 183.195 85.185 183.800 ;
        RECT 85.405 183.470 85.915 184.005 ;
        RECT 84.665 183.025 85.895 183.195 ;
        RECT 84.665 182.215 85.005 183.025 ;
        RECT 85.175 182.460 85.925 182.650 ;
        RECT 79.150 181.455 84.495 181.890 ;
        RECT 84.665 181.805 85.180 182.215 ;
        RECT 85.415 181.455 85.585 182.215 ;
        RECT 85.755 181.795 85.925 182.460 ;
        RECT 86.095 182.475 86.285 183.835 ;
        RECT 86.455 182.985 86.730 183.835 ;
        RECT 86.920 183.470 87.450 183.835 ;
        RECT 87.875 183.605 88.205 184.005 ;
        RECT 87.275 183.435 87.450 183.470 ;
        RECT 86.455 182.815 86.735 182.985 ;
        RECT 86.455 182.675 86.730 182.815 ;
        RECT 86.935 182.475 87.105 183.275 ;
        RECT 86.095 182.305 87.105 182.475 ;
        RECT 87.275 183.265 88.205 183.435 ;
        RECT 88.375 183.265 88.630 183.835 ;
        RECT 88.805 183.280 89.095 184.005 ;
        RECT 87.275 182.135 87.445 183.265 ;
        RECT 88.035 183.095 88.205 183.265 ;
        RECT 86.320 181.965 87.445 182.135 ;
        RECT 87.615 182.765 87.810 183.095 ;
        RECT 88.035 182.765 88.290 183.095 ;
        RECT 87.615 181.795 87.785 182.765 ;
        RECT 88.460 182.595 88.630 183.265 ;
        RECT 89.265 183.255 90.475 184.005 ;
        RECT 90.735 183.455 90.905 183.835 ;
        RECT 91.085 183.625 91.415 184.005 ;
        RECT 90.735 183.285 91.400 183.455 ;
        RECT 91.595 183.330 91.855 183.835 ;
        RECT 85.755 181.625 87.785 181.795 ;
        RECT 87.955 181.455 88.125 182.595 ;
        RECT 88.295 181.625 88.630 182.595 ;
        RECT 88.805 181.455 89.095 182.620 ;
        RECT 89.265 182.545 89.785 183.085 ;
        RECT 89.955 182.715 90.475 183.255 ;
        RECT 90.665 182.735 90.995 183.105 ;
        RECT 91.230 183.030 91.400 183.285 ;
        RECT 91.230 182.700 91.515 183.030 ;
        RECT 91.230 182.555 91.400 182.700 ;
        RECT 89.265 181.455 90.475 182.545 ;
        RECT 90.735 182.385 91.400 182.555 ;
        RECT 91.685 182.530 91.855 183.330 ;
        RECT 92.025 183.255 93.235 184.005 ;
        RECT 90.735 181.625 90.905 182.385 ;
        RECT 91.085 181.455 91.415 182.215 ;
        RECT 91.585 181.625 91.855 182.530 ;
        RECT 92.025 182.545 92.545 183.085 ;
        RECT 92.715 182.715 93.235 183.255 ;
        RECT 93.410 183.295 93.665 183.825 ;
        RECT 93.835 183.545 94.140 184.005 ;
        RECT 94.385 183.625 95.455 183.795 ;
        RECT 93.410 182.645 93.620 183.295 ;
        RECT 94.385 183.270 94.705 183.625 ;
        RECT 94.380 183.095 94.705 183.270 ;
        RECT 93.790 182.795 94.705 183.095 ;
        RECT 94.875 183.055 95.115 183.455 ;
        RECT 95.285 183.395 95.455 183.625 ;
        RECT 95.625 183.565 95.815 184.005 ;
        RECT 95.985 183.555 96.935 183.835 ;
        RECT 97.155 183.645 97.505 183.815 ;
        RECT 95.285 183.225 95.815 183.395 ;
        RECT 93.790 182.765 94.530 182.795 ;
        RECT 92.025 181.455 93.235 182.545 ;
        RECT 93.410 181.765 93.665 182.645 ;
        RECT 93.835 181.455 94.140 182.595 ;
        RECT 94.360 182.175 94.530 182.765 ;
        RECT 94.875 182.685 95.415 183.055 ;
        RECT 95.595 182.945 95.815 183.225 ;
        RECT 95.985 182.775 96.155 183.555 ;
        RECT 95.750 182.605 96.155 182.775 ;
        RECT 96.325 182.765 96.675 183.385 ;
        RECT 95.750 182.515 95.920 182.605 ;
        RECT 96.845 182.595 97.055 183.385 ;
        RECT 94.700 182.345 95.920 182.515 ;
        RECT 96.380 182.435 97.055 182.595 ;
        RECT 94.360 182.005 95.160 182.175 ;
        RECT 94.480 181.455 94.810 181.835 ;
        RECT 94.990 181.715 95.160 182.005 ;
        RECT 95.750 181.965 95.920 182.345 ;
        RECT 96.090 182.425 97.055 182.435 ;
        RECT 97.245 183.255 97.505 183.645 ;
        RECT 97.715 183.545 98.045 184.005 ;
        RECT 98.920 183.615 99.775 183.785 ;
        RECT 99.980 183.615 100.475 183.785 ;
        RECT 100.645 183.645 100.975 184.005 ;
        RECT 97.245 182.565 97.415 183.255 ;
        RECT 97.585 182.905 97.755 183.085 ;
        RECT 97.925 183.075 98.715 183.325 ;
        RECT 98.920 182.905 99.090 183.615 ;
        RECT 99.260 183.105 99.615 183.325 ;
        RECT 97.585 182.735 99.275 182.905 ;
        RECT 96.090 182.135 96.550 182.425 ;
        RECT 97.245 182.395 98.745 182.565 ;
        RECT 97.245 182.255 97.415 182.395 ;
        RECT 96.855 182.085 97.415 182.255 ;
        RECT 95.330 181.455 95.580 181.915 ;
        RECT 95.750 181.625 96.620 181.965 ;
        RECT 96.855 181.625 97.025 182.085 ;
        RECT 97.860 182.055 98.935 182.225 ;
        RECT 97.195 181.455 97.565 181.915 ;
        RECT 97.860 181.715 98.030 182.055 ;
        RECT 98.200 181.455 98.530 181.885 ;
        RECT 98.765 181.715 98.935 182.055 ;
        RECT 99.105 181.955 99.275 182.735 ;
        RECT 99.445 182.515 99.615 183.105 ;
        RECT 99.785 182.705 100.135 183.325 ;
        RECT 99.445 182.125 99.910 182.515 ;
        RECT 100.305 182.255 100.475 183.615 ;
        RECT 100.645 182.425 101.105 183.475 ;
        RECT 100.080 182.085 100.475 182.255 ;
        RECT 100.080 181.955 100.250 182.085 ;
        RECT 99.105 181.625 99.785 181.955 ;
        RECT 100.000 181.625 100.250 181.955 ;
        RECT 100.420 181.455 100.670 181.915 ;
        RECT 100.840 181.640 101.165 182.425 ;
        RECT 101.335 181.625 101.505 183.745 ;
        RECT 101.675 183.625 102.005 184.005 ;
        RECT 102.175 183.455 102.430 183.745 ;
        RECT 101.680 183.285 102.430 183.455 ;
        RECT 101.680 182.295 101.910 183.285 ;
        RECT 103.065 183.235 104.735 184.005 ;
        RECT 104.910 183.460 110.255 184.005 ;
        RECT 102.080 182.465 102.430 183.115 ;
        RECT 103.065 182.545 103.815 183.065 ;
        RECT 103.985 182.715 104.735 183.235 ;
        RECT 101.680 182.125 102.430 182.295 ;
        RECT 101.675 181.455 102.005 181.955 ;
        RECT 102.175 181.625 102.430 182.125 ;
        RECT 103.065 181.455 104.735 182.545 ;
        RECT 106.500 181.890 106.850 183.140 ;
        RECT 108.330 182.630 108.670 183.460 ;
        RECT 110.700 183.195 110.945 183.800 ;
        RECT 111.165 183.470 111.675 184.005 ;
        RECT 110.425 183.025 111.655 183.195 ;
        RECT 110.425 182.215 110.765 183.025 ;
        RECT 110.935 182.460 111.685 182.650 ;
        RECT 104.910 181.455 110.255 181.890 ;
        RECT 110.425 181.805 110.940 182.215 ;
        RECT 111.175 181.455 111.345 182.215 ;
        RECT 111.515 181.795 111.685 182.460 ;
        RECT 111.855 182.475 112.045 183.835 ;
        RECT 112.215 182.985 112.490 183.835 ;
        RECT 112.680 183.470 113.210 183.835 ;
        RECT 113.635 183.605 113.965 184.005 ;
        RECT 113.035 183.435 113.210 183.470 ;
        RECT 112.215 182.815 112.495 182.985 ;
        RECT 112.215 182.675 112.490 182.815 ;
        RECT 112.695 182.475 112.865 183.275 ;
        RECT 111.855 182.305 112.865 182.475 ;
        RECT 113.035 183.265 113.965 183.435 ;
        RECT 114.135 183.265 114.390 183.835 ;
        RECT 114.565 183.280 114.855 184.005 ;
        RECT 116.035 183.455 116.205 183.835 ;
        RECT 116.385 183.625 116.715 184.005 ;
        RECT 116.035 183.285 116.700 183.455 ;
        RECT 116.895 183.330 117.155 183.835 ;
        RECT 113.035 182.135 113.205 183.265 ;
        RECT 113.795 183.095 113.965 183.265 ;
        RECT 112.080 181.965 113.205 182.135 ;
        RECT 113.375 182.765 113.570 183.095 ;
        RECT 113.795 182.765 114.050 183.095 ;
        RECT 113.375 181.795 113.545 182.765 ;
        RECT 114.220 182.595 114.390 183.265 ;
        RECT 115.965 182.735 116.295 183.105 ;
        RECT 116.530 183.030 116.700 183.285 ;
        RECT 116.530 182.700 116.815 183.030 ;
        RECT 111.515 181.625 113.545 181.795 ;
        RECT 113.715 181.455 113.885 182.595 ;
        RECT 114.055 181.625 114.390 182.595 ;
        RECT 114.565 181.455 114.855 182.620 ;
        RECT 116.530 182.555 116.700 182.700 ;
        RECT 116.035 182.385 116.700 182.555 ;
        RECT 116.985 182.530 117.155 183.330 ;
        RECT 117.325 183.235 120.835 184.005 ;
        RECT 121.010 183.460 126.355 184.005 ;
        RECT 116.035 181.625 116.205 182.385 ;
        RECT 116.385 181.455 116.715 182.215 ;
        RECT 116.885 181.625 117.155 182.530 ;
        RECT 117.325 182.545 119.015 183.065 ;
        RECT 119.185 182.715 120.835 183.235 ;
        RECT 117.325 181.455 120.835 182.545 ;
        RECT 122.600 181.890 122.950 183.140 ;
        RECT 124.430 182.630 124.770 183.460 ;
        RECT 126.525 183.255 127.735 184.005 ;
        RECT 126.525 182.545 127.045 183.085 ;
        RECT 127.215 182.715 127.735 183.255 ;
        RECT 121.010 181.455 126.355 181.890 ;
        RECT 126.525 181.455 127.735 182.545 ;
        RECT 14.660 181.285 127.820 181.455 ;
        RECT 14.745 180.195 15.955 181.285 ;
        RECT 14.745 179.485 15.265 180.025 ;
        RECT 15.435 179.655 15.955 180.195 ;
        RECT 16.125 180.195 18.715 181.285 ;
        RECT 18.890 180.850 24.235 181.285 ;
        RECT 16.125 179.675 17.335 180.195 ;
        RECT 17.505 179.505 18.715 180.025 ;
        RECT 20.480 179.600 20.830 180.850 ;
        RECT 24.405 180.120 24.695 181.285 ;
        RECT 25.330 180.850 30.675 181.285 ;
        RECT 30.850 180.850 36.195 181.285 ;
        RECT 14.745 178.735 15.955 179.485 ;
        RECT 16.125 178.735 18.715 179.505 ;
        RECT 22.310 179.280 22.650 180.110 ;
        RECT 26.920 179.600 27.270 180.850 ;
        RECT 18.890 178.735 24.235 179.280 ;
        RECT 24.405 178.735 24.695 179.460 ;
        RECT 28.750 179.280 29.090 180.110 ;
        RECT 32.440 179.600 32.790 180.850 ;
        RECT 36.405 180.145 36.635 181.285 ;
        RECT 36.805 180.135 37.135 181.115 ;
        RECT 37.305 180.145 37.515 181.285 ;
        RECT 34.270 179.280 34.610 180.110 ;
        RECT 36.385 179.725 36.715 179.975 ;
        RECT 25.330 178.735 30.675 179.280 ;
        RECT 30.850 178.735 36.195 179.280 ;
        RECT 36.405 178.735 36.635 179.555 ;
        RECT 36.885 179.535 37.135 180.135 ;
        RECT 37.750 180.095 38.005 180.975 ;
        RECT 38.175 180.145 38.480 181.285 ;
        RECT 38.820 180.905 39.150 181.285 ;
        RECT 39.330 180.735 39.500 181.025 ;
        RECT 39.670 180.825 39.920 181.285 ;
        RECT 38.700 180.565 39.500 180.735 ;
        RECT 40.090 180.775 40.960 181.115 ;
        RECT 36.805 178.905 37.135 179.535 ;
        RECT 37.305 178.735 37.515 179.555 ;
        RECT 37.750 179.445 37.960 180.095 ;
        RECT 38.700 179.975 38.870 180.565 ;
        RECT 40.090 180.395 40.260 180.775 ;
        RECT 41.195 180.655 41.365 181.115 ;
        RECT 41.535 180.825 41.905 181.285 ;
        RECT 42.200 180.685 42.370 181.025 ;
        RECT 42.540 180.855 42.870 181.285 ;
        RECT 43.105 180.685 43.275 181.025 ;
        RECT 39.040 180.225 40.260 180.395 ;
        RECT 40.430 180.315 40.890 180.605 ;
        RECT 41.195 180.485 41.755 180.655 ;
        RECT 42.200 180.515 43.275 180.685 ;
        RECT 43.445 180.785 44.125 181.115 ;
        RECT 44.340 180.785 44.590 181.115 ;
        RECT 44.760 180.825 45.010 181.285 ;
        RECT 41.585 180.345 41.755 180.485 ;
        RECT 40.430 180.305 41.395 180.315 ;
        RECT 40.090 180.135 40.260 180.225 ;
        RECT 40.720 180.145 41.395 180.305 ;
        RECT 38.130 179.945 38.870 179.975 ;
        RECT 38.130 179.645 39.045 179.945 ;
        RECT 38.720 179.470 39.045 179.645 ;
        RECT 37.750 178.915 38.005 179.445 ;
        RECT 38.175 178.735 38.480 179.195 ;
        RECT 38.725 179.115 39.045 179.470 ;
        RECT 39.215 179.685 39.755 180.055 ;
        RECT 40.090 179.965 40.495 180.135 ;
        RECT 39.215 179.285 39.455 179.685 ;
        RECT 39.935 179.515 40.155 179.795 ;
        RECT 39.625 179.345 40.155 179.515 ;
        RECT 39.625 179.115 39.795 179.345 ;
        RECT 40.325 179.185 40.495 179.965 ;
        RECT 40.665 179.355 41.015 179.975 ;
        RECT 41.185 179.355 41.395 180.145 ;
        RECT 41.585 180.175 43.085 180.345 ;
        RECT 41.585 179.485 41.755 180.175 ;
        RECT 43.445 180.005 43.615 180.785 ;
        RECT 44.420 180.655 44.590 180.785 ;
        RECT 41.925 179.835 43.615 180.005 ;
        RECT 43.785 180.225 44.250 180.615 ;
        RECT 44.420 180.485 44.815 180.655 ;
        RECT 41.925 179.655 42.095 179.835 ;
        RECT 38.725 178.945 39.795 179.115 ;
        RECT 39.965 178.735 40.155 179.175 ;
        RECT 40.325 178.905 41.275 179.185 ;
        RECT 41.585 179.095 41.845 179.485 ;
        RECT 42.265 179.415 43.055 179.665 ;
        RECT 41.495 178.925 41.845 179.095 ;
        RECT 42.055 178.735 42.385 179.195 ;
        RECT 43.260 179.125 43.430 179.835 ;
        RECT 43.785 179.635 43.955 180.225 ;
        RECT 43.600 179.415 43.955 179.635 ;
        RECT 44.125 179.415 44.475 180.035 ;
        RECT 44.645 179.125 44.815 180.485 ;
        RECT 45.180 180.315 45.505 181.100 ;
        RECT 44.985 179.265 45.445 180.315 ;
        RECT 43.260 178.955 44.115 179.125 ;
        RECT 44.320 178.955 44.815 179.125 ;
        RECT 44.985 178.735 45.315 179.095 ;
        RECT 45.675 178.995 45.845 181.115 ;
        RECT 46.015 180.785 46.345 181.285 ;
        RECT 46.515 180.615 46.770 181.115 ;
        RECT 46.020 180.445 46.770 180.615 ;
        RECT 46.020 179.455 46.250 180.445 ;
        RECT 46.420 179.625 46.770 180.275 ;
        RECT 46.945 180.210 47.215 181.115 ;
        RECT 47.385 180.525 47.715 181.285 ;
        RECT 47.895 180.355 48.065 181.115 ;
        RECT 46.020 179.285 46.770 179.455 ;
        RECT 46.015 178.735 46.345 179.115 ;
        RECT 46.515 178.995 46.770 179.285 ;
        RECT 46.945 179.410 47.115 180.210 ;
        RECT 47.400 180.185 48.065 180.355 ;
        RECT 48.325 180.195 49.995 181.285 ;
        RECT 47.400 180.040 47.570 180.185 ;
        RECT 47.285 179.710 47.570 180.040 ;
        RECT 47.400 179.455 47.570 179.710 ;
        RECT 47.805 179.635 48.135 180.005 ;
        RECT 48.325 179.675 49.075 180.195 ;
        RECT 50.165 180.120 50.455 181.285 ;
        RECT 51.085 180.195 53.675 181.285 ;
        RECT 53.845 180.525 54.360 180.935 ;
        RECT 54.595 180.525 54.765 181.285 ;
        RECT 54.935 180.945 56.965 181.115 ;
        RECT 49.245 179.505 49.995 180.025 ;
        RECT 51.085 179.675 52.295 180.195 ;
        RECT 52.465 179.505 53.675 180.025 ;
        RECT 53.845 179.715 54.185 180.525 ;
        RECT 54.935 180.280 55.105 180.945 ;
        RECT 55.500 180.605 56.625 180.775 ;
        RECT 54.355 180.090 55.105 180.280 ;
        RECT 55.275 180.265 56.285 180.435 ;
        RECT 53.845 179.545 55.075 179.715 ;
        RECT 46.945 178.905 47.205 179.410 ;
        RECT 47.400 179.285 48.065 179.455 ;
        RECT 47.385 178.735 47.715 179.115 ;
        RECT 47.895 178.905 48.065 179.285 ;
        RECT 48.325 178.735 49.995 179.505 ;
        RECT 50.165 178.735 50.455 179.460 ;
        RECT 51.085 178.735 53.675 179.505 ;
        RECT 54.120 178.940 54.365 179.545 ;
        RECT 54.585 178.735 55.095 179.270 ;
        RECT 55.275 178.905 55.465 180.265 ;
        RECT 55.635 179.585 55.910 180.065 ;
        RECT 55.635 179.415 55.915 179.585 ;
        RECT 56.115 179.465 56.285 180.265 ;
        RECT 56.455 179.475 56.625 180.605 ;
        RECT 56.795 179.975 56.965 180.945 ;
        RECT 57.135 180.145 57.305 181.285 ;
        RECT 57.475 180.145 57.810 181.115 ;
        RECT 58.995 180.355 59.165 181.115 ;
        RECT 59.345 180.525 59.675 181.285 ;
        RECT 58.995 180.185 59.660 180.355 ;
        RECT 59.845 180.210 60.115 181.115 ;
        RECT 56.795 179.645 56.990 179.975 ;
        RECT 57.215 179.645 57.470 179.975 ;
        RECT 57.215 179.475 57.385 179.645 ;
        RECT 57.640 179.475 57.810 180.145 ;
        RECT 59.490 180.040 59.660 180.185 ;
        RECT 58.925 179.635 59.255 180.005 ;
        RECT 59.490 179.710 59.775 180.040 ;
        RECT 55.635 178.905 55.910 179.415 ;
        RECT 56.455 179.305 57.385 179.475 ;
        RECT 56.455 179.270 56.630 179.305 ;
        RECT 56.100 178.905 56.630 179.270 ;
        RECT 57.055 178.735 57.385 179.135 ;
        RECT 57.555 178.905 57.810 179.475 ;
        RECT 59.490 179.455 59.660 179.710 ;
        RECT 58.995 179.285 59.660 179.455 ;
        RECT 59.945 179.410 60.115 180.210 ;
        RECT 60.285 180.195 61.955 181.285 ;
        RECT 62.130 180.850 67.475 181.285 ;
        RECT 60.285 179.675 61.035 180.195 ;
        RECT 61.205 179.505 61.955 180.025 ;
        RECT 63.720 179.600 64.070 180.850 ;
        RECT 67.650 180.135 67.910 181.285 ;
        RECT 68.085 180.210 68.340 181.115 ;
        RECT 68.510 180.525 68.840 181.285 ;
        RECT 69.055 180.355 69.225 181.115 ;
        RECT 58.995 178.905 59.165 179.285 ;
        RECT 59.345 178.735 59.675 179.115 ;
        RECT 59.855 178.905 60.115 179.410 ;
        RECT 60.285 178.735 61.955 179.505 ;
        RECT 65.550 179.280 65.890 180.110 ;
        RECT 62.130 178.735 67.475 179.280 ;
        RECT 67.650 178.735 67.910 179.575 ;
        RECT 68.085 179.480 68.255 180.210 ;
        RECT 68.510 180.185 69.225 180.355 ;
        RECT 68.510 179.975 68.680 180.185 ;
        RECT 69.485 180.145 69.745 181.115 ;
        RECT 69.940 180.875 70.270 181.285 ;
        RECT 70.470 180.695 70.640 181.115 ;
        RECT 70.855 180.875 71.525 181.285 ;
        RECT 71.760 180.695 71.930 181.115 ;
        RECT 72.235 180.845 72.565 181.285 ;
        RECT 69.915 180.525 71.930 180.695 ;
        RECT 72.735 180.665 72.910 181.115 ;
        RECT 68.425 179.645 68.680 179.975 ;
        RECT 68.085 178.905 68.340 179.480 ;
        RECT 68.510 179.455 68.680 179.645 ;
        RECT 68.960 179.635 69.315 180.005 ;
        RECT 69.485 179.455 69.655 180.145 ;
        RECT 69.915 179.975 70.085 180.525 ;
        RECT 69.825 179.645 70.085 179.975 ;
        RECT 68.510 179.285 69.225 179.455 ;
        RECT 68.510 178.735 68.840 179.115 ;
        RECT 69.055 178.905 69.225 179.285 ;
        RECT 69.485 178.990 69.825 179.455 ;
        RECT 70.255 179.315 70.595 180.345 ;
        RECT 70.785 179.925 71.055 180.345 ;
        RECT 70.785 179.755 71.095 179.925 ;
        RECT 69.490 178.945 69.825 178.990 ;
        RECT 69.995 178.735 70.325 179.115 ;
        RECT 70.785 179.070 71.055 179.755 ;
        RECT 71.280 179.070 71.560 180.345 ;
        RECT 71.760 179.235 71.930 180.525 ;
        RECT 72.280 180.495 72.910 180.665 ;
        RECT 72.280 179.975 72.450 180.495 ;
        RECT 72.100 179.645 72.450 179.975 ;
        RECT 72.630 179.645 72.995 180.325 ;
        RECT 73.165 180.195 74.375 181.285 ;
        RECT 73.165 179.655 73.685 180.195 ;
        RECT 74.585 180.145 74.815 181.285 ;
        RECT 74.985 180.135 75.315 181.115 ;
        RECT 75.485 180.145 75.695 181.285 ;
        RECT 72.280 179.475 72.450 179.645 ;
        RECT 73.855 179.485 74.375 180.025 ;
        RECT 74.565 179.725 74.895 179.975 ;
        RECT 72.280 179.305 72.910 179.475 ;
        RECT 71.760 178.905 71.990 179.235 ;
        RECT 72.235 178.735 72.565 179.115 ;
        RECT 72.735 178.905 72.910 179.305 ;
        RECT 73.165 178.735 74.375 179.485 ;
        RECT 74.585 178.735 74.815 179.555 ;
        RECT 75.065 179.535 75.315 180.135 ;
        RECT 75.925 180.120 76.215 181.285 ;
        RECT 77.305 180.195 80.815 181.285 ;
        RECT 80.995 180.305 81.325 181.115 ;
        RECT 81.495 180.485 81.735 181.285 ;
        RECT 77.305 179.675 78.995 180.195 ;
        RECT 80.995 180.135 81.710 180.305 ;
        RECT 74.985 178.905 75.315 179.535 ;
        RECT 75.485 178.735 75.695 179.555 ;
        RECT 79.165 179.505 80.815 180.025 ;
        RECT 80.990 179.725 81.370 179.965 ;
        RECT 81.540 179.895 81.710 180.135 ;
        RECT 81.915 180.265 82.085 181.115 ;
        RECT 82.255 180.485 82.585 181.285 ;
        RECT 82.755 180.265 82.925 181.115 ;
        RECT 81.915 180.095 82.925 180.265 ;
        RECT 83.095 180.135 83.425 181.285 ;
        RECT 81.540 179.725 82.040 179.895 ;
        RECT 81.540 179.555 81.710 179.725 ;
        RECT 82.430 179.585 82.925 180.095 ;
        RECT 82.425 179.555 82.925 179.585 ;
        RECT 75.925 178.735 76.215 179.460 ;
        RECT 77.305 178.735 80.815 179.505 ;
        RECT 81.075 179.385 81.710 179.555 ;
        RECT 81.915 179.385 82.925 179.555 ;
        RECT 84.670 180.095 84.925 180.975 ;
        RECT 85.095 180.145 85.400 181.285 ;
        RECT 85.740 180.905 86.070 181.285 ;
        RECT 86.250 180.735 86.420 181.025 ;
        RECT 86.590 180.825 86.840 181.285 ;
        RECT 85.620 180.565 86.420 180.735 ;
        RECT 87.010 180.775 87.880 181.115 ;
        RECT 81.075 178.905 81.245 179.385 ;
        RECT 81.425 178.735 81.665 179.215 ;
        RECT 81.915 178.905 82.085 179.385 ;
        RECT 82.255 178.735 82.585 179.215 ;
        RECT 82.755 178.905 82.925 179.385 ;
        RECT 83.095 178.735 83.425 179.535 ;
        RECT 84.670 179.445 84.880 180.095 ;
        RECT 85.620 179.975 85.790 180.565 ;
        RECT 87.010 180.395 87.180 180.775 ;
        RECT 88.115 180.655 88.285 181.115 ;
        RECT 88.455 180.825 88.825 181.285 ;
        RECT 89.120 180.685 89.290 181.025 ;
        RECT 89.460 180.855 89.790 181.285 ;
        RECT 90.025 180.685 90.195 181.025 ;
        RECT 85.960 180.225 87.180 180.395 ;
        RECT 87.350 180.315 87.810 180.605 ;
        RECT 88.115 180.485 88.675 180.655 ;
        RECT 89.120 180.515 90.195 180.685 ;
        RECT 90.365 180.785 91.045 181.115 ;
        RECT 91.260 180.785 91.510 181.115 ;
        RECT 91.680 180.825 91.930 181.285 ;
        RECT 88.505 180.345 88.675 180.485 ;
        RECT 87.350 180.305 88.315 180.315 ;
        RECT 87.010 180.135 87.180 180.225 ;
        RECT 87.640 180.145 88.315 180.305 ;
        RECT 85.050 179.945 85.790 179.975 ;
        RECT 85.050 179.645 85.965 179.945 ;
        RECT 85.640 179.470 85.965 179.645 ;
        RECT 84.670 178.915 84.925 179.445 ;
        RECT 85.095 178.735 85.400 179.195 ;
        RECT 85.645 179.115 85.965 179.470 ;
        RECT 86.135 179.685 86.675 180.055 ;
        RECT 87.010 179.965 87.415 180.135 ;
        RECT 86.135 179.285 86.375 179.685 ;
        RECT 86.855 179.515 87.075 179.795 ;
        RECT 86.545 179.345 87.075 179.515 ;
        RECT 86.545 179.115 86.715 179.345 ;
        RECT 87.245 179.185 87.415 179.965 ;
        RECT 87.585 179.355 87.935 179.975 ;
        RECT 88.105 179.355 88.315 180.145 ;
        RECT 88.505 180.175 90.005 180.345 ;
        RECT 88.505 179.485 88.675 180.175 ;
        RECT 90.365 180.005 90.535 180.785 ;
        RECT 91.340 180.655 91.510 180.785 ;
        RECT 88.845 179.835 90.535 180.005 ;
        RECT 90.705 180.225 91.170 180.615 ;
        RECT 91.340 180.485 91.735 180.655 ;
        RECT 88.845 179.655 89.015 179.835 ;
        RECT 85.645 178.945 86.715 179.115 ;
        RECT 86.885 178.735 87.075 179.175 ;
        RECT 87.245 178.905 88.195 179.185 ;
        RECT 88.505 179.095 88.765 179.485 ;
        RECT 89.185 179.415 89.975 179.665 ;
        RECT 88.415 178.925 88.765 179.095 ;
        RECT 88.975 178.735 89.305 179.195 ;
        RECT 90.180 179.125 90.350 179.835 ;
        RECT 90.705 179.635 90.875 180.225 ;
        RECT 90.520 179.415 90.875 179.635 ;
        RECT 91.045 179.415 91.395 180.035 ;
        RECT 91.565 179.125 91.735 180.485 ;
        RECT 92.100 180.315 92.425 181.100 ;
        RECT 91.905 179.265 92.365 180.315 ;
        RECT 90.180 178.955 91.035 179.125 ;
        RECT 91.240 178.955 91.735 179.125 ;
        RECT 91.905 178.735 92.235 179.095 ;
        RECT 92.595 178.995 92.765 181.115 ;
        RECT 92.935 180.785 93.265 181.285 ;
        RECT 93.435 180.615 93.690 181.115 ;
        RECT 92.940 180.445 93.690 180.615 ;
        RECT 92.940 179.455 93.170 180.445 ;
        RECT 93.340 179.625 93.690 180.275 ;
        RECT 94.825 180.145 95.055 181.285 ;
        RECT 95.225 180.135 95.555 181.115 ;
        RECT 95.725 180.145 95.935 181.285 ;
        RECT 96.165 180.525 96.680 180.935 ;
        RECT 96.915 180.525 97.085 181.285 ;
        RECT 97.255 180.945 99.285 181.115 ;
        RECT 94.805 179.725 95.135 179.975 ;
        RECT 92.940 179.285 93.690 179.455 ;
        RECT 92.935 178.735 93.265 179.115 ;
        RECT 93.435 178.995 93.690 179.285 ;
        RECT 94.825 178.735 95.055 179.555 ;
        RECT 95.305 179.535 95.555 180.135 ;
        RECT 96.165 179.715 96.505 180.525 ;
        RECT 97.255 180.280 97.425 180.945 ;
        RECT 97.820 180.605 98.945 180.775 ;
        RECT 96.675 180.090 97.425 180.280 ;
        RECT 97.595 180.265 98.605 180.435 ;
        RECT 95.225 178.905 95.555 179.535 ;
        RECT 95.725 178.735 95.935 179.555 ;
        RECT 96.165 179.545 97.395 179.715 ;
        RECT 96.440 178.940 96.685 179.545 ;
        RECT 96.905 178.735 97.415 179.270 ;
        RECT 97.595 178.905 97.785 180.265 ;
        RECT 97.955 179.925 98.230 180.065 ;
        RECT 97.955 179.755 98.235 179.925 ;
        RECT 97.955 178.905 98.230 179.755 ;
        RECT 98.435 179.465 98.605 180.265 ;
        RECT 98.775 179.475 98.945 180.605 ;
        RECT 99.115 179.975 99.285 180.945 ;
        RECT 99.455 180.145 99.625 181.285 ;
        RECT 99.795 180.145 100.130 181.115 ;
        RECT 100.395 180.355 100.565 181.115 ;
        RECT 100.745 180.525 101.075 181.285 ;
        RECT 100.395 180.185 101.060 180.355 ;
        RECT 101.245 180.210 101.515 181.115 ;
        RECT 99.115 179.645 99.310 179.975 ;
        RECT 99.535 179.645 99.790 179.975 ;
        RECT 99.535 179.475 99.705 179.645 ;
        RECT 99.960 179.475 100.130 180.145 ;
        RECT 100.890 180.040 101.060 180.185 ;
        RECT 100.325 179.635 100.655 180.005 ;
        RECT 100.890 179.710 101.175 180.040 ;
        RECT 98.775 179.305 99.705 179.475 ;
        RECT 98.775 179.270 98.950 179.305 ;
        RECT 98.420 178.905 98.950 179.270 ;
        RECT 99.375 178.735 99.705 179.135 ;
        RECT 99.875 178.905 100.130 179.475 ;
        RECT 100.890 179.455 101.060 179.710 ;
        RECT 100.395 179.285 101.060 179.455 ;
        RECT 101.345 179.410 101.515 180.210 ;
        RECT 101.685 180.120 101.975 181.285 ;
        RECT 102.145 180.195 103.355 181.285 ;
        RECT 103.525 180.195 107.035 181.285 ;
        RECT 102.145 179.655 102.665 180.195 ;
        RECT 102.835 179.485 103.355 180.025 ;
        RECT 103.525 179.675 105.215 180.195 ;
        RECT 107.205 180.145 107.545 181.115 ;
        RECT 107.715 180.145 107.885 181.285 ;
        RECT 108.155 180.485 108.405 181.285 ;
        RECT 109.050 180.315 109.380 181.115 ;
        RECT 109.680 180.485 110.010 181.285 ;
        RECT 110.180 180.315 110.510 181.115 ;
        RECT 108.075 180.145 110.510 180.315 ;
        RECT 110.885 180.195 112.095 181.285 ;
        RECT 112.265 180.525 112.780 180.935 ;
        RECT 113.015 180.525 113.185 181.285 ;
        RECT 113.355 180.945 115.385 181.115 ;
        RECT 105.385 179.505 107.035 180.025 ;
        RECT 100.395 178.905 100.565 179.285 ;
        RECT 100.745 178.735 101.075 179.115 ;
        RECT 101.255 178.905 101.515 179.410 ;
        RECT 101.685 178.735 101.975 179.460 ;
        RECT 102.145 178.735 103.355 179.485 ;
        RECT 103.525 178.735 107.035 179.505 ;
        RECT 107.205 179.535 107.380 180.145 ;
        RECT 108.075 179.895 108.245 180.145 ;
        RECT 107.550 179.725 108.245 179.895 ;
        RECT 108.420 179.725 108.840 179.925 ;
        RECT 109.010 179.725 109.340 179.925 ;
        RECT 109.510 179.725 109.840 179.925 ;
        RECT 107.205 178.905 107.545 179.535 ;
        RECT 107.715 178.735 107.965 179.535 ;
        RECT 108.155 179.385 109.380 179.555 ;
        RECT 108.155 178.905 108.485 179.385 ;
        RECT 108.655 178.735 108.880 179.195 ;
        RECT 109.050 178.905 109.380 179.385 ;
        RECT 110.010 179.515 110.180 180.145 ;
        RECT 110.365 179.725 110.715 179.975 ;
        RECT 110.885 179.655 111.405 180.195 ;
        RECT 110.010 178.905 110.510 179.515 ;
        RECT 111.575 179.485 112.095 180.025 ;
        RECT 112.265 179.715 112.605 180.525 ;
        RECT 113.355 180.280 113.525 180.945 ;
        RECT 113.920 180.605 115.045 180.775 ;
        RECT 112.775 180.090 113.525 180.280 ;
        RECT 113.695 180.265 114.705 180.435 ;
        RECT 112.265 179.545 113.495 179.715 ;
        RECT 110.885 178.735 112.095 179.485 ;
        RECT 112.540 178.940 112.785 179.545 ;
        RECT 113.005 178.735 113.515 179.270 ;
        RECT 113.695 178.905 113.885 180.265 ;
        RECT 114.055 179.925 114.330 180.065 ;
        RECT 114.055 179.755 114.335 179.925 ;
        RECT 114.055 178.905 114.330 179.755 ;
        RECT 114.535 179.465 114.705 180.265 ;
        RECT 114.875 179.475 115.045 180.605 ;
        RECT 115.215 179.975 115.385 180.945 ;
        RECT 115.555 180.145 115.725 181.285 ;
        RECT 115.895 180.145 116.230 181.115 ;
        RECT 115.215 179.645 115.410 179.975 ;
        RECT 115.635 179.645 115.890 179.975 ;
        RECT 115.635 179.475 115.805 179.645 ;
        RECT 116.060 179.475 116.230 180.145 ;
        RECT 116.405 180.195 118.075 181.285 ;
        RECT 116.405 179.675 117.155 180.195 ;
        RECT 118.305 180.145 118.515 181.285 ;
        RECT 118.685 180.135 119.015 181.115 ;
        RECT 119.185 180.145 119.415 181.285 ;
        RECT 119.625 180.195 120.835 181.285 ;
        RECT 121.010 180.850 126.355 181.285 ;
        RECT 117.325 179.505 118.075 180.025 ;
        RECT 114.875 179.305 115.805 179.475 ;
        RECT 114.875 179.270 115.050 179.305 ;
        RECT 114.520 178.905 115.050 179.270 ;
        RECT 115.475 178.735 115.805 179.135 ;
        RECT 115.975 178.905 116.230 179.475 ;
        RECT 116.405 178.735 118.075 179.505 ;
        RECT 118.305 178.735 118.515 179.555 ;
        RECT 118.685 179.535 118.935 180.135 ;
        RECT 119.105 179.725 119.435 179.975 ;
        RECT 119.625 179.655 120.145 180.195 ;
        RECT 118.685 178.905 119.015 179.535 ;
        RECT 119.185 178.735 119.415 179.555 ;
        RECT 120.315 179.485 120.835 180.025 ;
        RECT 122.600 179.600 122.950 180.850 ;
        RECT 126.525 180.195 127.735 181.285 ;
        RECT 119.625 178.735 120.835 179.485 ;
        RECT 124.430 179.280 124.770 180.110 ;
        RECT 126.525 179.655 127.045 180.195 ;
        RECT 127.215 179.485 127.735 180.025 ;
        RECT 121.010 178.735 126.355 179.280 ;
        RECT 126.525 178.735 127.735 179.485 ;
        RECT 14.660 178.565 127.820 178.735 ;
        RECT 14.745 177.815 15.955 178.565 ;
        RECT 17.050 178.020 22.395 178.565 ;
        RECT 14.745 177.275 15.265 177.815 ;
        RECT 15.435 177.105 15.955 177.645 ;
        RECT 14.745 176.015 15.955 177.105 ;
        RECT 18.640 176.450 18.990 177.700 ;
        RECT 20.470 177.190 20.810 178.020 ;
        RECT 22.570 178.015 22.825 178.305 ;
        RECT 22.995 178.185 23.325 178.565 ;
        RECT 22.570 177.845 23.320 178.015 ;
        RECT 22.570 177.025 22.920 177.675 ;
        RECT 23.090 176.855 23.320 177.845 ;
        RECT 22.570 176.685 23.320 176.855 ;
        RECT 17.050 176.015 22.395 176.450 ;
        RECT 22.570 176.185 22.825 176.685 ;
        RECT 22.995 176.015 23.325 176.515 ;
        RECT 23.495 176.185 23.665 178.305 ;
        RECT 24.025 178.205 24.355 178.565 ;
        RECT 24.525 178.175 25.020 178.345 ;
        RECT 25.225 178.175 26.080 178.345 ;
        RECT 23.895 176.985 24.355 178.035 ;
        RECT 23.835 176.200 24.160 176.985 ;
        RECT 24.525 176.815 24.695 178.175 ;
        RECT 24.865 177.265 25.215 177.885 ;
        RECT 25.385 177.665 25.740 177.885 ;
        RECT 25.385 177.075 25.555 177.665 ;
        RECT 25.910 177.465 26.080 178.175 ;
        RECT 26.955 178.105 27.285 178.565 ;
        RECT 27.495 178.205 27.845 178.375 ;
        RECT 26.285 177.635 27.075 177.885 ;
        RECT 27.495 177.815 27.755 178.205 ;
        RECT 28.065 178.115 29.015 178.395 ;
        RECT 29.185 178.125 29.375 178.565 ;
        RECT 29.545 178.185 30.615 178.355 ;
        RECT 27.245 177.465 27.415 177.645 ;
        RECT 24.525 176.645 24.920 176.815 ;
        RECT 25.090 176.685 25.555 177.075 ;
        RECT 25.725 177.295 27.415 177.465 ;
        RECT 24.750 176.515 24.920 176.645 ;
        RECT 25.725 176.515 25.895 177.295 ;
        RECT 27.585 177.125 27.755 177.815 ;
        RECT 26.255 176.955 27.755 177.125 ;
        RECT 27.945 177.155 28.155 177.945 ;
        RECT 28.325 177.325 28.675 177.945 ;
        RECT 28.845 177.335 29.015 178.115 ;
        RECT 29.545 177.955 29.715 178.185 ;
        RECT 29.185 177.785 29.715 177.955 ;
        RECT 29.185 177.505 29.405 177.785 ;
        RECT 29.885 177.615 30.125 178.015 ;
        RECT 28.845 177.165 29.250 177.335 ;
        RECT 29.585 177.245 30.125 177.615 ;
        RECT 30.295 177.830 30.615 178.185 ;
        RECT 30.860 178.105 31.165 178.565 ;
        RECT 31.335 177.855 31.590 178.385 ;
        RECT 30.295 177.655 30.620 177.830 ;
        RECT 30.295 177.355 31.210 177.655 ;
        RECT 30.470 177.325 31.210 177.355 ;
        RECT 27.945 176.995 28.620 177.155 ;
        RECT 29.080 177.075 29.250 177.165 ;
        RECT 27.945 176.985 28.910 176.995 ;
        RECT 27.585 176.815 27.755 176.955 ;
        RECT 24.330 176.015 24.580 176.475 ;
        RECT 24.750 176.185 25.000 176.515 ;
        RECT 25.215 176.185 25.895 176.515 ;
        RECT 26.065 176.615 27.140 176.785 ;
        RECT 27.585 176.645 28.145 176.815 ;
        RECT 28.450 176.695 28.910 176.985 ;
        RECT 29.080 176.905 30.300 177.075 ;
        RECT 26.065 176.275 26.235 176.615 ;
        RECT 26.470 176.015 26.800 176.445 ;
        RECT 26.970 176.275 27.140 176.615 ;
        RECT 27.435 176.015 27.805 176.475 ;
        RECT 27.975 176.185 28.145 176.645 ;
        RECT 29.080 176.525 29.250 176.905 ;
        RECT 30.470 176.735 30.640 177.325 ;
        RECT 31.380 177.205 31.590 177.855 ;
        RECT 28.380 176.185 29.250 176.525 ;
        RECT 29.840 176.565 30.640 176.735 ;
        RECT 29.420 176.015 29.670 176.475 ;
        RECT 29.840 176.275 30.010 176.565 ;
        RECT 30.190 176.015 30.520 176.395 ;
        RECT 30.860 176.015 31.165 177.155 ;
        RECT 31.335 176.325 31.590 177.205 ;
        RECT 32.225 177.890 32.485 178.395 ;
        RECT 32.665 178.185 32.995 178.565 ;
        RECT 33.175 178.015 33.345 178.395 ;
        RECT 32.225 177.090 32.395 177.890 ;
        RECT 32.680 177.845 33.345 178.015 ;
        RECT 32.680 177.590 32.850 177.845 ;
        RECT 33.810 177.785 34.310 178.395 ;
        RECT 32.565 177.260 32.850 177.590 ;
        RECT 33.085 177.295 33.415 177.665 ;
        RECT 33.605 177.325 33.955 177.575 ;
        RECT 32.680 177.115 32.850 177.260 ;
        RECT 34.140 177.155 34.310 177.785 ;
        RECT 34.940 177.915 35.270 178.395 ;
        RECT 35.440 178.105 35.665 178.565 ;
        RECT 35.835 177.915 36.165 178.395 ;
        RECT 34.940 177.745 36.165 177.915 ;
        RECT 36.355 177.765 36.605 178.565 ;
        RECT 36.775 177.765 37.115 178.395 ;
        RECT 37.285 177.840 37.575 178.565 ;
        RECT 38.205 177.795 41.715 178.565 ;
        RECT 34.480 177.375 34.810 177.575 ;
        RECT 34.980 177.375 35.310 177.575 ;
        RECT 35.480 177.375 35.900 177.575 ;
        RECT 36.075 177.405 36.770 177.575 ;
        RECT 36.075 177.155 36.245 177.405 ;
        RECT 36.940 177.155 37.115 177.765 ;
        RECT 32.225 176.185 32.495 177.090 ;
        RECT 32.680 176.945 33.345 177.115 ;
        RECT 32.665 176.015 32.995 176.775 ;
        RECT 33.175 176.185 33.345 176.945 ;
        RECT 33.810 176.985 36.245 177.155 ;
        RECT 33.810 176.185 34.140 176.985 ;
        RECT 34.310 176.015 34.640 176.815 ;
        RECT 34.940 176.185 35.270 176.985 ;
        RECT 35.915 176.015 36.165 176.815 ;
        RECT 36.435 176.015 36.605 177.155 ;
        RECT 36.775 176.185 37.115 177.155 ;
        RECT 37.285 176.015 37.575 177.180 ;
        RECT 38.205 177.105 39.895 177.625 ;
        RECT 40.065 177.275 41.715 177.795 ;
        RECT 42.090 177.785 42.590 178.395 ;
        RECT 41.885 177.325 42.235 177.575 ;
        RECT 42.420 177.155 42.590 177.785 ;
        RECT 43.220 177.915 43.550 178.395 ;
        RECT 43.720 178.105 43.945 178.565 ;
        RECT 44.115 177.915 44.445 178.395 ;
        RECT 43.220 177.745 44.445 177.915 ;
        RECT 44.635 177.765 44.885 178.565 ;
        RECT 45.055 177.765 45.395 178.395 ;
        RECT 45.565 178.055 45.870 178.565 ;
        RECT 42.760 177.375 43.090 177.575 ;
        RECT 43.260 177.375 43.590 177.575 ;
        RECT 43.760 177.375 44.180 177.575 ;
        RECT 44.355 177.405 45.050 177.575 ;
        RECT 44.355 177.155 44.525 177.405 ;
        RECT 45.220 177.155 45.395 177.765 ;
        RECT 45.565 177.325 45.880 177.885 ;
        RECT 46.050 177.575 46.300 178.385 ;
        RECT 46.470 178.040 46.730 178.565 ;
        RECT 46.910 177.575 47.160 178.385 ;
        RECT 47.330 178.005 47.590 178.565 ;
        RECT 47.760 177.915 48.020 178.370 ;
        RECT 48.190 178.085 48.450 178.565 ;
        RECT 48.620 177.915 48.880 178.370 ;
        RECT 49.050 178.085 49.310 178.565 ;
        RECT 49.480 177.915 49.740 178.370 ;
        RECT 49.910 178.085 50.155 178.565 ;
        RECT 50.325 177.915 50.600 178.370 ;
        RECT 50.770 178.085 51.015 178.565 ;
        RECT 51.185 177.915 51.445 178.370 ;
        RECT 51.625 178.085 51.875 178.565 ;
        RECT 52.045 177.915 52.305 178.370 ;
        RECT 52.485 178.085 52.735 178.565 ;
        RECT 52.905 177.915 53.165 178.370 ;
        RECT 53.345 178.085 53.605 178.565 ;
        RECT 53.775 177.915 54.035 178.370 ;
        RECT 54.205 178.085 54.505 178.565 ;
        RECT 47.760 177.885 54.505 177.915 ;
        RECT 47.760 177.745 54.535 177.885 ;
        RECT 54.765 177.795 57.355 178.565 ;
        RECT 57.530 178.020 62.875 178.565 ;
        RECT 53.340 177.715 54.535 177.745 ;
        RECT 46.050 177.325 53.170 177.575 ;
        RECT 38.205 176.015 41.715 177.105 ;
        RECT 42.090 176.985 44.525 177.155 ;
        RECT 42.090 176.185 42.420 176.985 ;
        RECT 42.590 176.015 42.920 176.815 ;
        RECT 43.220 176.185 43.550 176.985 ;
        RECT 44.195 176.015 44.445 176.815 ;
        RECT 44.715 176.015 44.885 177.155 ;
        RECT 45.055 176.185 45.395 177.155 ;
        RECT 45.575 176.015 45.870 176.825 ;
        RECT 46.050 176.185 46.295 177.325 ;
        RECT 46.470 176.015 46.730 176.825 ;
        RECT 46.910 176.190 47.160 177.325 ;
        RECT 53.340 177.155 54.505 177.715 ;
        RECT 47.760 176.930 54.505 177.155 ;
        RECT 54.765 177.105 55.975 177.625 ;
        RECT 56.145 177.275 57.355 177.795 ;
        RECT 47.760 176.915 53.165 176.930 ;
        RECT 47.330 176.020 47.590 176.815 ;
        RECT 47.760 176.190 48.020 176.915 ;
        RECT 48.190 176.020 48.450 176.745 ;
        RECT 48.620 176.190 48.880 176.915 ;
        RECT 49.050 176.020 49.310 176.745 ;
        RECT 49.480 176.190 49.740 176.915 ;
        RECT 49.910 176.020 50.170 176.745 ;
        RECT 50.340 176.190 50.600 176.915 ;
        RECT 50.770 176.020 51.015 176.745 ;
        RECT 51.185 176.190 51.445 176.915 ;
        RECT 51.630 176.020 51.875 176.745 ;
        RECT 52.045 176.190 52.305 176.915 ;
        RECT 52.490 176.020 52.735 176.745 ;
        RECT 52.905 176.190 53.165 176.915 ;
        RECT 53.350 176.020 53.605 176.745 ;
        RECT 53.775 176.190 54.065 176.930 ;
        RECT 47.330 176.015 53.605 176.020 ;
        RECT 54.235 176.015 54.505 176.760 ;
        RECT 54.765 176.015 57.355 177.105 ;
        RECT 59.120 176.450 59.470 177.700 ;
        RECT 60.950 177.190 61.290 178.020 ;
        RECT 63.045 177.840 63.335 178.565 ;
        RECT 63.510 177.725 63.770 178.565 ;
        RECT 63.945 177.820 64.200 178.395 ;
        RECT 64.370 178.185 64.700 178.565 ;
        RECT 64.915 178.015 65.085 178.395 ;
        RECT 64.370 177.845 65.085 178.015 ;
        RECT 65.435 178.015 65.605 178.395 ;
        RECT 65.820 178.185 66.150 178.565 ;
        RECT 65.435 177.845 66.150 178.015 ;
        RECT 57.530 176.015 62.875 176.450 ;
        RECT 63.045 176.015 63.335 177.180 ;
        RECT 63.510 176.015 63.770 177.165 ;
        RECT 63.945 177.090 64.115 177.820 ;
        RECT 64.370 177.655 64.540 177.845 ;
        RECT 64.285 177.325 64.540 177.655 ;
        RECT 64.370 177.115 64.540 177.325 ;
        RECT 64.820 177.295 65.175 177.665 ;
        RECT 65.345 177.295 65.700 177.665 ;
        RECT 65.980 177.655 66.150 177.845 ;
        RECT 66.320 177.820 66.575 178.395 ;
        RECT 65.980 177.325 66.235 177.655 ;
        RECT 65.980 177.115 66.150 177.325 ;
        RECT 63.945 176.185 64.200 177.090 ;
        RECT 64.370 176.945 65.085 177.115 ;
        RECT 64.370 176.015 64.700 176.775 ;
        RECT 64.915 176.185 65.085 176.945 ;
        RECT 65.435 176.945 66.150 177.115 ;
        RECT 66.405 177.090 66.575 177.820 ;
        RECT 66.750 177.725 67.010 178.565 ;
        RECT 67.185 177.795 68.855 178.565 ;
        RECT 69.030 178.020 74.375 178.565 ;
        RECT 74.545 178.065 74.845 178.395 ;
        RECT 75.015 178.085 75.290 178.565 ;
        RECT 65.435 176.185 65.605 176.945 ;
        RECT 65.820 176.015 66.150 176.775 ;
        RECT 66.320 176.185 66.575 177.090 ;
        RECT 66.750 176.015 67.010 177.165 ;
        RECT 67.185 177.105 67.935 177.625 ;
        RECT 68.105 177.275 68.855 177.795 ;
        RECT 67.185 176.015 68.855 177.105 ;
        RECT 70.620 176.450 70.970 177.700 ;
        RECT 72.450 177.190 72.790 178.020 ;
        RECT 74.545 177.155 74.715 178.065 ;
        RECT 75.470 177.915 75.765 178.305 ;
        RECT 75.935 178.085 76.190 178.565 ;
        RECT 76.365 177.915 76.625 178.305 ;
        RECT 76.795 178.085 77.075 178.565 ;
        RECT 74.885 177.325 75.235 177.895 ;
        RECT 75.470 177.745 77.120 177.915 ;
        RECT 77.510 177.785 78.010 178.395 ;
        RECT 75.405 177.405 76.545 177.575 ;
        RECT 75.405 177.155 75.575 177.405 ;
        RECT 76.715 177.235 77.120 177.745 ;
        RECT 77.305 177.325 77.655 177.575 ;
        RECT 74.545 176.985 75.575 177.155 ;
        RECT 76.365 177.065 77.120 177.235 ;
        RECT 77.840 177.155 78.010 177.785 ;
        RECT 78.640 177.915 78.970 178.395 ;
        RECT 79.140 178.105 79.365 178.565 ;
        RECT 79.535 177.915 79.865 178.395 ;
        RECT 78.640 177.745 79.865 177.915 ;
        RECT 80.055 177.765 80.305 178.565 ;
        RECT 80.475 177.765 80.815 178.395 ;
        RECT 78.180 177.375 78.510 177.575 ;
        RECT 78.680 177.375 79.010 177.575 ;
        RECT 79.180 177.375 79.600 177.575 ;
        RECT 79.775 177.405 80.470 177.575 ;
        RECT 79.775 177.155 79.945 177.405 ;
        RECT 80.640 177.155 80.815 177.765 ;
        RECT 69.030 176.015 74.375 176.450 ;
        RECT 74.545 176.185 74.855 176.985 ;
        RECT 76.365 176.815 76.625 177.065 ;
        RECT 77.510 176.985 79.945 177.155 ;
        RECT 75.025 176.015 75.335 176.815 ;
        RECT 75.505 176.645 76.625 176.815 ;
        RECT 75.505 176.185 75.765 176.645 ;
        RECT 75.935 176.015 76.190 176.475 ;
        RECT 76.365 176.185 76.625 176.645 ;
        RECT 76.795 176.015 77.080 176.885 ;
        RECT 77.510 176.185 77.840 176.985 ;
        RECT 78.010 176.015 78.340 176.815 ;
        RECT 78.640 176.185 78.970 176.985 ;
        RECT 79.615 176.015 79.865 176.815 ;
        RECT 80.135 176.015 80.305 177.155 ;
        RECT 80.475 176.185 80.815 177.155 ;
        RECT 80.985 177.765 81.325 178.395 ;
        RECT 81.495 177.765 81.745 178.565 ;
        RECT 81.935 177.915 82.265 178.395 ;
        RECT 82.435 178.105 82.660 178.565 ;
        RECT 82.830 177.915 83.160 178.395 ;
        RECT 80.985 177.155 81.160 177.765 ;
        RECT 81.935 177.745 83.160 177.915 ;
        RECT 83.790 177.785 84.290 178.395 ;
        RECT 84.755 177.915 84.925 178.395 ;
        RECT 85.105 178.085 85.345 178.565 ;
        RECT 85.595 177.915 85.765 178.395 ;
        RECT 85.935 178.085 86.265 178.565 ;
        RECT 86.435 177.915 86.605 178.395 ;
        RECT 81.330 177.405 82.025 177.575 ;
        RECT 81.855 177.155 82.025 177.405 ;
        RECT 82.200 177.375 82.620 177.575 ;
        RECT 82.790 177.375 83.120 177.575 ;
        RECT 83.290 177.375 83.620 177.575 ;
        RECT 83.790 177.155 83.960 177.785 ;
        RECT 84.755 177.745 85.390 177.915 ;
        RECT 85.595 177.745 86.605 177.915 ;
        RECT 86.775 177.765 87.105 178.565 ;
        RECT 87.485 177.745 87.695 178.565 ;
        RECT 87.865 177.765 88.195 178.395 ;
        RECT 85.220 177.575 85.390 177.745 ;
        RECT 84.145 177.325 84.495 177.575 ;
        RECT 84.670 177.335 85.050 177.575 ;
        RECT 85.220 177.405 85.720 177.575 ;
        RECT 86.110 177.545 86.605 177.745 ;
        RECT 85.220 177.165 85.390 177.405 ;
        RECT 86.105 177.375 86.605 177.545 ;
        RECT 86.110 177.205 86.605 177.375 ;
        RECT 80.985 176.185 81.325 177.155 ;
        RECT 81.495 176.015 81.665 177.155 ;
        RECT 81.855 176.985 84.290 177.155 ;
        RECT 81.935 176.015 82.185 176.815 ;
        RECT 82.830 176.185 83.160 176.985 ;
        RECT 83.460 176.015 83.790 176.815 ;
        RECT 83.960 176.185 84.290 176.985 ;
        RECT 84.675 176.995 85.390 177.165 ;
        RECT 85.595 177.035 86.605 177.205 ;
        RECT 87.865 177.165 88.115 177.765 ;
        RECT 88.365 177.745 88.595 178.565 ;
        RECT 88.805 177.840 89.095 178.565 ;
        RECT 89.270 178.020 94.615 178.565 ;
        RECT 94.790 178.020 100.135 178.565 ;
        RECT 88.285 177.325 88.615 177.575 ;
        RECT 84.675 176.185 85.005 176.995 ;
        RECT 85.175 176.015 85.415 176.815 ;
        RECT 85.595 176.185 85.765 177.035 ;
        RECT 85.935 176.015 86.265 176.815 ;
        RECT 86.435 176.185 86.605 177.035 ;
        RECT 86.775 176.015 87.105 177.165 ;
        RECT 87.485 176.015 87.695 177.155 ;
        RECT 87.865 176.185 88.195 177.165 ;
        RECT 88.365 176.015 88.595 177.155 ;
        RECT 88.805 176.015 89.095 177.180 ;
        RECT 90.860 176.450 91.210 177.700 ;
        RECT 92.690 177.190 93.030 178.020 ;
        RECT 96.380 176.450 96.730 177.700 ;
        RECT 98.210 177.190 98.550 178.020 ;
        RECT 100.510 177.785 101.010 178.395 ;
        RECT 100.305 177.325 100.655 177.575 ;
        RECT 100.840 177.155 101.010 177.785 ;
        RECT 101.640 177.915 101.970 178.395 ;
        RECT 102.140 178.105 102.365 178.565 ;
        RECT 102.535 177.915 102.865 178.395 ;
        RECT 101.640 177.745 102.865 177.915 ;
        RECT 103.055 177.765 103.305 178.565 ;
        RECT 103.475 177.765 103.815 178.395 ;
        RECT 101.180 177.375 101.510 177.575 ;
        RECT 101.680 177.375 102.010 177.575 ;
        RECT 102.180 177.375 102.600 177.575 ;
        RECT 102.775 177.405 103.470 177.575 ;
        RECT 102.775 177.155 102.945 177.405 ;
        RECT 103.640 177.155 103.815 177.765 ;
        RECT 100.510 176.985 102.945 177.155 ;
        RECT 89.270 176.015 94.615 176.450 ;
        RECT 94.790 176.015 100.135 176.450 ;
        RECT 100.510 176.185 100.840 176.985 ;
        RECT 101.010 176.015 101.340 176.815 ;
        RECT 101.640 176.185 101.970 176.985 ;
        RECT 102.615 176.015 102.865 176.815 ;
        RECT 103.135 176.015 103.305 177.155 ;
        RECT 103.475 176.185 103.815 177.155 ;
        RECT 103.985 177.765 104.325 178.395 ;
        RECT 104.495 177.765 104.745 178.565 ;
        RECT 104.935 177.915 105.265 178.395 ;
        RECT 105.435 178.105 105.660 178.565 ;
        RECT 105.830 177.915 106.160 178.395 ;
        RECT 103.985 177.155 104.160 177.765 ;
        RECT 104.935 177.745 106.160 177.915 ;
        RECT 106.790 177.785 107.290 178.395 ;
        RECT 104.330 177.405 105.025 177.575 ;
        RECT 104.855 177.155 105.025 177.405 ;
        RECT 105.200 177.375 105.620 177.575 ;
        RECT 105.790 177.375 106.120 177.575 ;
        RECT 106.290 177.375 106.620 177.575 ;
        RECT 106.790 177.155 106.960 177.785 ;
        RECT 107.665 177.765 108.005 178.395 ;
        RECT 108.175 177.765 108.425 178.565 ;
        RECT 108.615 177.915 108.945 178.395 ;
        RECT 109.115 178.105 109.340 178.565 ;
        RECT 109.510 177.915 109.840 178.395 ;
        RECT 107.145 177.325 107.495 177.575 ;
        RECT 107.665 177.155 107.840 177.765 ;
        RECT 108.615 177.745 109.840 177.915 ;
        RECT 110.470 177.785 110.970 178.395 ;
        RECT 111.805 177.795 114.395 178.565 ;
        RECT 114.565 177.840 114.855 178.565 ;
        RECT 115.490 177.855 115.745 178.385 ;
        RECT 115.915 178.105 116.220 178.565 ;
        RECT 116.465 178.185 117.535 178.355 ;
        RECT 108.010 177.405 108.705 177.575 ;
        RECT 108.535 177.155 108.705 177.405 ;
        RECT 108.880 177.375 109.300 177.575 ;
        RECT 109.470 177.375 109.800 177.575 ;
        RECT 109.970 177.375 110.300 177.575 ;
        RECT 110.470 177.155 110.640 177.785 ;
        RECT 110.825 177.325 111.175 177.575 ;
        RECT 103.985 176.185 104.325 177.155 ;
        RECT 104.495 176.015 104.665 177.155 ;
        RECT 104.855 176.985 107.290 177.155 ;
        RECT 104.935 176.015 105.185 176.815 ;
        RECT 105.830 176.185 106.160 176.985 ;
        RECT 106.460 176.015 106.790 176.815 ;
        RECT 106.960 176.185 107.290 176.985 ;
        RECT 107.665 176.185 108.005 177.155 ;
        RECT 108.175 176.015 108.345 177.155 ;
        RECT 108.535 176.985 110.970 177.155 ;
        RECT 108.615 176.015 108.865 176.815 ;
        RECT 109.510 176.185 109.840 176.985 ;
        RECT 110.140 176.015 110.470 176.815 ;
        RECT 110.640 176.185 110.970 176.985 ;
        RECT 111.805 177.105 113.015 177.625 ;
        RECT 113.185 177.275 114.395 177.795 ;
        RECT 115.490 177.205 115.700 177.855 ;
        RECT 116.465 177.830 116.785 178.185 ;
        RECT 116.460 177.655 116.785 177.830 ;
        RECT 115.870 177.355 116.785 177.655 ;
        RECT 116.955 177.615 117.195 178.015 ;
        RECT 117.365 177.955 117.535 178.185 ;
        RECT 117.705 178.125 117.895 178.565 ;
        RECT 118.065 178.115 119.015 178.395 ;
        RECT 119.235 178.205 119.585 178.375 ;
        RECT 117.365 177.785 117.895 177.955 ;
        RECT 115.870 177.325 116.610 177.355 ;
        RECT 111.805 176.015 114.395 177.105 ;
        RECT 114.565 176.015 114.855 177.180 ;
        RECT 115.490 176.325 115.745 177.205 ;
        RECT 115.915 176.015 116.220 177.155 ;
        RECT 116.440 176.735 116.610 177.325 ;
        RECT 116.955 177.245 117.495 177.615 ;
        RECT 117.675 177.505 117.895 177.785 ;
        RECT 118.065 177.335 118.235 178.115 ;
        RECT 117.830 177.165 118.235 177.335 ;
        RECT 118.405 177.325 118.755 177.945 ;
        RECT 117.830 177.075 118.000 177.165 ;
        RECT 118.925 177.155 119.135 177.945 ;
        RECT 116.780 176.905 118.000 177.075 ;
        RECT 118.460 176.995 119.135 177.155 ;
        RECT 116.440 176.565 117.240 176.735 ;
        RECT 116.560 176.015 116.890 176.395 ;
        RECT 117.070 176.275 117.240 176.565 ;
        RECT 117.830 176.525 118.000 176.905 ;
        RECT 118.170 176.985 119.135 176.995 ;
        RECT 119.325 177.815 119.585 178.205 ;
        RECT 119.795 178.105 120.125 178.565 ;
        RECT 121.000 178.175 121.855 178.345 ;
        RECT 122.060 178.175 122.555 178.345 ;
        RECT 122.725 178.205 123.055 178.565 ;
        RECT 119.325 177.125 119.495 177.815 ;
        RECT 119.665 177.465 119.835 177.645 ;
        RECT 120.005 177.635 120.795 177.885 ;
        RECT 121.000 177.465 121.170 178.175 ;
        RECT 121.340 177.665 121.695 177.885 ;
        RECT 119.665 177.295 121.355 177.465 ;
        RECT 118.170 176.695 118.630 176.985 ;
        RECT 119.325 176.955 120.825 177.125 ;
        RECT 119.325 176.815 119.495 176.955 ;
        RECT 118.935 176.645 119.495 176.815 ;
        RECT 117.410 176.015 117.660 176.475 ;
        RECT 117.830 176.185 118.700 176.525 ;
        RECT 118.935 176.185 119.105 176.645 ;
        RECT 119.940 176.615 121.015 176.785 ;
        RECT 119.275 176.015 119.645 176.475 ;
        RECT 119.940 176.275 120.110 176.615 ;
        RECT 120.280 176.015 120.610 176.445 ;
        RECT 120.845 176.275 121.015 176.615 ;
        RECT 121.185 176.515 121.355 177.295 ;
        RECT 121.525 177.075 121.695 177.665 ;
        RECT 121.865 177.265 122.215 177.885 ;
        RECT 121.525 176.685 121.990 177.075 ;
        RECT 122.385 176.815 122.555 178.175 ;
        RECT 122.725 176.985 123.185 178.035 ;
        RECT 122.160 176.645 122.555 176.815 ;
        RECT 122.160 176.515 122.330 176.645 ;
        RECT 121.185 176.185 121.865 176.515 ;
        RECT 122.080 176.185 122.330 176.515 ;
        RECT 122.500 176.015 122.750 176.475 ;
        RECT 122.920 176.200 123.245 176.985 ;
        RECT 123.415 176.185 123.585 178.305 ;
        RECT 123.755 178.185 124.085 178.565 ;
        RECT 124.255 178.015 124.510 178.305 ;
        RECT 123.760 177.845 124.510 178.015 ;
        RECT 123.760 176.855 123.990 177.845 ;
        RECT 124.685 177.795 126.355 178.565 ;
        RECT 126.525 177.815 127.735 178.565 ;
        RECT 124.160 177.025 124.510 177.675 ;
        RECT 124.685 177.105 125.435 177.625 ;
        RECT 125.605 177.275 126.355 177.795 ;
        RECT 126.525 177.105 127.045 177.645 ;
        RECT 127.215 177.275 127.735 177.815 ;
        RECT 123.760 176.685 124.510 176.855 ;
        RECT 123.755 176.015 124.085 176.515 ;
        RECT 124.255 176.185 124.510 176.685 ;
        RECT 124.685 176.015 126.355 177.105 ;
        RECT 126.525 176.015 127.735 177.105 ;
        RECT 14.660 175.845 127.820 176.015 ;
        RECT 14.745 174.755 15.955 175.845 ;
        RECT 16.130 175.410 21.475 175.845 ;
        RECT 14.745 174.045 15.265 174.585 ;
        RECT 15.435 174.215 15.955 174.755 ;
        RECT 17.720 174.160 18.070 175.410 ;
        RECT 21.705 174.705 21.915 175.845 ;
        RECT 22.085 174.695 22.415 175.675 ;
        RECT 22.585 174.705 22.815 175.845 ;
        RECT 23.065 174.705 23.295 175.845 ;
        RECT 23.465 174.695 23.795 175.675 ;
        RECT 23.965 174.705 24.175 175.845 ;
        RECT 14.745 173.295 15.955 174.045 ;
        RECT 19.550 173.840 19.890 174.670 ;
        RECT 16.130 173.295 21.475 173.840 ;
        RECT 21.705 173.295 21.915 174.115 ;
        RECT 22.085 174.095 22.335 174.695 ;
        RECT 22.505 174.285 22.835 174.535 ;
        RECT 23.045 174.285 23.375 174.535 ;
        RECT 22.085 173.465 22.415 174.095 ;
        RECT 22.585 173.295 22.815 174.115 ;
        RECT 23.065 173.295 23.295 174.115 ;
        RECT 23.545 174.095 23.795 174.695 ;
        RECT 24.405 174.680 24.695 175.845 ;
        RECT 25.785 174.770 26.055 175.675 ;
        RECT 26.225 175.085 26.555 175.845 ;
        RECT 26.735 174.915 26.905 175.675 ;
        RECT 27.170 175.175 27.425 175.675 ;
        RECT 27.595 175.345 27.925 175.845 ;
        RECT 27.170 175.005 27.920 175.175 ;
        RECT 23.465 173.465 23.795 174.095 ;
        RECT 23.965 173.295 24.175 174.115 ;
        RECT 24.405 173.295 24.695 174.020 ;
        RECT 25.785 173.970 25.955 174.770 ;
        RECT 26.240 174.745 26.905 174.915 ;
        RECT 26.240 174.600 26.410 174.745 ;
        RECT 26.125 174.270 26.410 174.600 ;
        RECT 26.240 174.015 26.410 174.270 ;
        RECT 26.645 174.195 26.975 174.565 ;
        RECT 27.170 174.185 27.520 174.835 ;
        RECT 27.690 174.015 27.920 175.005 ;
        RECT 25.785 173.465 26.045 173.970 ;
        RECT 26.240 173.845 26.905 174.015 ;
        RECT 26.225 173.295 26.555 173.675 ;
        RECT 26.735 173.465 26.905 173.845 ;
        RECT 27.170 173.845 27.920 174.015 ;
        RECT 27.170 173.555 27.425 173.845 ;
        RECT 27.595 173.295 27.925 173.675 ;
        RECT 28.095 173.555 28.265 175.675 ;
        RECT 28.435 174.875 28.760 175.660 ;
        RECT 28.930 175.385 29.180 175.845 ;
        RECT 29.350 175.345 29.600 175.675 ;
        RECT 29.815 175.345 30.495 175.675 ;
        RECT 29.350 175.215 29.520 175.345 ;
        RECT 29.125 175.045 29.520 175.215 ;
        RECT 28.495 173.825 28.955 174.875 ;
        RECT 29.125 173.685 29.295 175.045 ;
        RECT 29.690 174.785 30.155 175.175 ;
        RECT 29.465 173.975 29.815 174.595 ;
        RECT 29.985 174.195 30.155 174.785 ;
        RECT 30.325 174.565 30.495 175.345 ;
        RECT 30.665 175.245 30.835 175.585 ;
        RECT 31.070 175.415 31.400 175.845 ;
        RECT 31.570 175.245 31.740 175.585 ;
        RECT 32.035 175.385 32.405 175.845 ;
        RECT 30.665 175.075 31.740 175.245 ;
        RECT 32.575 175.215 32.745 175.675 ;
        RECT 32.980 175.335 33.850 175.675 ;
        RECT 34.020 175.385 34.270 175.845 ;
        RECT 32.185 175.045 32.745 175.215 ;
        RECT 32.185 174.905 32.355 175.045 ;
        RECT 30.855 174.735 32.355 174.905 ;
        RECT 33.050 174.875 33.510 175.165 ;
        RECT 30.325 174.395 32.015 174.565 ;
        RECT 29.985 173.975 30.340 174.195 ;
        RECT 30.510 173.685 30.680 174.395 ;
        RECT 30.885 173.975 31.675 174.225 ;
        RECT 31.845 174.215 32.015 174.395 ;
        RECT 32.185 174.045 32.355 174.735 ;
        RECT 28.625 173.295 28.955 173.655 ;
        RECT 29.125 173.515 29.620 173.685 ;
        RECT 29.825 173.515 30.680 173.685 ;
        RECT 31.555 173.295 31.885 173.755 ;
        RECT 32.095 173.655 32.355 174.045 ;
        RECT 32.545 174.865 33.510 174.875 ;
        RECT 33.680 174.955 33.850 175.335 ;
        RECT 34.440 175.295 34.610 175.585 ;
        RECT 34.790 175.465 35.120 175.845 ;
        RECT 34.440 175.125 35.240 175.295 ;
        RECT 32.545 174.705 33.220 174.865 ;
        RECT 33.680 174.785 34.900 174.955 ;
        RECT 32.545 173.915 32.755 174.705 ;
        RECT 33.680 174.695 33.850 174.785 ;
        RECT 32.925 173.915 33.275 174.535 ;
        RECT 33.445 174.525 33.850 174.695 ;
        RECT 33.445 173.745 33.615 174.525 ;
        RECT 33.785 174.075 34.005 174.355 ;
        RECT 34.185 174.245 34.725 174.615 ;
        RECT 35.070 174.535 35.240 175.125 ;
        RECT 35.460 174.705 35.765 175.845 ;
        RECT 35.935 174.655 36.190 175.535 ;
        RECT 35.070 174.505 35.810 174.535 ;
        RECT 33.785 173.905 34.315 174.075 ;
        RECT 32.095 173.485 32.445 173.655 ;
        RECT 32.665 173.465 33.615 173.745 ;
        RECT 33.785 173.295 33.975 173.735 ;
        RECT 34.145 173.675 34.315 173.905 ;
        RECT 34.485 173.845 34.725 174.245 ;
        RECT 34.895 174.205 35.810 174.505 ;
        RECT 34.895 174.030 35.220 174.205 ;
        RECT 34.895 173.675 35.215 174.030 ;
        RECT 35.980 174.005 36.190 174.655 ;
        RECT 34.145 173.505 35.215 173.675 ;
        RECT 35.460 173.295 35.765 173.755 ;
        RECT 35.935 173.475 36.190 174.005 ;
        RECT 36.370 174.705 36.705 175.675 ;
        RECT 36.875 174.705 37.045 175.845 ;
        RECT 37.215 175.505 39.245 175.675 ;
        RECT 36.370 174.035 36.540 174.705 ;
        RECT 37.215 174.535 37.385 175.505 ;
        RECT 36.710 174.205 36.965 174.535 ;
        RECT 37.190 174.205 37.385 174.535 ;
        RECT 37.555 175.165 38.680 175.335 ;
        RECT 36.795 174.035 36.965 174.205 ;
        RECT 37.555 174.035 37.725 175.165 ;
        RECT 36.370 173.465 36.625 174.035 ;
        RECT 36.795 173.865 37.725 174.035 ;
        RECT 37.895 174.825 38.905 174.995 ;
        RECT 37.895 174.025 38.065 174.825 ;
        RECT 38.270 174.485 38.545 174.625 ;
        RECT 38.265 174.315 38.545 174.485 ;
        RECT 37.550 173.830 37.725 173.865 ;
        RECT 36.795 173.295 37.125 173.695 ;
        RECT 37.550 173.465 38.080 173.830 ;
        RECT 38.270 173.465 38.545 174.315 ;
        RECT 38.715 173.465 38.905 174.825 ;
        RECT 39.075 174.840 39.245 175.505 ;
        RECT 39.415 175.085 39.585 175.845 ;
        RECT 39.820 175.085 40.335 175.495 ;
        RECT 39.075 174.650 39.825 174.840 ;
        RECT 39.995 174.275 40.335 175.085 ;
        RECT 39.105 174.105 40.335 174.275 ;
        RECT 40.965 174.755 42.635 175.845 ;
        RECT 40.965 174.235 41.715 174.755 ;
        RECT 42.805 174.705 43.145 175.675 ;
        RECT 43.315 174.705 43.485 175.845 ;
        RECT 43.755 175.045 44.005 175.845 ;
        RECT 44.650 174.875 44.980 175.675 ;
        RECT 45.280 175.045 45.610 175.845 ;
        RECT 45.780 174.875 46.110 175.675 ;
        RECT 43.675 174.705 46.110 174.875 ;
        RECT 46.690 174.875 47.020 175.675 ;
        RECT 47.190 175.045 47.520 175.845 ;
        RECT 47.820 174.875 48.150 175.675 ;
        RECT 48.795 175.045 49.045 175.845 ;
        RECT 46.690 174.705 49.125 174.875 ;
        RECT 49.315 174.705 49.485 175.845 ;
        RECT 49.655 174.705 49.995 175.675 ;
        RECT 39.085 173.295 39.595 173.830 ;
        RECT 39.815 173.500 40.060 174.105 ;
        RECT 41.885 174.065 42.635 174.585 ;
        RECT 40.965 173.295 42.635 174.065 ;
        RECT 42.805 174.145 42.980 174.705 ;
        RECT 43.675 174.455 43.845 174.705 ;
        RECT 43.150 174.285 43.845 174.455 ;
        RECT 44.020 174.285 44.440 174.485 ;
        RECT 44.610 174.285 44.940 174.485 ;
        RECT 45.110 174.285 45.440 174.485 ;
        RECT 42.805 174.095 43.035 174.145 ;
        RECT 42.805 173.465 43.145 174.095 ;
        RECT 43.315 173.295 43.565 174.095 ;
        RECT 43.755 173.945 44.980 174.115 ;
        RECT 43.755 173.465 44.085 173.945 ;
        RECT 44.255 173.295 44.480 173.755 ;
        RECT 44.650 173.465 44.980 173.945 ;
        RECT 45.610 174.075 45.780 174.705 ;
        RECT 45.965 174.285 46.315 174.535 ;
        RECT 46.485 174.285 46.835 174.535 ;
        RECT 47.020 174.075 47.190 174.705 ;
        RECT 47.360 174.285 47.690 174.485 ;
        RECT 47.860 174.285 48.190 174.485 ;
        RECT 48.360 174.285 48.780 174.485 ;
        RECT 48.955 174.455 49.125 174.705 ;
        RECT 48.955 174.285 49.650 174.455 ;
        RECT 49.820 174.145 49.995 174.705 ;
        RECT 50.165 174.680 50.455 175.845 ;
        RECT 51.545 174.705 51.885 175.675 ;
        RECT 52.055 174.705 52.225 175.845 ;
        RECT 52.495 175.045 52.745 175.845 ;
        RECT 53.390 174.875 53.720 175.675 ;
        RECT 54.020 175.045 54.350 175.845 ;
        RECT 54.520 174.875 54.850 175.675 ;
        RECT 52.415 174.705 54.850 174.875 ;
        RECT 55.225 174.755 56.435 175.845 ;
        RECT 56.660 174.975 56.945 175.845 ;
        RECT 57.115 175.215 57.375 175.675 ;
        RECT 57.550 175.385 57.805 175.845 ;
        RECT 57.975 175.215 58.235 175.675 ;
        RECT 57.115 175.045 58.235 175.215 ;
        RECT 58.405 175.045 58.715 175.845 ;
        RECT 57.115 174.795 57.375 175.045 ;
        RECT 58.885 174.875 59.195 175.675 ;
        RECT 45.610 173.465 46.110 174.075 ;
        RECT 46.690 173.465 47.190 174.075 ;
        RECT 47.820 173.945 49.045 174.115 ;
        RECT 49.765 174.095 49.995 174.145 ;
        RECT 47.820 173.465 48.150 173.945 ;
        RECT 48.320 173.295 48.545 173.755 ;
        RECT 48.715 173.465 49.045 173.945 ;
        RECT 49.235 173.295 49.485 174.095 ;
        RECT 49.655 173.465 49.995 174.095 ;
        RECT 51.545 174.145 51.720 174.705 ;
        RECT 52.415 174.455 52.585 174.705 ;
        RECT 51.890 174.285 52.585 174.455 ;
        RECT 52.760 174.285 53.180 174.485 ;
        RECT 53.350 174.285 53.680 174.485 ;
        RECT 53.850 174.285 54.180 174.485 ;
        RECT 51.545 174.095 51.775 174.145 ;
        RECT 50.165 173.295 50.455 174.020 ;
        RECT 51.545 173.465 51.885 174.095 ;
        RECT 52.055 173.295 52.305 174.095 ;
        RECT 52.495 173.945 53.720 174.115 ;
        RECT 52.495 173.465 52.825 173.945 ;
        RECT 52.995 173.295 53.220 173.755 ;
        RECT 53.390 173.465 53.720 173.945 ;
        RECT 54.350 174.075 54.520 174.705 ;
        RECT 54.705 174.285 55.055 174.535 ;
        RECT 55.225 174.215 55.745 174.755 ;
        RECT 56.620 174.625 57.375 174.795 ;
        RECT 58.165 174.705 59.195 174.875 ;
        RECT 54.350 173.465 54.850 174.075 ;
        RECT 55.915 174.045 56.435 174.585 ;
        RECT 55.225 173.295 56.435 174.045 ;
        RECT 56.620 174.115 57.025 174.625 ;
        RECT 58.165 174.455 58.335 174.705 ;
        RECT 57.195 174.285 58.335 174.455 ;
        RECT 56.620 173.945 58.270 174.115 ;
        RECT 58.505 173.965 58.855 174.535 ;
        RECT 56.665 173.295 56.945 173.775 ;
        RECT 57.115 173.555 57.375 173.945 ;
        RECT 57.550 173.295 57.805 173.775 ;
        RECT 57.975 173.555 58.270 173.945 ;
        RECT 59.025 173.795 59.195 174.705 ;
        RECT 59.365 174.755 61.955 175.845 ;
        RECT 59.365 174.235 60.575 174.755 ;
        RECT 62.130 174.695 62.390 175.845 ;
        RECT 62.565 174.770 62.820 175.675 ;
        RECT 62.990 175.085 63.320 175.845 ;
        RECT 63.535 174.915 63.705 175.675 ;
        RECT 60.745 174.065 61.955 174.585 ;
        RECT 58.450 173.295 58.725 173.775 ;
        RECT 58.895 173.465 59.195 173.795 ;
        RECT 59.365 173.295 61.955 174.065 ;
        RECT 62.130 173.295 62.390 174.135 ;
        RECT 62.565 174.040 62.735 174.770 ;
        RECT 62.990 174.745 63.705 174.915 ;
        RECT 62.990 174.535 63.160 174.745 ;
        RECT 62.905 174.205 63.160 174.535 ;
        RECT 62.565 173.465 62.820 174.040 ;
        RECT 62.990 174.015 63.160 174.205 ;
        RECT 63.440 174.195 63.795 174.565 ;
        RECT 63.965 174.035 64.225 175.660 ;
        RECT 65.975 175.395 66.305 175.845 ;
        RECT 64.405 175.005 67.015 175.215 ;
        RECT 64.405 174.205 64.625 175.005 ;
        RECT 64.865 174.205 65.165 174.825 ;
        RECT 65.335 174.205 65.665 174.825 ;
        RECT 65.835 174.205 66.155 174.825 ;
        RECT 66.325 174.205 66.675 174.825 ;
        RECT 66.845 174.035 67.015 175.005 ;
        RECT 62.990 173.845 63.705 174.015 ;
        RECT 63.965 173.865 65.805 174.035 ;
        RECT 62.990 173.295 63.320 173.675 ;
        RECT 63.535 173.465 63.705 173.845 ;
        RECT 64.235 173.295 64.565 173.690 ;
        RECT 64.735 173.510 64.935 173.865 ;
        RECT 65.105 173.295 65.435 173.695 ;
        RECT 65.605 173.520 65.805 173.865 ;
        RECT 65.975 173.295 66.305 174.035 ;
        RECT 66.540 173.865 67.015 174.035 ;
        RECT 67.185 174.035 67.445 175.660 ;
        RECT 69.195 175.395 69.525 175.845 ;
        RECT 67.625 175.005 70.235 175.215 ;
        RECT 67.625 174.205 67.845 175.005 ;
        RECT 68.085 174.205 68.385 174.825 ;
        RECT 68.555 174.205 68.885 174.825 ;
        RECT 69.055 174.205 69.375 174.825 ;
        RECT 69.545 174.205 69.895 174.825 ;
        RECT 70.065 174.035 70.235 175.005 ;
        RECT 67.185 173.865 69.025 174.035 ;
        RECT 66.540 173.615 66.710 173.865 ;
        RECT 67.455 173.295 67.785 173.690 ;
        RECT 67.955 173.510 68.155 173.865 ;
        RECT 68.325 173.295 68.655 173.695 ;
        RECT 68.825 173.520 69.025 173.865 ;
        RECT 69.195 173.295 69.525 174.035 ;
        RECT 69.760 173.865 70.235 174.035 ;
        RECT 70.405 174.035 70.665 175.660 ;
        RECT 72.415 175.395 72.745 175.845 ;
        RECT 70.845 175.005 73.455 175.215 ;
        RECT 70.845 174.205 71.065 175.005 ;
        RECT 71.305 174.205 71.605 174.825 ;
        RECT 71.775 174.205 72.105 174.825 ;
        RECT 72.275 174.205 72.595 174.825 ;
        RECT 72.765 174.205 73.115 174.825 ;
        RECT 73.285 174.035 73.455 175.005 ;
        RECT 74.085 174.755 75.755 175.845 ;
        RECT 74.085 174.235 74.835 174.755 ;
        RECT 75.925 174.680 76.215 175.845 ;
        RECT 77.510 174.875 77.840 175.675 ;
        RECT 78.010 175.045 78.340 175.845 ;
        RECT 78.640 174.875 78.970 175.675 ;
        RECT 79.615 175.045 79.865 175.845 ;
        RECT 77.510 174.705 79.945 174.875 ;
        RECT 80.135 174.705 80.305 175.845 ;
        RECT 80.475 174.705 80.815 175.675 ;
        RECT 75.005 174.065 75.755 174.585 ;
        RECT 77.305 174.285 77.655 174.535 ;
        RECT 77.840 174.075 78.010 174.705 ;
        RECT 78.180 174.285 78.510 174.485 ;
        RECT 78.680 174.285 79.010 174.485 ;
        RECT 79.180 174.285 79.600 174.485 ;
        RECT 79.775 174.455 79.945 174.705 ;
        RECT 79.775 174.285 80.470 174.455 ;
        RECT 80.640 174.145 80.815 174.705 ;
        RECT 81.445 174.755 84.035 175.845 ;
        RECT 84.295 175.100 84.565 175.845 ;
        RECT 85.195 175.840 91.470 175.845 ;
        RECT 84.735 174.930 85.025 175.670 ;
        RECT 85.195 175.115 85.450 175.840 ;
        RECT 85.635 174.945 85.895 175.670 ;
        RECT 86.065 175.115 86.310 175.840 ;
        RECT 86.495 174.945 86.755 175.670 ;
        RECT 86.925 175.115 87.170 175.840 ;
        RECT 87.355 174.945 87.615 175.670 ;
        RECT 87.785 175.115 88.030 175.840 ;
        RECT 88.200 174.945 88.460 175.670 ;
        RECT 88.630 175.115 88.890 175.840 ;
        RECT 89.060 174.945 89.320 175.670 ;
        RECT 89.490 175.115 89.750 175.840 ;
        RECT 89.920 174.945 90.180 175.670 ;
        RECT 90.350 175.115 90.610 175.840 ;
        RECT 90.780 174.945 91.040 175.670 ;
        RECT 91.210 175.045 91.470 175.840 ;
        RECT 85.635 174.930 91.040 174.945 ;
        RECT 81.445 174.235 82.655 174.755 ;
        RECT 84.295 174.705 91.040 174.930 ;
        RECT 70.405 173.865 72.245 174.035 ;
        RECT 69.760 173.615 69.930 173.865 ;
        RECT 70.675 173.295 71.005 173.690 ;
        RECT 71.175 173.510 71.375 173.865 ;
        RECT 71.545 173.295 71.875 173.695 ;
        RECT 72.045 173.520 72.245 173.865 ;
        RECT 72.415 173.295 72.745 174.035 ;
        RECT 72.980 173.865 73.455 174.035 ;
        RECT 72.980 173.615 73.150 173.865 ;
        RECT 74.085 173.295 75.755 174.065 ;
        RECT 75.925 173.295 76.215 174.020 ;
        RECT 77.510 173.465 78.010 174.075 ;
        RECT 78.640 173.945 79.865 174.115 ;
        RECT 80.585 174.095 80.815 174.145 ;
        RECT 78.640 173.465 78.970 173.945 ;
        RECT 79.140 173.295 79.365 173.755 ;
        RECT 79.535 173.465 79.865 173.945 ;
        RECT 80.055 173.295 80.305 174.095 ;
        RECT 80.475 173.465 80.815 174.095 ;
        RECT 82.825 174.065 84.035 174.585 ;
        RECT 81.445 173.295 84.035 174.065 ;
        RECT 84.295 174.115 85.460 174.705 ;
        RECT 91.640 174.535 91.890 175.670 ;
        RECT 92.070 175.035 92.330 175.845 ;
        RECT 92.505 174.535 92.750 175.675 ;
        RECT 92.930 175.035 93.225 175.845 ;
        RECT 94.325 174.755 97.835 175.845 ;
        RECT 85.630 174.285 92.750 174.535 ;
        RECT 84.295 173.945 91.040 174.115 ;
        RECT 84.295 173.295 84.595 173.775 ;
        RECT 84.765 173.490 85.025 173.945 ;
        RECT 85.195 173.295 85.455 173.775 ;
        RECT 85.635 173.490 85.895 173.945 ;
        RECT 86.065 173.295 86.315 173.775 ;
        RECT 86.495 173.490 86.755 173.945 ;
        RECT 86.925 173.295 87.175 173.775 ;
        RECT 87.355 173.490 87.615 173.945 ;
        RECT 87.785 173.295 88.030 173.775 ;
        RECT 88.200 173.490 88.475 173.945 ;
        RECT 88.645 173.295 88.890 173.775 ;
        RECT 89.060 173.490 89.320 173.945 ;
        RECT 89.490 173.295 89.750 173.775 ;
        RECT 89.920 173.490 90.180 173.945 ;
        RECT 90.350 173.295 90.610 173.775 ;
        RECT 90.780 173.490 91.040 173.945 ;
        RECT 91.210 173.295 91.470 173.855 ;
        RECT 91.640 173.475 91.890 174.285 ;
        RECT 92.070 173.295 92.330 173.820 ;
        RECT 92.500 173.475 92.750 174.285 ;
        RECT 92.920 173.975 93.235 174.535 ;
        RECT 94.325 174.235 96.015 174.755 ;
        RECT 98.005 174.705 98.345 175.675 ;
        RECT 98.515 174.705 98.685 175.845 ;
        RECT 98.955 175.045 99.205 175.845 ;
        RECT 99.850 174.875 100.180 175.675 ;
        RECT 100.480 175.045 100.810 175.845 ;
        RECT 100.980 174.875 101.310 175.675 ;
        RECT 98.875 174.705 101.310 174.875 ;
        RECT 96.185 174.065 97.835 174.585 ;
        RECT 92.930 173.295 93.235 173.805 ;
        RECT 94.325 173.295 97.835 174.065 ;
        RECT 98.005 174.145 98.180 174.705 ;
        RECT 98.875 174.455 99.045 174.705 ;
        RECT 98.350 174.285 99.045 174.455 ;
        RECT 99.220 174.285 99.640 174.485 ;
        RECT 99.810 174.285 100.140 174.485 ;
        RECT 100.310 174.285 100.640 174.485 ;
        RECT 98.005 174.095 98.235 174.145 ;
        RECT 98.005 173.465 98.345 174.095 ;
        RECT 98.515 173.295 98.765 174.095 ;
        RECT 98.955 173.945 100.180 174.115 ;
        RECT 98.955 173.465 99.285 173.945 ;
        RECT 99.455 173.295 99.680 173.755 ;
        RECT 99.850 173.465 100.180 173.945 ;
        RECT 100.810 174.075 100.980 174.705 ;
        RECT 101.685 174.680 101.975 175.845 ;
        RECT 102.605 174.755 104.275 175.845 ;
        RECT 104.500 174.975 104.785 175.845 ;
        RECT 104.955 175.215 105.215 175.675 ;
        RECT 105.390 175.385 105.645 175.845 ;
        RECT 105.815 175.215 106.075 175.675 ;
        RECT 104.955 175.045 106.075 175.215 ;
        RECT 106.245 175.045 106.555 175.845 ;
        RECT 104.955 174.795 105.215 175.045 ;
        RECT 106.725 174.875 107.035 175.675 ;
        RECT 101.165 174.285 101.515 174.535 ;
        RECT 102.605 174.235 103.355 174.755 ;
        RECT 104.460 174.625 105.215 174.795 ;
        RECT 106.005 174.705 107.035 174.875 ;
        RECT 100.810 173.465 101.310 174.075 ;
        RECT 103.525 174.065 104.275 174.585 ;
        RECT 101.685 173.295 101.975 174.020 ;
        RECT 102.605 173.295 104.275 174.065 ;
        RECT 104.460 174.115 104.865 174.625 ;
        RECT 106.005 174.455 106.175 174.705 ;
        RECT 105.035 174.285 106.175 174.455 ;
        RECT 104.460 173.945 106.110 174.115 ;
        RECT 106.345 173.965 106.695 174.535 ;
        RECT 104.505 173.295 104.785 173.775 ;
        RECT 104.955 173.555 105.215 173.945 ;
        RECT 105.390 173.295 105.645 173.775 ;
        RECT 105.815 173.555 106.110 173.945 ;
        RECT 106.865 173.795 107.035 174.705 ;
        RECT 106.290 173.295 106.565 173.775 ;
        RECT 106.735 173.465 107.035 173.795 ;
        RECT 107.205 174.705 107.545 175.675 ;
        RECT 107.715 174.705 107.885 175.845 ;
        RECT 108.155 175.045 108.405 175.845 ;
        RECT 109.050 174.875 109.380 175.675 ;
        RECT 109.680 175.045 110.010 175.845 ;
        RECT 110.180 174.875 110.510 175.675 ;
        RECT 108.075 174.705 110.510 174.875 ;
        RECT 110.885 174.755 112.555 175.845 ;
        RECT 112.730 175.410 118.075 175.845 ;
        RECT 107.205 174.145 107.380 174.705 ;
        RECT 108.075 174.455 108.245 174.705 ;
        RECT 107.550 174.285 108.245 174.455 ;
        RECT 108.420 174.285 108.840 174.485 ;
        RECT 109.010 174.285 109.340 174.485 ;
        RECT 109.510 174.285 109.840 174.485 ;
        RECT 107.205 174.095 107.435 174.145 ;
        RECT 107.205 173.465 107.545 174.095 ;
        RECT 107.715 173.295 107.965 174.095 ;
        RECT 108.155 173.945 109.380 174.115 ;
        RECT 108.155 173.465 108.485 173.945 ;
        RECT 108.655 173.295 108.880 173.755 ;
        RECT 109.050 173.465 109.380 173.945 ;
        RECT 110.010 174.075 110.180 174.705 ;
        RECT 110.365 174.285 110.715 174.535 ;
        RECT 110.885 174.235 111.635 174.755 ;
        RECT 110.010 173.465 110.510 174.075 ;
        RECT 111.805 174.065 112.555 174.585 ;
        RECT 114.320 174.160 114.670 175.410 ;
        RECT 118.285 174.705 118.515 175.845 ;
        RECT 118.685 174.695 119.015 175.675 ;
        RECT 119.185 174.705 119.395 175.845 ;
        RECT 120.175 174.915 120.345 175.675 ;
        RECT 120.525 175.085 120.855 175.845 ;
        RECT 120.175 174.745 120.840 174.915 ;
        RECT 121.025 174.770 121.295 175.675 ;
        RECT 110.885 173.295 112.555 174.065 ;
        RECT 116.150 173.840 116.490 174.670 ;
        RECT 118.265 174.285 118.595 174.535 ;
        RECT 112.730 173.295 118.075 173.840 ;
        RECT 118.285 173.295 118.515 174.115 ;
        RECT 118.765 174.095 119.015 174.695 ;
        RECT 120.670 174.600 120.840 174.745 ;
        RECT 120.105 174.195 120.435 174.565 ;
        RECT 120.670 174.270 120.955 174.600 ;
        RECT 118.685 173.465 119.015 174.095 ;
        RECT 119.185 173.295 119.395 174.115 ;
        RECT 120.670 174.015 120.840 174.270 ;
        RECT 120.175 173.845 120.840 174.015 ;
        RECT 121.125 173.970 121.295 174.770 ;
        RECT 121.465 174.755 122.675 175.845 ;
        RECT 122.845 174.755 126.355 175.845 ;
        RECT 126.525 174.755 127.735 175.845 ;
        RECT 121.465 174.215 121.985 174.755 ;
        RECT 122.155 174.045 122.675 174.585 ;
        RECT 122.845 174.235 124.535 174.755 ;
        RECT 124.705 174.065 126.355 174.585 ;
        RECT 126.525 174.215 127.045 174.755 ;
        RECT 120.175 173.465 120.345 173.845 ;
        RECT 120.525 173.295 120.855 173.675 ;
        RECT 121.035 173.465 121.295 173.970 ;
        RECT 121.465 173.295 122.675 174.045 ;
        RECT 122.845 173.295 126.355 174.065 ;
        RECT 127.215 174.045 127.735 174.585 ;
        RECT 126.525 173.295 127.735 174.045 ;
        RECT 14.660 173.125 127.820 173.295 ;
        RECT 14.745 172.375 15.955 173.125 ;
        RECT 16.125 172.375 17.335 173.125 ;
        RECT 14.745 171.835 15.265 172.375 ;
        RECT 15.435 171.665 15.955 172.205 ;
        RECT 14.745 170.575 15.955 171.665 ;
        RECT 16.125 171.665 16.645 172.205 ;
        RECT 16.815 171.835 17.335 172.375 ;
        RECT 17.505 172.355 21.015 173.125 ;
        RECT 21.295 172.645 21.465 173.125 ;
        RECT 21.635 172.475 21.965 172.950 ;
        RECT 22.135 172.645 22.305 173.125 ;
        RECT 22.475 172.475 22.805 172.950 ;
        RECT 22.975 172.645 23.145 173.125 ;
        RECT 23.315 172.475 23.645 172.950 ;
        RECT 23.815 172.645 23.985 173.125 ;
        RECT 24.155 172.475 24.485 172.950 ;
        RECT 24.655 172.645 24.825 173.125 ;
        RECT 24.995 172.475 25.325 172.950 ;
        RECT 25.495 172.645 25.665 173.125 ;
        RECT 25.915 172.950 26.085 172.955 ;
        RECT 25.835 172.475 26.165 172.950 ;
        RECT 26.335 172.645 26.505 173.125 ;
        RECT 26.755 172.950 26.925 172.955 ;
        RECT 26.675 172.475 27.005 172.950 ;
        RECT 27.175 172.645 27.345 173.125 ;
        RECT 27.595 172.950 27.845 172.955 ;
        RECT 27.515 172.475 27.845 172.950 ;
        RECT 28.015 172.645 28.185 173.125 ;
        RECT 28.355 172.475 28.685 172.950 ;
        RECT 28.855 172.645 29.025 173.125 ;
        RECT 29.195 172.475 29.525 172.950 ;
        RECT 29.695 172.645 29.865 173.125 ;
        RECT 30.035 172.475 30.365 172.950 ;
        RECT 30.535 172.645 30.705 173.125 ;
        RECT 30.875 172.475 31.205 172.950 ;
        RECT 31.375 172.645 31.545 173.125 ;
        RECT 31.715 172.475 32.045 172.950 ;
        RECT 17.505 171.665 19.195 172.185 ;
        RECT 19.365 171.835 21.015 172.355 ;
        RECT 21.185 172.305 27.845 172.475 ;
        RECT 28.015 172.305 30.365 172.475 ;
        RECT 30.535 172.305 32.045 172.475 ;
        RECT 32.230 172.385 32.485 172.955 ;
        RECT 32.655 172.725 32.985 173.125 ;
        RECT 33.410 172.590 33.940 172.955 ;
        RECT 33.410 172.555 33.585 172.590 ;
        RECT 32.655 172.385 33.585 172.555 ;
        RECT 21.185 171.765 21.460 172.305 ;
        RECT 28.015 172.135 28.190 172.305 ;
        RECT 30.535 172.135 30.705 172.305 ;
        RECT 21.630 171.935 28.190 172.135 ;
        RECT 28.395 171.935 30.705 172.135 ;
        RECT 30.875 171.935 32.050 172.135 ;
        RECT 28.015 171.765 28.190 171.935 ;
        RECT 30.535 171.765 30.705 171.935 ;
        RECT 16.125 170.575 17.335 171.665 ;
        RECT 17.505 170.575 21.015 171.665 ;
        RECT 21.185 171.595 27.845 171.765 ;
        RECT 28.015 171.595 30.365 171.765 ;
        RECT 30.535 171.595 32.045 171.765 ;
        RECT 21.295 170.575 21.465 171.375 ;
        RECT 21.635 170.745 21.965 171.595 ;
        RECT 22.135 170.575 22.305 171.375 ;
        RECT 22.475 170.745 22.805 171.595 ;
        RECT 22.975 170.575 23.145 171.375 ;
        RECT 23.315 170.745 23.645 171.595 ;
        RECT 23.815 170.575 23.985 171.375 ;
        RECT 24.155 170.745 24.485 171.595 ;
        RECT 24.655 170.575 24.825 171.375 ;
        RECT 24.995 170.745 25.325 171.595 ;
        RECT 25.495 170.575 25.665 171.375 ;
        RECT 25.835 170.745 26.165 171.595 ;
        RECT 26.335 170.575 26.505 171.375 ;
        RECT 26.675 170.745 27.005 171.595 ;
        RECT 27.175 170.575 27.345 171.375 ;
        RECT 27.515 170.745 27.845 171.595 ;
        RECT 28.015 170.575 28.185 171.375 ;
        RECT 28.355 170.745 28.685 171.595 ;
        RECT 28.855 170.575 29.025 171.375 ;
        RECT 29.195 170.745 29.525 171.595 ;
        RECT 29.695 170.575 29.865 171.375 ;
        RECT 30.035 170.745 30.365 171.595 ;
        RECT 30.535 170.575 30.705 171.425 ;
        RECT 30.875 170.745 31.205 171.595 ;
        RECT 31.375 170.575 31.545 171.425 ;
        RECT 31.715 170.745 32.045 171.595 ;
        RECT 32.230 171.715 32.400 172.385 ;
        RECT 32.655 172.215 32.825 172.385 ;
        RECT 32.570 171.885 32.825 172.215 ;
        RECT 33.050 171.885 33.245 172.215 ;
        RECT 32.230 170.745 32.565 171.715 ;
        RECT 32.735 170.575 32.905 171.715 ;
        RECT 33.075 170.915 33.245 171.885 ;
        RECT 33.415 171.255 33.585 172.385 ;
        RECT 33.755 171.595 33.925 172.395 ;
        RECT 34.130 172.105 34.405 172.955 ;
        RECT 34.125 171.935 34.405 172.105 ;
        RECT 34.130 171.795 34.405 171.935 ;
        RECT 34.575 171.595 34.765 172.955 ;
        RECT 34.945 172.590 35.455 173.125 ;
        RECT 35.675 172.315 35.920 172.920 ;
        RECT 37.285 172.400 37.575 173.125 ;
        RECT 37.745 172.325 38.085 172.955 ;
        RECT 38.255 172.325 38.505 173.125 ;
        RECT 38.695 172.475 39.025 172.955 ;
        RECT 39.195 172.665 39.420 173.125 ;
        RECT 39.590 172.475 39.920 172.955 ;
        RECT 34.965 172.145 36.195 172.315 ;
        RECT 33.755 171.425 34.765 171.595 ;
        RECT 34.935 171.580 35.685 171.770 ;
        RECT 33.415 171.085 34.540 171.255 ;
        RECT 34.935 170.915 35.105 171.580 ;
        RECT 35.855 171.335 36.195 172.145 ;
        RECT 33.075 170.745 35.105 170.915 ;
        RECT 35.275 170.575 35.445 171.335 ;
        RECT 35.680 170.925 36.195 171.335 ;
        RECT 37.285 170.575 37.575 171.740 ;
        RECT 37.745 171.715 37.920 172.325 ;
        RECT 38.695 172.305 39.920 172.475 ;
        RECT 40.550 172.345 41.050 172.955 ;
        RECT 38.090 171.965 38.785 172.135 ;
        RECT 38.615 171.715 38.785 171.965 ;
        RECT 38.960 171.935 39.380 172.135 ;
        RECT 39.550 171.935 39.880 172.135 ;
        RECT 40.050 171.935 40.380 172.135 ;
        RECT 40.550 171.715 40.720 172.345 ;
        RECT 41.885 172.325 42.225 172.955 ;
        RECT 42.395 172.325 42.645 173.125 ;
        RECT 42.835 172.475 43.165 172.955 ;
        RECT 43.335 172.665 43.560 173.125 ;
        RECT 43.730 172.475 44.060 172.955 ;
        RECT 40.905 171.885 41.255 172.135 ;
        RECT 41.885 171.715 42.060 172.325 ;
        RECT 42.835 172.305 44.060 172.475 ;
        RECT 44.690 172.345 45.190 172.955 ;
        RECT 42.230 171.965 42.925 172.135 ;
        RECT 42.755 171.715 42.925 171.965 ;
        RECT 43.100 171.935 43.520 172.135 ;
        RECT 43.690 171.935 44.020 172.135 ;
        RECT 44.190 171.935 44.520 172.135 ;
        RECT 44.690 171.715 44.860 172.345 ;
        RECT 45.565 172.325 45.905 172.955 ;
        RECT 46.075 172.325 46.325 173.125 ;
        RECT 46.515 172.475 46.845 172.955 ;
        RECT 47.015 172.665 47.240 173.125 ;
        RECT 47.410 172.475 47.740 172.955 ;
        RECT 45.045 171.885 45.395 172.135 ;
        RECT 45.565 171.715 45.740 172.325 ;
        RECT 46.515 172.305 47.740 172.475 ;
        RECT 48.370 172.345 48.870 172.955 ;
        RECT 49.245 172.355 52.755 173.125 ;
        RECT 52.930 172.655 53.260 173.125 ;
        RECT 53.430 172.485 53.655 172.930 ;
        RECT 53.825 172.600 54.120 173.125 ;
        RECT 45.910 171.965 46.605 172.135 ;
        RECT 46.435 171.715 46.605 171.965 ;
        RECT 46.780 171.935 47.200 172.135 ;
        RECT 47.370 171.935 47.700 172.135 ;
        RECT 47.870 171.935 48.200 172.135 ;
        RECT 48.370 171.715 48.540 172.345 ;
        RECT 48.725 171.885 49.075 172.135 ;
        RECT 37.745 170.745 38.085 171.715 ;
        RECT 38.255 170.575 38.425 171.715 ;
        RECT 38.615 171.545 41.050 171.715 ;
        RECT 38.695 170.575 38.945 171.375 ;
        RECT 39.590 170.745 39.920 171.545 ;
        RECT 40.220 170.575 40.550 171.375 ;
        RECT 40.720 170.745 41.050 171.545 ;
        RECT 41.885 170.745 42.225 171.715 ;
        RECT 42.395 170.575 42.565 171.715 ;
        RECT 42.755 171.545 45.190 171.715 ;
        RECT 42.835 170.575 43.085 171.375 ;
        RECT 43.730 170.745 44.060 171.545 ;
        RECT 44.360 170.575 44.690 171.375 ;
        RECT 44.860 170.745 45.190 171.545 ;
        RECT 45.565 170.745 45.905 171.715 ;
        RECT 46.075 170.575 46.245 171.715 ;
        RECT 46.435 171.545 48.870 171.715 ;
        RECT 46.515 170.575 46.765 171.375 ;
        RECT 47.410 170.745 47.740 171.545 ;
        RECT 48.040 170.575 48.370 171.375 ;
        RECT 48.540 170.745 48.870 171.545 ;
        RECT 49.245 171.665 50.935 172.185 ;
        RECT 51.105 171.835 52.755 172.355 ;
        RECT 52.925 172.315 53.655 172.485 ;
        RECT 54.765 172.355 57.355 173.125 ;
        RECT 57.530 172.580 62.875 173.125 ;
        RECT 52.925 171.750 53.205 172.315 ;
        RECT 53.375 171.920 54.595 172.145 ;
        RECT 49.245 170.575 52.755 171.665 ;
        RECT 52.925 171.580 54.525 171.750 ;
        RECT 52.985 170.575 53.240 171.410 ;
        RECT 53.410 170.775 53.670 171.580 ;
        RECT 53.840 170.575 54.100 171.410 ;
        RECT 54.270 170.775 54.525 171.580 ;
        RECT 54.765 171.665 55.975 172.185 ;
        RECT 56.145 171.835 57.355 172.355 ;
        RECT 54.765 170.575 57.355 171.665 ;
        RECT 59.120 171.010 59.470 172.260 ;
        RECT 60.950 171.750 61.290 172.580 ;
        RECT 63.045 172.400 63.335 173.125 ;
        RECT 64.430 172.285 64.690 173.125 ;
        RECT 64.865 172.380 65.120 172.955 ;
        RECT 65.290 172.745 65.620 173.125 ;
        RECT 65.835 172.575 66.005 172.955 ;
        RECT 66.335 172.765 66.665 173.125 ;
        RECT 67.195 172.765 67.525 173.125 ;
        RECT 68.055 172.765 68.385 173.125 ;
        RECT 68.615 172.765 70.685 172.955 ;
        RECT 68.615 172.745 69.735 172.765 ;
        RECT 65.290 172.405 66.005 172.575 ;
        RECT 66.835 172.575 67.025 172.695 ;
        RECT 57.530 170.575 62.875 171.010 ;
        RECT 63.045 170.575 63.335 171.740 ;
        RECT 64.430 170.575 64.690 171.725 ;
        RECT 64.865 171.650 65.035 172.380 ;
        RECT 65.290 172.215 65.460 172.405 ;
        RECT 65.205 171.885 65.460 172.215 ;
        RECT 65.290 171.675 65.460 171.885 ;
        RECT 65.740 171.855 66.095 172.225 ;
        RECT 66.325 172.135 66.665 172.445 ;
        RECT 66.835 172.365 69.375 172.575 ;
        RECT 69.545 172.320 69.735 172.745 ;
        RECT 66.325 171.965 67.275 172.135 ;
        RECT 66.325 171.915 67.220 171.965 ;
        RECT 67.445 171.855 68.415 172.135 ;
        RECT 68.875 171.845 69.735 172.135 ;
        RECT 64.865 170.745 65.120 171.650 ;
        RECT 65.290 171.505 66.005 171.675 ;
        RECT 65.290 170.575 65.620 171.335 ;
        RECT 65.835 170.745 66.005 171.505 ;
        RECT 66.335 171.515 67.455 171.685 ;
        RECT 69.905 171.670 70.235 172.540 ;
        RECT 66.335 170.745 66.595 171.515 ;
        RECT 66.765 170.575 67.095 171.345 ;
        RECT 67.265 170.915 67.455 171.515 ;
        RECT 67.625 171.500 70.235 171.670 ;
        RECT 67.625 171.085 67.955 171.500 ;
        RECT 68.125 170.915 68.385 171.110 ;
        RECT 67.265 170.745 68.385 170.915 ;
        RECT 68.615 170.575 68.945 171.295 ;
        RECT 69.115 170.745 69.305 171.500 ;
        RECT 69.475 170.575 69.805 171.295 ;
        RECT 69.975 170.745 70.235 171.500 ;
        RECT 70.405 171.240 70.695 172.215 ;
        RECT 70.405 170.575 70.665 171.035 ;
        RECT 70.865 170.745 71.125 172.955 ;
        RECT 71.295 172.745 71.625 173.125 ;
        RECT 71.835 172.215 72.030 172.790 ;
        RECT 72.300 172.215 72.485 172.795 ;
        RECT 71.295 171.295 71.465 172.215 ;
        RECT 71.775 171.885 72.030 172.215 ;
        RECT 72.255 171.885 72.485 172.215 ;
        RECT 72.735 172.785 74.215 172.955 ;
        RECT 72.735 171.885 72.905 172.785 ;
        RECT 73.075 172.285 73.625 172.615 ;
        RECT 73.815 172.455 74.215 172.785 ;
        RECT 74.395 172.745 74.725 173.125 ;
        RECT 75.035 172.625 75.295 172.955 ;
        RECT 71.835 171.575 72.030 171.885 ;
        RECT 72.300 171.575 72.485 171.885 ;
        RECT 73.075 171.295 73.245 172.285 ;
        RECT 73.815 171.975 73.985 172.455 ;
        RECT 74.565 172.265 74.775 172.445 ;
        RECT 74.155 172.095 74.775 172.265 ;
        RECT 71.295 171.125 73.245 171.295 ;
        RECT 73.415 171.805 73.985 171.975 ;
        RECT 75.125 171.925 75.295 172.625 ;
        RECT 75.555 172.575 75.725 172.955 ;
        RECT 75.940 172.745 76.270 173.125 ;
        RECT 75.555 172.405 76.270 172.575 ;
        RECT 73.415 171.295 73.585 171.805 ;
        RECT 74.165 171.755 75.295 171.925 ;
        RECT 75.465 171.855 75.820 172.225 ;
        RECT 76.100 172.215 76.270 172.405 ;
        RECT 76.440 172.380 76.695 172.955 ;
        RECT 76.100 171.885 76.355 172.215 ;
        RECT 74.165 171.635 74.335 171.755 ;
        RECT 73.755 171.465 74.335 171.635 ;
        RECT 73.415 171.125 74.155 171.295 ;
        RECT 74.605 171.255 74.955 171.585 ;
        RECT 71.295 170.575 71.625 170.955 ;
        RECT 72.050 170.745 72.220 171.125 ;
        RECT 72.480 170.575 72.810 170.955 ;
        RECT 73.005 170.745 73.175 171.125 ;
        RECT 73.385 170.575 73.715 170.955 ;
        RECT 73.965 170.745 74.155 171.125 ;
        RECT 75.125 171.075 75.295 171.755 ;
        RECT 76.100 171.675 76.270 171.885 ;
        RECT 74.395 170.575 74.725 170.955 ;
        RECT 75.035 170.745 75.295 171.075 ;
        RECT 75.555 171.505 76.270 171.675 ;
        RECT 76.525 171.650 76.695 172.380 ;
        RECT 76.870 172.285 77.130 173.125 ;
        RECT 78.225 172.355 81.735 173.125 ;
        RECT 75.555 170.745 75.725 171.505 ;
        RECT 75.940 170.575 76.270 171.335 ;
        RECT 76.440 170.745 76.695 171.650 ;
        RECT 76.870 170.575 77.130 171.725 ;
        RECT 78.225 171.665 79.915 172.185 ;
        RECT 80.085 171.835 81.735 172.355 ;
        RECT 81.905 172.325 82.245 172.955 ;
        RECT 82.415 172.325 82.665 173.125 ;
        RECT 82.855 172.475 83.185 172.955 ;
        RECT 83.355 172.665 83.580 173.125 ;
        RECT 83.750 172.475 84.080 172.955 ;
        RECT 81.905 171.715 82.080 172.325 ;
        RECT 82.855 172.305 84.080 172.475 ;
        RECT 84.710 172.345 85.210 172.955 ;
        RECT 86.045 172.355 88.635 173.125 ;
        RECT 88.805 172.400 89.095 173.125 ;
        RECT 89.725 172.355 91.395 173.125 ;
        RECT 91.570 172.655 91.900 173.125 ;
        RECT 92.070 172.485 92.295 172.930 ;
        RECT 92.465 172.600 92.760 173.125 ;
        RECT 82.250 171.965 82.945 172.135 ;
        RECT 82.775 171.715 82.945 171.965 ;
        RECT 83.120 171.935 83.540 172.135 ;
        RECT 83.710 171.935 84.040 172.135 ;
        RECT 84.210 171.935 84.540 172.135 ;
        RECT 84.710 171.715 84.880 172.345 ;
        RECT 85.065 171.885 85.415 172.135 ;
        RECT 78.225 170.575 81.735 171.665 ;
        RECT 81.905 170.745 82.245 171.715 ;
        RECT 82.415 170.575 82.585 171.715 ;
        RECT 82.775 171.545 85.210 171.715 ;
        RECT 82.855 170.575 83.105 171.375 ;
        RECT 83.750 170.745 84.080 171.545 ;
        RECT 84.380 170.575 84.710 171.375 ;
        RECT 84.880 170.745 85.210 171.545 ;
        RECT 86.045 171.665 87.255 172.185 ;
        RECT 87.425 171.835 88.635 172.355 ;
        RECT 86.045 170.575 88.635 171.665 ;
        RECT 88.805 170.575 89.095 171.740 ;
        RECT 89.725 171.665 90.475 172.185 ;
        RECT 90.645 171.835 91.395 172.355 ;
        RECT 91.565 172.315 92.295 172.485 ;
        RECT 93.405 172.355 95.995 173.125 ;
        RECT 96.255 172.575 96.425 172.955 ;
        RECT 96.605 172.745 96.935 173.125 ;
        RECT 96.255 172.405 96.920 172.575 ;
        RECT 97.115 172.450 97.375 172.955 ;
        RECT 91.565 171.750 91.845 172.315 ;
        RECT 92.015 171.920 93.235 172.145 ;
        RECT 89.725 170.575 91.395 171.665 ;
        RECT 91.565 171.580 93.165 171.750 ;
        RECT 91.625 170.575 91.880 171.410 ;
        RECT 92.050 170.775 92.310 171.580 ;
        RECT 92.480 170.575 92.740 171.410 ;
        RECT 92.910 170.775 93.165 171.580 ;
        RECT 93.405 171.665 94.615 172.185 ;
        RECT 94.785 171.835 95.995 172.355 ;
        RECT 96.185 171.855 96.515 172.225 ;
        RECT 96.750 172.150 96.920 172.405 ;
        RECT 96.750 171.820 97.035 172.150 ;
        RECT 96.750 171.675 96.920 171.820 ;
        RECT 93.405 170.575 95.995 171.665 ;
        RECT 96.255 171.505 96.920 171.675 ;
        RECT 97.205 171.650 97.375 172.450 ;
        RECT 98.005 172.355 100.595 173.125 ;
        RECT 100.855 172.645 101.155 173.125 ;
        RECT 101.325 172.475 101.585 172.930 ;
        RECT 101.755 172.645 102.015 173.125 ;
        RECT 102.195 172.475 102.455 172.930 ;
        RECT 102.625 172.645 102.875 173.125 ;
        RECT 103.055 172.475 103.315 172.930 ;
        RECT 103.485 172.645 103.735 173.125 ;
        RECT 103.915 172.475 104.175 172.930 ;
        RECT 104.345 172.645 104.590 173.125 ;
        RECT 104.760 172.475 105.035 172.930 ;
        RECT 105.205 172.645 105.450 173.125 ;
        RECT 105.620 172.475 105.880 172.930 ;
        RECT 106.050 172.645 106.310 173.125 ;
        RECT 106.480 172.475 106.740 172.930 ;
        RECT 106.910 172.645 107.170 173.125 ;
        RECT 107.340 172.475 107.600 172.930 ;
        RECT 107.770 172.565 108.030 173.125 ;
        RECT 96.255 170.745 96.425 171.505 ;
        RECT 96.605 170.575 96.935 171.335 ;
        RECT 97.105 170.745 97.375 171.650 ;
        RECT 98.005 171.665 99.215 172.185 ;
        RECT 99.385 171.835 100.595 172.355 ;
        RECT 100.855 172.305 107.600 172.475 ;
        RECT 100.855 171.715 102.020 172.305 ;
        RECT 108.200 172.135 108.450 172.945 ;
        RECT 108.630 172.600 108.890 173.125 ;
        RECT 109.060 172.135 109.310 172.945 ;
        RECT 109.490 172.615 109.795 173.125 ;
        RECT 102.190 171.885 109.310 172.135 ;
        RECT 109.480 171.885 109.795 172.445 ;
        RECT 110.700 172.315 110.945 172.920 ;
        RECT 111.165 172.590 111.675 173.125 ;
        RECT 110.425 172.145 111.655 172.315 ;
        RECT 98.005 170.575 100.595 171.665 ;
        RECT 100.855 171.490 107.600 171.715 ;
        RECT 100.855 170.575 101.125 171.320 ;
        RECT 101.295 170.750 101.585 171.490 ;
        RECT 102.195 171.475 107.600 171.490 ;
        RECT 101.755 170.580 102.010 171.305 ;
        RECT 102.195 170.750 102.455 171.475 ;
        RECT 102.625 170.580 102.870 171.305 ;
        RECT 103.055 170.750 103.315 171.475 ;
        RECT 103.485 170.580 103.730 171.305 ;
        RECT 103.915 170.750 104.175 171.475 ;
        RECT 104.345 170.580 104.590 171.305 ;
        RECT 104.760 170.750 105.020 171.475 ;
        RECT 105.190 170.580 105.450 171.305 ;
        RECT 105.620 170.750 105.880 171.475 ;
        RECT 106.050 170.580 106.310 171.305 ;
        RECT 106.480 170.750 106.740 171.475 ;
        RECT 106.910 170.580 107.170 171.305 ;
        RECT 107.340 170.750 107.600 171.475 ;
        RECT 107.770 170.580 108.030 171.375 ;
        RECT 108.200 170.750 108.450 171.885 ;
        RECT 101.755 170.575 108.030 170.580 ;
        RECT 108.630 170.575 108.890 171.385 ;
        RECT 109.065 170.745 109.310 171.885 ;
        RECT 109.490 170.575 109.785 171.385 ;
        RECT 110.425 171.335 110.765 172.145 ;
        RECT 110.935 171.580 111.685 171.770 ;
        RECT 110.425 170.925 110.940 171.335 ;
        RECT 111.175 170.575 111.345 171.335 ;
        RECT 111.515 170.915 111.685 171.580 ;
        RECT 111.855 171.595 112.045 172.955 ;
        RECT 112.215 172.105 112.490 172.955 ;
        RECT 112.680 172.590 113.210 172.955 ;
        RECT 113.635 172.725 113.965 173.125 ;
        RECT 113.035 172.555 113.210 172.590 ;
        RECT 112.215 171.935 112.495 172.105 ;
        RECT 112.215 171.795 112.490 171.935 ;
        RECT 112.695 171.595 112.865 172.395 ;
        RECT 111.855 171.425 112.865 171.595 ;
        RECT 113.035 172.385 113.965 172.555 ;
        RECT 114.135 172.385 114.390 172.955 ;
        RECT 114.565 172.400 114.855 173.125 ;
        RECT 115.950 172.415 116.205 172.945 ;
        RECT 116.375 172.665 116.680 173.125 ;
        RECT 116.925 172.745 117.995 172.915 ;
        RECT 113.035 171.255 113.205 172.385 ;
        RECT 113.795 172.215 113.965 172.385 ;
        RECT 112.080 171.085 113.205 171.255 ;
        RECT 113.375 171.885 113.570 172.215 ;
        RECT 113.795 171.885 114.050 172.215 ;
        RECT 113.375 170.915 113.545 171.885 ;
        RECT 114.220 171.715 114.390 172.385 ;
        RECT 115.950 171.765 116.160 172.415 ;
        RECT 116.925 172.390 117.245 172.745 ;
        RECT 116.920 172.215 117.245 172.390 ;
        RECT 116.330 171.915 117.245 172.215 ;
        RECT 117.415 172.175 117.655 172.575 ;
        RECT 117.825 172.515 117.995 172.745 ;
        RECT 118.165 172.685 118.355 173.125 ;
        RECT 118.525 172.675 119.475 172.955 ;
        RECT 119.695 172.765 120.045 172.935 ;
        RECT 117.825 172.345 118.355 172.515 ;
        RECT 116.330 171.885 117.070 171.915 ;
        RECT 111.515 170.745 113.545 170.915 ;
        RECT 113.715 170.575 113.885 171.715 ;
        RECT 114.055 170.745 114.390 171.715 ;
        RECT 114.565 170.575 114.855 171.740 ;
        RECT 115.950 170.885 116.205 171.765 ;
        RECT 116.375 170.575 116.680 171.715 ;
        RECT 116.900 171.295 117.070 171.885 ;
        RECT 117.415 171.805 117.955 172.175 ;
        RECT 118.135 172.065 118.355 172.345 ;
        RECT 118.525 171.895 118.695 172.675 ;
        RECT 118.290 171.725 118.695 171.895 ;
        RECT 118.865 171.885 119.215 172.505 ;
        RECT 118.290 171.635 118.460 171.725 ;
        RECT 119.385 171.715 119.595 172.505 ;
        RECT 117.240 171.465 118.460 171.635 ;
        RECT 118.920 171.555 119.595 171.715 ;
        RECT 116.900 171.125 117.700 171.295 ;
        RECT 117.020 170.575 117.350 170.955 ;
        RECT 117.530 170.835 117.700 171.125 ;
        RECT 118.290 171.085 118.460 171.465 ;
        RECT 118.630 171.545 119.595 171.555 ;
        RECT 119.785 172.375 120.045 172.765 ;
        RECT 120.255 172.665 120.585 173.125 ;
        RECT 121.460 172.735 122.315 172.905 ;
        RECT 122.520 172.735 123.015 172.905 ;
        RECT 123.185 172.765 123.515 173.125 ;
        RECT 119.785 171.685 119.955 172.375 ;
        RECT 120.125 172.025 120.295 172.205 ;
        RECT 120.465 172.195 121.255 172.445 ;
        RECT 121.460 172.025 121.630 172.735 ;
        RECT 121.800 172.225 122.155 172.445 ;
        RECT 120.125 171.855 121.815 172.025 ;
        RECT 118.630 171.255 119.090 171.545 ;
        RECT 119.785 171.515 121.285 171.685 ;
        RECT 119.785 171.375 119.955 171.515 ;
        RECT 119.395 171.205 119.955 171.375 ;
        RECT 117.870 170.575 118.120 171.035 ;
        RECT 118.290 170.745 119.160 171.085 ;
        RECT 119.395 170.745 119.565 171.205 ;
        RECT 120.400 171.175 121.475 171.345 ;
        RECT 119.735 170.575 120.105 171.035 ;
        RECT 120.400 170.835 120.570 171.175 ;
        RECT 120.740 170.575 121.070 171.005 ;
        RECT 121.305 170.835 121.475 171.175 ;
        RECT 121.645 171.075 121.815 171.855 ;
        RECT 121.985 171.635 122.155 172.225 ;
        RECT 122.325 171.825 122.675 172.445 ;
        RECT 121.985 171.245 122.450 171.635 ;
        RECT 122.845 171.375 123.015 172.735 ;
        RECT 123.185 171.545 123.645 172.595 ;
        RECT 122.620 171.205 123.015 171.375 ;
        RECT 122.620 171.075 122.790 171.205 ;
        RECT 121.645 170.745 122.325 171.075 ;
        RECT 122.540 170.745 122.790 171.075 ;
        RECT 122.960 170.575 123.210 171.035 ;
        RECT 123.380 170.760 123.705 171.545 ;
        RECT 123.875 170.745 124.045 172.865 ;
        RECT 124.215 172.745 124.545 173.125 ;
        RECT 124.715 172.575 124.970 172.865 ;
        RECT 124.220 172.405 124.970 172.575 ;
        RECT 124.220 171.415 124.450 172.405 ;
        RECT 125.145 172.375 126.355 173.125 ;
        RECT 126.525 172.375 127.735 173.125 ;
        RECT 124.620 171.585 124.970 172.235 ;
        RECT 125.145 171.665 125.665 172.205 ;
        RECT 125.835 171.835 126.355 172.375 ;
        RECT 126.525 171.665 127.045 172.205 ;
        RECT 127.215 171.835 127.735 172.375 ;
        RECT 124.220 171.245 124.970 171.415 ;
        RECT 124.215 170.575 124.545 171.075 ;
        RECT 124.715 170.745 124.970 171.245 ;
        RECT 125.145 170.575 126.355 171.665 ;
        RECT 126.525 170.575 127.735 171.665 ;
        RECT 14.660 170.405 127.820 170.575 ;
        RECT 14.745 169.315 15.955 170.405 ;
        RECT 14.745 168.605 15.265 169.145 ;
        RECT 15.435 168.775 15.955 169.315 ;
        RECT 16.125 169.315 18.715 170.405 ;
        RECT 18.890 169.970 24.235 170.405 ;
        RECT 16.125 168.795 17.335 169.315 ;
        RECT 17.505 168.625 18.715 169.145 ;
        RECT 20.480 168.720 20.830 169.970 ;
        RECT 24.405 169.240 24.695 170.405 ;
        RECT 24.955 169.660 25.225 170.405 ;
        RECT 25.855 170.400 32.130 170.405 ;
        RECT 25.395 169.490 25.685 170.230 ;
        RECT 25.855 169.675 26.110 170.400 ;
        RECT 26.295 169.505 26.555 170.230 ;
        RECT 26.725 169.675 26.970 170.400 ;
        RECT 27.155 169.505 27.415 170.230 ;
        RECT 27.585 169.675 27.830 170.400 ;
        RECT 28.015 169.505 28.275 170.230 ;
        RECT 28.445 169.675 28.690 170.400 ;
        RECT 28.860 169.505 29.120 170.230 ;
        RECT 29.290 169.675 29.550 170.400 ;
        RECT 29.720 169.505 29.980 170.230 ;
        RECT 30.150 169.675 30.410 170.400 ;
        RECT 30.580 169.505 30.840 170.230 ;
        RECT 31.010 169.675 31.270 170.400 ;
        RECT 31.440 169.505 31.700 170.230 ;
        RECT 31.870 169.605 32.130 170.400 ;
        RECT 26.295 169.490 31.700 169.505 ;
        RECT 24.955 169.385 31.700 169.490 ;
        RECT 24.925 169.265 31.700 169.385 ;
        RECT 14.745 167.855 15.955 168.605 ;
        RECT 16.125 167.855 18.715 168.625 ;
        RECT 22.310 168.400 22.650 169.230 ;
        RECT 24.925 169.215 26.120 169.265 ;
        RECT 24.955 168.675 26.120 169.215 ;
        RECT 32.300 169.095 32.550 170.230 ;
        RECT 32.730 169.595 32.990 170.405 ;
        RECT 33.165 169.095 33.410 170.235 ;
        RECT 33.590 169.595 33.885 170.405 ;
        RECT 34.270 169.435 34.600 170.235 ;
        RECT 34.770 169.605 35.100 170.405 ;
        RECT 35.400 169.435 35.730 170.235 ;
        RECT 36.375 169.605 36.625 170.405 ;
        RECT 34.270 169.265 36.705 169.435 ;
        RECT 36.895 169.265 37.065 170.405 ;
        RECT 37.235 169.265 37.575 170.235 ;
        RECT 26.290 168.845 33.410 169.095 ;
        RECT 18.890 167.855 24.235 168.400 ;
        RECT 24.405 167.855 24.695 168.580 ;
        RECT 24.955 168.505 31.700 168.675 ;
        RECT 24.955 167.855 25.255 168.335 ;
        RECT 25.425 168.050 25.685 168.505 ;
        RECT 25.855 167.855 26.115 168.335 ;
        RECT 26.295 168.050 26.555 168.505 ;
        RECT 26.725 167.855 26.975 168.335 ;
        RECT 27.155 168.050 27.415 168.505 ;
        RECT 27.585 167.855 27.835 168.335 ;
        RECT 28.015 168.050 28.275 168.505 ;
        RECT 28.445 167.855 28.690 168.335 ;
        RECT 28.860 168.050 29.135 168.505 ;
        RECT 29.305 167.855 29.550 168.335 ;
        RECT 29.720 168.050 29.980 168.505 ;
        RECT 30.150 167.855 30.410 168.335 ;
        RECT 30.580 168.050 30.840 168.505 ;
        RECT 31.010 167.855 31.270 168.335 ;
        RECT 31.440 168.050 31.700 168.505 ;
        RECT 31.870 167.855 32.130 168.415 ;
        RECT 32.300 168.035 32.550 168.845 ;
        RECT 32.730 167.855 32.990 168.380 ;
        RECT 33.160 168.035 33.410 168.845 ;
        RECT 33.580 168.535 33.895 169.095 ;
        RECT 34.065 168.845 34.415 169.095 ;
        RECT 34.600 168.635 34.770 169.265 ;
        RECT 34.940 168.845 35.270 169.045 ;
        RECT 35.440 168.845 35.770 169.045 ;
        RECT 35.940 168.845 36.360 169.045 ;
        RECT 36.535 169.015 36.705 169.265 ;
        RECT 36.535 168.845 37.230 169.015 ;
        RECT 33.590 167.855 33.895 168.365 ;
        RECT 34.270 168.025 34.770 168.635 ;
        RECT 35.400 168.505 36.625 168.675 ;
        RECT 37.400 168.655 37.575 169.265 ;
        RECT 37.745 169.315 38.955 170.405 ;
        RECT 39.130 169.970 44.475 170.405 ;
        RECT 44.650 169.970 49.995 170.405 ;
        RECT 37.745 168.775 38.265 169.315 ;
        RECT 35.400 168.025 35.730 168.505 ;
        RECT 35.900 167.855 36.125 168.315 ;
        RECT 36.295 168.025 36.625 168.505 ;
        RECT 36.815 167.855 37.065 168.655 ;
        RECT 37.235 168.025 37.575 168.655 ;
        RECT 38.435 168.605 38.955 169.145 ;
        RECT 40.720 168.720 41.070 169.970 ;
        RECT 37.745 167.855 38.955 168.605 ;
        RECT 42.550 168.400 42.890 169.230 ;
        RECT 46.240 168.720 46.590 169.970 ;
        RECT 50.165 169.240 50.455 170.405 ;
        RECT 51.545 169.315 55.055 170.405 ;
        RECT 48.070 168.400 48.410 169.230 ;
        RECT 51.545 168.795 53.235 169.315 ;
        RECT 55.285 169.265 55.495 170.405 ;
        RECT 55.665 169.255 55.995 170.235 ;
        RECT 56.165 169.265 56.395 170.405 ;
        RECT 57.615 169.475 57.785 170.235 ;
        RECT 57.965 169.645 58.295 170.405 ;
        RECT 57.615 169.305 58.280 169.475 ;
        RECT 58.465 169.330 58.735 170.235 ;
        RECT 53.405 168.625 55.055 169.145 ;
        RECT 39.130 167.855 44.475 168.400 ;
        RECT 44.650 167.855 49.995 168.400 ;
        RECT 50.165 167.855 50.455 168.580 ;
        RECT 51.545 167.855 55.055 168.625 ;
        RECT 55.285 167.855 55.495 168.675 ;
        RECT 55.665 168.655 55.915 169.255 ;
        RECT 58.110 169.160 58.280 169.305 ;
        RECT 56.085 168.845 56.415 169.095 ;
        RECT 57.545 168.755 57.875 169.125 ;
        RECT 58.110 168.830 58.395 169.160 ;
        RECT 55.665 168.025 55.995 168.655 ;
        RECT 56.165 167.855 56.395 168.675 ;
        RECT 58.110 168.575 58.280 168.830 ;
        RECT 57.615 168.405 58.280 168.575 ;
        RECT 58.565 168.530 58.735 169.330 ;
        RECT 59.055 169.255 59.385 170.405 ;
        RECT 59.555 169.385 59.725 170.235 ;
        RECT 59.895 169.605 60.225 170.405 ;
        RECT 60.395 169.385 60.565 170.235 ;
        RECT 60.745 169.605 60.985 170.405 ;
        RECT 61.155 169.425 61.485 170.235 ;
        RECT 59.555 169.215 60.565 169.385 ;
        RECT 60.770 169.255 61.485 169.425 ;
        RECT 61.665 169.315 62.875 170.405 ;
        RECT 63.050 169.970 68.395 170.405 ;
        RECT 59.555 168.675 60.050 169.215 ;
        RECT 60.770 169.015 60.940 169.255 ;
        RECT 60.440 168.845 60.940 169.015 ;
        RECT 61.110 168.845 61.490 169.085 ;
        RECT 60.770 168.675 60.940 168.845 ;
        RECT 61.665 168.775 62.185 169.315 ;
        RECT 57.615 168.025 57.785 168.405 ;
        RECT 57.965 167.855 58.295 168.235 ;
        RECT 58.475 168.025 58.735 168.530 ;
        RECT 59.055 167.855 59.385 168.655 ;
        RECT 59.555 168.505 60.565 168.675 ;
        RECT 60.770 168.505 61.405 168.675 ;
        RECT 62.355 168.605 62.875 169.145 ;
        RECT 64.640 168.720 64.990 169.970 ;
        RECT 68.605 169.265 68.835 170.405 ;
        RECT 69.005 169.255 69.335 170.235 ;
        RECT 69.505 169.265 69.715 170.405 ;
        RECT 59.555 168.025 59.725 168.505 ;
        RECT 59.895 167.855 60.225 168.335 ;
        RECT 60.395 168.025 60.565 168.505 ;
        RECT 60.815 167.855 61.055 168.335 ;
        RECT 61.235 168.025 61.405 168.505 ;
        RECT 61.665 167.855 62.875 168.605 ;
        RECT 66.470 168.400 66.810 169.230 ;
        RECT 68.585 168.845 68.915 169.095 ;
        RECT 63.050 167.855 68.395 168.400 ;
        RECT 68.605 167.855 68.835 168.675 ;
        RECT 69.085 168.655 69.335 169.255 ;
        RECT 69.005 168.025 69.335 168.655 ;
        RECT 69.505 167.855 69.715 168.675 ;
        RECT 69.945 168.595 70.205 170.220 ;
        RECT 71.955 169.955 72.285 170.405 ;
        RECT 70.385 169.565 72.995 169.775 ;
        RECT 70.385 168.765 70.605 169.565 ;
        RECT 70.845 168.765 71.145 169.385 ;
        RECT 71.315 168.765 71.645 169.385 ;
        RECT 71.815 168.765 72.135 169.385 ;
        RECT 72.305 168.765 72.655 169.385 ;
        RECT 72.825 168.595 72.995 169.565 ;
        RECT 73.165 169.315 75.755 170.405 ;
        RECT 73.165 168.795 74.375 169.315 ;
        RECT 75.925 169.240 76.215 170.405 ;
        RECT 76.850 169.970 82.195 170.405 ;
        RECT 74.545 168.625 75.755 169.145 ;
        RECT 78.440 168.720 78.790 169.970 ;
        RECT 82.365 169.645 82.880 170.055 ;
        RECT 83.115 169.645 83.285 170.405 ;
        RECT 83.455 170.065 85.485 170.235 ;
        RECT 69.945 168.425 71.785 168.595 ;
        RECT 70.215 167.855 70.545 168.250 ;
        RECT 70.715 168.070 70.915 168.425 ;
        RECT 71.085 167.855 71.415 168.255 ;
        RECT 71.585 168.080 71.785 168.425 ;
        RECT 71.955 167.855 72.285 168.595 ;
        RECT 72.520 168.425 72.995 168.595 ;
        RECT 72.520 168.175 72.690 168.425 ;
        RECT 73.165 167.855 75.755 168.625 ;
        RECT 75.925 167.855 76.215 168.580 ;
        RECT 80.270 168.400 80.610 169.230 ;
        RECT 82.365 168.835 82.705 169.645 ;
        RECT 83.455 169.400 83.625 170.065 ;
        RECT 84.020 169.725 85.145 169.895 ;
        RECT 82.875 169.210 83.625 169.400 ;
        RECT 83.795 169.385 84.805 169.555 ;
        RECT 82.365 168.665 83.595 168.835 ;
        RECT 76.850 167.855 82.195 168.400 ;
        RECT 82.640 168.060 82.885 168.665 ;
        RECT 83.105 167.855 83.615 168.390 ;
        RECT 83.795 168.025 83.985 169.385 ;
        RECT 84.155 168.365 84.430 169.185 ;
        RECT 84.635 168.585 84.805 169.385 ;
        RECT 84.975 168.595 85.145 169.725 ;
        RECT 85.315 169.095 85.485 170.065 ;
        RECT 85.655 169.265 85.825 170.405 ;
        RECT 85.995 169.265 86.330 170.235 ;
        RECT 86.565 169.265 86.775 170.405 ;
        RECT 85.315 168.765 85.510 169.095 ;
        RECT 85.735 168.765 85.990 169.095 ;
        RECT 85.735 168.595 85.905 168.765 ;
        RECT 86.160 168.595 86.330 169.265 ;
        RECT 86.945 169.255 87.275 170.235 ;
        RECT 87.445 169.265 87.675 170.405 ;
        RECT 88.345 169.315 90.015 170.405 ;
        RECT 84.975 168.425 85.905 168.595 ;
        RECT 84.975 168.390 85.150 168.425 ;
        RECT 84.155 168.195 84.435 168.365 ;
        RECT 84.155 168.025 84.430 168.195 ;
        RECT 84.620 168.025 85.150 168.390 ;
        RECT 85.575 167.855 85.905 168.255 ;
        RECT 86.075 168.025 86.330 168.595 ;
        RECT 86.565 167.855 86.775 168.675 ;
        RECT 86.945 168.655 87.195 169.255 ;
        RECT 87.365 168.845 87.695 169.095 ;
        RECT 88.345 168.795 89.095 169.315 ;
        RECT 90.225 169.265 90.455 170.405 ;
        RECT 90.625 169.255 90.955 170.235 ;
        RECT 91.125 169.265 91.335 170.405 ;
        RECT 86.945 168.025 87.275 168.655 ;
        RECT 87.445 167.855 87.675 168.675 ;
        RECT 89.265 168.625 90.015 169.145 ;
        RECT 90.205 168.845 90.535 169.095 ;
        RECT 88.345 167.855 90.015 168.625 ;
        RECT 90.225 167.855 90.455 168.675 ;
        RECT 90.705 168.655 90.955 169.255 ;
        RECT 91.570 169.215 91.825 170.095 ;
        RECT 91.995 169.265 92.300 170.405 ;
        RECT 92.640 170.025 92.970 170.405 ;
        RECT 93.150 169.855 93.320 170.145 ;
        RECT 93.490 169.945 93.740 170.405 ;
        RECT 92.520 169.685 93.320 169.855 ;
        RECT 93.910 169.895 94.780 170.235 ;
        RECT 90.625 168.025 90.955 168.655 ;
        RECT 91.125 167.855 91.335 168.675 ;
        RECT 91.570 168.565 91.780 169.215 ;
        RECT 92.520 169.095 92.690 169.685 ;
        RECT 93.910 169.515 94.080 169.895 ;
        RECT 95.015 169.775 95.185 170.235 ;
        RECT 95.355 169.945 95.725 170.405 ;
        RECT 96.020 169.805 96.190 170.145 ;
        RECT 96.360 169.975 96.690 170.405 ;
        RECT 96.925 169.805 97.095 170.145 ;
        RECT 92.860 169.345 94.080 169.515 ;
        RECT 94.250 169.435 94.710 169.725 ;
        RECT 95.015 169.605 95.575 169.775 ;
        RECT 96.020 169.635 97.095 169.805 ;
        RECT 97.265 169.905 97.945 170.235 ;
        RECT 98.160 169.905 98.410 170.235 ;
        RECT 98.580 169.945 98.830 170.405 ;
        RECT 95.405 169.465 95.575 169.605 ;
        RECT 94.250 169.425 95.215 169.435 ;
        RECT 93.910 169.255 94.080 169.345 ;
        RECT 94.540 169.265 95.215 169.425 ;
        RECT 91.950 169.065 92.690 169.095 ;
        RECT 91.950 168.765 92.865 169.065 ;
        RECT 92.540 168.590 92.865 168.765 ;
        RECT 91.570 168.035 91.825 168.565 ;
        RECT 91.995 167.855 92.300 168.315 ;
        RECT 92.545 168.235 92.865 168.590 ;
        RECT 93.035 168.805 93.575 169.175 ;
        RECT 93.910 169.085 94.315 169.255 ;
        RECT 93.035 168.405 93.275 168.805 ;
        RECT 93.755 168.635 93.975 168.915 ;
        RECT 93.445 168.465 93.975 168.635 ;
        RECT 93.445 168.235 93.615 168.465 ;
        RECT 94.145 168.305 94.315 169.085 ;
        RECT 94.485 168.475 94.835 169.095 ;
        RECT 95.005 168.475 95.215 169.265 ;
        RECT 95.405 169.295 96.905 169.465 ;
        RECT 95.405 168.605 95.575 169.295 ;
        RECT 97.265 169.125 97.435 169.905 ;
        RECT 98.240 169.775 98.410 169.905 ;
        RECT 95.745 168.955 97.435 169.125 ;
        RECT 97.605 169.345 98.070 169.735 ;
        RECT 98.240 169.605 98.635 169.775 ;
        RECT 95.745 168.775 95.915 168.955 ;
        RECT 92.545 168.065 93.615 168.235 ;
        RECT 93.785 167.855 93.975 168.295 ;
        RECT 94.145 168.025 95.095 168.305 ;
        RECT 95.405 168.215 95.665 168.605 ;
        RECT 96.085 168.535 96.875 168.785 ;
        RECT 95.315 168.045 95.665 168.215 ;
        RECT 95.875 167.855 96.205 168.315 ;
        RECT 97.080 168.245 97.250 168.955 ;
        RECT 97.605 168.755 97.775 169.345 ;
        RECT 97.420 168.535 97.775 168.755 ;
        RECT 97.945 168.535 98.295 169.155 ;
        RECT 98.465 168.245 98.635 169.605 ;
        RECT 99.000 169.435 99.325 170.220 ;
        RECT 98.805 168.385 99.265 169.435 ;
        RECT 97.080 168.075 97.935 168.245 ;
        RECT 98.140 168.075 98.635 168.245 ;
        RECT 98.805 167.855 99.135 168.215 ;
        RECT 99.495 168.115 99.665 170.235 ;
        RECT 99.835 169.905 100.165 170.405 ;
        RECT 100.335 169.735 100.590 170.235 ;
        RECT 99.840 169.565 100.590 169.735 ;
        RECT 99.840 168.575 100.070 169.565 ;
        RECT 100.240 168.745 100.590 169.395 ;
        RECT 101.685 169.240 101.975 170.405 ;
        RECT 102.645 169.265 102.875 170.405 ;
        RECT 103.045 169.255 103.375 170.235 ;
        RECT 103.545 169.265 103.755 170.405 ;
        RECT 102.625 168.845 102.955 169.095 ;
        RECT 99.840 168.405 100.590 168.575 ;
        RECT 99.835 167.855 100.165 168.235 ;
        RECT 100.335 168.115 100.590 168.405 ;
        RECT 101.685 167.855 101.975 168.580 ;
        RECT 102.645 167.855 102.875 168.675 ;
        RECT 103.125 168.655 103.375 169.255 ;
        RECT 103.990 169.215 104.245 170.095 ;
        RECT 104.415 169.265 104.720 170.405 ;
        RECT 105.060 170.025 105.390 170.405 ;
        RECT 105.570 169.855 105.740 170.145 ;
        RECT 105.910 169.945 106.160 170.405 ;
        RECT 104.940 169.685 105.740 169.855 ;
        RECT 106.330 169.895 107.200 170.235 ;
        RECT 103.045 168.025 103.375 168.655 ;
        RECT 103.545 167.855 103.755 168.675 ;
        RECT 103.990 168.565 104.200 169.215 ;
        RECT 104.940 169.095 105.110 169.685 ;
        RECT 106.330 169.515 106.500 169.895 ;
        RECT 107.435 169.775 107.605 170.235 ;
        RECT 107.775 169.945 108.145 170.405 ;
        RECT 108.440 169.805 108.610 170.145 ;
        RECT 108.780 169.975 109.110 170.405 ;
        RECT 109.345 169.805 109.515 170.145 ;
        RECT 105.280 169.345 106.500 169.515 ;
        RECT 106.670 169.435 107.130 169.725 ;
        RECT 107.435 169.605 107.995 169.775 ;
        RECT 108.440 169.635 109.515 169.805 ;
        RECT 109.685 169.905 110.365 170.235 ;
        RECT 110.580 169.905 110.830 170.235 ;
        RECT 111.000 169.945 111.250 170.405 ;
        RECT 107.825 169.465 107.995 169.605 ;
        RECT 106.670 169.425 107.635 169.435 ;
        RECT 106.330 169.255 106.500 169.345 ;
        RECT 106.960 169.265 107.635 169.425 ;
        RECT 104.370 169.065 105.110 169.095 ;
        RECT 104.370 168.765 105.285 169.065 ;
        RECT 104.960 168.590 105.285 168.765 ;
        RECT 103.990 168.035 104.245 168.565 ;
        RECT 104.415 167.855 104.720 168.315 ;
        RECT 104.965 168.235 105.285 168.590 ;
        RECT 105.455 168.805 105.995 169.175 ;
        RECT 106.330 169.085 106.735 169.255 ;
        RECT 105.455 168.405 105.695 168.805 ;
        RECT 106.175 168.635 106.395 168.915 ;
        RECT 105.865 168.465 106.395 168.635 ;
        RECT 105.865 168.235 106.035 168.465 ;
        RECT 106.565 168.305 106.735 169.085 ;
        RECT 106.905 168.475 107.255 169.095 ;
        RECT 107.425 168.475 107.635 169.265 ;
        RECT 107.825 169.295 109.325 169.465 ;
        RECT 107.825 168.605 107.995 169.295 ;
        RECT 109.685 169.125 109.855 169.905 ;
        RECT 110.660 169.775 110.830 169.905 ;
        RECT 108.165 168.955 109.855 169.125 ;
        RECT 110.025 169.345 110.490 169.735 ;
        RECT 110.660 169.605 111.055 169.775 ;
        RECT 108.165 168.775 108.335 168.955 ;
        RECT 104.965 168.065 106.035 168.235 ;
        RECT 106.205 167.855 106.395 168.295 ;
        RECT 106.565 168.025 107.515 168.305 ;
        RECT 107.825 168.215 108.085 168.605 ;
        RECT 108.505 168.535 109.295 168.785 ;
        RECT 107.735 168.045 108.085 168.215 ;
        RECT 108.295 167.855 108.625 168.315 ;
        RECT 109.500 168.245 109.670 168.955 ;
        RECT 110.025 168.755 110.195 169.345 ;
        RECT 109.840 168.535 110.195 168.755 ;
        RECT 110.365 168.535 110.715 169.155 ;
        RECT 110.885 168.245 111.055 169.605 ;
        RECT 111.420 169.435 111.745 170.220 ;
        RECT 111.225 168.385 111.685 169.435 ;
        RECT 109.500 168.075 110.355 168.245 ;
        RECT 110.560 168.075 111.055 168.245 ;
        RECT 111.225 167.855 111.555 168.215 ;
        RECT 111.915 168.115 112.085 170.235 ;
        RECT 112.255 169.905 112.585 170.405 ;
        RECT 112.755 169.735 113.010 170.235 ;
        RECT 112.260 169.565 113.010 169.735 ;
        RECT 112.260 168.575 112.490 169.565 ;
        RECT 112.660 168.745 113.010 169.395 ;
        RECT 113.185 169.315 114.855 170.405 ;
        RECT 115.030 169.970 120.375 170.405 ;
        RECT 113.185 168.795 113.935 169.315 ;
        RECT 114.105 168.625 114.855 169.145 ;
        RECT 116.620 168.720 116.970 169.970 ;
        RECT 120.635 169.475 120.805 170.235 ;
        RECT 120.985 169.645 121.315 170.405 ;
        RECT 120.635 169.305 121.300 169.475 ;
        RECT 121.485 169.330 121.755 170.235 ;
        RECT 121.930 169.980 122.265 170.405 ;
        RECT 122.435 169.800 122.620 170.205 ;
        RECT 112.260 168.405 113.010 168.575 ;
        RECT 112.255 167.855 112.585 168.235 ;
        RECT 112.755 168.115 113.010 168.405 ;
        RECT 113.185 167.855 114.855 168.625 ;
        RECT 118.450 168.400 118.790 169.230 ;
        RECT 121.130 169.160 121.300 169.305 ;
        RECT 120.565 168.755 120.895 169.125 ;
        RECT 121.130 168.830 121.415 169.160 ;
        RECT 121.130 168.575 121.300 168.830 ;
        RECT 120.635 168.405 121.300 168.575 ;
        RECT 121.585 168.530 121.755 169.330 ;
        RECT 115.030 167.855 120.375 168.400 ;
        RECT 120.635 168.025 120.805 168.405 ;
        RECT 120.985 167.855 121.315 168.235 ;
        RECT 121.495 168.025 121.755 168.530 ;
        RECT 121.955 169.625 122.620 169.800 ;
        RECT 122.825 169.625 123.155 170.405 ;
        RECT 121.955 168.595 122.295 169.625 ;
        RECT 123.325 169.435 123.595 170.205 ;
        RECT 122.465 169.265 123.595 169.435 ;
        RECT 122.465 168.765 122.715 169.265 ;
        RECT 121.955 168.425 122.640 168.595 ;
        RECT 122.895 168.515 123.255 169.095 ;
        RECT 121.930 167.855 122.265 168.255 ;
        RECT 122.435 168.025 122.640 168.425 ;
        RECT 123.425 168.355 123.595 169.265 ;
        RECT 123.765 169.315 126.355 170.405 ;
        RECT 126.525 169.315 127.735 170.405 ;
        RECT 123.765 168.795 124.975 169.315 ;
        RECT 125.145 168.625 126.355 169.145 ;
        RECT 126.525 168.775 127.045 169.315 ;
        RECT 122.850 167.855 123.125 168.335 ;
        RECT 123.335 168.025 123.595 168.355 ;
        RECT 123.765 167.855 126.355 168.625 ;
        RECT 127.215 168.605 127.735 169.145 ;
        RECT 126.525 167.855 127.735 168.605 ;
        RECT 14.660 167.685 127.820 167.855 ;
        RECT 14.745 166.935 15.955 167.685 ;
        RECT 16.500 166.975 16.755 167.505 ;
        RECT 16.935 167.225 17.220 167.685 ;
        RECT 14.745 166.395 15.265 166.935 ;
        RECT 15.435 166.225 15.955 166.765 ;
        RECT 14.745 165.135 15.955 166.225 ;
        RECT 16.500 166.115 16.680 166.975 ;
        RECT 17.400 166.775 17.650 167.425 ;
        RECT 16.850 166.445 17.650 166.775 ;
        RECT 16.500 165.645 16.755 166.115 ;
        RECT 16.415 165.475 16.755 165.645 ;
        RECT 16.500 165.445 16.755 165.475 ;
        RECT 16.935 165.135 17.220 165.935 ;
        RECT 17.400 165.855 17.650 166.445 ;
        RECT 17.850 167.090 18.170 167.420 ;
        RECT 18.350 167.205 19.010 167.685 ;
        RECT 19.210 167.295 20.060 167.465 ;
        RECT 17.850 166.195 18.040 167.090 ;
        RECT 18.360 166.765 19.020 167.035 ;
        RECT 18.690 166.705 19.020 166.765 ;
        RECT 18.210 166.535 18.540 166.595 ;
        RECT 19.210 166.535 19.380 167.295 ;
        RECT 20.620 167.225 20.940 167.685 ;
        RECT 21.140 167.045 21.390 167.475 ;
        RECT 21.680 167.245 22.090 167.685 ;
        RECT 22.260 167.305 23.275 167.505 ;
        RECT 19.550 166.875 20.800 167.045 ;
        RECT 19.550 166.755 19.880 166.875 ;
        RECT 18.210 166.365 20.110 166.535 ;
        RECT 17.850 166.025 19.770 166.195 ;
        RECT 17.850 166.005 18.170 166.025 ;
        RECT 17.400 165.345 17.730 165.855 ;
        RECT 18.000 165.395 18.170 166.005 ;
        RECT 19.940 165.855 20.110 166.365 ;
        RECT 20.280 166.295 20.460 166.705 ;
        RECT 20.630 166.115 20.800 166.875 ;
        RECT 18.340 165.135 18.670 165.825 ;
        RECT 18.900 165.685 20.110 165.855 ;
        RECT 20.280 165.805 20.800 166.115 ;
        RECT 20.970 166.705 21.390 167.045 ;
        RECT 21.680 166.705 22.090 167.035 ;
        RECT 20.970 165.935 21.160 166.705 ;
        RECT 22.260 166.575 22.430 167.305 ;
        RECT 23.575 167.135 23.745 167.465 ;
        RECT 23.915 167.305 24.245 167.685 ;
        RECT 22.600 166.755 22.950 167.125 ;
        RECT 22.260 166.535 22.680 166.575 ;
        RECT 21.330 166.365 22.680 166.535 ;
        RECT 21.330 166.205 21.580 166.365 ;
        RECT 22.090 165.935 22.340 166.195 ;
        RECT 20.970 165.685 22.340 165.935 ;
        RECT 18.900 165.395 19.140 165.685 ;
        RECT 19.940 165.605 20.110 165.685 ;
        RECT 19.340 165.135 19.760 165.515 ;
        RECT 19.940 165.355 20.570 165.605 ;
        RECT 21.040 165.135 21.370 165.515 ;
        RECT 21.540 165.395 21.710 165.685 ;
        RECT 22.510 165.520 22.680 166.365 ;
        RECT 23.130 166.195 23.350 167.065 ;
        RECT 23.575 166.945 24.270 167.135 ;
        RECT 22.850 165.815 23.350 166.195 ;
        RECT 23.520 166.145 23.930 166.765 ;
        RECT 24.100 165.975 24.270 166.945 ;
        RECT 23.575 165.805 24.270 165.975 ;
        RECT 21.890 165.135 22.270 165.515 ;
        RECT 22.510 165.350 23.340 165.520 ;
        RECT 23.575 165.305 23.745 165.805 ;
        RECT 23.915 165.135 24.245 165.635 ;
        RECT 24.460 165.305 24.685 167.425 ;
        RECT 24.855 167.305 25.185 167.685 ;
        RECT 25.355 167.135 25.525 167.425 ;
        RECT 26.250 167.140 31.595 167.685 ;
        RECT 31.770 167.140 37.115 167.685 ;
        RECT 24.860 166.965 25.525 167.135 ;
        RECT 24.860 165.975 25.090 166.965 ;
        RECT 25.260 166.145 25.610 166.795 ;
        RECT 24.860 165.805 25.525 165.975 ;
        RECT 24.855 165.135 25.185 165.635 ;
        RECT 25.355 165.305 25.525 165.805 ;
        RECT 27.840 165.570 28.190 166.820 ;
        RECT 29.670 166.310 30.010 167.140 ;
        RECT 33.360 165.570 33.710 166.820 ;
        RECT 35.190 166.310 35.530 167.140 ;
        RECT 37.285 166.960 37.575 167.685 ;
        RECT 38.205 166.915 40.795 167.685 ;
        RECT 40.970 167.140 46.315 167.685 ;
        RECT 46.490 167.140 51.835 167.685 ;
        RECT 26.250 165.135 31.595 165.570 ;
        RECT 31.770 165.135 37.115 165.570 ;
        RECT 37.285 165.135 37.575 166.300 ;
        RECT 38.205 166.225 39.415 166.745 ;
        RECT 39.585 166.395 40.795 166.915 ;
        RECT 38.205 165.135 40.795 166.225 ;
        RECT 42.560 165.570 42.910 166.820 ;
        RECT 44.390 166.310 44.730 167.140 ;
        RECT 48.080 165.570 48.430 166.820 ;
        RECT 49.910 166.310 50.250 167.140 ;
        RECT 52.010 166.975 52.265 167.505 ;
        RECT 52.435 167.225 52.740 167.685 ;
        RECT 52.985 167.305 54.055 167.475 ;
        RECT 52.010 166.325 52.220 166.975 ;
        RECT 52.985 166.950 53.305 167.305 ;
        RECT 52.980 166.775 53.305 166.950 ;
        RECT 52.390 166.475 53.305 166.775 ;
        RECT 53.475 166.735 53.715 167.135 ;
        RECT 53.885 167.075 54.055 167.305 ;
        RECT 54.225 167.245 54.415 167.685 ;
        RECT 54.585 167.235 55.535 167.515 ;
        RECT 55.755 167.325 56.105 167.495 ;
        RECT 53.885 166.905 54.415 167.075 ;
        RECT 52.390 166.445 53.130 166.475 ;
        RECT 40.970 165.135 46.315 165.570 ;
        RECT 46.490 165.135 51.835 165.570 ;
        RECT 52.010 165.445 52.265 166.325 ;
        RECT 52.435 165.135 52.740 166.275 ;
        RECT 52.960 165.855 53.130 166.445 ;
        RECT 53.475 166.365 54.015 166.735 ;
        RECT 54.195 166.625 54.415 166.905 ;
        RECT 54.585 166.455 54.755 167.235 ;
        RECT 54.350 166.285 54.755 166.455 ;
        RECT 54.925 166.445 55.275 167.065 ;
        RECT 54.350 166.195 54.520 166.285 ;
        RECT 55.445 166.275 55.655 167.065 ;
        RECT 53.300 166.025 54.520 166.195 ;
        RECT 54.980 166.115 55.655 166.275 ;
        RECT 52.960 165.685 53.760 165.855 ;
        RECT 53.080 165.135 53.410 165.515 ;
        RECT 53.590 165.395 53.760 165.685 ;
        RECT 54.350 165.645 54.520 166.025 ;
        RECT 54.690 166.105 55.655 166.115 ;
        RECT 55.845 166.935 56.105 167.325 ;
        RECT 56.315 167.225 56.645 167.685 ;
        RECT 57.520 167.295 58.375 167.465 ;
        RECT 58.580 167.295 59.075 167.465 ;
        RECT 59.245 167.325 59.575 167.685 ;
        RECT 55.845 166.245 56.015 166.935 ;
        RECT 56.185 166.585 56.355 166.765 ;
        RECT 56.525 166.755 57.315 167.005 ;
        RECT 57.520 166.585 57.690 167.295 ;
        RECT 57.860 166.785 58.215 167.005 ;
        RECT 56.185 166.415 57.875 166.585 ;
        RECT 54.690 165.815 55.150 166.105 ;
        RECT 55.845 166.075 57.345 166.245 ;
        RECT 55.845 165.935 56.015 166.075 ;
        RECT 55.455 165.765 56.015 165.935 ;
        RECT 53.930 165.135 54.180 165.595 ;
        RECT 54.350 165.305 55.220 165.645 ;
        RECT 55.455 165.305 55.625 165.765 ;
        RECT 56.460 165.735 57.535 165.905 ;
        RECT 55.795 165.135 56.165 165.595 ;
        RECT 56.460 165.395 56.630 165.735 ;
        RECT 56.800 165.135 57.130 165.565 ;
        RECT 57.365 165.395 57.535 165.735 ;
        RECT 57.705 165.635 57.875 166.415 ;
        RECT 58.045 166.195 58.215 166.785 ;
        RECT 58.385 166.385 58.735 167.005 ;
        RECT 58.045 165.805 58.510 166.195 ;
        RECT 58.905 165.935 59.075 167.295 ;
        RECT 59.245 166.105 59.705 167.155 ;
        RECT 58.680 165.765 59.075 165.935 ;
        RECT 58.680 165.635 58.850 165.765 ;
        RECT 57.705 165.305 58.385 165.635 ;
        RECT 58.600 165.305 58.850 165.635 ;
        RECT 59.020 165.135 59.270 165.595 ;
        RECT 59.440 165.320 59.765 166.105 ;
        RECT 59.935 165.305 60.105 167.425 ;
        RECT 60.275 167.305 60.605 167.685 ;
        RECT 60.775 167.135 61.030 167.425 ;
        RECT 60.280 166.965 61.030 167.135 ;
        RECT 60.280 165.975 60.510 166.965 ;
        RECT 61.205 166.915 62.875 167.685 ;
        RECT 63.045 166.960 63.335 167.685 ;
        RECT 63.505 166.935 64.715 167.685 ;
        RECT 64.890 167.140 70.235 167.685 ;
        RECT 60.680 166.145 61.030 166.795 ;
        RECT 61.205 166.225 61.955 166.745 ;
        RECT 62.125 166.395 62.875 166.915 ;
        RECT 60.280 165.805 61.030 165.975 ;
        RECT 60.275 165.135 60.605 165.635 ;
        RECT 60.775 165.305 61.030 165.805 ;
        RECT 61.205 165.135 62.875 166.225 ;
        RECT 63.045 165.135 63.335 166.300 ;
        RECT 63.505 166.225 64.025 166.765 ;
        RECT 64.195 166.395 64.715 166.935 ;
        RECT 63.505 165.135 64.715 166.225 ;
        RECT 66.480 165.570 66.830 166.820 ;
        RECT 68.310 166.310 68.650 167.140 ;
        RECT 70.410 166.845 70.670 167.685 ;
        RECT 70.845 166.940 71.100 167.515 ;
        RECT 71.270 167.305 71.600 167.685 ;
        RECT 71.815 167.135 71.985 167.515 ;
        RECT 71.270 166.965 71.985 167.135 ;
        RECT 64.890 165.135 70.235 165.570 ;
        RECT 70.410 165.135 70.670 166.285 ;
        RECT 70.845 166.210 71.015 166.940 ;
        RECT 71.270 166.775 71.440 166.965 ;
        RECT 72.245 166.935 73.455 167.685 ;
        RECT 73.630 167.140 78.975 167.685 ;
        RECT 71.185 166.445 71.440 166.775 ;
        RECT 71.270 166.235 71.440 166.445 ;
        RECT 71.720 166.415 72.075 166.785 ;
        RECT 70.845 165.305 71.100 166.210 ;
        RECT 71.270 166.065 71.985 166.235 ;
        RECT 71.270 165.135 71.600 165.895 ;
        RECT 71.815 165.305 71.985 166.065 ;
        RECT 72.245 166.225 72.765 166.765 ;
        RECT 72.935 166.395 73.455 166.935 ;
        RECT 72.245 165.135 73.455 166.225 ;
        RECT 75.220 165.570 75.570 166.820 ;
        RECT 77.050 166.310 77.390 167.140 ;
        RECT 79.235 167.135 79.405 167.425 ;
        RECT 79.575 167.305 79.905 167.685 ;
        RECT 79.235 166.965 79.900 167.135 ;
        RECT 79.150 166.145 79.500 166.795 ;
        RECT 79.670 165.975 79.900 166.965 ;
        RECT 79.235 165.805 79.900 165.975 ;
        RECT 73.630 165.135 78.975 165.570 ;
        RECT 79.235 165.305 79.405 165.805 ;
        RECT 79.575 165.135 79.905 165.635 ;
        RECT 80.075 165.305 80.300 167.425 ;
        RECT 80.515 167.305 80.845 167.685 ;
        RECT 81.015 167.135 81.185 167.465 ;
        RECT 81.485 167.305 82.500 167.505 ;
        RECT 80.490 166.945 81.185 167.135 ;
        RECT 80.490 165.975 80.660 166.945 ;
        RECT 80.830 166.145 81.240 166.765 ;
        RECT 81.410 166.195 81.630 167.065 ;
        RECT 81.810 166.755 82.160 167.125 ;
        RECT 82.330 166.575 82.500 167.305 ;
        RECT 82.670 167.245 83.080 167.685 ;
        RECT 83.370 167.045 83.620 167.475 ;
        RECT 83.820 167.225 84.140 167.685 ;
        RECT 84.700 167.295 85.550 167.465 ;
        RECT 82.670 166.705 83.080 167.035 ;
        RECT 83.370 166.705 83.790 167.045 ;
        RECT 82.080 166.535 82.500 166.575 ;
        RECT 82.080 166.365 83.430 166.535 ;
        RECT 80.490 165.805 81.185 165.975 ;
        RECT 81.410 165.815 81.910 166.195 ;
        RECT 80.515 165.135 80.845 165.635 ;
        RECT 81.015 165.305 81.185 165.805 ;
        RECT 82.080 165.520 82.250 166.365 ;
        RECT 83.180 166.205 83.430 166.365 ;
        RECT 82.420 165.935 82.670 166.195 ;
        RECT 83.600 165.935 83.790 166.705 ;
        RECT 82.420 165.685 83.790 165.935 ;
        RECT 83.960 166.875 85.210 167.045 ;
        RECT 83.960 166.115 84.130 166.875 ;
        RECT 84.880 166.755 85.210 166.875 ;
        RECT 84.300 166.295 84.480 166.705 ;
        RECT 85.380 166.535 85.550 167.295 ;
        RECT 85.750 167.205 86.410 167.685 ;
        RECT 86.590 167.090 86.910 167.420 ;
        RECT 85.740 166.765 86.400 167.035 ;
        RECT 85.740 166.705 86.070 166.765 ;
        RECT 86.220 166.535 86.550 166.595 ;
        RECT 84.650 166.365 86.550 166.535 ;
        RECT 83.960 165.805 84.480 166.115 ;
        RECT 84.650 165.855 84.820 166.365 ;
        RECT 86.720 166.195 86.910 167.090 ;
        RECT 84.990 166.025 86.910 166.195 ;
        RECT 86.590 166.005 86.910 166.025 ;
        RECT 87.110 166.775 87.360 167.425 ;
        RECT 87.540 167.225 87.825 167.685 ;
        RECT 88.005 167.005 88.260 167.505 ;
        RECT 88.005 166.975 88.345 167.005 ;
        RECT 88.080 166.835 88.345 166.975 ;
        RECT 88.805 166.960 89.095 167.685 ;
        RECT 89.265 167.010 89.525 167.515 ;
        RECT 89.705 167.305 90.035 167.685 ;
        RECT 90.215 167.135 90.385 167.515 ;
        RECT 87.110 166.445 87.910 166.775 ;
        RECT 84.650 165.685 85.860 165.855 ;
        RECT 81.420 165.350 82.250 165.520 ;
        RECT 82.490 165.135 82.870 165.515 ;
        RECT 83.050 165.395 83.220 165.685 ;
        RECT 84.650 165.605 84.820 165.685 ;
        RECT 83.390 165.135 83.720 165.515 ;
        RECT 84.190 165.355 84.820 165.605 ;
        RECT 85.000 165.135 85.420 165.515 ;
        RECT 85.620 165.395 85.860 165.685 ;
        RECT 86.090 165.135 86.420 165.825 ;
        RECT 86.590 165.395 86.760 166.005 ;
        RECT 87.110 165.855 87.360 166.445 ;
        RECT 88.080 166.115 88.260 166.835 ;
        RECT 87.030 165.345 87.360 165.855 ;
        RECT 87.540 165.135 87.825 165.935 ;
        RECT 88.005 165.445 88.260 166.115 ;
        RECT 88.805 165.135 89.095 166.300 ;
        RECT 89.265 166.210 89.435 167.010 ;
        RECT 89.720 166.965 90.385 167.135 ;
        RECT 89.720 166.710 89.890 166.965 ;
        RECT 91.840 166.875 92.085 167.480 ;
        RECT 92.305 167.150 92.815 167.685 ;
        RECT 89.605 166.380 89.890 166.710 ;
        RECT 90.125 166.415 90.455 166.785 ;
        RECT 91.565 166.705 92.795 166.875 ;
        RECT 89.720 166.235 89.890 166.380 ;
        RECT 89.265 165.305 89.535 166.210 ;
        RECT 89.720 166.065 90.385 166.235 ;
        RECT 89.705 165.135 90.035 165.895 ;
        RECT 90.215 165.305 90.385 166.065 ;
        RECT 91.565 165.895 91.905 166.705 ;
        RECT 92.075 166.140 92.825 166.330 ;
        RECT 91.565 165.485 92.080 165.895 ;
        RECT 92.315 165.135 92.485 165.895 ;
        RECT 92.655 165.475 92.825 166.140 ;
        RECT 92.995 166.155 93.185 167.515 ;
        RECT 93.355 167.005 93.630 167.515 ;
        RECT 93.820 167.150 94.350 167.515 ;
        RECT 94.775 167.285 95.105 167.685 ;
        RECT 94.175 167.115 94.350 167.150 ;
        RECT 93.355 166.835 93.635 167.005 ;
        RECT 93.355 166.355 93.630 166.835 ;
        RECT 93.835 166.155 94.005 166.955 ;
        RECT 92.995 165.985 94.005 166.155 ;
        RECT 94.175 166.945 95.105 167.115 ;
        RECT 95.275 166.945 95.530 167.515 ;
        RECT 94.175 165.815 94.345 166.945 ;
        RECT 94.935 166.775 95.105 166.945 ;
        RECT 93.220 165.645 94.345 165.815 ;
        RECT 94.515 166.445 94.710 166.775 ;
        RECT 94.935 166.445 95.190 166.775 ;
        RECT 94.515 165.475 94.685 166.445 ;
        RECT 95.360 166.275 95.530 166.945 ;
        RECT 95.705 166.935 96.915 167.685 ;
        RECT 97.090 167.140 102.435 167.685 ;
        RECT 92.655 165.305 94.685 165.475 ;
        RECT 94.855 165.135 95.025 166.275 ;
        RECT 95.195 165.305 95.530 166.275 ;
        RECT 95.705 166.225 96.225 166.765 ;
        RECT 96.395 166.395 96.915 166.935 ;
        RECT 95.705 165.135 96.915 166.225 ;
        RECT 98.680 165.570 99.030 166.820 ;
        RECT 100.510 166.310 100.850 167.140 ;
        RECT 102.880 166.875 103.125 167.480 ;
        RECT 103.345 167.150 103.855 167.685 ;
        RECT 102.605 166.705 103.835 166.875 ;
        RECT 102.605 165.895 102.945 166.705 ;
        RECT 103.115 166.140 103.865 166.330 ;
        RECT 97.090 165.135 102.435 165.570 ;
        RECT 102.605 165.485 103.120 165.895 ;
        RECT 103.355 165.135 103.525 165.895 ;
        RECT 103.695 165.475 103.865 166.140 ;
        RECT 104.035 166.155 104.225 167.515 ;
        RECT 104.395 166.665 104.670 167.515 ;
        RECT 104.860 167.150 105.390 167.515 ;
        RECT 105.815 167.285 106.145 167.685 ;
        RECT 105.215 167.115 105.390 167.150 ;
        RECT 104.395 166.495 104.675 166.665 ;
        RECT 104.395 166.355 104.670 166.495 ;
        RECT 104.875 166.155 105.045 166.955 ;
        RECT 104.035 165.985 105.045 166.155 ;
        RECT 105.215 166.945 106.145 167.115 ;
        RECT 106.315 166.945 106.570 167.515 ;
        RECT 105.215 165.815 105.385 166.945 ;
        RECT 105.975 166.775 106.145 166.945 ;
        RECT 104.260 165.645 105.385 165.815 ;
        RECT 105.555 166.445 105.750 166.775 ;
        RECT 105.975 166.445 106.230 166.775 ;
        RECT 105.555 165.475 105.725 166.445 ;
        RECT 106.400 166.275 106.570 166.945 ;
        RECT 107.480 166.875 107.725 167.480 ;
        RECT 107.945 167.150 108.455 167.685 ;
        RECT 103.695 165.305 105.725 165.475 ;
        RECT 105.895 165.135 106.065 166.275 ;
        RECT 106.235 165.305 106.570 166.275 ;
        RECT 107.205 166.705 108.435 166.875 ;
        RECT 107.205 165.895 107.545 166.705 ;
        RECT 107.715 166.140 108.465 166.330 ;
        RECT 107.205 165.485 107.720 165.895 ;
        RECT 107.955 165.135 108.125 165.895 ;
        RECT 108.295 165.475 108.465 166.140 ;
        RECT 108.635 166.155 108.825 167.515 ;
        RECT 108.995 166.665 109.270 167.515 ;
        RECT 109.460 167.150 109.990 167.515 ;
        RECT 110.415 167.285 110.745 167.685 ;
        RECT 109.815 167.115 109.990 167.150 ;
        RECT 108.995 166.495 109.275 166.665 ;
        RECT 108.995 166.355 109.270 166.495 ;
        RECT 109.475 166.155 109.645 166.955 ;
        RECT 108.635 165.985 109.645 166.155 ;
        RECT 109.815 166.945 110.745 167.115 ;
        RECT 110.915 166.945 111.170 167.515 ;
        RECT 109.815 165.815 109.985 166.945 ;
        RECT 110.575 166.775 110.745 166.945 ;
        RECT 108.860 165.645 109.985 165.815 ;
        RECT 110.155 166.445 110.350 166.775 ;
        RECT 110.575 166.445 110.830 166.775 ;
        RECT 110.155 165.475 110.325 166.445 ;
        RECT 111.000 166.275 111.170 166.945 ;
        RECT 108.295 165.305 110.325 165.475 ;
        RECT 110.495 165.135 110.665 166.275 ;
        RECT 110.835 165.305 111.170 166.275 ;
        RECT 111.345 167.010 111.605 167.515 ;
        RECT 111.785 167.305 112.115 167.685 ;
        RECT 112.295 167.135 112.465 167.515 ;
        RECT 111.345 166.210 111.515 167.010 ;
        RECT 111.800 166.965 112.465 167.135 ;
        RECT 111.800 166.710 111.970 166.965 ;
        RECT 112.725 166.915 114.395 167.685 ;
        RECT 114.565 166.960 114.855 167.685 ;
        RECT 111.685 166.380 111.970 166.710 ;
        RECT 112.205 166.415 112.535 166.785 ;
        RECT 111.800 166.235 111.970 166.380 ;
        RECT 111.345 165.305 111.615 166.210 ;
        RECT 111.800 166.065 112.465 166.235 ;
        RECT 111.785 165.135 112.115 165.895 ;
        RECT 112.295 165.305 112.465 166.065 ;
        RECT 112.725 166.225 113.475 166.745 ;
        RECT 113.645 166.395 114.395 166.915 ;
        RECT 115.300 166.875 115.545 167.480 ;
        RECT 115.765 167.150 116.275 167.685 ;
        RECT 115.025 166.705 116.255 166.875 ;
        RECT 112.725 165.135 114.395 166.225 ;
        RECT 114.565 165.135 114.855 166.300 ;
        RECT 115.025 165.895 115.365 166.705 ;
        RECT 115.535 166.140 116.285 166.330 ;
        RECT 115.025 165.485 115.540 165.895 ;
        RECT 115.775 165.135 115.945 165.895 ;
        RECT 116.115 165.475 116.285 166.140 ;
        RECT 116.455 166.155 116.645 167.515 ;
        RECT 116.815 166.665 117.090 167.515 ;
        RECT 117.280 167.150 117.810 167.515 ;
        RECT 118.235 167.285 118.565 167.685 ;
        RECT 117.635 167.115 117.810 167.150 ;
        RECT 116.815 166.495 117.095 166.665 ;
        RECT 116.815 166.355 117.090 166.495 ;
        RECT 117.295 166.155 117.465 166.955 ;
        RECT 116.455 165.985 117.465 166.155 ;
        RECT 117.635 166.945 118.565 167.115 ;
        RECT 118.735 166.945 118.990 167.515 ;
        RECT 117.635 165.815 117.805 166.945 ;
        RECT 118.395 166.775 118.565 166.945 ;
        RECT 116.680 165.645 117.805 165.815 ;
        RECT 117.975 166.445 118.170 166.775 ;
        RECT 118.395 166.445 118.650 166.775 ;
        RECT 117.975 165.475 118.145 166.445 ;
        RECT 118.820 166.275 118.990 166.945 ;
        RECT 119.205 166.865 119.435 167.685 ;
        RECT 119.605 166.885 119.935 167.515 ;
        RECT 119.185 166.445 119.515 166.695 ;
        RECT 119.685 166.285 119.935 166.885 ;
        RECT 120.105 166.865 120.315 167.685 ;
        RECT 121.095 167.135 121.265 167.515 ;
        RECT 121.445 167.305 121.775 167.685 ;
        RECT 121.095 166.965 121.760 167.135 ;
        RECT 121.955 167.010 122.215 167.515 ;
        RECT 121.025 166.415 121.355 166.785 ;
        RECT 121.590 166.710 121.760 166.965 ;
        RECT 116.115 165.305 118.145 165.475 ;
        RECT 118.315 165.135 118.485 166.275 ;
        RECT 118.655 165.305 118.990 166.275 ;
        RECT 119.205 165.135 119.435 166.275 ;
        RECT 119.605 165.305 119.935 166.285 ;
        RECT 121.590 166.380 121.875 166.710 ;
        RECT 120.105 165.135 120.315 166.275 ;
        RECT 121.590 166.235 121.760 166.380 ;
        RECT 121.095 166.065 121.760 166.235 ;
        RECT 122.045 166.210 122.215 167.010 ;
        RECT 122.845 166.915 126.355 167.685 ;
        RECT 126.525 166.935 127.735 167.685 ;
        RECT 121.095 165.305 121.265 166.065 ;
        RECT 121.445 165.135 121.775 165.895 ;
        RECT 121.945 165.305 122.215 166.210 ;
        RECT 122.845 166.225 124.535 166.745 ;
        RECT 124.705 166.395 126.355 166.915 ;
        RECT 126.525 166.225 127.045 166.765 ;
        RECT 127.215 166.395 127.735 166.935 ;
        RECT 122.845 165.135 126.355 166.225 ;
        RECT 126.525 165.135 127.735 166.225 ;
        RECT 14.660 164.965 127.820 165.135 ;
        RECT 14.745 163.875 15.955 164.965 ;
        RECT 14.745 163.165 15.265 163.705 ;
        RECT 15.435 163.335 15.955 163.875 ;
        RECT 16.125 163.875 18.715 164.965 ;
        RECT 16.125 163.355 17.335 163.875 ;
        RECT 18.925 163.825 19.155 164.965 ;
        RECT 19.325 163.815 19.655 164.795 ;
        RECT 19.825 163.825 20.035 164.965 ;
        RECT 20.265 164.205 20.780 164.615 ;
        RECT 21.015 164.205 21.185 164.965 ;
        RECT 21.355 164.625 23.385 164.795 ;
        RECT 17.505 163.185 18.715 163.705 ;
        RECT 18.905 163.405 19.235 163.655 ;
        RECT 14.745 162.415 15.955 163.165 ;
        RECT 16.125 162.415 18.715 163.185 ;
        RECT 18.925 162.415 19.155 163.235 ;
        RECT 19.405 163.215 19.655 163.815 ;
        RECT 20.265 163.395 20.605 164.205 ;
        RECT 21.355 163.960 21.525 164.625 ;
        RECT 21.920 164.285 23.045 164.455 ;
        RECT 20.775 163.770 21.525 163.960 ;
        RECT 21.695 163.945 22.705 164.115 ;
        RECT 19.325 162.585 19.655 163.215 ;
        RECT 19.825 162.415 20.035 163.235 ;
        RECT 20.265 163.225 21.495 163.395 ;
        RECT 20.540 162.620 20.785 163.225 ;
        RECT 21.005 162.415 21.515 162.950 ;
        RECT 21.695 162.585 21.885 163.945 ;
        RECT 22.055 162.925 22.330 163.745 ;
        RECT 22.535 163.145 22.705 163.945 ;
        RECT 22.875 163.155 23.045 164.285 ;
        RECT 23.215 163.655 23.385 164.625 ;
        RECT 23.555 163.825 23.725 164.965 ;
        RECT 23.895 163.825 24.230 164.795 ;
        RECT 23.215 163.325 23.410 163.655 ;
        RECT 23.635 163.325 23.890 163.655 ;
        RECT 23.635 163.155 23.805 163.325 ;
        RECT 24.060 163.155 24.230 163.825 ;
        RECT 24.405 163.800 24.695 164.965 ;
        RECT 25.415 164.035 25.585 164.795 ;
        RECT 25.765 164.205 26.095 164.965 ;
        RECT 25.415 163.865 26.080 164.035 ;
        RECT 26.265 163.890 26.535 164.795 ;
        RECT 25.910 163.720 26.080 163.865 ;
        RECT 25.345 163.315 25.675 163.685 ;
        RECT 25.910 163.390 26.195 163.720 ;
        RECT 22.875 162.985 23.805 163.155 ;
        RECT 22.875 162.950 23.050 162.985 ;
        RECT 22.055 162.755 22.335 162.925 ;
        RECT 22.055 162.585 22.330 162.755 ;
        RECT 22.520 162.585 23.050 162.950 ;
        RECT 23.475 162.415 23.805 162.815 ;
        RECT 23.975 162.585 24.230 163.155 ;
        RECT 24.405 162.415 24.695 163.140 ;
        RECT 25.910 163.135 26.080 163.390 ;
        RECT 25.415 162.965 26.080 163.135 ;
        RECT 26.365 163.090 26.535 163.890 ;
        RECT 26.705 163.875 28.375 164.965 ;
        RECT 26.705 163.355 27.455 163.875 ;
        RECT 28.585 163.825 28.815 164.965 ;
        RECT 28.985 163.815 29.315 164.795 ;
        RECT 29.485 163.825 29.695 164.965 ;
        RECT 27.625 163.185 28.375 163.705 ;
        RECT 28.565 163.405 28.895 163.655 ;
        RECT 25.415 162.585 25.585 162.965 ;
        RECT 25.765 162.415 26.095 162.795 ;
        RECT 26.275 162.585 26.535 163.090 ;
        RECT 26.705 162.415 28.375 163.185 ;
        RECT 28.585 162.415 28.815 163.235 ;
        RECT 29.065 163.215 29.315 163.815 ;
        RECT 29.930 163.775 30.185 164.655 ;
        RECT 30.355 163.825 30.660 164.965 ;
        RECT 31.000 164.585 31.330 164.965 ;
        RECT 31.510 164.415 31.680 164.705 ;
        RECT 31.850 164.505 32.100 164.965 ;
        RECT 30.880 164.245 31.680 164.415 ;
        RECT 32.270 164.455 33.140 164.795 ;
        RECT 28.985 162.585 29.315 163.215 ;
        RECT 29.485 162.415 29.695 163.235 ;
        RECT 29.930 163.125 30.140 163.775 ;
        RECT 30.880 163.655 31.050 164.245 ;
        RECT 32.270 164.075 32.440 164.455 ;
        RECT 33.375 164.335 33.545 164.795 ;
        RECT 33.715 164.505 34.085 164.965 ;
        RECT 34.380 164.365 34.550 164.705 ;
        RECT 34.720 164.535 35.050 164.965 ;
        RECT 35.285 164.365 35.455 164.705 ;
        RECT 31.220 163.905 32.440 164.075 ;
        RECT 32.610 163.995 33.070 164.285 ;
        RECT 33.375 164.165 33.935 164.335 ;
        RECT 34.380 164.195 35.455 164.365 ;
        RECT 35.625 164.465 36.305 164.795 ;
        RECT 36.520 164.465 36.770 164.795 ;
        RECT 36.940 164.505 37.190 164.965 ;
        RECT 33.765 164.025 33.935 164.165 ;
        RECT 32.610 163.985 33.575 163.995 ;
        RECT 32.270 163.815 32.440 163.905 ;
        RECT 32.900 163.825 33.575 163.985 ;
        RECT 30.310 163.625 31.050 163.655 ;
        RECT 30.310 163.325 31.225 163.625 ;
        RECT 30.900 163.150 31.225 163.325 ;
        RECT 29.930 162.595 30.185 163.125 ;
        RECT 30.355 162.415 30.660 162.875 ;
        RECT 30.905 162.795 31.225 163.150 ;
        RECT 31.395 163.365 31.935 163.735 ;
        RECT 32.270 163.645 32.675 163.815 ;
        RECT 31.395 162.965 31.635 163.365 ;
        RECT 32.115 163.195 32.335 163.475 ;
        RECT 31.805 163.025 32.335 163.195 ;
        RECT 31.805 162.795 31.975 163.025 ;
        RECT 32.505 162.865 32.675 163.645 ;
        RECT 32.845 163.035 33.195 163.655 ;
        RECT 33.365 163.035 33.575 163.825 ;
        RECT 33.765 163.855 35.265 164.025 ;
        RECT 33.765 163.165 33.935 163.855 ;
        RECT 35.625 163.685 35.795 164.465 ;
        RECT 36.600 164.335 36.770 164.465 ;
        RECT 34.105 163.515 35.795 163.685 ;
        RECT 35.965 163.905 36.430 164.295 ;
        RECT 36.600 164.165 36.995 164.335 ;
        RECT 34.105 163.335 34.275 163.515 ;
        RECT 30.905 162.625 31.975 162.795 ;
        RECT 32.145 162.415 32.335 162.855 ;
        RECT 32.505 162.585 33.455 162.865 ;
        RECT 33.765 162.775 34.025 163.165 ;
        RECT 34.445 163.095 35.235 163.345 ;
        RECT 33.675 162.605 34.025 162.775 ;
        RECT 34.235 162.415 34.565 162.875 ;
        RECT 35.440 162.805 35.610 163.515 ;
        RECT 35.965 163.315 36.135 163.905 ;
        RECT 35.780 163.095 36.135 163.315 ;
        RECT 36.305 163.095 36.655 163.715 ;
        RECT 36.825 162.805 36.995 164.165 ;
        RECT 37.360 163.995 37.685 164.780 ;
        RECT 37.165 162.945 37.625 163.995 ;
        RECT 35.440 162.635 36.295 162.805 ;
        RECT 36.500 162.635 36.995 162.805 ;
        RECT 37.165 162.415 37.495 162.775 ;
        RECT 37.855 162.675 38.025 164.795 ;
        RECT 38.195 164.465 38.525 164.965 ;
        RECT 38.695 164.295 38.950 164.795 ;
        RECT 38.200 164.125 38.950 164.295 ;
        RECT 38.200 163.135 38.430 164.125 ;
        RECT 38.600 163.305 38.950 163.955 ;
        RECT 39.130 163.825 39.465 164.795 ;
        RECT 39.635 163.825 39.805 164.965 ;
        RECT 39.975 164.625 42.005 164.795 ;
        RECT 39.130 163.155 39.300 163.825 ;
        RECT 39.975 163.655 40.145 164.625 ;
        RECT 39.470 163.325 39.725 163.655 ;
        RECT 39.950 163.325 40.145 163.655 ;
        RECT 40.315 164.285 41.440 164.455 ;
        RECT 39.555 163.155 39.725 163.325 ;
        RECT 40.315 163.155 40.485 164.285 ;
        RECT 38.200 162.965 38.950 163.135 ;
        RECT 38.195 162.415 38.525 162.795 ;
        RECT 38.695 162.675 38.950 162.965 ;
        RECT 39.130 162.585 39.385 163.155 ;
        RECT 39.555 162.985 40.485 163.155 ;
        RECT 40.655 163.945 41.665 164.115 ;
        RECT 40.655 163.145 40.825 163.945 ;
        RECT 41.030 163.605 41.305 163.745 ;
        RECT 41.025 163.435 41.305 163.605 ;
        RECT 40.310 162.950 40.485 162.985 ;
        RECT 39.555 162.415 39.885 162.815 ;
        RECT 40.310 162.585 40.840 162.950 ;
        RECT 41.030 162.585 41.305 163.435 ;
        RECT 41.475 162.585 41.665 163.945 ;
        RECT 41.835 163.960 42.005 164.625 ;
        RECT 42.175 164.205 42.345 164.965 ;
        RECT 42.580 164.205 43.095 164.615 ;
        RECT 41.835 163.770 42.585 163.960 ;
        RECT 42.755 163.395 43.095 164.205 ;
        RECT 43.325 163.825 43.535 164.965 ;
        RECT 41.865 163.225 43.095 163.395 ;
        RECT 43.705 163.815 44.035 164.795 ;
        RECT 44.205 163.825 44.435 164.965 ;
        RECT 44.645 163.875 45.855 164.965 ;
        RECT 46.025 164.205 46.540 164.615 ;
        RECT 46.775 164.205 46.945 164.965 ;
        RECT 47.115 164.625 49.145 164.795 ;
        RECT 41.845 162.415 42.355 162.950 ;
        RECT 42.575 162.620 42.820 163.225 ;
        RECT 43.325 162.415 43.535 163.235 ;
        RECT 43.705 163.215 43.955 163.815 ;
        RECT 44.125 163.405 44.455 163.655 ;
        RECT 44.645 163.335 45.165 163.875 ;
        RECT 43.705 162.585 44.035 163.215 ;
        RECT 44.205 162.415 44.435 163.235 ;
        RECT 45.335 163.165 45.855 163.705 ;
        RECT 46.025 163.395 46.365 164.205 ;
        RECT 47.115 163.960 47.285 164.625 ;
        RECT 47.680 164.285 48.805 164.455 ;
        RECT 46.535 163.770 47.285 163.960 ;
        RECT 47.455 163.945 48.465 164.115 ;
        RECT 46.025 163.225 47.255 163.395 ;
        RECT 44.645 162.415 45.855 163.165 ;
        RECT 46.300 162.620 46.545 163.225 ;
        RECT 46.765 162.415 47.275 162.950 ;
        RECT 47.455 162.585 47.645 163.945 ;
        RECT 47.815 162.925 48.090 163.745 ;
        RECT 48.295 163.145 48.465 163.945 ;
        RECT 48.635 163.155 48.805 164.285 ;
        RECT 48.975 163.655 49.145 164.625 ;
        RECT 49.315 163.825 49.485 164.965 ;
        RECT 49.655 163.825 49.990 164.795 ;
        RECT 48.975 163.325 49.170 163.655 ;
        RECT 49.395 163.325 49.650 163.655 ;
        RECT 49.395 163.155 49.565 163.325 ;
        RECT 49.820 163.155 49.990 163.825 ;
        RECT 50.165 163.800 50.455 164.965 ;
        RECT 50.625 163.875 52.295 164.965 ;
        RECT 50.625 163.355 51.375 163.875 ;
        RECT 52.505 163.825 52.735 164.965 ;
        RECT 52.905 163.815 53.235 164.795 ;
        RECT 53.405 163.825 53.615 164.965 ;
        RECT 51.545 163.185 52.295 163.705 ;
        RECT 52.485 163.405 52.815 163.655 ;
        RECT 48.635 162.985 49.565 163.155 ;
        RECT 48.635 162.950 48.810 162.985 ;
        RECT 47.815 162.755 48.095 162.925 ;
        RECT 47.815 162.585 48.090 162.755 ;
        RECT 48.280 162.585 48.810 162.950 ;
        RECT 49.235 162.415 49.565 162.815 ;
        RECT 49.735 162.585 49.990 163.155 ;
        RECT 50.165 162.415 50.455 163.140 ;
        RECT 50.625 162.415 52.295 163.185 ;
        RECT 52.505 162.415 52.735 163.235 ;
        RECT 52.985 163.215 53.235 163.815 ;
        RECT 53.850 163.775 54.105 164.655 ;
        RECT 54.275 163.825 54.580 164.965 ;
        RECT 54.920 164.585 55.250 164.965 ;
        RECT 55.430 164.415 55.600 164.705 ;
        RECT 55.770 164.505 56.020 164.965 ;
        RECT 54.800 164.245 55.600 164.415 ;
        RECT 56.190 164.455 57.060 164.795 ;
        RECT 52.905 162.585 53.235 163.215 ;
        RECT 53.405 162.415 53.615 163.235 ;
        RECT 53.850 163.125 54.060 163.775 ;
        RECT 54.800 163.655 54.970 164.245 ;
        RECT 56.190 164.075 56.360 164.455 ;
        RECT 57.295 164.335 57.465 164.795 ;
        RECT 57.635 164.505 58.005 164.965 ;
        RECT 58.300 164.365 58.470 164.705 ;
        RECT 58.640 164.535 58.970 164.965 ;
        RECT 59.205 164.365 59.375 164.705 ;
        RECT 55.140 163.905 56.360 164.075 ;
        RECT 56.530 163.995 56.990 164.285 ;
        RECT 57.295 164.165 57.855 164.335 ;
        RECT 58.300 164.195 59.375 164.365 ;
        RECT 59.545 164.465 60.225 164.795 ;
        RECT 60.440 164.465 60.690 164.795 ;
        RECT 60.860 164.505 61.110 164.965 ;
        RECT 57.685 164.025 57.855 164.165 ;
        RECT 56.530 163.985 57.495 163.995 ;
        RECT 56.190 163.815 56.360 163.905 ;
        RECT 56.820 163.825 57.495 163.985 ;
        RECT 54.230 163.625 54.970 163.655 ;
        RECT 54.230 163.325 55.145 163.625 ;
        RECT 54.820 163.150 55.145 163.325 ;
        RECT 53.850 162.595 54.105 163.125 ;
        RECT 54.275 162.415 54.580 162.875 ;
        RECT 54.825 162.795 55.145 163.150 ;
        RECT 55.315 163.365 55.855 163.735 ;
        RECT 56.190 163.645 56.595 163.815 ;
        RECT 55.315 162.965 55.555 163.365 ;
        RECT 56.035 163.195 56.255 163.475 ;
        RECT 55.725 163.025 56.255 163.195 ;
        RECT 55.725 162.795 55.895 163.025 ;
        RECT 56.425 162.865 56.595 163.645 ;
        RECT 56.765 163.035 57.115 163.655 ;
        RECT 57.285 163.035 57.495 163.825 ;
        RECT 57.685 163.855 59.185 164.025 ;
        RECT 57.685 163.165 57.855 163.855 ;
        RECT 59.545 163.685 59.715 164.465 ;
        RECT 60.520 164.335 60.690 164.465 ;
        RECT 58.025 163.515 59.715 163.685 ;
        RECT 59.885 163.905 60.350 164.295 ;
        RECT 60.520 164.165 60.915 164.335 ;
        RECT 58.025 163.335 58.195 163.515 ;
        RECT 54.825 162.625 55.895 162.795 ;
        RECT 56.065 162.415 56.255 162.855 ;
        RECT 56.425 162.585 57.375 162.865 ;
        RECT 57.685 162.775 57.945 163.165 ;
        RECT 58.365 163.095 59.155 163.345 ;
        RECT 57.595 162.605 57.945 162.775 ;
        RECT 58.155 162.415 58.485 162.875 ;
        RECT 59.360 162.805 59.530 163.515 ;
        RECT 59.885 163.315 60.055 163.905 ;
        RECT 59.700 163.095 60.055 163.315 ;
        RECT 60.225 163.095 60.575 163.715 ;
        RECT 60.745 162.805 60.915 164.165 ;
        RECT 61.280 163.995 61.605 164.780 ;
        RECT 61.085 162.945 61.545 163.995 ;
        RECT 59.360 162.635 60.215 162.805 ;
        RECT 60.420 162.635 60.915 162.805 ;
        RECT 61.085 162.415 61.415 162.775 ;
        RECT 61.775 162.675 61.945 164.795 ;
        RECT 62.115 164.465 62.445 164.965 ;
        RECT 62.615 164.295 62.870 164.795 ;
        RECT 62.120 164.125 62.870 164.295 ;
        RECT 62.120 163.135 62.350 164.125 ;
        RECT 62.520 163.305 62.870 163.955 ;
        RECT 63.045 163.875 64.255 164.965 ;
        RECT 63.045 163.335 63.565 163.875 ;
        RECT 64.575 163.815 64.905 164.965 ;
        RECT 65.075 163.945 65.245 164.795 ;
        RECT 65.415 164.165 65.745 164.965 ;
        RECT 65.915 163.945 66.085 164.795 ;
        RECT 66.265 164.165 66.505 164.965 ;
        RECT 66.675 163.985 67.005 164.795 ;
        RECT 65.075 163.775 66.085 163.945 ;
        RECT 66.290 163.815 67.005 163.985 ;
        RECT 67.335 163.815 67.665 164.965 ;
        RECT 67.835 163.945 68.005 164.795 ;
        RECT 68.175 164.165 68.505 164.965 ;
        RECT 68.675 163.945 68.845 164.795 ;
        RECT 69.025 164.165 69.265 164.965 ;
        RECT 69.435 163.985 69.765 164.795 ;
        RECT 63.735 163.165 64.255 163.705 ;
        RECT 65.075 163.235 65.570 163.775 ;
        RECT 66.290 163.575 66.460 163.815 ;
        RECT 67.835 163.775 68.845 163.945 ;
        RECT 69.050 163.815 69.765 163.985 ;
        RECT 70.415 163.905 70.745 164.965 ;
        RECT 65.960 163.405 66.460 163.575 ;
        RECT 66.630 163.405 67.010 163.645 ;
        RECT 66.290 163.235 66.460 163.405 ;
        RECT 67.835 163.235 68.330 163.775 ;
        RECT 69.050 163.575 69.220 163.815 ;
        RECT 70.925 163.655 71.095 164.625 ;
        RECT 71.265 164.375 71.595 164.775 ;
        RECT 71.765 164.605 72.095 164.965 ;
        RECT 72.295 164.375 72.995 164.795 ;
        RECT 71.265 164.145 72.995 164.375 ;
        RECT 71.265 163.925 71.595 164.145 ;
        RECT 71.790 163.655 72.115 163.945 ;
        RECT 68.720 163.405 69.220 163.575 ;
        RECT 69.390 163.405 69.770 163.645 ;
        RECT 69.050 163.235 69.220 163.405 ;
        RECT 70.405 163.325 70.715 163.655 ;
        RECT 70.925 163.325 71.300 163.655 ;
        RECT 71.620 163.325 72.115 163.655 ;
        RECT 72.290 163.405 72.620 163.945 ;
        RECT 62.120 162.965 62.870 163.135 ;
        RECT 62.115 162.415 62.445 162.795 ;
        RECT 62.615 162.675 62.870 162.965 ;
        RECT 63.045 162.415 64.255 163.165 ;
        RECT 64.575 162.415 64.905 163.215 ;
        RECT 65.075 163.065 66.085 163.235 ;
        RECT 66.290 163.065 66.925 163.235 ;
        RECT 65.075 162.585 65.245 163.065 ;
        RECT 65.415 162.415 65.745 162.895 ;
        RECT 65.915 162.585 66.085 163.065 ;
        RECT 66.335 162.415 66.575 162.895 ;
        RECT 66.755 162.585 66.925 163.065 ;
        RECT 67.335 162.415 67.665 163.215 ;
        RECT 67.835 163.065 68.845 163.235 ;
        RECT 69.050 163.065 69.685 163.235 ;
        RECT 72.790 163.175 72.995 164.145 ;
        RECT 67.835 162.585 68.005 163.065 ;
        RECT 68.175 162.415 68.505 162.895 ;
        RECT 68.675 162.585 68.845 163.065 ;
        RECT 69.095 162.415 69.335 162.895 ;
        RECT 69.515 162.585 69.685 163.065 ;
        RECT 70.415 162.945 71.775 163.155 ;
        RECT 70.415 162.585 70.745 162.945 ;
        RECT 70.915 162.415 71.245 162.775 ;
        RECT 71.445 162.585 71.775 162.945 ;
        RECT 72.285 162.585 72.995 163.175 ;
        RECT 73.165 163.995 73.475 164.795 ;
        RECT 73.645 164.165 73.955 164.965 ;
        RECT 74.125 164.335 74.385 164.795 ;
        RECT 74.555 164.505 74.810 164.965 ;
        RECT 74.985 164.335 75.245 164.795 ;
        RECT 74.125 164.165 75.245 164.335 ;
        RECT 73.165 163.825 74.195 163.995 ;
        RECT 73.165 162.915 73.335 163.825 ;
        RECT 73.505 163.085 73.855 163.655 ;
        RECT 74.025 163.575 74.195 163.825 ;
        RECT 74.985 163.915 75.245 164.165 ;
        RECT 75.415 164.095 75.700 164.965 ;
        RECT 74.985 163.745 75.740 163.915 ;
        RECT 75.925 163.800 76.215 164.965 ;
        RECT 77.220 163.985 77.475 164.655 ;
        RECT 77.655 164.165 77.940 164.965 ;
        RECT 78.120 164.245 78.450 164.755 ;
        RECT 74.025 163.405 75.165 163.575 ;
        RECT 75.335 163.235 75.740 163.745 ;
        RECT 74.090 163.065 75.740 163.235 ;
        RECT 73.165 162.585 73.465 162.915 ;
        RECT 73.635 162.415 73.910 162.895 ;
        RECT 74.090 162.675 74.385 163.065 ;
        RECT 74.555 162.415 74.810 162.895 ;
        RECT 74.985 162.675 75.245 163.065 ;
        RECT 75.415 162.415 75.695 162.895 ;
        RECT 75.925 162.415 76.215 163.140 ;
        RECT 77.220 163.125 77.400 163.985 ;
        RECT 78.120 163.655 78.370 164.245 ;
        RECT 78.720 164.095 78.890 164.705 ;
        RECT 79.060 164.275 79.390 164.965 ;
        RECT 79.620 164.415 79.860 164.705 ;
        RECT 80.060 164.585 80.480 164.965 ;
        RECT 80.660 164.495 81.290 164.745 ;
        RECT 81.760 164.585 82.090 164.965 ;
        RECT 80.660 164.415 80.830 164.495 ;
        RECT 82.260 164.415 82.430 164.705 ;
        RECT 82.610 164.585 82.990 164.965 ;
        RECT 83.230 164.580 84.060 164.750 ;
        RECT 79.620 164.245 80.830 164.415 ;
        RECT 77.570 163.325 78.370 163.655 ;
        RECT 77.220 162.925 77.475 163.125 ;
        RECT 77.135 162.755 77.475 162.925 ;
        RECT 77.220 162.595 77.475 162.755 ;
        RECT 77.655 162.415 77.940 162.875 ;
        RECT 78.120 162.675 78.370 163.325 ;
        RECT 78.570 164.075 78.890 164.095 ;
        RECT 78.570 163.905 80.490 164.075 ;
        RECT 78.570 163.010 78.760 163.905 ;
        RECT 80.660 163.735 80.830 164.245 ;
        RECT 81.000 163.985 81.520 164.295 ;
        RECT 78.930 163.565 80.830 163.735 ;
        RECT 78.930 163.505 79.260 163.565 ;
        RECT 79.410 163.335 79.740 163.395 ;
        RECT 79.080 163.065 79.740 163.335 ;
        RECT 78.570 162.680 78.890 163.010 ;
        RECT 79.070 162.415 79.730 162.895 ;
        RECT 79.930 162.805 80.100 163.565 ;
        RECT 81.000 163.395 81.180 163.805 ;
        RECT 80.270 163.225 80.600 163.345 ;
        RECT 81.350 163.225 81.520 163.985 ;
        RECT 80.270 163.055 81.520 163.225 ;
        RECT 81.690 164.165 83.060 164.415 ;
        RECT 81.690 163.395 81.880 164.165 ;
        RECT 82.810 163.905 83.060 164.165 ;
        RECT 82.050 163.735 82.300 163.895 ;
        RECT 83.230 163.735 83.400 164.580 ;
        RECT 84.295 164.295 84.465 164.795 ;
        RECT 84.635 164.465 84.965 164.965 ;
        RECT 83.570 163.905 84.070 164.285 ;
        RECT 84.295 164.125 84.990 164.295 ;
        RECT 82.050 163.565 83.400 163.735 ;
        RECT 82.980 163.525 83.400 163.565 ;
        RECT 81.690 163.055 82.110 163.395 ;
        RECT 82.400 163.065 82.810 163.395 ;
        RECT 79.930 162.635 80.780 162.805 ;
        RECT 81.340 162.415 81.660 162.875 ;
        RECT 81.860 162.625 82.110 163.055 ;
        RECT 82.400 162.415 82.810 162.855 ;
        RECT 82.980 162.795 83.150 163.525 ;
        RECT 83.320 162.975 83.670 163.345 ;
        RECT 83.850 163.035 84.070 163.905 ;
        RECT 84.240 163.335 84.650 163.955 ;
        RECT 84.820 163.155 84.990 164.125 ;
        RECT 84.295 162.965 84.990 163.155 ;
        RECT 82.980 162.595 83.995 162.795 ;
        RECT 84.295 162.635 84.465 162.965 ;
        RECT 84.635 162.415 84.965 162.795 ;
        RECT 85.180 162.675 85.405 164.795 ;
        RECT 85.575 164.465 85.905 164.965 ;
        RECT 86.075 164.295 86.245 164.795 ;
        RECT 85.580 164.125 86.245 164.295 ;
        RECT 85.580 163.135 85.810 164.125 ;
        RECT 85.980 163.305 86.330 163.955 ;
        RECT 86.505 163.890 86.775 164.795 ;
        RECT 86.945 164.205 87.275 164.965 ;
        RECT 87.455 164.035 87.625 164.795 ;
        RECT 85.580 162.965 86.245 163.135 ;
        RECT 85.575 162.415 85.905 162.795 ;
        RECT 86.075 162.675 86.245 162.965 ;
        RECT 86.505 163.090 86.675 163.890 ;
        RECT 86.960 163.865 87.625 164.035 ;
        RECT 86.960 163.720 87.130 163.865 ;
        RECT 87.945 163.825 88.155 164.965 ;
        RECT 86.845 163.390 87.130 163.720 ;
        RECT 88.325 163.815 88.655 164.795 ;
        RECT 88.825 163.825 89.055 164.965 ;
        RECT 89.730 164.530 95.075 164.965 ;
        RECT 86.960 163.135 87.130 163.390 ;
        RECT 87.365 163.315 87.695 163.685 ;
        RECT 86.505 162.585 86.765 163.090 ;
        RECT 86.960 162.965 87.625 163.135 ;
        RECT 86.945 162.415 87.275 162.795 ;
        RECT 87.455 162.585 87.625 162.965 ;
        RECT 87.945 162.415 88.155 163.235 ;
        RECT 88.325 163.215 88.575 163.815 ;
        RECT 88.745 163.405 89.075 163.655 ;
        RECT 91.320 163.280 91.670 164.530 ;
        RECT 95.245 164.205 95.760 164.615 ;
        RECT 95.995 164.205 96.165 164.965 ;
        RECT 96.335 164.625 98.365 164.795 ;
        RECT 88.325 162.585 88.655 163.215 ;
        RECT 88.825 162.415 89.055 163.235 ;
        RECT 93.150 162.960 93.490 163.790 ;
        RECT 95.245 163.395 95.585 164.205 ;
        RECT 96.335 163.960 96.505 164.625 ;
        RECT 96.900 164.285 98.025 164.455 ;
        RECT 95.755 163.770 96.505 163.960 ;
        RECT 96.675 163.945 97.685 164.115 ;
        RECT 95.245 163.225 96.475 163.395 ;
        RECT 89.730 162.415 95.075 162.960 ;
        RECT 95.520 162.620 95.765 163.225 ;
        RECT 95.985 162.415 96.495 162.950 ;
        RECT 96.675 162.585 96.865 163.945 ;
        RECT 97.035 163.605 97.310 163.745 ;
        RECT 97.035 163.435 97.315 163.605 ;
        RECT 97.035 162.585 97.310 163.435 ;
        RECT 97.515 163.145 97.685 163.945 ;
        RECT 97.855 163.155 98.025 164.285 ;
        RECT 98.195 163.655 98.365 164.625 ;
        RECT 98.535 163.825 98.705 164.965 ;
        RECT 98.875 163.825 99.210 164.795 ;
        RECT 100.345 163.825 100.575 164.965 ;
        RECT 98.195 163.325 98.390 163.655 ;
        RECT 98.615 163.325 98.870 163.655 ;
        RECT 98.615 163.155 98.785 163.325 ;
        RECT 99.040 163.155 99.210 163.825 ;
        RECT 100.745 163.815 101.075 164.795 ;
        RECT 101.245 163.825 101.455 164.965 ;
        RECT 100.325 163.405 100.655 163.655 ;
        RECT 97.855 162.985 98.785 163.155 ;
        RECT 97.855 162.950 98.030 162.985 ;
        RECT 97.500 162.585 98.030 162.950 ;
        RECT 98.455 162.415 98.785 162.815 ;
        RECT 98.955 162.585 99.210 163.155 ;
        RECT 100.345 162.415 100.575 163.235 ;
        RECT 100.825 163.215 101.075 163.815 ;
        RECT 101.685 163.800 101.975 164.965 ;
        RECT 102.520 163.985 102.775 164.655 ;
        RECT 102.955 164.165 103.240 164.965 ;
        RECT 103.420 164.245 103.750 164.755 ;
        RECT 102.520 163.945 102.700 163.985 ;
        RECT 102.435 163.775 102.700 163.945 ;
        RECT 100.745 162.585 101.075 163.215 ;
        RECT 101.245 162.415 101.455 163.235 ;
        RECT 101.685 162.415 101.975 163.140 ;
        RECT 102.520 163.125 102.700 163.775 ;
        RECT 103.420 163.655 103.670 164.245 ;
        RECT 104.020 164.095 104.190 164.705 ;
        RECT 104.360 164.275 104.690 164.965 ;
        RECT 104.920 164.415 105.160 164.705 ;
        RECT 105.360 164.585 105.780 164.965 ;
        RECT 105.960 164.495 106.590 164.745 ;
        RECT 107.060 164.585 107.390 164.965 ;
        RECT 105.960 164.415 106.130 164.495 ;
        RECT 107.560 164.415 107.730 164.705 ;
        RECT 107.910 164.585 108.290 164.965 ;
        RECT 108.530 164.580 109.360 164.750 ;
        RECT 104.920 164.245 106.130 164.415 ;
        RECT 102.870 163.325 103.670 163.655 ;
        RECT 102.520 162.595 102.775 163.125 ;
        RECT 102.955 162.415 103.240 162.875 ;
        RECT 103.420 162.675 103.670 163.325 ;
        RECT 103.870 164.075 104.190 164.095 ;
        RECT 103.870 163.905 105.790 164.075 ;
        RECT 103.870 163.010 104.060 163.905 ;
        RECT 105.960 163.735 106.130 164.245 ;
        RECT 106.300 163.985 106.820 164.295 ;
        RECT 104.230 163.565 106.130 163.735 ;
        RECT 104.230 163.505 104.560 163.565 ;
        RECT 104.710 163.335 105.040 163.395 ;
        RECT 104.380 163.065 105.040 163.335 ;
        RECT 103.870 162.680 104.190 163.010 ;
        RECT 104.370 162.415 105.030 162.895 ;
        RECT 105.230 162.805 105.400 163.565 ;
        RECT 106.300 163.395 106.480 163.805 ;
        RECT 105.570 163.225 105.900 163.345 ;
        RECT 106.650 163.225 106.820 163.985 ;
        RECT 105.570 163.055 106.820 163.225 ;
        RECT 106.990 164.165 108.360 164.415 ;
        RECT 106.990 163.395 107.180 164.165 ;
        RECT 108.110 163.905 108.360 164.165 ;
        RECT 107.350 163.735 107.600 163.895 ;
        RECT 108.530 163.735 108.700 164.580 ;
        RECT 109.595 164.295 109.765 164.795 ;
        RECT 109.935 164.465 110.265 164.965 ;
        RECT 108.870 163.905 109.370 164.285 ;
        RECT 109.595 164.125 110.290 164.295 ;
        RECT 107.350 163.565 108.700 163.735 ;
        RECT 108.280 163.525 108.700 163.565 ;
        RECT 106.990 163.055 107.410 163.395 ;
        RECT 107.700 163.065 108.110 163.395 ;
        RECT 105.230 162.635 106.080 162.805 ;
        RECT 106.640 162.415 106.960 162.875 ;
        RECT 107.160 162.625 107.410 163.055 ;
        RECT 107.700 162.415 108.110 162.855 ;
        RECT 108.280 162.795 108.450 163.525 ;
        RECT 108.620 162.975 108.970 163.345 ;
        RECT 109.150 163.035 109.370 163.905 ;
        RECT 109.540 163.335 109.950 163.955 ;
        RECT 110.120 163.155 110.290 164.125 ;
        RECT 109.595 162.965 110.290 163.155 ;
        RECT 108.280 162.595 109.295 162.795 ;
        RECT 109.595 162.635 109.765 162.965 ;
        RECT 109.935 162.415 110.265 162.795 ;
        RECT 110.480 162.675 110.705 164.795 ;
        RECT 110.875 164.465 111.205 164.965 ;
        RECT 111.375 164.295 111.545 164.795 ;
        RECT 110.880 164.125 111.545 164.295 ;
        RECT 112.265 164.205 112.780 164.615 ;
        RECT 113.015 164.205 113.185 164.965 ;
        RECT 113.355 164.625 115.385 164.795 ;
        RECT 110.880 163.135 111.110 164.125 ;
        RECT 111.280 163.305 111.630 163.955 ;
        RECT 112.265 163.395 112.605 164.205 ;
        RECT 113.355 163.960 113.525 164.625 ;
        RECT 113.920 164.285 115.045 164.455 ;
        RECT 112.775 163.770 113.525 163.960 ;
        RECT 113.695 163.945 114.705 164.115 ;
        RECT 112.265 163.225 113.495 163.395 ;
        RECT 110.880 162.965 111.545 163.135 ;
        RECT 110.875 162.415 111.205 162.795 ;
        RECT 111.375 162.675 111.545 162.965 ;
        RECT 112.540 162.620 112.785 163.225 ;
        RECT 113.005 162.415 113.515 162.950 ;
        RECT 113.695 162.585 113.885 163.945 ;
        RECT 114.055 162.925 114.330 163.745 ;
        RECT 114.535 163.145 114.705 163.945 ;
        RECT 114.875 163.155 115.045 164.285 ;
        RECT 115.215 163.655 115.385 164.625 ;
        RECT 115.555 163.825 115.725 164.965 ;
        RECT 115.895 163.825 116.230 164.795 ;
        RECT 115.215 163.325 115.410 163.655 ;
        RECT 115.635 163.325 115.890 163.655 ;
        RECT 115.635 163.155 115.805 163.325 ;
        RECT 116.060 163.155 116.230 163.825 ;
        RECT 114.875 162.985 115.805 163.155 ;
        RECT 114.875 162.950 115.050 162.985 ;
        RECT 114.055 162.755 114.335 162.925 ;
        RECT 114.055 162.585 114.330 162.755 ;
        RECT 114.520 162.585 115.050 162.950 ;
        RECT 115.475 162.415 115.805 162.815 ;
        RECT 115.975 162.585 116.230 163.155 ;
        RECT 116.410 163.775 116.665 164.655 ;
        RECT 116.835 163.825 117.140 164.965 ;
        RECT 117.480 164.585 117.810 164.965 ;
        RECT 117.990 164.415 118.160 164.705 ;
        RECT 118.330 164.505 118.580 164.965 ;
        RECT 117.360 164.245 118.160 164.415 ;
        RECT 118.750 164.455 119.620 164.795 ;
        RECT 116.410 163.125 116.620 163.775 ;
        RECT 117.360 163.655 117.530 164.245 ;
        RECT 118.750 164.075 118.920 164.455 ;
        RECT 119.855 164.335 120.025 164.795 ;
        RECT 120.195 164.505 120.565 164.965 ;
        RECT 120.860 164.365 121.030 164.705 ;
        RECT 121.200 164.535 121.530 164.965 ;
        RECT 121.765 164.365 121.935 164.705 ;
        RECT 117.700 163.905 118.920 164.075 ;
        RECT 119.090 163.995 119.550 164.285 ;
        RECT 119.855 164.165 120.415 164.335 ;
        RECT 120.860 164.195 121.935 164.365 ;
        RECT 122.105 164.465 122.785 164.795 ;
        RECT 123.000 164.465 123.250 164.795 ;
        RECT 123.420 164.505 123.670 164.965 ;
        RECT 120.245 164.025 120.415 164.165 ;
        RECT 119.090 163.985 120.055 163.995 ;
        RECT 118.750 163.815 118.920 163.905 ;
        RECT 119.380 163.825 120.055 163.985 ;
        RECT 116.790 163.625 117.530 163.655 ;
        RECT 116.790 163.325 117.705 163.625 ;
        RECT 117.380 163.150 117.705 163.325 ;
        RECT 116.410 162.595 116.665 163.125 ;
        RECT 116.835 162.415 117.140 162.875 ;
        RECT 117.385 162.795 117.705 163.150 ;
        RECT 117.875 163.365 118.415 163.735 ;
        RECT 118.750 163.645 119.155 163.815 ;
        RECT 117.875 162.965 118.115 163.365 ;
        RECT 118.595 163.195 118.815 163.475 ;
        RECT 118.285 163.025 118.815 163.195 ;
        RECT 118.285 162.795 118.455 163.025 ;
        RECT 118.985 162.865 119.155 163.645 ;
        RECT 119.325 163.035 119.675 163.655 ;
        RECT 119.845 163.035 120.055 163.825 ;
        RECT 120.245 163.855 121.745 164.025 ;
        RECT 120.245 163.165 120.415 163.855 ;
        RECT 122.105 163.685 122.275 164.465 ;
        RECT 123.080 164.335 123.250 164.465 ;
        RECT 120.585 163.515 122.275 163.685 ;
        RECT 122.445 163.905 122.910 164.295 ;
        RECT 123.080 164.165 123.475 164.335 ;
        RECT 120.585 163.335 120.755 163.515 ;
        RECT 117.385 162.625 118.455 162.795 ;
        RECT 118.625 162.415 118.815 162.855 ;
        RECT 118.985 162.585 119.935 162.865 ;
        RECT 120.245 162.775 120.505 163.165 ;
        RECT 120.925 163.095 121.715 163.345 ;
        RECT 120.155 162.605 120.505 162.775 ;
        RECT 120.715 162.415 121.045 162.875 ;
        RECT 121.920 162.805 122.090 163.515 ;
        RECT 122.445 163.315 122.615 163.905 ;
        RECT 122.260 163.095 122.615 163.315 ;
        RECT 122.785 163.095 123.135 163.715 ;
        RECT 123.305 162.805 123.475 164.165 ;
        RECT 123.840 163.995 124.165 164.780 ;
        RECT 123.645 162.945 124.105 163.995 ;
        RECT 121.920 162.635 122.775 162.805 ;
        RECT 122.980 162.635 123.475 162.805 ;
        RECT 123.645 162.415 123.975 162.775 ;
        RECT 124.335 162.675 124.505 164.795 ;
        RECT 124.675 164.465 125.005 164.965 ;
        RECT 125.175 164.295 125.430 164.795 ;
        RECT 124.680 164.125 125.430 164.295 ;
        RECT 124.680 163.135 124.910 164.125 ;
        RECT 125.080 163.305 125.430 163.955 ;
        RECT 126.525 163.875 127.735 164.965 ;
        RECT 126.525 163.335 127.045 163.875 ;
        RECT 127.215 163.165 127.735 163.705 ;
        RECT 124.680 162.965 125.430 163.135 ;
        RECT 124.675 162.415 125.005 162.795 ;
        RECT 125.175 162.675 125.430 162.965 ;
        RECT 126.525 162.415 127.735 163.165 ;
        RECT 14.660 162.245 127.820 162.415 ;
        RECT 14.745 161.495 15.955 162.245 ;
        RECT 14.745 160.955 15.265 161.495 ;
        RECT 16.645 161.425 16.855 162.245 ;
        RECT 17.025 161.445 17.355 162.075 ;
        RECT 15.435 160.785 15.955 161.325 ;
        RECT 17.025 160.845 17.275 161.445 ;
        RECT 17.525 161.425 17.755 162.245 ;
        RECT 18.340 161.905 18.595 162.065 ;
        RECT 18.255 161.735 18.595 161.905 ;
        RECT 18.775 161.785 19.060 162.245 ;
        RECT 18.340 161.535 18.595 161.735 ;
        RECT 17.445 161.005 17.775 161.255 ;
        RECT 14.745 159.695 15.955 160.785 ;
        RECT 16.645 159.695 16.855 160.835 ;
        RECT 17.025 159.865 17.355 160.845 ;
        RECT 17.525 159.695 17.755 160.835 ;
        RECT 18.340 160.675 18.520 161.535 ;
        RECT 19.240 161.335 19.490 161.985 ;
        RECT 18.690 161.005 19.490 161.335 ;
        RECT 18.340 160.005 18.595 160.675 ;
        RECT 18.775 159.695 19.060 160.495 ;
        RECT 19.240 160.415 19.490 161.005 ;
        RECT 19.690 161.650 20.010 161.980 ;
        RECT 20.190 161.765 20.850 162.245 ;
        RECT 21.050 161.855 21.900 162.025 ;
        RECT 19.690 160.755 19.880 161.650 ;
        RECT 20.200 161.325 20.860 161.595 ;
        RECT 20.530 161.265 20.860 161.325 ;
        RECT 20.050 161.095 20.380 161.155 ;
        RECT 21.050 161.095 21.220 161.855 ;
        RECT 22.460 161.785 22.780 162.245 ;
        RECT 22.980 161.605 23.230 162.035 ;
        RECT 23.520 161.805 23.930 162.245 ;
        RECT 24.100 161.865 25.115 162.065 ;
        RECT 21.390 161.435 22.640 161.605 ;
        RECT 21.390 161.315 21.720 161.435 ;
        RECT 20.050 160.925 21.950 161.095 ;
        RECT 19.690 160.585 21.610 160.755 ;
        RECT 19.690 160.565 20.010 160.585 ;
        RECT 19.240 159.905 19.570 160.415 ;
        RECT 19.840 159.955 20.010 160.565 ;
        RECT 21.780 160.415 21.950 160.925 ;
        RECT 22.120 160.855 22.300 161.265 ;
        RECT 22.470 160.675 22.640 161.435 ;
        RECT 20.180 159.695 20.510 160.385 ;
        RECT 20.740 160.245 21.950 160.415 ;
        RECT 22.120 160.365 22.640 160.675 ;
        RECT 22.810 161.265 23.230 161.605 ;
        RECT 23.520 161.265 23.930 161.595 ;
        RECT 22.810 160.495 23.000 161.265 ;
        RECT 24.100 161.135 24.270 161.865 ;
        RECT 25.415 161.695 25.585 162.025 ;
        RECT 25.755 161.865 26.085 162.245 ;
        RECT 24.440 161.315 24.790 161.685 ;
        RECT 24.100 161.095 24.520 161.135 ;
        RECT 23.170 160.925 24.520 161.095 ;
        RECT 23.170 160.765 23.420 160.925 ;
        RECT 23.930 160.495 24.180 160.755 ;
        RECT 22.810 160.245 24.180 160.495 ;
        RECT 20.740 159.955 20.980 160.245 ;
        RECT 21.780 160.165 21.950 160.245 ;
        RECT 21.180 159.695 21.600 160.075 ;
        RECT 21.780 159.915 22.410 160.165 ;
        RECT 22.880 159.695 23.210 160.075 ;
        RECT 23.380 159.955 23.550 160.245 ;
        RECT 24.350 160.080 24.520 160.925 ;
        RECT 24.970 160.755 25.190 161.625 ;
        RECT 25.415 161.505 26.110 161.695 ;
        RECT 24.690 160.375 25.190 160.755 ;
        RECT 25.360 160.705 25.770 161.325 ;
        RECT 25.940 160.535 26.110 161.505 ;
        RECT 25.415 160.365 26.110 160.535 ;
        RECT 23.730 159.695 24.110 160.075 ;
        RECT 24.350 159.910 25.180 160.080 ;
        RECT 25.415 159.865 25.585 160.365 ;
        RECT 25.755 159.695 26.085 160.195 ;
        RECT 26.300 159.865 26.525 161.985 ;
        RECT 26.695 161.865 27.025 162.245 ;
        RECT 27.195 161.695 27.365 161.985 ;
        RECT 26.700 161.525 27.365 161.695 ;
        RECT 27.715 161.695 27.885 161.985 ;
        RECT 28.055 161.865 28.385 162.245 ;
        RECT 27.715 161.525 28.380 161.695 ;
        RECT 26.700 160.535 26.930 161.525 ;
        RECT 27.100 160.705 27.450 161.355 ;
        RECT 27.630 160.705 27.980 161.355 ;
        RECT 28.150 160.535 28.380 161.525 ;
        RECT 26.700 160.365 27.365 160.535 ;
        RECT 26.695 159.695 27.025 160.195 ;
        RECT 27.195 159.865 27.365 160.365 ;
        RECT 27.715 160.365 28.380 160.535 ;
        RECT 27.715 159.865 27.885 160.365 ;
        RECT 28.055 159.695 28.385 160.195 ;
        RECT 28.555 159.865 28.780 161.985 ;
        RECT 28.995 161.865 29.325 162.245 ;
        RECT 29.495 161.695 29.665 162.025 ;
        RECT 29.965 161.865 30.980 162.065 ;
        RECT 28.970 161.505 29.665 161.695 ;
        RECT 28.970 160.535 29.140 161.505 ;
        RECT 29.310 160.705 29.720 161.325 ;
        RECT 29.890 160.755 30.110 161.625 ;
        RECT 30.290 161.315 30.640 161.685 ;
        RECT 30.810 161.135 30.980 161.865 ;
        RECT 31.150 161.805 31.560 162.245 ;
        RECT 31.850 161.605 32.100 162.035 ;
        RECT 32.300 161.785 32.620 162.245 ;
        RECT 33.180 161.855 34.030 162.025 ;
        RECT 31.150 161.265 31.560 161.595 ;
        RECT 31.850 161.265 32.270 161.605 ;
        RECT 30.560 161.095 30.980 161.135 ;
        RECT 30.560 160.925 31.910 161.095 ;
        RECT 28.970 160.365 29.665 160.535 ;
        RECT 29.890 160.375 30.390 160.755 ;
        RECT 28.995 159.695 29.325 160.195 ;
        RECT 29.495 159.865 29.665 160.365 ;
        RECT 30.560 160.080 30.730 160.925 ;
        RECT 31.660 160.765 31.910 160.925 ;
        RECT 30.900 160.495 31.150 160.755 ;
        RECT 32.080 160.495 32.270 161.265 ;
        RECT 30.900 160.245 32.270 160.495 ;
        RECT 32.440 161.435 33.690 161.605 ;
        RECT 32.440 160.675 32.610 161.435 ;
        RECT 33.360 161.315 33.690 161.435 ;
        RECT 32.780 160.855 32.960 161.265 ;
        RECT 33.860 161.095 34.030 161.855 ;
        RECT 34.230 161.765 34.890 162.245 ;
        RECT 35.070 161.650 35.390 161.980 ;
        RECT 34.220 161.325 34.880 161.595 ;
        RECT 34.220 161.265 34.550 161.325 ;
        RECT 34.700 161.095 35.030 161.155 ;
        RECT 33.130 160.925 35.030 161.095 ;
        RECT 32.440 160.365 32.960 160.675 ;
        RECT 33.130 160.415 33.300 160.925 ;
        RECT 35.200 160.755 35.390 161.650 ;
        RECT 33.470 160.585 35.390 160.755 ;
        RECT 35.070 160.565 35.390 160.585 ;
        RECT 35.590 161.335 35.840 161.985 ;
        RECT 36.020 161.785 36.305 162.245 ;
        RECT 36.485 161.535 36.740 162.065 ;
        RECT 35.590 161.005 36.390 161.335 ;
        RECT 33.130 160.245 34.340 160.415 ;
        RECT 29.900 159.910 30.730 160.080 ;
        RECT 30.970 159.695 31.350 160.075 ;
        RECT 31.530 159.955 31.700 160.245 ;
        RECT 33.130 160.165 33.300 160.245 ;
        RECT 31.870 159.695 32.200 160.075 ;
        RECT 32.670 159.915 33.300 160.165 ;
        RECT 33.480 159.695 33.900 160.075 ;
        RECT 34.100 159.955 34.340 160.245 ;
        RECT 34.570 159.695 34.900 160.385 ;
        RECT 35.070 159.955 35.240 160.565 ;
        RECT 35.590 160.415 35.840 161.005 ;
        RECT 36.560 160.675 36.740 161.535 ;
        RECT 37.285 161.520 37.575 162.245 ;
        RECT 37.745 161.570 38.005 162.075 ;
        RECT 38.185 161.865 38.515 162.245 ;
        RECT 38.695 161.695 38.865 162.075 ;
        RECT 35.510 159.905 35.840 160.415 ;
        RECT 36.020 159.695 36.305 160.495 ;
        RECT 36.485 160.205 36.740 160.675 ;
        RECT 36.485 160.035 36.825 160.205 ;
        RECT 36.485 160.005 36.740 160.035 ;
        RECT 37.285 159.695 37.575 160.860 ;
        RECT 37.745 160.770 37.915 161.570 ;
        RECT 38.200 161.525 38.865 161.695 ;
        RECT 39.125 161.570 39.385 162.075 ;
        RECT 39.565 161.865 39.895 162.245 ;
        RECT 40.075 161.695 40.245 162.075 ;
        RECT 38.200 161.270 38.370 161.525 ;
        RECT 38.085 160.940 38.370 161.270 ;
        RECT 38.605 160.975 38.935 161.345 ;
        RECT 38.200 160.795 38.370 160.940 ;
        RECT 37.745 159.865 38.015 160.770 ;
        RECT 38.200 160.625 38.865 160.795 ;
        RECT 38.185 159.695 38.515 160.455 ;
        RECT 38.695 159.865 38.865 160.625 ;
        RECT 39.125 160.770 39.295 161.570 ;
        RECT 39.580 161.525 40.245 161.695 ;
        RECT 40.510 161.535 40.765 162.065 ;
        RECT 40.935 161.785 41.240 162.245 ;
        RECT 41.485 161.865 42.555 162.035 ;
        RECT 39.580 161.270 39.750 161.525 ;
        RECT 39.465 160.940 39.750 161.270 ;
        RECT 39.985 160.975 40.315 161.345 ;
        RECT 39.580 160.795 39.750 160.940 ;
        RECT 40.510 160.885 40.720 161.535 ;
        RECT 41.485 161.510 41.805 161.865 ;
        RECT 41.480 161.335 41.805 161.510 ;
        RECT 40.890 161.035 41.805 161.335 ;
        RECT 41.975 161.295 42.215 161.695 ;
        RECT 42.385 161.635 42.555 161.865 ;
        RECT 42.725 161.805 42.915 162.245 ;
        RECT 43.085 161.795 44.035 162.075 ;
        RECT 44.255 161.885 44.605 162.055 ;
        RECT 42.385 161.465 42.915 161.635 ;
        RECT 40.890 161.005 41.630 161.035 ;
        RECT 39.125 159.865 39.395 160.770 ;
        RECT 39.580 160.625 40.245 160.795 ;
        RECT 39.565 159.695 39.895 160.455 ;
        RECT 40.075 159.865 40.245 160.625 ;
        RECT 40.510 160.005 40.765 160.885 ;
        RECT 40.935 159.695 41.240 160.835 ;
        RECT 41.460 160.415 41.630 161.005 ;
        RECT 41.975 160.925 42.515 161.295 ;
        RECT 42.695 161.185 42.915 161.465 ;
        RECT 43.085 161.015 43.255 161.795 ;
        RECT 42.850 160.845 43.255 161.015 ;
        RECT 43.425 161.005 43.775 161.625 ;
        RECT 42.850 160.755 43.020 160.845 ;
        RECT 43.945 160.835 44.155 161.625 ;
        RECT 41.800 160.585 43.020 160.755 ;
        RECT 43.480 160.675 44.155 160.835 ;
        RECT 41.460 160.245 42.260 160.415 ;
        RECT 41.580 159.695 41.910 160.075 ;
        RECT 42.090 159.955 42.260 160.245 ;
        RECT 42.850 160.205 43.020 160.585 ;
        RECT 43.190 160.665 44.155 160.675 ;
        RECT 44.345 161.495 44.605 161.885 ;
        RECT 44.815 161.785 45.145 162.245 ;
        RECT 46.020 161.855 46.875 162.025 ;
        RECT 47.080 161.855 47.575 162.025 ;
        RECT 47.745 161.885 48.075 162.245 ;
        RECT 44.345 160.805 44.515 161.495 ;
        RECT 44.685 161.145 44.855 161.325 ;
        RECT 45.025 161.315 45.815 161.565 ;
        RECT 46.020 161.145 46.190 161.855 ;
        RECT 46.360 161.345 46.715 161.565 ;
        RECT 44.685 160.975 46.375 161.145 ;
        RECT 43.190 160.375 43.650 160.665 ;
        RECT 44.345 160.635 45.845 160.805 ;
        RECT 44.345 160.495 44.515 160.635 ;
        RECT 43.955 160.325 44.515 160.495 ;
        RECT 42.430 159.695 42.680 160.155 ;
        RECT 42.850 159.865 43.720 160.205 ;
        RECT 43.955 159.865 44.125 160.325 ;
        RECT 44.960 160.295 46.035 160.465 ;
        RECT 44.295 159.695 44.665 160.155 ;
        RECT 44.960 159.955 45.130 160.295 ;
        RECT 45.300 159.695 45.630 160.125 ;
        RECT 45.865 159.955 46.035 160.295 ;
        RECT 46.205 160.195 46.375 160.975 ;
        RECT 46.545 160.755 46.715 161.345 ;
        RECT 46.885 160.945 47.235 161.565 ;
        RECT 46.545 160.365 47.010 160.755 ;
        RECT 47.405 160.495 47.575 161.855 ;
        RECT 47.745 160.665 48.205 161.715 ;
        RECT 47.180 160.325 47.575 160.495 ;
        RECT 47.180 160.195 47.350 160.325 ;
        RECT 46.205 159.865 46.885 160.195 ;
        RECT 47.100 159.865 47.350 160.195 ;
        RECT 47.520 159.695 47.770 160.155 ;
        RECT 47.940 159.880 48.265 160.665 ;
        RECT 48.435 159.865 48.605 161.985 ;
        RECT 48.775 161.865 49.105 162.245 ;
        RECT 49.275 161.695 49.530 161.985 ;
        RECT 48.780 161.525 49.530 161.695 ;
        RECT 49.705 161.570 49.965 162.075 ;
        RECT 50.145 161.865 50.475 162.245 ;
        RECT 50.655 161.695 50.825 162.075 ;
        RECT 48.780 160.535 49.010 161.525 ;
        RECT 49.180 160.705 49.530 161.355 ;
        RECT 49.705 160.770 49.875 161.570 ;
        RECT 50.160 161.525 50.825 161.695 ;
        RECT 50.160 161.270 50.330 161.525 ;
        RECT 52.045 161.425 52.275 162.245 ;
        RECT 52.445 161.445 52.775 162.075 ;
        RECT 50.045 160.940 50.330 161.270 ;
        RECT 50.565 160.975 50.895 161.345 ;
        RECT 52.025 161.005 52.355 161.255 ;
        RECT 50.160 160.795 50.330 160.940 ;
        RECT 52.525 160.845 52.775 161.445 ;
        RECT 52.945 161.425 53.155 162.245 ;
        RECT 53.660 161.435 53.905 162.040 ;
        RECT 54.125 161.710 54.635 162.245 ;
        RECT 48.780 160.365 49.530 160.535 ;
        RECT 48.775 159.695 49.105 160.195 ;
        RECT 49.275 159.865 49.530 160.365 ;
        RECT 49.705 159.865 49.975 160.770 ;
        RECT 50.160 160.625 50.825 160.795 ;
        RECT 50.145 159.695 50.475 160.455 ;
        RECT 50.655 159.865 50.825 160.625 ;
        RECT 52.045 159.695 52.275 160.835 ;
        RECT 52.445 159.865 52.775 160.845 ;
        RECT 53.385 161.265 54.615 161.435 ;
        RECT 52.945 159.695 53.155 160.835 ;
        RECT 53.385 160.455 53.725 161.265 ;
        RECT 53.895 160.700 54.645 160.890 ;
        RECT 53.385 160.045 53.900 160.455 ;
        RECT 54.135 159.695 54.305 160.455 ;
        RECT 54.475 160.035 54.645 160.700 ;
        RECT 54.815 160.715 55.005 162.075 ;
        RECT 55.175 161.225 55.450 162.075 ;
        RECT 55.640 161.710 56.170 162.075 ;
        RECT 56.595 161.845 56.925 162.245 ;
        RECT 55.995 161.675 56.170 161.710 ;
        RECT 55.175 161.055 55.455 161.225 ;
        RECT 55.175 160.915 55.450 161.055 ;
        RECT 55.655 160.715 55.825 161.515 ;
        RECT 54.815 160.545 55.825 160.715 ;
        RECT 55.995 161.505 56.925 161.675 ;
        RECT 57.095 161.505 57.350 162.075 ;
        RECT 55.995 160.375 56.165 161.505 ;
        RECT 56.755 161.335 56.925 161.505 ;
        RECT 55.040 160.205 56.165 160.375 ;
        RECT 56.335 161.005 56.530 161.335 ;
        RECT 56.755 161.005 57.010 161.335 ;
        RECT 56.335 160.035 56.505 161.005 ;
        RECT 57.180 160.835 57.350 161.505 ;
        RECT 57.525 161.495 58.735 162.245 ;
        RECT 58.995 161.695 59.165 162.075 ;
        RECT 59.345 161.865 59.675 162.245 ;
        RECT 58.995 161.525 59.660 161.695 ;
        RECT 59.855 161.570 60.115 162.075 ;
        RECT 54.475 159.865 56.505 160.035 ;
        RECT 56.675 159.695 56.845 160.835 ;
        RECT 57.015 159.865 57.350 160.835 ;
        RECT 57.525 160.785 58.045 161.325 ;
        RECT 58.215 160.955 58.735 161.495 ;
        RECT 58.925 160.975 59.255 161.345 ;
        RECT 59.490 161.270 59.660 161.525 ;
        RECT 59.490 160.940 59.775 161.270 ;
        RECT 59.490 160.795 59.660 160.940 ;
        RECT 57.525 159.695 58.735 160.785 ;
        RECT 58.995 160.625 59.660 160.795 ;
        RECT 59.945 160.770 60.115 161.570 ;
        RECT 60.435 161.445 60.765 162.245 ;
        RECT 60.935 161.595 61.105 162.075 ;
        RECT 61.275 161.765 61.605 162.245 ;
        RECT 61.775 161.595 61.945 162.075 ;
        RECT 62.195 161.765 62.435 162.245 ;
        RECT 62.615 161.595 62.785 162.075 ;
        RECT 60.935 161.425 61.945 161.595 ;
        RECT 62.150 161.425 62.785 161.595 ;
        RECT 63.045 161.520 63.335 162.245 ;
        RECT 63.965 161.475 65.635 162.245 ;
        RECT 65.865 161.765 66.145 162.245 ;
        RECT 66.315 161.595 66.575 161.985 ;
        RECT 66.750 161.765 67.005 162.245 ;
        RECT 67.175 161.595 67.470 161.985 ;
        RECT 67.650 161.765 67.925 162.245 ;
        RECT 68.095 161.745 68.395 162.075 ;
        RECT 60.935 160.885 61.430 161.425 ;
        RECT 62.150 161.255 62.320 161.425 ;
        RECT 61.820 161.085 62.320 161.255 ;
        RECT 58.995 159.865 59.165 160.625 ;
        RECT 59.345 159.695 59.675 160.455 ;
        RECT 59.845 159.865 60.115 160.770 ;
        RECT 60.435 159.695 60.765 160.845 ;
        RECT 60.935 160.715 61.945 160.885 ;
        RECT 60.935 159.865 61.105 160.715 ;
        RECT 61.275 159.695 61.605 160.495 ;
        RECT 61.775 159.865 61.945 160.715 ;
        RECT 62.150 160.845 62.320 161.085 ;
        RECT 62.490 161.015 62.870 161.255 ;
        RECT 62.150 160.675 62.865 160.845 ;
        RECT 62.125 159.695 62.365 160.495 ;
        RECT 62.535 159.865 62.865 160.675 ;
        RECT 63.045 159.695 63.335 160.860 ;
        RECT 63.965 160.785 64.715 161.305 ;
        RECT 64.885 160.955 65.635 161.475 ;
        RECT 65.820 161.425 67.470 161.595 ;
        RECT 65.820 160.915 66.225 161.425 ;
        RECT 66.395 161.085 67.535 161.255 ;
        RECT 63.965 159.695 65.635 160.785 ;
        RECT 65.820 160.745 66.575 160.915 ;
        RECT 65.860 159.695 66.145 160.565 ;
        RECT 66.315 160.495 66.575 160.745 ;
        RECT 67.365 160.835 67.535 161.085 ;
        RECT 67.705 161.005 68.055 161.575 ;
        RECT 68.225 160.835 68.395 161.745 ;
        RECT 68.565 161.495 69.775 162.245 ;
        RECT 67.365 160.665 68.395 160.835 ;
        RECT 66.315 160.325 67.435 160.495 ;
        RECT 66.315 159.865 66.575 160.325 ;
        RECT 66.750 159.695 67.005 160.155 ;
        RECT 67.175 159.865 67.435 160.325 ;
        RECT 67.605 159.695 67.915 160.495 ;
        RECT 68.085 159.865 68.395 160.665 ;
        RECT 68.565 160.785 69.085 161.325 ;
        RECT 69.255 160.955 69.775 161.495 ;
        RECT 69.950 161.405 70.210 162.245 ;
        RECT 70.385 161.500 70.640 162.075 ;
        RECT 70.810 161.865 71.140 162.245 ;
        RECT 71.355 161.695 71.525 162.075 ;
        RECT 70.810 161.525 71.525 161.695 ;
        RECT 68.565 159.695 69.775 160.785 ;
        RECT 69.950 159.695 70.210 160.845 ;
        RECT 70.385 160.770 70.555 161.500 ;
        RECT 70.810 161.335 70.980 161.525 ;
        RECT 72.245 161.475 73.915 162.245 ;
        RECT 74.090 161.700 79.435 162.245 ;
        RECT 70.725 161.005 70.980 161.335 ;
        RECT 70.810 160.795 70.980 161.005 ;
        RECT 71.260 160.975 71.615 161.345 ;
        RECT 70.385 159.865 70.640 160.770 ;
        RECT 70.810 160.625 71.525 160.795 ;
        RECT 70.810 159.695 71.140 160.455 ;
        RECT 71.355 159.865 71.525 160.625 ;
        RECT 72.245 160.785 72.995 161.305 ;
        RECT 73.165 160.955 73.915 161.475 ;
        RECT 72.245 159.695 73.915 160.785 ;
        RECT 75.680 160.130 76.030 161.380 ;
        RECT 77.510 160.870 77.850 161.700 ;
        RECT 79.880 161.435 80.125 162.040 ;
        RECT 80.345 161.710 80.855 162.245 ;
        RECT 79.605 161.265 80.835 161.435 ;
        RECT 79.605 160.455 79.945 161.265 ;
        RECT 80.115 160.700 80.865 160.890 ;
        RECT 74.090 159.695 79.435 160.130 ;
        RECT 79.605 160.045 80.120 160.455 ;
        RECT 80.355 159.695 80.525 160.455 ;
        RECT 80.695 160.035 80.865 160.700 ;
        RECT 81.035 160.715 81.225 162.075 ;
        RECT 81.395 161.225 81.670 162.075 ;
        RECT 81.860 161.710 82.390 162.075 ;
        RECT 82.815 161.845 83.145 162.245 ;
        RECT 82.215 161.675 82.390 161.710 ;
        RECT 81.395 161.055 81.675 161.225 ;
        RECT 81.395 160.915 81.670 161.055 ;
        RECT 81.875 160.715 82.045 161.515 ;
        RECT 81.035 160.545 82.045 160.715 ;
        RECT 82.215 161.505 83.145 161.675 ;
        RECT 83.315 161.505 83.570 162.075 ;
        RECT 82.215 160.375 82.385 161.505 ;
        RECT 82.975 161.335 83.145 161.505 ;
        RECT 81.260 160.205 82.385 160.375 ;
        RECT 82.555 161.005 82.750 161.335 ;
        RECT 82.975 161.005 83.230 161.335 ;
        RECT 82.555 160.035 82.725 161.005 ;
        RECT 83.400 160.835 83.570 161.505 ;
        RECT 84.725 161.425 84.935 162.245 ;
        RECT 85.105 161.445 85.435 162.075 ;
        RECT 85.105 160.845 85.355 161.445 ;
        RECT 85.605 161.425 85.835 162.245 ;
        RECT 87.055 161.695 87.225 162.075 ;
        RECT 87.405 161.865 87.735 162.245 ;
        RECT 87.055 161.525 87.720 161.695 ;
        RECT 87.915 161.570 88.175 162.075 ;
        RECT 85.525 161.005 85.855 161.255 ;
        RECT 86.985 160.975 87.315 161.345 ;
        RECT 87.550 161.270 87.720 161.525 ;
        RECT 87.550 160.940 87.835 161.270 ;
        RECT 80.695 159.865 82.725 160.035 ;
        RECT 82.895 159.695 83.065 160.835 ;
        RECT 83.235 159.865 83.570 160.835 ;
        RECT 84.725 159.695 84.935 160.835 ;
        RECT 85.105 159.865 85.435 160.845 ;
        RECT 85.605 159.695 85.835 160.835 ;
        RECT 87.550 160.795 87.720 160.940 ;
        RECT 87.055 160.625 87.720 160.795 ;
        RECT 88.005 160.770 88.175 161.570 ;
        RECT 88.805 161.520 89.095 162.245 ;
        RECT 89.265 161.495 90.475 162.245 ;
        RECT 87.055 159.865 87.225 160.625 ;
        RECT 87.405 159.695 87.735 160.455 ;
        RECT 87.905 159.865 88.175 160.770 ;
        RECT 88.805 159.695 89.095 160.860 ;
        RECT 89.265 160.785 89.785 161.325 ;
        RECT 89.955 160.955 90.475 161.495 ;
        RECT 91.020 161.535 91.275 162.065 ;
        RECT 91.455 161.785 91.740 162.245 ;
        RECT 89.265 159.695 90.475 160.785 ;
        RECT 91.020 160.675 91.200 161.535 ;
        RECT 91.920 161.335 92.170 161.985 ;
        RECT 91.370 161.005 92.170 161.335 ;
        RECT 91.020 160.545 91.275 160.675 ;
        RECT 90.935 160.375 91.275 160.545 ;
        RECT 91.020 160.005 91.275 160.375 ;
        RECT 91.455 159.695 91.740 160.495 ;
        RECT 91.920 160.415 92.170 161.005 ;
        RECT 92.370 161.650 92.690 161.980 ;
        RECT 92.870 161.765 93.530 162.245 ;
        RECT 93.730 161.855 94.580 162.025 ;
        RECT 92.370 160.755 92.560 161.650 ;
        RECT 92.880 161.325 93.540 161.595 ;
        RECT 93.210 161.265 93.540 161.325 ;
        RECT 92.730 161.095 93.060 161.155 ;
        RECT 93.730 161.095 93.900 161.855 ;
        RECT 95.140 161.785 95.460 162.245 ;
        RECT 95.660 161.605 95.910 162.035 ;
        RECT 96.200 161.805 96.610 162.245 ;
        RECT 96.780 161.865 97.795 162.065 ;
        RECT 94.070 161.435 95.320 161.605 ;
        RECT 94.070 161.315 94.400 161.435 ;
        RECT 92.730 160.925 94.630 161.095 ;
        RECT 92.370 160.585 94.290 160.755 ;
        RECT 92.370 160.565 92.690 160.585 ;
        RECT 91.920 159.905 92.250 160.415 ;
        RECT 92.520 159.955 92.690 160.565 ;
        RECT 94.460 160.415 94.630 160.925 ;
        RECT 94.800 160.855 94.980 161.265 ;
        RECT 95.150 160.675 95.320 161.435 ;
        RECT 92.860 159.695 93.190 160.385 ;
        RECT 93.420 160.245 94.630 160.415 ;
        RECT 94.800 160.365 95.320 160.675 ;
        RECT 95.490 161.265 95.910 161.605 ;
        RECT 96.200 161.265 96.610 161.595 ;
        RECT 95.490 160.495 95.680 161.265 ;
        RECT 96.780 161.135 96.950 161.865 ;
        RECT 98.095 161.695 98.265 162.025 ;
        RECT 98.435 161.865 98.765 162.245 ;
        RECT 97.120 161.315 97.470 161.685 ;
        RECT 96.780 161.095 97.200 161.135 ;
        RECT 95.850 160.925 97.200 161.095 ;
        RECT 95.850 160.765 96.100 160.925 ;
        RECT 96.610 160.495 96.860 160.755 ;
        RECT 95.490 160.245 96.860 160.495 ;
        RECT 93.420 159.955 93.660 160.245 ;
        RECT 94.460 160.165 94.630 160.245 ;
        RECT 93.860 159.695 94.280 160.075 ;
        RECT 94.460 159.915 95.090 160.165 ;
        RECT 95.560 159.695 95.890 160.075 ;
        RECT 96.060 159.955 96.230 160.245 ;
        RECT 97.030 160.080 97.200 160.925 ;
        RECT 97.650 160.755 97.870 161.625 ;
        RECT 98.095 161.505 98.790 161.695 ;
        RECT 97.370 160.375 97.870 160.755 ;
        RECT 98.040 160.705 98.450 161.325 ;
        RECT 98.620 160.535 98.790 161.505 ;
        RECT 98.095 160.365 98.790 160.535 ;
        RECT 96.410 159.695 96.790 160.075 ;
        RECT 97.030 159.910 97.860 160.080 ;
        RECT 98.095 159.865 98.265 160.365 ;
        RECT 98.435 159.695 98.765 160.195 ;
        RECT 98.980 159.865 99.205 161.985 ;
        RECT 99.375 161.865 99.705 162.245 ;
        RECT 99.875 161.695 100.045 161.985 ;
        RECT 99.380 161.525 100.045 161.695 ;
        RECT 100.305 161.570 100.565 162.075 ;
        RECT 100.745 161.865 101.075 162.245 ;
        RECT 101.255 161.695 101.425 162.075 ;
        RECT 99.380 160.535 99.610 161.525 ;
        RECT 99.780 160.705 100.130 161.355 ;
        RECT 100.305 160.770 100.475 161.570 ;
        RECT 100.760 161.525 101.425 161.695 ;
        RECT 100.760 161.270 100.930 161.525 ;
        RECT 102.605 161.475 106.115 162.245 ;
        RECT 106.375 161.695 106.545 162.075 ;
        RECT 106.725 161.865 107.055 162.245 ;
        RECT 106.375 161.525 107.040 161.695 ;
        RECT 107.235 161.570 107.495 162.075 ;
        RECT 100.645 160.940 100.930 161.270 ;
        RECT 101.165 160.975 101.495 161.345 ;
        RECT 100.760 160.795 100.930 160.940 ;
        RECT 99.380 160.365 100.045 160.535 ;
        RECT 99.375 159.695 99.705 160.195 ;
        RECT 99.875 159.865 100.045 160.365 ;
        RECT 100.305 159.865 100.575 160.770 ;
        RECT 100.760 160.625 101.425 160.795 ;
        RECT 100.745 159.695 101.075 160.455 ;
        RECT 101.255 159.865 101.425 160.625 ;
        RECT 102.605 160.785 104.295 161.305 ;
        RECT 104.465 160.955 106.115 161.475 ;
        RECT 106.305 160.975 106.635 161.345 ;
        RECT 106.870 161.270 107.040 161.525 ;
        RECT 106.870 160.940 107.155 161.270 ;
        RECT 106.870 160.795 107.040 160.940 ;
        RECT 102.605 159.695 106.115 160.785 ;
        RECT 106.375 160.625 107.040 160.795 ;
        RECT 107.325 160.770 107.495 161.570 ;
        RECT 107.665 161.495 108.875 162.245 ;
        RECT 109.050 161.700 114.395 162.245 ;
        RECT 106.375 159.865 106.545 160.625 ;
        RECT 106.725 159.695 107.055 160.455 ;
        RECT 107.225 159.865 107.495 160.770 ;
        RECT 107.665 160.785 108.185 161.325 ;
        RECT 108.355 160.955 108.875 161.495 ;
        RECT 107.665 159.695 108.875 160.785 ;
        RECT 110.640 160.130 110.990 161.380 ;
        RECT 112.470 160.870 112.810 161.700 ;
        RECT 114.565 161.520 114.855 162.245 ;
        RECT 115.485 161.475 117.155 162.245 ;
        RECT 109.050 159.695 114.395 160.130 ;
        RECT 114.565 159.695 114.855 160.860 ;
        RECT 115.485 160.785 116.235 161.305 ;
        RECT 116.405 160.955 117.155 161.475 ;
        RECT 117.475 161.445 117.805 162.245 ;
        RECT 117.975 161.595 118.145 162.075 ;
        RECT 118.315 161.765 118.645 162.245 ;
        RECT 118.815 161.595 118.985 162.075 ;
        RECT 119.235 161.765 119.475 162.245 ;
        RECT 119.655 161.595 119.825 162.075 ;
        RECT 121.010 161.700 126.355 162.245 ;
        RECT 117.975 161.425 118.985 161.595 ;
        RECT 119.190 161.425 119.825 161.595 ;
        RECT 117.975 160.885 118.470 161.425 ;
        RECT 119.190 161.255 119.360 161.425 ;
        RECT 118.860 161.085 119.360 161.255 ;
        RECT 115.485 159.695 117.155 160.785 ;
        RECT 117.475 159.695 117.805 160.845 ;
        RECT 117.975 160.715 118.985 160.885 ;
        RECT 117.975 159.865 118.145 160.715 ;
        RECT 118.315 159.695 118.645 160.495 ;
        RECT 118.815 159.865 118.985 160.715 ;
        RECT 119.190 160.845 119.360 161.085 ;
        RECT 119.530 161.015 119.910 161.255 ;
        RECT 119.190 160.675 119.905 160.845 ;
        RECT 119.165 159.695 119.405 160.495 ;
        RECT 119.575 159.865 119.905 160.675 ;
        RECT 122.600 160.130 122.950 161.380 ;
        RECT 124.430 160.870 124.770 161.700 ;
        RECT 126.525 161.495 127.735 162.245 ;
        RECT 126.525 160.785 127.045 161.325 ;
        RECT 127.215 160.955 127.735 161.495 ;
        RECT 121.010 159.695 126.355 160.130 ;
        RECT 126.525 159.695 127.735 160.785 ;
        RECT 14.660 159.525 127.820 159.695 ;
        RECT 14.745 158.435 15.955 159.525 ;
        RECT 14.745 157.725 15.265 158.265 ;
        RECT 15.435 157.895 15.955 158.435 ;
        RECT 16.125 158.435 18.715 159.525 ;
        RECT 18.975 158.595 19.145 159.355 ;
        RECT 19.325 158.765 19.655 159.525 ;
        RECT 16.125 157.915 17.335 158.435 ;
        RECT 18.975 158.425 19.640 158.595 ;
        RECT 19.825 158.450 20.095 159.355 ;
        RECT 19.470 158.280 19.640 158.425 ;
        RECT 17.505 157.745 18.715 158.265 ;
        RECT 18.905 157.875 19.235 158.245 ;
        RECT 19.470 157.950 19.755 158.280 ;
        RECT 14.745 156.975 15.955 157.725 ;
        RECT 16.125 156.975 18.715 157.745 ;
        RECT 19.470 157.695 19.640 157.950 ;
        RECT 18.975 157.525 19.640 157.695 ;
        RECT 19.925 157.650 20.095 158.450 ;
        RECT 18.975 157.145 19.145 157.525 ;
        RECT 19.325 156.975 19.655 157.355 ;
        RECT 19.835 157.145 20.095 157.650 ;
        RECT 20.270 158.385 20.605 159.355 ;
        RECT 20.775 158.385 20.945 159.525 ;
        RECT 21.115 159.185 23.145 159.355 ;
        RECT 20.270 157.715 20.440 158.385 ;
        RECT 21.115 158.215 21.285 159.185 ;
        RECT 20.610 157.885 20.865 158.215 ;
        RECT 21.090 157.885 21.285 158.215 ;
        RECT 21.455 158.845 22.580 159.015 ;
        RECT 20.695 157.715 20.865 157.885 ;
        RECT 21.455 157.715 21.625 158.845 ;
        RECT 20.270 157.145 20.525 157.715 ;
        RECT 20.695 157.545 21.625 157.715 ;
        RECT 21.795 158.505 22.805 158.675 ;
        RECT 21.795 157.705 21.965 158.505 ;
        RECT 21.450 157.510 21.625 157.545 ;
        RECT 20.695 156.975 21.025 157.375 ;
        RECT 21.450 157.145 21.980 157.510 ;
        RECT 22.170 157.485 22.445 158.305 ;
        RECT 22.165 157.315 22.445 157.485 ;
        RECT 22.170 157.145 22.445 157.315 ;
        RECT 22.615 157.145 22.805 158.505 ;
        RECT 22.975 158.520 23.145 159.185 ;
        RECT 23.315 158.765 23.485 159.525 ;
        RECT 23.720 158.765 24.235 159.175 ;
        RECT 22.975 158.330 23.725 158.520 ;
        RECT 23.895 157.955 24.235 158.765 ;
        RECT 24.405 158.360 24.695 159.525 ;
        RECT 24.865 158.435 26.075 159.525 ;
        RECT 26.250 159.090 31.595 159.525 ;
        RECT 23.005 157.785 24.235 157.955 ;
        RECT 24.865 157.895 25.385 158.435 ;
        RECT 22.985 156.975 23.495 157.510 ;
        RECT 23.715 157.180 23.960 157.785 ;
        RECT 25.555 157.725 26.075 158.265 ;
        RECT 27.840 157.840 28.190 159.090 ;
        RECT 31.805 158.385 32.035 159.525 ;
        RECT 32.205 158.375 32.535 159.355 ;
        RECT 32.705 158.385 32.915 159.525 ;
        RECT 33.145 158.765 33.660 159.175 ;
        RECT 33.895 158.765 34.065 159.525 ;
        RECT 34.235 159.185 36.265 159.355 ;
        RECT 24.405 156.975 24.695 157.700 ;
        RECT 24.865 156.975 26.075 157.725 ;
        RECT 29.670 157.520 30.010 158.350 ;
        RECT 31.785 157.965 32.115 158.215 ;
        RECT 26.250 156.975 31.595 157.520 ;
        RECT 31.805 156.975 32.035 157.795 ;
        RECT 32.285 157.775 32.535 158.375 ;
        RECT 33.145 157.955 33.485 158.765 ;
        RECT 34.235 158.520 34.405 159.185 ;
        RECT 34.800 158.845 35.925 159.015 ;
        RECT 33.655 158.330 34.405 158.520 ;
        RECT 34.575 158.505 35.585 158.675 ;
        RECT 32.205 157.145 32.535 157.775 ;
        RECT 32.705 156.975 32.915 157.795 ;
        RECT 33.145 157.785 34.375 157.955 ;
        RECT 33.420 157.180 33.665 157.785 ;
        RECT 33.885 156.975 34.395 157.510 ;
        RECT 34.575 157.145 34.765 158.505 ;
        RECT 34.935 157.825 35.210 158.305 ;
        RECT 34.935 157.655 35.215 157.825 ;
        RECT 35.415 157.705 35.585 158.505 ;
        RECT 35.755 157.715 35.925 158.845 ;
        RECT 36.095 158.215 36.265 159.185 ;
        RECT 36.435 158.385 36.605 159.525 ;
        RECT 36.775 158.385 37.110 159.355 ;
        RECT 36.095 157.885 36.290 158.215 ;
        RECT 36.515 157.885 36.770 158.215 ;
        RECT 36.515 157.715 36.685 157.885 ;
        RECT 36.940 157.715 37.110 158.385 ;
        RECT 37.285 158.435 39.875 159.525 ;
        RECT 37.285 157.915 38.495 158.435 ;
        RECT 40.045 158.385 40.385 159.355 ;
        RECT 40.555 158.385 40.725 159.525 ;
        RECT 40.995 158.725 41.245 159.525 ;
        RECT 41.890 158.555 42.220 159.355 ;
        RECT 42.520 158.725 42.850 159.525 ;
        RECT 43.020 158.555 43.350 159.355 ;
        RECT 40.915 158.385 43.350 158.555 ;
        RECT 44.185 158.435 45.855 159.525 ;
        RECT 46.025 158.765 46.540 159.175 ;
        RECT 46.775 158.765 46.945 159.525 ;
        RECT 47.115 159.185 49.145 159.355 ;
        RECT 38.665 157.745 39.875 158.265 ;
        RECT 34.935 157.145 35.210 157.655 ;
        RECT 35.755 157.545 36.685 157.715 ;
        RECT 35.755 157.510 35.930 157.545 ;
        RECT 35.400 157.145 35.930 157.510 ;
        RECT 36.355 156.975 36.685 157.375 ;
        RECT 36.855 157.145 37.110 157.715 ;
        RECT 37.285 156.975 39.875 157.745 ;
        RECT 40.045 157.775 40.220 158.385 ;
        RECT 40.915 158.135 41.085 158.385 ;
        RECT 40.390 157.965 41.085 158.135 ;
        RECT 41.260 157.965 41.680 158.165 ;
        RECT 41.850 157.965 42.180 158.165 ;
        RECT 42.350 157.965 42.680 158.165 ;
        RECT 40.045 157.145 40.385 157.775 ;
        RECT 40.555 156.975 40.805 157.775 ;
        RECT 40.995 157.625 42.220 157.795 ;
        RECT 40.995 157.145 41.325 157.625 ;
        RECT 41.495 156.975 41.720 157.435 ;
        RECT 41.890 157.145 42.220 157.625 ;
        RECT 42.850 157.755 43.020 158.385 ;
        RECT 43.205 157.965 43.555 158.215 ;
        RECT 44.185 157.915 44.935 158.435 ;
        RECT 42.850 157.145 43.350 157.755 ;
        RECT 45.105 157.745 45.855 158.265 ;
        RECT 46.025 157.955 46.365 158.765 ;
        RECT 47.115 158.520 47.285 159.185 ;
        RECT 47.680 158.845 48.805 159.015 ;
        RECT 46.535 158.330 47.285 158.520 ;
        RECT 47.455 158.505 48.465 158.675 ;
        RECT 46.025 157.785 47.255 157.955 ;
        RECT 44.185 156.975 45.855 157.745 ;
        RECT 46.300 157.180 46.545 157.785 ;
        RECT 46.765 156.975 47.275 157.510 ;
        RECT 47.455 157.145 47.645 158.505 ;
        RECT 47.815 157.485 48.090 158.305 ;
        RECT 48.295 157.705 48.465 158.505 ;
        RECT 48.635 157.715 48.805 158.845 ;
        RECT 48.975 158.215 49.145 159.185 ;
        RECT 49.315 158.385 49.485 159.525 ;
        RECT 49.655 158.385 49.990 159.355 ;
        RECT 48.975 157.885 49.170 158.215 ;
        RECT 49.395 157.885 49.650 158.215 ;
        RECT 49.395 157.715 49.565 157.885 ;
        RECT 49.820 157.715 49.990 158.385 ;
        RECT 50.165 158.360 50.455 159.525 ;
        RECT 50.625 158.435 51.835 159.525 ;
        RECT 50.625 157.895 51.145 158.435 ;
        RECT 52.010 158.335 52.265 159.215 ;
        RECT 52.435 158.385 52.740 159.525 ;
        RECT 53.080 159.145 53.410 159.525 ;
        RECT 53.590 158.975 53.760 159.265 ;
        RECT 53.930 159.065 54.180 159.525 ;
        RECT 52.960 158.805 53.760 158.975 ;
        RECT 54.350 159.015 55.220 159.355 ;
        RECT 51.315 157.725 51.835 158.265 ;
        RECT 48.635 157.545 49.565 157.715 ;
        RECT 48.635 157.510 48.810 157.545 ;
        RECT 47.815 157.315 48.095 157.485 ;
        RECT 47.815 157.145 48.090 157.315 ;
        RECT 48.280 157.145 48.810 157.510 ;
        RECT 49.235 156.975 49.565 157.375 ;
        RECT 49.735 157.145 49.990 157.715 ;
        RECT 50.165 156.975 50.455 157.700 ;
        RECT 50.625 156.975 51.835 157.725 ;
        RECT 52.010 157.685 52.220 158.335 ;
        RECT 52.960 158.215 53.130 158.805 ;
        RECT 54.350 158.635 54.520 159.015 ;
        RECT 55.455 158.895 55.625 159.355 ;
        RECT 55.795 159.065 56.165 159.525 ;
        RECT 56.460 158.925 56.630 159.265 ;
        RECT 56.800 159.095 57.130 159.525 ;
        RECT 57.365 158.925 57.535 159.265 ;
        RECT 53.300 158.465 54.520 158.635 ;
        RECT 54.690 158.555 55.150 158.845 ;
        RECT 55.455 158.725 56.015 158.895 ;
        RECT 56.460 158.755 57.535 158.925 ;
        RECT 57.705 159.025 58.385 159.355 ;
        RECT 58.600 159.025 58.850 159.355 ;
        RECT 59.020 159.065 59.270 159.525 ;
        RECT 55.845 158.585 56.015 158.725 ;
        RECT 54.690 158.545 55.655 158.555 ;
        RECT 54.350 158.375 54.520 158.465 ;
        RECT 54.980 158.385 55.655 158.545 ;
        RECT 52.390 158.185 53.130 158.215 ;
        RECT 52.390 157.885 53.305 158.185 ;
        RECT 52.980 157.710 53.305 157.885 ;
        RECT 52.010 157.155 52.265 157.685 ;
        RECT 52.435 156.975 52.740 157.435 ;
        RECT 52.985 157.355 53.305 157.710 ;
        RECT 53.475 157.925 54.015 158.295 ;
        RECT 54.350 158.205 54.755 158.375 ;
        RECT 53.475 157.525 53.715 157.925 ;
        RECT 54.195 157.755 54.415 158.035 ;
        RECT 53.885 157.585 54.415 157.755 ;
        RECT 53.885 157.355 54.055 157.585 ;
        RECT 54.585 157.425 54.755 158.205 ;
        RECT 54.925 157.595 55.275 158.215 ;
        RECT 55.445 157.595 55.655 158.385 ;
        RECT 55.845 158.415 57.345 158.585 ;
        RECT 55.845 157.725 56.015 158.415 ;
        RECT 57.705 158.245 57.875 159.025 ;
        RECT 58.680 158.895 58.850 159.025 ;
        RECT 56.185 158.075 57.875 158.245 ;
        RECT 58.045 158.465 58.510 158.855 ;
        RECT 58.680 158.725 59.075 158.895 ;
        RECT 56.185 157.895 56.355 158.075 ;
        RECT 52.985 157.185 54.055 157.355 ;
        RECT 54.225 156.975 54.415 157.415 ;
        RECT 54.585 157.145 55.535 157.425 ;
        RECT 55.845 157.335 56.105 157.725 ;
        RECT 56.525 157.655 57.315 157.905 ;
        RECT 55.755 157.165 56.105 157.335 ;
        RECT 56.315 156.975 56.645 157.435 ;
        RECT 57.520 157.365 57.690 158.075 ;
        RECT 58.045 157.875 58.215 158.465 ;
        RECT 57.860 157.655 58.215 157.875 ;
        RECT 58.385 157.655 58.735 158.275 ;
        RECT 58.905 157.365 59.075 158.725 ;
        RECT 59.440 158.555 59.765 159.340 ;
        RECT 59.245 157.505 59.705 158.555 ;
        RECT 57.520 157.195 58.375 157.365 ;
        RECT 58.580 157.195 59.075 157.365 ;
        RECT 59.245 156.975 59.575 157.335 ;
        RECT 59.935 157.235 60.105 159.355 ;
        RECT 60.275 159.025 60.605 159.525 ;
        RECT 60.775 158.855 61.030 159.355 ;
        RECT 60.280 158.685 61.030 158.855 ;
        RECT 60.280 157.695 60.510 158.685 ;
        RECT 60.680 157.865 61.030 158.515 ;
        RECT 61.665 158.435 64.255 159.525 ;
        RECT 61.665 157.915 62.875 158.435 ;
        RECT 64.430 158.375 64.690 159.525 ;
        RECT 64.865 158.450 65.120 159.355 ;
        RECT 65.290 158.765 65.620 159.525 ;
        RECT 65.835 158.595 66.005 159.355 ;
        RECT 63.045 157.745 64.255 158.265 ;
        RECT 60.280 157.525 61.030 157.695 ;
        RECT 60.275 156.975 60.605 157.355 ;
        RECT 60.775 157.235 61.030 157.525 ;
        RECT 61.665 156.975 64.255 157.745 ;
        RECT 64.430 156.975 64.690 157.815 ;
        RECT 64.865 157.720 65.035 158.450 ;
        RECT 65.290 158.425 66.005 158.595 ;
        RECT 65.290 158.215 65.460 158.425 ;
        RECT 66.270 158.375 66.530 159.525 ;
        RECT 66.705 158.450 66.960 159.355 ;
        RECT 67.130 158.765 67.460 159.525 ;
        RECT 67.675 158.595 67.845 159.355 ;
        RECT 65.205 157.885 65.460 158.215 ;
        RECT 64.865 157.145 65.120 157.720 ;
        RECT 65.290 157.695 65.460 157.885 ;
        RECT 65.740 157.875 66.095 158.245 ;
        RECT 65.290 157.525 66.005 157.695 ;
        RECT 65.290 156.975 65.620 157.355 ;
        RECT 65.835 157.145 66.005 157.525 ;
        RECT 66.270 156.975 66.530 157.815 ;
        RECT 66.705 157.720 66.875 158.450 ;
        RECT 67.130 158.425 67.845 158.595 ;
        RECT 68.195 158.595 68.365 159.355 ;
        RECT 68.580 158.765 68.910 159.525 ;
        RECT 68.195 158.425 68.910 158.595 ;
        RECT 69.080 158.450 69.335 159.355 ;
        RECT 67.130 158.215 67.300 158.425 ;
        RECT 67.045 157.885 67.300 158.215 ;
        RECT 66.705 157.145 66.960 157.720 ;
        RECT 67.130 157.695 67.300 157.885 ;
        RECT 67.580 157.875 67.935 158.245 ;
        RECT 68.105 157.875 68.460 158.245 ;
        RECT 68.740 158.215 68.910 158.425 ;
        RECT 68.740 157.885 68.995 158.215 ;
        RECT 68.740 157.695 68.910 157.885 ;
        RECT 69.165 157.720 69.335 158.450 ;
        RECT 69.510 158.375 69.770 159.525 ;
        RECT 70.035 158.595 70.205 159.355 ;
        RECT 70.420 158.765 70.750 159.525 ;
        RECT 70.035 158.425 70.750 158.595 ;
        RECT 70.920 158.450 71.175 159.355 ;
        RECT 69.945 157.875 70.300 158.245 ;
        RECT 70.580 158.215 70.750 158.425 ;
        RECT 70.580 157.885 70.835 158.215 ;
        RECT 67.130 157.525 67.845 157.695 ;
        RECT 67.130 156.975 67.460 157.355 ;
        RECT 67.675 157.145 67.845 157.525 ;
        RECT 68.195 157.525 68.910 157.695 ;
        RECT 68.195 157.145 68.365 157.525 ;
        RECT 68.580 156.975 68.910 157.355 ;
        RECT 69.080 157.145 69.335 157.720 ;
        RECT 69.510 156.975 69.770 157.815 ;
        RECT 70.580 157.695 70.750 157.885 ;
        RECT 71.005 157.720 71.175 158.450 ;
        RECT 71.350 158.375 71.610 159.525 ;
        RECT 72.245 158.435 75.755 159.525 ;
        RECT 72.245 157.915 73.935 158.435 ;
        RECT 75.925 158.360 76.215 159.525 ;
        RECT 77.305 158.435 80.815 159.525 ;
        RECT 81.360 158.545 81.615 159.215 ;
        RECT 81.795 158.725 82.080 159.525 ;
        RECT 82.260 158.805 82.590 159.315 ;
        RECT 70.035 157.525 70.750 157.695 ;
        RECT 70.035 157.145 70.205 157.525 ;
        RECT 70.420 156.975 70.750 157.355 ;
        RECT 70.920 157.145 71.175 157.720 ;
        RECT 71.350 156.975 71.610 157.815 ;
        RECT 74.105 157.745 75.755 158.265 ;
        RECT 77.305 157.915 78.995 158.435 ;
        RECT 79.165 157.745 80.815 158.265 ;
        RECT 81.360 157.825 81.540 158.545 ;
        RECT 82.260 158.215 82.510 158.805 ;
        RECT 82.860 158.655 83.030 159.265 ;
        RECT 83.200 158.835 83.530 159.525 ;
        RECT 83.760 158.975 84.000 159.265 ;
        RECT 84.200 159.145 84.620 159.525 ;
        RECT 84.800 159.055 85.430 159.305 ;
        RECT 85.900 159.145 86.230 159.525 ;
        RECT 84.800 158.975 84.970 159.055 ;
        RECT 86.400 158.975 86.570 159.265 ;
        RECT 86.750 159.145 87.130 159.525 ;
        RECT 87.370 159.140 88.200 159.310 ;
        RECT 83.760 158.805 84.970 158.975 ;
        RECT 81.710 157.885 82.510 158.215 ;
        RECT 72.245 156.975 75.755 157.745 ;
        RECT 75.925 156.975 76.215 157.700 ;
        RECT 77.305 156.975 80.815 157.745 ;
        RECT 81.275 157.685 81.540 157.825 ;
        RECT 81.275 157.655 81.615 157.685 ;
        RECT 81.360 157.155 81.615 157.655 ;
        RECT 81.795 156.975 82.080 157.435 ;
        RECT 82.260 157.235 82.510 157.885 ;
        RECT 82.710 158.635 83.030 158.655 ;
        RECT 82.710 158.465 84.630 158.635 ;
        RECT 82.710 157.570 82.900 158.465 ;
        RECT 84.800 158.295 84.970 158.805 ;
        RECT 85.140 158.545 85.660 158.855 ;
        RECT 83.070 158.125 84.970 158.295 ;
        RECT 83.070 158.065 83.400 158.125 ;
        RECT 83.550 157.895 83.880 157.955 ;
        RECT 83.220 157.625 83.880 157.895 ;
        RECT 82.710 157.240 83.030 157.570 ;
        RECT 83.210 156.975 83.870 157.455 ;
        RECT 84.070 157.365 84.240 158.125 ;
        RECT 85.140 157.955 85.320 158.365 ;
        RECT 84.410 157.785 84.740 157.905 ;
        RECT 85.490 157.785 85.660 158.545 ;
        RECT 84.410 157.615 85.660 157.785 ;
        RECT 85.830 158.725 87.200 158.975 ;
        RECT 85.830 157.955 86.020 158.725 ;
        RECT 86.950 158.465 87.200 158.725 ;
        RECT 86.190 158.295 86.440 158.455 ;
        RECT 87.370 158.295 87.540 159.140 ;
        RECT 88.435 158.855 88.605 159.355 ;
        RECT 88.775 159.025 89.105 159.525 ;
        RECT 87.710 158.465 88.210 158.845 ;
        RECT 88.435 158.685 89.130 158.855 ;
        RECT 86.190 158.125 87.540 158.295 ;
        RECT 87.120 158.085 87.540 158.125 ;
        RECT 85.830 157.615 86.250 157.955 ;
        RECT 86.540 157.625 86.950 157.955 ;
        RECT 84.070 157.195 84.920 157.365 ;
        RECT 85.480 156.975 85.800 157.435 ;
        RECT 86.000 157.185 86.250 157.615 ;
        RECT 86.540 156.975 86.950 157.415 ;
        RECT 87.120 157.355 87.290 158.085 ;
        RECT 87.460 157.535 87.810 157.905 ;
        RECT 87.990 157.595 88.210 158.465 ;
        RECT 88.380 157.895 88.790 158.515 ;
        RECT 88.960 157.715 89.130 158.685 ;
        RECT 88.435 157.525 89.130 157.715 ;
        RECT 87.120 157.155 88.135 157.355 ;
        RECT 88.435 157.195 88.605 157.525 ;
        RECT 88.775 156.975 89.105 157.355 ;
        RECT 89.320 157.235 89.545 159.355 ;
        RECT 89.715 159.025 90.045 159.525 ;
        RECT 90.215 158.855 90.385 159.355 ;
        RECT 89.720 158.685 90.385 158.855 ;
        RECT 89.720 157.695 89.950 158.685 ;
        RECT 90.120 157.865 90.470 158.515 ;
        RECT 90.645 158.435 94.155 159.525 ;
        RECT 90.645 157.915 92.335 158.435 ;
        RECT 94.385 158.385 94.595 159.525 ;
        RECT 94.765 158.375 95.095 159.355 ;
        RECT 95.265 158.385 95.495 159.525 ;
        RECT 96.170 159.090 101.515 159.525 ;
        RECT 92.505 157.745 94.155 158.265 ;
        RECT 89.720 157.525 90.385 157.695 ;
        RECT 89.715 156.975 90.045 157.355 ;
        RECT 90.215 157.235 90.385 157.525 ;
        RECT 90.645 156.975 94.155 157.745 ;
        RECT 94.385 156.975 94.595 157.795 ;
        RECT 94.765 157.775 95.015 158.375 ;
        RECT 95.185 157.965 95.515 158.215 ;
        RECT 97.760 157.840 98.110 159.090 ;
        RECT 101.685 158.360 101.975 159.525 ;
        RECT 102.605 158.435 104.275 159.525 ;
        RECT 94.765 157.145 95.095 157.775 ;
        RECT 95.265 156.975 95.495 157.795 ;
        RECT 99.590 157.520 99.930 158.350 ;
        RECT 102.605 157.915 103.355 158.435 ;
        RECT 104.445 158.385 104.785 159.355 ;
        RECT 104.955 158.385 105.125 159.525 ;
        RECT 105.395 158.725 105.645 159.525 ;
        RECT 106.290 158.555 106.620 159.355 ;
        RECT 106.920 158.725 107.250 159.525 ;
        RECT 107.420 158.555 107.750 159.355 ;
        RECT 105.315 158.385 107.750 158.555 ;
        RECT 108.585 158.435 110.255 159.525 ;
        RECT 110.430 159.090 115.775 159.525 ;
        RECT 103.525 157.745 104.275 158.265 ;
        RECT 96.170 156.975 101.515 157.520 ;
        RECT 101.685 156.975 101.975 157.700 ;
        RECT 102.605 156.975 104.275 157.745 ;
        RECT 104.445 157.775 104.620 158.385 ;
        RECT 105.315 158.135 105.485 158.385 ;
        RECT 104.790 157.965 105.485 158.135 ;
        RECT 105.660 157.965 106.080 158.165 ;
        RECT 106.250 157.965 106.580 158.165 ;
        RECT 106.750 157.965 107.080 158.165 ;
        RECT 104.445 157.145 104.785 157.775 ;
        RECT 104.955 156.975 105.205 157.775 ;
        RECT 105.395 157.625 106.620 157.795 ;
        RECT 105.395 157.145 105.725 157.625 ;
        RECT 105.895 156.975 106.120 157.435 ;
        RECT 106.290 157.145 106.620 157.625 ;
        RECT 107.250 157.755 107.420 158.385 ;
        RECT 107.605 157.965 107.955 158.215 ;
        RECT 108.585 157.915 109.335 158.435 ;
        RECT 107.250 157.145 107.750 157.755 ;
        RECT 109.505 157.745 110.255 158.265 ;
        RECT 112.020 157.840 112.370 159.090 ;
        RECT 115.955 158.545 116.285 159.355 ;
        RECT 116.455 158.725 116.695 159.525 ;
        RECT 115.955 158.375 116.670 158.545 ;
        RECT 108.585 156.975 110.255 157.745 ;
        RECT 113.850 157.520 114.190 158.350 ;
        RECT 115.950 157.965 116.330 158.205 ;
        RECT 116.500 158.135 116.670 158.375 ;
        RECT 116.875 158.505 117.045 159.355 ;
        RECT 117.215 158.725 117.545 159.525 ;
        RECT 117.715 158.505 117.885 159.355 ;
        RECT 116.875 158.335 117.885 158.505 ;
        RECT 118.055 158.375 118.385 159.525 ;
        RECT 119.165 158.435 120.835 159.525 ;
        RECT 121.010 159.090 126.355 159.525 ;
        RECT 116.500 157.965 117.000 158.135 ;
        RECT 116.500 157.795 116.670 157.965 ;
        RECT 117.390 157.795 117.885 158.335 ;
        RECT 119.165 157.915 119.915 158.435 ;
        RECT 116.035 157.625 116.670 157.795 ;
        RECT 116.875 157.625 117.885 157.795 ;
        RECT 110.430 156.975 115.775 157.520 ;
        RECT 116.035 157.145 116.205 157.625 ;
        RECT 116.385 156.975 116.625 157.455 ;
        RECT 116.875 157.145 117.045 157.625 ;
        RECT 117.215 156.975 117.545 157.455 ;
        RECT 117.715 157.145 117.885 157.625 ;
        RECT 118.055 156.975 118.385 157.775 ;
        RECT 120.085 157.745 120.835 158.265 ;
        RECT 122.600 157.840 122.950 159.090 ;
        RECT 126.525 158.435 127.735 159.525 ;
        RECT 119.165 156.975 120.835 157.745 ;
        RECT 124.430 157.520 124.770 158.350 ;
        RECT 126.525 157.895 127.045 158.435 ;
        RECT 127.215 157.725 127.735 158.265 ;
        RECT 121.010 156.975 126.355 157.520 ;
        RECT 126.525 156.975 127.735 157.725 ;
        RECT 14.660 156.805 127.820 156.975 ;
        RECT 14.745 156.055 15.955 156.805 ;
        RECT 17.420 156.095 17.675 156.625 ;
        RECT 17.855 156.345 18.140 156.805 ;
        RECT 14.745 155.515 15.265 156.055 ;
        RECT 15.435 155.345 15.955 155.885 ;
        RECT 14.745 154.255 15.955 155.345 ;
        RECT 17.420 155.235 17.600 156.095 ;
        RECT 18.320 155.895 18.570 156.545 ;
        RECT 17.770 155.565 18.570 155.895 ;
        RECT 17.420 154.765 17.675 155.235 ;
        RECT 17.335 154.595 17.675 154.765 ;
        RECT 17.420 154.565 17.675 154.595 ;
        RECT 17.855 154.255 18.140 155.055 ;
        RECT 18.320 154.975 18.570 155.565 ;
        RECT 18.770 156.210 19.090 156.540 ;
        RECT 19.270 156.325 19.930 156.805 ;
        RECT 20.130 156.415 20.980 156.585 ;
        RECT 18.770 155.315 18.960 156.210 ;
        RECT 19.280 155.885 19.940 156.155 ;
        RECT 19.610 155.825 19.940 155.885 ;
        RECT 19.130 155.655 19.460 155.715 ;
        RECT 20.130 155.655 20.300 156.415 ;
        RECT 21.540 156.345 21.860 156.805 ;
        RECT 22.060 156.165 22.310 156.595 ;
        RECT 22.600 156.365 23.010 156.805 ;
        RECT 23.180 156.425 24.195 156.625 ;
        RECT 20.470 155.995 21.720 156.165 ;
        RECT 20.470 155.875 20.800 155.995 ;
        RECT 19.130 155.485 21.030 155.655 ;
        RECT 18.770 155.145 20.690 155.315 ;
        RECT 18.770 155.125 19.090 155.145 ;
        RECT 18.320 154.465 18.650 154.975 ;
        RECT 18.920 154.515 19.090 155.125 ;
        RECT 20.860 154.975 21.030 155.485 ;
        RECT 21.200 155.415 21.380 155.825 ;
        RECT 21.550 155.235 21.720 155.995 ;
        RECT 19.260 154.255 19.590 154.945 ;
        RECT 19.820 154.805 21.030 154.975 ;
        RECT 21.200 154.925 21.720 155.235 ;
        RECT 21.890 155.825 22.310 156.165 ;
        RECT 22.600 155.825 23.010 156.155 ;
        RECT 21.890 155.055 22.080 155.825 ;
        RECT 23.180 155.695 23.350 156.425 ;
        RECT 24.495 156.255 24.665 156.585 ;
        RECT 24.835 156.425 25.165 156.805 ;
        RECT 23.520 155.875 23.870 156.245 ;
        RECT 23.180 155.655 23.600 155.695 ;
        RECT 22.250 155.485 23.600 155.655 ;
        RECT 22.250 155.325 22.500 155.485 ;
        RECT 23.010 155.055 23.260 155.315 ;
        RECT 21.890 154.805 23.260 155.055 ;
        RECT 19.820 154.515 20.060 154.805 ;
        RECT 20.860 154.725 21.030 154.805 ;
        RECT 20.260 154.255 20.680 154.635 ;
        RECT 20.860 154.475 21.490 154.725 ;
        RECT 21.960 154.255 22.290 154.635 ;
        RECT 22.460 154.515 22.630 154.805 ;
        RECT 23.430 154.640 23.600 155.485 ;
        RECT 24.050 155.315 24.270 156.185 ;
        RECT 24.495 156.065 25.190 156.255 ;
        RECT 23.770 154.935 24.270 155.315 ;
        RECT 24.440 155.265 24.850 155.885 ;
        RECT 25.020 155.095 25.190 156.065 ;
        RECT 24.495 154.925 25.190 155.095 ;
        RECT 22.810 154.255 23.190 154.635 ;
        RECT 23.430 154.470 24.260 154.640 ;
        RECT 24.495 154.425 24.665 154.925 ;
        RECT 24.835 154.255 25.165 154.755 ;
        RECT 25.380 154.425 25.605 156.545 ;
        RECT 25.775 156.425 26.105 156.805 ;
        RECT 26.275 156.255 26.445 156.545 ;
        RECT 25.780 156.085 26.445 156.255 ;
        RECT 25.780 155.095 26.010 156.085 ;
        RECT 26.705 156.055 27.915 156.805 ;
        RECT 26.180 155.265 26.530 155.915 ;
        RECT 26.705 155.345 27.225 155.885 ;
        RECT 27.395 155.515 27.915 156.055 ;
        RECT 28.085 156.035 31.595 156.805 ;
        RECT 31.770 156.260 37.115 156.805 ;
        RECT 28.085 155.345 29.775 155.865 ;
        RECT 29.945 155.515 31.595 156.035 ;
        RECT 25.780 154.925 26.445 155.095 ;
        RECT 25.775 154.255 26.105 154.755 ;
        RECT 26.275 154.425 26.445 154.925 ;
        RECT 26.705 154.255 27.915 155.345 ;
        RECT 28.085 154.255 31.595 155.345 ;
        RECT 33.360 154.690 33.710 155.940 ;
        RECT 35.190 155.430 35.530 156.260 ;
        RECT 37.285 156.080 37.575 156.805 ;
        RECT 38.205 156.035 39.875 156.805 ;
        RECT 40.050 156.260 45.395 156.805 ;
        RECT 45.570 156.260 50.915 156.805 ;
        RECT 31.770 154.255 37.115 154.690 ;
        RECT 37.285 154.255 37.575 155.420 ;
        RECT 38.205 155.345 38.955 155.865 ;
        RECT 39.125 155.515 39.875 156.035 ;
        RECT 38.205 154.255 39.875 155.345 ;
        RECT 41.640 154.690 41.990 155.940 ;
        RECT 43.470 155.430 43.810 156.260 ;
        RECT 47.160 154.690 47.510 155.940 ;
        RECT 48.990 155.430 49.330 156.260 ;
        RECT 51.360 155.995 51.605 156.600 ;
        RECT 51.825 156.270 52.335 156.805 ;
        RECT 51.085 155.825 52.315 155.995 ;
        RECT 51.085 155.015 51.425 155.825 ;
        RECT 51.595 155.260 52.345 155.450 ;
        RECT 40.050 154.255 45.395 154.690 ;
        RECT 45.570 154.255 50.915 154.690 ;
        RECT 51.085 154.605 51.600 155.015 ;
        RECT 51.835 154.255 52.005 155.015 ;
        RECT 52.175 154.595 52.345 155.260 ;
        RECT 52.515 155.275 52.705 156.635 ;
        RECT 52.875 156.465 53.150 156.635 ;
        RECT 52.875 156.295 53.155 156.465 ;
        RECT 52.875 155.475 53.150 156.295 ;
        RECT 53.340 156.270 53.870 156.635 ;
        RECT 54.295 156.405 54.625 156.805 ;
        RECT 53.695 156.235 53.870 156.270 ;
        RECT 53.355 155.275 53.525 156.075 ;
        RECT 52.515 155.105 53.525 155.275 ;
        RECT 53.695 156.065 54.625 156.235 ;
        RECT 54.795 156.065 55.050 156.635 ;
        RECT 53.695 154.935 53.865 156.065 ;
        RECT 54.455 155.895 54.625 156.065 ;
        RECT 52.740 154.765 53.865 154.935 ;
        RECT 54.035 155.565 54.230 155.895 ;
        RECT 54.455 155.565 54.710 155.895 ;
        RECT 54.035 154.595 54.205 155.565 ;
        RECT 54.880 155.395 55.050 156.065 ;
        RECT 55.225 156.055 56.435 156.805 ;
        RECT 56.695 156.255 56.865 156.635 ;
        RECT 57.045 156.425 57.375 156.805 ;
        RECT 56.695 156.085 57.360 156.255 ;
        RECT 57.555 156.130 57.815 156.635 ;
        RECT 52.175 154.425 54.205 154.595 ;
        RECT 54.375 154.255 54.545 155.395 ;
        RECT 54.715 154.425 55.050 155.395 ;
        RECT 55.225 155.345 55.745 155.885 ;
        RECT 55.915 155.515 56.435 156.055 ;
        RECT 56.625 155.535 56.955 155.905 ;
        RECT 57.190 155.830 57.360 156.085 ;
        RECT 57.190 155.500 57.475 155.830 ;
        RECT 57.190 155.355 57.360 155.500 ;
        RECT 55.225 154.255 56.435 155.345 ;
        RECT 56.695 155.185 57.360 155.355 ;
        RECT 57.645 155.330 57.815 156.130 ;
        RECT 57.985 156.055 59.195 156.805 ;
        RECT 56.695 154.425 56.865 155.185 ;
        RECT 57.045 154.255 57.375 155.015 ;
        RECT 57.545 154.425 57.815 155.330 ;
        RECT 57.985 155.345 58.505 155.885 ;
        RECT 58.675 155.515 59.195 156.055 ;
        RECT 59.365 156.035 62.875 156.805 ;
        RECT 63.045 156.080 63.335 156.805 ;
        RECT 63.505 156.035 66.095 156.805 ;
        RECT 59.365 155.345 61.055 155.865 ;
        RECT 61.225 155.515 62.875 156.035 ;
        RECT 57.985 154.255 59.195 155.345 ;
        RECT 59.365 154.255 62.875 155.345 ;
        RECT 63.045 154.255 63.335 155.420 ;
        RECT 63.505 155.345 64.715 155.865 ;
        RECT 64.885 155.515 66.095 156.035 ;
        RECT 66.270 155.965 66.530 156.805 ;
        RECT 66.705 156.060 66.960 156.635 ;
        RECT 67.130 156.425 67.460 156.805 ;
        RECT 67.675 156.255 67.845 156.635 ;
        RECT 67.130 156.085 67.845 156.255 ;
        RECT 68.195 156.255 68.365 156.635 ;
        RECT 68.580 156.425 68.910 156.805 ;
        RECT 68.195 156.085 68.910 156.255 ;
        RECT 63.505 154.255 66.095 155.345 ;
        RECT 66.270 154.255 66.530 155.405 ;
        RECT 66.705 155.330 66.875 156.060 ;
        RECT 67.130 155.895 67.300 156.085 ;
        RECT 67.045 155.565 67.300 155.895 ;
        RECT 67.130 155.355 67.300 155.565 ;
        RECT 67.580 155.535 67.935 155.905 ;
        RECT 68.105 155.535 68.460 155.905 ;
        RECT 68.740 155.895 68.910 156.085 ;
        RECT 69.080 156.060 69.335 156.635 ;
        RECT 68.740 155.565 68.995 155.895 ;
        RECT 68.740 155.355 68.910 155.565 ;
        RECT 66.705 154.425 66.960 155.330 ;
        RECT 67.130 155.185 67.845 155.355 ;
        RECT 67.130 154.255 67.460 155.015 ;
        RECT 67.675 154.425 67.845 155.185 ;
        RECT 68.195 155.185 68.910 155.355 ;
        RECT 69.165 155.330 69.335 156.060 ;
        RECT 69.510 155.965 69.770 156.805 ;
        RECT 70.035 156.255 70.205 156.635 ;
        RECT 70.420 156.425 70.750 156.805 ;
        RECT 70.035 156.085 70.750 156.255 ;
        RECT 69.945 155.535 70.300 155.905 ;
        RECT 70.580 155.895 70.750 156.085 ;
        RECT 70.920 156.060 71.175 156.635 ;
        RECT 70.580 155.565 70.835 155.895 ;
        RECT 68.195 154.425 68.365 155.185 ;
        RECT 68.580 154.255 68.910 155.015 ;
        RECT 69.080 154.425 69.335 155.330 ;
        RECT 69.510 154.255 69.770 155.405 ;
        RECT 70.580 155.355 70.750 155.565 ;
        RECT 70.035 155.185 70.750 155.355 ;
        RECT 71.005 155.330 71.175 156.060 ;
        RECT 71.350 155.965 71.610 156.805 ;
        RECT 71.790 155.965 72.050 156.805 ;
        RECT 72.225 156.060 72.480 156.635 ;
        RECT 72.650 156.425 72.980 156.805 ;
        RECT 73.195 156.255 73.365 156.635 ;
        RECT 72.650 156.085 73.365 156.255 ;
        RECT 70.035 154.425 70.205 155.185 ;
        RECT 70.420 154.255 70.750 155.015 ;
        RECT 70.920 154.425 71.175 155.330 ;
        RECT 71.350 154.255 71.610 155.405 ;
        RECT 71.790 154.255 72.050 155.405 ;
        RECT 72.225 155.330 72.395 156.060 ;
        RECT 72.650 155.895 72.820 156.085 ;
        RECT 73.625 156.055 74.835 156.805 ;
        RECT 72.565 155.565 72.820 155.895 ;
        RECT 72.650 155.355 72.820 155.565 ;
        RECT 73.100 155.535 73.455 155.905 ;
        RECT 72.225 154.425 72.480 155.330 ;
        RECT 72.650 155.185 73.365 155.355 ;
        RECT 72.650 154.255 72.980 155.015 ;
        RECT 73.195 154.425 73.365 155.185 ;
        RECT 73.625 155.345 74.145 155.885 ;
        RECT 74.315 155.515 74.835 156.055 ;
        RECT 75.005 156.035 78.515 156.805 ;
        RECT 75.005 155.345 76.695 155.865 ;
        RECT 76.865 155.515 78.515 156.035 ;
        RECT 78.685 156.005 79.025 156.635 ;
        RECT 79.195 156.005 79.445 156.805 ;
        RECT 79.635 156.155 79.965 156.635 ;
        RECT 80.135 156.345 80.360 156.805 ;
        RECT 80.530 156.155 80.860 156.635 ;
        RECT 78.685 155.395 78.860 156.005 ;
        RECT 79.635 155.985 80.860 156.155 ;
        RECT 81.490 156.025 81.990 156.635 ;
        RECT 79.030 155.645 79.725 155.815 ;
        RECT 79.555 155.395 79.725 155.645 ;
        RECT 79.900 155.615 80.320 155.815 ;
        RECT 80.490 155.615 80.820 155.815 ;
        RECT 80.990 155.615 81.320 155.815 ;
        RECT 81.490 155.395 81.660 156.025 ;
        RECT 83.100 155.995 83.345 156.600 ;
        RECT 83.565 156.270 84.075 156.805 ;
        RECT 82.825 155.825 84.055 155.995 ;
        RECT 81.845 155.565 82.195 155.815 ;
        RECT 73.625 154.255 74.835 155.345 ;
        RECT 75.005 154.255 78.515 155.345 ;
        RECT 78.685 154.425 79.025 155.395 ;
        RECT 79.195 154.255 79.365 155.395 ;
        RECT 79.555 155.225 81.990 155.395 ;
        RECT 79.635 154.255 79.885 155.055 ;
        RECT 80.530 154.425 80.860 155.225 ;
        RECT 81.160 154.255 81.490 155.055 ;
        RECT 81.660 154.425 81.990 155.225 ;
        RECT 82.825 155.015 83.165 155.825 ;
        RECT 83.335 155.260 84.085 155.450 ;
        RECT 82.825 154.605 83.340 155.015 ;
        RECT 83.575 154.255 83.745 155.015 ;
        RECT 83.915 154.595 84.085 155.260 ;
        RECT 84.255 155.275 84.445 156.635 ;
        RECT 84.615 155.785 84.890 156.635 ;
        RECT 85.080 156.270 85.610 156.635 ;
        RECT 86.035 156.405 86.365 156.805 ;
        RECT 85.435 156.235 85.610 156.270 ;
        RECT 84.615 155.615 84.895 155.785 ;
        RECT 84.615 155.475 84.890 155.615 ;
        RECT 85.095 155.275 85.265 156.075 ;
        RECT 84.255 155.105 85.265 155.275 ;
        RECT 85.435 156.065 86.365 156.235 ;
        RECT 86.535 156.065 86.790 156.635 ;
        RECT 85.435 154.935 85.605 156.065 ;
        RECT 86.195 155.895 86.365 156.065 ;
        RECT 84.480 154.765 85.605 154.935 ;
        RECT 85.775 155.565 85.970 155.895 ;
        RECT 86.195 155.565 86.450 155.895 ;
        RECT 85.775 154.595 85.945 155.565 ;
        RECT 86.620 155.395 86.790 156.065 ;
        RECT 86.965 156.035 88.635 156.805 ;
        RECT 88.805 156.080 89.095 156.805 ;
        RECT 89.725 156.035 92.315 156.805 ;
        RECT 92.490 156.260 97.835 156.805 ;
        RECT 83.915 154.425 85.945 154.595 ;
        RECT 86.115 154.255 86.285 155.395 ;
        RECT 86.455 154.425 86.790 155.395 ;
        RECT 86.965 155.345 87.715 155.865 ;
        RECT 87.885 155.515 88.635 156.035 ;
        RECT 86.965 154.255 88.635 155.345 ;
        RECT 88.805 154.255 89.095 155.420 ;
        RECT 89.725 155.345 90.935 155.865 ;
        RECT 91.105 155.515 92.315 156.035 ;
        RECT 89.725 154.255 92.315 155.345 ;
        RECT 94.080 154.690 94.430 155.940 ;
        RECT 95.910 155.430 96.250 156.260 ;
        RECT 98.005 156.005 98.345 156.635 ;
        RECT 98.515 156.005 98.765 156.805 ;
        RECT 98.955 156.155 99.285 156.635 ;
        RECT 99.455 156.345 99.680 156.805 ;
        RECT 99.850 156.155 100.180 156.635 ;
        RECT 98.005 155.395 98.180 156.005 ;
        RECT 98.955 155.985 100.180 156.155 ;
        RECT 100.810 156.025 101.310 156.635 ;
        RECT 101.685 156.035 103.355 156.805 ;
        RECT 98.350 155.645 99.045 155.815 ;
        RECT 98.875 155.395 99.045 155.645 ;
        RECT 99.220 155.615 99.640 155.815 ;
        RECT 99.810 155.615 100.140 155.815 ;
        RECT 100.310 155.615 100.640 155.815 ;
        RECT 100.810 155.395 100.980 156.025 ;
        RECT 101.165 155.565 101.515 155.815 ;
        RECT 92.490 154.255 97.835 154.690 ;
        RECT 98.005 154.425 98.345 155.395 ;
        RECT 98.515 154.255 98.685 155.395 ;
        RECT 98.875 155.225 101.310 155.395 ;
        RECT 98.955 154.255 99.205 155.055 ;
        RECT 99.850 154.425 100.180 155.225 ;
        RECT 100.480 154.255 100.810 155.055 ;
        RECT 100.980 154.425 101.310 155.225 ;
        RECT 101.685 155.345 102.435 155.865 ;
        RECT 102.605 155.515 103.355 156.035 ;
        RECT 103.525 156.005 103.865 156.635 ;
        RECT 104.035 156.005 104.285 156.805 ;
        RECT 104.475 156.155 104.805 156.635 ;
        RECT 104.975 156.345 105.200 156.805 ;
        RECT 105.370 156.155 105.700 156.635 ;
        RECT 103.525 155.395 103.700 156.005 ;
        RECT 104.475 155.985 105.700 156.155 ;
        RECT 106.330 156.025 106.830 156.635 ;
        RECT 103.870 155.645 104.565 155.815 ;
        RECT 104.395 155.395 104.565 155.645 ;
        RECT 104.740 155.615 105.160 155.815 ;
        RECT 105.330 155.615 105.660 155.815 ;
        RECT 105.830 155.615 106.160 155.815 ;
        RECT 106.330 155.395 106.500 156.025 ;
        RECT 107.205 156.005 107.545 156.635 ;
        RECT 107.715 156.005 107.965 156.805 ;
        RECT 108.155 156.155 108.485 156.635 ;
        RECT 108.655 156.345 108.880 156.805 ;
        RECT 109.050 156.155 109.380 156.635 ;
        RECT 106.685 155.565 107.035 155.815 ;
        RECT 107.205 155.395 107.380 156.005 ;
        RECT 108.155 155.985 109.380 156.155 ;
        RECT 110.010 156.025 110.510 156.635 ;
        RECT 107.550 155.645 108.245 155.815 ;
        RECT 108.075 155.395 108.245 155.645 ;
        RECT 108.420 155.615 108.840 155.815 ;
        RECT 109.010 155.615 109.340 155.815 ;
        RECT 109.510 155.615 109.840 155.815 ;
        RECT 110.010 155.395 110.180 156.025 ;
        RECT 110.885 156.005 111.225 156.635 ;
        RECT 111.395 156.005 111.645 156.805 ;
        RECT 111.835 156.155 112.165 156.635 ;
        RECT 112.335 156.345 112.560 156.805 ;
        RECT 112.730 156.155 113.060 156.635 ;
        RECT 110.365 155.565 110.715 155.815 ;
        RECT 110.885 155.395 111.060 156.005 ;
        RECT 111.835 155.985 113.060 156.155 ;
        RECT 113.690 156.025 114.190 156.635 ;
        RECT 114.565 156.080 114.855 156.805 ;
        RECT 111.230 155.645 111.925 155.815 ;
        RECT 111.755 155.395 111.925 155.645 ;
        RECT 112.100 155.615 112.520 155.815 ;
        RECT 112.690 155.615 113.020 155.815 ;
        RECT 113.190 155.615 113.520 155.815 ;
        RECT 113.690 155.395 113.860 156.025 ;
        RECT 115.065 155.985 115.295 156.805 ;
        RECT 115.465 156.005 115.795 156.635 ;
        RECT 114.045 155.565 114.395 155.815 ;
        RECT 115.045 155.565 115.375 155.815 ;
        RECT 101.685 154.255 103.355 155.345 ;
        RECT 103.525 154.425 103.865 155.395 ;
        RECT 104.035 154.255 104.205 155.395 ;
        RECT 104.395 155.225 106.830 155.395 ;
        RECT 104.475 154.255 104.725 155.055 ;
        RECT 105.370 154.425 105.700 155.225 ;
        RECT 106.000 154.255 106.330 155.055 ;
        RECT 106.500 154.425 106.830 155.225 ;
        RECT 107.205 154.425 107.545 155.395 ;
        RECT 107.715 154.255 107.885 155.395 ;
        RECT 108.075 155.225 110.510 155.395 ;
        RECT 108.155 154.255 108.405 155.055 ;
        RECT 109.050 154.425 109.380 155.225 ;
        RECT 109.680 154.255 110.010 155.055 ;
        RECT 110.180 154.425 110.510 155.225 ;
        RECT 110.885 154.425 111.225 155.395 ;
        RECT 111.395 154.255 111.565 155.395 ;
        RECT 111.755 155.225 114.190 155.395 ;
        RECT 111.835 154.255 112.085 155.055 ;
        RECT 112.730 154.425 113.060 155.225 ;
        RECT 113.360 154.255 113.690 155.055 ;
        RECT 113.860 154.425 114.190 155.225 ;
        RECT 114.565 154.255 114.855 155.420 ;
        RECT 115.545 155.405 115.795 156.005 ;
        RECT 115.965 155.985 116.175 156.805 ;
        RECT 116.410 156.095 116.665 156.625 ;
        RECT 116.835 156.345 117.140 156.805 ;
        RECT 117.385 156.425 118.455 156.595 ;
        RECT 115.065 154.255 115.295 155.395 ;
        RECT 115.465 154.425 115.795 155.405 ;
        RECT 116.410 155.445 116.620 156.095 ;
        RECT 117.385 156.070 117.705 156.425 ;
        RECT 117.380 155.895 117.705 156.070 ;
        RECT 116.790 155.595 117.705 155.895 ;
        RECT 117.875 155.855 118.115 156.255 ;
        RECT 118.285 156.195 118.455 156.425 ;
        RECT 118.625 156.365 118.815 156.805 ;
        RECT 118.985 156.355 119.935 156.635 ;
        RECT 120.155 156.445 120.505 156.615 ;
        RECT 118.285 156.025 118.815 156.195 ;
        RECT 116.790 155.565 117.530 155.595 ;
        RECT 115.965 154.255 116.175 155.395 ;
        RECT 116.410 154.565 116.665 155.445 ;
        RECT 116.835 154.255 117.140 155.395 ;
        RECT 117.360 154.975 117.530 155.565 ;
        RECT 117.875 155.485 118.415 155.855 ;
        RECT 118.595 155.745 118.815 156.025 ;
        RECT 118.985 155.575 119.155 156.355 ;
        RECT 118.750 155.405 119.155 155.575 ;
        RECT 119.325 155.565 119.675 156.185 ;
        RECT 118.750 155.315 118.920 155.405 ;
        RECT 119.845 155.395 120.055 156.185 ;
        RECT 117.700 155.145 118.920 155.315 ;
        RECT 119.380 155.235 120.055 155.395 ;
        RECT 117.360 154.805 118.160 154.975 ;
        RECT 117.480 154.255 117.810 154.635 ;
        RECT 117.990 154.515 118.160 154.805 ;
        RECT 118.750 154.765 118.920 155.145 ;
        RECT 119.090 155.225 120.055 155.235 ;
        RECT 120.245 156.055 120.505 156.445 ;
        RECT 120.715 156.345 121.045 156.805 ;
        RECT 121.920 156.415 122.775 156.585 ;
        RECT 122.980 156.415 123.475 156.585 ;
        RECT 123.645 156.445 123.975 156.805 ;
        RECT 120.245 155.365 120.415 156.055 ;
        RECT 120.585 155.705 120.755 155.885 ;
        RECT 120.925 155.875 121.715 156.125 ;
        RECT 121.920 155.705 122.090 156.415 ;
        RECT 122.260 155.905 122.615 156.125 ;
        RECT 120.585 155.535 122.275 155.705 ;
        RECT 119.090 154.935 119.550 155.225 ;
        RECT 120.245 155.195 121.745 155.365 ;
        RECT 120.245 155.055 120.415 155.195 ;
        RECT 119.855 154.885 120.415 155.055 ;
        RECT 118.330 154.255 118.580 154.715 ;
        RECT 118.750 154.425 119.620 154.765 ;
        RECT 119.855 154.425 120.025 154.885 ;
        RECT 120.860 154.855 121.935 155.025 ;
        RECT 120.195 154.255 120.565 154.715 ;
        RECT 120.860 154.515 121.030 154.855 ;
        RECT 121.200 154.255 121.530 154.685 ;
        RECT 121.765 154.515 121.935 154.855 ;
        RECT 122.105 154.755 122.275 155.535 ;
        RECT 122.445 155.315 122.615 155.905 ;
        RECT 122.785 155.505 123.135 156.125 ;
        RECT 122.445 154.925 122.910 155.315 ;
        RECT 123.305 155.055 123.475 156.415 ;
        RECT 123.645 155.225 124.105 156.275 ;
        RECT 123.080 154.885 123.475 155.055 ;
        RECT 123.080 154.755 123.250 154.885 ;
        RECT 122.105 154.425 122.785 154.755 ;
        RECT 123.000 154.425 123.250 154.755 ;
        RECT 123.420 154.255 123.670 154.715 ;
        RECT 123.840 154.440 124.165 155.225 ;
        RECT 124.335 154.425 124.505 156.545 ;
        RECT 124.675 156.425 125.005 156.805 ;
        RECT 125.175 156.255 125.430 156.545 ;
        RECT 124.680 156.085 125.430 156.255 ;
        RECT 124.680 155.095 124.910 156.085 ;
        RECT 126.525 156.055 127.735 156.805 ;
        RECT 125.080 155.265 125.430 155.915 ;
        RECT 126.525 155.345 127.045 155.885 ;
        RECT 127.215 155.515 127.735 156.055 ;
        RECT 124.680 154.925 125.430 155.095 ;
        RECT 124.675 154.255 125.005 154.755 ;
        RECT 125.175 154.425 125.430 154.925 ;
        RECT 126.525 154.255 127.735 155.345 ;
        RECT 14.660 154.085 127.820 154.255 ;
        RECT 14.745 152.995 15.955 154.085 ;
        RECT 14.745 152.285 15.265 152.825 ;
        RECT 15.435 152.455 15.955 152.995 ;
        RECT 16.585 152.995 20.095 154.085 ;
        RECT 20.265 153.325 20.780 153.735 ;
        RECT 21.015 153.325 21.185 154.085 ;
        RECT 21.355 153.745 23.385 153.915 ;
        RECT 16.585 152.475 18.275 152.995 ;
        RECT 18.445 152.305 20.095 152.825 ;
        RECT 20.265 152.515 20.605 153.325 ;
        RECT 21.355 153.080 21.525 153.745 ;
        RECT 21.920 153.405 23.045 153.575 ;
        RECT 20.775 152.890 21.525 153.080 ;
        RECT 21.695 153.065 22.705 153.235 ;
        RECT 20.265 152.345 21.495 152.515 ;
        RECT 14.745 151.535 15.955 152.285 ;
        RECT 16.585 151.535 20.095 152.305 ;
        RECT 20.540 151.740 20.785 152.345 ;
        RECT 21.005 151.535 21.515 152.070 ;
        RECT 21.695 151.705 21.885 153.065 ;
        RECT 22.055 152.385 22.330 152.865 ;
        RECT 22.055 152.215 22.335 152.385 ;
        RECT 22.535 152.265 22.705 153.065 ;
        RECT 22.875 152.275 23.045 153.405 ;
        RECT 23.215 152.775 23.385 153.745 ;
        RECT 23.555 152.945 23.725 154.085 ;
        RECT 23.895 152.945 24.230 153.915 ;
        RECT 23.215 152.445 23.410 152.775 ;
        RECT 23.635 152.445 23.890 152.775 ;
        RECT 23.635 152.275 23.805 152.445 ;
        RECT 24.060 152.275 24.230 152.945 ;
        RECT 24.405 152.920 24.695 154.085 ;
        RECT 24.865 152.995 26.535 154.085 ;
        RECT 26.705 153.325 27.220 153.735 ;
        RECT 27.455 153.325 27.625 154.085 ;
        RECT 27.795 153.745 29.825 153.915 ;
        RECT 24.865 152.475 25.615 152.995 ;
        RECT 25.785 152.305 26.535 152.825 ;
        RECT 26.705 152.515 27.045 153.325 ;
        RECT 27.795 153.080 27.965 153.745 ;
        RECT 28.360 153.405 29.485 153.575 ;
        RECT 27.215 152.890 27.965 153.080 ;
        RECT 28.135 153.065 29.145 153.235 ;
        RECT 26.705 152.345 27.935 152.515 ;
        RECT 22.055 151.705 22.330 152.215 ;
        RECT 22.875 152.105 23.805 152.275 ;
        RECT 22.875 152.070 23.050 152.105 ;
        RECT 22.520 151.705 23.050 152.070 ;
        RECT 23.475 151.535 23.805 151.935 ;
        RECT 23.975 151.705 24.230 152.275 ;
        RECT 24.405 151.535 24.695 152.260 ;
        RECT 24.865 151.535 26.535 152.305 ;
        RECT 26.980 151.740 27.225 152.345 ;
        RECT 27.445 151.535 27.955 152.070 ;
        RECT 28.135 151.705 28.325 153.065 ;
        RECT 28.495 152.725 28.770 152.865 ;
        RECT 28.495 152.555 28.775 152.725 ;
        RECT 28.495 151.705 28.770 152.555 ;
        RECT 28.975 152.265 29.145 153.065 ;
        RECT 29.315 152.275 29.485 153.405 ;
        RECT 29.655 152.775 29.825 153.745 ;
        RECT 29.995 152.945 30.165 154.085 ;
        RECT 30.335 152.945 30.670 153.915 ;
        RECT 31.510 153.115 31.840 153.915 ;
        RECT 32.010 153.285 32.340 154.085 ;
        RECT 32.640 153.115 32.970 153.915 ;
        RECT 33.615 153.285 33.865 154.085 ;
        RECT 31.510 152.945 33.945 153.115 ;
        RECT 34.135 152.945 34.305 154.085 ;
        RECT 34.475 152.945 34.815 153.915 ;
        RECT 29.655 152.445 29.850 152.775 ;
        RECT 30.075 152.445 30.330 152.775 ;
        RECT 30.075 152.275 30.245 152.445 ;
        RECT 30.500 152.275 30.670 152.945 ;
        RECT 31.305 152.525 31.655 152.775 ;
        RECT 31.840 152.315 32.010 152.945 ;
        RECT 32.180 152.525 32.510 152.725 ;
        RECT 32.680 152.525 33.010 152.725 ;
        RECT 33.180 152.525 33.600 152.725 ;
        RECT 33.775 152.695 33.945 152.945 ;
        RECT 33.775 152.525 34.470 152.695 ;
        RECT 29.315 152.105 30.245 152.275 ;
        RECT 29.315 152.070 29.490 152.105 ;
        RECT 28.960 151.705 29.490 152.070 ;
        RECT 29.915 151.535 30.245 151.935 ;
        RECT 30.415 151.705 30.670 152.275 ;
        RECT 31.510 151.705 32.010 152.315 ;
        RECT 32.640 152.185 33.865 152.355 ;
        RECT 34.640 152.335 34.815 152.945 ;
        RECT 32.640 151.705 32.970 152.185 ;
        RECT 33.140 151.535 33.365 151.995 ;
        RECT 33.535 151.705 33.865 152.185 ;
        RECT 34.055 151.535 34.305 152.335 ;
        RECT 34.475 151.705 34.815 152.335 ;
        RECT 34.985 152.945 35.325 153.915 ;
        RECT 35.495 152.945 35.665 154.085 ;
        RECT 35.935 153.285 36.185 154.085 ;
        RECT 36.830 153.115 37.160 153.915 ;
        RECT 37.460 153.285 37.790 154.085 ;
        RECT 37.960 153.115 38.290 153.915 ;
        RECT 35.855 152.945 38.290 153.115 ;
        RECT 39.125 152.995 42.635 154.085 ;
        RECT 43.010 153.115 43.340 153.915 ;
        RECT 43.510 153.285 43.840 154.085 ;
        RECT 44.140 153.115 44.470 153.915 ;
        RECT 45.115 153.285 45.365 154.085 ;
        RECT 34.985 152.335 35.160 152.945 ;
        RECT 35.855 152.695 36.025 152.945 ;
        RECT 35.330 152.525 36.025 152.695 ;
        RECT 36.200 152.525 36.620 152.725 ;
        RECT 36.790 152.525 37.120 152.725 ;
        RECT 37.290 152.525 37.620 152.725 ;
        RECT 34.985 151.705 35.325 152.335 ;
        RECT 35.495 151.535 35.745 152.335 ;
        RECT 35.935 152.185 37.160 152.355 ;
        RECT 35.935 151.705 36.265 152.185 ;
        RECT 36.435 151.535 36.660 151.995 ;
        RECT 36.830 151.705 37.160 152.185 ;
        RECT 37.790 152.315 37.960 152.945 ;
        RECT 38.145 152.525 38.495 152.775 ;
        RECT 39.125 152.475 40.815 152.995 ;
        RECT 43.010 152.945 45.445 153.115 ;
        RECT 45.635 152.945 45.805 154.085 ;
        RECT 45.975 152.945 46.315 153.915 ;
        RECT 46.690 153.115 47.020 153.915 ;
        RECT 47.190 153.285 47.520 154.085 ;
        RECT 47.820 153.115 48.150 153.915 ;
        RECT 48.795 153.285 49.045 154.085 ;
        RECT 46.690 152.945 49.125 153.115 ;
        RECT 49.315 152.945 49.485 154.085 ;
        RECT 49.655 152.945 49.995 153.915 ;
        RECT 37.790 151.705 38.290 152.315 ;
        RECT 40.985 152.305 42.635 152.825 ;
        RECT 42.805 152.525 43.155 152.775 ;
        RECT 43.340 152.315 43.510 152.945 ;
        RECT 43.680 152.525 44.010 152.725 ;
        RECT 44.180 152.525 44.510 152.725 ;
        RECT 44.680 152.525 45.100 152.725 ;
        RECT 45.275 152.695 45.445 152.945 ;
        RECT 45.275 152.525 45.970 152.695 ;
        RECT 39.125 151.535 42.635 152.305 ;
        RECT 43.010 151.705 43.510 152.315 ;
        RECT 44.140 152.185 45.365 152.355 ;
        RECT 46.140 152.335 46.315 152.945 ;
        RECT 46.485 152.525 46.835 152.775 ;
        RECT 44.140 151.705 44.470 152.185 ;
        RECT 44.640 151.535 44.865 151.995 ;
        RECT 45.035 151.705 45.365 152.185 ;
        RECT 45.555 151.535 45.805 152.335 ;
        RECT 45.975 151.705 46.315 152.335 ;
        RECT 47.020 152.315 47.190 152.945 ;
        RECT 47.360 152.525 47.690 152.725 ;
        RECT 47.860 152.525 48.190 152.725 ;
        RECT 48.360 152.525 48.780 152.725 ;
        RECT 48.955 152.695 49.125 152.945 ;
        RECT 48.955 152.525 49.650 152.695 ;
        RECT 46.690 151.705 47.190 152.315 ;
        RECT 47.820 152.185 49.045 152.355 ;
        RECT 49.820 152.335 49.995 152.945 ;
        RECT 50.165 152.920 50.455 154.085 ;
        RECT 50.625 152.945 50.965 153.915 ;
        RECT 51.135 152.945 51.305 154.085 ;
        RECT 51.575 153.285 51.825 154.085 ;
        RECT 52.470 153.115 52.800 153.915 ;
        RECT 53.100 153.285 53.430 154.085 ;
        RECT 53.600 153.115 53.930 153.915 ;
        RECT 51.495 152.945 53.930 153.115 ;
        RECT 54.765 152.995 56.435 154.085 ;
        RECT 56.610 153.650 61.955 154.085 ;
        RECT 47.820 151.705 48.150 152.185 ;
        RECT 48.320 151.535 48.545 151.995 ;
        RECT 48.715 151.705 49.045 152.185 ;
        RECT 49.235 151.535 49.485 152.335 ;
        RECT 49.655 151.705 49.995 152.335 ;
        RECT 50.625 152.895 50.855 152.945 ;
        RECT 50.625 152.335 50.800 152.895 ;
        RECT 51.495 152.695 51.665 152.945 ;
        RECT 50.970 152.525 51.665 152.695 ;
        RECT 51.840 152.525 52.260 152.725 ;
        RECT 52.430 152.525 52.760 152.725 ;
        RECT 52.930 152.525 53.260 152.725 ;
        RECT 50.165 151.535 50.455 152.260 ;
        RECT 50.625 151.705 50.965 152.335 ;
        RECT 51.135 151.535 51.385 152.335 ;
        RECT 51.575 152.185 52.800 152.355 ;
        RECT 51.575 151.705 51.905 152.185 ;
        RECT 52.075 151.535 52.300 151.995 ;
        RECT 52.470 151.705 52.800 152.185 ;
        RECT 53.430 152.315 53.600 152.945 ;
        RECT 53.785 152.525 54.135 152.775 ;
        RECT 54.765 152.475 55.515 152.995 ;
        RECT 53.430 151.705 53.930 152.315 ;
        RECT 55.685 152.305 56.435 152.825 ;
        RECT 58.200 152.400 58.550 153.650 ;
        RECT 62.165 152.945 62.395 154.085 ;
        RECT 62.565 152.935 62.895 153.915 ;
        RECT 63.065 152.945 63.275 154.085 ;
        RECT 63.510 152.935 63.770 154.085 ;
        RECT 63.945 153.010 64.200 153.915 ;
        RECT 64.370 153.325 64.700 154.085 ;
        RECT 64.915 153.155 65.085 153.915 ;
        RECT 54.765 151.535 56.435 152.305 ;
        RECT 60.030 152.080 60.370 152.910 ;
        RECT 62.145 152.525 62.475 152.775 ;
        RECT 56.610 151.535 61.955 152.080 ;
        RECT 62.165 151.535 62.395 152.355 ;
        RECT 62.645 152.335 62.895 152.935 ;
        RECT 62.565 151.705 62.895 152.335 ;
        RECT 63.065 151.535 63.275 152.355 ;
        RECT 63.510 151.535 63.770 152.375 ;
        RECT 63.945 152.280 64.115 153.010 ;
        RECT 64.370 152.985 65.085 153.155 ;
        RECT 64.370 152.775 64.540 152.985 ;
        RECT 65.345 152.945 65.685 153.915 ;
        RECT 65.855 152.945 66.025 154.085 ;
        RECT 66.295 153.285 66.545 154.085 ;
        RECT 67.190 153.115 67.520 153.915 ;
        RECT 67.820 153.285 68.150 154.085 ;
        RECT 68.320 153.115 68.650 153.915 ;
        RECT 70.000 153.215 70.285 154.085 ;
        RECT 70.455 153.455 70.715 153.915 ;
        RECT 70.890 153.625 71.145 154.085 ;
        RECT 71.315 153.455 71.575 153.915 ;
        RECT 70.455 153.285 71.575 153.455 ;
        RECT 71.745 153.285 72.055 154.085 ;
        RECT 66.215 152.945 68.650 153.115 ;
        RECT 70.455 153.035 70.715 153.285 ;
        RECT 72.225 153.115 72.535 153.915 ;
        RECT 64.285 152.445 64.540 152.775 ;
        RECT 63.945 151.705 64.200 152.280 ;
        RECT 64.370 152.255 64.540 152.445 ;
        RECT 64.820 152.435 65.175 152.805 ;
        RECT 65.345 152.335 65.520 152.945 ;
        RECT 66.215 152.695 66.385 152.945 ;
        RECT 65.690 152.525 66.385 152.695 ;
        RECT 66.560 152.525 66.980 152.725 ;
        RECT 67.150 152.525 67.480 152.725 ;
        RECT 67.650 152.525 67.980 152.725 ;
        RECT 64.370 152.085 65.085 152.255 ;
        RECT 64.370 151.535 64.700 151.915 ;
        RECT 64.915 151.705 65.085 152.085 ;
        RECT 65.345 151.705 65.685 152.335 ;
        RECT 65.855 151.535 66.105 152.335 ;
        RECT 66.295 152.185 67.520 152.355 ;
        RECT 66.295 151.705 66.625 152.185 ;
        RECT 66.795 151.535 67.020 151.995 ;
        RECT 67.190 151.705 67.520 152.185 ;
        RECT 68.150 152.315 68.320 152.945 ;
        RECT 69.960 152.865 70.715 153.035 ;
        RECT 71.505 152.945 72.535 153.115 ;
        RECT 72.715 153.025 73.045 154.085 ;
        RECT 68.505 152.525 68.855 152.775 ;
        RECT 69.960 152.355 70.365 152.865 ;
        RECT 71.505 152.695 71.675 152.945 ;
        RECT 70.535 152.525 71.675 152.695 ;
        RECT 68.150 151.705 68.650 152.315 ;
        RECT 69.960 152.185 71.610 152.355 ;
        RECT 71.845 152.205 72.195 152.775 ;
        RECT 70.005 151.535 70.285 152.015 ;
        RECT 70.455 151.795 70.715 152.185 ;
        RECT 70.890 151.535 71.145 152.015 ;
        RECT 71.315 151.795 71.610 152.185 ;
        RECT 72.365 152.035 72.535 152.945 ;
        RECT 73.225 152.775 73.395 153.745 ;
        RECT 73.565 153.495 73.895 153.895 ;
        RECT 74.065 153.725 74.395 154.085 ;
        RECT 74.595 153.495 75.295 153.915 ;
        RECT 73.565 153.265 75.295 153.495 ;
        RECT 73.565 153.045 73.895 153.265 ;
        RECT 74.090 152.775 74.415 153.065 ;
        RECT 72.705 152.445 73.015 152.775 ;
        RECT 73.225 152.445 73.600 152.775 ;
        RECT 73.920 152.445 74.415 152.775 ;
        RECT 74.590 152.525 74.920 153.065 ;
        RECT 75.090 152.295 75.295 153.265 ;
        RECT 75.925 152.920 76.215 154.085 ;
        RECT 76.385 152.995 77.595 154.085 ;
        RECT 76.385 152.455 76.905 152.995 ;
        RECT 77.765 152.945 78.105 153.915 ;
        RECT 78.275 152.945 78.445 154.085 ;
        RECT 78.715 153.285 78.965 154.085 ;
        RECT 79.610 153.115 79.940 153.915 ;
        RECT 80.240 153.285 80.570 154.085 ;
        RECT 80.740 153.115 81.070 153.915 ;
        RECT 78.635 152.945 81.070 153.115 ;
        RECT 81.445 152.945 81.785 153.915 ;
        RECT 81.955 152.945 82.125 154.085 ;
        RECT 82.395 153.285 82.645 154.085 ;
        RECT 83.290 153.115 83.620 153.915 ;
        RECT 83.920 153.285 84.250 154.085 ;
        RECT 84.420 153.115 84.750 153.915 ;
        RECT 82.315 152.945 84.750 153.115 ;
        RECT 86.045 152.995 89.555 154.085 ;
        RECT 89.730 153.650 95.075 154.085 ;
        RECT 71.790 151.535 72.065 152.015 ;
        RECT 72.235 151.705 72.535 152.035 ;
        RECT 72.715 152.065 74.075 152.275 ;
        RECT 72.715 151.705 73.045 152.065 ;
        RECT 73.215 151.535 73.545 151.895 ;
        RECT 73.745 151.705 74.075 152.065 ;
        RECT 74.585 151.705 75.295 152.295 ;
        RECT 77.075 152.285 77.595 152.825 ;
        RECT 75.925 151.535 76.215 152.260 ;
        RECT 76.385 151.535 77.595 152.285 ;
        RECT 77.765 152.335 77.940 152.945 ;
        RECT 78.635 152.695 78.805 152.945 ;
        RECT 78.110 152.525 78.805 152.695 ;
        RECT 78.980 152.525 79.400 152.725 ;
        RECT 79.570 152.525 79.900 152.725 ;
        RECT 80.070 152.525 80.400 152.725 ;
        RECT 77.765 151.705 78.105 152.335 ;
        RECT 78.275 151.535 78.525 152.335 ;
        RECT 78.715 152.185 79.940 152.355 ;
        RECT 78.715 151.705 79.045 152.185 ;
        RECT 79.215 151.535 79.440 151.995 ;
        RECT 79.610 151.705 79.940 152.185 ;
        RECT 80.570 152.315 80.740 152.945 ;
        RECT 80.925 152.525 81.275 152.775 ;
        RECT 81.445 152.335 81.620 152.945 ;
        RECT 82.315 152.695 82.485 152.945 ;
        RECT 81.790 152.525 82.485 152.695 ;
        RECT 82.660 152.525 83.080 152.725 ;
        RECT 83.250 152.525 83.580 152.725 ;
        RECT 83.750 152.525 84.080 152.725 ;
        RECT 80.570 151.705 81.070 152.315 ;
        RECT 81.445 151.705 81.785 152.335 ;
        RECT 81.955 151.535 82.205 152.335 ;
        RECT 82.395 152.185 83.620 152.355 ;
        RECT 82.395 151.705 82.725 152.185 ;
        RECT 82.895 151.535 83.120 151.995 ;
        RECT 83.290 151.705 83.620 152.185 ;
        RECT 84.250 152.315 84.420 152.945 ;
        RECT 84.605 152.525 84.955 152.775 ;
        RECT 86.045 152.475 87.735 152.995 ;
        RECT 84.250 151.705 84.750 152.315 ;
        RECT 87.905 152.305 89.555 152.825 ;
        RECT 91.320 152.400 91.670 153.650 ;
        RECT 95.305 152.945 95.515 154.085 ;
        RECT 95.685 152.935 96.015 153.915 ;
        RECT 96.185 152.945 96.415 154.085 ;
        RECT 97.635 153.155 97.805 153.915 ;
        RECT 97.985 153.325 98.315 154.085 ;
        RECT 97.635 152.985 98.300 153.155 ;
        RECT 98.485 153.010 98.755 153.915 ;
        RECT 86.045 151.535 89.555 152.305 ;
        RECT 93.150 152.080 93.490 152.910 ;
        RECT 89.730 151.535 95.075 152.080 ;
        RECT 95.305 151.535 95.515 152.355 ;
        RECT 95.685 152.335 95.935 152.935 ;
        RECT 98.130 152.840 98.300 152.985 ;
        RECT 96.105 152.525 96.435 152.775 ;
        RECT 97.565 152.435 97.895 152.805 ;
        RECT 98.130 152.510 98.415 152.840 ;
        RECT 95.685 151.705 96.015 152.335 ;
        RECT 96.185 151.535 96.415 152.355 ;
        RECT 98.130 152.255 98.300 152.510 ;
        RECT 97.635 152.085 98.300 152.255 ;
        RECT 98.585 152.210 98.755 153.010 ;
        RECT 98.925 152.995 101.515 154.085 ;
        RECT 98.925 152.475 100.135 152.995 ;
        RECT 101.685 152.920 101.975 154.085 ;
        RECT 102.150 153.650 107.495 154.085 ;
        RECT 100.305 152.305 101.515 152.825 ;
        RECT 103.740 152.400 104.090 153.650 ;
        RECT 107.665 152.945 108.005 153.915 ;
        RECT 108.175 152.945 108.345 154.085 ;
        RECT 108.615 153.285 108.865 154.085 ;
        RECT 109.510 153.115 109.840 153.915 ;
        RECT 110.140 153.285 110.470 154.085 ;
        RECT 110.640 153.115 110.970 153.915 ;
        RECT 108.535 152.945 110.970 153.115 ;
        RECT 111.345 152.995 114.855 154.085 ;
        RECT 115.025 153.325 115.540 153.735 ;
        RECT 115.775 153.325 115.945 154.085 ;
        RECT 116.115 153.745 118.145 153.915 ;
        RECT 97.635 151.705 97.805 152.085 ;
        RECT 97.985 151.535 98.315 151.915 ;
        RECT 98.495 151.705 98.755 152.210 ;
        RECT 98.925 151.535 101.515 152.305 ;
        RECT 101.685 151.535 101.975 152.260 ;
        RECT 105.570 152.080 105.910 152.910 ;
        RECT 107.665 152.335 107.840 152.945 ;
        RECT 108.535 152.695 108.705 152.945 ;
        RECT 108.010 152.525 108.705 152.695 ;
        RECT 108.880 152.525 109.300 152.725 ;
        RECT 109.470 152.525 109.800 152.725 ;
        RECT 109.970 152.525 110.300 152.725 ;
        RECT 102.150 151.535 107.495 152.080 ;
        RECT 107.665 151.705 108.005 152.335 ;
        RECT 108.175 151.535 108.425 152.335 ;
        RECT 108.615 152.185 109.840 152.355 ;
        RECT 108.615 151.705 108.945 152.185 ;
        RECT 109.115 151.535 109.340 151.995 ;
        RECT 109.510 151.705 109.840 152.185 ;
        RECT 110.470 152.315 110.640 152.945 ;
        RECT 110.825 152.525 111.175 152.775 ;
        RECT 111.345 152.475 113.035 152.995 ;
        RECT 110.470 151.705 110.970 152.315 ;
        RECT 113.205 152.305 114.855 152.825 ;
        RECT 115.025 152.515 115.365 153.325 ;
        RECT 116.115 153.080 116.285 153.745 ;
        RECT 116.680 153.405 117.805 153.575 ;
        RECT 115.535 152.890 116.285 153.080 ;
        RECT 116.455 153.065 117.465 153.235 ;
        RECT 115.025 152.345 116.255 152.515 ;
        RECT 111.345 151.535 114.855 152.305 ;
        RECT 115.300 151.740 115.545 152.345 ;
        RECT 115.765 151.535 116.275 152.070 ;
        RECT 116.455 151.705 116.645 153.065 ;
        RECT 116.815 152.045 117.090 152.865 ;
        RECT 117.295 152.265 117.465 153.065 ;
        RECT 117.635 152.275 117.805 153.405 ;
        RECT 117.975 152.775 118.145 153.745 ;
        RECT 118.315 152.945 118.485 154.085 ;
        RECT 118.655 152.945 118.990 153.915 ;
        RECT 119.665 152.945 119.895 154.085 ;
        RECT 117.975 152.445 118.170 152.775 ;
        RECT 118.395 152.445 118.650 152.775 ;
        RECT 118.395 152.275 118.565 152.445 ;
        RECT 118.820 152.275 118.990 152.945 ;
        RECT 120.065 152.935 120.395 153.915 ;
        RECT 120.565 152.945 120.775 154.085 ;
        RECT 121.555 153.155 121.725 153.915 ;
        RECT 121.905 153.325 122.235 154.085 ;
        RECT 121.555 152.985 122.220 153.155 ;
        RECT 122.405 153.010 122.675 153.915 ;
        RECT 119.645 152.525 119.975 152.775 ;
        RECT 117.635 152.105 118.565 152.275 ;
        RECT 117.635 152.070 117.810 152.105 ;
        RECT 116.815 151.875 117.095 152.045 ;
        RECT 116.815 151.705 117.090 151.875 ;
        RECT 117.280 151.705 117.810 152.070 ;
        RECT 118.235 151.535 118.565 151.935 ;
        RECT 118.735 151.705 118.990 152.275 ;
        RECT 119.665 151.535 119.895 152.355 ;
        RECT 120.145 152.335 120.395 152.935 ;
        RECT 122.050 152.840 122.220 152.985 ;
        RECT 121.485 152.435 121.815 152.805 ;
        RECT 122.050 152.510 122.335 152.840 ;
        RECT 120.065 151.705 120.395 152.335 ;
        RECT 120.565 151.535 120.775 152.355 ;
        RECT 122.050 152.255 122.220 152.510 ;
        RECT 121.555 152.085 122.220 152.255 ;
        RECT 122.505 152.210 122.675 153.010 ;
        RECT 122.935 153.155 123.105 153.915 ;
        RECT 123.285 153.325 123.615 154.085 ;
        RECT 122.935 152.985 123.600 153.155 ;
        RECT 123.785 153.010 124.055 153.915 ;
        RECT 123.430 152.840 123.600 152.985 ;
        RECT 122.865 152.435 123.195 152.805 ;
        RECT 123.430 152.510 123.715 152.840 ;
        RECT 123.430 152.255 123.600 152.510 ;
        RECT 121.555 151.705 121.725 152.085 ;
        RECT 121.905 151.535 122.235 151.915 ;
        RECT 122.415 151.705 122.675 152.210 ;
        RECT 122.935 152.085 123.600 152.255 ;
        RECT 123.885 152.210 124.055 153.010 ;
        RECT 124.685 152.995 126.355 154.085 ;
        RECT 126.525 152.995 127.735 154.085 ;
        RECT 124.685 152.475 125.435 152.995 ;
        RECT 125.605 152.305 126.355 152.825 ;
        RECT 126.525 152.455 127.045 152.995 ;
        RECT 122.935 151.705 123.105 152.085 ;
        RECT 123.285 151.535 123.615 151.915 ;
        RECT 123.795 151.705 124.055 152.210 ;
        RECT 124.685 151.535 126.355 152.305 ;
        RECT 127.215 152.285 127.735 152.825 ;
        RECT 126.525 151.535 127.735 152.285 ;
        RECT 14.660 151.365 127.820 151.535 ;
        RECT 14.745 150.615 15.955 151.365 ;
        RECT 14.745 150.075 15.265 150.615 ;
        RECT 17.105 150.545 17.315 151.365 ;
        RECT 17.485 150.565 17.815 151.195 ;
        RECT 15.435 149.905 15.955 150.445 ;
        RECT 17.485 149.965 17.735 150.565 ;
        RECT 17.985 150.545 18.215 151.365 ;
        RECT 18.465 150.545 18.695 151.365 ;
        RECT 18.865 150.565 19.195 151.195 ;
        RECT 17.905 150.125 18.235 150.375 ;
        RECT 18.445 150.125 18.775 150.375 ;
        RECT 18.945 149.965 19.195 150.565 ;
        RECT 19.365 150.545 19.575 151.365 ;
        RECT 20.180 150.655 20.435 151.185 ;
        RECT 20.615 150.905 20.900 151.365 ;
        RECT 20.180 150.005 20.360 150.655 ;
        RECT 21.080 150.455 21.330 151.105 ;
        RECT 20.530 150.125 21.330 150.455 ;
        RECT 14.745 148.815 15.955 149.905 ;
        RECT 17.105 148.815 17.315 149.955 ;
        RECT 17.485 148.985 17.815 149.965 ;
        RECT 17.985 148.815 18.215 149.955 ;
        RECT 18.465 148.815 18.695 149.955 ;
        RECT 18.865 148.985 19.195 149.965 ;
        RECT 19.365 148.815 19.575 149.955 ;
        RECT 20.095 149.835 20.360 150.005 ;
        RECT 20.180 149.795 20.360 149.835 ;
        RECT 20.180 149.125 20.435 149.795 ;
        RECT 20.615 148.815 20.900 149.615 ;
        RECT 21.080 149.535 21.330 150.125 ;
        RECT 21.530 150.770 21.850 151.100 ;
        RECT 22.030 150.885 22.690 151.365 ;
        RECT 22.890 150.975 23.740 151.145 ;
        RECT 21.530 149.875 21.720 150.770 ;
        RECT 22.040 150.445 22.700 150.715 ;
        RECT 22.370 150.385 22.700 150.445 ;
        RECT 21.890 150.215 22.220 150.275 ;
        RECT 22.890 150.215 23.060 150.975 ;
        RECT 24.300 150.905 24.620 151.365 ;
        RECT 24.820 150.725 25.070 151.155 ;
        RECT 25.360 150.925 25.770 151.365 ;
        RECT 25.940 150.985 26.955 151.185 ;
        RECT 23.230 150.555 24.480 150.725 ;
        RECT 23.230 150.435 23.560 150.555 ;
        RECT 21.890 150.045 23.790 150.215 ;
        RECT 21.530 149.705 23.450 149.875 ;
        RECT 21.530 149.685 21.850 149.705 ;
        RECT 21.080 149.025 21.410 149.535 ;
        RECT 21.680 149.075 21.850 149.685 ;
        RECT 23.620 149.535 23.790 150.045 ;
        RECT 23.960 149.975 24.140 150.385 ;
        RECT 24.310 149.795 24.480 150.555 ;
        RECT 22.020 148.815 22.350 149.505 ;
        RECT 22.580 149.365 23.790 149.535 ;
        RECT 23.960 149.485 24.480 149.795 ;
        RECT 24.650 150.385 25.070 150.725 ;
        RECT 25.360 150.385 25.770 150.715 ;
        RECT 24.650 149.615 24.840 150.385 ;
        RECT 25.940 150.255 26.110 150.985 ;
        RECT 27.255 150.815 27.425 151.145 ;
        RECT 27.595 150.985 27.925 151.365 ;
        RECT 26.280 150.435 26.630 150.805 ;
        RECT 25.940 150.215 26.360 150.255 ;
        RECT 25.010 150.045 26.360 150.215 ;
        RECT 25.010 149.885 25.260 150.045 ;
        RECT 25.770 149.615 26.020 149.875 ;
        RECT 24.650 149.365 26.020 149.615 ;
        RECT 22.580 149.075 22.820 149.365 ;
        RECT 23.620 149.285 23.790 149.365 ;
        RECT 23.020 148.815 23.440 149.195 ;
        RECT 23.620 149.035 24.250 149.285 ;
        RECT 24.720 148.815 25.050 149.195 ;
        RECT 25.220 149.075 25.390 149.365 ;
        RECT 26.190 149.200 26.360 150.045 ;
        RECT 26.810 149.875 27.030 150.745 ;
        RECT 27.255 150.625 27.950 150.815 ;
        RECT 26.530 149.495 27.030 149.875 ;
        RECT 27.200 149.825 27.610 150.445 ;
        RECT 27.780 149.655 27.950 150.625 ;
        RECT 27.255 149.485 27.950 149.655 ;
        RECT 25.570 148.815 25.950 149.195 ;
        RECT 26.190 149.030 27.020 149.200 ;
        RECT 27.255 148.985 27.425 149.485 ;
        RECT 27.595 148.815 27.925 149.315 ;
        RECT 28.140 148.985 28.365 151.105 ;
        RECT 28.535 150.985 28.865 151.365 ;
        RECT 29.035 150.815 29.205 151.105 ;
        RECT 28.540 150.645 29.205 150.815 ;
        RECT 29.465 150.690 29.725 151.195 ;
        RECT 29.905 150.985 30.235 151.365 ;
        RECT 30.415 150.815 30.585 151.195 ;
        RECT 28.540 149.655 28.770 150.645 ;
        RECT 28.940 149.825 29.290 150.475 ;
        RECT 29.465 149.890 29.635 150.690 ;
        RECT 29.920 150.645 30.585 150.815 ;
        RECT 29.920 150.390 30.090 150.645 ;
        RECT 30.845 150.595 33.435 151.365 ;
        RECT 29.805 150.060 30.090 150.390 ;
        RECT 30.325 150.095 30.655 150.465 ;
        RECT 29.920 149.915 30.090 150.060 ;
        RECT 28.540 149.485 29.205 149.655 ;
        RECT 28.535 148.815 28.865 149.315 ;
        RECT 29.035 148.985 29.205 149.485 ;
        RECT 29.465 148.985 29.735 149.890 ;
        RECT 29.920 149.745 30.585 149.915 ;
        RECT 29.905 148.815 30.235 149.575 ;
        RECT 30.415 148.985 30.585 149.745 ;
        RECT 30.845 149.905 32.055 150.425 ;
        RECT 32.225 150.075 33.435 150.595 ;
        RECT 33.810 150.585 34.310 151.195 ;
        RECT 33.605 150.125 33.955 150.375 ;
        RECT 34.140 149.955 34.310 150.585 ;
        RECT 34.940 150.715 35.270 151.195 ;
        RECT 35.440 150.905 35.665 151.365 ;
        RECT 35.835 150.715 36.165 151.195 ;
        RECT 34.940 150.545 36.165 150.715 ;
        RECT 36.355 150.565 36.605 151.365 ;
        RECT 36.775 150.565 37.115 151.195 ;
        RECT 37.285 150.640 37.575 151.365 ;
        RECT 34.480 150.175 34.810 150.375 ;
        RECT 34.980 150.175 35.310 150.375 ;
        RECT 35.480 150.175 35.900 150.375 ;
        RECT 36.075 150.205 36.770 150.375 ;
        RECT 36.075 149.955 36.245 150.205 ;
        RECT 36.940 149.955 37.115 150.565 ;
        RECT 38.665 150.565 39.005 151.195 ;
        RECT 39.175 150.565 39.425 151.365 ;
        RECT 39.615 150.715 39.945 151.195 ;
        RECT 40.115 150.905 40.340 151.365 ;
        RECT 40.510 150.715 40.840 151.195 ;
        RECT 30.845 148.815 33.435 149.905 ;
        RECT 33.810 149.785 36.245 149.955 ;
        RECT 33.810 148.985 34.140 149.785 ;
        RECT 34.310 148.815 34.640 149.615 ;
        RECT 34.940 148.985 35.270 149.785 ;
        RECT 35.915 148.815 36.165 149.615 ;
        RECT 36.435 148.815 36.605 149.955 ;
        RECT 36.775 148.985 37.115 149.955 ;
        RECT 37.285 148.815 37.575 149.980 ;
        RECT 38.665 149.955 38.840 150.565 ;
        RECT 39.615 150.545 40.840 150.715 ;
        RECT 41.470 150.585 41.970 151.195 ;
        RECT 39.010 150.205 39.705 150.375 ;
        RECT 39.535 149.955 39.705 150.205 ;
        RECT 39.880 150.175 40.300 150.375 ;
        RECT 40.470 150.175 40.800 150.375 ;
        RECT 40.970 150.175 41.300 150.375 ;
        RECT 41.470 149.955 41.640 150.585 ;
        RECT 42.345 150.565 42.685 151.195 ;
        RECT 42.855 150.565 43.105 151.365 ;
        RECT 43.295 150.715 43.625 151.195 ;
        RECT 43.795 150.905 44.020 151.365 ;
        RECT 44.190 150.715 44.520 151.195 ;
        RECT 41.825 150.125 42.175 150.375 ;
        RECT 42.345 149.955 42.520 150.565 ;
        RECT 43.295 150.545 44.520 150.715 ;
        RECT 45.150 150.585 45.650 151.195 ;
        RECT 46.025 150.595 48.615 151.365 ;
        RECT 42.690 150.205 43.385 150.375 ;
        RECT 43.215 149.955 43.385 150.205 ;
        RECT 43.560 150.175 43.980 150.375 ;
        RECT 44.150 150.175 44.480 150.375 ;
        RECT 44.650 150.175 44.980 150.375 ;
        RECT 45.150 149.955 45.320 150.585 ;
        RECT 45.505 150.125 45.855 150.375 ;
        RECT 38.665 148.985 39.005 149.955 ;
        RECT 39.175 148.815 39.345 149.955 ;
        RECT 39.535 149.785 41.970 149.955 ;
        RECT 39.615 148.815 39.865 149.615 ;
        RECT 40.510 148.985 40.840 149.785 ;
        RECT 41.140 148.815 41.470 149.615 ;
        RECT 41.640 148.985 41.970 149.785 ;
        RECT 42.345 148.985 42.685 149.955 ;
        RECT 42.855 148.815 43.025 149.955 ;
        RECT 43.215 149.785 45.650 149.955 ;
        RECT 43.295 148.815 43.545 149.615 ;
        RECT 44.190 148.985 44.520 149.785 ;
        RECT 44.820 148.815 45.150 149.615 ;
        RECT 45.320 148.985 45.650 149.785 ;
        RECT 46.025 149.905 47.235 150.425 ;
        RECT 47.405 150.075 48.615 150.595 ;
        RECT 48.785 150.565 49.125 151.195 ;
        RECT 49.295 150.565 49.545 151.365 ;
        RECT 49.735 150.715 50.065 151.195 ;
        RECT 50.235 150.905 50.460 151.365 ;
        RECT 50.630 150.715 50.960 151.195 ;
        RECT 48.785 149.955 48.960 150.565 ;
        RECT 49.735 150.545 50.960 150.715 ;
        RECT 51.590 150.585 52.090 151.195 ;
        RECT 52.465 150.615 53.675 151.365 ;
        RECT 53.850 150.820 59.195 151.365 ;
        RECT 49.130 150.205 49.825 150.375 ;
        RECT 49.655 149.955 49.825 150.205 ;
        RECT 50.000 150.175 50.420 150.375 ;
        RECT 50.590 150.175 50.920 150.375 ;
        RECT 51.090 150.175 51.420 150.375 ;
        RECT 51.590 149.955 51.760 150.585 ;
        RECT 51.945 150.125 52.295 150.375 ;
        RECT 46.025 148.815 48.615 149.905 ;
        RECT 48.785 148.985 49.125 149.955 ;
        RECT 49.295 148.815 49.465 149.955 ;
        RECT 49.655 149.785 52.090 149.955 ;
        RECT 49.735 148.815 49.985 149.615 ;
        RECT 50.630 148.985 50.960 149.785 ;
        RECT 51.260 148.815 51.590 149.615 ;
        RECT 51.760 148.985 52.090 149.785 ;
        RECT 52.465 149.905 52.985 150.445 ;
        RECT 53.155 150.075 53.675 150.615 ;
        RECT 52.465 148.815 53.675 149.905 ;
        RECT 55.440 149.250 55.790 150.500 ;
        RECT 57.270 149.990 57.610 150.820 ;
        RECT 59.365 150.565 59.705 151.195 ;
        RECT 59.875 150.565 60.125 151.365 ;
        RECT 60.315 150.715 60.645 151.195 ;
        RECT 60.815 150.905 61.040 151.365 ;
        RECT 61.210 150.715 61.540 151.195 ;
        RECT 59.365 149.955 59.540 150.565 ;
        RECT 60.315 150.545 61.540 150.715 ;
        RECT 62.170 150.585 62.670 151.195 ;
        RECT 63.045 150.640 63.335 151.365 ;
        RECT 63.595 150.885 63.895 151.365 ;
        RECT 64.065 150.715 64.325 151.170 ;
        RECT 64.495 150.885 64.755 151.365 ;
        RECT 64.935 150.715 65.195 151.170 ;
        RECT 65.365 150.885 65.615 151.365 ;
        RECT 65.795 150.715 66.055 151.170 ;
        RECT 66.225 150.885 66.475 151.365 ;
        RECT 66.655 150.715 66.915 151.170 ;
        RECT 67.085 150.885 67.330 151.365 ;
        RECT 67.500 150.715 67.775 151.170 ;
        RECT 67.945 150.885 68.190 151.365 ;
        RECT 68.360 150.715 68.620 151.170 ;
        RECT 68.790 150.885 69.050 151.365 ;
        RECT 69.220 150.715 69.480 151.170 ;
        RECT 69.650 150.885 69.910 151.365 ;
        RECT 70.080 150.715 70.340 151.170 ;
        RECT 70.510 150.805 70.770 151.365 ;
        RECT 59.710 150.205 60.405 150.375 ;
        RECT 60.235 149.955 60.405 150.205 ;
        RECT 60.580 150.175 61.000 150.375 ;
        RECT 61.170 150.175 61.500 150.375 ;
        RECT 61.670 150.175 62.000 150.375 ;
        RECT 62.170 149.955 62.340 150.585 ;
        RECT 63.595 150.545 70.340 150.715 ;
        RECT 62.525 150.125 62.875 150.375 ;
        RECT 53.850 148.815 59.195 149.250 ;
        RECT 59.365 148.985 59.705 149.955 ;
        RECT 59.875 148.815 60.045 149.955 ;
        RECT 60.235 149.785 62.670 149.955 ;
        RECT 60.315 148.815 60.565 149.615 ;
        RECT 61.210 148.985 61.540 149.785 ;
        RECT 61.840 148.815 62.170 149.615 ;
        RECT 62.340 148.985 62.670 149.785 ;
        RECT 63.045 148.815 63.335 149.980 ;
        RECT 63.595 149.955 64.760 150.545 ;
        RECT 70.940 150.375 71.190 151.185 ;
        RECT 71.370 150.840 71.630 151.365 ;
        RECT 71.800 150.375 72.050 151.185 ;
        RECT 72.230 150.855 72.535 151.365 ;
        RECT 72.795 150.815 72.965 151.195 ;
        RECT 73.180 150.985 73.510 151.365 ;
        RECT 64.930 150.125 72.050 150.375 ;
        RECT 72.220 150.125 72.535 150.685 ;
        RECT 72.795 150.645 73.510 150.815 ;
        RECT 63.595 149.730 70.340 149.955 ;
        RECT 63.595 148.815 63.865 149.560 ;
        RECT 64.035 148.990 64.325 149.730 ;
        RECT 64.935 149.715 70.340 149.730 ;
        RECT 64.495 148.820 64.750 149.545 ;
        RECT 64.935 148.990 65.195 149.715 ;
        RECT 65.365 148.820 65.610 149.545 ;
        RECT 65.795 148.990 66.055 149.715 ;
        RECT 66.225 148.820 66.470 149.545 ;
        RECT 66.655 148.990 66.915 149.715 ;
        RECT 67.085 148.820 67.330 149.545 ;
        RECT 67.500 148.990 67.760 149.715 ;
        RECT 67.930 148.820 68.190 149.545 ;
        RECT 68.360 148.990 68.620 149.715 ;
        RECT 68.790 148.820 69.050 149.545 ;
        RECT 69.220 148.990 69.480 149.715 ;
        RECT 69.650 148.820 69.910 149.545 ;
        RECT 70.080 148.990 70.340 149.715 ;
        RECT 70.510 148.820 70.770 149.615 ;
        RECT 70.940 148.990 71.190 150.125 ;
        RECT 64.495 148.815 70.770 148.820 ;
        RECT 71.370 148.815 71.630 149.625 ;
        RECT 71.805 148.985 72.050 150.125 ;
        RECT 72.705 150.095 73.060 150.465 ;
        RECT 73.340 150.455 73.510 150.645 ;
        RECT 73.680 150.620 73.935 151.195 ;
        RECT 73.340 150.125 73.595 150.455 ;
        RECT 73.340 149.915 73.510 150.125 ;
        RECT 72.795 149.745 73.510 149.915 ;
        RECT 73.765 149.890 73.935 150.620 ;
        RECT 74.110 150.525 74.370 151.365 ;
        RECT 74.635 150.815 74.805 151.195 ;
        RECT 75.020 150.985 75.350 151.365 ;
        RECT 74.635 150.645 75.350 150.815 ;
        RECT 74.545 150.095 74.900 150.465 ;
        RECT 75.180 150.455 75.350 150.645 ;
        RECT 75.520 150.620 75.775 151.195 ;
        RECT 75.180 150.125 75.435 150.455 ;
        RECT 72.230 148.815 72.525 149.625 ;
        RECT 72.795 148.985 72.965 149.745 ;
        RECT 73.180 148.815 73.510 149.575 ;
        RECT 73.680 148.985 73.935 149.890 ;
        RECT 74.110 148.815 74.370 149.965 ;
        RECT 75.180 149.915 75.350 150.125 ;
        RECT 74.635 149.745 75.350 149.915 ;
        RECT 75.605 149.890 75.775 150.620 ;
        RECT 75.950 150.525 76.210 151.365 ;
        RECT 76.385 150.865 76.685 151.195 ;
        RECT 76.855 150.885 77.130 151.365 ;
        RECT 74.635 148.985 74.805 149.745 ;
        RECT 75.020 148.815 75.350 149.575 ;
        RECT 75.520 148.985 75.775 149.890 ;
        RECT 75.950 148.815 76.210 149.965 ;
        RECT 76.385 149.955 76.555 150.865 ;
        RECT 77.310 150.715 77.605 151.105 ;
        RECT 77.775 150.885 78.030 151.365 ;
        RECT 78.205 150.715 78.465 151.105 ;
        RECT 78.635 150.885 78.915 151.365 ;
        RECT 76.725 150.125 77.075 150.695 ;
        RECT 77.310 150.545 78.960 150.715 ;
        RECT 77.245 150.205 78.385 150.375 ;
        RECT 77.245 149.955 77.415 150.205 ;
        RECT 78.555 150.035 78.960 150.545 ;
        RECT 76.385 149.785 77.415 149.955 ;
        RECT 78.205 149.865 78.960 150.035 ;
        RECT 79.605 150.565 79.945 151.195 ;
        RECT 80.115 150.565 80.365 151.365 ;
        RECT 80.555 150.715 80.885 151.195 ;
        RECT 81.055 150.905 81.280 151.365 ;
        RECT 81.450 150.715 81.780 151.195 ;
        RECT 79.605 149.955 79.780 150.565 ;
        RECT 80.555 150.545 81.780 150.715 ;
        RECT 82.410 150.585 82.910 151.195 ;
        RECT 83.290 150.820 88.635 151.365 ;
        RECT 79.950 150.205 80.645 150.375 ;
        RECT 80.475 149.955 80.645 150.205 ;
        RECT 80.820 150.175 81.240 150.375 ;
        RECT 81.410 150.175 81.740 150.375 ;
        RECT 81.910 150.175 82.240 150.375 ;
        RECT 82.410 149.955 82.580 150.585 ;
        RECT 82.765 150.125 83.115 150.375 ;
        RECT 76.385 148.985 76.695 149.785 ;
        RECT 78.205 149.615 78.465 149.865 ;
        RECT 76.865 148.815 77.175 149.615 ;
        RECT 77.345 149.445 78.465 149.615 ;
        RECT 77.345 148.985 77.605 149.445 ;
        RECT 77.775 148.815 78.030 149.275 ;
        RECT 78.205 148.985 78.465 149.445 ;
        RECT 78.635 148.815 78.920 149.685 ;
        RECT 79.605 148.985 79.945 149.955 ;
        RECT 80.115 148.815 80.285 149.955 ;
        RECT 80.475 149.785 82.910 149.955 ;
        RECT 80.555 148.815 80.805 149.615 ;
        RECT 81.450 148.985 81.780 149.785 ;
        RECT 82.080 148.815 82.410 149.615 ;
        RECT 82.580 148.985 82.910 149.785 ;
        RECT 84.880 149.250 85.230 150.500 ;
        RECT 86.710 149.990 87.050 150.820 ;
        RECT 88.805 150.640 89.095 151.365 ;
        RECT 89.785 150.545 89.995 151.365 ;
        RECT 90.165 150.565 90.495 151.195 ;
        RECT 83.290 148.815 88.635 149.250 ;
        RECT 88.805 148.815 89.095 149.980 ;
        RECT 90.165 149.965 90.415 150.565 ;
        RECT 90.665 150.545 90.895 151.365 ;
        RECT 91.195 150.815 91.365 151.195 ;
        RECT 91.545 150.985 91.875 151.365 ;
        RECT 91.195 150.645 91.860 150.815 ;
        RECT 92.055 150.690 92.315 151.195 ;
        RECT 90.585 150.125 90.915 150.375 ;
        RECT 91.125 150.095 91.455 150.465 ;
        RECT 91.690 150.390 91.860 150.645 ;
        RECT 91.690 150.060 91.975 150.390 ;
        RECT 89.785 148.815 89.995 149.955 ;
        RECT 90.165 148.985 90.495 149.965 ;
        RECT 90.665 148.815 90.895 149.955 ;
        RECT 91.690 149.915 91.860 150.060 ;
        RECT 91.195 149.745 91.860 149.915 ;
        RECT 92.145 149.890 92.315 150.690 ;
        RECT 91.195 148.985 91.365 149.745 ;
        RECT 91.545 148.815 91.875 149.575 ;
        RECT 92.045 148.985 92.315 149.890 ;
        RECT 92.490 150.655 92.745 151.185 ;
        RECT 92.915 150.905 93.220 151.365 ;
        RECT 93.465 150.985 94.535 151.155 ;
        RECT 92.490 150.005 92.700 150.655 ;
        RECT 93.465 150.630 93.785 150.985 ;
        RECT 93.460 150.455 93.785 150.630 ;
        RECT 92.870 150.155 93.785 150.455 ;
        RECT 93.955 150.415 94.195 150.815 ;
        RECT 94.365 150.755 94.535 150.985 ;
        RECT 94.705 150.925 94.895 151.365 ;
        RECT 95.065 150.915 96.015 151.195 ;
        RECT 96.235 151.005 96.585 151.175 ;
        RECT 94.365 150.585 94.895 150.755 ;
        RECT 92.870 150.125 93.610 150.155 ;
        RECT 92.490 149.125 92.745 150.005 ;
        RECT 92.915 148.815 93.220 149.955 ;
        RECT 93.440 149.535 93.610 150.125 ;
        RECT 93.955 150.045 94.495 150.415 ;
        RECT 94.675 150.305 94.895 150.585 ;
        RECT 95.065 150.135 95.235 150.915 ;
        RECT 94.830 149.965 95.235 150.135 ;
        RECT 95.405 150.125 95.755 150.745 ;
        RECT 94.830 149.875 95.000 149.965 ;
        RECT 95.925 149.955 96.135 150.745 ;
        RECT 93.780 149.705 95.000 149.875 ;
        RECT 95.460 149.795 96.135 149.955 ;
        RECT 93.440 149.365 94.240 149.535 ;
        RECT 93.560 148.815 93.890 149.195 ;
        RECT 94.070 149.075 94.240 149.365 ;
        RECT 94.830 149.325 95.000 149.705 ;
        RECT 95.170 149.785 96.135 149.795 ;
        RECT 96.325 150.615 96.585 151.005 ;
        RECT 96.795 150.905 97.125 151.365 ;
        RECT 98.000 150.975 98.855 151.145 ;
        RECT 99.060 150.975 99.555 151.145 ;
        RECT 99.725 151.005 100.055 151.365 ;
        RECT 96.325 149.925 96.495 150.615 ;
        RECT 96.665 150.265 96.835 150.445 ;
        RECT 97.005 150.435 97.795 150.685 ;
        RECT 98.000 150.265 98.170 150.975 ;
        RECT 98.340 150.465 98.695 150.685 ;
        RECT 96.665 150.095 98.355 150.265 ;
        RECT 95.170 149.495 95.630 149.785 ;
        RECT 96.325 149.755 97.825 149.925 ;
        RECT 96.325 149.615 96.495 149.755 ;
        RECT 95.935 149.445 96.495 149.615 ;
        RECT 94.410 148.815 94.660 149.275 ;
        RECT 94.830 148.985 95.700 149.325 ;
        RECT 95.935 148.985 96.105 149.445 ;
        RECT 96.940 149.415 98.015 149.585 ;
        RECT 96.275 148.815 96.645 149.275 ;
        RECT 96.940 149.075 97.110 149.415 ;
        RECT 97.280 148.815 97.610 149.245 ;
        RECT 97.845 149.075 98.015 149.415 ;
        RECT 98.185 149.315 98.355 150.095 ;
        RECT 98.525 149.875 98.695 150.465 ;
        RECT 98.865 150.065 99.215 150.685 ;
        RECT 98.525 149.485 98.990 149.875 ;
        RECT 99.385 149.615 99.555 150.975 ;
        RECT 99.725 149.785 100.185 150.835 ;
        RECT 99.160 149.445 99.555 149.615 ;
        RECT 99.160 149.315 99.330 149.445 ;
        RECT 98.185 148.985 98.865 149.315 ;
        RECT 99.080 148.985 99.330 149.315 ;
        RECT 99.500 148.815 99.750 149.275 ;
        RECT 99.920 149.000 100.245 149.785 ;
        RECT 100.415 148.985 100.585 151.105 ;
        RECT 100.755 150.985 101.085 151.365 ;
        RECT 101.255 150.815 101.510 151.105 ;
        RECT 100.760 150.645 101.510 150.815 ;
        RECT 100.760 149.655 100.990 150.645 ;
        RECT 101.685 150.595 103.355 151.365 ;
        RECT 101.160 149.825 101.510 150.475 ;
        RECT 101.685 149.905 102.435 150.425 ;
        RECT 102.605 150.075 103.355 150.595 ;
        RECT 103.525 150.690 103.795 151.035 ;
        RECT 103.985 150.965 104.365 151.365 ;
        RECT 104.535 150.795 104.705 151.145 ;
        RECT 104.875 150.965 105.205 151.365 ;
        RECT 105.405 150.795 105.575 151.145 ;
        RECT 105.775 150.865 106.105 151.365 ;
        RECT 106.295 150.865 106.625 151.365 ;
        RECT 103.525 149.955 103.695 150.690 ;
        RECT 103.965 150.625 105.575 150.795 ;
        RECT 106.825 150.795 106.995 151.145 ;
        RECT 107.195 150.965 107.525 151.365 ;
        RECT 107.695 150.795 107.865 151.145 ;
        RECT 108.035 150.965 108.415 151.365 ;
        RECT 103.965 150.455 104.135 150.625 ;
        RECT 103.865 150.125 104.135 150.455 ;
        RECT 104.305 150.125 104.710 150.455 ;
        RECT 103.965 149.955 104.135 150.125 ;
        RECT 100.760 149.485 101.510 149.655 ;
        RECT 100.755 148.815 101.085 149.315 ;
        RECT 101.255 148.985 101.510 149.485 ;
        RECT 101.685 148.815 103.355 149.905 ;
        RECT 103.525 148.985 103.795 149.955 ;
        RECT 103.965 149.785 104.690 149.955 ;
        RECT 104.880 149.835 105.590 150.455 ;
        RECT 105.760 150.125 106.110 150.695 ;
        RECT 106.290 150.125 106.640 150.695 ;
        RECT 106.825 150.625 108.435 150.795 ;
        RECT 108.605 150.690 108.875 151.035 ;
        RECT 108.265 150.455 108.435 150.625 ;
        RECT 104.520 149.665 104.690 149.785 ;
        RECT 105.790 149.665 106.110 149.955 ;
        RECT 104.005 148.815 104.285 149.615 ;
        RECT 104.520 149.495 106.110 149.665 ;
        RECT 106.290 149.665 106.610 149.955 ;
        RECT 106.810 149.835 107.520 150.455 ;
        RECT 107.690 150.125 108.095 150.455 ;
        RECT 108.265 150.125 108.535 150.455 ;
        RECT 108.265 149.955 108.435 150.125 ;
        RECT 108.705 149.955 108.875 150.690 ;
        RECT 107.710 149.785 108.435 149.955 ;
        RECT 107.710 149.665 107.880 149.785 ;
        RECT 106.290 149.495 107.880 149.665 ;
        RECT 104.455 149.035 106.110 149.325 ;
        RECT 106.290 149.035 107.945 149.325 ;
        RECT 108.115 148.815 108.395 149.615 ;
        RECT 108.605 148.985 108.875 149.955 ;
        RECT 109.045 150.565 109.385 151.195 ;
        RECT 109.555 150.565 109.805 151.365 ;
        RECT 109.995 150.715 110.325 151.195 ;
        RECT 110.495 150.905 110.720 151.365 ;
        RECT 110.890 150.715 111.220 151.195 ;
        RECT 109.045 149.955 109.220 150.565 ;
        RECT 109.995 150.545 111.220 150.715 ;
        RECT 111.850 150.585 112.350 151.195 ;
        RECT 112.725 150.595 114.395 151.365 ;
        RECT 114.565 150.640 114.855 151.365 ;
        RECT 115.025 150.615 116.235 151.365 ;
        RECT 109.390 150.205 110.085 150.375 ;
        RECT 109.915 149.955 110.085 150.205 ;
        RECT 110.260 150.175 110.680 150.375 ;
        RECT 110.850 150.175 111.180 150.375 ;
        RECT 111.350 150.175 111.680 150.375 ;
        RECT 111.850 149.955 112.020 150.585 ;
        RECT 112.205 150.125 112.555 150.375 ;
        RECT 109.045 148.985 109.385 149.955 ;
        RECT 109.555 148.815 109.725 149.955 ;
        RECT 109.915 149.785 112.350 149.955 ;
        RECT 109.995 148.815 110.245 149.615 ;
        RECT 110.890 148.985 111.220 149.785 ;
        RECT 111.520 148.815 111.850 149.615 ;
        RECT 112.020 148.985 112.350 149.785 ;
        RECT 112.725 149.905 113.475 150.425 ;
        RECT 113.645 150.075 114.395 150.595 ;
        RECT 112.725 148.815 114.395 149.905 ;
        RECT 114.565 148.815 114.855 149.980 ;
        RECT 115.025 149.905 115.545 150.445 ;
        RECT 115.715 150.075 116.235 150.615 ;
        RECT 116.780 150.655 117.035 151.185 ;
        RECT 117.215 150.905 117.500 151.365 ;
        RECT 115.025 148.815 116.235 149.905 ;
        RECT 116.780 149.795 116.960 150.655 ;
        RECT 117.680 150.455 117.930 151.105 ;
        RECT 117.130 150.125 117.930 150.455 ;
        RECT 116.780 149.325 117.035 149.795 ;
        RECT 116.695 149.155 117.035 149.325 ;
        RECT 116.780 149.125 117.035 149.155 ;
        RECT 117.215 148.815 117.500 149.615 ;
        RECT 117.680 149.535 117.930 150.125 ;
        RECT 118.130 150.770 118.450 151.100 ;
        RECT 118.630 150.885 119.290 151.365 ;
        RECT 119.490 150.975 120.340 151.145 ;
        RECT 118.130 149.875 118.320 150.770 ;
        RECT 118.640 150.445 119.300 150.715 ;
        RECT 118.970 150.385 119.300 150.445 ;
        RECT 118.490 150.215 118.820 150.275 ;
        RECT 119.490 150.215 119.660 150.975 ;
        RECT 120.900 150.905 121.220 151.365 ;
        RECT 121.420 150.725 121.670 151.155 ;
        RECT 121.960 150.925 122.370 151.365 ;
        RECT 122.540 150.985 123.555 151.185 ;
        RECT 119.830 150.555 121.080 150.725 ;
        RECT 119.830 150.435 120.160 150.555 ;
        RECT 118.490 150.045 120.390 150.215 ;
        RECT 118.130 149.705 120.050 149.875 ;
        RECT 118.130 149.685 118.450 149.705 ;
        RECT 117.680 149.025 118.010 149.535 ;
        RECT 118.280 149.075 118.450 149.685 ;
        RECT 120.220 149.535 120.390 150.045 ;
        RECT 120.560 149.975 120.740 150.385 ;
        RECT 120.910 149.795 121.080 150.555 ;
        RECT 118.620 148.815 118.950 149.505 ;
        RECT 119.180 149.365 120.390 149.535 ;
        RECT 120.560 149.485 121.080 149.795 ;
        RECT 121.250 150.385 121.670 150.725 ;
        RECT 121.960 150.385 122.370 150.715 ;
        RECT 121.250 149.615 121.440 150.385 ;
        RECT 122.540 150.255 122.710 150.985 ;
        RECT 123.855 150.815 124.025 151.145 ;
        RECT 124.195 150.985 124.525 151.365 ;
        RECT 122.880 150.435 123.230 150.805 ;
        RECT 122.540 150.215 122.960 150.255 ;
        RECT 121.610 150.045 122.960 150.215 ;
        RECT 121.610 149.885 121.860 150.045 ;
        RECT 122.370 149.615 122.620 149.875 ;
        RECT 121.250 149.365 122.620 149.615 ;
        RECT 119.180 149.075 119.420 149.365 ;
        RECT 120.220 149.285 120.390 149.365 ;
        RECT 119.620 148.815 120.040 149.195 ;
        RECT 120.220 149.035 120.850 149.285 ;
        RECT 121.320 148.815 121.650 149.195 ;
        RECT 121.820 149.075 121.990 149.365 ;
        RECT 122.790 149.200 122.960 150.045 ;
        RECT 123.410 149.875 123.630 150.745 ;
        RECT 123.855 150.625 124.550 150.815 ;
        RECT 123.130 149.495 123.630 149.875 ;
        RECT 123.800 149.825 124.210 150.445 ;
        RECT 124.380 149.655 124.550 150.625 ;
        RECT 123.855 149.485 124.550 149.655 ;
        RECT 122.170 148.815 122.550 149.195 ;
        RECT 122.790 149.030 123.620 149.200 ;
        RECT 123.855 148.985 124.025 149.485 ;
        RECT 124.195 148.815 124.525 149.315 ;
        RECT 124.740 148.985 124.965 151.105 ;
        RECT 125.135 150.985 125.465 151.365 ;
        RECT 125.635 150.815 125.805 151.105 ;
        RECT 125.140 150.645 125.805 150.815 ;
        RECT 125.140 149.655 125.370 150.645 ;
        RECT 126.525 150.615 127.735 151.365 ;
        RECT 125.540 149.825 125.890 150.475 ;
        RECT 126.525 149.905 127.045 150.445 ;
        RECT 127.215 150.075 127.735 150.615 ;
        RECT 125.140 149.485 125.805 149.655 ;
        RECT 125.135 148.815 125.465 149.315 ;
        RECT 125.635 148.985 125.805 149.485 ;
        RECT 126.525 148.815 127.735 149.905 ;
        RECT 14.660 148.645 127.820 148.815 ;
        RECT 14.745 147.555 15.955 148.645 ;
        RECT 14.745 146.845 15.265 147.385 ;
        RECT 15.435 147.015 15.955 147.555 ;
        RECT 16.125 147.555 17.335 148.645 ;
        RECT 17.510 148.210 22.855 148.645 ;
        RECT 16.125 147.015 16.645 147.555 ;
        RECT 16.815 146.845 17.335 147.385 ;
        RECT 19.100 146.960 19.450 148.210 ;
        RECT 23.115 147.715 23.285 148.475 ;
        RECT 23.465 147.885 23.795 148.645 ;
        RECT 23.115 147.545 23.780 147.715 ;
        RECT 23.965 147.570 24.235 148.475 ;
        RECT 14.745 146.095 15.955 146.845 ;
        RECT 16.125 146.095 17.335 146.845 ;
        RECT 20.930 146.640 21.270 147.470 ;
        RECT 23.610 147.400 23.780 147.545 ;
        RECT 23.045 146.995 23.375 147.365 ;
        RECT 23.610 147.070 23.895 147.400 ;
        RECT 23.610 146.815 23.780 147.070 ;
        RECT 23.115 146.645 23.780 146.815 ;
        RECT 24.065 146.770 24.235 147.570 ;
        RECT 24.405 147.480 24.695 148.645 ;
        RECT 25.325 147.555 27.915 148.645 ;
        RECT 28.090 148.210 33.435 148.645 ;
        RECT 25.325 147.035 26.535 147.555 ;
        RECT 26.705 146.865 27.915 147.385 ;
        RECT 29.680 146.960 30.030 148.210 ;
        RECT 33.605 147.505 33.875 148.475 ;
        RECT 34.085 147.845 34.365 148.645 ;
        RECT 34.535 148.135 36.190 148.425 ;
        RECT 34.600 147.795 36.190 147.965 ;
        RECT 34.600 147.675 34.770 147.795 ;
        RECT 34.045 147.505 34.770 147.675 ;
        RECT 17.510 146.095 22.855 146.640 ;
        RECT 23.115 146.265 23.285 146.645 ;
        RECT 23.465 146.095 23.795 146.475 ;
        RECT 23.975 146.265 24.235 146.770 ;
        RECT 24.405 146.095 24.695 146.820 ;
        RECT 25.325 146.095 27.915 146.865 ;
        RECT 31.510 146.640 31.850 147.470 ;
        RECT 33.605 146.770 33.775 147.505 ;
        RECT 34.045 147.335 34.215 147.505 ;
        RECT 34.960 147.455 35.675 147.625 ;
        RECT 35.870 147.505 36.190 147.795 ;
        RECT 36.365 147.555 38.035 148.645 ;
        RECT 33.945 147.005 34.215 147.335 ;
        RECT 34.385 147.005 34.790 147.335 ;
        RECT 34.960 147.005 35.670 147.455 ;
        RECT 34.045 146.835 34.215 147.005 ;
        RECT 28.090 146.095 33.435 146.640 ;
        RECT 33.605 146.425 33.875 146.770 ;
        RECT 34.045 146.665 35.655 146.835 ;
        RECT 35.840 146.765 36.190 147.335 ;
        RECT 36.365 147.035 37.115 147.555 ;
        RECT 38.205 147.505 38.475 148.475 ;
        RECT 38.685 147.845 38.965 148.645 ;
        RECT 39.135 148.135 40.790 148.425 ;
        RECT 39.200 147.795 40.790 147.965 ;
        RECT 39.200 147.675 39.370 147.795 ;
        RECT 38.645 147.505 39.370 147.675 ;
        RECT 37.285 146.865 38.035 147.385 ;
        RECT 34.065 146.095 34.445 146.495 ;
        RECT 34.615 146.315 34.785 146.665 ;
        RECT 34.955 146.095 35.285 146.495 ;
        RECT 35.485 146.315 35.655 146.665 ;
        RECT 35.855 146.095 36.185 146.595 ;
        RECT 36.365 146.095 38.035 146.865 ;
        RECT 38.205 146.770 38.375 147.505 ;
        RECT 38.645 147.335 38.815 147.505 ;
        RECT 39.560 147.455 40.275 147.625 ;
        RECT 40.470 147.505 40.790 147.795 ;
        RECT 40.965 147.555 44.475 148.645 ;
        RECT 44.650 148.210 49.995 148.645 ;
        RECT 38.545 147.005 38.815 147.335 ;
        RECT 38.985 147.005 39.390 147.335 ;
        RECT 39.560 147.005 40.270 147.455 ;
        RECT 38.645 146.835 38.815 147.005 ;
        RECT 38.205 146.425 38.475 146.770 ;
        RECT 38.645 146.665 40.255 146.835 ;
        RECT 40.440 146.765 40.790 147.335 ;
        RECT 40.965 147.035 42.655 147.555 ;
        RECT 42.825 146.865 44.475 147.385 ;
        RECT 46.240 146.960 46.590 148.210 ;
        RECT 50.165 147.480 50.455 148.645 ;
        RECT 50.625 147.555 53.215 148.645 ;
        RECT 38.665 146.095 39.045 146.495 ;
        RECT 39.215 146.315 39.385 146.665 ;
        RECT 39.555 146.095 39.885 146.495 ;
        RECT 40.085 146.315 40.255 146.665 ;
        RECT 40.455 146.095 40.785 146.595 ;
        RECT 40.965 146.095 44.475 146.865 ;
        RECT 48.070 146.640 48.410 147.470 ;
        RECT 50.625 147.035 51.835 147.555 ;
        RECT 53.425 147.505 53.655 148.645 ;
        RECT 53.825 147.495 54.155 148.475 ;
        RECT 54.325 147.505 54.535 148.645 ;
        RECT 55.685 147.555 59.195 148.645 ;
        RECT 59.740 147.665 59.995 148.335 ;
        RECT 60.175 147.845 60.460 148.645 ;
        RECT 60.640 147.925 60.970 148.435 ;
        RECT 59.740 147.625 59.920 147.665 ;
        RECT 52.005 146.865 53.215 147.385 ;
        RECT 53.405 147.085 53.735 147.335 ;
        RECT 44.650 146.095 49.995 146.640 ;
        RECT 50.165 146.095 50.455 146.820 ;
        RECT 50.625 146.095 53.215 146.865 ;
        RECT 53.425 146.095 53.655 146.915 ;
        RECT 53.905 146.895 54.155 147.495 ;
        RECT 55.685 147.035 57.375 147.555 ;
        RECT 59.655 147.455 59.920 147.625 ;
        RECT 53.825 146.265 54.155 146.895 ;
        RECT 54.325 146.095 54.535 146.915 ;
        RECT 57.545 146.865 59.195 147.385 ;
        RECT 55.685 146.095 59.195 146.865 ;
        RECT 59.740 146.805 59.920 147.455 ;
        RECT 60.640 147.335 60.890 147.925 ;
        RECT 61.240 147.775 61.410 148.385 ;
        RECT 61.580 147.955 61.910 148.645 ;
        RECT 62.140 148.095 62.380 148.385 ;
        RECT 62.580 148.265 63.000 148.645 ;
        RECT 63.180 148.175 63.810 148.425 ;
        RECT 64.280 148.265 64.610 148.645 ;
        RECT 63.180 148.095 63.350 148.175 ;
        RECT 64.780 148.095 64.950 148.385 ;
        RECT 65.130 148.265 65.510 148.645 ;
        RECT 65.750 148.260 66.580 148.430 ;
        RECT 62.140 147.925 63.350 148.095 ;
        RECT 60.090 147.005 60.890 147.335 ;
        RECT 59.740 146.275 59.995 146.805 ;
        RECT 60.175 146.095 60.460 146.555 ;
        RECT 60.640 146.355 60.890 147.005 ;
        RECT 61.090 147.755 61.410 147.775 ;
        RECT 61.090 147.585 63.010 147.755 ;
        RECT 61.090 146.690 61.280 147.585 ;
        RECT 63.180 147.415 63.350 147.925 ;
        RECT 63.520 147.665 64.040 147.975 ;
        RECT 61.450 147.245 63.350 147.415 ;
        RECT 61.450 147.185 61.780 147.245 ;
        RECT 61.930 147.015 62.260 147.075 ;
        RECT 61.600 146.745 62.260 147.015 ;
        RECT 61.090 146.360 61.410 146.690 ;
        RECT 61.590 146.095 62.250 146.575 ;
        RECT 62.450 146.485 62.620 147.245 ;
        RECT 63.520 147.075 63.700 147.485 ;
        RECT 62.790 146.905 63.120 147.025 ;
        RECT 63.870 146.905 64.040 147.665 ;
        RECT 62.790 146.735 64.040 146.905 ;
        RECT 64.210 147.845 65.580 148.095 ;
        RECT 64.210 147.075 64.400 147.845 ;
        RECT 65.330 147.585 65.580 147.845 ;
        RECT 64.570 147.415 64.820 147.575 ;
        RECT 65.750 147.415 65.920 148.260 ;
        RECT 66.815 147.975 66.985 148.475 ;
        RECT 67.155 148.145 67.485 148.645 ;
        RECT 66.090 147.585 66.590 147.965 ;
        RECT 66.815 147.805 67.510 147.975 ;
        RECT 64.570 147.245 65.920 147.415 ;
        RECT 65.500 147.205 65.920 147.245 ;
        RECT 64.210 146.735 64.630 147.075 ;
        RECT 64.920 146.745 65.330 147.075 ;
        RECT 62.450 146.315 63.300 146.485 ;
        RECT 63.860 146.095 64.180 146.555 ;
        RECT 64.380 146.305 64.630 146.735 ;
        RECT 64.920 146.095 65.330 146.535 ;
        RECT 65.500 146.475 65.670 147.205 ;
        RECT 65.840 146.655 66.190 147.025 ;
        RECT 66.370 146.715 66.590 147.585 ;
        RECT 66.760 147.015 67.170 147.635 ;
        RECT 67.340 146.835 67.510 147.805 ;
        RECT 66.815 146.645 67.510 146.835 ;
        RECT 65.500 146.275 66.515 146.475 ;
        RECT 66.815 146.315 66.985 146.645 ;
        RECT 67.155 146.095 67.485 146.475 ;
        RECT 67.700 146.355 67.925 148.475 ;
        RECT 68.095 148.145 68.425 148.645 ;
        RECT 68.595 147.975 68.765 148.475 ;
        RECT 68.100 147.805 68.765 147.975 ;
        RECT 68.100 146.815 68.330 147.805 ;
        RECT 69.025 147.795 69.285 148.475 ;
        RECT 69.455 147.865 69.705 148.645 ;
        RECT 69.955 148.095 70.205 148.475 ;
        RECT 70.375 148.265 70.730 148.645 ;
        RECT 71.735 148.255 72.070 148.475 ;
        RECT 71.335 148.095 71.565 148.135 ;
        RECT 69.955 147.895 71.565 148.095 ;
        RECT 69.955 147.885 70.790 147.895 ;
        RECT 71.380 147.805 71.565 147.895 ;
        RECT 68.500 146.985 68.850 147.635 ;
        RECT 68.100 146.645 68.765 146.815 ;
        RECT 68.095 146.095 68.425 146.475 ;
        RECT 68.595 146.355 68.765 146.645 ;
        RECT 69.025 146.595 69.195 147.795 ;
        RECT 70.895 147.695 71.225 147.725 ;
        RECT 69.425 147.635 71.225 147.695 ;
        RECT 71.815 147.635 72.070 148.255 ;
        RECT 69.365 147.525 72.070 147.635 ;
        RECT 69.365 147.490 69.565 147.525 ;
        RECT 69.365 146.915 69.535 147.490 ;
        RECT 70.895 147.465 72.070 147.525 ;
        RECT 72.245 147.555 75.755 148.645 ;
        RECT 69.765 147.050 70.175 147.355 ;
        RECT 70.345 147.085 70.675 147.295 ;
        RECT 69.365 146.795 69.635 146.915 ;
        RECT 69.365 146.750 70.210 146.795 ;
        RECT 69.455 146.625 70.210 146.750 ;
        RECT 70.465 146.685 70.675 147.085 ;
        RECT 70.920 147.085 71.395 147.295 ;
        RECT 71.585 147.085 72.075 147.285 ;
        RECT 70.920 146.685 71.140 147.085 ;
        RECT 72.245 147.035 73.935 147.555 ;
        RECT 75.925 147.480 76.215 148.645 ;
        RECT 76.845 147.555 80.355 148.645 ;
        RECT 80.530 148.210 85.875 148.645 ;
        RECT 74.105 146.865 75.755 147.385 ;
        RECT 76.845 147.035 78.535 147.555 ;
        RECT 78.705 146.865 80.355 147.385 ;
        RECT 82.120 146.960 82.470 148.210 ;
        RECT 86.420 147.665 86.675 148.335 ;
        RECT 86.855 147.845 87.140 148.645 ;
        RECT 87.320 147.925 87.650 148.435 ;
        RECT 69.025 146.265 69.285 146.595 ;
        RECT 70.040 146.475 70.210 146.625 ;
        RECT 69.455 146.095 69.785 146.455 ;
        RECT 70.040 146.265 71.340 146.475 ;
        RECT 71.615 146.095 72.070 146.860 ;
        RECT 72.245 146.095 75.755 146.865 ;
        RECT 75.925 146.095 76.215 146.820 ;
        RECT 76.845 146.095 80.355 146.865 ;
        RECT 83.950 146.640 84.290 147.470 ;
        RECT 86.420 146.805 86.600 147.665 ;
        RECT 87.320 147.335 87.570 147.925 ;
        RECT 87.920 147.775 88.090 148.385 ;
        RECT 88.260 147.955 88.590 148.645 ;
        RECT 88.820 148.095 89.060 148.385 ;
        RECT 89.260 148.265 89.680 148.645 ;
        RECT 89.860 148.175 90.490 148.425 ;
        RECT 90.960 148.265 91.290 148.645 ;
        RECT 89.860 148.095 90.030 148.175 ;
        RECT 91.460 148.095 91.630 148.385 ;
        RECT 91.810 148.265 92.190 148.645 ;
        RECT 92.430 148.260 93.260 148.430 ;
        RECT 88.820 147.925 90.030 148.095 ;
        RECT 86.770 147.005 87.570 147.335 ;
        RECT 80.530 146.095 85.875 146.640 ;
        RECT 86.420 146.605 86.675 146.805 ;
        RECT 86.335 146.435 86.675 146.605 ;
        RECT 86.420 146.275 86.675 146.435 ;
        RECT 86.855 146.095 87.140 146.555 ;
        RECT 87.320 146.355 87.570 147.005 ;
        RECT 87.770 147.755 88.090 147.775 ;
        RECT 87.770 147.585 89.690 147.755 ;
        RECT 87.770 146.690 87.960 147.585 ;
        RECT 89.860 147.415 90.030 147.925 ;
        RECT 90.200 147.665 90.720 147.975 ;
        RECT 88.130 147.245 90.030 147.415 ;
        RECT 88.130 147.185 88.460 147.245 ;
        RECT 88.610 147.015 88.940 147.075 ;
        RECT 88.280 146.745 88.940 147.015 ;
        RECT 87.770 146.360 88.090 146.690 ;
        RECT 88.270 146.095 88.930 146.575 ;
        RECT 89.130 146.485 89.300 147.245 ;
        RECT 90.200 147.075 90.380 147.485 ;
        RECT 89.470 146.905 89.800 147.025 ;
        RECT 90.550 146.905 90.720 147.665 ;
        RECT 89.470 146.735 90.720 146.905 ;
        RECT 90.890 147.845 92.260 148.095 ;
        RECT 90.890 147.075 91.080 147.845 ;
        RECT 92.010 147.585 92.260 147.845 ;
        RECT 91.250 147.415 91.500 147.575 ;
        RECT 92.430 147.415 92.600 148.260 ;
        RECT 93.495 147.975 93.665 148.475 ;
        RECT 93.835 148.145 94.165 148.645 ;
        RECT 92.770 147.585 93.270 147.965 ;
        RECT 93.495 147.805 94.190 147.975 ;
        RECT 91.250 147.245 92.600 147.415 ;
        RECT 92.180 147.205 92.600 147.245 ;
        RECT 90.890 146.735 91.310 147.075 ;
        RECT 91.600 146.745 92.010 147.075 ;
        RECT 89.130 146.315 89.980 146.485 ;
        RECT 90.540 146.095 90.860 146.555 ;
        RECT 91.060 146.305 91.310 146.735 ;
        RECT 91.600 146.095 92.010 146.535 ;
        RECT 92.180 146.475 92.350 147.205 ;
        RECT 92.520 146.655 92.870 147.025 ;
        RECT 93.050 146.715 93.270 147.585 ;
        RECT 93.440 147.015 93.850 147.635 ;
        RECT 94.020 146.835 94.190 147.805 ;
        RECT 93.495 146.645 94.190 146.835 ;
        RECT 92.180 146.275 93.195 146.475 ;
        RECT 93.495 146.315 93.665 146.645 ;
        RECT 93.835 146.095 94.165 146.475 ;
        RECT 94.380 146.355 94.605 148.475 ;
        RECT 94.775 148.145 95.105 148.645 ;
        RECT 95.275 147.975 95.445 148.475 ;
        RECT 96.170 148.210 101.515 148.645 ;
        RECT 94.780 147.805 95.445 147.975 ;
        RECT 94.780 146.815 95.010 147.805 ;
        RECT 95.180 146.985 95.530 147.635 ;
        RECT 97.760 146.960 98.110 148.210 ;
        RECT 101.685 147.480 101.975 148.645 ;
        RECT 102.605 147.505 102.875 148.475 ;
        RECT 103.085 147.845 103.365 148.645 ;
        RECT 103.535 148.135 105.190 148.425 ;
        RECT 103.600 147.795 105.190 147.965 ;
        RECT 103.600 147.675 103.770 147.795 ;
        RECT 103.045 147.505 103.770 147.675 ;
        RECT 94.780 146.645 95.445 146.815 ;
        RECT 94.775 146.095 95.105 146.475 ;
        RECT 95.275 146.355 95.445 146.645 ;
        RECT 99.590 146.640 99.930 147.470 ;
        RECT 96.170 146.095 101.515 146.640 ;
        RECT 101.685 146.095 101.975 146.820 ;
        RECT 102.605 146.770 102.775 147.505 ;
        RECT 103.045 147.335 103.215 147.505 ;
        RECT 102.945 147.005 103.215 147.335 ;
        RECT 103.385 147.005 103.790 147.335 ;
        RECT 103.960 147.005 104.670 147.625 ;
        RECT 104.870 147.505 105.190 147.795 ;
        RECT 105.365 147.505 105.705 148.475 ;
        RECT 105.875 147.505 106.045 148.645 ;
        RECT 106.315 147.845 106.565 148.645 ;
        RECT 107.210 147.675 107.540 148.475 ;
        RECT 107.840 147.845 108.170 148.645 ;
        RECT 108.340 147.675 108.670 148.475 ;
        RECT 106.235 147.505 108.670 147.675 ;
        RECT 109.045 147.505 109.385 148.475 ;
        RECT 109.555 147.505 109.725 148.645 ;
        RECT 109.995 147.845 110.245 148.645 ;
        RECT 110.890 147.675 111.220 148.475 ;
        RECT 111.520 147.845 111.850 148.645 ;
        RECT 112.020 147.675 112.350 148.475 ;
        RECT 109.915 147.505 112.350 147.675 ;
        RECT 112.725 147.555 116.235 148.645 ;
        RECT 116.405 147.885 116.920 148.295 ;
        RECT 117.155 147.885 117.325 148.645 ;
        RECT 117.495 148.305 119.525 148.475 ;
        RECT 103.045 146.835 103.215 147.005 ;
        RECT 102.605 146.425 102.875 146.770 ;
        RECT 103.045 146.665 104.655 146.835 ;
        RECT 104.840 146.765 105.190 147.335 ;
        RECT 105.365 146.945 105.540 147.505 ;
        RECT 106.235 147.255 106.405 147.505 ;
        RECT 105.710 147.085 106.405 147.255 ;
        RECT 106.580 147.085 107.000 147.285 ;
        RECT 107.170 147.085 107.500 147.285 ;
        RECT 107.670 147.085 108.000 147.285 ;
        RECT 105.365 146.895 105.595 146.945 ;
        RECT 103.065 146.095 103.445 146.495 ;
        RECT 103.615 146.315 103.785 146.665 ;
        RECT 103.955 146.095 104.285 146.495 ;
        RECT 104.485 146.315 104.655 146.665 ;
        RECT 104.855 146.095 105.185 146.595 ;
        RECT 105.365 146.265 105.705 146.895 ;
        RECT 105.875 146.095 106.125 146.895 ;
        RECT 106.315 146.745 107.540 146.915 ;
        RECT 106.315 146.265 106.645 146.745 ;
        RECT 106.815 146.095 107.040 146.555 ;
        RECT 107.210 146.265 107.540 146.745 ;
        RECT 108.170 146.875 108.340 147.505 ;
        RECT 108.525 147.085 108.875 147.335 ;
        RECT 109.045 146.895 109.220 147.505 ;
        RECT 109.915 147.255 110.085 147.505 ;
        RECT 109.390 147.085 110.085 147.255 ;
        RECT 110.260 147.085 110.680 147.285 ;
        RECT 110.850 147.085 111.180 147.285 ;
        RECT 111.350 147.085 111.680 147.285 ;
        RECT 108.170 146.265 108.670 146.875 ;
        RECT 109.045 146.265 109.385 146.895 ;
        RECT 109.555 146.095 109.805 146.895 ;
        RECT 109.995 146.745 111.220 146.915 ;
        RECT 109.995 146.265 110.325 146.745 ;
        RECT 110.495 146.095 110.720 146.555 ;
        RECT 110.890 146.265 111.220 146.745 ;
        RECT 111.850 146.875 112.020 147.505 ;
        RECT 112.205 147.085 112.555 147.335 ;
        RECT 112.725 147.035 114.415 147.555 ;
        RECT 111.850 146.265 112.350 146.875 ;
        RECT 114.585 146.865 116.235 147.385 ;
        RECT 116.405 147.075 116.745 147.885 ;
        RECT 117.495 147.640 117.665 148.305 ;
        RECT 118.060 147.965 119.185 148.135 ;
        RECT 116.915 147.450 117.665 147.640 ;
        RECT 117.835 147.625 118.845 147.795 ;
        RECT 116.405 146.905 117.635 147.075 ;
        RECT 112.725 146.095 116.235 146.865 ;
        RECT 116.680 146.300 116.925 146.905 ;
        RECT 117.145 146.095 117.655 146.630 ;
        RECT 117.835 146.265 118.025 147.625 ;
        RECT 118.195 147.285 118.470 147.425 ;
        RECT 118.195 147.115 118.475 147.285 ;
        RECT 118.195 146.265 118.470 147.115 ;
        RECT 118.675 146.825 118.845 147.625 ;
        RECT 119.015 146.835 119.185 147.965 ;
        RECT 119.355 147.335 119.525 148.305 ;
        RECT 119.695 147.505 119.865 148.645 ;
        RECT 120.035 147.505 120.370 148.475 ;
        RECT 121.010 148.210 126.355 148.645 ;
        RECT 119.355 147.005 119.550 147.335 ;
        RECT 119.775 147.005 120.030 147.335 ;
        RECT 119.775 146.835 119.945 147.005 ;
        RECT 120.200 146.835 120.370 147.505 ;
        RECT 122.600 146.960 122.950 148.210 ;
        RECT 126.525 147.555 127.735 148.645 ;
        RECT 119.015 146.665 119.945 146.835 ;
        RECT 119.015 146.630 119.190 146.665 ;
        RECT 118.660 146.265 119.190 146.630 ;
        RECT 119.615 146.095 119.945 146.495 ;
        RECT 120.115 146.265 120.370 146.835 ;
        RECT 124.430 146.640 124.770 147.470 ;
        RECT 126.525 147.015 127.045 147.555 ;
        RECT 127.215 146.845 127.735 147.385 ;
        RECT 121.010 146.095 126.355 146.640 ;
        RECT 126.525 146.095 127.735 146.845 ;
        RECT 14.660 145.925 127.820 146.095 ;
        RECT 14.745 145.175 15.955 145.925 ;
        RECT 16.500 145.215 16.755 145.745 ;
        RECT 16.935 145.465 17.220 145.925 ;
        RECT 14.745 144.635 15.265 145.175 ;
        RECT 15.435 144.465 15.955 145.005 ;
        RECT 14.745 143.375 15.955 144.465 ;
        RECT 16.500 144.355 16.680 145.215 ;
        RECT 17.400 145.015 17.650 145.665 ;
        RECT 16.850 144.685 17.650 145.015 ;
        RECT 16.500 143.885 16.755 144.355 ;
        RECT 16.415 143.715 16.755 143.885 ;
        RECT 16.500 143.685 16.755 143.715 ;
        RECT 16.935 143.375 17.220 144.175 ;
        RECT 17.400 144.095 17.650 144.685 ;
        RECT 17.850 145.330 18.170 145.660 ;
        RECT 18.350 145.445 19.010 145.925 ;
        RECT 19.210 145.535 20.060 145.705 ;
        RECT 17.850 144.435 18.040 145.330 ;
        RECT 18.360 145.005 19.020 145.275 ;
        RECT 18.690 144.945 19.020 145.005 ;
        RECT 18.210 144.775 18.540 144.835 ;
        RECT 19.210 144.775 19.380 145.535 ;
        RECT 20.620 145.465 20.940 145.925 ;
        RECT 21.140 145.285 21.390 145.715 ;
        RECT 21.680 145.485 22.090 145.925 ;
        RECT 22.260 145.545 23.275 145.745 ;
        RECT 19.550 145.115 20.800 145.285 ;
        RECT 19.550 144.995 19.880 145.115 ;
        RECT 18.210 144.605 20.110 144.775 ;
        RECT 17.850 144.265 19.770 144.435 ;
        RECT 17.850 144.245 18.170 144.265 ;
        RECT 17.400 143.585 17.730 144.095 ;
        RECT 18.000 143.635 18.170 144.245 ;
        RECT 19.940 144.095 20.110 144.605 ;
        RECT 20.280 144.535 20.460 144.945 ;
        RECT 20.630 144.355 20.800 145.115 ;
        RECT 18.340 143.375 18.670 144.065 ;
        RECT 18.900 143.925 20.110 144.095 ;
        RECT 20.280 144.045 20.800 144.355 ;
        RECT 20.970 144.945 21.390 145.285 ;
        RECT 21.680 144.945 22.090 145.275 ;
        RECT 20.970 144.175 21.160 144.945 ;
        RECT 22.260 144.815 22.430 145.545 ;
        RECT 23.575 145.375 23.745 145.705 ;
        RECT 23.915 145.545 24.245 145.925 ;
        RECT 22.600 144.995 22.950 145.365 ;
        RECT 22.260 144.775 22.680 144.815 ;
        RECT 21.330 144.605 22.680 144.775 ;
        RECT 21.330 144.445 21.580 144.605 ;
        RECT 22.090 144.175 22.340 144.435 ;
        RECT 20.970 143.925 22.340 144.175 ;
        RECT 18.900 143.635 19.140 143.925 ;
        RECT 19.940 143.845 20.110 143.925 ;
        RECT 19.340 143.375 19.760 143.755 ;
        RECT 19.940 143.595 20.570 143.845 ;
        RECT 21.040 143.375 21.370 143.755 ;
        RECT 21.540 143.635 21.710 143.925 ;
        RECT 22.510 143.760 22.680 144.605 ;
        RECT 23.130 144.435 23.350 145.305 ;
        RECT 23.575 145.185 24.270 145.375 ;
        RECT 22.850 144.055 23.350 144.435 ;
        RECT 23.520 144.385 23.930 145.005 ;
        RECT 24.100 144.215 24.270 145.185 ;
        RECT 23.575 144.045 24.270 144.215 ;
        RECT 21.890 143.375 22.270 143.755 ;
        RECT 22.510 143.590 23.340 143.760 ;
        RECT 23.575 143.545 23.745 144.045 ;
        RECT 23.915 143.375 24.245 143.875 ;
        RECT 24.460 143.545 24.685 145.665 ;
        RECT 24.855 145.545 25.185 145.925 ;
        RECT 25.355 145.375 25.525 145.665 ;
        RECT 24.860 145.205 25.525 145.375 ;
        RECT 24.860 144.215 25.090 145.205 ;
        RECT 25.785 145.155 27.455 145.925 ;
        RECT 27.630 145.380 32.975 145.925 ;
        RECT 25.260 144.385 25.610 145.035 ;
        RECT 25.785 144.465 26.535 144.985 ;
        RECT 26.705 144.635 27.455 145.155 ;
        RECT 24.860 144.045 25.525 144.215 ;
        RECT 24.855 143.375 25.185 143.875 ;
        RECT 25.355 143.545 25.525 144.045 ;
        RECT 25.785 143.375 27.455 144.465 ;
        RECT 29.220 143.810 29.570 145.060 ;
        RECT 31.050 144.550 31.390 145.380 ;
        RECT 33.145 145.250 33.415 145.595 ;
        RECT 33.605 145.525 33.985 145.925 ;
        RECT 34.155 145.355 34.325 145.705 ;
        RECT 34.495 145.525 34.825 145.925 ;
        RECT 35.025 145.355 35.195 145.705 ;
        RECT 35.395 145.425 35.725 145.925 ;
        RECT 33.145 144.515 33.315 145.250 ;
        RECT 33.585 145.185 35.195 145.355 ;
        RECT 33.585 145.015 33.755 145.185 ;
        RECT 33.485 144.685 33.755 145.015 ;
        RECT 33.925 144.685 34.330 145.015 ;
        RECT 33.585 144.515 33.755 144.685 ;
        RECT 27.630 143.375 32.975 143.810 ;
        RECT 33.145 143.545 33.415 144.515 ;
        RECT 33.585 144.345 34.310 144.515 ;
        RECT 34.500 144.395 35.210 145.015 ;
        RECT 35.380 144.685 35.730 145.255 ;
        RECT 35.905 145.175 37.115 145.925 ;
        RECT 37.285 145.200 37.575 145.925 ;
        RECT 37.745 145.175 38.955 145.925 ;
        RECT 39.130 145.380 44.475 145.925 ;
        RECT 44.655 145.425 44.985 145.925 ;
        RECT 34.140 144.225 34.310 144.345 ;
        RECT 35.410 144.225 35.730 144.515 ;
        RECT 33.625 143.375 33.905 144.175 ;
        RECT 34.140 144.055 35.730 144.225 ;
        RECT 35.905 144.465 36.425 145.005 ;
        RECT 36.595 144.635 37.115 145.175 ;
        RECT 34.075 143.595 35.730 143.885 ;
        RECT 35.905 143.375 37.115 144.465 ;
        RECT 37.285 143.375 37.575 144.540 ;
        RECT 37.745 144.465 38.265 145.005 ;
        RECT 38.435 144.635 38.955 145.175 ;
        RECT 37.745 143.375 38.955 144.465 ;
        RECT 40.720 143.810 41.070 145.060 ;
        RECT 42.550 144.550 42.890 145.380 ;
        RECT 45.185 145.355 45.355 145.705 ;
        RECT 45.555 145.525 45.885 145.925 ;
        RECT 46.055 145.355 46.225 145.705 ;
        RECT 46.395 145.525 46.775 145.925 ;
        RECT 44.650 144.685 45.000 145.255 ;
        RECT 45.185 145.185 46.795 145.355 ;
        RECT 46.965 145.250 47.235 145.595 ;
        RECT 46.625 145.015 46.795 145.185 ;
        RECT 45.170 144.565 45.880 145.015 ;
        RECT 46.050 144.685 46.455 145.015 ;
        RECT 46.625 144.685 46.895 145.015 ;
        RECT 44.650 144.225 44.970 144.515 ;
        RECT 45.165 144.395 45.880 144.565 ;
        RECT 46.625 144.515 46.795 144.685 ;
        RECT 47.065 144.515 47.235 145.250 ;
        RECT 46.070 144.345 46.795 144.515 ;
        RECT 46.070 144.225 46.240 144.345 ;
        RECT 44.650 144.055 46.240 144.225 ;
        RECT 39.130 143.375 44.475 143.810 ;
        RECT 44.650 143.595 46.305 143.885 ;
        RECT 46.475 143.375 46.755 144.175 ;
        RECT 46.965 143.545 47.235 144.515 ;
        RECT 47.405 145.125 47.745 145.755 ;
        RECT 47.915 145.125 48.165 145.925 ;
        RECT 48.355 145.275 48.685 145.755 ;
        RECT 48.855 145.465 49.080 145.925 ;
        RECT 49.250 145.275 49.580 145.755 ;
        RECT 47.405 145.075 47.635 145.125 ;
        RECT 48.355 145.105 49.580 145.275 ;
        RECT 50.210 145.145 50.710 145.755 ;
        RECT 51.090 145.215 51.345 145.745 ;
        RECT 51.515 145.465 51.820 145.925 ;
        RECT 52.065 145.545 53.135 145.715 ;
        RECT 47.405 144.515 47.580 145.075 ;
        RECT 47.750 144.765 48.445 144.935 ;
        RECT 48.275 144.515 48.445 144.765 ;
        RECT 48.620 144.735 49.040 144.935 ;
        RECT 49.210 144.735 49.540 144.935 ;
        RECT 49.710 144.735 50.040 144.935 ;
        RECT 50.210 144.515 50.380 145.145 ;
        RECT 50.565 144.685 50.915 144.935 ;
        RECT 51.090 144.565 51.300 145.215 ;
        RECT 52.065 145.190 52.385 145.545 ;
        RECT 52.060 145.015 52.385 145.190 ;
        RECT 51.470 144.715 52.385 145.015 ;
        RECT 52.555 144.975 52.795 145.375 ;
        RECT 52.965 145.315 53.135 145.545 ;
        RECT 53.305 145.485 53.495 145.925 ;
        RECT 53.665 145.475 54.615 145.755 ;
        RECT 54.835 145.565 55.185 145.735 ;
        RECT 52.965 145.145 53.495 145.315 ;
        RECT 51.470 144.685 52.210 144.715 ;
        RECT 47.405 143.545 47.745 144.515 ;
        RECT 47.915 143.375 48.085 144.515 ;
        RECT 48.275 144.345 50.710 144.515 ;
        RECT 48.355 143.375 48.605 144.175 ;
        RECT 49.250 143.545 49.580 144.345 ;
        RECT 49.880 143.375 50.210 144.175 ;
        RECT 50.380 143.545 50.710 144.345 ;
        RECT 51.090 143.685 51.345 144.565 ;
        RECT 51.515 143.375 51.820 144.515 ;
        RECT 52.040 144.095 52.210 144.685 ;
        RECT 52.555 144.605 53.095 144.975 ;
        RECT 53.275 144.865 53.495 145.145 ;
        RECT 53.665 144.695 53.835 145.475 ;
        RECT 53.430 144.525 53.835 144.695 ;
        RECT 54.005 144.685 54.355 145.305 ;
        RECT 53.430 144.435 53.600 144.525 ;
        RECT 54.525 144.515 54.735 145.305 ;
        RECT 52.380 144.265 53.600 144.435 ;
        RECT 54.060 144.355 54.735 144.515 ;
        RECT 52.040 143.925 52.840 144.095 ;
        RECT 52.160 143.375 52.490 143.755 ;
        RECT 52.670 143.635 52.840 143.925 ;
        RECT 53.430 143.885 53.600 144.265 ;
        RECT 53.770 144.345 54.735 144.355 ;
        RECT 54.925 145.175 55.185 145.565 ;
        RECT 55.395 145.465 55.725 145.925 ;
        RECT 56.600 145.535 57.455 145.705 ;
        RECT 57.660 145.535 58.155 145.705 ;
        RECT 58.325 145.565 58.655 145.925 ;
        RECT 54.925 144.485 55.095 145.175 ;
        RECT 55.265 144.825 55.435 145.005 ;
        RECT 55.605 144.995 56.395 145.245 ;
        RECT 56.600 144.825 56.770 145.535 ;
        RECT 56.940 145.025 57.295 145.245 ;
        RECT 55.265 144.655 56.955 144.825 ;
        RECT 53.770 144.055 54.230 144.345 ;
        RECT 54.925 144.315 56.425 144.485 ;
        RECT 54.925 144.175 55.095 144.315 ;
        RECT 54.535 144.005 55.095 144.175 ;
        RECT 53.010 143.375 53.260 143.835 ;
        RECT 53.430 143.545 54.300 143.885 ;
        RECT 54.535 143.545 54.705 144.005 ;
        RECT 55.540 143.975 56.615 144.145 ;
        RECT 54.875 143.375 55.245 143.835 ;
        RECT 55.540 143.635 55.710 143.975 ;
        RECT 55.880 143.375 56.210 143.805 ;
        RECT 56.445 143.635 56.615 143.975 ;
        RECT 56.785 143.875 56.955 144.655 ;
        RECT 57.125 144.435 57.295 145.025 ;
        RECT 57.465 144.625 57.815 145.245 ;
        RECT 57.125 144.045 57.590 144.435 ;
        RECT 57.985 144.175 58.155 145.535 ;
        RECT 58.325 144.345 58.785 145.395 ;
        RECT 57.760 144.005 58.155 144.175 ;
        RECT 57.760 143.875 57.930 144.005 ;
        RECT 56.785 143.545 57.465 143.875 ;
        RECT 57.680 143.545 57.930 143.875 ;
        RECT 58.100 143.375 58.350 143.835 ;
        RECT 58.520 143.560 58.845 144.345 ;
        RECT 59.015 143.545 59.185 145.665 ;
        RECT 59.355 145.545 59.685 145.925 ;
        RECT 59.855 145.375 60.110 145.665 ;
        RECT 59.360 145.205 60.110 145.375 ;
        RECT 60.285 145.250 60.545 145.755 ;
        RECT 60.725 145.545 61.055 145.925 ;
        RECT 61.235 145.375 61.405 145.755 ;
        RECT 59.360 144.215 59.590 145.205 ;
        RECT 59.760 144.385 60.110 145.035 ;
        RECT 60.285 144.450 60.455 145.250 ;
        RECT 60.740 145.205 61.405 145.375 ;
        RECT 60.740 144.950 60.910 145.205 ;
        RECT 61.665 145.175 62.875 145.925 ;
        RECT 63.045 145.200 63.335 145.925 ;
        RECT 60.625 144.620 60.910 144.950 ;
        RECT 61.145 144.655 61.475 145.025 ;
        RECT 60.740 144.475 60.910 144.620 ;
        RECT 59.360 144.045 60.110 144.215 ;
        RECT 59.355 143.375 59.685 143.875 ;
        RECT 59.855 143.545 60.110 144.045 ;
        RECT 60.285 143.545 60.555 144.450 ;
        RECT 60.740 144.305 61.405 144.475 ;
        RECT 60.725 143.375 61.055 144.135 ;
        RECT 61.235 143.545 61.405 144.305 ;
        RECT 61.665 144.465 62.185 145.005 ;
        RECT 62.355 144.635 62.875 145.175 ;
        RECT 63.965 145.125 64.305 145.755 ;
        RECT 64.475 145.125 64.725 145.925 ;
        RECT 64.915 145.275 65.245 145.755 ;
        RECT 65.415 145.465 65.640 145.925 ;
        RECT 65.810 145.275 66.140 145.755 ;
        RECT 61.665 143.375 62.875 144.465 ;
        RECT 63.045 143.375 63.335 144.540 ;
        RECT 63.965 144.515 64.140 145.125 ;
        RECT 64.915 145.105 66.140 145.275 ;
        RECT 66.770 145.145 67.270 145.755 ;
        RECT 64.310 144.765 65.005 144.935 ;
        RECT 64.835 144.515 65.005 144.765 ;
        RECT 65.180 144.735 65.600 144.935 ;
        RECT 65.770 144.735 66.100 144.935 ;
        RECT 66.270 144.735 66.600 144.935 ;
        RECT 66.770 144.515 66.940 145.145 ;
        RECT 68.840 145.115 69.085 145.720 ;
        RECT 69.305 145.390 69.815 145.925 ;
        RECT 68.565 144.945 69.795 145.115 ;
        RECT 67.125 144.685 67.475 144.935 ;
        RECT 63.965 143.545 64.305 144.515 ;
        RECT 64.475 143.375 64.645 144.515 ;
        RECT 64.835 144.345 67.270 144.515 ;
        RECT 64.915 143.375 65.165 144.175 ;
        RECT 65.810 143.545 66.140 144.345 ;
        RECT 66.440 143.375 66.770 144.175 ;
        RECT 66.940 143.545 67.270 144.345 ;
        RECT 68.565 144.135 68.905 144.945 ;
        RECT 69.075 144.380 69.825 144.570 ;
        RECT 68.565 143.725 69.080 144.135 ;
        RECT 69.315 143.375 69.485 144.135 ;
        RECT 69.655 143.715 69.825 144.380 ;
        RECT 69.995 144.395 70.185 145.755 ;
        RECT 70.355 145.245 70.630 145.755 ;
        RECT 70.820 145.390 71.350 145.755 ;
        RECT 71.775 145.525 72.105 145.925 ;
        RECT 71.175 145.355 71.350 145.390 ;
        RECT 70.355 145.075 70.635 145.245 ;
        RECT 70.355 144.595 70.630 145.075 ;
        RECT 70.835 144.395 71.005 145.195 ;
        RECT 69.995 144.225 71.005 144.395 ;
        RECT 71.175 145.185 72.105 145.355 ;
        RECT 72.275 145.185 72.530 145.755 ;
        RECT 73.715 145.375 73.885 145.755 ;
        RECT 74.065 145.545 74.395 145.925 ;
        RECT 73.715 145.205 74.380 145.375 ;
        RECT 74.575 145.250 74.835 145.755 ;
        RECT 71.175 144.055 71.345 145.185 ;
        RECT 71.935 145.015 72.105 145.185 ;
        RECT 70.220 143.885 71.345 144.055 ;
        RECT 71.515 144.685 71.710 145.015 ;
        RECT 71.935 144.685 72.190 145.015 ;
        RECT 71.515 143.715 71.685 144.685 ;
        RECT 72.360 144.515 72.530 145.185 ;
        RECT 73.645 144.655 73.975 145.025 ;
        RECT 74.210 144.950 74.380 145.205 ;
        RECT 69.655 143.545 71.685 143.715 ;
        RECT 71.855 143.375 72.025 144.515 ;
        RECT 72.195 143.545 72.530 144.515 ;
        RECT 74.210 144.620 74.495 144.950 ;
        RECT 74.210 144.475 74.380 144.620 ;
        RECT 73.715 144.305 74.380 144.475 ;
        RECT 74.665 144.450 74.835 145.250 ;
        RECT 75.465 145.155 78.055 145.925 ;
        RECT 73.715 143.545 73.885 144.305 ;
        RECT 74.065 143.375 74.395 144.135 ;
        RECT 74.565 143.545 74.835 144.450 ;
        RECT 75.465 144.465 76.675 144.985 ;
        RECT 76.845 144.635 78.055 145.155 ;
        RECT 78.225 145.250 78.495 145.595 ;
        RECT 78.685 145.525 79.065 145.925 ;
        RECT 79.235 145.355 79.405 145.705 ;
        RECT 79.575 145.525 79.905 145.925 ;
        RECT 80.105 145.355 80.275 145.705 ;
        RECT 80.475 145.425 80.805 145.925 ;
        RECT 78.225 144.515 78.395 145.250 ;
        RECT 78.665 145.185 80.275 145.355 ;
        RECT 78.665 145.015 78.835 145.185 ;
        RECT 78.565 144.685 78.835 145.015 ;
        RECT 79.005 144.685 79.410 145.015 ;
        RECT 78.665 144.515 78.835 144.685 ;
        RECT 79.580 144.565 80.290 145.015 ;
        RECT 80.460 144.685 80.810 145.255 ;
        RECT 80.985 145.125 81.325 145.755 ;
        RECT 81.495 145.125 81.745 145.925 ;
        RECT 81.935 145.275 82.265 145.755 ;
        RECT 82.435 145.465 82.660 145.925 ;
        RECT 82.830 145.275 83.160 145.755 ;
        RECT 80.985 145.075 81.215 145.125 ;
        RECT 81.935 145.105 83.160 145.275 ;
        RECT 83.790 145.145 84.290 145.755 ;
        RECT 75.465 143.375 78.055 144.465 ;
        RECT 78.225 143.545 78.495 144.515 ;
        RECT 78.665 144.345 79.390 144.515 ;
        RECT 79.580 144.395 80.295 144.565 ;
        RECT 80.985 144.515 81.160 145.075 ;
        RECT 81.330 144.765 82.025 144.935 ;
        RECT 81.855 144.515 82.025 144.765 ;
        RECT 82.200 144.735 82.620 144.935 ;
        RECT 82.790 144.735 83.120 144.935 ;
        RECT 83.290 144.735 83.620 144.935 ;
        RECT 83.790 144.515 83.960 145.145 ;
        RECT 84.940 145.115 85.185 145.720 ;
        RECT 85.405 145.390 85.915 145.925 ;
        RECT 84.665 144.945 85.895 145.115 ;
        RECT 84.145 144.685 84.495 144.935 ;
        RECT 79.220 144.225 79.390 144.345 ;
        RECT 80.490 144.225 80.810 144.515 ;
        RECT 78.705 143.375 78.985 144.175 ;
        RECT 79.220 144.055 80.810 144.225 ;
        RECT 79.155 143.595 80.810 143.885 ;
        RECT 80.985 143.545 81.325 144.515 ;
        RECT 81.495 143.375 81.665 144.515 ;
        RECT 81.855 144.345 84.290 144.515 ;
        RECT 81.935 143.375 82.185 144.175 ;
        RECT 82.830 143.545 83.160 144.345 ;
        RECT 83.460 143.375 83.790 144.175 ;
        RECT 83.960 143.545 84.290 144.345 ;
        RECT 84.665 144.135 85.005 144.945 ;
        RECT 85.175 144.380 85.925 144.570 ;
        RECT 84.665 143.725 85.180 144.135 ;
        RECT 85.415 143.375 85.585 144.135 ;
        RECT 85.755 143.715 85.925 144.380 ;
        RECT 86.095 144.395 86.285 145.755 ;
        RECT 86.455 145.585 86.730 145.755 ;
        RECT 86.455 145.415 86.735 145.585 ;
        RECT 86.455 144.595 86.730 145.415 ;
        RECT 86.920 145.390 87.450 145.755 ;
        RECT 87.875 145.525 88.205 145.925 ;
        RECT 87.275 145.355 87.450 145.390 ;
        RECT 86.935 144.395 87.105 145.195 ;
        RECT 86.095 144.225 87.105 144.395 ;
        RECT 87.275 145.185 88.205 145.355 ;
        RECT 88.375 145.185 88.630 145.755 ;
        RECT 88.805 145.200 89.095 145.925 ;
        RECT 87.275 144.055 87.445 145.185 ;
        RECT 88.035 145.015 88.205 145.185 ;
        RECT 86.320 143.885 87.445 144.055 ;
        RECT 87.615 144.685 87.810 145.015 ;
        RECT 88.035 144.685 88.290 145.015 ;
        RECT 87.615 143.715 87.785 144.685 ;
        RECT 88.460 144.515 88.630 145.185 ;
        RECT 89.265 145.155 92.775 145.925 ;
        RECT 85.755 143.545 87.785 143.715 ;
        RECT 87.955 143.375 88.125 144.515 ;
        RECT 88.295 143.545 88.630 144.515 ;
        RECT 88.805 143.375 89.095 144.540 ;
        RECT 89.265 144.465 90.955 144.985 ;
        RECT 91.125 144.635 92.775 145.155 ;
        RECT 93.220 145.115 93.465 145.720 ;
        RECT 93.685 145.390 94.195 145.925 ;
        RECT 92.945 144.945 94.175 145.115 ;
        RECT 89.265 143.375 92.775 144.465 ;
        RECT 92.945 144.135 93.285 144.945 ;
        RECT 93.455 144.380 94.205 144.570 ;
        RECT 92.945 143.725 93.460 144.135 ;
        RECT 93.695 143.375 93.865 144.135 ;
        RECT 94.035 143.715 94.205 144.380 ;
        RECT 94.375 144.395 94.565 145.755 ;
        RECT 94.735 145.245 95.010 145.755 ;
        RECT 95.200 145.390 95.730 145.755 ;
        RECT 96.155 145.525 96.485 145.925 ;
        RECT 95.555 145.355 95.730 145.390 ;
        RECT 94.735 145.075 95.015 145.245 ;
        RECT 94.735 144.595 95.010 145.075 ;
        RECT 95.215 144.395 95.385 145.195 ;
        RECT 94.375 144.225 95.385 144.395 ;
        RECT 95.555 145.185 96.485 145.355 ;
        RECT 96.655 145.185 96.910 145.755 ;
        RECT 97.550 145.380 102.895 145.925 ;
        RECT 103.070 145.380 108.415 145.925 ;
        RECT 95.555 144.055 95.725 145.185 ;
        RECT 96.315 145.015 96.485 145.185 ;
        RECT 94.600 143.885 95.725 144.055 ;
        RECT 95.895 144.685 96.090 145.015 ;
        RECT 96.315 144.685 96.570 145.015 ;
        RECT 95.895 143.715 96.065 144.685 ;
        RECT 96.740 144.515 96.910 145.185 ;
        RECT 94.035 143.545 96.065 143.715 ;
        RECT 96.235 143.375 96.405 144.515 ;
        RECT 96.575 143.545 96.910 144.515 ;
        RECT 99.140 143.810 99.490 145.060 ;
        RECT 100.970 144.550 101.310 145.380 ;
        RECT 104.660 143.810 105.010 145.060 ;
        RECT 106.490 144.550 106.830 145.380 ;
        RECT 108.585 145.125 108.925 145.755 ;
        RECT 109.095 145.125 109.345 145.925 ;
        RECT 109.535 145.275 109.865 145.755 ;
        RECT 110.035 145.465 110.260 145.925 ;
        RECT 110.430 145.275 110.760 145.755 ;
        RECT 108.585 144.515 108.760 145.125 ;
        RECT 109.535 145.105 110.760 145.275 ;
        RECT 111.390 145.145 111.890 145.755 ;
        RECT 112.725 145.155 114.395 145.925 ;
        RECT 114.565 145.200 114.855 145.925 ;
        RECT 115.490 145.380 120.835 145.925 ;
        RECT 121.010 145.380 126.355 145.925 ;
        RECT 108.930 144.765 109.625 144.935 ;
        RECT 109.455 144.515 109.625 144.765 ;
        RECT 109.800 144.735 110.220 144.935 ;
        RECT 110.390 144.735 110.720 144.935 ;
        RECT 110.890 144.735 111.220 144.935 ;
        RECT 111.390 144.515 111.560 145.145 ;
        RECT 111.745 144.685 112.095 144.935 ;
        RECT 97.550 143.375 102.895 143.810 ;
        RECT 103.070 143.375 108.415 143.810 ;
        RECT 108.585 143.545 108.925 144.515 ;
        RECT 109.095 143.375 109.265 144.515 ;
        RECT 109.455 144.345 111.890 144.515 ;
        RECT 109.535 143.375 109.785 144.175 ;
        RECT 110.430 143.545 110.760 144.345 ;
        RECT 111.060 143.375 111.390 144.175 ;
        RECT 111.560 143.545 111.890 144.345 ;
        RECT 112.725 144.465 113.475 144.985 ;
        RECT 113.645 144.635 114.395 145.155 ;
        RECT 112.725 143.375 114.395 144.465 ;
        RECT 114.565 143.375 114.855 144.540 ;
        RECT 117.080 143.810 117.430 145.060 ;
        RECT 118.910 144.550 119.250 145.380 ;
        RECT 122.600 143.810 122.950 145.060 ;
        RECT 124.430 144.550 124.770 145.380 ;
        RECT 126.525 145.175 127.735 145.925 ;
        RECT 126.525 144.465 127.045 145.005 ;
        RECT 127.215 144.635 127.735 145.175 ;
        RECT 115.490 143.375 120.835 143.810 ;
        RECT 121.010 143.375 126.355 143.810 ;
        RECT 126.525 143.375 127.735 144.465 ;
        RECT 14.660 143.205 127.820 143.375 ;
        RECT 14.745 142.115 15.955 143.205 ;
        RECT 14.745 141.405 15.265 141.945 ;
        RECT 15.435 141.575 15.955 142.115 ;
        RECT 16.125 142.115 18.715 143.205 ;
        RECT 18.890 142.770 24.235 143.205 ;
        RECT 16.125 141.595 17.335 142.115 ;
        RECT 17.505 141.425 18.715 141.945 ;
        RECT 20.480 141.520 20.830 142.770 ;
        RECT 24.405 142.040 24.695 143.205 ;
        RECT 24.865 142.115 26.535 143.205 ;
        RECT 26.710 142.770 32.055 143.205 ;
        RECT 14.745 140.655 15.955 141.405 ;
        RECT 16.125 140.655 18.715 141.425 ;
        RECT 22.310 141.200 22.650 142.030 ;
        RECT 24.865 141.595 25.615 142.115 ;
        RECT 25.785 141.425 26.535 141.945 ;
        RECT 28.300 141.520 28.650 142.770 ;
        RECT 32.425 142.535 32.705 143.205 ;
        RECT 32.875 142.315 33.175 142.865 ;
        RECT 33.375 142.485 33.705 143.205 ;
        RECT 33.895 142.485 34.355 143.035 ;
        RECT 18.890 140.655 24.235 141.200 ;
        RECT 24.405 140.655 24.695 141.380 ;
        RECT 24.865 140.655 26.535 141.425 ;
        RECT 30.130 141.200 30.470 142.030 ;
        RECT 32.240 141.895 32.505 142.255 ;
        RECT 32.875 142.145 33.815 142.315 ;
        RECT 33.645 141.895 33.815 142.145 ;
        RECT 32.240 141.645 32.915 141.895 ;
        RECT 33.135 141.645 33.475 141.895 ;
        RECT 33.645 141.565 33.935 141.895 ;
        RECT 33.645 141.475 33.815 141.565 ;
        RECT 32.425 141.285 33.815 141.475 ;
        RECT 26.710 140.655 32.055 141.200 ;
        RECT 32.425 140.925 32.755 141.285 ;
        RECT 34.105 141.115 34.355 142.485 ;
        RECT 33.375 140.655 33.625 141.115 ;
        RECT 33.795 140.825 34.355 141.115 ;
        RECT 34.525 142.065 34.795 143.035 ;
        RECT 35.005 142.405 35.285 143.205 ;
        RECT 35.455 142.695 37.110 142.985 ;
        RECT 35.520 142.355 37.110 142.525 ;
        RECT 35.520 142.235 35.690 142.355 ;
        RECT 34.965 142.065 35.690 142.235 ;
        RECT 34.525 141.330 34.695 142.065 ;
        RECT 34.965 141.895 35.135 142.065 ;
        RECT 35.880 142.015 36.595 142.185 ;
        RECT 36.790 142.065 37.110 142.355 ;
        RECT 37.285 142.115 38.955 143.205 ;
        RECT 39.130 142.770 44.475 143.205 ;
        RECT 44.650 142.770 49.995 143.205 ;
        RECT 34.865 141.565 35.135 141.895 ;
        RECT 35.305 141.565 35.710 141.895 ;
        RECT 35.880 141.565 36.590 142.015 ;
        RECT 34.965 141.395 35.135 141.565 ;
        RECT 34.525 140.985 34.795 141.330 ;
        RECT 34.965 141.225 36.575 141.395 ;
        RECT 36.760 141.325 37.110 141.895 ;
        RECT 37.285 141.595 38.035 142.115 ;
        RECT 38.205 141.425 38.955 141.945 ;
        RECT 40.720 141.520 41.070 142.770 ;
        RECT 34.985 140.655 35.365 141.055 ;
        RECT 35.535 140.875 35.705 141.225 ;
        RECT 35.875 140.655 36.205 141.055 ;
        RECT 36.405 140.875 36.575 141.225 ;
        RECT 36.775 140.655 37.105 141.155 ;
        RECT 37.285 140.655 38.955 141.425 ;
        RECT 42.550 141.200 42.890 142.030 ;
        RECT 46.240 141.520 46.590 142.770 ;
        RECT 50.165 142.040 50.455 143.205 ;
        RECT 51.090 142.770 56.435 143.205 ;
        RECT 48.070 141.200 48.410 142.030 ;
        RECT 52.680 141.520 53.030 142.770 ;
        RECT 56.605 142.445 57.120 142.855 ;
        RECT 57.355 142.445 57.525 143.205 ;
        RECT 57.695 142.865 59.725 143.035 ;
        RECT 39.130 140.655 44.475 141.200 ;
        RECT 44.650 140.655 49.995 141.200 ;
        RECT 50.165 140.655 50.455 141.380 ;
        RECT 54.510 141.200 54.850 142.030 ;
        RECT 56.605 141.635 56.945 142.445 ;
        RECT 57.695 142.200 57.865 142.865 ;
        RECT 58.260 142.525 59.385 142.695 ;
        RECT 57.115 142.010 57.865 142.200 ;
        RECT 58.035 142.185 59.045 142.355 ;
        RECT 56.605 141.465 57.835 141.635 ;
        RECT 51.090 140.655 56.435 141.200 ;
        RECT 56.880 140.860 57.125 141.465 ;
        RECT 57.345 140.655 57.855 141.190 ;
        RECT 58.035 140.825 58.225 142.185 ;
        RECT 58.395 141.845 58.670 141.985 ;
        RECT 58.395 141.675 58.675 141.845 ;
        RECT 58.395 140.825 58.670 141.675 ;
        RECT 58.875 141.385 59.045 142.185 ;
        RECT 59.215 141.395 59.385 142.525 ;
        RECT 59.555 141.895 59.725 142.865 ;
        RECT 59.895 142.065 60.065 143.205 ;
        RECT 60.235 142.065 60.570 143.035 ;
        RECT 59.555 141.565 59.750 141.895 ;
        RECT 59.975 141.565 60.230 141.895 ;
        RECT 59.975 141.395 60.145 141.565 ;
        RECT 60.400 141.395 60.570 142.065 ;
        RECT 60.745 142.115 62.415 143.205 ;
        RECT 60.745 141.595 61.495 142.115 ;
        RECT 62.585 142.065 62.925 143.035 ;
        RECT 63.095 142.065 63.265 143.205 ;
        RECT 63.535 142.405 63.785 143.205 ;
        RECT 64.430 142.235 64.760 143.035 ;
        RECT 65.060 142.405 65.390 143.205 ;
        RECT 65.560 142.235 65.890 143.035 ;
        RECT 66.640 142.865 66.895 142.895 ;
        RECT 66.555 142.695 66.895 142.865 ;
        RECT 63.455 142.065 65.890 142.235 ;
        RECT 66.640 142.225 66.895 142.695 ;
        RECT 67.075 142.405 67.360 143.205 ;
        RECT 67.540 142.485 67.870 142.995 ;
        RECT 61.665 141.425 62.415 141.945 ;
        RECT 59.215 141.225 60.145 141.395 ;
        RECT 59.215 141.190 59.390 141.225 ;
        RECT 58.860 140.825 59.390 141.190 ;
        RECT 59.815 140.655 60.145 141.055 ;
        RECT 60.315 140.825 60.570 141.395 ;
        RECT 60.745 140.655 62.415 141.425 ;
        RECT 62.585 141.455 62.760 142.065 ;
        RECT 63.455 141.815 63.625 142.065 ;
        RECT 62.930 141.645 63.625 141.815 ;
        RECT 63.800 141.645 64.220 141.845 ;
        RECT 64.390 141.645 64.720 141.845 ;
        RECT 64.890 141.645 65.220 141.845 ;
        RECT 62.585 140.825 62.925 141.455 ;
        RECT 63.095 140.655 63.345 141.455 ;
        RECT 63.535 141.305 64.760 141.475 ;
        RECT 63.535 140.825 63.865 141.305 ;
        RECT 64.035 140.655 64.260 141.115 ;
        RECT 64.430 140.825 64.760 141.305 ;
        RECT 65.390 141.435 65.560 142.065 ;
        RECT 65.745 141.645 66.095 141.895 ;
        RECT 65.390 140.825 65.890 141.435 ;
        RECT 66.640 141.365 66.820 142.225 ;
        RECT 67.540 141.895 67.790 142.485 ;
        RECT 68.140 142.335 68.310 142.945 ;
        RECT 68.480 142.515 68.810 143.205 ;
        RECT 69.040 142.655 69.280 142.945 ;
        RECT 69.480 142.825 69.900 143.205 ;
        RECT 70.080 142.735 70.710 142.985 ;
        RECT 71.180 142.825 71.510 143.205 ;
        RECT 70.080 142.655 70.250 142.735 ;
        RECT 71.680 142.655 71.850 142.945 ;
        RECT 72.030 142.825 72.410 143.205 ;
        RECT 72.650 142.820 73.480 142.990 ;
        RECT 69.040 142.485 70.250 142.655 ;
        RECT 66.990 141.565 67.790 141.895 ;
        RECT 66.640 140.835 66.895 141.365 ;
        RECT 67.075 140.655 67.360 141.115 ;
        RECT 67.540 140.915 67.790 141.565 ;
        RECT 67.990 142.315 68.310 142.335 ;
        RECT 67.990 142.145 69.910 142.315 ;
        RECT 67.990 141.250 68.180 142.145 ;
        RECT 70.080 141.975 70.250 142.485 ;
        RECT 70.420 142.225 70.940 142.535 ;
        RECT 68.350 141.805 70.250 141.975 ;
        RECT 68.350 141.745 68.680 141.805 ;
        RECT 68.830 141.575 69.160 141.635 ;
        RECT 68.500 141.305 69.160 141.575 ;
        RECT 67.990 140.920 68.310 141.250 ;
        RECT 68.490 140.655 69.150 141.135 ;
        RECT 69.350 141.045 69.520 141.805 ;
        RECT 70.420 141.635 70.600 142.045 ;
        RECT 69.690 141.465 70.020 141.585 ;
        RECT 70.770 141.465 70.940 142.225 ;
        RECT 69.690 141.295 70.940 141.465 ;
        RECT 71.110 142.405 72.480 142.655 ;
        RECT 71.110 141.635 71.300 142.405 ;
        RECT 72.230 142.145 72.480 142.405 ;
        RECT 71.470 141.975 71.720 142.135 ;
        RECT 72.650 141.975 72.820 142.820 ;
        RECT 73.715 142.535 73.885 143.035 ;
        RECT 74.055 142.705 74.385 143.205 ;
        RECT 72.990 142.145 73.490 142.525 ;
        RECT 73.715 142.365 74.410 142.535 ;
        RECT 71.470 141.805 72.820 141.975 ;
        RECT 72.400 141.765 72.820 141.805 ;
        RECT 71.110 141.295 71.530 141.635 ;
        RECT 71.820 141.305 72.230 141.635 ;
        RECT 69.350 140.875 70.200 141.045 ;
        RECT 70.760 140.655 71.080 141.115 ;
        RECT 71.280 140.865 71.530 141.295 ;
        RECT 71.820 140.655 72.230 141.095 ;
        RECT 72.400 141.035 72.570 141.765 ;
        RECT 72.740 141.215 73.090 141.585 ;
        RECT 73.270 141.275 73.490 142.145 ;
        RECT 73.660 141.575 74.070 142.195 ;
        RECT 74.240 141.395 74.410 142.365 ;
        RECT 73.715 141.205 74.410 141.395 ;
        RECT 72.400 140.835 73.415 141.035 ;
        RECT 73.715 140.875 73.885 141.205 ;
        RECT 74.055 140.655 74.385 141.035 ;
        RECT 74.600 140.915 74.825 143.035 ;
        RECT 74.995 142.705 75.325 143.205 ;
        RECT 75.495 142.535 75.665 143.035 ;
        RECT 75.000 142.365 75.665 142.535 ;
        RECT 75.000 141.375 75.230 142.365 ;
        RECT 75.400 141.545 75.750 142.195 ;
        RECT 75.925 142.040 76.215 143.205 ;
        RECT 76.385 142.115 77.595 143.205 ;
        RECT 77.770 142.695 79.425 142.985 ;
        RECT 77.770 142.355 79.360 142.525 ;
        RECT 79.595 142.405 79.875 143.205 ;
        RECT 76.385 141.575 76.905 142.115 ;
        RECT 77.770 142.065 78.090 142.355 ;
        RECT 79.190 142.235 79.360 142.355 ;
        RECT 77.075 141.405 77.595 141.945 ;
        RECT 75.000 141.205 75.665 141.375 ;
        RECT 74.995 140.655 75.325 141.035 ;
        RECT 75.495 140.915 75.665 141.205 ;
        RECT 75.925 140.655 76.215 141.380 ;
        RECT 76.385 140.655 77.595 141.405 ;
        RECT 77.770 141.325 78.120 141.895 ;
        RECT 78.290 141.565 79.000 142.185 ;
        RECT 79.190 142.065 79.915 142.235 ;
        RECT 80.085 142.065 80.355 143.035 ;
        RECT 79.745 141.895 79.915 142.065 ;
        RECT 79.170 141.565 79.575 141.895 ;
        RECT 79.745 141.565 80.015 141.895 ;
        RECT 79.745 141.395 79.915 141.565 ;
        RECT 78.305 141.225 79.915 141.395 ;
        RECT 80.185 141.330 80.355 142.065 ;
        RECT 77.775 140.655 78.105 141.155 ;
        RECT 78.305 140.875 78.475 141.225 ;
        RECT 78.675 140.655 79.005 141.055 ;
        RECT 79.175 140.875 79.345 141.225 ;
        RECT 79.515 140.655 79.895 141.055 ;
        RECT 80.085 140.985 80.355 141.330 ;
        RECT 80.525 142.065 80.865 143.035 ;
        RECT 81.035 142.065 81.205 143.205 ;
        RECT 81.475 142.405 81.725 143.205 ;
        RECT 82.370 142.235 82.700 143.035 ;
        RECT 83.000 142.405 83.330 143.205 ;
        RECT 83.500 142.235 83.830 143.035 ;
        RECT 81.395 142.065 83.830 142.235 ;
        RECT 84.665 142.445 85.180 142.855 ;
        RECT 85.415 142.445 85.585 143.205 ;
        RECT 85.755 142.865 87.785 143.035 ;
        RECT 80.525 141.505 80.700 142.065 ;
        RECT 81.395 141.815 81.565 142.065 ;
        RECT 80.870 141.645 81.565 141.815 ;
        RECT 81.740 141.645 82.160 141.845 ;
        RECT 82.330 141.645 82.660 141.845 ;
        RECT 82.830 141.645 83.160 141.845 ;
        RECT 80.525 141.455 80.755 141.505 ;
        RECT 80.525 140.825 80.865 141.455 ;
        RECT 81.035 140.655 81.285 141.455 ;
        RECT 81.475 141.305 82.700 141.475 ;
        RECT 81.475 140.825 81.805 141.305 ;
        RECT 81.975 140.655 82.200 141.115 ;
        RECT 82.370 140.825 82.700 141.305 ;
        RECT 83.330 141.435 83.500 142.065 ;
        RECT 83.685 141.645 84.035 141.895 ;
        RECT 84.665 141.635 85.005 142.445 ;
        RECT 85.755 142.200 85.925 142.865 ;
        RECT 86.320 142.525 87.445 142.695 ;
        RECT 85.175 142.010 85.925 142.200 ;
        RECT 86.095 142.185 87.105 142.355 ;
        RECT 84.665 141.465 85.895 141.635 ;
        RECT 83.330 140.825 83.830 141.435 ;
        RECT 84.940 140.860 85.185 141.465 ;
        RECT 85.405 140.655 85.915 141.190 ;
        RECT 86.095 140.825 86.285 142.185 ;
        RECT 86.455 141.165 86.730 141.985 ;
        RECT 86.935 141.385 87.105 142.185 ;
        RECT 87.275 141.395 87.445 142.525 ;
        RECT 87.615 141.895 87.785 142.865 ;
        RECT 87.955 142.065 88.125 143.205 ;
        RECT 88.295 142.065 88.630 143.035 ;
        RECT 88.865 142.065 89.075 143.205 ;
        RECT 87.615 141.565 87.810 141.895 ;
        RECT 88.035 141.565 88.290 141.895 ;
        RECT 88.035 141.395 88.205 141.565 ;
        RECT 88.460 141.395 88.630 142.065 ;
        RECT 89.245 142.055 89.575 143.035 ;
        RECT 89.745 142.065 89.975 143.205 ;
        RECT 90.650 142.770 95.995 143.205 ;
        RECT 96.170 142.770 101.515 143.205 ;
        RECT 87.275 141.225 88.205 141.395 ;
        RECT 87.275 141.190 87.450 141.225 ;
        RECT 86.455 140.995 86.735 141.165 ;
        RECT 86.455 140.825 86.730 140.995 ;
        RECT 86.920 140.825 87.450 141.190 ;
        RECT 87.875 140.655 88.205 141.055 ;
        RECT 88.375 140.825 88.630 141.395 ;
        RECT 88.865 140.655 89.075 141.475 ;
        RECT 89.245 141.455 89.495 142.055 ;
        RECT 89.665 141.645 89.995 141.895 ;
        RECT 92.240 141.520 92.590 142.770 ;
        RECT 89.245 140.825 89.575 141.455 ;
        RECT 89.745 140.655 89.975 141.475 ;
        RECT 94.070 141.200 94.410 142.030 ;
        RECT 97.760 141.520 98.110 142.770 ;
        RECT 101.685 142.040 101.975 143.205 ;
        RECT 102.145 142.115 103.355 143.205 ;
        RECT 99.590 141.200 99.930 142.030 ;
        RECT 102.145 141.575 102.665 142.115 ;
        RECT 103.525 142.065 103.795 143.035 ;
        RECT 104.005 142.405 104.285 143.205 ;
        RECT 104.455 142.695 106.110 142.985 ;
        RECT 104.520 142.355 106.110 142.525 ;
        RECT 104.520 142.235 104.690 142.355 ;
        RECT 103.965 142.065 104.690 142.235 ;
        RECT 102.835 141.405 103.355 141.945 ;
        RECT 90.650 140.655 95.995 141.200 ;
        RECT 96.170 140.655 101.515 141.200 ;
        RECT 101.685 140.655 101.975 141.380 ;
        RECT 102.145 140.655 103.355 141.405 ;
        RECT 103.525 141.330 103.695 142.065 ;
        RECT 103.965 141.895 104.135 142.065 ;
        RECT 104.880 142.015 105.595 142.185 ;
        RECT 105.790 142.065 106.110 142.355 ;
        RECT 106.285 142.065 106.625 143.035 ;
        RECT 106.795 142.065 106.965 143.205 ;
        RECT 107.235 142.405 107.485 143.205 ;
        RECT 108.130 142.235 108.460 143.035 ;
        RECT 108.760 142.405 109.090 143.205 ;
        RECT 109.260 142.235 109.590 143.035 ;
        RECT 107.155 142.065 109.590 142.235 ;
        RECT 110.425 142.115 112.095 143.205 ;
        RECT 112.265 142.445 112.780 142.855 ;
        RECT 113.015 142.445 113.185 143.205 ;
        RECT 113.355 142.865 115.385 143.035 ;
        RECT 103.865 141.565 104.135 141.895 ;
        RECT 104.305 141.565 104.710 141.895 ;
        RECT 104.880 141.565 105.590 142.015 ;
        RECT 103.965 141.395 104.135 141.565 ;
        RECT 103.525 140.985 103.795 141.330 ;
        RECT 103.965 141.225 105.575 141.395 ;
        RECT 105.760 141.325 106.110 141.895 ;
        RECT 106.285 141.455 106.460 142.065 ;
        RECT 107.155 141.815 107.325 142.065 ;
        RECT 106.630 141.645 107.325 141.815 ;
        RECT 107.500 141.645 107.920 141.845 ;
        RECT 108.090 141.645 108.420 141.845 ;
        RECT 108.590 141.645 108.920 141.845 ;
        RECT 103.985 140.655 104.365 141.055 ;
        RECT 104.535 140.875 104.705 141.225 ;
        RECT 104.875 140.655 105.205 141.055 ;
        RECT 105.405 140.875 105.575 141.225 ;
        RECT 105.775 140.655 106.105 141.155 ;
        RECT 106.285 140.825 106.625 141.455 ;
        RECT 106.795 140.655 107.045 141.455 ;
        RECT 107.235 141.305 108.460 141.475 ;
        RECT 107.235 140.825 107.565 141.305 ;
        RECT 107.735 140.655 107.960 141.115 ;
        RECT 108.130 140.825 108.460 141.305 ;
        RECT 109.090 141.435 109.260 142.065 ;
        RECT 109.445 141.645 109.795 141.895 ;
        RECT 110.425 141.595 111.175 142.115 ;
        RECT 109.090 140.825 109.590 141.435 ;
        RECT 111.345 141.425 112.095 141.945 ;
        RECT 112.265 141.635 112.605 142.445 ;
        RECT 113.355 142.200 113.525 142.865 ;
        RECT 113.920 142.525 115.045 142.695 ;
        RECT 112.775 142.010 113.525 142.200 ;
        RECT 113.695 142.185 114.705 142.355 ;
        RECT 112.265 141.465 113.495 141.635 ;
        RECT 110.425 140.655 112.095 141.425 ;
        RECT 112.540 140.860 112.785 141.465 ;
        RECT 113.005 140.655 113.515 141.190 ;
        RECT 113.695 140.825 113.885 142.185 ;
        RECT 114.055 141.845 114.330 141.985 ;
        RECT 114.055 141.675 114.335 141.845 ;
        RECT 114.055 140.825 114.330 141.675 ;
        RECT 114.535 141.385 114.705 142.185 ;
        RECT 114.875 141.395 115.045 142.525 ;
        RECT 115.215 141.895 115.385 142.865 ;
        RECT 115.555 142.065 115.725 143.205 ;
        RECT 115.895 142.065 116.230 143.035 ;
        RECT 115.215 141.565 115.410 141.895 ;
        RECT 115.635 141.565 115.890 141.895 ;
        RECT 115.635 141.395 115.805 141.565 ;
        RECT 116.060 141.395 116.230 142.065 ;
        RECT 114.875 141.225 115.805 141.395 ;
        RECT 114.875 141.190 115.050 141.225 ;
        RECT 114.520 140.825 115.050 141.190 ;
        RECT 115.475 140.655 115.805 141.055 ;
        RECT 115.975 140.825 116.230 141.395 ;
        RECT 116.410 142.065 116.745 143.035 ;
        RECT 116.915 142.065 117.085 143.205 ;
        RECT 117.255 142.865 119.285 143.035 ;
        RECT 116.410 141.395 116.580 142.065 ;
        RECT 117.255 141.895 117.425 142.865 ;
        RECT 116.750 141.565 117.005 141.895 ;
        RECT 117.230 141.565 117.425 141.895 ;
        RECT 117.595 142.525 118.720 142.695 ;
        RECT 116.835 141.395 117.005 141.565 ;
        RECT 117.595 141.395 117.765 142.525 ;
        RECT 116.410 140.825 116.665 141.395 ;
        RECT 116.835 141.225 117.765 141.395 ;
        RECT 117.935 142.185 118.945 142.355 ;
        RECT 117.935 141.385 118.105 142.185 ;
        RECT 118.310 141.845 118.585 141.985 ;
        RECT 118.305 141.675 118.585 141.845 ;
        RECT 117.590 141.190 117.765 141.225 ;
        RECT 116.835 140.655 117.165 141.055 ;
        RECT 117.590 140.825 118.120 141.190 ;
        RECT 118.310 140.825 118.585 141.675 ;
        RECT 118.755 140.825 118.945 142.185 ;
        RECT 119.115 142.200 119.285 142.865 ;
        RECT 119.455 142.445 119.625 143.205 ;
        RECT 119.860 142.445 120.375 142.855 ;
        RECT 119.115 142.010 119.865 142.200 ;
        RECT 120.035 141.635 120.375 142.445 ;
        RECT 120.585 142.065 120.815 143.205 ;
        RECT 120.985 142.055 121.315 143.035 ;
        RECT 121.485 142.065 121.695 143.205 ;
        RECT 122.845 142.115 126.355 143.205 ;
        RECT 126.525 142.115 127.735 143.205 ;
        RECT 120.565 141.645 120.895 141.895 ;
        RECT 119.145 141.465 120.375 141.635 ;
        RECT 119.125 140.655 119.635 141.190 ;
        RECT 119.855 140.860 120.100 141.465 ;
        RECT 120.585 140.655 120.815 141.475 ;
        RECT 121.065 141.455 121.315 142.055 ;
        RECT 122.845 141.595 124.535 142.115 ;
        RECT 120.985 140.825 121.315 141.455 ;
        RECT 121.485 140.655 121.695 141.475 ;
        RECT 124.705 141.425 126.355 141.945 ;
        RECT 126.525 141.575 127.045 142.115 ;
        RECT 122.845 140.655 126.355 141.425 ;
        RECT 127.215 141.405 127.735 141.945 ;
        RECT 126.525 140.655 127.735 141.405 ;
        RECT 14.660 140.485 127.820 140.655 ;
        RECT 14.745 139.735 15.955 140.485 ;
        RECT 16.960 139.775 17.215 140.305 ;
        RECT 17.395 140.025 17.680 140.485 ;
        RECT 14.745 139.195 15.265 139.735 ;
        RECT 15.435 139.025 15.955 139.565 ;
        RECT 14.745 137.935 15.955 139.025 ;
        RECT 16.960 138.915 17.140 139.775 ;
        RECT 17.860 139.575 18.110 140.225 ;
        RECT 17.310 139.245 18.110 139.575 ;
        RECT 16.960 138.445 17.215 138.915 ;
        RECT 16.875 138.275 17.215 138.445 ;
        RECT 16.960 138.245 17.215 138.275 ;
        RECT 17.395 137.935 17.680 138.735 ;
        RECT 17.860 138.655 18.110 139.245 ;
        RECT 18.310 139.890 18.630 140.220 ;
        RECT 18.810 140.005 19.470 140.485 ;
        RECT 19.670 140.095 20.520 140.265 ;
        RECT 18.310 138.995 18.500 139.890 ;
        RECT 18.820 139.565 19.480 139.835 ;
        RECT 19.150 139.505 19.480 139.565 ;
        RECT 18.670 139.335 19.000 139.395 ;
        RECT 19.670 139.335 19.840 140.095 ;
        RECT 21.080 140.025 21.400 140.485 ;
        RECT 21.600 139.845 21.850 140.275 ;
        RECT 22.140 140.045 22.550 140.485 ;
        RECT 22.720 140.105 23.735 140.305 ;
        RECT 20.010 139.675 21.260 139.845 ;
        RECT 20.010 139.555 20.340 139.675 ;
        RECT 18.670 139.165 20.570 139.335 ;
        RECT 18.310 138.825 20.230 138.995 ;
        RECT 18.310 138.805 18.630 138.825 ;
        RECT 17.860 138.145 18.190 138.655 ;
        RECT 18.460 138.195 18.630 138.805 ;
        RECT 20.400 138.655 20.570 139.165 ;
        RECT 20.740 139.095 20.920 139.505 ;
        RECT 21.090 138.915 21.260 139.675 ;
        RECT 18.800 137.935 19.130 138.625 ;
        RECT 19.360 138.485 20.570 138.655 ;
        RECT 20.740 138.605 21.260 138.915 ;
        RECT 21.430 139.505 21.850 139.845 ;
        RECT 22.140 139.505 22.550 139.835 ;
        RECT 21.430 138.735 21.620 139.505 ;
        RECT 22.720 139.375 22.890 140.105 ;
        RECT 24.035 139.935 24.205 140.265 ;
        RECT 24.375 140.105 24.705 140.485 ;
        RECT 23.060 139.555 23.410 139.925 ;
        RECT 22.720 139.335 23.140 139.375 ;
        RECT 21.790 139.165 23.140 139.335 ;
        RECT 21.790 139.005 22.040 139.165 ;
        RECT 22.550 138.735 22.800 138.995 ;
        RECT 21.430 138.485 22.800 138.735 ;
        RECT 19.360 138.195 19.600 138.485 ;
        RECT 20.400 138.405 20.570 138.485 ;
        RECT 19.800 137.935 20.220 138.315 ;
        RECT 20.400 138.155 21.030 138.405 ;
        RECT 21.500 137.935 21.830 138.315 ;
        RECT 22.000 138.195 22.170 138.485 ;
        RECT 22.970 138.320 23.140 139.165 ;
        RECT 23.590 138.995 23.810 139.865 ;
        RECT 24.035 139.745 24.730 139.935 ;
        RECT 23.310 138.615 23.810 138.995 ;
        RECT 23.980 138.945 24.390 139.565 ;
        RECT 24.560 138.775 24.730 139.745 ;
        RECT 24.035 138.605 24.730 138.775 ;
        RECT 22.350 137.935 22.730 138.315 ;
        RECT 22.970 138.150 23.800 138.320 ;
        RECT 24.035 138.105 24.205 138.605 ;
        RECT 24.375 137.935 24.705 138.435 ;
        RECT 24.920 138.105 25.145 140.225 ;
        RECT 25.315 140.105 25.645 140.485 ;
        RECT 25.815 139.935 25.985 140.225 ;
        RECT 25.320 139.765 25.985 139.935 ;
        RECT 25.320 138.775 25.550 139.765 ;
        RECT 26.705 139.715 30.215 140.485 ;
        RECT 25.720 138.945 26.070 139.595 ;
        RECT 26.705 139.025 28.395 139.545 ;
        RECT 28.565 139.195 30.215 139.715 ;
        RECT 30.585 139.855 30.915 140.215 ;
        RECT 31.535 140.025 31.785 140.485 ;
        RECT 31.955 140.025 32.515 140.315 ;
        RECT 30.585 139.665 31.975 139.855 ;
        RECT 31.805 139.575 31.975 139.665 ;
        RECT 30.400 139.245 31.075 139.495 ;
        RECT 31.295 139.245 31.635 139.495 ;
        RECT 31.805 139.245 32.095 139.575 ;
        RECT 25.320 138.605 25.985 138.775 ;
        RECT 25.315 137.935 25.645 138.435 ;
        RECT 25.815 138.105 25.985 138.605 ;
        RECT 26.705 137.935 30.215 139.025 ;
        RECT 30.400 138.885 30.665 139.245 ;
        RECT 31.805 138.995 31.975 139.245 ;
        RECT 31.035 138.825 31.975 138.995 ;
        RECT 30.585 137.935 30.865 138.605 ;
        RECT 31.035 138.275 31.335 138.825 ;
        RECT 32.265 138.655 32.515 140.025 ;
        RECT 32.885 139.855 33.215 140.215 ;
        RECT 33.835 140.025 34.085 140.485 ;
        RECT 34.255 140.025 34.815 140.315 ;
        RECT 32.885 139.665 34.275 139.855 ;
        RECT 34.105 139.575 34.275 139.665 ;
        RECT 32.700 139.245 33.375 139.495 ;
        RECT 33.595 139.245 33.935 139.495 ;
        RECT 34.105 139.245 34.395 139.575 ;
        RECT 32.700 138.885 32.965 139.245 ;
        RECT 34.105 138.995 34.275 139.245 ;
        RECT 31.535 137.935 31.865 138.655 ;
        RECT 32.055 138.105 32.515 138.655 ;
        RECT 33.335 138.825 34.275 138.995 ;
        RECT 32.885 137.935 33.165 138.605 ;
        RECT 33.335 138.275 33.635 138.825 ;
        RECT 34.565 138.655 34.815 140.025 ;
        RECT 35.185 139.855 35.515 140.215 ;
        RECT 36.135 140.025 36.385 140.485 ;
        RECT 36.555 140.025 37.115 140.315 ;
        RECT 35.185 139.665 36.575 139.855 ;
        RECT 36.405 139.575 36.575 139.665 ;
        RECT 35.000 139.245 35.675 139.495 ;
        RECT 35.895 139.245 36.235 139.495 ;
        RECT 36.405 139.245 36.695 139.575 ;
        RECT 35.000 138.885 35.265 139.245 ;
        RECT 36.405 138.995 36.575 139.245 ;
        RECT 33.835 137.935 34.165 138.655 ;
        RECT 34.355 138.105 34.815 138.655 ;
        RECT 35.635 138.825 36.575 138.995 ;
        RECT 35.185 137.935 35.465 138.605 ;
        RECT 35.635 138.275 35.935 138.825 ;
        RECT 36.865 138.655 37.115 140.025 ;
        RECT 37.285 139.760 37.575 140.485 ;
        RECT 38.205 139.715 39.875 140.485 ;
        RECT 40.050 139.940 45.395 140.485 ;
        RECT 36.135 137.935 36.465 138.655 ;
        RECT 36.655 138.105 37.115 138.655 ;
        RECT 37.285 137.935 37.575 139.100 ;
        RECT 38.205 139.025 38.955 139.545 ;
        RECT 39.125 139.195 39.875 139.715 ;
        RECT 38.205 137.935 39.875 139.025 ;
        RECT 41.640 138.370 41.990 139.620 ;
        RECT 43.470 139.110 43.810 139.940 ;
        RECT 45.765 139.855 46.095 140.215 ;
        RECT 46.715 140.025 46.965 140.485 ;
        RECT 47.135 140.025 47.695 140.315 ;
        RECT 45.765 139.665 47.155 139.855 ;
        RECT 46.985 139.575 47.155 139.665 ;
        RECT 45.580 139.245 46.255 139.495 ;
        RECT 46.475 139.245 46.815 139.495 ;
        RECT 46.985 139.245 47.275 139.575 ;
        RECT 45.580 138.885 45.845 139.245 ;
        RECT 46.985 138.995 47.155 139.245 ;
        RECT 46.215 138.825 47.155 138.995 ;
        RECT 40.050 137.935 45.395 138.370 ;
        RECT 45.765 137.935 46.045 138.605 ;
        RECT 46.215 138.275 46.515 138.825 ;
        RECT 47.445 138.655 47.695 140.025 ;
        RECT 47.865 139.735 49.075 140.485 ;
        RECT 49.255 139.985 49.585 140.485 ;
        RECT 49.785 139.915 49.955 140.265 ;
        RECT 50.155 140.085 50.485 140.485 ;
        RECT 50.655 139.915 50.825 140.265 ;
        RECT 50.995 140.085 51.375 140.485 ;
        RECT 46.715 137.935 47.045 138.655 ;
        RECT 47.235 138.105 47.695 138.655 ;
        RECT 47.865 139.025 48.385 139.565 ;
        RECT 48.555 139.195 49.075 139.735 ;
        RECT 49.250 139.245 49.600 139.815 ;
        RECT 49.785 139.745 51.395 139.915 ;
        RECT 51.565 139.810 51.835 140.155 ;
        RECT 51.225 139.575 51.395 139.745 ;
        RECT 49.770 139.125 50.480 139.575 ;
        RECT 50.650 139.245 51.055 139.575 ;
        RECT 51.225 139.245 51.495 139.575 ;
        RECT 47.865 137.935 49.075 139.025 ;
        RECT 49.250 138.785 49.570 139.075 ;
        RECT 49.765 138.955 50.480 139.125 ;
        RECT 51.225 139.075 51.395 139.245 ;
        RECT 51.665 139.075 51.835 139.810 ;
        RECT 50.670 138.905 51.395 139.075 ;
        RECT 50.670 138.785 50.840 138.905 ;
        RECT 49.250 138.615 50.840 138.785 ;
        RECT 49.250 138.155 50.905 138.445 ;
        RECT 51.075 137.935 51.355 138.735 ;
        RECT 51.565 138.105 51.835 139.075 ;
        RECT 52.005 139.685 52.345 140.315 ;
        RECT 52.515 139.685 52.765 140.485 ;
        RECT 52.955 139.835 53.285 140.315 ;
        RECT 53.455 140.025 53.680 140.485 ;
        RECT 53.850 139.835 54.180 140.315 ;
        RECT 52.005 139.635 52.235 139.685 ;
        RECT 52.955 139.665 54.180 139.835 ;
        RECT 54.810 139.705 55.310 140.315 ;
        RECT 52.005 139.075 52.180 139.635 ;
        RECT 52.350 139.325 53.045 139.495 ;
        RECT 52.875 139.075 53.045 139.325 ;
        RECT 53.220 139.295 53.640 139.495 ;
        RECT 53.810 139.295 54.140 139.495 ;
        RECT 54.310 139.295 54.640 139.495 ;
        RECT 54.810 139.075 54.980 139.705 ;
        RECT 56.420 139.675 56.665 140.280 ;
        RECT 56.885 139.950 57.395 140.485 ;
        RECT 56.145 139.505 57.375 139.675 ;
        RECT 55.165 139.245 55.515 139.495 ;
        RECT 52.005 138.105 52.345 139.075 ;
        RECT 52.515 137.935 52.685 139.075 ;
        RECT 52.875 138.905 55.310 139.075 ;
        RECT 52.955 137.935 53.205 138.735 ;
        RECT 53.850 138.105 54.180 138.905 ;
        RECT 54.480 137.935 54.810 138.735 ;
        RECT 54.980 138.105 55.310 138.905 ;
        RECT 56.145 138.695 56.485 139.505 ;
        RECT 56.655 138.940 57.405 139.130 ;
        RECT 56.145 138.285 56.660 138.695 ;
        RECT 56.895 137.935 57.065 138.695 ;
        RECT 57.235 138.275 57.405 138.940 ;
        RECT 57.575 138.955 57.765 140.315 ;
        RECT 57.935 140.145 58.210 140.315 ;
        RECT 57.935 139.975 58.215 140.145 ;
        RECT 57.935 139.155 58.210 139.975 ;
        RECT 58.400 139.950 58.930 140.315 ;
        RECT 59.355 140.085 59.685 140.485 ;
        RECT 58.755 139.915 58.930 139.950 ;
        RECT 58.415 138.955 58.585 139.755 ;
        RECT 57.575 138.785 58.585 138.955 ;
        RECT 58.755 139.745 59.685 139.915 ;
        RECT 59.855 139.745 60.110 140.315 ;
        RECT 60.375 139.935 60.545 140.315 ;
        RECT 60.725 140.105 61.055 140.485 ;
        RECT 60.375 139.765 61.040 139.935 ;
        RECT 61.235 139.810 61.495 140.315 ;
        RECT 58.755 138.615 58.925 139.745 ;
        RECT 59.515 139.575 59.685 139.745 ;
        RECT 57.800 138.445 58.925 138.615 ;
        RECT 59.095 139.245 59.290 139.575 ;
        RECT 59.515 139.245 59.770 139.575 ;
        RECT 59.095 138.275 59.265 139.245 ;
        RECT 59.940 139.075 60.110 139.745 ;
        RECT 60.305 139.215 60.635 139.585 ;
        RECT 60.870 139.510 61.040 139.765 ;
        RECT 57.235 138.105 59.265 138.275 ;
        RECT 59.435 137.935 59.605 139.075 ;
        RECT 59.775 138.105 60.110 139.075 ;
        RECT 60.870 139.180 61.155 139.510 ;
        RECT 60.870 139.035 61.040 139.180 ;
        RECT 60.375 138.865 61.040 139.035 ;
        RECT 61.325 139.010 61.495 139.810 ;
        RECT 61.665 139.735 62.875 140.485 ;
        RECT 63.045 139.760 63.335 140.485 ;
        RECT 60.375 138.105 60.545 138.865 ;
        RECT 60.725 137.935 61.055 138.695 ;
        RECT 61.225 138.105 61.495 139.010 ;
        RECT 61.665 139.025 62.185 139.565 ;
        RECT 62.355 139.195 62.875 139.735 ;
        RECT 63.965 139.715 66.555 140.485 ;
        RECT 66.730 139.940 72.075 140.485 ;
        RECT 61.665 137.935 62.875 139.025 ;
        RECT 63.045 137.935 63.335 139.100 ;
        RECT 63.965 139.025 65.175 139.545 ;
        RECT 65.345 139.195 66.555 139.715 ;
        RECT 63.965 137.935 66.555 139.025 ;
        RECT 68.320 138.370 68.670 139.620 ;
        RECT 70.150 139.110 70.490 139.940 ;
        RECT 72.305 139.665 72.515 140.485 ;
        RECT 72.685 139.685 73.015 140.315 ;
        RECT 72.685 139.085 72.935 139.685 ;
        RECT 73.185 139.665 73.415 140.485 ;
        RECT 73.630 139.940 78.975 140.485 ;
        RECT 79.520 140.145 79.775 140.305 ;
        RECT 79.435 139.975 79.775 140.145 ;
        RECT 79.955 140.025 80.240 140.485 ;
        RECT 73.105 139.245 73.435 139.495 ;
        RECT 66.730 137.935 72.075 138.370 ;
        RECT 72.305 137.935 72.515 139.075 ;
        RECT 72.685 138.105 73.015 139.085 ;
        RECT 73.185 137.935 73.415 139.075 ;
        RECT 75.220 138.370 75.570 139.620 ;
        RECT 77.050 139.110 77.390 139.940 ;
        RECT 79.520 139.775 79.775 139.975 ;
        RECT 79.520 138.915 79.700 139.775 ;
        RECT 80.420 139.575 80.670 140.225 ;
        RECT 79.870 139.245 80.670 139.575 ;
        RECT 73.630 137.935 78.975 138.370 ;
        RECT 79.520 138.245 79.775 138.915 ;
        RECT 79.955 137.935 80.240 138.735 ;
        RECT 80.420 138.655 80.670 139.245 ;
        RECT 80.870 139.890 81.190 140.220 ;
        RECT 81.370 140.005 82.030 140.485 ;
        RECT 82.230 140.095 83.080 140.265 ;
        RECT 80.870 138.995 81.060 139.890 ;
        RECT 81.380 139.565 82.040 139.835 ;
        RECT 81.710 139.505 82.040 139.565 ;
        RECT 81.230 139.335 81.560 139.395 ;
        RECT 82.230 139.335 82.400 140.095 ;
        RECT 83.640 140.025 83.960 140.485 ;
        RECT 84.160 139.845 84.410 140.275 ;
        RECT 84.700 140.045 85.110 140.485 ;
        RECT 85.280 140.105 86.295 140.305 ;
        RECT 82.570 139.675 83.820 139.845 ;
        RECT 82.570 139.555 82.900 139.675 ;
        RECT 81.230 139.165 83.130 139.335 ;
        RECT 80.870 138.825 82.790 138.995 ;
        RECT 80.870 138.805 81.190 138.825 ;
        RECT 80.420 138.145 80.750 138.655 ;
        RECT 81.020 138.195 81.190 138.805 ;
        RECT 82.960 138.655 83.130 139.165 ;
        RECT 83.300 139.095 83.480 139.505 ;
        RECT 83.650 138.915 83.820 139.675 ;
        RECT 81.360 137.935 81.690 138.625 ;
        RECT 81.920 138.485 83.130 138.655 ;
        RECT 83.300 138.605 83.820 138.915 ;
        RECT 83.990 139.505 84.410 139.845 ;
        RECT 84.700 139.505 85.110 139.835 ;
        RECT 83.990 138.735 84.180 139.505 ;
        RECT 85.280 139.375 85.450 140.105 ;
        RECT 86.595 139.935 86.765 140.265 ;
        RECT 86.935 140.105 87.265 140.485 ;
        RECT 85.620 139.555 85.970 139.925 ;
        RECT 85.280 139.335 85.700 139.375 ;
        RECT 84.350 139.165 85.700 139.335 ;
        RECT 84.350 139.005 84.600 139.165 ;
        RECT 85.110 138.735 85.360 138.995 ;
        RECT 83.990 138.485 85.360 138.735 ;
        RECT 81.920 138.195 82.160 138.485 ;
        RECT 82.960 138.405 83.130 138.485 ;
        RECT 82.360 137.935 82.780 138.315 ;
        RECT 82.960 138.155 83.590 138.405 ;
        RECT 84.060 137.935 84.390 138.315 ;
        RECT 84.560 138.195 84.730 138.485 ;
        RECT 85.530 138.320 85.700 139.165 ;
        RECT 86.150 138.995 86.370 139.865 ;
        RECT 86.595 139.745 87.290 139.935 ;
        RECT 85.870 138.615 86.370 138.995 ;
        RECT 86.540 138.945 86.950 139.565 ;
        RECT 87.120 138.775 87.290 139.745 ;
        RECT 86.595 138.605 87.290 138.775 ;
        RECT 84.910 137.935 85.290 138.315 ;
        RECT 85.530 138.150 86.360 138.320 ;
        RECT 86.595 138.105 86.765 138.605 ;
        RECT 86.935 137.935 87.265 138.435 ;
        RECT 87.480 138.105 87.705 140.225 ;
        RECT 87.875 140.105 88.205 140.485 ;
        RECT 88.375 139.935 88.545 140.225 ;
        RECT 87.880 139.765 88.545 139.935 ;
        RECT 87.880 138.775 88.110 139.765 ;
        RECT 88.805 139.760 89.095 140.485 ;
        RECT 89.265 139.810 89.525 140.315 ;
        RECT 89.705 140.105 90.035 140.485 ;
        RECT 90.215 139.935 90.385 140.315 ;
        RECT 91.110 139.940 96.455 140.485 ;
        RECT 96.635 139.985 96.965 140.485 ;
        RECT 88.280 138.945 88.630 139.595 ;
        RECT 87.880 138.605 88.545 138.775 ;
        RECT 87.875 137.935 88.205 138.435 ;
        RECT 88.375 138.105 88.545 138.605 ;
        RECT 88.805 137.935 89.095 139.100 ;
        RECT 89.265 139.010 89.435 139.810 ;
        RECT 89.720 139.765 90.385 139.935 ;
        RECT 89.720 139.510 89.890 139.765 ;
        RECT 89.605 139.180 89.890 139.510 ;
        RECT 90.125 139.215 90.455 139.585 ;
        RECT 89.720 139.035 89.890 139.180 ;
        RECT 89.265 138.105 89.535 139.010 ;
        RECT 89.720 138.865 90.385 139.035 ;
        RECT 89.705 137.935 90.035 138.695 ;
        RECT 90.215 138.105 90.385 138.865 ;
        RECT 92.700 138.370 93.050 139.620 ;
        RECT 94.530 139.110 94.870 139.940 ;
        RECT 97.165 139.915 97.335 140.265 ;
        RECT 97.535 140.085 97.865 140.485 ;
        RECT 98.035 139.915 98.205 140.265 ;
        RECT 98.375 140.085 98.755 140.485 ;
        RECT 96.630 139.245 96.980 139.815 ;
        RECT 97.165 139.745 98.775 139.915 ;
        RECT 98.945 139.810 99.215 140.155 ;
        RECT 98.605 139.575 98.775 139.745 ;
        RECT 97.150 139.125 97.860 139.575 ;
        RECT 98.030 139.245 98.435 139.575 ;
        RECT 98.605 139.245 98.875 139.575 ;
        RECT 96.630 138.785 96.950 139.075 ;
        RECT 97.145 138.955 97.860 139.125 ;
        RECT 98.605 139.075 98.775 139.245 ;
        RECT 99.045 139.075 99.215 139.810 ;
        RECT 98.050 138.905 98.775 139.075 ;
        RECT 98.050 138.785 98.220 138.905 ;
        RECT 96.630 138.615 98.220 138.785 ;
        RECT 91.110 137.935 96.455 138.370 ;
        RECT 96.630 138.155 98.285 138.445 ;
        RECT 98.455 137.935 98.735 138.735 ;
        RECT 98.945 138.105 99.215 139.075 ;
        RECT 99.385 139.685 99.725 140.315 ;
        RECT 99.895 139.685 100.145 140.485 ;
        RECT 100.335 139.835 100.665 140.315 ;
        RECT 100.835 140.025 101.060 140.485 ;
        RECT 101.230 139.835 101.560 140.315 ;
        RECT 99.385 139.635 99.615 139.685 ;
        RECT 100.335 139.665 101.560 139.835 ;
        RECT 102.190 139.705 102.690 140.315 ;
        RECT 103.525 139.810 103.795 140.155 ;
        RECT 103.985 140.085 104.365 140.485 ;
        RECT 104.535 139.915 104.705 140.265 ;
        RECT 104.875 140.085 105.205 140.485 ;
        RECT 105.405 139.915 105.575 140.265 ;
        RECT 105.775 139.985 106.105 140.485 ;
        RECT 99.385 139.075 99.560 139.635 ;
        RECT 99.730 139.325 100.425 139.495 ;
        RECT 100.255 139.075 100.425 139.325 ;
        RECT 100.600 139.295 101.020 139.495 ;
        RECT 101.190 139.295 101.520 139.495 ;
        RECT 101.690 139.295 102.020 139.495 ;
        RECT 102.190 139.075 102.360 139.705 ;
        RECT 102.545 139.245 102.895 139.495 ;
        RECT 103.525 139.075 103.695 139.810 ;
        RECT 103.965 139.745 105.575 139.915 ;
        RECT 103.965 139.575 104.135 139.745 ;
        RECT 103.865 139.245 104.135 139.575 ;
        RECT 104.305 139.245 104.710 139.575 ;
        RECT 103.965 139.075 104.135 139.245 ;
        RECT 99.385 138.105 99.725 139.075 ;
        RECT 99.895 137.935 100.065 139.075 ;
        RECT 100.255 138.905 102.690 139.075 ;
        RECT 100.335 137.935 100.585 138.735 ;
        RECT 101.230 138.105 101.560 138.905 ;
        RECT 101.860 137.935 102.190 138.735 ;
        RECT 102.360 138.105 102.690 138.905 ;
        RECT 103.525 138.105 103.795 139.075 ;
        RECT 103.965 138.905 104.690 139.075 ;
        RECT 104.880 138.955 105.590 139.575 ;
        RECT 105.760 139.245 106.110 139.815 ;
        RECT 106.285 139.735 107.495 140.485 ;
        RECT 104.520 138.785 104.690 138.905 ;
        RECT 105.790 138.785 106.110 139.075 ;
        RECT 104.005 137.935 104.285 138.735 ;
        RECT 104.520 138.615 106.110 138.785 ;
        RECT 106.285 139.025 106.805 139.565 ;
        RECT 106.975 139.195 107.495 139.735 ;
        RECT 107.940 139.675 108.185 140.280 ;
        RECT 108.405 139.950 108.915 140.485 ;
        RECT 107.665 139.505 108.895 139.675 ;
        RECT 104.455 138.155 106.110 138.445 ;
        RECT 106.285 137.935 107.495 139.025 ;
        RECT 107.665 138.695 108.005 139.505 ;
        RECT 108.175 138.940 108.925 139.130 ;
        RECT 107.665 138.285 108.180 138.695 ;
        RECT 108.415 137.935 108.585 138.695 ;
        RECT 108.755 138.275 108.925 138.940 ;
        RECT 109.095 138.955 109.285 140.315 ;
        RECT 109.455 139.805 109.730 140.315 ;
        RECT 109.920 139.950 110.450 140.315 ;
        RECT 110.875 140.085 111.205 140.485 ;
        RECT 110.275 139.915 110.450 139.950 ;
        RECT 109.455 139.635 109.735 139.805 ;
        RECT 109.455 139.155 109.730 139.635 ;
        RECT 109.935 138.955 110.105 139.755 ;
        RECT 109.095 138.785 110.105 138.955 ;
        RECT 110.275 139.745 111.205 139.915 ;
        RECT 111.375 139.745 111.630 140.315 ;
        RECT 110.275 138.615 110.445 139.745 ;
        RECT 111.035 139.575 111.205 139.745 ;
        RECT 109.320 138.445 110.445 138.615 ;
        RECT 110.615 139.245 110.810 139.575 ;
        RECT 111.035 139.245 111.290 139.575 ;
        RECT 110.615 138.275 110.785 139.245 ;
        RECT 111.460 139.075 111.630 139.745 ;
        RECT 111.805 139.735 113.015 140.485 ;
        RECT 113.275 139.935 113.445 140.315 ;
        RECT 113.625 140.105 113.955 140.485 ;
        RECT 113.275 139.765 113.940 139.935 ;
        RECT 114.135 139.810 114.395 140.315 ;
        RECT 108.755 138.105 110.785 138.275 ;
        RECT 110.955 137.935 111.125 139.075 ;
        RECT 111.295 138.105 111.630 139.075 ;
        RECT 111.805 139.025 112.325 139.565 ;
        RECT 112.495 139.195 113.015 139.735 ;
        RECT 113.205 139.215 113.535 139.585 ;
        RECT 113.770 139.510 113.940 139.765 ;
        RECT 113.770 139.180 114.055 139.510 ;
        RECT 113.770 139.035 113.940 139.180 ;
        RECT 111.805 137.935 113.015 139.025 ;
        RECT 113.275 138.865 113.940 139.035 ;
        RECT 114.225 139.010 114.395 139.810 ;
        RECT 114.565 139.760 114.855 140.485 ;
        RECT 115.065 139.665 115.295 140.485 ;
        RECT 115.465 139.685 115.795 140.315 ;
        RECT 115.045 139.245 115.375 139.495 ;
        RECT 113.275 138.105 113.445 138.865 ;
        RECT 113.625 137.935 113.955 138.695 ;
        RECT 114.125 138.105 114.395 139.010 ;
        RECT 114.565 137.935 114.855 139.100 ;
        RECT 115.545 139.085 115.795 139.685 ;
        RECT 115.965 139.665 116.175 140.485 ;
        RECT 116.780 140.145 117.035 140.305 ;
        RECT 116.695 139.975 117.035 140.145 ;
        RECT 117.215 140.025 117.500 140.485 ;
        RECT 116.780 139.775 117.035 139.975 ;
        RECT 115.065 137.935 115.295 139.075 ;
        RECT 115.465 138.105 115.795 139.085 ;
        RECT 115.965 137.935 116.175 139.075 ;
        RECT 116.780 138.915 116.960 139.775 ;
        RECT 117.680 139.575 117.930 140.225 ;
        RECT 117.130 139.245 117.930 139.575 ;
        RECT 116.780 138.245 117.035 138.915 ;
        RECT 117.215 137.935 117.500 138.735 ;
        RECT 117.680 138.655 117.930 139.245 ;
        RECT 118.130 139.890 118.450 140.220 ;
        RECT 118.630 140.005 119.290 140.485 ;
        RECT 119.490 140.095 120.340 140.265 ;
        RECT 118.130 138.995 118.320 139.890 ;
        RECT 118.640 139.565 119.300 139.835 ;
        RECT 118.970 139.505 119.300 139.565 ;
        RECT 118.490 139.335 118.820 139.395 ;
        RECT 119.490 139.335 119.660 140.095 ;
        RECT 120.900 140.025 121.220 140.485 ;
        RECT 121.420 139.845 121.670 140.275 ;
        RECT 121.960 140.045 122.370 140.485 ;
        RECT 122.540 140.105 123.555 140.305 ;
        RECT 119.830 139.675 121.080 139.845 ;
        RECT 119.830 139.555 120.160 139.675 ;
        RECT 118.490 139.165 120.390 139.335 ;
        RECT 118.130 138.825 120.050 138.995 ;
        RECT 118.130 138.805 118.450 138.825 ;
        RECT 117.680 138.145 118.010 138.655 ;
        RECT 118.280 138.195 118.450 138.805 ;
        RECT 120.220 138.655 120.390 139.165 ;
        RECT 120.560 139.095 120.740 139.505 ;
        RECT 120.910 138.915 121.080 139.675 ;
        RECT 118.620 137.935 118.950 138.625 ;
        RECT 119.180 138.485 120.390 138.655 ;
        RECT 120.560 138.605 121.080 138.915 ;
        RECT 121.250 139.505 121.670 139.845 ;
        RECT 121.960 139.505 122.370 139.835 ;
        RECT 121.250 138.735 121.440 139.505 ;
        RECT 122.540 139.375 122.710 140.105 ;
        RECT 123.855 139.935 124.025 140.265 ;
        RECT 124.195 140.105 124.525 140.485 ;
        RECT 122.880 139.555 123.230 139.925 ;
        RECT 122.540 139.335 122.960 139.375 ;
        RECT 121.610 139.165 122.960 139.335 ;
        RECT 121.610 139.005 121.860 139.165 ;
        RECT 122.370 138.735 122.620 138.995 ;
        RECT 121.250 138.485 122.620 138.735 ;
        RECT 119.180 138.195 119.420 138.485 ;
        RECT 120.220 138.405 120.390 138.485 ;
        RECT 119.620 137.935 120.040 138.315 ;
        RECT 120.220 138.155 120.850 138.405 ;
        RECT 121.320 137.935 121.650 138.315 ;
        RECT 121.820 138.195 121.990 138.485 ;
        RECT 122.790 138.320 122.960 139.165 ;
        RECT 123.410 138.995 123.630 139.865 ;
        RECT 123.855 139.745 124.550 139.935 ;
        RECT 123.130 138.615 123.630 138.995 ;
        RECT 123.800 138.945 124.210 139.565 ;
        RECT 124.380 138.775 124.550 139.745 ;
        RECT 123.855 138.605 124.550 138.775 ;
        RECT 122.170 137.935 122.550 138.315 ;
        RECT 122.790 138.150 123.620 138.320 ;
        RECT 123.855 138.105 124.025 138.605 ;
        RECT 124.195 137.935 124.525 138.435 ;
        RECT 124.740 138.105 124.965 140.225 ;
        RECT 125.135 140.105 125.465 140.485 ;
        RECT 125.635 139.935 125.805 140.225 ;
        RECT 125.140 139.765 125.805 139.935 ;
        RECT 125.140 138.775 125.370 139.765 ;
        RECT 126.525 139.735 127.735 140.485 ;
        RECT 125.540 138.945 125.890 139.595 ;
        RECT 126.525 139.025 127.045 139.565 ;
        RECT 127.215 139.195 127.735 139.735 ;
        RECT 125.140 138.605 125.805 138.775 ;
        RECT 125.135 137.935 125.465 138.435 ;
        RECT 125.635 138.105 125.805 138.605 ;
        RECT 126.525 137.935 127.735 139.025 ;
        RECT 14.660 137.765 127.820 137.935 ;
        RECT 14.745 136.675 15.955 137.765 ;
        RECT 14.745 135.965 15.265 136.505 ;
        RECT 15.435 136.135 15.955 136.675 ;
        RECT 16.125 136.675 17.335 137.765 ;
        RECT 16.125 136.135 16.645 136.675 ;
        RECT 17.545 136.625 17.775 137.765 ;
        RECT 17.945 136.615 18.275 137.595 ;
        RECT 18.445 136.625 18.655 137.765 ;
        RECT 18.925 136.625 19.155 137.765 ;
        RECT 19.325 136.615 19.655 137.595 ;
        RECT 19.825 136.625 20.035 137.765 ;
        RECT 20.265 137.005 20.780 137.415 ;
        RECT 21.015 137.005 21.185 137.765 ;
        RECT 21.355 137.425 23.385 137.595 ;
        RECT 16.815 135.965 17.335 136.505 ;
        RECT 17.525 136.205 17.855 136.455 ;
        RECT 14.745 135.215 15.955 135.965 ;
        RECT 16.125 135.215 17.335 135.965 ;
        RECT 17.545 135.215 17.775 136.035 ;
        RECT 18.025 136.015 18.275 136.615 ;
        RECT 18.905 136.205 19.235 136.455 ;
        RECT 17.945 135.385 18.275 136.015 ;
        RECT 18.445 135.215 18.655 136.035 ;
        RECT 18.925 135.215 19.155 136.035 ;
        RECT 19.405 136.015 19.655 136.615 ;
        RECT 20.265 136.195 20.605 137.005 ;
        RECT 21.355 136.760 21.525 137.425 ;
        RECT 21.920 137.085 23.045 137.255 ;
        RECT 20.775 136.570 21.525 136.760 ;
        RECT 21.695 136.745 22.705 136.915 ;
        RECT 19.325 135.385 19.655 136.015 ;
        RECT 19.825 135.215 20.035 136.035 ;
        RECT 20.265 136.025 21.495 136.195 ;
        RECT 20.540 135.420 20.785 136.025 ;
        RECT 21.005 135.215 21.515 135.750 ;
        RECT 21.695 135.385 21.885 136.745 ;
        RECT 22.055 136.405 22.330 136.545 ;
        RECT 22.055 136.235 22.335 136.405 ;
        RECT 22.055 135.385 22.330 136.235 ;
        RECT 22.535 135.945 22.705 136.745 ;
        RECT 22.875 135.955 23.045 137.085 ;
        RECT 23.215 136.455 23.385 137.425 ;
        RECT 23.555 136.625 23.725 137.765 ;
        RECT 23.895 136.625 24.230 137.595 ;
        RECT 23.215 136.125 23.410 136.455 ;
        RECT 23.635 136.125 23.890 136.455 ;
        RECT 23.635 135.955 23.805 136.125 ;
        RECT 24.060 135.955 24.230 136.625 ;
        RECT 24.405 136.600 24.695 137.765 ;
        RECT 24.865 136.690 25.135 137.595 ;
        RECT 25.305 137.005 25.635 137.765 ;
        RECT 25.815 136.835 25.985 137.595 ;
        RECT 22.875 135.785 23.805 135.955 ;
        RECT 22.875 135.750 23.050 135.785 ;
        RECT 22.520 135.385 23.050 135.750 ;
        RECT 23.475 135.215 23.805 135.615 ;
        RECT 23.975 135.385 24.230 135.955 ;
        RECT 24.405 135.215 24.695 135.940 ;
        RECT 24.865 135.890 25.035 136.690 ;
        RECT 25.320 136.665 25.985 136.835 ;
        RECT 25.320 136.520 25.490 136.665 ;
        RECT 26.745 136.625 26.975 137.765 ;
        RECT 27.145 136.615 27.475 137.595 ;
        RECT 27.645 136.625 27.855 137.765 ;
        RECT 28.085 137.005 28.600 137.415 ;
        RECT 28.835 137.005 29.005 137.765 ;
        RECT 29.175 137.425 31.205 137.595 ;
        RECT 25.205 136.190 25.490 136.520 ;
        RECT 25.320 135.935 25.490 136.190 ;
        RECT 25.725 136.115 26.055 136.485 ;
        RECT 26.725 136.205 27.055 136.455 ;
        RECT 24.865 135.385 25.125 135.890 ;
        RECT 25.320 135.765 25.985 135.935 ;
        RECT 25.305 135.215 25.635 135.595 ;
        RECT 25.815 135.385 25.985 135.765 ;
        RECT 26.745 135.215 26.975 136.035 ;
        RECT 27.225 136.015 27.475 136.615 ;
        RECT 28.085 136.195 28.425 137.005 ;
        RECT 29.175 136.760 29.345 137.425 ;
        RECT 29.740 137.085 30.865 137.255 ;
        RECT 28.595 136.570 29.345 136.760 ;
        RECT 29.515 136.745 30.525 136.915 ;
        RECT 27.145 135.385 27.475 136.015 ;
        RECT 27.645 135.215 27.855 136.035 ;
        RECT 28.085 136.025 29.315 136.195 ;
        RECT 28.360 135.420 28.605 136.025 ;
        RECT 28.825 135.215 29.335 135.750 ;
        RECT 29.515 135.385 29.705 136.745 ;
        RECT 29.875 135.725 30.150 136.545 ;
        RECT 30.355 135.945 30.525 136.745 ;
        RECT 30.695 135.955 30.865 137.085 ;
        RECT 31.035 136.455 31.205 137.425 ;
        RECT 31.375 136.625 31.545 137.765 ;
        RECT 31.715 136.625 32.050 137.595 ;
        RECT 31.035 136.125 31.230 136.455 ;
        RECT 31.455 136.125 31.710 136.455 ;
        RECT 31.455 135.955 31.625 136.125 ;
        RECT 31.880 135.955 32.050 136.625 ;
        RECT 30.695 135.785 31.625 135.955 ;
        RECT 30.695 135.750 30.870 135.785 ;
        RECT 29.875 135.555 30.155 135.725 ;
        RECT 29.875 135.385 30.150 135.555 ;
        RECT 30.340 135.385 30.870 135.750 ;
        RECT 31.295 135.215 31.625 135.615 ;
        RECT 31.795 135.385 32.050 135.955 ;
        RECT 32.600 136.785 32.855 137.455 ;
        RECT 33.035 136.965 33.320 137.765 ;
        RECT 33.500 137.045 33.830 137.555 ;
        RECT 32.600 135.925 32.780 136.785 ;
        RECT 33.500 136.455 33.750 137.045 ;
        RECT 34.100 136.895 34.270 137.505 ;
        RECT 34.440 137.075 34.770 137.765 ;
        RECT 35.000 137.215 35.240 137.505 ;
        RECT 35.440 137.385 35.860 137.765 ;
        RECT 36.040 137.295 36.670 137.545 ;
        RECT 37.140 137.385 37.470 137.765 ;
        RECT 36.040 137.215 36.210 137.295 ;
        RECT 37.640 137.215 37.810 137.505 ;
        RECT 37.990 137.385 38.370 137.765 ;
        RECT 38.610 137.380 39.440 137.550 ;
        RECT 35.000 137.045 36.210 137.215 ;
        RECT 32.950 136.125 33.750 136.455 ;
        RECT 32.600 135.725 32.855 135.925 ;
        RECT 32.515 135.555 32.855 135.725 ;
        RECT 32.600 135.395 32.855 135.555 ;
        RECT 33.035 135.215 33.320 135.675 ;
        RECT 33.500 135.475 33.750 136.125 ;
        RECT 33.950 136.875 34.270 136.895 ;
        RECT 33.950 136.705 35.870 136.875 ;
        RECT 33.950 135.810 34.140 136.705 ;
        RECT 36.040 136.535 36.210 137.045 ;
        RECT 36.380 136.785 36.900 137.095 ;
        RECT 34.310 136.365 36.210 136.535 ;
        RECT 34.310 136.305 34.640 136.365 ;
        RECT 34.790 136.135 35.120 136.195 ;
        RECT 34.460 135.865 35.120 136.135 ;
        RECT 33.950 135.480 34.270 135.810 ;
        RECT 34.450 135.215 35.110 135.695 ;
        RECT 35.310 135.605 35.480 136.365 ;
        RECT 36.380 136.195 36.560 136.605 ;
        RECT 35.650 136.025 35.980 136.145 ;
        RECT 36.730 136.025 36.900 136.785 ;
        RECT 35.650 135.855 36.900 136.025 ;
        RECT 37.070 136.965 38.440 137.215 ;
        RECT 37.070 136.195 37.260 136.965 ;
        RECT 38.190 136.705 38.440 136.965 ;
        RECT 37.430 136.535 37.680 136.695 ;
        RECT 38.610 136.535 38.780 137.380 ;
        RECT 39.675 137.095 39.845 137.595 ;
        RECT 40.015 137.265 40.345 137.765 ;
        RECT 38.950 136.705 39.450 137.085 ;
        RECT 39.675 136.925 40.370 137.095 ;
        RECT 37.430 136.365 38.780 136.535 ;
        RECT 38.360 136.325 38.780 136.365 ;
        RECT 37.070 135.855 37.490 136.195 ;
        RECT 37.780 135.865 38.190 136.195 ;
        RECT 35.310 135.435 36.160 135.605 ;
        RECT 36.720 135.215 37.040 135.675 ;
        RECT 37.240 135.425 37.490 135.855 ;
        RECT 37.780 135.215 38.190 135.655 ;
        RECT 38.360 135.595 38.530 136.325 ;
        RECT 38.700 135.775 39.050 136.145 ;
        RECT 39.230 135.835 39.450 136.705 ;
        RECT 39.620 136.135 40.030 136.755 ;
        RECT 40.200 135.955 40.370 136.925 ;
        RECT 39.675 135.765 40.370 135.955 ;
        RECT 38.360 135.395 39.375 135.595 ;
        RECT 39.675 135.435 39.845 135.765 ;
        RECT 40.015 135.215 40.345 135.595 ;
        RECT 40.560 135.475 40.785 137.595 ;
        RECT 40.955 137.265 41.285 137.765 ;
        RECT 41.455 137.095 41.625 137.595 ;
        RECT 40.960 136.925 41.625 137.095 ;
        RECT 42.805 137.005 43.320 137.415 ;
        RECT 43.555 137.005 43.725 137.765 ;
        RECT 43.895 137.425 45.925 137.595 ;
        RECT 40.960 135.935 41.190 136.925 ;
        RECT 41.360 136.105 41.710 136.755 ;
        RECT 42.805 136.195 43.145 137.005 ;
        RECT 43.895 136.760 44.065 137.425 ;
        RECT 44.460 137.085 45.585 137.255 ;
        RECT 43.315 136.570 44.065 136.760 ;
        RECT 44.235 136.745 45.245 136.915 ;
        RECT 42.805 136.025 44.035 136.195 ;
        RECT 40.960 135.765 41.625 135.935 ;
        RECT 40.955 135.215 41.285 135.595 ;
        RECT 41.455 135.475 41.625 135.765 ;
        RECT 43.080 135.420 43.325 136.025 ;
        RECT 43.545 135.215 44.055 135.750 ;
        RECT 44.235 135.385 44.425 136.745 ;
        RECT 44.595 136.405 44.870 136.545 ;
        RECT 44.595 136.235 44.875 136.405 ;
        RECT 44.595 135.385 44.870 136.235 ;
        RECT 45.075 135.945 45.245 136.745 ;
        RECT 45.415 135.955 45.585 137.085 ;
        RECT 45.755 136.455 45.925 137.425 ;
        RECT 46.095 136.625 46.265 137.765 ;
        RECT 46.435 136.625 46.770 137.595 ;
        RECT 45.755 136.125 45.950 136.455 ;
        RECT 46.175 136.125 46.430 136.455 ;
        RECT 46.175 135.955 46.345 136.125 ;
        RECT 46.600 135.955 46.770 136.625 ;
        RECT 45.415 135.785 46.345 135.955 ;
        RECT 45.415 135.750 45.590 135.785 ;
        RECT 45.060 135.385 45.590 135.750 ;
        RECT 46.015 135.215 46.345 135.615 ;
        RECT 46.515 135.385 46.770 135.955 ;
        RECT 46.945 137.045 47.405 137.595 ;
        RECT 47.595 137.045 47.925 137.765 ;
        RECT 46.945 135.675 47.195 137.045 ;
        RECT 48.125 136.875 48.425 137.425 ;
        RECT 48.595 137.095 48.875 137.765 ;
        RECT 47.485 136.705 48.425 136.875 ;
        RECT 47.485 136.455 47.655 136.705 ;
        RECT 48.795 136.455 49.060 136.815 ;
        RECT 50.165 136.600 50.455 137.765 ;
        RECT 50.625 136.675 54.135 137.765 ;
        RECT 54.680 136.785 54.935 137.455 ;
        RECT 55.115 136.965 55.400 137.765 ;
        RECT 55.580 137.045 55.910 137.555 ;
        RECT 47.365 136.125 47.655 136.455 ;
        RECT 47.825 136.205 48.165 136.455 ;
        RECT 48.385 136.205 49.060 136.455 ;
        RECT 50.625 136.155 52.315 136.675 ;
        RECT 47.485 136.035 47.655 136.125 ;
        RECT 47.485 135.845 48.875 136.035 ;
        RECT 52.485 135.985 54.135 136.505 ;
        RECT 46.945 135.385 47.505 135.675 ;
        RECT 47.675 135.215 47.925 135.675 ;
        RECT 48.545 135.485 48.875 135.845 ;
        RECT 50.165 135.215 50.455 135.940 ;
        RECT 50.625 135.215 54.135 135.985 ;
        RECT 54.680 135.925 54.860 136.785 ;
        RECT 55.580 136.455 55.830 137.045 ;
        RECT 56.180 136.895 56.350 137.505 ;
        RECT 56.520 137.075 56.850 137.765 ;
        RECT 57.080 137.215 57.320 137.505 ;
        RECT 57.520 137.385 57.940 137.765 ;
        RECT 58.120 137.295 58.750 137.545 ;
        RECT 59.220 137.385 59.550 137.765 ;
        RECT 58.120 137.215 58.290 137.295 ;
        RECT 59.720 137.215 59.890 137.505 ;
        RECT 60.070 137.385 60.450 137.765 ;
        RECT 60.690 137.380 61.520 137.550 ;
        RECT 57.080 137.045 58.290 137.215 ;
        RECT 55.030 136.125 55.830 136.455 ;
        RECT 54.680 135.725 54.935 135.925 ;
        RECT 54.595 135.555 54.935 135.725 ;
        RECT 54.680 135.395 54.935 135.555 ;
        RECT 55.115 135.215 55.400 135.675 ;
        RECT 55.580 135.475 55.830 136.125 ;
        RECT 56.030 136.875 56.350 136.895 ;
        RECT 56.030 136.705 57.950 136.875 ;
        RECT 56.030 135.810 56.220 136.705 ;
        RECT 58.120 136.535 58.290 137.045 ;
        RECT 58.460 136.785 58.980 137.095 ;
        RECT 56.390 136.365 58.290 136.535 ;
        RECT 56.390 136.305 56.720 136.365 ;
        RECT 56.870 136.135 57.200 136.195 ;
        RECT 56.540 135.865 57.200 136.135 ;
        RECT 56.030 135.480 56.350 135.810 ;
        RECT 56.530 135.215 57.190 135.695 ;
        RECT 57.390 135.605 57.560 136.365 ;
        RECT 58.460 136.195 58.640 136.605 ;
        RECT 57.730 136.025 58.060 136.145 ;
        RECT 58.810 136.025 58.980 136.785 ;
        RECT 57.730 135.855 58.980 136.025 ;
        RECT 59.150 136.965 60.520 137.215 ;
        RECT 59.150 136.195 59.340 136.965 ;
        RECT 60.270 136.705 60.520 136.965 ;
        RECT 59.510 136.535 59.760 136.695 ;
        RECT 60.690 136.535 60.860 137.380 ;
        RECT 61.755 137.095 61.925 137.595 ;
        RECT 62.095 137.265 62.425 137.765 ;
        RECT 61.030 136.705 61.530 137.085 ;
        RECT 61.755 136.925 62.450 137.095 ;
        RECT 59.510 136.365 60.860 136.535 ;
        RECT 60.440 136.325 60.860 136.365 ;
        RECT 59.150 135.855 59.570 136.195 ;
        RECT 59.860 135.865 60.270 136.195 ;
        RECT 57.390 135.435 58.240 135.605 ;
        RECT 58.800 135.215 59.120 135.675 ;
        RECT 59.320 135.425 59.570 135.855 ;
        RECT 59.860 135.215 60.270 135.655 ;
        RECT 60.440 135.595 60.610 136.325 ;
        RECT 60.780 135.775 61.130 136.145 ;
        RECT 61.310 135.835 61.530 136.705 ;
        RECT 61.700 136.135 62.110 136.755 ;
        RECT 62.280 135.955 62.450 136.925 ;
        RECT 61.755 135.765 62.450 135.955 ;
        RECT 60.440 135.395 61.455 135.595 ;
        RECT 61.755 135.435 61.925 135.765 ;
        RECT 62.095 135.215 62.425 135.595 ;
        RECT 62.640 135.475 62.865 137.595 ;
        RECT 63.035 137.265 63.365 137.765 ;
        RECT 63.535 137.095 63.705 137.595 ;
        RECT 64.890 137.330 70.235 137.765 ;
        RECT 70.410 137.330 75.755 137.765 ;
        RECT 63.040 136.925 63.705 137.095 ;
        RECT 63.040 135.935 63.270 136.925 ;
        RECT 63.440 136.105 63.790 136.755 ;
        RECT 66.480 136.080 66.830 137.330 ;
        RECT 63.040 135.765 63.705 135.935 ;
        RECT 63.035 135.215 63.365 135.595 ;
        RECT 63.535 135.475 63.705 135.765 ;
        RECT 68.310 135.760 68.650 136.590 ;
        RECT 72.000 136.080 72.350 137.330 ;
        RECT 75.925 136.600 76.215 137.765 ;
        RECT 76.390 137.330 81.735 137.765 ;
        RECT 73.830 135.760 74.170 136.590 ;
        RECT 77.980 136.080 78.330 137.330 ;
        RECT 81.905 136.625 82.245 137.595 ;
        RECT 82.415 136.625 82.585 137.765 ;
        RECT 82.855 136.965 83.105 137.765 ;
        RECT 83.750 136.795 84.080 137.595 ;
        RECT 84.380 136.965 84.710 137.765 ;
        RECT 84.880 136.795 85.210 137.595 ;
        RECT 85.590 137.330 90.935 137.765 ;
        RECT 91.110 137.330 96.455 137.765 ;
        RECT 82.775 136.625 85.210 136.795 ;
        RECT 64.890 135.215 70.235 135.760 ;
        RECT 70.410 135.215 75.755 135.760 ;
        RECT 75.925 135.215 76.215 135.940 ;
        RECT 79.810 135.760 80.150 136.590 ;
        RECT 81.905 136.015 82.080 136.625 ;
        RECT 82.775 136.375 82.945 136.625 ;
        RECT 82.250 136.205 82.945 136.375 ;
        RECT 83.120 136.205 83.540 136.405 ;
        RECT 83.710 136.205 84.040 136.405 ;
        RECT 84.210 136.205 84.540 136.405 ;
        RECT 76.390 135.215 81.735 135.760 ;
        RECT 81.905 135.385 82.245 136.015 ;
        RECT 82.415 135.215 82.665 136.015 ;
        RECT 82.855 135.865 84.080 136.035 ;
        RECT 82.855 135.385 83.185 135.865 ;
        RECT 83.355 135.215 83.580 135.675 ;
        RECT 83.750 135.385 84.080 135.865 ;
        RECT 84.710 135.995 84.880 136.625 ;
        RECT 85.065 136.205 85.415 136.455 ;
        RECT 87.180 136.080 87.530 137.330 ;
        RECT 84.710 135.385 85.210 135.995 ;
        RECT 89.010 135.760 89.350 136.590 ;
        RECT 92.700 136.080 93.050 137.330 ;
        RECT 96.625 137.005 97.140 137.415 ;
        RECT 97.375 137.005 97.545 137.765 ;
        RECT 97.715 137.425 99.745 137.595 ;
        RECT 94.530 135.760 94.870 136.590 ;
        RECT 96.625 136.195 96.965 137.005 ;
        RECT 97.715 136.760 97.885 137.425 ;
        RECT 98.280 137.085 99.405 137.255 ;
        RECT 97.135 136.570 97.885 136.760 ;
        RECT 98.055 136.745 99.065 136.915 ;
        RECT 96.625 136.025 97.855 136.195 ;
        RECT 85.590 135.215 90.935 135.760 ;
        RECT 91.110 135.215 96.455 135.760 ;
        RECT 96.900 135.420 97.145 136.025 ;
        RECT 97.365 135.215 97.875 135.750 ;
        RECT 98.055 135.385 98.245 136.745 ;
        RECT 98.415 136.405 98.690 136.545 ;
        RECT 98.415 136.235 98.695 136.405 ;
        RECT 98.415 135.385 98.690 136.235 ;
        RECT 98.895 135.945 99.065 136.745 ;
        RECT 99.235 135.955 99.405 137.085 ;
        RECT 99.575 136.455 99.745 137.425 ;
        RECT 99.915 136.625 100.085 137.765 ;
        RECT 100.255 136.625 100.590 137.595 ;
        RECT 99.575 136.125 99.770 136.455 ;
        RECT 99.995 136.125 100.250 136.455 ;
        RECT 99.995 135.955 100.165 136.125 ;
        RECT 100.420 135.955 100.590 136.625 ;
        RECT 101.685 136.600 101.975 137.765 ;
        RECT 102.145 136.675 104.735 137.765 ;
        RECT 105.280 136.785 105.535 137.455 ;
        RECT 105.715 136.965 106.000 137.765 ;
        RECT 106.180 137.045 106.510 137.555 ;
        RECT 102.145 136.155 103.355 136.675 ;
        RECT 103.525 135.985 104.735 136.505 ;
        RECT 105.280 136.405 105.460 136.785 ;
        RECT 106.180 136.455 106.430 137.045 ;
        RECT 106.780 136.895 106.950 137.505 ;
        RECT 107.120 137.075 107.450 137.765 ;
        RECT 107.680 137.215 107.920 137.505 ;
        RECT 108.120 137.385 108.540 137.765 ;
        RECT 108.720 137.295 109.350 137.545 ;
        RECT 109.820 137.385 110.150 137.765 ;
        RECT 108.720 137.215 108.890 137.295 ;
        RECT 110.320 137.215 110.490 137.505 ;
        RECT 110.670 137.385 111.050 137.765 ;
        RECT 111.290 137.380 112.120 137.550 ;
        RECT 107.680 137.045 108.890 137.215 ;
        RECT 105.195 136.235 105.460 136.405 ;
        RECT 99.235 135.785 100.165 135.955 ;
        RECT 99.235 135.750 99.410 135.785 ;
        RECT 98.880 135.385 99.410 135.750 ;
        RECT 99.835 135.215 100.165 135.615 ;
        RECT 100.335 135.385 100.590 135.955 ;
        RECT 101.685 135.215 101.975 135.940 ;
        RECT 102.145 135.215 104.735 135.985 ;
        RECT 105.280 135.925 105.460 136.235 ;
        RECT 105.630 136.125 106.430 136.455 ;
        RECT 105.280 135.395 105.535 135.925 ;
        RECT 105.715 135.215 106.000 135.675 ;
        RECT 106.180 135.475 106.430 136.125 ;
        RECT 106.630 136.875 106.950 136.895 ;
        RECT 106.630 136.705 108.550 136.875 ;
        RECT 106.630 135.810 106.820 136.705 ;
        RECT 108.720 136.535 108.890 137.045 ;
        RECT 109.060 136.785 109.580 137.095 ;
        RECT 106.990 136.365 108.890 136.535 ;
        RECT 106.990 136.305 107.320 136.365 ;
        RECT 107.470 136.135 107.800 136.195 ;
        RECT 107.140 135.865 107.800 136.135 ;
        RECT 106.630 135.480 106.950 135.810 ;
        RECT 107.130 135.215 107.790 135.695 ;
        RECT 107.990 135.605 108.160 136.365 ;
        RECT 109.060 136.195 109.240 136.605 ;
        RECT 108.330 136.025 108.660 136.145 ;
        RECT 109.410 136.025 109.580 136.785 ;
        RECT 108.330 135.855 109.580 136.025 ;
        RECT 109.750 136.965 111.120 137.215 ;
        RECT 109.750 136.195 109.940 136.965 ;
        RECT 110.870 136.705 111.120 136.965 ;
        RECT 110.110 136.535 110.360 136.695 ;
        RECT 111.290 136.535 111.460 137.380 ;
        RECT 112.355 137.095 112.525 137.595 ;
        RECT 112.695 137.265 113.025 137.765 ;
        RECT 111.630 136.705 112.130 137.085 ;
        RECT 112.355 136.925 113.050 137.095 ;
        RECT 110.110 136.365 111.460 136.535 ;
        RECT 111.040 136.325 111.460 136.365 ;
        RECT 109.750 135.855 110.170 136.195 ;
        RECT 110.460 135.865 110.870 136.195 ;
        RECT 107.990 135.435 108.840 135.605 ;
        RECT 109.400 135.215 109.720 135.675 ;
        RECT 109.920 135.425 110.170 135.855 ;
        RECT 110.460 135.215 110.870 135.655 ;
        RECT 111.040 135.595 111.210 136.325 ;
        RECT 111.380 135.775 111.730 136.145 ;
        RECT 111.910 135.835 112.130 136.705 ;
        RECT 112.300 136.135 112.710 136.755 ;
        RECT 112.880 135.955 113.050 136.925 ;
        RECT 112.355 135.765 113.050 135.955 ;
        RECT 111.040 135.395 112.055 135.595 ;
        RECT 112.355 135.435 112.525 135.765 ;
        RECT 112.695 135.215 113.025 135.595 ;
        RECT 113.240 135.475 113.465 137.595 ;
        RECT 113.635 137.265 113.965 137.765 ;
        RECT 114.135 137.095 114.305 137.595 ;
        RECT 113.640 136.925 114.305 137.095 ;
        RECT 113.640 135.935 113.870 136.925 ;
        RECT 114.040 136.105 114.390 136.755 ;
        RECT 114.565 136.675 115.775 137.765 ;
        RECT 116.320 137.425 116.575 137.455 ;
        RECT 116.235 137.255 116.575 137.425 ;
        RECT 116.320 136.785 116.575 137.255 ;
        RECT 116.755 136.965 117.040 137.765 ;
        RECT 117.220 137.045 117.550 137.555 ;
        RECT 114.565 136.135 115.085 136.675 ;
        RECT 115.255 135.965 115.775 136.505 ;
        RECT 113.640 135.765 114.305 135.935 ;
        RECT 113.635 135.215 113.965 135.595 ;
        RECT 114.135 135.475 114.305 135.765 ;
        RECT 114.565 135.215 115.775 135.965 ;
        RECT 116.320 135.925 116.500 136.785 ;
        RECT 117.220 136.455 117.470 137.045 ;
        RECT 117.820 136.895 117.990 137.505 ;
        RECT 118.160 137.075 118.490 137.765 ;
        RECT 118.720 137.215 118.960 137.505 ;
        RECT 119.160 137.385 119.580 137.765 ;
        RECT 119.760 137.295 120.390 137.545 ;
        RECT 120.860 137.385 121.190 137.765 ;
        RECT 119.760 137.215 119.930 137.295 ;
        RECT 121.360 137.215 121.530 137.505 ;
        RECT 121.710 137.385 122.090 137.765 ;
        RECT 122.330 137.380 123.160 137.550 ;
        RECT 118.720 137.045 119.930 137.215 ;
        RECT 116.670 136.125 117.470 136.455 ;
        RECT 116.320 135.395 116.575 135.925 ;
        RECT 116.755 135.215 117.040 135.675 ;
        RECT 117.220 135.475 117.470 136.125 ;
        RECT 117.670 136.875 117.990 136.895 ;
        RECT 117.670 136.705 119.590 136.875 ;
        RECT 117.670 135.810 117.860 136.705 ;
        RECT 119.760 136.535 119.930 137.045 ;
        RECT 120.100 136.785 120.620 137.095 ;
        RECT 118.030 136.365 119.930 136.535 ;
        RECT 118.030 136.305 118.360 136.365 ;
        RECT 118.510 136.135 118.840 136.195 ;
        RECT 118.180 135.865 118.840 136.135 ;
        RECT 117.670 135.480 117.990 135.810 ;
        RECT 118.170 135.215 118.830 135.695 ;
        RECT 119.030 135.605 119.200 136.365 ;
        RECT 120.100 136.195 120.280 136.605 ;
        RECT 119.370 136.025 119.700 136.145 ;
        RECT 120.450 136.025 120.620 136.785 ;
        RECT 119.370 135.855 120.620 136.025 ;
        RECT 120.790 136.965 122.160 137.215 ;
        RECT 120.790 136.195 120.980 136.965 ;
        RECT 121.910 136.705 122.160 136.965 ;
        RECT 121.150 136.535 121.400 136.695 ;
        RECT 122.330 136.535 122.500 137.380 ;
        RECT 123.395 137.095 123.565 137.595 ;
        RECT 123.735 137.265 124.065 137.765 ;
        RECT 122.670 136.705 123.170 137.085 ;
        RECT 123.395 136.925 124.090 137.095 ;
        RECT 121.150 136.365 122.500 136.535 ;
        RECT 122.080 136.325 122.500 136.365 ;
        RECT 120.790 135.855 121.210 136.195 ;
        RECT 121.500 135.865 121.910 136.195 ;
        RECT 119.030 135.435 119.880 135.605 ;
        RECT 120.440 135.215 120.760 135.675 ;
        RECT 120.960 135.425 121.210 135.855 ;
        RECT 121.500 135.215 121.910 135.655 ;
        RECT 122.080 135.595 122.250 136.325 ;
        RECT 122.420 135.775 122.770 136.145 ;
        RECT 122.950 135.835 123.170 136.705 ;
        RECT 123.340 136.135 123.750 136.755 ;
        RECT 123.920 135.955 124.090 136.925 ;
        RECT 123.395 135.765 124.090 135.955 ;
        RECT 122.080 135.395 123.095 135.595 ;
        RECT 123.395 135.435 123.565 135.765 ;
        RECT 123.735 135.215 124.065 135.595 ;
        RECT 124.280 135.475 124.505 137.595 ;
        RECT 124.675 137.265 125.005 137.765 ;
        RECT 125.175 137.095 125.345 137.595 ;
        RECT 124.680 136.925 125.345 137.095 ;
        RECT 124.680 135.935 124.910 136.925 ;
        RECT 125.080 136.105 125.430 136.755 ;
        RECT 126.525 136.675 127.735 137.765 ;
        RECT 126.525 136.135 127.045 136.675 ;
        RECT 127.215 135.965 127.735 136.505 ;
        RECT 124.680 135.765 125.345 135.935 ;
        RECT 124.675 135.215 125.005 135.595 ;
        RECT 125.175 135.475 125.345 135.765 ;
        RECT 126.525 135.215 127.735 135.965 ;
        RECT 14.660 135.045 127.820 135.215 ;
        RECT 14.745 134.295 15.955 135.045 ;
        RECT 14.745 133.755 15.265 134.295 ;
        RECT 16.585 134.275 18.255 135.045 ;
        RECT 18.515 134.495 18.685 134.875 ;
        RECT 18.865 134.665 19.195 135.045 ;
        RECT 18.515 134.325 19.180 134.495 ;
        RECT 19.375 134.370 19.635 134.875 ;
        RECT 15.435 133.585 15.955 134.125 ;
        RECT 14.745 132.495 15.955 133.585 ;
        RECT 16.585 133.585 17.335 134.105 ;
        RECT 17.505 133.755 18.255 134.275 ;
        RECT 18.445 133.775 18.775 134.145 ;
        RECT 19.010 134.070 19.180 134.325 ;
        RECT 19.010 133.740 19.295 134.070 ;
        RECT 19.010 133.595 19.180 133.740 ;
        RECT 16.585 132.495 18.255 133.585 ;
        RECT 18.515 133.425 19.180 133.595 ;
        RECT 19.465 133.570 19.635 134.370 ;
        RECT 18.515 132.665 18.685 133.425 ;
        RECT 18.865 132.495 19.195 133.255 ;
        RECT 19.365 132.665 19.635 133.570 ;
        RECT 19.810 134.305 20.065 134.875 ;
        RECT 20.235 134.645 20.565 135.045 ;
        RECT 20.990 134.510 21.520 134.875 ;
        RECT 21.710 134.705 21.985 134.875 ;
        RECT 21.705 134.535 21.985 134.705 ;
        RECT 20.990 134.475 21.165 134.510 ;
        RECT 20.235 134.305 21.165 134.475 ;
        RECT 19.810 133.635 19.980 134.305 ;
        RECT 20.235 134.135 20.405 134.305 ;
        RECT 20.150 133.805 20.405 134.135 ;
        RECT 20.630 133.805 20.825 134.135 ;
        RECT 19.810 132.665 20.145 133.635 ;
        RECT 20.315 132.495 20.485 133.635 ;
        RECT 20.655 132.835 20.825 133.805 ;
        RECT 20.995 133.175 21.165 134.305 ;
        RECT 21.335 133.515 21.505 134.315 ;
        RECT 21.710 133.715 21.985 134.535 ;
        RECT 22.155 133.515 22.345 134.875 ;
        RECT 22.525 134.510 23.035 135.045 ;
        RECT 23.255 134.235 23.500 134.840 ;
        RECT 24.320 134.705 24.575 134.865 ;
        RECT 24.235 134.535 24.575 134.705 ;
        RECT 24.755 134.585 25.040 135.045 ;
        RECT 24.320 134.335 24.575 134.535 ;
        RECT 22.545 134.065 23.775 134.235 ;
        RECT 21.335 133.345 22.345 133.515 ;
        RECT 22.515 133.500 23.265 133.690 ;
        RECT 20.995 133.005 22.120 133.175 ;
        RECT 22.515 132.835 22.685 133.500 ;
        RECT 23.435 133.255 23.775 134.065 ;
        RECT 20.655 132.665 22.685 132.835 ;
        RECT 22.855 132.495 23.025 133.255 ;
        RECT 23.260 132.845 23.775 133.255 ;
        RECT 24.320 133.475 24.500 134.335 ;
        RECT 25.220 134.135 25.470 134.785 ;
        RECT 24.670 133.805 25.470 134.135 ;
        RECT 24.320 132.805 24.575 133.475 ;
        RECT 24.755 132.495 25.040 133.295 ;
        RECT 25.220 133.215 25.470 133.805 ;
        RECT 25.670 134.450 25.990 134.780 ;
        RECT 26.170 134.565 26.830 135.045 ;
        RECT 27.030 134.655 27.880 134.825 ;
        RECT 25.670 133.555 25.860 134.450 ;
        RECT 26.180 134.125 26.840 134.395 ;
        RECT 26.510 134.065 26.840 134.125 ;
        RECT 26.030 133.895 26.360 133.955 ;
        RECT 27.030 133.895 27.200 134.655 ;
        RECT 28.440 134.585 28.760 135.045 ;
        RECT 28.960 134.405 29.210 134.835 ;
        RECT 29.500 134.605 29.910 135.045 ;
        RECT 30.080 134.665 31.095 134.865 ;
        RECT 27.370 134.235 28.620 134.405 ;
        RECT 27.370 134.115 27.700 134.235 ;
        RECT 26.030 133.725 27.930 133.895 ;
        RECT 25.670 133.385 27.590 133.555 ;
        RECT 25.670 133.365 25.990 133.385 ;
        RECT 25.220 132.705 25.550 133.215 ;
        RECT 25.820 132.755 25.990 133.365 ;
        RECT 27.760 133.215 27.930 133.725 ;
        RECT 28.100 133.655 28.280 134.065 ;
        RECT 28.450 133.475 28.620 134.235 ;
        RECT 26.160 132.495 26.490 133.185 ;
        RECT 26.720 133.045 27.930 133.215 ;
        RECT 28.100 133.165 28.620 133.475 ;
        RECT 28.790 134.065 29.210 134.405 ;
        RECT 29.500 134.065 29.910 134.395 ;
        RECT 28.790 133.295 28.980 134.065 ;
        RECT 30.080 133.935 30.250 134.665 ;
        RECT 31.395 134.495 31.565 134.825 ;
        RECT 31.735 134.665 32.065 135.045 ;
        RECT 30.420 134.115 30.770 134.485 ;
        RECT 30.080 133.895 30.500 133.935 ;
        RECT 29.150 133.725 30.500 133.895 ;
        RECT 29.150 133.565 29.400 133.725 ;
        RECT 29.910 133.295 30.160 133.555 ;
        RECT 28.790 133.045 30.160 133.295 ;
        RECT 26.720 132.755 26.960 133.045 ;
        RECT 27.760 132.965 27.930 133.045 ;
        RECT 27.160 132.495 27.580 132.875 ;
        RECT 27.760 132.715 28.390 132.965 ;
        RECT 28.860 132.495 29.190 132.875 ;
        RECT 29.360 132.755 29.530 133.045 ;
        RECT 30.330 132.880 30.500 133.725 ;
        RECT 30.950 133.555 31.170 134.425 ;
        RECT 31.395 134.305 32.090 134.495 ;
        RECT 30.670 133.175 31.170 133.555 ;
        RECT 31.340 133.505 31.750 134.125 ;
        RECT 31.920 133.335 32.090 134.305 ;
        RECT 31.395 133.165 32.090 133.335 ;
        RECT 29.710 132.495 30.090 132.875 ;
        RECT 30.330 132.710 31.160 132.880 ;
        RECT 31.395 132.665 31.565 133.165 ;
        RECT 31.735 132.495 32.065 132.995 ;
        RECT 32.280 132.665 32.505 134.785 ;
        RECT 32.675 134.665 33.005 135.045 ;
        RECT 33.175 134.495 33.345 134.785 ;
        RECT 32.680 134.325 33.345 134.495 ;
        RECT 32.680 133.335 32.910 134.325 ;
        RECT 33.605 134.275 35.275 135.045 ;
        RECT 33.080 133.505 33.430 134.155 ;
        RECT 33.605 133.585 34.355 134.105 ;
        RECT 34.525 133.755 35.275 134.275 ;
        RECT 35.485 134.225 35.715 135.045 ;
        RECT 35.885 134.245 36.215 134.875 ;
        RECT 35.465 133.805 35.795 134.055 ;
        RECT 35.965 133.645 36.215 134.245 ;
        RECT 36.385 134.225 36.595 135.045 ;
        RECT 37.285 134.320 37.575 135.045 ;
        RECT 38.295 134.495 38.465 134.875 ;
        RECT 38.645 134.665 38.975 135.045 ;
        RECT 38.295 134.325 38.960 134.495 ;
        RECT 39.155 134.370 39.415 134.875 ;
        RECT 38.225 133.775 38.555 134.145 ;
        RECT 38.790 134.070 38.960 134.325 ;
        RECT 38.790 133.740 39.075 134.070 ;
        RECT 32.680 133.165 33.345 133.335 ;
        RECT 32.675 132.495 33.005 132.995 ;
        RECT 33.175 132.665 33.345 133.165 ;
        RECT 33.605 132.495 35.275 133.585 ;
        RECT 35.485 132.495 35.715 133.635 ;
        RECT 35.885 132.665 36.215 133.645 ;
        RECT 36.385 132.495 36.595 133.635 ;
        RECT 37.285 132.495 37.575 133.660 ;
        RECT 38.790 133.595 38.960 133.740 ;
        RECT 38.295 133.425 38.960 133.595 ;
        RECT 39.245 133.570 39.415 134.370 ;
        RECT 38.295 132.665 38.465 133.425 ;
        RECT 38.645 132.495 38.975 133.255 ;
        RECT 39.145 132.665 39.415 133.570 ;
        RECT 39.960 134.335 40.215 134.865 ;
        RECT 40.395 134.585 40.680 135.045 ;
        RECT 39.960 133.475 40.140 134.335 ;
        RECT 40.860 134.135 41.110 134.785 ;
        RECT 40.310 133.805 41.110 134.135 ;
        RECT 39.960 133.005 40.215 133.475 ;
        RECT 39.875 132.835 40.215 133.005 ;
        RECT 39.960 132.805 40.215 132.835 ;
        RECT 40.395 132.495 40.680 133.295 ;
        RECT 40.860 133.215 41.110 133.805 ;
        RECT 41.310 134.450 41.630 134.780 ;
        RECT 41.810 134.565 42.470 135.045 ;
        RECT 42.670 134.655 43.520 134.825 ;
        RECT 41.310 133.555 41.500 134.450 ;
        RECT 41.820 134.125 42.480 134.395 ;
        RECT 42.150 134.065 42.480 134.125 ;
        RECT 41.670 133.895 42.000 133.955 ;
        RECT 42.670 133.895 42.840 134.655 ;
        RECT 44.080 134.585 44.400 135.045 ;
        RECT 44.600 134.405 44.850 134.835 ;
        RECT 45.140 134.605 45.550 135.045 ;
        RECT 45.720 134.665 46.735 134.865 ;
        RECT 43.010 134.235 44.260 134.405 ;
        RECT 43.010 134.115 43.340 134.235 ;
        RECT 41.670 133.725 43.570 133.895 ;
        RECT 41.310 133.385 43.230 133.555 ;
        RECT 41.310 133.365 41.630 133.385 ;
        RECT 40.860 132.705 41.190 133.215 ;
        RECT 41.460 132.755 41.630 133.365 ;
        RECT 43.400 133.215 43.570 133.725 ;
        RECT 43.740 133.655 43.920 134.065 ;
        RECT 44.090 133.475 44.260 134.235 ;
        RECT 41.800 132.495 42.130 133.185 ;
        RECT 42.360 133.045 43.570 133.215 ;
        RECT 43.740 133.165 44.260 133.475 ;
        RECT 44.430 134.065 44.850 134.405 ;
        RECT 45.140 134.065 45.550 134.395 ;
        RECT 44.430 133.295 44.620 134.065 ;
        RECT 45.720 133.935 45.890 134.665 ;
        RECT 47.035 134.495 47.205 134.825 ;
        RECT 47.375 134.665 47.705 135.045 ;
        RECT 46.060 134.115 46.410 134.485 ;
        RECT 45.720 133.895 46.140 133.935 ;
        RECT 44.790 133.725 46.140 133.895 ;
        RECT 44.790 133.565 45.040 133.725 ;
        RECT 45.550 133.295 45.800 133.555 ;
        RECT 44.430 133.045 45.800 133.295 ;
        RECT 42.360 132.755 42.600 133.045 ;
        RECT 43.400 132.965 43.570 133.045 ;
        RECT 42.800 132.495 43.220 132.875 ;
        RECT 43.400 132.715 44.030 132.965 ;
        RECT 44.500 132.495 44.830 132.875 ;
        RECT 45.000 132.755 45.170 133.045 ;
        RECT 45.970 132.880 46.140 133.725 ;
        RECT 46.590 133.555 46.810 134.425 ;
        RECT 47.035 134.305 47.730 134.495 ;
        RECT 46.310 133.175 46.810 133.555 ;
        RECT 46.980 133.505 47.390 134.125 ;
        RECT 47.560 133.335 47.730 134.305 ;
        RECT 47.035 133.165 47.730 133.335 ;
        RECT 45.350 132.495 45.730 132.875 ;
        RECT 45.970 132.710 46.800 132.880 ;
        RECT 47.035 132.665 47.205 133.165 ;
        RECT 47.375 132.495 47.705 132.995 ;
        RECT 47.920 132.665 48.145 134.785 ;
        RECT 48.315 134.665 48.645 135.045 ;
        RECT 48.815 134.495 48.985 134.785 ;
        RECT 48.320 134.325 48.985 134.495 ;
        RECT 48.320 133.335 48.550 134.325 ;
        RECT 49.245 134.275 51.835 135.045 ;
        RECT 52.010 134.500 57.355 135.045 ;
        RECT 48.720 133.505 49.070 134.155 ;
        RECT 49.245 133.585 50.455 134.105 ;
        RECT 50.625 133.755 51.835 134.275 ;
        RECT 48.320 133.165 48.985 133.335 ;
        RECT 48.315 132.495 48.645 132.995 ;
        RECT 48.815 132.665 48.985 133.165 ;
        RECT 49.245 132.495 51.835 133.585 ;
        RECT 53.600 132.930 53.950 134.180 ;
        RECT 55.430 133.670 55.770 134.500 ;
        RECT 57.565 134.225 57.795 135.045 ;
        RECT 57.965 134.245 58.295 134.875 ;
        RECT 57.545 133.805 57.875 134.055 ;
        RECT 58.045 133.645 58.295 134.245 ;
        RECT 58.465 134.225 58.675 135.045 ;
        RECT 59.365 134.275 62.875 135.045 ;
        RECT 63.045 134.320 63.335 135.045 ;
        RECT 63.505 134.275 66.095 135.045 ;
        RECT 66.270 134.645 66.605 135.045 ;
        RECT 66.775 134.475 66.980 134.875 ;
        RECT 67.190 134.565 67.465 135.045 ;
        RECT 67.675 134.545 67.935 134.875 ;
        RECT 52.010 132.495 57.355 132.930 ;
        RECT 57.565 132.495 57.795 133.635 ;
        RECT 57.965 132.665 58.295 133.645 ;
        RECT 58.465 132.495 58.675 133.635 ;
        RECT 59.365 133.585 61.055 134.105 ;
        RECT 61.225 133.755 62.875 134.275 ;
        RECT 59.365 132.495 62.875 133.585 ;
        RECT 63.045 132.495 63.335 133.660 ;
        RECT 63.505 133.585 64.715 134.105 ;
        RECT 64.885 133.755 66.095 134.275 ;
        RECT 66.295 134.305 66.980 134.475 ;
        RECT 63.505 132.495 66.095 133.585 ;
        RECT 66.295 133.275 66.635 134.305 ;
        RECT 66.805 133.635 67.055 134.135 ;
        RECT 67.235 133.805 67.595 134.385 ;
        RECT 67.765 133.635 67.935 134.545 ;
        RECT 68.380 134.235 68.625 134.840 ;
        RECT 68.845 134.510 69.355 135.045 ;
        RECT 66.805 133.465 67.935 133.635 ;
        RECT 66.295 133.100 66.960 133.275 ;
        RECT 66.270 132.495 66.605 132.920 ;
        RECT 66.775 132.695 66.960 133.100 ;
        RECT 67.165 132.495 67.495 133.275 ;
        RECT 67.665 132.695 67.935 133.465 ;
        RECT 68.105 134.065 69.335 134.235 ;
        RECT 68.105 133.255 68.445 134.065 ;
        RECT 68.615 133.500 69.365 133.690 ;
        RECT 68.105 132.845 68.620 133.255 ;
        RECT 68.855 132.495 69.025 133.255 ;
        RECT 69.195 132.835 69.365 133.500 ;
        RECT 69.535 133.515 69.725 134.875 ;
        RECT 69.895 134.025 70.170 134.875 ;
        RECT 70.360 134.510 70.890 134.875 ;
        RECT 71.315 134.645 71.645 135.045 ;
        RECT 70.715 134.475 70.890 134.510 ;
        RECT 69.895 133.855 70.175 134.025 ;
        RECT 69.895 133.715 70.170 133.855 ;
        RECT 70.375 133.515 70.545 134.315 ;
        RECT 69.535 133.345 70.545 133.515 ;
        RECT 70.715 134.305 71.645 134.475 ;
        RECT 71.815 134.305 72.070 134.875 ;
        RECT 70.715 133.175 70.885 134.305 ;
        RECT 71.475 134.135 71.645 134.305 ;
        RECT 69.760 133.005 70.885 133.175 ;
        RECT 71.055 133.805 71.250 134.135 ;
        RECT 71.475 133.805 71.730 134.135 ;
        RECT 71.055 132.835 71.225 133.805 ;
        RECT 71.900 133.635 72.070 134.305 ;
        RECT 69.195 132.665 71.225 132.835 ;
        RECT 71.395 132.495 71.565 133.635 ;
        RECT 71.735 132.665 72.070 133.635 ;
        RECT 72.245 134.545 72.505 134.875 ;
        RECT 72.715 134.565 72.990 135.045 ;
        RECT 72.245 133.635 72.415 134.545 ;
        RECT 73.200 134.475 73.405 134.875 ;
        RECT 73.575 134.645 73.910 135.045 ;
        RECT 72.585 133.805 72.945 134.385 ;
        RECT 73.200 134.305 73.885 134.475 ;
        RECT 73.125 133.635 73.375 134.135 ;
        RECT 72.245 133.465 73.375 133.635 ;
        RECT 72.245 132.695 72.515 133.465 ;
        RECT 73.545 133.275 73.885 134.305 ;
        RECT 74.545 134.275 78.055 135.045 ;
        RECT 72.685 132.495 73.015 133.275 ;
        RECT 73.220 133.100 73.885 133.275 ;
        RECT 74.545 133.585 76.235 134.105 ;
        RECT 76.405 133.755 78.055 134.275 ;
        RECT 78.225 134.370 78.495 134.715 ;
        RECT 78.685 134.645 79.065 135.045 ;
        RECT 79.235 134.475 79.405 134.825 ;
        RECT 79.575 134.645 79.905 135.045 ;
        RECT 80.105 134.475 80.275 134.825 ;
        RECT 80.475 134.545 80.805 135.045 ;
        RECT 78.225 133.635 78.395 134.370 ;
        RECT 78.665 134.305 80.275 134.475 ;
        RECT 78.665 134.135 78.835 134.305 ;
        RECT 78.565 133.805 78.835 134.135 ;
        RECT 79.005 133.805 79.410 134.135 ;
        RECT 78.665 133.635 78.835 133.805 ;
        RECT 79.580 133.685 80.290 134.135 ;
        RECT 80.460 133.805 80.810 134.375 ;
        RECT 80.985 134.245 81.325 134.875 ;
        RECT 81.495 134.245 81.745 135.045 ;
        RECT 81.935 134.395 82.265 134.875 ;
        RECT 82.435 134.585 82.660 135.045 ;
        RECT 82.830 134.395 83.160 134.875 ;
        RECT 73.220 132.695 73.405 133.100 ;
        RECT 73.575 132.495 73.910 132.920 ;
        RECT 74.545 132.495 78.055 133.585 ;
        RECT 78.225 132.665 78.495 133.635 ;
        RECT 78.665 133.465 79.390 133.635 ;
        RECT 79.580 133.515 80.295 133.685 ;
        RECT 80.985 133.635 81.160 134.245 ;
        RECT 81.935 134.225 83.160 134.395 ;
        RECT 83.790 134.265 84.290 134.875 ;
        RECT 81.330 133.885 82.025 134.055 ;
        RECT 81.855 133.635 82.025 133.885 ;
        RECT 82.200 133.855 82.620 134.055 ;
        RECT 82.790 133.855 83.120 134.055 ;
        RECT 83.290 133.855 83.620 134.055 ;
        RECT 83.790 133.635 83.960 134.265 ;
        RECT 84.940 134.235 85.185 134.840 ;
        RECT 85.405 134.510 85.915 135.045 ;
        RECT 84.665 134.065 85.895 134.235 ;
        RECT 84.145 133.805 84.495 134.055 ;
        RECT 79.220 133.345 79.390 133.465 ;
        RECT 80.490 133.345 80.810 133.635 ;
        RECT 78.705 132.495 78.985 133.295 ;
        RECT 79.220 133.175 80.810 133.345 ;
        RECT 79.155 132.715 80.810 133.005 ;
        RECT 80.985 132.665 81.325 133.635 ;
        RECT 81.495 132.495 81.665 133.635 ;
        RECT 81.855 133.465 84.290 133.635 ;
        RECT 81.935 132.495 82.185 133.295 ;
        RECT 82.830 132.665 83.160 133.465 ;
        RECT 83.460 132.495 83.790 133.295 ;
        RECT 83.960 132.665 84.290 133.465 ;
        RECT 84.665 133.255 85.005 134.065 ;
        RECT 85.175 133.500 85.925 133.690 ;
        RECT 84.665 132.845 85.180 133.255 ;
        RECT 85.415 132.495 85.585 133.255 ;
        RECT 85.755 132.835 85.925 133.500 ;
        RECT 86.095 133.515 86.285 134.875 ;
        RECT 86.455 134.365 86.730 134.875 ;
        RECT 86.920 134.510 87.450 134.875 ;
        RECT 87.875 134.645 88.205 135.045 ;
        RECT 87.275 134.475 87.450 134.510 ;
        RECT 86.455 134.195 86.735 134.365 ;
        RECT 86.455 133.715 86.730 134.195 ;
        RECT 86.935 133.515 87.105 134.315 ;
        RECT 86.095 133.345 87.105 133.515 ;
        RECT 87.275 134.305 88.205 134.475 ;
        RECT 88.375 134.305 88.630 134.875 ;
        RECT 88.805 134.320 89.095 135.045 ;
        RECT 87.275 133.175 87.445 134.305 ;
        RECT 88.035 134.135 88.205 134.305 ;
        RECT 86.320 133.005 87.445 133.175 ;
        RECT 87.615 133.805 87.810 134.135 ;
        RECT 88.035 133.805 88.290 134.135 ;
        RECT 87.615 132.835 87.785 133.805 ;
        RECT 88.460 133.635 88.630 134.305 ;
        RECT 89.325 134.225 89.535 135.045 ;
        RECT 89.705 134.245 90.035 134.875 ;
        RECT 85.755 132.665 87.785 132.835 ;
        RECT 87.955 132.495 88.125 133.635 ;
        RECT 88.295 132.665 88.630 133.635 ;
        RECT 88.805 132.495 89.095 133.660 ;
        RECT 89.705 133.645 89.955 134.245 ;
        RECT 90.205 134.225 90.435 135.045 ;
        RECT 90.735 134.495 90.905 134.875 ;
        RECT 91.085 134.665 91.415 135.045 ;
        RECT 90.735 134.325 91.400 134.495 ;
        RECT 91.595 134.370 91.855 134.875 ;
        RECT 90.125 133.805 90.455 134.055 ;
        RECT 90.665 133.775 90.995 134.145 ;
        RECT 91.230 134.070 91.400 134.325 ;
        RECT 91.230 133.740 91.515 134.070 ;
        RECT 89.325 132.495 89.535 133.635 ;
        RECT 89.705 132.665 90.035 133.645 ;
        RECT 90.205 132.495 90.435 133.635 ;
        RECT 91.230 133.595 91.400 133.740 ;
        RECT 90.735 133.425 91.400 133.595 ;
        RECT 91.685 133.570 91.855 134.370 ;
        RECT 92.860 134.335 93.115 134.865 ;
        RECT 93.295 134.585 93.580 135.045 ;
        RECT 92.860 133.685 93.040 134.335 ;
        RECT 93.760 134.135 94.010 134.785 ;
        RECT 93.210 133.805 94.010 134.135 ;
        RECT 90.735 132.665 90.905 133.425 ;
        RECT 91.085 132.495 91.415 133.255 ;
        RECT 91.585 132.665 91.855 133.570 ;
        RECT 92.775 133.515 93.040 133.685 ;
        RECT 92.860 133.475 93.040 133.515 ;
        RECT 92.860 132.805 93.115 133.475 ;
        RECT 93.295 132.495 93.580 133.295 ;
        RECT 93.760 133.215 94.010 133.805 ;
        RECT 94.210 134.450 94.530 134.780 ;
        RECT 94.710 134.565 95.370 135.045 ;
        RECT 95.570 134.655 96.420 134.825 ;
        RECT 94.210 133.555 94.400 134.450 ;
        RECT 94.720 134.125 95.380 134.395 ;
        RECT 95.050 134.065 95.380 134.125 ;
        RECT 94.570 133.895 94.900 133.955 ;
        RECT 95.570 133.895 95.740 134.655 ;
        RECT 96.980 134.585 97.300 135.045 ;
        RECT 97.500 134.405 97.750 134.835 ;
        RECT 98.040 134.605 98.450 135.045 ;
        RECT 98.620 134.665 99.635 134.865 ;
        RECT 95.910 134.235 97.160 134.405 ;
        RECT 95.910 134.115 96.240 134.235 ;
        RECT 94.570 133.725 96.470 133.895 ;
        RECT 94.210 133.385 96.130 133.555 ;
        RECT 94.210 133.365 94.530 133.385 ;
        RECT 93.760 132.705 94.090 133.215 ;
        RECT 94.360 132.755 94.530 133.365 ;
        RECT 96.300 133.215 96.470 133.725 ;
        RECT 96.640 133.655 96.820 134.065 ;
        RECT 96.990 133.475 97.160 134.235 ;
        RECT 94.700 132.495 95.030 133.185 ;
        RECT 95.260 133.045 96.470 133.215 ;
        RECT 96.640 133.165 97.160 133.475 ;
        RECT 97.330 134.065 97.750 134.405 ;
        RECT 98.040 134.065 98.450 134.395 ;
        RECT 97.330 133.295 97.520 134.065 ;
        RECT 98.620 133.935 98.790 134.665 ;
        RECT 99.935 134.495 100.105 134.825 ;
        RECT 100.275 134.665 100.605 135.045 ;
        RECT 98.960 134.115 99.310 134.485 ;
        RECT 98.620 133.895 99.040 133.935 ;
        RECT 97.690 133.725 99.040 133.895 ;
        RECT 97.690 133.565 97.940 133.725 ;
        RECT 98.450 133.295 98.700 133.555 ;
        RECT 97.330 133.045 98.700 133.295 ;
        RECT 95.260 132.755 95.500 133.045 ;
        RECT 96.300 132.965 96.470 133.045 ;
        RECT 95.700 132.495 96.120 132.875 ;
        RECT 96.300 132.715 96.930 132.965 ;
        RECT 97.400 132.495 97.730 132.875 ;
        RECT 97.900 132.755 98.070 133.045 ;
        RECT 98.870 132.880 99.040 133.725 ;
        RECT 99.490 133.555 99.710 134.425 ;
        RECT 99.935 134.305 100.630 134.495 ;
        RECT 99.210 133.175 99.710 133.555 ;
        RECT 99.880 133.505 100.290 134.125 ;
        RECT 100.460 133.335 100.630 134.305 ;
        RECT 99.935 133.165 100.630 133.335 ;
        RECT 98.250 132.495 98.630 132.875 ;
        RECT 98.870 132.710 99.700 132.880 ;
        RECT 99.935 132.665 100.105 133.165 ;
        RECT 100.275 132.495 100.605 132.995 ;
        RECT 100.820 132.665 101.045 134.785 ;
        RECT 101.215 134.665 101.545 135.045 ;
        RECT 101.715 134.495 101.885 134.785 ;
        RECT 101.220 134.325 101.885 134.495 ;
        RECT 102.145 134.370 102.405 134.875 ;
        RECT 102.585 134.665 102.915 135.045 ;
        RECT 103.095 134.495 103.265 134.875 ;
        RECT 101.220 133.335 101.450 134.325 ;
        RECT 101.620 133.505 101.970 134.155 ;
        RECT 102.145 133.570 102.315 134.370 ;
        RECT 102.600 134.325 103.265 134.495 ;
        RECT 102.600 134.070 102.770 134.325 ;
        RECT 103.525 134.295 104.735 135.045 ;
        RECT 102.485 133.740 102.770 134.070 ;
        RECT 103.005 133.775 103.335 134.145 ;
        RECT 102.600 133.595 102.770 133.740 ;
        RECT 101.220 133.165 101.885 133.335 ;
        RECT 101.215 132.495 101.545 132.995 ;
        RECT 101.715 132.665 101.885 133.165 ;
        RECT 102.145 132.665 102.415 133.570 ;
        RECT 102.600 133.425 103.265 133.595 ;
        RECT 102.585 132.495 102.915 133.255 ;
        RECT 103.095 132.665 103.265 133.425 ;
        RECT 103.525 133.585 104.045 134.125 ;
        RECT 104.215 133.755 104.735 134.295 ;
        RECT 104.905 134.275 108.415 135.045 ;
        RECT 104.905 133.585 106.595 134.105 ;
        RECT 106.765 133.755 108.415 134.275 ;
        RECT 108.645 134.225 108.855 135.045 ;
        RECT 109.025 134.245 109.355 134.875 ;
        RECT 109.025 133.645 109.275 134.245 ;
        RECT 109.525 134.225 109.755 135.045 ;
        RECT 109.965 134.295 111.175 135.045 ;
        RECT 111.435 134.495 111.605 134.875 ;
        RECT 111.785 134.665 112.115 135.045 ;
        RECT 111.435 134.325 112.100 134.495 ;
        RECT 112.295 134.370 112.555 134.875 ;
        RECT 109.445 133.805 109.775 134.055 ;
        RECT 103.525 132.495 104.735 133.585 ;
        RECT 104.905 132.495 108.415 133.585 ;
        RECT 108.645 132.495 108.855 133.635 ;
        RECT 109.025 132.665 109.355 133.645 ;
        RECT 109.525 132.495 109.755 133.635 ;
        RECT 109.965 133.585 110.485 134.125 ;
        RECT 110.655 133.755 111.175 134.295 ;
        RECT 111.365 133.775 111.695 134.145 ;
        RECT 111.930 134.070 112.100 134.325 ;
        RECT 111.930 133.740 112.215 134.070 ;
        RECT 111.930 133.595 112.100 133.740 ;
        RECT 109.965 132.495 111.175 133.585 ;
        RECT 111.435 133.425 112.100 133.595 ;
        RECT 112.385 133.570 112.555 134.370 ;
        RECT 112.725 134.275 114.395 135.045 ;
        RECT 114.565 134.320 114.855 135.045 ;
        RECT 115.490 134.500 120.835 135.045 ;
        RECT 111.435 132.665 111.605 133.425 ;
        RECT 111.785 132.495 112.115 133.255 ;
        RECT 112.285 132.665 112.555 133.570 ;
        RECT 112.725 133.585 113.475 134.105 ;
        RECT 113.645 133.755 114.395 134.275 ;
        RECT 112.725 132.495 114.395 133.585 ;
        RECT 114.565 132.495 114.855 133.660 ;
        RECT 117.080 132.930 117.430 134.180 ;
        RECT 118.910 133.670 119.250 134.500 ;
        RECT 121.095 134.495 121.265 134.875 ;
        RECT 121.445 134.665 121.775 135.045 ;
        RECT 121.095 134.325 121.760 134.495 ;
        RECT 121.955 134.370 122.215 134.875 ;
        RECT 121.025 133.775 121.355 134.145 ;
        RECT 121.590 134.070 121.760 134.325 ;
        RECT 121.590 133.740 121.875 134.070 ;
        RECT 121.590 133.595 121.760 133.740 ;
        RECT 121.095 133.425 121.760 133.595 ;
        RECT 122.045 133.570 122.215 134.370 ;
        RECT 122.845 134.275 126.355 135.045 ;
        RECT 126.525 134.295 127.735 135.045 ;
        RECT 115.490 132.495 120.835 132.930 ;
        RECT 121.095 132.665 121.265 133.425 ;
        RECT 121.445 132.495 121.775 133.255 ;
        RECT 121.945 132.665 122.215 133.570 ;
        RECT 122.845 133.585 124.535 134.105 ;
        RECT 124.705 133.755 126.355 134.275 ;
        RECT 126.525 133.585 127.045 134.125 ;
        RECT 127.215 133.755 127.735 134.295 ;
        RECT 122.845 132.495 126.355 133.585 ;
        RECT 126.525 132.495 127.735 133.585 ;
        RECT 14.660 132.325 127.820 132.495 ;
        RECT 14.745 131.235 15.955 132.325 ;
        RECT 14.745 130.525 15.265 131.065 ;
        RECT 15.435 130.695 15.955 131.235 ;
        RECT 16.125 131.235 18.715 132.325 ;
        RECT 18.890 131.890 24.235 132.325 ;
        RECT 16.125 130.715 17.335 131.235 ;
        RECT 17.505 130.545 18.715 131.065 ;
        RECT 20.480 130.640 20.830 131.890 ;
        RECT 24.405 131.160 24.695 132.325 ;
        RECT 25.330 131.890 30.675 132.325 ;
        RECT 14.745 129.775 15.955 130.525 ;
        RECT 16.125 129.775 18.715 130.545 ;
        RECT 22.310 130.320 22.650 131.150 ;
        RECT 26.920 130.640 27.270 131.890 ;
        RECT 30.845 131.250 31.115 132.155 ;
        RECT 31.285 131.565 31.615 132.325 ;
        RECT 31.795 131.395 31.965 132.155 ;
        RECT 18.890 129.775 24.235 130.320 ;
        RECT 24.405 129.775 24.695 130.500 ;
        RECT 28.750 130.320 29.090 131.150 ;
        RECT 30.845 130.450 31.015 131.250 ;
        RECT 31.300 131.225 31.965 131.395 ;
        RECT 32.225 131.235 34.815 132.325 ;
        RECT 34.985 131.565 35.500 131.975 ;
        RECT 35.735 131.565 35.905 132.325 ;
        RECT 36.075 131.985 38.105 132.155 ;
        RECT 31.300 131.080 31.470 131.225 ;
        RECT 31.185 130.750 31.470 131.080 ;
        RECT 31.300 130.495 31.470 130.750 ;
        RECT 31.705 130.675 32.035 131.045 ;
        RECT 32.225 130.715 33.435 131.235 ;
        RECT 33.605 130.545 34.815 131.065 ;
        RECT 34.985 130.755 35.325 131.565 ;
        RECT 36.075 131.320 36.245 131.985 ;
        RECT 36.640 131.645 37.765 131.815 ;
        RECT 35.495 131.130 36.245 131.320 ;
        RECT 36.415 131.305 37.425 131.475 ;
        RECT 34.985 130.585 36.215 130.755 ;
        RECT 25.330 129.775 30.675 130.320 ;
        RECT 30.845 129.945 31.105 130.450 ;
        RECT 31.300 130.325 31.965 130.495 ;
        RECT 31.285 129.775 31.615 130.155 ;
        RECT 31.795 129.945 31.965 130.325 ;
        RECT 32.225 129.775 34.815 130.545 ;
        RECT 35.260 129.980 35.505 130.585 ;
        RECT 35.725 129.775 36.235 130.310 ;
        RECT 36.415 129.945 36.605 131.305 ;
        RECT 36.775 130.965 37.050 131.105 ;
        RECT 36.775 130.795 37.055 130.965 ;
        RECT 36.775 129.945 37.050 130.795 ;
        RECT 37.255 130.505 37.425 131.305 ;
        RECT 37.595 130.515 37.765 131.645 ;
        RECT 37.935 131.015 38.105 131.985 ;
        RECT 38.275 131.185 38.445 132.325 ;
        RECT 38.615 131.185 38.950 132.155 ;
        RECT 37.935 130.685 38.130 131.015 ;
        RECT 38.355 130.685 38.610 131.015 ;
        RECT 38.355 130.515 38.525 130.685 ;
        RECT 38.780 130.515 38.950 131.185 ;
        RECT 39.125 131.235 42.635 132.325 ;
        RECT 39.125 130.715 40.815 131.235 ;
        RECT 42.845 131.185 43.075 132.325 ;
        RECT 43.245 131.175 43.575 132.155 ;
        RECT 43.745 131.185 43.955 132.325 ;
        RECT 44.185 131.235 45.395 132.325 ;
        RECT 45.655 131.395 45.825 132.155 ;
        RECT 46.005 131.565 46.335 132.325 ;
        RECT 40.985 130.545 42.635 131.065 ;
        RECT 42.825 130.765 43.155 131.015 ;
        RECT 37.595 130.345 38.525 130.515 ;
        RECT 37.595 130.310 37.770 130.345 ;
        RECT 37.240 129.945 37.770 130.310 ;
        RECT 38.195 129.775 38.525 130.175 ;
        RECT 38.695 129.945 38.950 130.515 ;
        RECT 39.125 129.775 42.635 130.545 ;
        RECT 42.845 129.775 43.075 130.595 ;
        RECT 43.325 130.575 43.575 131.175 ;
        RECT 44.185 130.695 44.705 131.235 ;
        RECT 45.655 131.225 46.320 131.395 ;
        RECT 46.505 131.250 46.775 132.155 ;
        RECT 46.150 131.080 46.320 131.225 ;
        RECT 43.245 129.945 43.575 130.575 ;
        RECT 43.745 129.775 43.955 130.595 ;
        RECT 44.875 130.525 45.395 131.065 ;
        RECT 45.585 130.675 45.915 131.045 ;
        RECT 46.150 130.750 46.435 131.080 ;
        RECT 44.185 129.775 45.395 130.525 ;
        RECT 46.150 130.495 46.320 130.750 ;
        RECT 45.655 130.325 46.320 130.495 ;
        RECT 46.605 130.450 46.775 131.250 ;
        RECT 47.405 131.235 49.995 132.325 ;
        RECT 47.405 130.715 48.615 131.235 ;
        RECT 50.165 131.160 50.455 132.325 ;
        RECT 50.625 131.235 51.835 132.325 ;
        RECT 52.005 131.235 55.515 132.325 ;
        RECT 48.785 130.545 49.995 131.065 ;
        RECT 50.625 130.695 51.145 131.235 ;
        RECT 45.655 129.945 45.825 130.325 ;
        RECT 46.005 129.775 46.335 130.155 ;
        RECT 46.515 129.945 46.775 130.450 ;
        RECT 47.405 129.775 49.995 130.545 ;
        RECT 51.315 130.525 51.835 131.065 ;
        RECT 52.005 130.715 53.695 131.235 ;
        RECT 55.725 131.185 55.955 132.325 ;
        RECT 56.125 131.175 56.455 132.155 ;
        RECT 56.625 131.185 56.835 132.325 ;
        RECT 57.065 131.565 57.580 131.975 ;
        RECT 57.815 131.565 57.985 132.325 ;
        RECT 58.155 131.985 60.185 132.155 ;
        RECT 53.865 130.545 55.515 131.065 ;
        RECT 55.705 130.765 56.035 131.015 ;
        RECT 50.165 129.775 50.455 130.500 ;
        RECT 50.625 129.775 51.835 130.525 ;
        RECT 52.005 129.775 55.515 130.545 ;
        RECT 55.725 129.775 55.955 130.595 ;
        RECT 56.205 130.575 56.455 131.175 ;
        RECT 57.065 130.755 57.405 131.565 ;
        RECT 58.155 131.320 58.325 131.985 ;
        RECT 58.720 131.645 59.845 131.815 ;
        RECT 57.575 131.130 58.325 131.320 ;
        RECT 58.495 131.305 59.505 131.475 ;
        RECT 56.125 129.945 56.455 130.575 ;
        RECT 56.625 129.775 56.835 130.595 ;
        RECT 57.065 130.585 58.295 130.755 ;
        RECT 57.340 129.980 57.585 130.585 ;
        RECT 57.805 129.775 58.315 130.310 ;
        RECT 58.495 129.945 58.685 131.305 ;
        RECT 58.855 130.965 59.130 131.105 ;
        RECT 58.855 130.795 59.135 130.965 ;
        RECT 58.855 129.945 59.130 130.795 ;
        RECT 59.335 130.505 59.505 131.305 ;
        RECT 59.675 130.515 59.845 131.645 ;
        RECT 60.015 131.015 60.185 131.985 ;
        RECT 60.355 131.185 60.525 132.325 ;
        RECT 60.695 131.185 61.030 132.155 ;
        RECT 60.015 130.685 60.210 131.015 ;
        RECT 60.435 130.685 60.690 131.015 ;
        RECT 60.435 130.515 60.605 130.685 ;
        RECT 60.860 130.515 61.030 131.185 ;
        RECT 61.205 131.235 62.415 132.325 ;
        RECT 62.585 131.235 66.095 132.325 ;
        RECT 66.640 131.985 66.895 132.015 ;
        RECT 66.555 131.815 66.895 131.985 ;
        RECT 66.640 131.345 66.895 131.815 ;
        RECT 67.075 131.525 67.360 132.325 ;
        RECT 67.540 131.605 67.870 132.115 ;
        RECT 61.205 130.695 61.725 131.235 ;
        RECT 61.895 130.525 62.415 131.065 ;
        RECT 62.585 130.715 64.275 131.235 ;
        RECT 64.445 130.545 66.095 131.065 ;
        RECT 59.675 130.345 60.605 130.515 ;
        RECT 59.675 130.310 59.850 130.345 ;
        RECT 59.320 129.945 59.850 130.310 ;
        RECT 60.275 129.775 60.605 130.175 ;
        RECT 60.775 129.945 61.030 130.515 ;
        RECT 61.205 129.775 62.415 130.525 ;
        RECT 62.585 129.775 66.095 130.545 ;
        RECT 66.640 130.485 66.820 131.345 ;
        RECT 67.540 131.015 67.790 131.605 ;
        RECT 68.140 131.455 68.310 132.065 ;
        RECT 68.480 131.635 68.810 132.325 ;
        RECT 69.040 131.775 69.280 132.065 ;
        RECT 69.480 131.945 69.900 132.325 ;
        RECT 70.080 131.855 70.710 132.105 ;
        RECT 71.180 131.945 71.510 132.325 ;
        RECT 70.080 131.775 70.250 131.855 ;
        RECT 71.680 131.775 71.850 132.065 ;
        RECT 72.030 131.945 72.410 132.325 ;
        RECT 72.650 131.940 73.480 132.110 ;
        RECT 69.040 131.605 70.250 131.775 ;
        RECT 66.990 130.685 67.790 131.015 ;
        RECT 66.640 129.955 66.895 130.485 ;
        RECT 67.075 129.775 67.360 130.235 ;
        RECT 67.540 130.035 67.790 130.685 ;
        RECT 67.990 131.435 68.310 131.455 ;
        RECT 67.990 131.265 69.910 131.435 ;
        RECT 67.990 130.370 68.180 131.265 ;
        RECT 70.080 131.095 70.250 131.605 ;
        RECT 70.420 131.345 70.940 131.655 ;
        RECT 68.350 130.925 70.250 131.095 ;
        RECT 68.350 130.865 68.680 130.925 ;
        RECT 68.830 130.695 69.160 130.755 ;
        RECT 68.500 130.425 69.160 130.695 ;
        RECT 67.990 130.040 68.310 130.370 ;
        RECT 68.490 129.775 69.150 130.255 ;
        RECT 69.350 130.165 69.520 130.925 ;
        RECT 70.420 130.755 70.600 131.165 ;
        RECT 69.690 130.585 70.020 130.705 ;
        RECT 70.770 130.585 70.940 131.345 ;
        RECT 69.690 130.415 70.940 130.585 ;
        RECT 71.110 131.525 72.480 131.775 ;
        RECT 71.110 130.755 71.300 131.525 ;
        RECT 72.230 131.265 72.480 131.525 ;
        RECT 71.470 131.095 71.720 131.255 ;
        RECT 72.650 131.095 72.820 131.940 ;
        RECT 73.715 131.655 73.885 132.155 ;
        RECT 74.055 131.825 74.385 132.325 ;
        RECT 72.990 131.265 73.490 131.645 ;
        RECT 73.715 131.485 74.410 131.655 ;
        RECT 71.470 130.925 72.820 131.095 ;
        RECT 72.400 130.885 72.820 130.925 ;
        RECT 71.110 130.415 71.530 130.755 ;
        RECT 71.820 130.425 72.230 130.755 ;
        RECT 69.350 129.995 70.200 130.165 ;
        RECT 70.760 129.775 71.080 130.235 ;
        RECT 71.280 129.985 71.530 130.415 ;
        RECT 71.820 129.775 72.230 130.215 ;
        RECT 72.400 130.155 72.570 130.885 ;
        RECT 72.740 130.335 73.090 130.705 ;
        RECT 73.270 130.395 73.490 131.265 ;
        RECT 73.660 130.695 74.070 131.315 ;
        RECT 74.240 130.515 74.410 131.485 ;
        RECT 73.715 130.325 74.410 130.515 ;
        RECT 72.400 129.955 73.415 130.155 ;
        RECT 73.715 129.995 73.885 130.325 ;
        RECT 74.055 129.775 74.385 130.155 ;
        RECT 74.600 130.035 74.825 132.155 ;
        RECT 74.995 131.825 75.325 132.325 ;
        RECT 75.495 131.655 75.665 132.155 ;
        RECT 75.000 131.485 75.665 131.655 ;
        RECT 75.000 130.495 75.230 131.485 ;
        RECT 75.400 130.665 75.750 131.315 ;
        RECT 75.925 131.160 76.215 132.325 ;
        RECT 76.385 131.250 76.655 132.155 ;
        RECT 76.825 131.565 77.155 132.325 ;
        RECT 77.335 131.395 77.505 132.155 ;
        RECT 75.000 130.325 75.665 130.495 ;
        RECT 74.995 129.775 75.325 130.155 ;
        RECT 75.495 130.035 75.665 130.325 ;
        RECT 75.925 129.775 76.215 130.500 ;
        RECT 76.385 130.450 76.555 131.250 ;
        RECT 76.840 131.225 77.505 131.395 ;
        RECT 77.765 131.235 79.435 132.325 ;
        RECT 79.610 131.815 81.265 132.105 ;
        RECT 79.610 131.475 81.200 131.645 ;
        RECT 81.435 131.525 81.715 132.325 ;
        RECT 76.840 131.080 77.010 131.225 ;
        RECT 76.725 130.750 77.010 131.080 ;
        RECT 76.840 130.495 77.010 130.750 ;
        RECT 77.245 130.675 77.575 131.045 ;
        RECT 77.765 130.715 78.515 131.235 ;
        RECT 79.610 131.185 79.930 131.475 ;
        RECT 81.030 131.355 81.200 131.475 ;
        RECT 78.685 130.545 79.435 131.065 ;
        RECT 76.385 129.945 76.645 130.450 ;
        RECT 76.840 130.325 77.505 130.495 ;
        RECT 76.825 129.775 77.155 130.155 ;
        RECT 77.335 129.945 77.505 130.325 ;
        RECT 77.765 129.775 79.435 130.545 ;
        RECT 79.610 130.445 79.960 131.015 ;
        RECT 80.130 130.685 80.840 131.305 ;
        RECT 81.030 131.185 81.755 131.355 ;
        RECT 81.925 131.185 82.195 132.155 ;
        RECT 81.585 131.015 81.755 131.185 ;
        RECT 81.010 130.685 81.415 131.015 ;
        RECT 81.585 130.685 81.855 131.015 ;
        RECT 81.585 130.515 81.755 130.685 ;
        RECT 80.145 130.345 81.755 130.515 ;
        RECT 82.025 130.450 82.195 131.185 ;
        RECT 82.365 131.235 84.955 132.325 ;
        RECT 85.500 131.985 85.755 132.015 ;
        RECT 85.415 131.815 85.755 131.985 ;
        RECT 85.500 131.345 85.755 131.815 ;
        RECT 85.935 131.525 86.220 132.325 ;
        RECT 86.400 131.605 86.730 132.115 ;
        RECT 82.365 130.715 83.575 131.235 ;
        RECT 83.745 130.545 84.955 131.065 ;
        RECT 79.615 129.775 79.945 130.275 ;
        RECT 80.145 129.995 80.315 130.345 ;
        RECT 80.515 129.775 80.845 130.175 ;
        RECT 81.015 129.995 81.185 130.345 ;
        RECT 81.355 129.775 81.735 130.175 ;
        RECT 81.925 130.105 82.195 130.450 ;
        RECT 82.365 129.775 84.955 130.545 ;
        RECT 85.500 130.485 85.680 131.345 ;
        RECT 86.400 131.015 86.650 131.605 ;
        RECT 87.000 131.455 87.170 132.065 ;
        RECT 87.340 131.635 87.670 132.325 ;
        RECT 87.900 131.775 88.140 132.065 ;
        RECT 88.340 131.945 88.760 132.325 ;
        RECT 88.940 131.855 89.570 132.105 ;
        RECT 90.040 131.945 90.370 132.325 ;
        RECT 88.940 131.775 89.110 131.855 ;
        RECT 90.540 131.775 90.710 132.065 ;
        RECT 90.890 131.945 91.270 132.325 ;
        RECT 91.510 131.940 92.340 132.110 ;
        RECT 87.900 131.605 89.110 131.775 ;
        RECT 85.850 130.685 86.650 131.015 ;
        RECT 85.500 129.955 85.755 130.485 ;
        RECT 85.935 129.775 86.220 130.235 ;
        RECT 86.400 130.035 86.650 130.685 ;
        RECT 86.850 131.435 87.170 131.455 ;
        RECT 86.850 131.265 88.770 131.435 ;
        RECT 86.850 130.370 87.040 131.265 ;
        RECT 88.940 131.095 89.110 131.605 ;
        RECT 89.280 131.345 89.800 131.655 ;
        RECT 87.210 130.925 89.110 131.095 ;
        RECT 87.210 130.865 87.540 130.925 ;
        RECT 87.690 130.695 88.020 130.755 ;
        RECT 87.360 130.425 88.020 130.695 ;
        RECT 86.850 130.040 87.170 130.370 ;
        RECT 87.350 129.775 88.010 130.255 ;
        RECT 88.210 130.165 88.380 130.925 ;
        RECT 89.280 130.755 89.460 131.165 ;
        RECT 88.550 130.585 88.880 130.705 ;
        RECT 89.630 130.585 89.800 131.345 ;
        RECT 88.550 130.415 89.800 130.585 ;
        RECT 89.970 131.525 91.340 131.775 ;
        RECT 89.970 130.755 90.160 131.525 ;
        RECT 91.090 131.265 91.340 131.525 ;
        RECT 90.330 131.095 90.580 131.255 ;
        RECT 91.510 131.095 91.680 131.940 ;
        RECT 92.575 131.655 92.745 132.155 ;
        RECT 92.915 131.825 93.245 132.325 ;
        RECT 91.850 131.265 92.350 131.645 ;
        RECT 92.575 131.485 93.270 131.655 ;
        RECT 90.330 130.925 91.680 131.095 ;
        RECT 91.260 130.885 91.680 130.925 ;
        RECT 89.970 130.415 90.390 130.755 ;
        RECT 90.680 130.425 91.090 130.755 ;
        RECT 88.210 129.995 89.060 130.165 ;
        RECT 89.620 129.775 89.940 130.235 ;
        RECT 90.140 129.985 90.390 130.415 ;
        RECT 90.680 129.775 91.090 130.215 ;
        RECT 91.260 130.155 91.430 130.885 ;
        RECT 91.600 130.335 91.950 130.705 ;
        RECT 92.130 130.395 92.350 131.265 ;
        RECT 92.520 130.695 92.930 131.315 ;
        RECT 93.100 130.515 93.270 131.485 ;
        RECT 92.575 130.325 93.270 130.515 ;
        RECT 91.260 129.955 92.275 130.155 ;
        RECT 92.575 129.995 92.745 130.325 ;
        RECT 92.915 129.775 93.245 130.155 ;
        RECT 93.460 130.035 93.685 132.155 ;
        RECT 93.855 131.825 94.185 132.325 ;
        RECT 94.355 131.655 94.525 132.155 ;
        RECT 93.860 131.485 94.525 131.655 ;
        RECT 93.860 130.495 94.090 131.485 ;
        RECT 94.260 130.665 94.610 131.315 ;
        RECT 95.745 131.185 95.975 132.325 ;
        RECT 96.145 131.175 96.475 132.155 ;
        RECT 96.645 131.185 96.855 132.325 ;
        RECT 97.545 131.605 98.005 132.155 ;
        RECT 98.195 131.605 98.525 132.325 ;
        RECT 95.725 130.765 96.055 131.015 ;
        RECT 93.860 130.325 94.525 130.495 ;
        RECT 93.855 129.775 94.185 130.155 ;
        RECT 94.355 130.035 94.525 130.325 ;
        RECT 95.745 129.775 95.975 130.595 ;
        RECT 96.225 130.575 96.475 131.175 ;
        RECT 96.145 129.945 96.475 130.575 ;
        RECT 96.645 129.775 96.855 130.595 ;
        RECT 97.545 130.235 97.795 131.605 ;
        RECT 98.725 131.435 99.025 131.985 ;
        RECT 99.195 131.655 99.475 132.325 ;
        RECT 98.085 131.265 99.025 131.435 ;
        RECT 98.085 131.015 98.255 131.265 ;
        RECT 99.395 131.015 99.660 131.375 ;
        RECT 97.965 130.685 98.255 131.015 ;
        RECT 98.425 130.765 98.765 131.015 ;
        RECT 98.985 130.765 99.660 131.015 ;
        RECT 99.845 131.235 101.515 132.325 ;
        RECT 99.845 130.715 100.595 131.235 ;
        RECT 101.685 131.160 101.975 132.325 ;
        RECT 102.145 131.235 103.355 132.325 ;
        RECT 103.725 131.655 104.005 132.325 ;
        RECT 104.175 131.435 104.475 131.985 ;
        RECT 104.675 131.605 105.005 132.325 ;
        RECT 105.195 131.605 105.655 132.155 ;
        RECT 98.085 130.595 98.255 130.685 ;
        RECT 98.085 130.405 99.475 130.595 ;
        RECT 100.765 130.545 101.515 131.065 ;
        RECT 102.145 130.695 102.665 131.235 ;
        RECT 97.545 129.945 98.105 130.235 ;
        RECT 98.275 129.775 98.525 130.235 ;
        RECT 99.145 130.045 99.475 130.405 ;
        RECT 99.845 129.775 101.515 130.545 ;
        RECT 102.835 130.525 103.355 131.065 ;
        RECT 103.540 131.015 103.805 131.375 ;
        RECT 104.175 131.265 105.115 131.435 ;
        RECT 104.945 131.015 105.115 131.265 ;
        RECT 103.540 130.765 104.215 131.015 ;
        RECT 104.435 130.765 104.775 131.015 ;
        RECT 104.945 130.685 105.235 131.015 ;
        RECT 104.945 130.595 105.115 130.685 ;
        RECT 101.685 129.775 101.975 130.500 ;
        RECT 102.145 129.775 103.355 130.525 ;
        RECT 103.725 130.405 105.115 130.595 ;
        RECT 103.725 130.045 104.055 130.405 ;
        RECT 105.405 130.235 105.655 131.605 ;
        RECT 105.825 131.235 107.495 132.325 ;
        RECT 107.665 131.605 108.125 132.155 ;
        RECT 108.315 131.605 108.645 132.325 ;
        RECT 105.825 130.715 106.575 131.235 ;
        RECT 106.745 130.545 107.495 131.065 ;
        RECT 104.675 129.775 104.925 130.235 ;
        RECT 105.095 129.945 105.655 130.235 ;
        RECT 105.825 129.775 107.495 130.545 ;
        RECT 107.665 130.235 107.915 131.605 ;
        RECT 108.845 131.435 109.145 131.985 ;
        RECT 109.315 131.655 109.595 132.325 ;
        RECT 109.970 131.890 115.315 132.325 ;
        RECT 115.490 131.890 120.835 132.325 ;
        RECT 121.010 131.890 126.355 132.325 ;
        RECT 108.205 131.265 109.145 131.435 ;
        RECT 108.205 131.015 108.375 131.265 ;
        RECT 109.515 131.015 109.780 131.375 ;
        RECT 108.085 130.685 108.375 131.015 ;
        RECT 108.545 130.765 108.885 131.015 ;
        RECT 109.105 130.765 109.780 131.015 ;
        RECT 108.205 130.595 108.375 130.685 ;
        RECT 111.560 130.640 111.910 131.890 ;
        RECT 108.205 130.405 109.595 130.595 ;
        RECT 107.665 129.945 108.225 130.235 ;
        RECT 108.395 129.775 108.645 130.235 ;
        RECT 109.265 130.045 109.595 130.405 ;
        RECT 113.390 130.320 113.730 131.150 ;
        RECT 117.080 130.640 117.430 131.890 ;
        RECT 118.910 130.320 119.250 131.150 ;
        RECT 122.600 130.640 122.950 131.890 ;
        RECT 126.525 131.235 127.735 132.325 ;
        RECT 124.430 130.320 124.770 131.150 ;
        RECT 126.525 130.695 127.045 131.235 ;
        RECT 127.215 130.525 127.735 131.065 ;
        RECT 109.970 129.775 115.315 130.320 ;
        RECT 115.490 129.775 120.835 130.320 ;
        RECT 121.010 129.775 126.355 130.320 ;
        RECT 126.525 129.775 127.735 130.525 ;
        RECT 14.660 129.605 127.820 129.775 ;
        RECT 14.745 128.855 15.955 129.605 ;
        RECT 16.500 128.895 16.755 129.425 ;
        RECT 16.935 129.145 17.220 129.605 ;
        RECT 14.745 128.315 15.265 128.855 ;
        RECT 15.435 128.145 15.955 128.685 ;
        RECT 14.745 127.055 15.955 128.145 ;
        RECT 16.500 128.035 16.680 128.895 ;
        RECT 17.400 128.695 17.650 129.345 ;
        RECT 16.850 128.365 17.650 128.695 ;
        RECT 16.500 127.565 16.755 128.035 ;
        RECT 16.415 127.395 16.755 127.565 ;
        RECT 16.500 127.365 16.755 127.395 ;
        RECT 16.935 127.055 17.220 127.855 ;
        RECT 17.400 127.775 17.650 128.365 ;
        RECT 17.850 129.010 18.170 129.340 ;
        RECT 18.350 129.125 19.010 129.605 ;
        RECT 19.210 129.215 20.060 129.385 ;
        RECT 17.850 128.115 18.040 129.010 ;
        RECT 18.360 128.685 19.020 128.955 ;
        RECT 18.690 128.625 19.020 128.685 ;
        RECT 18.210 128.455 18.540 128.515 ;
        RECT 19.210 128.455 19.380 129.215 ;
        RECT 20.620 129.145 20.940 129.605 ;
        RECT 21.140 128.965 21.390 129.395 ;
        RECT 21.680 129.165 22.090 129.605 ;
        RECT 22.260 129.225 23.275 129.425 ;
        RECT 19.550 128.795 20.800 128.965 ;
        RECT 19.550 128.675 19.880 128.795 ;
        RECT 18.210 128.285 20.110 128.455 ;
        RECT 17.850 127.945 19.770 128.115 ;
        RECT 17.850 127.925 18.170 127.945 ;
        RECT 17.400 127.265 17.730 127.775 ;
        RECT 18.000 127.315 18.170 127.925 ;
        RECT 19.940 127.775 20.110 128.285 ;
        RECT 20.280 128.215 20.460 128.625 ;
        RECT 20.630 128.035 20.800 128.795 ;
        RECT 18.340 127.055 18.670 127.745 ;
        RECT 18.900 127.605 20.110 127.775 ;
        RECT 20.280 127.725 20.800 128.035 ;
        RECT 20.970 128.625 21.390 128.965 ;
        RECT 21.680 128.625 22.090 128.955 ;
        RECT 20.970 127.855 21.160 128.625 ;
        RECT 22.260 128.495 22.430 129.225 ;
        RECT 23.575 129.055 23.745 129.385 ;
        RECT 23.915 129.225 24.245 129.605 ;
        RECT 22.600 128.675 22.950 129.045 ;
        RECT 22.260 128.455 22.680 128.495 ;
        RECT 21.330 128.285 22.680 128.455 ;
        RECT 21.330 128.125 21.580 128.285 ;
        RECT 22.090 127.855 22.340 128.115 ;
        RECT 20.970 127.605 22.340 127.855 ;
        RECT 18.900 127.315 19.140 127.605 ;
        RECT 19.940 127.525 20.110 127.605 ;
        RECT 19.340 127.055 19.760 127.435 ;
        RECT 19.940 127.275 20.570 127.525 ;
        RECT 21.040 127.055 21.370 127.435 ;
        RECT 21.540 127.315 21.710 127.605 ;
        RECT 22.510 127.440 22.680 128.285 ;
        RECT 23.130 128.115 23.350 128.985 ;
        RECT 23.575 128.865 24.270 129.055 ;
        RECT 22.850 127.735 23.350 128.115 ;
        RECT 23.520 128.065 23.930 128.685 ;
        RECT 24.100 127.895 24.270 128.865 ;
        RECT 23.575 127.725 24.270 127.895 ;
        RECT 21.890 127.055 22.270 127.435 ;
        RECT 22.510 127.270 23.340 127.440 ;
        RECT 23.575 127.225 23.745 127.725 ;
        RECT 23.915 127.055 24.245 127.555 ;
        RECT 24.460 127.225 24.685 129.345 ;
        RECT 24.855 129.225 25.185 129.605 ;
        RECT 25.355 129.055 25.525 129.345 ;
        RECT 26.250 129.060 31.595 129.605 ;
        RECT 31.770 129.060 37.115 129.605 ;
        RECT 24.860 128.885 25.525 129.055 ;
        RECT 24.860 127.895 25.090 128.885 ;
        RECT 25.260 128.065 25.610 128.715 ;
        RECT 24.860 127.725 25.525 127.895 ;
        RECT 24.855 127.055 25.185 127.555 ;
        RECT 25.355 127.225 25.525 127.725 ;
        RECT 27.840 127.490 28.190 128.740 ;
        RECT 29.670 128.230 30.010 129.060 ;
        RECT 33.360 127.490 33.710 128.740 ;
        RECT 35.190 128.230 35.530 129.060 ;
        RECT 37.285 128.880 37.575 129.605 ;
        RECT 38.670 129.060 44.015 129.605 ;
        RECT 44.245 129.125 44.525 129.605 ;
        RECT 26.250 127.055 31.595 127.490 ;
        RECT 31.770 127.055 37.115 127.490 ;
        RECT 37.285 127.055 37.575 128.220 ;
        RECT 40.260 127.490 40.610 128.740 ;
        RECT 42.090 128.230 42.430 129.060 ;
        RECT 44.695 128.955 44.955 129.345 ;
        RECT 45.130 129.125 45.385 129.605 ;
        RECT 45.555 128.955 45.850 129.345 ;
        RECT 46.030 129.125 46.305 129.605 ;
        RECT 46.475 129.105 46.775 129.435 ;
        RECT 46.955 129.105 47.285 129.605 ;
        RECT 44.200 128.785 45.850 128.955 ;
        RECT 44.200 128.275 44.605 128.785 ;
        RECT 44.775 128.445 45.915 128.615 ;
        RECT 44.200 128.105 44.955 128.275 ;
        RECT 38.670 127.055 44.015 127.490 ;
        RECT 44.240 127.055 44.525 127.925 ;
        RECT 44.695 127.855 44.955 128.105 ;
        RECT 45.745 128.195 45.915 128.445 ;
        RECT 46.085 128.365 46.435 128.935 ;
        RECT 46.605 128.195 46.775 129.105 ;
        RECT 47.485 129.035 47.655 129.385 ;
        RECT 47.855 129.205 48.185 129.605 ;
        RECT 48.355 129.035 48.525 129.385 ;
        RECT 48.695 129.205 49.075 129.605 ;
        RECT 46.950 128.365 47.300 128.935 ;
        RECT 47.485 128.865 49.095 129.035 ;
        RECT 49.265 128.930 49.535 129.275 ;
        RECT 48.925 128.695 49.095 128.865 ;
        RECT 45.745 128.025 46.775 128.195 ;
        RECT 44.695 127.685 45.815 127.855 ;
        RECT 44.695 127.225 44.955 127.685 ;
        RECT 45.130 127.055 45.385 127.515 ;
        RECT 45.555 127.225 45.815 127.685 ;
        RECT 45.985 127.055 46.295 127.855 ;
        RECT 46.465 127.225 46.775 128.025 ;
        RECT 46.950 127.905 47.270 128.195 ;
        RECT 47.470 128.075 48.180 128.695 ;
        RECT 48.350 128.365 48.755 128.695 ;
        RECT 48.925 128.365 49.195 128.695 ;
        RECT 48.925 128.195 49.095 128.365 ;
        RECT 49.365 128.195 49.535 128.930 ;
        RECT 48.370 128.025 49.095 128.195 ;
        RECT 48.370 127.905 48.540 128.025 ;
        RECT 46.950 127.735 48.540 127.905 ;
        RECT 46.950 127.275 48.605 127.565 ;
        RECT 48.775 127.055 49.055 127.855 ;
        RECT 49.265 127.225 49.535 128.195 ;
        RECT 49.705 128.805 50.045 129.435 ;
        RECT 50.215 128.805 50.465 129.605 ;
        RECT 50.655 128.955 50.985 129.435 ;
        RECT 51.155 129.145 51.380 129.605 ;
        RECT 51.550 128.955 51.880 129.435 ;
        RECT 49.705 128.755 49.935 128.805 ;
        RECT 50.655 128.785 51.880 128.955 ;
        RECT 52.510 128.825 53.010 129.435 ;
        RECT 53.760 129.265 54.015 129.425 ;
        RECT 53.675 129.095 54.015 129.265 ;
        RECT 54.195 129.145 54.480 129.605 ;
        RECT 53.760 128.895 54.015 129.095 ;
        RECT 49.705 128.195 49.880 128.755 ;
        RECT 50.050 128.445 50.745 128.615 ;
        RECT 50.575 128.195 50.745 128.445 ;
        RECT 50.920 128.415 51.340 128.615 ;
        RECT 51.510 128.415 51.840 128.615 ;
        RECT 52.010 128.415 52.340 128.615 ;
        RECT 52.510 128.195 52.680 128.825 ;
        RECT 52.865 128.365 53.215 128.615 ;
        RECT 49.705 127.225 50.045 128.195 ;
        RECT 50.215 127.055 50.385 128.195 ;
        RECT 50.575 128.025 53.010 128.195 ;
        RECT 50.655 127.055 50.905 127.855 ;
        RECT 51.550 127.225 51.880 128.025 ;
        RECT 52.180 127.055 52.510 127.855 ;
        RECT 52.680 127.225 53.010 128.025 ;
        RECT 53.760 128.035 53.940 128.895 ;
        RECT 54.660 128.695 54.910 129.345 ;
        RECT 54.110 128.365 54.910 128.695 ;
        RECT 53.760 127.365 54.015 128.035 ;
        RECT 54.195 127.055 54.480 127.855 ;
        RECT 54.660 127.775 54.910 128.365 ;
        RECT 55.110 129.010 55.430 129.340 ;
        RECT 55.610 129.125 56.270 129.605 ;
        RECT 56.470 129.215 57.320 129.385 ;
        RECT 55.110 128.115 55.300 129.010 ;
        RECT 55.620 128.685 56.280 128.955 ;
        RECT 55.950 128.625 56.280 128.685 ;
        RECT 55.470 128.455 55.800 128.515 ;
        RECT 56.470 128.455 56.640 129.215 ;
        RECT 57.880 129.145 58.200 129.605 ;
        RECT 58.400 128.965 58.650 129.395 ;
        RECT 58.940 129.165 59.350 129.605 ;
        RECT 59.520 129.225 60.535 129.425 ;
        RECT 56.810 128.795 58.060 128.965 ;
        RECT 56.810 128.675 57.140 128.795 ;
        RECT 55.470 128.285 57.370 128.455 ;
        RECT 55.110 127.945 57.030 128.115 ;
        RECT 55.110 127.925 55.430 127.945 ;
        RECT 54.660 127.265 54.990 127.775 ;
        RECT 55.260 127.315 55.430 127.925 ;
        RECT 57.200 127.775 57.370 128.285 ;
        RECT 57.540 128.215 57.720 128.625 ;
        RECT 57.890 128.035 58.060 128.795 ;
        RECT 55.600 127.055 55.930 127.745 ;
        RECT 56.160 127.605 57.370 127.775 ;
        RECT 57.540 127.725 58.060 128.035 ;
        RECT 58.230 128.625 58.650 128.965 ;
        RECT 58.940 128.625 59.350 128.955 ;
        RECT 58.230 127.855 58.420 128.625 ;
        RECT 59.520 128.495 59.690 129.225 ;
        RECT 60.835 129.055 61.005 129.385 ;
        RECT 61.175 129.225 61.505 129.605 ;
        RECT 59.860 128.675 60.210 129.045 ;
        RECT 59.520 128.455 59.940 128.495 ;
        RECT 58.590 128.285 59.940 128.455 ;
        RECT 58.590 128.125 58.840 128.285 ;
        RECT 59.350 127.855 59.600 128.115 ;
        RECT 58.230 127.605 59.600 127.855 ;
        RECT 56.160 127.315 56.400 127.605 ;
        RECT 57.200 127.525 57.370 127.605 ;
        RECT 56.600 127.055 57.020 127.435 ;
        RECT 57.200 127.275 57.830 127.525 ;
        RECT 58.300 127.055 58.630 127.435 ;
        RECT 58.800 127.315 58.970 127.605 ;
        RECT 59.770 127.440 59.940 128.285 ;
        RECT 60.390 128.115 60.610 128.985 ;
        RECT 60.835 128.865 61.530 129.055 ;
        RECT 60.110 127.735 60.610 128.115 ;
        RECT 60.780 128.065 61.190 128.685 ;
        RECT 61.360 127.895 61.530 128.865 ;
        RECT 60.835 127.725 61.530 127.895 ;
        RECT 59.150 127.055 59.530 127.435 ;
        RECT 59.770 127.270 60.600 127.440 ;
        RECT 60.835 127.225 61.005 127.725 ;
        RECT 61.175 127.055 61.505 127.555 ;
        RECT 61.720 127.225 61.945 129.345 ;
        RECT 62.115 129.225 62.445 129.605 ;
        RECT 62.615 129.055 62.785 129.345 ;
        RECT 62.120 128.885 62.785 129.055 ;
        RECT 62.120 127.895 62.350 128.885 ;
        RECT 63.045 128.880 63.335 129.605 ;
        RECT 63.505 128.930 63.765 129.435 ;
        RECT 63.945 129.225 64.275 129.605 ;
        RECT 64.455 129.055 64.625 129.435 ;
        RECT 62.520 128.065 62.870 128.715 ;
        RECT 62.120 127.725 62.785 127.895 ;
        RECT 62.115 127.055 62.445 127.555 ;
        RECT 62.615 127.225 62.785 127.725 ;
        RECT 63.045 127.055 63.335 128.220 ;
        RECT 63.505 128.130 63.675 128.930 ;
        RECT 63.960 128.885 64.625 129.055 ;
        RECT 63.960 128.630 64.130 128.885 ;
        RECT 65.345 128.835 67.935 129.605 ;
        RECT 63.845 128.300 64.130 128.630 ;
        RECT 64.365 128.335 64.695 128.705 ;
        RECT 63.960 128.155 64.130 128.300 ;
        RECT 63.505 127.225 63.775 128.130 ;
        RECT 63.960 127.985 64.625 128.155 ;
        RECT 63.945 127.055 64.275 127.815 ;
        RECT 64.455 127.225 64.625 127.985 ;
        RECT 65.345 128.145 66.555 128.665 ;
        RECT 66.725 128.315 67.935 128.835 ;
        RECT 68.145 128.785 68.375 129.605 ;
        RECT 68.545 128.805 68.875 129.435 ;
        RECT 68.125 128.365 68.455 128.615 ;
        RECT 68.625 128.205 68.875 128.805 ;
        RECT 69.045 128.785 69.255 129.605 ;
        RECT 69.685 128.975 70.015 129.335 ;
        RECT 70.635 129.145 70.885 129.605 ;
        RECT 71.055 129.145 71.615 129.435 ;
        RECT 69.685 128.785 71.075 128.975 ;
        RECT 70.905 128.695 71.075 128.785 ;
        RECT 65.345 127.055 67.935 128.145 ;
        RECT 68.145 127.055 68.375 128.195 ;
        RECT 68.545 127.225 68.875 128.205 ;
        RECT 69.500 128.365 70.175 128.615 ;
        RECT 70.395 128.365 70.735 128.615 ;
        RECT 70.905 128.365 71.195 128.695 ;
        RECT 69.045 127.055 69.255 128.195 ;
        RECT 69.500 128.005 69.765 128.365 ;
        RECT 70.905 128.115 71.075 128.365 ;
        RECT 70.135 127.945 71.075 128.115 ;
        RECT 69.685 127.055 69.965 127.725 ;
        RECT 70.135 127.395 70.435 127.945 ;
        RECT 71.365 127.775 71.615 129.145 ;
        RECT 70.635 127.055 70.965 127.775 ;
        RECT 71.155 127.225 71.615 127.775 ;
        RECT 71.785 129.105 72.085 129.435 ;
        RECT 72.255 129.125 72.530 129.605 ;
        RECT 71.785 128.195 71.955 129.105 ;
        RECT 72.710 128.955 73.005 129.345 ;
        RECT 73.175 129.125 73.430 129.605 ;
        RECT 73.605 128.955 73.865 129.345 ;
        RECT 74.035 129.125 74.315 129.605 ;
        RECT 72.125 128.365 72.475 128.935 ;
        RECT 72.710 128.785 74.360 128.955 ;
        RECT 74.545 128.855 75.755 129.605 ;
        RECT 72.645 128.445 73.785 128.615 ;
        RECT 72.645 128.195 72.815 128.445 ;
        RECT 73.955 128.275 74.360 128.785 ;
        RECT 71.785 128.025 72.815 128.195 ;
        RECT 73.605 128.105 74.360 128.275 ;
        RECT 74.545 128.145 75.065 128.685 ;
        RECT 75.235 128.315 75.755 128.855 ;
        RECT 75.925 128.835 79.435 129.605 ;
        RECT 75.925 128.145 77.615 128.665 ;
        RECT 77.785 128.315 79.435 128.835 ;
        RECT 79.605 129.145 80.165 129.435 ;
        RECT 80.335 129.145 80.585 129.605 ;
        RECT 71.785 127.225 72.095 128.025 ;
        RECT 73.605 127.855 73.865 128.105 ;
        RECT 72.265 127.055 72.575 127.855 ;
        RECT 72.745 127.685 73.865 127.855 ;
        RECT 72.745 127.225 73.005 127.685 ;
        RECT 73.175 127.055 73.430 127.515 ;
        RECT 73.605 127.225 73.865 127.685 ;
        RECT 74.035 127.055 74.320 127.925 ;
        RECT 74.545 127.055 75.755 128.145 ;
        RECT 75.925 127.055 79.435 128.145 ;
        RECT 79.605 127.775 79.855 129.145 ;
        RECT 81.205 128.975 81.535 129.335 ;
        RECT 80.145 128.785 81.535 128.975 ;
        RECT 81.905 129.145 82.465 129.435 ;
        RECT 82.635 129.145 82.885 129.605 ;
        RECT 80.145 128.695 80.315 128.785 ;
        RECT 80.025 128.365 80.315 128.695 ;
        RECT 80.485 128.365 80.825 128.615 ;
        RECT 81.045 128.365 81.720 128.615 ;
        RECT 80.145 128.115 80.315 128.365 ;
        RECT 80.145 127.945 81.085 128.115 ;
        RECT 81.455 128.005 81.720 128.365 ;
        RECT 79.605 127.225 80.065 127.775 ;
        RECT 80.255 127.055 80.585 127.775 ;
        RECT 80.785 127.395 81.085 127.945 ;
        RECT 81.905 127.775 82.155 129.145 ;
        RECT 83.505 128.975 83.835 129.335 ;
        RECT 82.445 128.785 83.835 128.975 ;
        RECT 85.125 128.835 88.635 129.605 ;
        RECT 88.805 128.880 89.095 129.605 ;
        RECT 89.265 128.855 90.475 129.605 ;
        RECT 82.445 128.695 82.615 128.785 ;
        RECT 82.325 128.365 82.615 128.695 ;
        RECT 82.785 128.365 83.125 128.615 ;
        RECT 83.345 128.365 84.020 128.615 ;
        RECT 82.445 128.115 82.615 128.365 ;
        RECT 82.445 127.945 83.385 128.115 ;
        RECT 83.755 128.005 84.020 128.365 ;
        RECT 85.125 128.145 86.815 128.665 ;
        RECT 86.985 128.315 88.635 128.835 ;
        RECT 81.255 127.055 81.535 127.725 ;
        RECT 81.905 127.225 82.365 127.775 ;
        RECT 82.555 127.055 82.885 127.775 ;
        RECT 83.085 127.395 83.385 127.945 ;
        RECT 83.555 127.055 83.835 127.725 ;
        RECT 85.125 127.055 88.635 128.145 ;
        RECT 88.805 127.055 89.095 128.220 ;
        RECT 89.265 128.145 89.785 128.685 ;
        RECT 89.955 128.315 90.475 128.855 ;
        RECT 90.645 128.835 94.155 129.605 ;
        RECT 94.330 129.060 99.675 129.605 ;
        RECT 99.850 129.060 105.195 129.605 ;
        RECT 105.365 129.145 105.925 129.435 ;
        RECT 106.095 129.145 106.345 129.605 ;
        RECT 90.645 128.145 92.335 128.665 ;
        RECT 92.505 128.315 94.155 128.835 ;
        RECT 89.265 127.055 90.475 128.145 ;
        RECT 90.645 127.055 94.155 128.145 ;
        RECT 95.920 127.490 96.270 128.740 ;
        RECT 97.750 128.230 98.090 129.060 ;
        RECT 101.440 127.490 101.790 128.740 ;
        RECT 103.270 128.230 103.610 129.060 ;
        RECT 105.365 127.775 105.615 129.145 ;
        RECT 106.965 128.975 107.295 129.335 ;
        RECT 105.905 128.785 107.295 128.975 ;
        RECT 107.665 129.145 108.225 129.435 ;
        RECT 108.395 129.145 108.645 129.605 ;
        RECT 105.905 128.695 106.075 128.785 ;
        RECT 105.785 128.365 106.075 128.695 ;
        RECT 106.245 128.365 106.585 128.615 ;
        RECT 106.805 128.365 107.480 128.615 ;
        RECT 105.905 128.115 106.075 128.365 ;
        RECT 105.905 127.945 106.845 128.115 ;
        RECT 107.215 128.005 107.480 128.365 ;
        RECT 94.330 127.055 99.675 127.490 ;
        RECT 99.850 127.055 105.195 127.490 ;
        RECT 105.365 127.225 105.825 127.775 ;
        RECT 106.015 127.055 106.345 127.775 ;
        RECT 106.545 127.395 106.845 127.945 ;
        RECT 107.665 127.775 107.915 129.145 ;
        RECT 109.265 128.975 109.595 129.335 ;
        RECT 108.205 128.785 109.595 128.975 ;
        RECT 109.965 129.145 110.525 129.435 ;
        RECT 110.695 129.145 110.945 129.605 ;
        RECT 108.205 128.695 108.375 128.785 ;
        RECT 108.085 128.365 108.375 128.695 ;
        RECT 108.545 128.365 108.885 128.615 ;
        RECT 109.105 128.365 109.780 128.615 ;
        RECT 108.205 128.115 108.375 128.365 ;
        RECT 108.205 127.945 109.145 128.115 ;
        RECT 109.515 128.005 109.780 128.365 ;
        RECT 107.015 127.055 107.295 127.725 ;
        RECT 107.665 127.225 108.125 127.775 ;
        RECT 108.315 127.055 108.645 127.775 ;
        RECT 108.845 127.395 109.145 127.945 ;
        RECT 109.965 127.775 110.215 129.145 ;
        RECT 111.565 128.975 111.895 129.335 ;
        RECT 110.505 128.785 111.895 128.975 ;
        RECT 112.725 128.835 114.395 129.605 ;
        RECT 114.565 128.880 114.855 129.605 ;
        RECT 110.505 128.695 110.675 128.785 ;
        RECT 110.385 128.365 110.675 128.695 ;
        RECT 110.845 128.365 111.185 128.615 ;
        RECT 111.405 128.365 112.080 128.615 ;
        RECT 110.505 128.115 110.675 128.365 ;
        RECT 110.505 127.945 111.445 128.115 ;
        RECT 111.815 128.005 112.080 128.365 ;
        RECT 112.725 128.145 113.475 128.665 ;
        RECT 113.645 128.315 114.395 128.835 ;
        RECT 115.300 128.795 115.545 129.400 ;
        RECT 115.765 129.070 116.275 129.605 ;
        RECT 115.025 128.625 116.255 128.795 ;
        RECT 109.315 127.055 109.595 127.725 ;
        RECT 109.965 127.225 110.425 127.775 ;
        RECT 110.615 127.055 110.945 127.775 ;
        RECT 111.145 127.395 111.445 127.945 ;
        RECT 111.615 127.055 111.895 127.725 ;
        RECT 112.725 127.055 114.395 128.145 ;
        RECT 114.565 127.055 114.855 128.220 ;
        RECT 115.025 127.815 115.365 128.625 ;
        RECT 115.535 128.060 116.285 128.250 ;
        RECT 115.025 127.405 115.540 127.815 ;
        RECT 115.775 127.055 115.945 127.815 ;
        RECT 116.115 127.395 116.285 128.060 ;
        RECT 116.455 128.075 116.645 129.435 ;
        RECT 116.815 128.585 117.090 129.435 ;
        RECT 117.280 129.070 117.810 129.435 ;
        RECT 118.235 129.205 118.565 129.605 ;
        RECT 117.635 129.035 117.810 129.070 ;
        RECT 116.815 128.415 117.095 128.585 ;
        RECT 116.815 128.275 117.090 128.415 ;
        RECT 117.295 128.075 117.465 128.875 ;
        RECT 116.455 127.905 117.465 128.075 ;
        RECT 117.635 128.865 118.565 129.035 ;
        RECT 118.735 128.865 118.990 129.435 ;
        RECT 117.635 127.735 117.805 128.865 ;
        RECT 118.395 128.695 118.565 128.865 ;
        RECT 116.680 127.565 117.805 127.735 ;
        RECT 117.975 128.365 118.170 128.695 ;
        RECT 118.395 128.365 118.650 128.695 ;
        RECT 117.975 127.395 118.145 128.365 ;
        RECT 118.820 128.195 118.990 128.865 ;
        RECT 119.165 128.835 120.835 129.605 ;
        RECT 121.010 129.060 126.355 129.605 ;
        RECT 116.115 127.225 118.145 127.395 ;
        RECT 118.315 127.055 118.485 128.195 ;
        RECT 118.655 127.225 118.990 128.195 ;
        RECT 119.165 128.145 119.915 128.665 ;
        RECT 120.085 128.315 120.835 128.835 ;
        RECT 119.165 127.055 120.835 128.145 ;
        RECT 122.600 127.490 122.950 128.740 ;
        RECT 124.430 128.230 124.770 129.060 ;
        RECT 126.525 128.855 127.735 129.605 ;
        RECT 126.525 128.145 127.045 128.685 ;
        RECT 127.215 128.315 127.735 128.855 ;
        RECT 121.010 127.055 126.355 127.490 ;
        RECT 126.525 127.055 127.735 128.145 ;
        RECT 14.660 126.885 127.820 127.055 ;
        RECT 14.745 125.795 15.955 126.885 ;
        RECT 14.745 125.085 15.265 125.625 ;
        RECT 15.435 125.255 15.955 125.795 ;
        RECT 16.125 125.795 18.715 126.885 ;
        RECT 18.890 126.450 24.235 126.885 ;
        RECT 16.125 125.275 17.335 125.795 ;
        RECT 17.505 125.105 18.715 125.625 ;
        RECT 20.480 125.200 20.830 126.450 ;
        RECT 24.405 125.720 24.695 126.885 ;
        RECT 25.785 125.795 29.295 126.885 ;
        RECT 29.555 125.955 29.725 126.715 ;
        RECT 29.905 126.125 30.235 126.885 ;
        RECT 14.745 124.335 15.955 125.085 ;
        RECT 16.125 124.335 18.715 125.105 ;
        RECT 22.310 124.880 22.650 125.710 ;
        RECT 25.785 125.275 27.475 125.795 ;
        RECT 29.555 125.785 30.220 125.955 ;
        RECT 30.405 125.810 30.675 126.715 ;
        RECT 30.900 126.015 31.185 126.885 ;
        RECT 31.355 126.255 31.615 126.715 ;
        RECT 31.790 126.425 32.045 126.885 ;
        RECT 32.215 126.255 32.475 126.715 ;
        RECT 31.355 126.085 32.475 126.255 ;
        RECT 32.645 126.085 32.955 126.885 ;
        RECT 31.355 125.835 31.615 126.085 ;
        RECT 33.125 125.915 33.435 126.715 ;
        RECT 30.050 125.640 30.220 125.785 ;
        RECT 27.645 125.105 29.295 125.625 ;
        RECT 29.485 125.235 29.815 125.605 ;
        RECT 30.050 125.310 30.335 125.640 ;
        RECT 18.890 124.335 24.235 124.880 ;
        RECT 24.405 124.335 24.695 125.060 ;
        RECT 25.785 124.335 29.295 125.105 ;
        RECT 30.050 125.055 30.220 125.310 ;
        RECT 29.555 124.885 30.220 125.055 ;
        RECT 30.505 125.010 30.675 125.810 ;
        RECT 29.555 124.505 29.725 124.885 ;
        RECT 29.905 124.335 30.235 124.715 ;
        RECT 30.415 124.505 30.675 125.010 ;
        RECT 30.860 125.665 31.615 125.835 ;
        RECT 32.405 125.745 33.435 125.915 ;
        RECT 30.860 125.155 31.265 125.665 ;
        RECT 32.405 125.495 32.575 125.745 ;
        RECT 31.435 125.325 32.575 125.495 ;
        RECT 30.860 124.985 32.510 125.155 ;
        RECT 32.745 125.005 33.095 125.575 ;
        RECT 30.905 124.335 31.185 124.815 ;
        RECT 31.355 124.595 31.615 124.985 ;
        RECT 31.790 124.335 32.045 124.815 ;
        RECT 32.215 124.595 32.510 124.985 ;
        RECT 33.265 124.835 33.435 125.745 ;
        RECT 34.525 125.795 38.035 126.885 ;
        RECT 34.525 125.275 36.215 125.795 ;
        RECT 38.205 125.745 38.475 126.715 ;
        RECT 38.685 126.085 38.965 126.885 ;
        RECT 39.135 126.375 40.790 126.665 ;
        RECT 39.200 126.035 40.790 126.205 ;
        RECT 39.200 125.915 39.370 126.035 ;
        RECT 38.645 125.745 39.370 125.915 ;
        RECT 36.385 125.105 38.035 125.625 ;
        RECT 32.690 124.335 32.965 124.815 ;
        RECT 33.135 124.505 33.435 124.835 ;
        RECT 34.525 124.335 38.035 125.105 ;
        RECT 38.205 125.010 38.375 125.745 ;
        RECT 38.645 125.575 38.815 125.745 ;
        RECT 38.545 125.245 38.815 125.575 ;
        RECT 38.985 125.245 39.390 125.575 ;
        RECT 39.560 125.245 40.270 125.865 ;
        RECT 40.470 125.745 40.790 126.035 ;
        RECT 40.965 125.745 41.235 126.715 ;
        RECT 41.445 126.085 41.725 126.885 ;
        RECT 41.895 126.375 43.550 126.665 ;
        RECT 43.730 126.375 45.385 126.665 ;
        RECT 41.960 126.035 43.550 126.205 ;
        RECT 41.960 125.915 42.130 126.035 ;
        RECT 41.405 125.745 42.130 125.915 ;
        RECT 38.645 125.075 38.815 125.245 ;
        RECT 38.205 124.665 38.475 125.010 ;
        RECT 38.645 124.905 40.255 125.075 ;
        RECT 40.440 125.005 40.790 125.575 ;
        RECT 40.965 125.010 41.135 125.745 ;
        RECT 41.405 125.575 41.575 125.745 ;
        RECT 41.305 125.245 41.575 125.575 ;
        RECT 41.745 125.245 42.150 125.575 ;
        RECT 42.320 125.245 43.030 125.865 ;
        RECT 43.230 125.745 43.550 126.035 ;
        RECT 43.730 126.035 45.320 126.205 ;
        RECT 45.555 126.085 45.835 126.885 ;
        RECT 43.730 125.745 44.050 126.035 ;
        RECT 45.150 125.915 45.320 126.035 ;
        RECT 41.405 125.075 41.575 125.245 ;
        RECT 38.665 124.335 39.045 124.735 ;
        RECT 39.215 124.555 39.385 124.905 ;
        RECT 39.555 124.335 39.885 124.735 ;
        RECT 40.085 124.555 40.255 124.905 ;
        RECT 40.455 124.335 40.785 124.835 ;
        RECT 40.965 124.665 41.235 125.010 ;
        RECT 41.405 124.905 43.015 125.075 ;
        RECT 43.200 125.005 43.550 125.575 ;
        RECT 43.730 125.005 44.080 125.575 ;
        RECT 44.250 125.245 44.960 125.865 ;
        RECT 45.150 125.745 45.875 125.915 ;
        RECT 46.045 125.745 46.315 126.715 ;
        RECT 45.705 125.575 45.875 125.745 ;
        RECT 45.130 125.245 45.535 125.575 ;
        RECT 45.705 125.245 45.975 125.575 ;
        RECT 45.705 125.075 45.875 125.245 ;
        RECT 41.425 124.335 41.805 124.735 ;
        RECT 41.975 124.555 42.145 124.905 ;
        RECT 42.315 124.335 42.645 124.735 ;
        RECT 42.845 124.555 43.015 124.905 ;
        RECT 44.265 124.905 45.875 125.075 ;
        RECT 46.145 125.010 46.315 125.745 ;
        RECT 43.215 124.335 43.545 124.835 ;
        RECT 43.735 124.335 44.065 124.835 ;
        RECT 44.265 124.555 44.435 124.905 ;
        RECT 44.635 124.335 44.965 124.735 ;
        RECT 45.135 124.555 45.305 124.905 ;
        RECT 45.475 124.335 45.855 124.735 ;
        RECT 46.045 124.665 46.315 125.010 ;
        RECT 46.485 125.745 46.825 126.715 ;
        RECT 46.995 125.745 47.165 126.885 ;
        RECT 47.435 126.085 47.685 126.885 ;
        RECT 48.330 125.915 48.660 126.715 ;
        RECT 48.960 126.085 49.290 126.885 ;
        RECT 49.460 125.915 49.790 126.715 ;
        RECT 47.355 125.745 49.790 125.915 ;
        RECT 46.485 125.185 46.660 125.745 ;
        RECT 47.355 125.495 47.525 125.745 ;
        RECT 46.830 125.325 47.525 125.495 ;
        RECT 47.700 125.325 48.120 125.525 ;
        RECT 48.290 125.325 48.620 125.525 ;
        RECT 48.790 125.325 49.120 125.525 ;
        RECT 46.485 125.135 46.715 125.185 ;
        RECT 46.485 124.505 46.825 125.135 ;
        RECT 46.995 124.335 47.245 125.135 ;
        RECT 47.435 124.985 48.660 125.155 ;
        RECT 47.435 124.505 47.765 124.985 ;
        RECT 47.935 124.335 48.160 124.795 ;
        RECT 48.330 124.505 48.660 124.985 ;
        RECT 49.290 125.115 49.460 125.745 ;
        RECT 50.165 125.720 50.455 126.885 ;
        RECT 50.625 125.745 50.965 126.715 ;
        RECT 51.135 125.745 51.305 126.885 ;
        RECT 51.575 126.085 51.825 126.885 ;
        RECT 52.470 125.915 52.800 126.715 ;
        RECT 53.100 126.085 53.430 126.885 ;
        RECT 53.600 125.915 53.930 126.715 ;
        RECT 51.495 125.745 53.930 125.915 ;
        RECT 54.305 126.125 54.820 126.535 ;
        RECT 55.055 126.125 55.225 126.885 ;
        RECT 55.395 126.545 57.425 126.715 ;
        RECT 49.645 125.325 49.995 125.575 ;
        RECT 50.625 125.185 50.800 125.745 ;
        RECT 51.495 125.495 51.665 125.745 ;
        RECT 50.970 125.325 51.665 125.495 ;
        RECT 51.840 125.325 52.260 125.525 ;
        RECT 52.430 125.325 52.760 125.525 ;
        RECT 52.930 125.325 53.260 125.525 ;
        RECT 50.625 125.135 50.855 125.185 ;
        RECT 49.290 124.505 49.790 125.115 ;
        RECT 50.165 124.335 50.455 125.060 ;
        RECT 50.625 124.505 50.965 125.135 ;
        RECT 51.135 124.335 51.385 125.135 ;
        RECT 51.575 124.985 52.800 125.155 ;
        RECT 51.575 124.505 51.905 124.985 ;
        RECT 52.075 124.335 52.300 124.795 ;
        RECT 52.470 124.505 52.800 124.985 ;
        RECT 53.430 125.115 53.600 125.745 ;
        RECT 53.785 125.325 54.135 125.575 ;
        RECT 54.305 125.315 54.645 126.125 ;
        RECT 55.395 125.880 55.565 126.545 ;
        RECT 55.960 126.205 57.085 126.375 ;
        RECT 54.815 125.690 55.565 125.880 ;
        RECT 55.735 125.865 56.745 126.035 ;
        RECT 54.305 125.145 55.535 125.315 ;
        RECT 53.430 124.505 53.930 125.115 ;
        RECT 54.580 124.540 54.825 125.145 ;
        RECT 55.045 124.335 55.555 124.870 ;
        RECT 55.735 124.505 55.925 125.865 ;
        RECT 56.095 125.525 56.370 125.665 ;
        RECT 56.095 125.355 56.375 125.525 ;
        RECT 56.095 124.505 56.370 125.355 ;
        RECT 56.575 125.065 56.745 125.865 ;
        RECT 56.915 125.075 57.085 126.205 ;
        RECT 57.255 125.575 57.425 126.545 ;
        RECT 57.595 125.745 57.765 126.885 ;
        RECT 57.935 125.745 58.270 126.715 ;
        RECT 57.255 125.245 57.450 125.575 ;
        RECT 57.675 125.245 57.930 125.575 ;
        RECT 57.675 125.075 57.845 125.245 ;
        RECT 58.100 125.075 58.270 125.745 ;
        RECT 58.820 125.905 59.075 126.575 ;
        RECT 59.255 126.085 59.540 126.885 ;
        RECT 59.720 126.165 60.050 126.675 ;
        RECT 58.820 125.185 59.000 125.905 ;
        RECT 59.720 125.575 59.970 126.165 ;
        RECT 60.320 126.015 60.490 126.625 ;
        RECT 60.660 126.195 60.990 126.885 ;
        RECT 61.220 126.335 61.460 126.625 ;
        RECT 61.660 126.505 62.080 126.885 ;
        RECT 62.260 126.415 62.890 126.665 ;
        RECT 63.360 126.505 63.690 126.885 ;
        RECT 62.260 126.335 62.430 126.415 ;
        RECT 63.860 126.335 64.030 126.625 ;
        RECT 64.210 126.505 64.590 126.885 ;
        RECT 64.830 126.500 65.660 126.670 ;
        RECT 61.220 126.165 62.430 126.335 ;
        RECT 59.170 125.245 59.970 125.575 ;
        RECT 56.915 124.905 57.845 125.075 ;
        RECT 56.915 124.870 57.090 124.905 ;
        RECT 56.560 124.505 57.090 124.870 ;
        RECT 57.515 124.335 57.845 124.735 ;
        RECT 58.015 124.505 58.270 125.075 ;
        RECT 58.735 125.045 59.000 125.185 ;
        RECT 58.735 125.015 59.075 125.045 ;
        RECT 58.820 124.515 59.075 125.015 ;
        RECT 59.255 124.335 59.540 124.795 ;
        RECT 59.720 124.595 59.970 125.245 ;
        RECT 60.170 125.995 60.490 126.015 ;
        RECT 60.170 125.825 62.090 125.995 ;
        RECT 60.170 124.930 60.360 125.825 ;
        RECT 62.260 125.655 62.430 126.165 ;
        RECT 62.600 125.905 63.120 126.215 ;
        RECT 60.530 125.485 62.430 125.655 ;
        RECT 60.530 125.425 60.860 125.485 ;
        RECT 61.010 125.255 61.340 125.315 ;
        RECT 60.680 124.985 61.340 125.255 ;
        RECT 60.170 124.600 60.490 124.930 ;
        RECT 60.670 124.335 61.330 124.815 ;
        RECT 61.530 124.725 61.700 125.485 ;
        RECT 62.600 125.315 62.780 125.725 ;
        RECT 61.870 125.145 62.200 125.265 ;
        RECT 62.950 125.145 63.120 125.905 ;
        RECT 61.870 124.975 63.120 125.145 ;
        RECT 63.290 126.085 64.660 126.335 ;
        RECT 63.290 125.315 63.480 126.085 ;
        RECT 64.410 125.825 64.660 126.085 ;
        RECT 63.650 125.655 63.900 125.815 ;
        RECT 64.830 125.655 65.000 126.500 ;
        RECT 65.895 126.215 66.065 126.715 ;
        RECT 66.235 126.385 66.565 126.885 ;
        RECT 65.170 125.825 65.670 126.205 ;
        RECT 65.895 126.045 66.590 126.215 ;
        RECT 63.650 125.485 65.000 125.655 ;
        RECT 64.580 125.445 65.000 125.485 ;
        RECT 63.290 124.975 63.710 125.315 ;
        RECT 64.000 124.985 64.410 125.315 ;
        RECT 61.530 124.555 62.380 124.725 ;
        RECT 62.940 124.335 63.260 124.795 ;
        RECT 63.460 124.545 63.710 124.975 ;
        RECT 64.000 124.335 64.410 124.775 ;
        RECT 64.580 124.715 64.750 125.445 ;
        RECT 64.920 124.895 65.270 125.265 ;
        RECT 65.450 124.955 65.670 125.825 ;
        RECT 65.840 125.255 66.250 125.875 ;
        RECT 66.420 125.075 66.590 126.045 ;
        RECT 65.895 124.885 66.590 125.075 ;
        RECT 64.580 124.515 65.595 124.715 ;
        RECT 65.895 124.555 66.065 124.885 ;
        RECT 66.235 124.335 66.565 124.715 ;
        RECT 66.780 124.595 67.005 126.715 ;
        RECT 67.175 126.385 67.505 126.885 ;
        RECT 67.675 126.215 67.845 126.715 ;
        RECT 67.180 126.045 67.845 126.215 ;
        RECT 67.180 125.055 67.410 126.045 ;
        RECT 67.580 125.225 67.930 125.875 ;
        RECT 68.565 125.795 70.235 126.885 ;
        RECT 70.410 126.450 75.755 126.885 ;
        RECT 68.565 125.275 69.315 125.795 ;
        RECT 69.485 125.105 70.235 125.625 ;
        RECT 72.000 125.200 72.350 126.450 ;
        RECT 75.925 125.720 76.215 126.885 ;
        RECT 77.505 126.215 77.785 126.885 ;
        RECT 77.955 125.995 78.255 126.545 ;
        RECT 78.455 126.165 78.785 126.885 ;
        RECT 78.975 126.165 79.435 126.715 ;
        RECT 67.180 124.885 67.845 125.055 ;
        RECT 67.175 124.335 67.505 124.715 ;
        RECT 67.675 124.595 67.845 124.885 ;
        RECT 68.565 124.335 70.235 125.105 ;
        RECT 73.830 124.880 74.170 125.710 ;
        RECT 77.320 125.575 77.585 125.935 ;
        RECT 77.955 125.825 78.895 125.995 ;
        RECT 78.725 125.575 78.895 125.825 ;
        RECT 77.320 125.325 77.995 125.575 ;
        RECT 78.215 125.325 78.555 125.575 ;
        RECT 78.725 125.245 79.015 125.575 ;
        RECT 78.725 125.155 78.895 125.245 ;
        RECT 70.410 124.335 75.755 124.880 ;
        RECT 75.925 124.335 76.215 125.060 ;
        RECT 77.505 124.965 78.895 125.155 ;
        RECT 77.505 124.605 77.835 124.965 ;
        RECT 79.185 124.795 79.435 126.165 ;
        RECT 79.605 125.795 81.275 126.885 ;
        RECT 81.445 126.125 81.960 126.535 ;
        RECT 82.195 126.125 82.365 126.885 ;
        RECT 82.535 126.545 84.565 126.715 ;
        RECT 79.605 125.275 80.355 125.795 ;
        RECT 80.525 125.105 81.275 125.625 ;
        RECT 81.445 125.315 81.785 126.125 ;
        RECT 82.535 125.880 82.705 126.545 ;
        RECT 83.100 126.205 84.225 126.375 ;
        RECT 81.955 125.690 82.705 125.880 ;
        RECT 82.875 125.865 83.885 126.035 ;
        RECT 81.445 125.145 82.675 125.315 ;
        RECT 78.455 124.335 78.705 124.795 ;
        RECT 78.875 124.505 79.435 124.795 ;
        RECT 79.605 124.335 81.275 125.105 ;
        RECT 81.720 124.540 81.965 125.145 ;
        RECT 82.185 124.335 82.695 124.870 ;
        RECT 82.875 124.505 83.065 125.865 ;
        RECT 83.235 124.845 83.510 125.665 ;
        RECT 83.715 125.065 83.885 125.865 ;
        RECT 84.055 125.075 84.225 126.205 ;
        RECT 84.395 125.575 84.565 126.545 ;
        RECT 84.735 125.745 84.905 126.885 ;
        RECT 85.075 125.745 85.410 126.715 ;
        RECT 84.395 125.245 84.590 125.575 ;
        RECT 84.815 125.245 85.070 125.575 ;
        RECT 84.815 125.075 84.985 125.245 ;
        RECT 85.240 125.075 85.410 125.745 ;
        RECT 84.055 124.905 84.985 125.075 ;
        RECT 84.055 124.870 84.230 124.905 ;
        RECT 83.235 124.675 83.515 124.845 ;
        RECT 83.235 124.505 83.510 124.675 ;
        RECT 83.700 124.505 84.230 124.870 ;
        RECT 84.655 124.335 84.985 124.735 ;
        RECT 85.155 124.505 85.410 125.075 ;
        RECT 85.585 126.165 86.045 126.715 ;
        RECT 86.235 126.165 86.565 126.885 ;
        RECT 85.585 124.795 85.835 126.165 ;
        RECT 86.765 125.995 87.065 126.545 ;
        RECT 87.235 126.215 87.515 126.885 ;
        RECT 86.125 125.825 87.065 125.995 ;
        RECT 86.125 125.575 86.295 125.825 ;
        RECT 87.435 125.575 87.700 125.935 ;
        RECT 86.005 125.245 86.295 125.575 ;
        RECT 86.465 125.325 86.805 125.575 ;
        RECT 87.025 125.325 87.700 125.575 ;
        RECT 88.345 125.795 91.855 126.885 ;
        RECT 92.030 126.450 97.375 126.885 ;
        RECT 88.345 125.275 90.035 125.795 ;
        RECT 86.125 125.155 86.295 125.245 ;
        RECT 86.125 124.965 87.515 125.155 ;
        RECT 90.205 125.105 91.855 125.625 ;
        RECT 93.620 125.200 93.970 126.450 ;
        RECT 97.545 126.125 98.060 126.535 ;
        RECT 98.295 126.125 98.465 126.885 ;
        RECT 98.635 126.545 100.665 126.715 ;
        RECT 85.585 124.505 86.145 124.795 ;
        RECT 86.315 124.335 86.565 124.795 ;
        RECT 87.185 124.605 87.515 124.965 ;
        RECT 88.345 124.335 91.855 125.105 ;
        RECT 95.450 124.880 95.790 125.710 ;
        RECT 97.545 125.315 97.885 126.125 ;
        RECT 98.635 125.880 98.805 126.545 ;
        RECT 99.200 126.205 100.325 126.375 ;
        RECT 98.055 125.690 98.805 125.880 ;
        RECT 98.975 125.865 99.985 126.035 ;
        RECT 97.545 125.145 98.775 125.315 ;
        RECT 92.030 124.335 97.375 124.880 ;
        RECT 97.820 124.540 98.065 125.145 ;
        RECT 98.285 124.335 98.795 124.870 ;
        RECT 98.975 124.505 99.165 125.865 ;
        RECT 99.335 124.845 99.610 125.665 ;
        RECT 99.815 125.065 99.985 125.865 ;
        RECT 100.155 125.075 100.325 126.205 ;
        RECT 100.495 125.575 100.665 126.545 ;
        RECT 100.835 125.745 101.005 126.885 ;
        RECT 101.175 125.745 101.510 126.715 ;
        RECT 100.495 125.245 100.690 125.575 ;
        RECT 100.915 125.245 101.170 125.575 ;
        RECT 100.915 125.075 101.085 125.245 ;
        RECT 101.340 125.075 101.510 125.745 ;
        RECT 101.685 125.720 101.975 126.885 ;
        RECT 102.145 125.795 103.815 126.885 ;
        RECT 102.145 125.275 102.895 125.795 ;
        RECT 104.025 125.745 104.255 126.885 ;
        RECT 104.425 125.735 104.755 126.715 ;
        RECT 104.925 125.745 105.135 126.885 ;
        RECT 105.365 126.125 105.880 126.535 ;
        RECT 106.115 126.125 106.285 126.885 ;
        RECT 106.455 126.545 108.485 126.715 ;
        RECT 103.065 125.105 103.815 125.625 ;
        RECT 104.005 125.325 104.335 125.575 ;
        RECT 100.155 124.905 101.085 125.075 ;
        RECT 100.155 124.870 100.330 124.905 ;
        RECT 99.335 124.675 99.615 124.845 ;
        RECT 99.335 124.505 99.610 124.675 ;
        RECT 99.800 124.505 100.330 124.870 ;
        RECT 100.755 124.335 101.085 124.735 ;
        RECT 101.255 124.505 101.510 125.075 ;
        RECT 101.685 124.335 101.975 125.060 ;
        RECT 102.145 124.335 103.815 125.105 ;
        RECT 104.025 124.335 104.255 125.155 ;
        RECT 104.505 125.135 104.755 125.735 ;
        RECT 105.365 125.315 105.705 126.125 ;
        RECT 106.455 125.880 106.625 126.545 ;
        RECT 107.020 126.205 108.145 126.375 ;
        RECT 105.875 125.690 106.625 125.880 ;
        RECT 106.795 125.865 107.805 126.035 ;
        RECT 104.425 124.505 104.755 125.135 ;
        RECT 104.925 124.335 105.135 125.155 ;
        RECT 105.365 125.145 106.595 125.315 ;
        RECT 105.640 124.540 105.885 125.145 ;
        RECT 106.105 124.335 106.615 124.870 ;
        RECT 106.795 124.505 106.985 125.865 ;
        RECT 107.155 124.845 107.430 125.665 ;
        RECT 107.635 125.065 107.805 125.865 ;
        RECT 107.975 125.075 108.145 126.205 ;
        RECT 108.315 125.575 108.485 126.545 ;
        RECT 108.655 125.745 108.825 126.885 ;
        RECT 108.995 125.745 109.330 126.715 ;
        RECT 108.315 125.245 108.510 125.575 ;
        RECT 108.735 125.245 108.990 125.575 ;
        RECT 108.735 125.075 108.905 125.245 ;
        RECT 109.160 125.075 109.330 125.745 ;
        RECT 109.965 125.795 112.555 126.885 ;
        RECT 109.965 125.275 111.175 125.795 ;
        RECT 112.765 125.745 112.995 126.885 ;
        RECT 113.165 125.735 113.495 126.715 ;
        RECT 113.665 125.745 113.875 126.885 ;
        RECT 114.480 125.905 114.735 126.575 ;
        RECT 114.915 126.085 115.200 126.885 ;
        RECT 115.380 126.165 115.710 126.675 ;
        RECT 114.480 125.865 114.660 125.905 ;
        RECT 111.345 125.105 112.555 125.625 ;
        RECT 112.745 125.325 113.075 125.575 ;
        RECT 107.975 124.905 108.905 125.075 ;
        RECT 107.975 124.870 108.150 124.905 ;
        RECT 107.155 124.675 107.435 124.845 ;
        RECT 107.155 124.505 107.430 124.675 ;
        RECT 107.620 124.505 108.150 124.870 ;
        RECT 108.575 124.335 108.905 124.735 ;
        RECT 109.075 124.505 109.330 125.075 ;
        RECT 109.965 124.335 112.555 125.105 ;
        RECT 112.765 124.335 112.995 125.155 ;
        RECT 113.245 125.135 113.495 125.735 ;
        RECT 114.395 125.695 114.660 125.865 ;
        RECT 113.165 124.505 113.495 125.135 ;
        RECT 113.665 124.335 113.875 125.155 ;
        RECT 114.480 125.045 114.660 125.695 ;
        RECT 115.380 125.575 115.630 126.165 ;
        RECT 115.980 126.015 116.150 126.625 ;
        RECT 116.320 126.195 116.650 126.885 ;
        RECT 116.880 126.335 117.120 126.625 ;
        RECT 117.320 126.505 117.740 126.885 ;
        RECT 117.920 126.415 118.550 126.665 ;
        RECT 119.020 126.505 119.350 126.885 ;
        RECT 117.920 126.335 118.090 126.415 ;
        RECT 119.520 126.335 119.690 126.625 ;
        RECT 119.870 126.505 120.250 126.885 ;
        RECT 120.490 126.500 121.320 126.670 ;
        RECT 116.880 126.165 118.090 126.335 ;
        RECT 114.830 125.245 115.630 125.575 ;
        RECT 114.480 124.515 114.735 125.045 ;
        RECT 114.915 124.335 115.200 124.795 ;
        RECT 115.380 124.595 115.630 125.245 ;
        RECT 115.830 125.995 116.150 126.015 ;
        RECT 115.830 125.825 117.750 125.995 ;
        RECT 115.830 124.930 116.020 125.825 ;
        RECT 117.920 125.655 118.090 126.165 ;
        RECT 118.260 125.905 118.780 126.215 ;
        RECT 116.190 125.485 118.090 125.655 ;
        RECT 116.190 125.425 116.520 125.485 ;
        RECT 116.670 125.255 117.000 125.315 ;
        RECT 116.340 124.985 117.000 125.255 ;
        RECT 115.830 124.600 116.150 124.930 ;
        RECT 116.330 124.335 116.990 124.815 ;
        RECT 117.190 124.725 117.360 125.485 ;
        RECT 118.260 125.315 118.440 125.725 ;
        RECT 117.530 125.145 117.860 125.265 ;
        RECT 118.610 125.145 118.780 125.905 ;
        RECT 117.530 124.975 118.780 125.145 ;
        RECT 118.950 126.085 120.320 126.335 ;
        RECT 118.950 125.315 119.140 126.085 ;
        RECT 120.070 125.825 120.320 126.085 ;
        RECT 119.310 125.655 119.560 125.815 ;
        RECT 120.490 125.655 120.660 126.500 ;
        RECT 121.555 126.215 121.725 126.715 ;
        RECT 121.895 126.385 122.225 126.885 ;
        RECT 120.830 125.825 121.330 126.205 ;
        RECT 121.555 126.045 122.250 126.215 ;
        RECT 119.310 125.485 120.660 125.655 ;
        RECT 120.240 125.445 120.660 125.485 ;
        RECT 118.950 124.975 119.370 125.315 ;
        RECT 119.660 124.985 120.070 125.315 ;
        RECT 117.190 124.555 118.040 124.725 ;
        RECT 118.600 124.335 118.920 124.795 ;
        RECT 119.120 124.545 119.370 124.975 ;
        RECT 119.660 124.335 120.070 124.775 ;
        RECT 120.240 124.715 120.410 125.445 ;
        RECT 120.580 124.895 120.930 125.265 ;
        RECT 121.110 124.955 121.330 125.825 ;
        RECT 121.500 125.255 121.910 125.875 ;
        RECT 122.080 125.075 122.250 126.045 ;
        RECT 121.555 124.885 122.250 125.075 ;
        RECT 120.240 124.515 121.255 124.715 ;
        RECT 121.555 124.555 121.725 124.885 ;
        RECT 121.895 124.335 122.225 124.715 ;
        RECT 122.440 124.595 122.665 126.715 ;
        RECT 122.835 126.385 123.165 126.885 ;
        RECT 123.335 126.215 123.505 126.715 ;
        RECT 122.840 126.045 123.505 126.215 ;
        RECT 122.840 125.055 123.070 126.045 ;
        RECT 123.240 125.225 123.590 125.875 ;
        RECT 123.765 125.795 126.355 126.885 ;
        RECT 126.525 125.795 127.735 126.885 ;
        RECT 123.765 125.275 124.975 125.795 ;
        RECT 125.145 125.105 126.355 125.625 ;
        RECT 126.525 125.255 127.045 125.795 ;
        RECT 122.840 124.885 123.505 125.055 ;
        RECT 122.835 124.335 123.165 124.715 ;
        RECT 123.335 124.595 123.505 124.885 ;
        RECT 123.765 124.335 126.355 125.105 ;
        RECT 127.215 125.085 127.735 125.625 ;
        RECT 126.525 124.335 127.735 125.085 ;
        RECT 14.660 124.165 127.820 124.335 ;
        RECT 14.745 123.415 15.955 124.165 ;
        RECT 16.590 123.620 21.935 124.165 ;
        RECT 14.745 122.875 15.265 123.415 ;
        RECT 15.435 122.705 15.955 123.245 ;
        RECT 14.745 121.615 15.955 122.705 ;
        RECT 18.180 122.050 18.530 123.300 ;
        RECT 20.010 122.790 20.350 123.620 ;
        RECT 22.195 123.615 22.365 123.995 ;
        RECT 22.545 123.785 22.875 124.165 ;
        RECT 22.195 123.445 22.860 123.615 ;
        RECT 23.055 123.490 23.315 123.995 ;
        RECT 22.125 122.895 22.455 123.265 ;
        RECT 22.690 123.190 22.860 123.445 ;
        RECT 22.690 122.860 22.975 123.190 ;
        RECT 22.690 122.715 22.860 122.860 ;
        RECT 22.195 122.545 22.860 122.715 ;
        RECT 23.145 122.690 23.315 123.490 ;
        RECT 16.590 121.615 21.935 122.050 ;
        RECT 22.195 121.785 22.365 122.545 ;
        RECT 22.545 121.615 22.875 122.375 ;
        RECT 23.045 121.785 23.315 122.690 ;
        RECT 23.860 123.455 24.115 123.985 ;
        RECT 24.295 123.705 24.580 124.165 ;
        RECT 23.860 122.595 24.040 123.455 ;
        RECT 24.760 123.255 25.010 123.905 ;
        RECT 24.210 122.925 25.010 123.255 ;
        RECT 23.860 122.125 24.115 122.595 ;
        RECT 23.775 121.955 24.115 122.125 ;
        RECT 23.860 121.925 24.115 121.955 ;
        RECT 24.295 121.615 24.580 122.415 ;
        RECT 24.760 122.335 25.010 122.925 ;
        RECT 25.210 123.570 25.530 123.900 ;
        RECT 25.710 123.685 26.370 124.165 ;
        RECT 26.570 123.775 27.420 123.945 ;
        RECT 25.210 122.675 25.400 123.570 ;
        RECT 25.720 123.245 26.380 123.515 ;
        RECT 26.050 123.185 26.380 123.245 ;
        RECT 25.570 123.015 25.900 123.075 ;
        RECT 26.570 123.015 26.740 123.775 ;
        RECT 27.980 123.705 28.300 124.165 ;
        RECT 28.500 123.525 28.750 123.955 ;
        RECT 29.040 123.725 29.450 124.165 ;
        RECT 29.620 123.785 30.635 123.985 ;
        RECT 26.910 123.355 28.160 123.525 ;
        RECT 26.910 123.235 27.240 123.355 ;
        RECT 25.570 122.845 27.470 123.015 ;
        RECT 25.210 122.505 27.130 122.675 ;
        RECT 25.210 122.485 25.530 122.505 ;
        RECT 24.760 121.825 25.090 122.335 ;
        RECT 25.360 121.875 25.530 122.485 ;
        RECT 27.300 122.335 27.470 122.845 ;
        RECT 27.640 122.775 27.820 123.185 ;
        RECT 27.990 122.595 28.160 123.355 ;
        RECT 25.700 121.615 26.030 122.305 ;
        RECT 26.260 122.165 27.470 122.335 ;
        RECT 27.640 122.285 28.160 122.595 ;
        RECT 28.330 123.185 28.750 123.525 ;
        RECT 29.040 123.185 29.450 123.515 ;
        RECT 28.330 122.415 28.520 123.185 ;
        RECT 29.620 123.055 29.790 123.785 ;
        RECT 30.935 123.615 31.105 123.945 ;
        RECT 31.275 123.785 31.605 124.165 ;
        RECT 29.960 123.235 30.310 123.605 ;
        RECT 29.620 123.015 30.040 123.055 ;
        RECT 28.690 122.845 30.040 123.015 ;
        RECT 28.690 122.685 28.940 122.845 ;
        RECT 29.450 122.415 29.700 122.675 ;
        RECT 28.330 122.165 29.700 122.415 ;
        RECT 26.260 121.875 26.500 122.165 ;
        RECT 27.300 122.085 27.470 122.165 ;
        RECT 26.700 121.615 27.120 121.995 ;
        RECT 27.300 121.835 27.930 122.085 ;
        RECT 28.400 121.615 28.730 121.995 ;
        RECT 28.900 121.875 29.070 122.165 ;
        RECT 29.870 122.000 30.040 122.845 ;
        RECT 30.490 122.675 30.710 123.545 ;
        RECT 30.935 123.425 31.630 123.615 ;
        RECT 30.210 122.295 30.710 122.675 ;
        RECT 30.880 122.625 31.290 123.245 ;
        RECT 31.460 122.455 31.630 123.425 ;
        RECT 30.935 122.285 31.630 122.455 ;
        RECT 29.250 121.615 29.630 121.995 ;
        RECT 29.870 121.830 30.700 122.000 ;
        RECT 30.935 121.785 31.105 122.285 ;
        RECT 31.275 121.615 31.605 122.115 ;
        RECT 31.820 121.785 32.045 123.905 ;
        RECT 32.215 123.785 32.545 124.165 ;
        RECT 32.715 123.615 32.885 123.905 ;
        RECT 32.220 123.445 32.885 123.615 ;
        RECT 32.220 122.455 32.450 123.445 ;
        RECT 33.150 123.425 33.405 123.995 ;
        RECT 33.575 123.765 33.905 124.165 ;
        RECT 34.330 123.630 34.860 123.995 ;
        RECT 34.330 123.595 34.505 123.630 ;
        RECT 33.575 123.425 34.505 123.595 ;
        RECT 32.620 122.625 32.970 123.275 ;
        RECT 33.150 122.755 33.320 123.425 ;
        RECT 33.575 123.255 33.745 123.425 ;
        RECT 33.490 122.925 33.745 123.255 ;
        RECT 33.970 122.925 34.165 123.255 ;
        RECT 32.220 122.285 32.885 122.455 ;
        RECT 32.215 121.615 32.545 122.115 ;
        RECT 32.715 121.785 32.885 122.285 ;
        RECT 33.150 121.785 33.485 122.755 ;
        RECT 33.655 121.615 33.825 122.755 ;
        RECT 33.995 121.955 34.165 122.925 ;
        RECT 34.335 122.295 34.505 123.425 ;
        RECT 34.675 122.635 34.845 123.435 ;
        RECT 35.050 123.145 35.325 123.995 ;
        RECT 35.045 122.975 35.325 123.145 ;
        RECT 35.050 122.835 35.325 122.975 ;
        RECT 35.495 122.635 35.685 123.995 ;
        RECT 35.865 123.630 36.375 124.165 ;
        RECT 36.595 123.355 36.840 123.960 ;
        RECT 37.285 123.440 37.575 124.165 ;
        RECT 37.945 123.535 38.275 123.895 ;
        RECT 38.895 123.705 39.145 124.165 ;
        RECT 39.315 123.705 39.875 123.995 ;
        RECT 35.885 123.185 37.115 123.355 ;
        RECT 37.945 123.345 39.335 123.535 ;
        RECT 34.675 122.465 35.685 122.635 ;
        RECT 35.855 122.620 36.605 122.810 ;
        RECT 34.335 122.125 35.460 122.295 ;
        RECT 35.855 121.955 36.025 122.620 ;
        RECT 36.775 122.375 37.115 123.185 ;
        RECT 39.165 123.255 39.335 123.345 ;
        RECT 37.760 122.925 38.435 123.175 ;
        RECT 38.655 122.925 38.995 123.175 ;
        RECT 39.165 122.925 39.455 123.255 ;
        RECT 33.995 121.785 36.025 121.955 ;
        RECT 36.195 121.615 36.365 122.375 ;
        RECT 36.600 121.965 37.115 122.375 ;
        RECT 37.285 121.615 37.575 122.780 ;
        RECT 37.760 122.565 38.025 122.925 ;
        RECT 39.165 122.675 39.335 122.925 ;
        RECT 38.395 122.505 39.335 122.675 ;
        RECT 37.945 121.615 38.225 122.285 ;
        RECT 38.395 121.955 38.695 122.505 ;
        RECT 39.625 122.335 39.875 123.705 ;
        RECT 40.245 123.535 40.575 123.895 ;
        RECT 41.195 123.705 41.445 124.165 ;
        RECT 41.615 123.705 42.175 123.995 ;
        RECT 40.245 123.345 41.635 123.535 ;
        RECT 41.465 123.255 41.635 123.345 ;
        RECT 40.060 122.925 40.735 123.175 ;
        RECT 40.955 122.925 41.295 123.175 ;
        RECT 41.465 122.925 41.755 123.255 ;
        RECT 40.060 122.565 40.325 122.925 ;
        RECT 41.465 122.675 41.635 122.925 ;
        RECT 38.895 121.615 39.225 122.335 ;
        RECT 39.415 121.785 39.875 122.335 ;
        RECT 40.695 122.505 41.635 122.675 ;
        RECT 40.245 121.615 40.525 122.285 ;
        RECT 40.695 121.955 40.995 122.505 ;
        RECT 41.925 122.335 42.175 123.705 ;
        RECT 42.545 123.535 42.875 123.895 ;
        RECT 43.495 123.705 43.745 124.165 ;
        RECT 43.915 123.705 44.475 123.995 ;
        RECT 42.545 123.345 43.935 123.535 ;
        RECT 43.765 123.255 43.935 123.345 ;
        RECT 42.360 122.925 43.035 123.175 ;
        RECT 43.255 122.925 43.595 123.175 ;
        RECT 43.765 122.925 44.055 123.255 ;
        RECT 42.360 122.565 42.625 122.925 ;
        RECT 43.765 122.675 43.935 122.925 ;
        RECT 41.195 121.615 41.525 122.335 ;
        RECT 41.715 121.785 42.175 122.335 ;
        RECT 42.995 122.505 43.935 122.675 ;
        RECT 42.545 121.615 42.825 122.285 ;
        RECT 42.995 121.955 43.295 122.505 ;
        RECT 44.225 122.335 44.475 123.705 ;
        RECT 44.845 123.535 45.175 123.895 ;
        RECT 45.795 123.705 46.045 124.165 ;
        RECT 46.215 123.705 46.775 123.995 ;
        RECT 44.845 123.345 46.235 123.535 ;
        RECT 46.065 123.255 46.235 123.345 ;
        RECT 44.660 122.925 45.335 123.175 ;
        RECT 45.555 122.925 45.895 123.175 ;
        RECT 46.065 122.925 46.355 123.255 ;
        RECT 44.660 122.565 44.925 122.925 ;
        RECT 46.065 122.675 46.235 122.925 ;
        RECT 43.495 121.615 43.825 122.335 ;
        RECT 44.015 121.785 44.475 122.335 ;
        RECT 45.295 122.505 46.235 122.675 ;
        RECT 44.845 121.615 45.125 122.285 ;
        RECT 45.295 121.955 45.595 122.505 ;
        RECT 46.525 122.335 46.775 123.705 ;
        RECT 47.495 123.685 47.795 124.165 ;
        RECT 47.965 123.515 48.225 123.970 ;
        RECT 48.395 123.685 48.655 124.165 ;
        RECT 48.835 123.515 49.095 123.970 ;
        RECT 49.265 123.685 49.515 124.165 ;
        RECT 49.695 123.515 49.955 123.970 ;
        RECT 50.125 123.685 50.375 124.165 ;
        RECT 50.555 123.515 50.815 123.970 ;
        RECT 50.985 123.685 51.230 124.165 ;
        RECT 51.400 123.515 51.675 123.970 ;
        RECT 51.845 123.685 52.090 124.165 ;
        RECT 52.260 123.515 52.520 123.970 ;
        RECT 52.690 123.685 52.950 124.165 ;
        RECT 53.120 123.515 53.380 123.970 ;
        RECT 53.550 123.685 53.810 124.165 ;
        RECT 53.980 123.515 54.240 123.970 ;
        RECT 54.410 123.605 54.670 124.165 ;
        RECT 47.495 123.345 54.240 123.515 ;
        RECT 47.495 122.755 48.660 123.345 ;
        RECT 54.840 123.175 55.090 123.985 ;
        RECT 55.270 123.640 55.530 124.165 ;
        RECT 55.700 123.175 55.950 123.985 ;
        RECT 56.130 123.655 56.435 124.165 ;
        RECT 48.830 122.925 55.950 123.175 ;
        RECT 56.120 122.925 56.435 123.485 ;
        RECT 57.525 123.395 61.035 124.165 ;
        RECT 47.495 122.530 54.240 122.755 ;
        RECT 45.795 121.615 46.125 122.335 ;
        RECT 46.315 121.785 46.775 122.335 ;
        RECT 47.495 121.615 47.765 122.360 ;
        RECT 47.935 121.790 48.225 122.530 ;
        RECT 48.835 122.515 54.240 122.530 ;
        RECT 48.395 121.620 48.650 122.345 ;
        RECT 48.835 121.790 49.095 122.515 ;
        RECT 49.265 121.620 49.510 122.345 ;
        RECT 49.695 121.790 49.955 122.515 ;
        RECT 50.125 121.620 50.370 122.345 ;
        RECT 50.555 121.790 50.815 122.515 ;
        RECT 50.985 121.620 51.230 122.345 ;
        RECT 51.400 121.790 51.660 122.515 ;
        RECT 51.830 121.620 52.090 122.345 ;
        RECT 52.260 121.790 52.520 122.515 ;
        RECT 52.690 121.620 52.950 122.345 ;
        RECT 53.120 121.790 53.380 122.515 ;
        RECT 53.550 121.620 53.810 122.345 ;
        RECT 53.980 121.790 54.240 122.515 ;
        RECT 54.410 121.620 54.670 122.415 ;
        RECT 54.840 121.790 55.090 122.925 ;
        RECT 48.395 121.615 54.670 121.620 ;
        RECT 55.270 121.615 55.530 122.425 ;
        RECT 55.705 121.785 55.950 122.925 ;
        RECT 57.525 122.705 59.215 123.225 ;
        RECT 59.385 122.875 61.035 123.395 ;
        RECT 61.245 123.345 61.475 124.165 ;
        RECT 61.645 123.365 61.975 123.995 ;
        RECT 61.225 122.925 61.555 123.175 ;
        RECT 61.725 122.765 61.975 123.365 ;
        RECT 62.145 123.345 62.355 124.165 ;
        RECT 63.045 123.440 63.335 124.165 ;
        RECT 64.055 123.615 64.225 123.995 ;
        RECT 64.405 123.785 64.735 124.165 ;
        RECT 64.055 123.445 64.720 123.615 ;
        RECT 64.915 123.490 65.175 123.995 ;
        RECT 63.985 122.895 64.315 123.265 ;
        RECT 64.550 123.190 64.720 123.445 ;
        RECT 64.550 122.860 64.835 123.190 ;
        RECT 56.130 121.615 56.425 122.425 ;
        RECT 57.525 121.615 61.035 122.705 ;
        RECT 61.245 121.615 61.475 122.755 ;
        RECT 61.645 121.785 61.975 122.765 ;
        RECT 62.145 121.615 62.355 122.755 ;
        RECT 63.045 121.615 63.335 122.780 ;
        RECT 64.550 122.715 64.720 122.860 ;
        RECT 64.055 122.545 64.720 122.715 ;
        RECT 65.005 122.690 65.175 123.490 ;
        RECT 65.805 123.395 67.475 124.165 ;
        RECT 67.650 123.620 72.995 124.165 ;
        RECT 64.055 121.785 64.225 122.545 ;
        RECT 64.405 121.615 64.735 122.375 ;
        RECT 64.905 121.785 65.175 122.690 ;
        RECT 65.805 122.705 66.555 123.225 ;
        RECT 66.725 122.875 67.475 123.395 ;
        RECT 65.805 121.615 67.475 122.705 ;
        RECT 69.240 122.050 69.590 123.300 ;
        RECT 71.070 122.790 71.410 123.620 ;
        RECT 73.225 123.345 73.435 124.165 ;
        RECT 73.605 123.365 73.935 123.995 ;
        RECT 73.605 122.765 73.855 123.365 ;
        RECT 74.105 123.345 74.335 124.165 ;
        RECT 75.740 123.355 75.985 123.960 ;
        RECT 76.205 123.630 76.715 124.165 ;
        RECT 75.465 123.185 76.695 123.355 ;
        RECT 74.025 122.925 74.355 123.175 ;
        RECT 67.650 121.615 72.995 122.050 ;
        RECT 73.225 121.615 73.435 122.755 ;
        RECT 73.605 121.785 73.935 122.765 ;
        RECT 74.105 121.615 74.335 122.755 ;
        RECT 75.465 122.375 75.805 123.185 ;
        RECT 75.975 122.620 76.725 122.810 ;
        RECT 75.465 121.965 75.980 122.375 ;
        RECT 76.215 121.615 76.385 122.375 ;
        RECT 76.555 121.955 76.725 122.620 ;
        RECT 76.895 122.635 77.085 123.995 ;
        RECT 77.255 123.145 77.530 123.995 ;
        RECT 77.720 123.630 78.250 123.995 ;
        RECT 78.675 123.765 79.005 124.165 ;
        RECT 78.075 123.595 78.250 123.630 ;
        RECT 77.255 122.975 77.535 123.145 ;
        RECT 77.255 122.835 77.530 122.975 ;
        RECT 77.735 122.635 77.905 123.435 ;
        RECT 76.895 122.465 77.905 122.635 ;
        RECT 78.075 123.425 79.005 123.595 ;
        RECT 79.175 123.425 79.430 123.995 ;
        RECT 79.695 123.685 79.995 124.165 ;
        RECT 80.165 123.515 80.425 123.970 ;
        RECT 80.595 123.685 80.855 124.165 ;
        RECT 81.035 123.515 81.295 123.970 ;
        RECT 81.465 123.685 81.715 124.165 ;
        RECT 81.895 123.515 82.155 123.970 ;
        RECT 82.325 123.685 82.575 124.165 ;
        RECT 82.755 123.515 83.015 123.970 ;
        RECT 83.185 123.685 83.430 124.165 ;
        RECT 83.600 123.515 83.875 123.970 ;
        RECT 84.045 123.685 84.290 124.165 ;
        RECT 84.460 123.515 84.720 123.970 ;
        RECT 84.890 123.685 85.150 124.165 ;
        RECT 85.320 123.515 85.580 123.970 ;
        RECT 85.750 123.685 86.010 124.165 ;
        RECT 86.180 123.515 86.440 123.970 ;
        RECT 86.610 123.605 86.870 124.165 ;
        RECT 78.075 122.295 78.245 123.425 ;
        RECT 78.835 123.255 79.005 123.425 ;
        RECT 77.120 122.125 78.245 122.295 ;
        RECT 78.415 122.925 78.610 123.255 ;
        RECT 78.835 122.925 79.090 123.255 ;
        RECT 78.415 121.955 78.585 122.925 ;
        RECT 79.260 122.755 79.430 123.425 ;
        RECT 76.555 121.785 78.585 121.955 ;
        RECT 78.755 121.615 78.925 122.755 ;
        RECT 79.095 121.785 79.430 122.755 ;
        RECT 79.695 123.345 86.440 123.515 ;
        RECT 79.695 122.755 80.860 123.345 ;
        RECT 87.040 123.175 87.290 123.985 ;
        RECT 87.470 123.640 87.730 124.165 ;
        RECT 87.900 123.175 88.150 123.985 ;
        RECT 88.330 123.655 88.635 124.165 ;
        RECT 81.030 122.925 88.150 123.175 ;
        RECT 88.320 122.925 88.635 123.485 ;
        RECT 88.805 123.440 89.095 124.165 ;
        RECT 89.265 123.395 90.935 124.165 ;
        RECT 79.695 122.530 86.440 122.755 ;
        RECT 79.695 121.615 79.965 122.360 ;
        RECT 80.135 121.790 80.425 122.530 ;
        RECT 81.035 122.515 86.440 122.530 ;
        RECT 80.595 121.620 80.850 122.345 ;
        RECT 81.035 121.790 81.295 122.515 ;
        RECT 81.465 121.620 81.710 122.345 ;
        RECT 81.895 121.790 82.155 122.515 ;
        RECT 82.325 121.620 82.570 122.345 ;
        RECT 82.755 121.790 83.015 122.515 ;
        RECT 83.185 121.620 83.430 122.345 ;
        RECT 83.600 121.790 83.860 122.515 ;
        RECT 84.030 121.620 84.290 122.345 ;
        RECT 84.460 121.790 84.720 122.515 ;
        RECT 84.890 121.620 85.150 122.345 ;
        RECT 85.320 121.790 85.580 122.515 ;
        RECT 85.750 121.620 86.010 122.345 ;
        RECT 86.180 121.790 86.440 122.515 ;
        RECT 86.610 121.620 86.870 122.415 ;
        RECT 87.040 121.790 87.290 122.925 ;
        RECT 80.595 121.615 86.870 121.620 ;
        RECT 87.470 121.615 87.730 122.425 ;
        RECT 87.905 121.785 88.150 122.925 ;
        RECT 88.330 121.615 88.625 122.425 ;
        RECT 88.805 121.615 89.095 122.780 ;
        RECT 89.265 122.705 90.015 123.225 ;
        RECT 90.185 122.875 90.935 123.395 ;
        RECT 91.145 123.345 91.375 124.165 ;
        RECT 91.545 123.365 91.875 123.995 ;
        RECT 91.125 122.925 91.455 123.175 ;
        RECT 91.625 122.765 91.875 123.365 ;
        RECT 92.045 123.345 92.255 124.165 ;
        RECT 92.860 123.455 93.115 123.985 ;
        RECT 93.295 123.705 93.580 124.165 ;
        RECT 89.265 121.615 90.935 122.705 ;
        RECT 91.145 121.615 91.375 122.755 ;
        RECT 91.545 121.785 91.875 122.765 ;
        RECT 92.045 121.615 92.255 122.755 ;
        RECT 92.860 122.595 93.040 123.455 ;
        RECT 93.760 123.255 94.010 123.905 ;
        RECT 93.210 122.925 94.010 123.255 ;
        RECT 92.860 122.125 93.115 122.595 ;
        RECT 92.775 121.955 93.115 122.125 ;
        RECT 92.860 121.925 93.115 121.955 ;
        RECT 93.295 121.615 93.580 122.415 ;
        RECT 93.760 122.335 94.010 122.925 ;
        RECT 94.210 123.570 94.530 123.900 ;
        RECT 94.710 123.685 95.370 124.165 ;
        RECT 95.570 123.775 96.420 123.945 ;
        RECT 94.210 122.675 94.400 123.570 ;
        RECT 94.720 123.245 95.380 123.515 ;
        RECT 95.050 123.185 95.380 123.245 ;
        RECT 94.570 123.015 94.900 123.075 ;
        RECT 95.570 123.015 95.740 123.775 ;
        RECT 96.980 123.705 97.300 124.165 ;
        RECT 97.500 123.525 97.750 123.955 ;
        RECT 98.040 123.725 98.450 124.165 ;
        RECT 98.620 123.785 99.635 123.985 ;
        RECT 95.910 123.355 97.160 123.525 ;
        RECT 95.910 123.235 96.240 123.355 ;
        RECT 94.570 122.845 96.470 123.015 ;
        RECT 94.210 122.505 96.130 122.675 ;
        RECT 94.210 122.485 94.530 122.505 ;
        RECT 93.760 121.825 94.090 122.335 ;
        RECT 94.360 121.875 94.530 122.485 ;
        RECT 96.300 122.335 96.470 122.845 ;
        RECT 96.640 122.775 96.820 123.185 ;
        RECT 96.990 122.595 97.160 123.355 ;
        RECT 94.700 121.615 95.030 122.305 ;
        RECT 95.260 122.165 96.470 122.335 ;
        RECT 96.640 122.285 97.160 122.595 ;
        RECT 97.330 123.185 97.750 123.525 ;
        RECT 98.040 123.185 98.450 123.515 ;
        RECT 97.330 122.415 97.520 123.185 ;
        RECT 98.620 123.055 98.790 123.785 ;
        RECT 99.935 123.615 100.105 123.945 ;
        RECT 100.275 123.785 100.605 124.165 ;
        RECT 98.960 123.235 99.310 123.605 ;
        RECT 98.620 123.015 99.040 123.055 ;
        RECT 97.690 122.845 99.040 123.015 ;
        RECT 97.690 122.685 97.940 122.845 ;
        RECT 98.450 122.415 98.700 122.675 ;
        RECT 97.330 122.165 98.700 122.415 ;
        RECT 95.260 121.875 95.500 122.165 ;
        RECT 96.300 122.085 96.470 122.165 ;
        RECT 95.700 121.615 96.120 121.995 ;
        RECT 96.300 121.835 96.930 122.085 ;
        RECT 97.400 121.615 97.730 121.995 ;
        RECT 97.900 121.875 98.070 122.165 ;
        RECT 98.870 122.000 99.040 122.845 ;
        RECT 99.490 122.675 99.710 123.545 ;
        RECT 99.935 123.425 100.630 123.615 ;
        RECT 99.210 122.295 99.710 122.675 ;
        RECT 99.880 122.625 100.290 123.245 ;
        RECT 100.460 122.455 100.630 123.425 ;
        RECT 99.935 122.285 100.630 122.455 ;
        RECT 98.250 121.615 98.630 121.995 ;
        RECT 98.870 121.830 99.700 122.000 ;
        RECT 99.935 121.785 100.105 122.285 ;
        RECT 100.275 121.615 100.605 122.115 ;
        RECT 100.820 121.785 101.045 123.905 ;
        RECT 101.215 123.785 101.545 124.165 ;
        RECT 101.715 123.615 101.885 123.905 ;
        RECT 102.520 123.825 102.775 123.985 ;
        RECT 102.435 123.655 102.775 123.825 ;
        RECT 102.955 123.705 103.240 124.165 ;
        RECT 101.220 123.445 101.885 123.615 ;
        RECT 102.520 123.455 102.775 123.655 ;
        RECT 101.220 122.455 101.450 123.445 ;
        RECT 101.620 122.625 101.970 123.275 ;
        RECT 102.520 122.595 102.700 123.455 ;
        RECT 103.420 123.255 103.670 123.905 ;
        RECT 102.870 122.925 103.670 123.255 ;
        RECT 101.220 122.285 101.885 122.455 ;
        RECT 101.215 121.615 101.545 122.115 ;
        RECT 101.715 121.785 101.885 122.285 ;
        RECT 102.520 121.925 102.775 122.595 ;
        RECT 102.955 121.615 103.240 122.415 ;
        RECT 103.420 122.335 103.670 122.925 ;
        RECT 103.870 123.570 104.190 123.900 ;
        RECT 104.370 123.685 105.030 124.165 ;
        RECT 105.230 123.775 106.080 123.945 ;
        RECT 103.870 122.675 104.060 123.570 ;
        RECT 104.380 123.245 105.040 123.515 ;
        RECT 104.710 123.185 105.040 123.245 ;
        RECT 104.230 123.015 104.560 123.075 ;
        RECT 105.230 123.015 105.400 123.775 ;
        RECT 106.640 123.705 106.960 124.165 ;
        RECT 107.160 123.525 107.410 123.955 ;
        RECT 107.700 123.725 108.110 124.165 ;
        RECT 108.280 123.785 109.295 123.985 ;
        RECT 105.570 123.355 106.820 123.525 ;
        RECT 105.570 123.235 105.900 123.355 ;
        RECT 104.230 122.845 106.130 123.015 ;
        RECT 103.870 122.505 105.790 122.675 ;
        RECT 103.870 122.485 104.190 122.505 ;
        RECT 103.420 121.825 103.750 122.335 ;
        RECT 104.020 121.875 104.190 122.485 ;
        RECT 105.960 122.335 106.130 122.845 ;
        RECT 106.300 122.775 106.480 123.185 ;
        RECT 106.650 122.595 106.820 123.355 ;
        RECT 104.360 121.615 104.690 122.305 ;
        RECT 104.920 122.165 106.130 122.335 ;
        RECT 106.300 122.285 106.820 122.595 ;
        RECT 106.990 123.185 107.410 123.525 ;
        RECT 107.700 123.185 108.110 123.515 ;
        RECT 106.990 122.415 107.180 123.185 ;
        RECT 108.280 123.055 108.450 123.785 ;
        RECT 109.595 123.615 109.765 123.945 ;
        RECT 109.935 123.785 110.265 124.165 ;
        RECT 108.620 123.235 108.970 123.605 ;
        RECT 108.280 123.015 108.700 123.055 ;
        RECT 107.350 122.845 108.700 123.015 ;
        RECT 107.350 122.685 107.600 122.845 ;
        RECT 108.110 122.415 108.360 122.675 ;
        RECT 106.990 122.165 108.360 122.415 ;
        RECT 104.920 121.875 105.160 122.165 ;
        RECT 105.960 122.085 106.130 122.165 ;
        RECT 105.360 121.615 105.780 121.995 ;
        RECT 105.960 121.835 106.590 122.085 ;
        RECT 107.060 121.615 107.390 121.995 ;
        RECT 107.560 121.875 107.730 122.165 ;
        RECT 108.530 122.000 108.700 122.845 ;
        RECT 109.150 122.675 109.370 123.545 ;
        RECT 109.595 123.425 110.290 123.615 ;
        RECT 108.870 122.295 109.370 122.675 ;
        RECT 109.540 122.625 109.950 123.245 ;
        RECT 110.120 122.455 110.290 123.425 ;
        RECT 109.595 122.285 110.290 122.455 ;
        RECT 107.910 121.615 108.290 121.995 ;
        RECT 108.530 121.830 109.360 122.000 ;
        RECT 109.595 121.785 109.765 122.285 ;
        RECT 109.935 121.615 110.265 122.115 ;
        RECT 110.480 121.785 110.705 123.905 ;
        RECT 110.875 123.785 111.205 124.165 ;
        RECT 111.375 123.615 111.545 123.905 ;
        RECT 110.880 123.445 111.545 123.615 ;
        RECT 110.880 122.455 111.110 123.445 ;
        RECT 111.805 123.415 113.015 124.165 ;
        RECT 111.280 122.625 111.630 123.275 ;
        RECT 111.805 122.705 112.325 123.245 ;
        RECT 112.495 122.875 113.015 123.415 ;
        RECT 113.225 123.345 113.455 124.165 ;
        RECT 113.625 123.365 113.955 123.995 ;
        RECT 113.205 122.925 113.535 123.175 ;
        RECT 113.705 122.765 113.955 123.365 ;
        RECT 114.125 123.345 114.335 124.165 ;
        RECT 114.565 123.440 114.855 124.165 ;
        RECT 116.320 123.825 116.575 123.985 ;
        RECT 116.235 123.655 116.575 123.825 ;
        RECT 116.755 123.705 117.040 124.165 ;
        RECT 116.320 123.455 116.575 123.655 ;
        RECT 110.880 122.285 111.545 122.455 ;
        RECT 110.875 121.615 111.205 122.115 ;
        RECT 111.375 121.785 111.545 122.285 ;
        RECT 111.805 121.615 113.015 122.705 ;
        RECT 113.225 121.615 113.455 122.755 ;
        RECT 113.625 121.785 113.955 122.765 ;
        RECT 114.125 121.615 114.335 122.755 ;
        RECT 114.565 121.615 114.855 122.780 ;
        RECT 116.320 122.595 116.500 123.455 ;
        RECT 117.220 123.255 117.470 123.905 ;
        RECT 116.670 122.925 117.470 123.255 ;
        RECT 116.320 121.925 116.575 122.595 ;
        RECT 116.755 121.615 117.040 122.415 ;
        RECT 117.220 122.335 117.470 122.925 ;
        RECT 117.670 123.570 117.990 123.900 ;
        RECT 118.170 123.685 118.830 124.165 ;
        RECT 119.030 123.775 119.880 123.945 ;
        RECT 117.670 122.675 117.860 123.570 ;
        RECT 118.180 123.245 118.840 123.515 ;
        RECT 118.510 123.185 118.840 123.245 ;
        RECT 118.030 123.015 118.360 123.075 ;
        RECT 119.030 123.015 119.200 123.775 ;
        RECT 120.440 123.705 120.760 124.165 ;
        RECT 120.960 123.525 121.210 123.955 ;
        RECT 121.500 123.725 121.910 124.165 ;
        RECT 122.080 123.785 123.095 123.985 ;
        RECT 119.370 123.355 120.620 123.525 ;
        RECT 119.370 123.235 119.700 123.355 ;
        RECT 118.030 122.845 119.930 123.015 ;
        RECT 117.670 122.505 119.590 122.675 ;
        RECT 117.670 122.485 117.990 122.505 ;
        RECT 117.220 121.825 117.550 122.335 ;
        RECT 117.820 121.875 117.990 122.485 ;
        RECT 119.760 122.335 119.930 122.845 ;
        RECT 120.100 122.775 120.280 123.185 ;
        RECT 120.450 122.595 120.620 123.355 ;
        RECT 118.160 121.615 118.490 122.305 ;
        RECT 118.720 122.165 119.930 122.335 ;
        RECT 120.100 122.285 120.620 122.595 ;
        RECT 120.790 123.185 121.210 123.525 ;
        RECT 121.500 123.185 121.910 123.515 ;
        RECT 120.790 122.415 120.980 123.185 ;
        RECT 122.080 123.055 122.250 123.785 ;
        RECT 123.395 123.615 123.565 123.945 ;
        RECT 123.735 123.785 124.065 124.165 ;
        RECT 122.420 123.235 122.770 123.605 ;
        RECT 122.080 123.015 122.500 123.055 ;
        RECT 121.150 122.845 122.500 123.015 ;
        RECT 121.150 122.685 121.400 122.845 ;
        RECT 121.910 122.415 122.160 122.675 ;
        RECT 120.790 122.165 122.160 122.415 ;
        RECT 118.720 121.875 118.960 122.165 ;
        RECT 119.760 122.085 119.930 122.165 ;
        RECT 119.160 121.615 119.580 121.995 ;
        RECT 119.760 121.835 120.390 122.085 ;
        RECT 120.860 121.615 121.190 121.995 ;
        RECT 121.360 121.875 121.530 122.165 ;
        RECT 122.330 122.000 122.500 122.845 ;
        RECT 122.950 122.675 123.170 123.545 ;
        RECT 123.395 123.425 124.090 123.615 ;
        RECT 122.670 122.295 123.170 122.675 ;
        RECT 123.340 122.625 123.750 123.245 ;
        RECT 123.920 122.455 124.090 123.425 ;
        RECT 123.395 122.285 124.090 122.455 ;
        RECT 121.710 121.615 122.090 121.995 ;
        RECT 122.330 121.830 123.160 122.000 ;
        RECT 123.395 121.785 123.565 122.285 ;
        RECT 123.735 121.615 124.065 122.115 ;
        RECT 124.280 121.785 124.505 123.905 ;
        RECT 124.675 123.785 125.005 124.165 ;
        RECT 125.175 123.615 125.345 123.905 ;
        RECT 124.680 123.445 125.345 123.615 ;
        RECT 124.680 122.455 124.910 123.445 ;
        RECT 126.525 123.415 127.735 124.165 ;
        RECT 125.080 122.625 125.430 123.275 ;
        RECT 126.525 122.705 127.045 123.245 ;
        RECT 127.215 122.875 127.735 123.415 ;
        RECT 124.680 122.285 125.345 122.455 ;
        RECT 124.675 121.615 125.005 122.115 ;
        RECT 125.175 121.785 125.345 122.285 ;
        RECT 126.525 121.615 127.735 122.705 ;
        RECT 14.660 121.445 127.820 121.615 ;
        RECT 14.745 120.355 15.955 121.445 ;
        RECT 14.745 119.645 15.265 120.185 ;
        RECT 15.435 119.815 15.955 120.355 ;
        RECT 16.185 120.305 16.395 121.445 ;
        RECT 16.565 120.295 16.895 121.275 ;
        RECT 17.065 120.305 17.295 121.445 ;
        RECT 17.545 120.305 17.775 121.445 ;
        RECT 17.945 120.295 18.275 121.275 ;
        RECT 18.445 120.305 18.655 121.445 ;
        RECT 18.925 120.305 19.155 121.445 ;
        RECT 19.325 120.295 19.655 121.275 ;
        RECT 19.825 120.305 20.035 121.445 ;
        RECT 20.265 120.685 20.780 121.095 ;
        RECT 21.015 120.685 21.185 121.445 ;
        RECT 21.355 121.105 23.385 121.275 ;
        RECT 14.745 118.895 15.955 119.645 ;
        RECT 16.185 118.895 16.395 119.715 ;
        RECT 16.565 119.695 16.815 120.295 ;
        RECT 16.985 119.885 17.315 120.135 ;
        RECT 17.525 119.885 17.855 120.135 ;
        RECT 16.565 119.065 16.895 119.695 ;
        RECT 17.065 118.895 17.295 119.715 ;
        RECT 17.545 118.895 17.775 119.715 ;
        RECT 18.025 119.695 18.275 120.295 ;
        RECT 18.905 119.885 19.235 120.135 ;
        RECT 17.945 119.065 18.275 119.695 ;
        RECT 18.445 118.895 18.655 119.715 ;
        RECT 18.925 118.895 19.155 119.715 ;
        RECT 19.405 119.695 19.655 120.295 ;
        RECT 20.265 119.875 20.605 120.685 ;
        RECT 21.355 120.440 21.525 121.105 ;
        RECT 21.920 120.765 23.045 120.935 ;
        RECT 20.775 120.250 21.525 120.440 ;
        RECT 21.695 120.425 22.705 120.595 ;
        RECT 19.325 119.065 19.655 119.695 ;
        RECT 19.825 118.895 20.035 119.715 ;
        RECT 20.265 119.705 21.495 119.875 ;
        RECT 20.540 119.100 20.785 119.705 ;
        RECT 21.005 118.895 21.515 119.430 ;
        RECT 21.695 119.065 21.885 120.425 ;
        RECT 22.055 119.405 22.330 120.225 ;
        RECT 22.535 119.625 22.705 120.425 ;
        RECT 22.875 119.635 23.045 120.765 ;
        RECT 23.215 120.135 23.385 121.105 ;
        RECT 23.555 120.305 23.725 121.445 ;
        RECT 23.895 120.305 24.230 121.275 ;
        RECT 23.215 119.805 23.410 120.135 ;
        RECT 23.635 119.805 23.890 120.135 ;
        RECT 23.635 119.635 23.805 119.805 ;
        RECT 24.060 119.635 24.230 120.305 ;
        RECT 24.405 120.280 24.695 121.445 ;
        RECT 24.870 120.305 25.205 121.275 ;
        RECT 25.375 120.305 25.545 121.445 ;
        RECT 25.715 121.105 27.745 121.275 ;
        RECT 22.875 119.465 23.805 119.635 ;
        RECT 22.875 119.430 23.050 119.465 ;
        RECT 22.055 119.235 22.335 119.405 ;
        RECT 22.055 119.065 22.330 119.235 ;
        RECT 22.520 119.065 23.050 119.430 ;
        RECT 23.475 118.895 23.805 119.295 ;
        RECT 23.975 119.065 24.230 119.635 ;
        RECT 24.870 119.635 25.040 120.305 ;
        RECT 25.715 120.135 25.885 121.105 ;
        RECT 25.210 119.805 25.465 120.135 ;
        RECT 25.690 119.805 25.885 120.135 ;
        RECT 26.055 120.765 27.180 120.935 ;
        RECT 25.295 119.635 25.465 119.805 ;
        RECT 26.055 119.635 26.225 120.765 ;
        RECT 24.405 118.895 24.695 119.620 ;
        RECT 24.870 119.065 25.125 119.635 ;
        RECT 25.295 119.465 26.225 119.635 ;
        RECT 26.395 120.425 27.405 120.595 ;
        RECT 26.395 119.625 26.565 120.425 ;
        RECT 26.770 120.085 27.045 120.225 ;
        RECT 26.765 119.915 27.045 120.085 ;
        RECT 26.050 119.430 26.225 119.465 ;
        RECT 25.295 118.895 25.625 119.295 ;
        RECT 26.050 119.065 26.580 119.430 ;
        RECT 26.770 119.065 27.045 119.915 ;
        RECT 27.215 119.065 27.405 120.425 ;
        RECT 27.575 120.440 27.745 121.105 ;
        RECT 27.915 120.685 28.085 121.445 ;
        RECT 28.320 120.685 28.835 121.095 ;
        RECT 27.575 120.250 28.325 120.440 ;
        RECT 28.495 119.875 28.835 120.685 ;
        RECT 27.605 119.705 28.835 119.875 ;
        RECT 29.380 120.465 29.635 121.135 ;
        RECT 29.815 120.645 30.100 121.445 ;
        RECT 30.280 120.725 30.610 121.235 ;
        RECT 27.585 118.895 28.095 119.430 ;
        RECT 28.315 119.100 28.560 119.705 ;
        RECT 29.380 119.605 29.560 120.465 ;
        RECT 30.280 120.135 30.530 120.725 ;
        RECT 30.880 120.575 31.050 121.185 ;
        RECT 31.220 120.755 31.550 121.445 ;
        RECT 31.780 120.895 32.020 121.185 ;
        RECT 32.220 121.065 32.640 121.445 ;
        RECT 32.820 120.975 33.450 121.225 ;
        RECT 33.920 121.065 34.250 121.445 ;
        RECT 32.820 120.895 32.990 120.975 ;
        RECT 34.420 120.895 34.590 121.185 ;
        RECT 34.770 121.065 35.150 121.445 ;
        RECT 35.390 121.060 36.220 121.230 ;
        RECT 31.780 120.725 32.990 120.895 ;
        RECT 29.730 119.805 30.530 120.135 ;
        RECT 29.380 119.405 29.635 119.605 ;
        RECT 29.295 119.235 29.635 119.405 ;
        RECT 29.380 119.075 29.635 119.235 ;
        RECT 29.815 118.895 30.100 119.355 ;
        RECT 30.280 119.155 30.530 119.805 ;
        RECT 30.730 120.555 31.050 120.575 ;
        RECT 30.730 120.385 32.650 120.555 ;
        RECT 30.730 119.490 30.920 120.385 ;
        RECT 32.820 120.215 32.990 120.725 ;
        RECT 33.160 120.465 33.680 120.775 ;
        RECT 31.090 120.045 32.990 120.215 ;
        RECT 31.090 119.985 31.420 120.045 ;
        RECT 31.570 119.815 31.900 119.875 ;
        RECT 31.240 119.545 31.900 119.815 ;
        RECT 30.730 119.160 31.050 119.490 ;
        RECT 31.230 118.895 31.890 119.375 ;
        RECT 32.090 119.285 32.260 120.045 ;
        RECT 33.160 119.875 33.340 120.285 ;
        RECT 32.430 119.705 32.760 119.825 ;
        RECT 33.510 119.705 33.680 120.465 ;
        RECT 32.430 119.535 33.680 119.705 ;
        RECT 33.850 120.645 35.220 120.895 ;
        RECT 33.850 119.875 34.040 120.645 ;
        RECT 34.970 120.385 35.220 120.645 ;
        RECT 34.210 120.215 34.460 120.375 ;
        RECT 35.390 120.215 35.560 121.060 ;
        RECT 36.455 120.775 36.625 121.275 ;
        RECT 36.795 120.945 37.125 121.445 ;
        RECT 35.730 120.385 36.230 120.765 ;
        RECT 36.455 120.605 37.150 120.775 ;
        RECT 34.210 120.045 35.560 120.215 ;
        RECT 35.140 120.005 35.560 120.045 ;
        RECT 33.850 119.535 34.270 119.875 ;
        RECT 34.560 119.545 34.970 119.875 ;
        RECT 32.090 119.115 32.940 119.285 ;
        RECT 33.500 118.895 33.820 119.355 ;
        RECT 34.020 119.105 34.270 119.535 ;
        RECT 34.560 118.895 34.970 119.335 ;
        RECT 35.140 119.275 35.310 120.005 ;
        RECT 35.480 119.455 35.830 119.825 ;
        RECT 36.010 119.515 36.230 120.385 ;
        RECT 36.400 119.815 36.810 120.435 ;
        RECT 36.980 119.635 37.150 120.605 ;
        RECT 36.455 119.445 37.150 119.635 ;
        RECT 35.140 119.075 36.155 119.275 ;
        RECT 36.455 119.115 36.625 119.445 ;
        RECT 36.795 118.895 37.125 119.275 ;
        RECT 37.340 119.155 37.565 121.275 ;
        RECT 37.735 120.945 38.065 121.445 ;
        RECT 38.235 120.775 38.405 121.275 ;
        RECT 37.740 120.605 38.405 120.775 ;
        RECT 37.740 119.615 37.970 120.605 ;
        RECT 38.140 119.785 38.490 120.435 ;
        RECT 38.665 120.355 41.255 121.445 ;
        RECT 41.425 120.685 41.940 121.095 ;
        RECT 42.175 120.685 42.345 121.445 ;
        RECT 42.515 121.105 44.545 121.275 ;
        RECT 38.665 119.835 39.875 120.355 ;
        RECT 40.045 119.665 41.255 120.185 ;
        RECT 41.425 119.875 41.765 120.685 ;
        RECT 42.515 120.440 42.685 121.105 ;
        RECT 43.080 120.765 44.205 120.935 ;
        RECT 41.935 120.250 42.685 120.440 ;
        RECT 42.855 120.425 43.865 120.595 ;
        RECT 41.425 119.705 42.655 119.875 ;
        RECT 37.740 119.445 38.405 119.615 ;
        RECT 37.735 118.895 38.065 119.275 ;
        RECT 38.235 119.155 38.405 119.445 ;
        RECT 38.665 118.895 41.255 119.665 ;
        RECT 41.700 119.100 41.945 119.705 ;
        RECT 42.165 118.895 42.675 119.430 ;
        RECT 42.855 119.065 43.045 120.425 ;
        RECT 43.215 119.745 43.490 120.225 ;
        RECT 43.215 119.575 43.495 119.745 ;
        RECT 43.695 119.625 43.865 120.425 ;
        RECT 44.035 119.635 44.205 120.765 ;
        RECT 44.375 120.135 44.545 121.105 ;
        RECT 44.715 120.305 44.885 121.445 ;
        RECT 45.055 120.305 45.390 121.275 ;
        RECT 44.375 119.805 44.570 120.135 ;
        RECT 44.795 119.805 45.050 120.135 ;
        RECT 44.795 119.635 44.965 119.805 ;
        RECT 45.220 119.635 45.390 120.305 ;
        RECT 45.565 120.355 48.155 121.445 ;
        RECT 48.385 120.610 48.640 121.445 ;
        RECT 48.810 120.440 49.070 121.245 ;
        RECT 49.240 120.610 49.500 121.445 ;
        RECT 49.670 120.440 49.925 121.245 ;
        RECT 45.565 119.835 46.775 120.355 ;
        RECT 48.325 120.270 49.925 120.440 ;
        RECT 50.165 120.280 50.455 121.445 ;
        RECT 50.625 120.305 50.965 121.275 ;
        RECT 51.135 120.305 51.305 121.445 ;
        RECT 51.575 120.645 51.825 121.445 ;
        RECT 52.470 120.475 52.800 121.275 ;
        RECT 53.100 120.645 53.430 121.445 ;
        RECT 53.600 120.475 53.930 121.275 ;
        RECT 51.495 120.305 53.930 120.475 ;
        RECT 54.345 120.305 54.575 121.445 ;
        RECT 46.945 119.665 48.155 120.185 ;
        RECT 43.215 119.065 43.490 119.575 ;
        RECT 44.035 119.465 44.965 119.635 ;
        RECT 44.035 119.430 44.210 119.465 ;
        RECT 43.680 119.065 44.210 119.430 ;
        RECT 44.635 118.895 44.965 119.295 ;
        RECT 45.135 119.065 45.390 119.635 ;
        RECT 45.565 118.895 48.155 119.665 ;
        RECT 48.325 119.705 48.605 120.270 ;
        RECT 48.775 119.875 49.995 120.100 ;
        RECT 48.325 119.535 49.055 119.705 ;
        RECT 50.625 119.695 50.800 120.305 ;
        RECT 51.495 120.055 51.665 120.305 ;
        RECT 50.970 119.885 51.665 120.055 ;
        RECT 51.840 119.885 52.260 120.085 ;
        RECT 52.430 119.885 52.760 120.085 ;
        RECT 52.930 119.885 53.260 120.085 ;
        RECT 48.330 118.895 48.660 119.365 ;
        RECT 48.830 119.090 49.055 119.535 ;
        RECT 49.225 118.895 49.520 119.420 ;
        RECT 50.165 118.895 50.455 119.620 ;
        RECT 50.625 119.065 50.965 119.695 ;
        RECT 51.135 118.895 51.385 119.695 ;
        RECT 51.575 119.545 52.800 119.715 ;
        RECT 51.575 119.065 51.905 119.545 ;
        RECT 52.075 118.895 52.300 119.355 ;
        RECT 52.470 119.065 52.800 119.545 ;
        RECT 53.430 119.675 53.600 120.305 ;
        RECT 54.745 120.295 55.075 121.275 ;
        RECT 55.245 120.305 55.455 121.445 ;
        RECT 55.685 120.685 56.200 121.095 ;
        RECT 56.435 120.685 56.605 121.445 ;
        RECT 56.775 121.105 58.805 121.275 ;
        RECT 53.785 119.885 54.135 120.135 ;
        RECT 54.325 119.885 54.655 120.135 ;
        RECT 53.430 119.065 53.930 119.675 ;
        RECT 54.345 118.895 54.575 119.715 ;
        RECT 54.825 119.695 55.075 120.295 ;
        RECT 55.685 119.875 56.025 120.685 ;
        RECT 56.775 120.440 56.945 121.105 ;
        RECT 57.340 120.765 58.465 120.935 ;
        RECT 56.195 120.250 56.945 120.440 ;
        RECT 57.115 120.425 58.125 120.595 ;
        RECT 54.745 119.065 55.075 119.695 ;
        RECT 55.245 118.895 55.455 119.715 ;
        RECT 55.685 119.705 56.915 119.875 ;
        RECT 55.960 119.100 56.205 119.705 ;
        RECT 56.425 118.895 56.935 119.430 ;
        RECT 57.115 119.065 57.305 120.425 ;
        RECT 57.475 120.085 57.750 120.225 ;
        RECT 57.475 119.915 57.755 120.085 ;
        RECT 57.475 119.065 57.750 119.915 ;
        RECT 57.955 119.625 58.125 120.425 ;
        RECT 58.295 119.635 58.465 120.765 ;
        RECT 58.635 120.135 58.805 121.105 ;
        RECT 58.975 120.305 59.145 121.445 ;
        RECT 59.315 120.305 59.650 121.275 ;
        RECT 60.750 121.010 66.095 121.445 ;
        RECT 58.635 119.805 58.830 120.135 ;
        RECT 59.055 119.805 59.310 120.135 ;
        RECT 59.055 119.635 59.225 119.805 ;
        RECT 59.480 119.635 59.650 120.305 ;
        RECT 62.340 119.760 62.690 121.010 ;
        RECT 66.355 120.775 66.525 121.275 ;
        RECT 66.695 120.945 67.025 121.445 ;
        RECT 66.355 120.605 67.020 120.775 ;
        RECT 58.295 119.465 59.225 119.635 ;
        RECT 58.295 119.430 58.470 119.465 ;
        RECT 57.940 119.065 58.470 119.430 ;
        RECT 58.895 118.895 59.225 119.295 ;
        RECT 59.395 119.065 59.650 119.635 ;
        RECT 64.170 119.440 64.510 120.270 ;
        RECT 66.270 119.785 66.620 120.435 ;
        RECT 66.790 119.615 67.020 120.605 ;
        RECT 66.355 119.445 67.020 119.615 ;
        RECT 60.750 118.895 66.095 119.440 ;
        RECT 66.355 119.155 66.525 119.445 ;
        RECT 66.695 118.895 67.025 119.275 ;
        RECT 67.195 119.155 67.420 121.275 ;
        RECT 67.635 120.945 67.965 121.445 ;
        RECT 68.135 120.775 68.305 121.275 ;
        RECT 68.540 121.060 69.370 121.230 ;
        RECT 69.610 121.065 69.990 121.445 ;
        RECT 67.610 120.605 68.305 120.775 ;
        RECT 67.610 119.635 67.780 120.605 ;
        RECT 67.950 119.815 68.360 120.435 ;
        RECT 68.530 120.385 69.030 120.765 ;
        RECT 67.610 119.445 68.305 119.635 ;
        RECT 68.530 119.515 68.750 120.385 ;
        RECT 69.200 120.215 69.370 121.060 ;
        RECT 70.170 120.895 70.340 121.185 ;
        RECT 70.510 121.065 70.840 121.445 ;
        RECT 71.310 120.975 71.940 121.225 ;
        RECT 72.120 121.065 72.540 121.445 ;
        RECT 71.770 120.895 71.940 120.975 ;
        RECT 72.740 120.895 72.980 121.185 ;
        RECT 69.540 120.645 70.910 120.895 ;
        RECT 69.540 120.385 69.790 120.645 ;
        RECT 70.300 120.215 70.550 120.375 ;
        RECT 69.200 120.045 70.550 120.215 ;
        RECT 69.200 120.005 69.620 120.045 ;
        RECT 68.930 119.455 69.280 119.825 ;
        RECT 67.635 118.895 67.965 119.275 ;
        RECT 68.135 119.115 68.305 119.445 ;
        RECT 69.450 119.275 69.620 120.005 ;
        RECT 70.720 119.875 70.910 120.645 ;
        RECT 69.790 119.545 70.200 119.875 ;
        RECT 70.490 119.535 70.910 119.875 ;
        RECT 71.080 120.465 71.600 120.775 ;
        RECT 71.770 120.725 72.980 120.895 ;
        RECT 73.210 120.755 73.540 121.445 ;
        RECT 71.080 119.705 71.250 120.465 ;
        RECT 71.420 119.875 71.600 120.285 ;
        RECT 71.770 120.215 71.940 120.725 ;
        RECT 73.710 120.575 73.880 121.185 ;
        RECT 74.150 120.725 74.480 121.235 ;
        RECT 73.710 120.555 74.030 120.575 ;
        RECT 72.110 120.385 74.030 120.555 ;
        RECT 71.770 120.045 73.670 120.215 ;
        RECT 72.000 119.705 72.330 119.825 ;
        RECT 71.080 119.535 72.330 119.705 ;
        RECT 68.605 119.075 69.620 119.275 ;
        RECT 69.790 118.895 70.200 119.335 ;
        RECT 70.490 119.105 70.740 119.535 ;
        RECT 70.940 118.895 71.260 119.355 ;
        RECT 72.500 119.285 72.670 120.045 ;
        RECT 73.340 119.985 73.670 120.045 ;
        RECT 72.860 119.815 73.190 119.875 ;
        RECT 72.860 119.545 73.520 119.815 ;
        RECT 73.840 119.490 74.030 120.385 ;
        RECT 71.820 119.115 72.670 119.285 ;
        RECT 72.870 118.895 73.530 119.375 ;
        RECT 73.710 119.160 74.030 119.490 ;
        RECT 74.230 120.135 74.480 120.725 ;
        RECT 74.660 120.645 74.945 121.445 ;
        RECT 75.125 121.105 75.380 121.135 ;
        RECT 75.125 120.935 75.465 121.105 ;
        RECT 75.125 120.465 75.380 120.935 ;
        RECT 74.230 119.805 75.030 120.135 ;
        RECT 74.230 119.155 74.480 119.805 ;
        RECT 75.200 119.605 75.380 120.465 ;
        RECT 75.925 120.280 76.215 121.445 ;
        RECT 76.760 121.105 77.015 121.135 ;
        RECT 76.675 120.935 77.015 121.105 ;
        RECT 76.760 120.465 77.015 120.935 ;
        RECT 77.195 120.645 77.480 121.445 ;
        RECT 77.660 120.725 77.990 121.235 ;
        RECT 74.660 118.895 74.945 119.355 ;
        RECT 75.125 119.075 75.380 119.605 ;
        RECT 75.925 118.895 76.215 119.620 ;
        RECT 76.760 119.605 76.940 120.465 ;
        RECT 77.660 120.135 77.910 120.725 ;
        RECT 78.260 120.575 78.430 121.185 ;
        RECT 78.600 120.755 78.930 121.445 ;
        RECT 79.160 120.895 79.400 121.185 ;
        RECT 79.600 121.065 80.020 121.445 ;
        RECT 80.200 120.975 80.830 121.225 ;
        RECT 81.300 121.065 81.630 121.445 ;
        RECT 80.200 120.895 80.370 120.975 ;
        RECT 81.800 120.895 81.970 121.185 ;
        RECT 82.150 121.065 82.530 121.445 ;
        RECT 82.770 121.060 83.600 121.230 ;
        RECT 79.160 120.725 80.370 120.895 ;
        RECT 77.110 119.805 77.910 120.135 ;
        RECT 76.760 119.075 77.015 119.605 ;
        RECT 77.195 118.895 77.480 119.355 ;
        RECT 77.660 119.155 77.910 119.805 ;
        RECT 78.110 120.555 78.430 120.575 ;
        RECT 78.110 120.385 80.030 120.555 ;
        RECT 78.110 119.490 78.300 120.385 ;
        RECT 80.200 120.215 80.370 120.725 ;
        RECT 80.540 120.465 81.060 120.775 ;
        RECT 78.470 120.045 80.370 120.215 ;
        RECT 78.470 119.985 78.800 120.045 ;
        RECT 78.950 119.815 79.280 119.875 ;
        RECT 78.620 119.545 79.280 119.815 ;
        RECT 78.110 119.160 78.430 119.490 ;
        RECT 78.610 118.895 79.270 119.375 ;
        RECT 79.470 119.285 79.640 120.045 ;
        RECT 80.540 119.875 80.720 120.285 ;
        RECT 79.810 119.705 80.140 119.825 ;
        RECT 80.890 119.705 81.060 120.465 ;
        RECT 79.810 119.535 81.060 119.705 ;
        RECT 81.230 120.645 82.600 120.895 ;
        RECT 81.230 119.875 81.420 120.645 ;
        RECT 82.350 120.385 82.600 120.645 ;
        RECT 81.590 120.215 81.840 120.375 ;
        RECT 82.770 120.215 82.940 121.060 ;
        RECT 83.835 120.775 84.005 121.275 ;
        RECT 84.175 120.945 84.505 121.445 ;
        RECT 83.110 120.385 83.610 120.765 ;
        RECT 83.835 120.605 84.530 120.775 ;
        RECT 81.590 120.045 82.940 120.215 ;
        RECT 82.520 120.005 82.940 120.045 ;
        RECT 81.230 119.535 81.650 119.875 ;
        RECT 81.940 119.545 82.350 119.875 ;
        RECT 79.470 119.115 80.320 119.285 ;
        RECT 80.880 118.895 81.200 119.355 ;
        RECT 81.400 119.105 81.650 119.535 ;
        RECT 81.940 118.895 82.350 119.335 ;
        RECT 82.520 119.275 82.690 120.005 ;
        RECT 82.860 119.455 83.210 119.825 ;
        RECT 83.390 119.515 83.610 120.385 ;
        RECT 83.780 119.815 84.190 120.435 ;
        RECT 84.360 119.635 84.530 120.605 ;
        RECT 83.835 119.445 84.530 119.635 ;
        RECT 82.520 119.075 83.535 119.275 ;
        RECT 83.835 119.115 84.005 119.445 ;
        RECT 84.175 118.895 84.505 119.275 ;
        RECT 84.720 119.155 84.945 121.275 ;
        RECT 85.115 120.945 85.445 121.445 ;
        RECT 85.615 120.775 85.785 121.275 ;
        RECT 85.120 120.605 85.785 120.775 ;
        RECT 85.120 119.615 85.350 120.605 ;
        RECT 85.520 119.785 85.870 120.435 ;
        RECT 86.045 120.370 86.315 121.275 ;
        RECT 86.485 120.685 86.815 121.445 ;
        RECT 86.995 120.515 87.165 121.275 ;
        RECT 85.120 119.445 85.785 119.615 ;
        RECT 85.115 118.895 85.445 119.275 ;
        RECT 85.615 119.155 85.785 119.445 ;
        RECT 86.045 119.570 86.215 120.370 ;
        RECT 86.500 120.345 87.165 120.515 ;
        RECT 88.260 120.465 88.515 121.135 ;
        RECT 88.695 120.645 88.980 121.445 ;
        RECT 89.160 120.725 89.490 121.235 ;
        RECT 86.500 120.200 86.670 120.345 ;
        RECT 86.385 119.870 86.670 120.200 ;
        RECT 86.500 119.615 86.670 119.870 ;
        RECT 86.905 119.795 87.235 120.165 ;
        RECT 86.045 119.065 86.305 119.570 ;
        RECT 86.500 119.445 87.165 119.615 ;
        RECT 86.485 118.895 86.815 119.275 ;
        RECT 86.995 119.065 87.165 119.445 ;
        RECT 88.260 119.605 88.440 120.465 ;
        RECT 89.160 120.135 89.410 120.725 ;
        RECT 89.760 120.575 89.930 121.185 ;
        RECT 90.100 120.755 90.430 121.445 ;
        RECT 90.660 120.895 90.900 121.185 ;
        RECT 91.100 121.065 91.520 121.445 ;
        RECT 91.700 120.975 92.330 121.225 ;
        RECT 92.800 121.065 93.130 121.445 ;
        RECT 91.700 120.895 91.870 120.975 ;
        RECT 93.300 120.895 93.470 121.185 ;
        RECT 93.650 121.065 94.030 121.445 ;
        RECT 94.270 121.060 95.100 121.230 ;
        RECT 90.660 120.725 91.870 120.895 ;
        RECT 88.610 119.805 89.410 120.135 ;
        RECT 88.260 119.405 88.515 119.605 ;
        RECT 88.175 119.235 88.515 119.405 ;
        RECT 88.260 119.075 88.515 119.235 ;
        RECT 88.695 118.895 88.980 119.355 ;
        RECT 89.160 119.155 89.410 119.805 ;
        RECT 89.610 120.555 89.930 120.575 ;
        RECT 89.610 120.385 91.530 120.555 ;
        RECT 89.610 119.490 89.800 120.385 ;
        RECT 91.700 120.215 91.870 120.725 ;
        RECT 92.040 120.465 92.560 120.775 ;
        RECT 89.970 120.045 91.870 120.215 ;
        RECT 89.970 119.985 90.300 120.045 ;
        RECT 90.450 119.815 90.780 119.875 ;
        RECT 90.120 119.545 90.780 119.815 ;
        RECT 89.610 119.160 89.930 119.490 ;
        RECT 90.110 118.895 90.770 119.375 ;
        RECT 90.970 119.285 91.140 120.045 ;
        RECT 92.040 119.875 92.220 120.285 ;
        RECT 91.310 119.705 91.640 119.825 ;
        RECT 92.390 119.705 92.560 120.465 ;
        RECT 91.310 119.535 92.560 119.705 ;
        RECT 92.730 120.645 94.100 120.895 ;
        RECT 92.730 119.875 92.920 120.645 ;
        RECT 93.850 120.385 94.100 120.645 ;
        RECT 93.090 120.215 93.340 120.375 ;
        RECT 94.270 120.215 94.440 121.060 ;
        RECT 95.335 120.775 95.505 121.275 ;
        RECT 95.675 120.945 96.005 121.445 ;
        RECT 94.610 120.385 95.110 120.765 ;
        RECT 95.335 120.605 96.030 120.775 ;
        RECT 93.090 120.045 94.440 120.215 ;
        RECT 94.020 120.005 94.440 120.045 ;
        RECT 92.730 119.535 93.150 119.875 ;
        RECT 93.440 119.545 93.850 119.875 ;
        RECT 90.970 119.115 91.820 119.285 ;
        RECT 92.380 118.895 92.700 119.355 ;
        RECT 92.900 119.105 93.150 119.535 ;
        RECT 93.440 118.895 93.850 119.335 ;
        RECT 94.020 119.275 94.190 120.005 ;
        RECT 94.360 119.455 94.710 119.825 ;
        RECT 94.890 119.515 95.110 120.385 ;
        RECT 95.280 119.815 95.690 120.435 ;
        RECT 95.860 119.635 96.030 120.605 ;
        RECT 95.335 119.445 96.030 119.635 ;
        RECT 94.020 119.075 95.035 119.275 ;
        RECT 95.335 119.115 95.505 119.445 ;
        RECT 95.675 118.895 96.005 119.275 ;
        RECT 96.220 119.155 96.445 121.275 ;
        RECT 96.615 120.945 96.945 121.445 ;
        RECT 97.115 120.775 97.285 121.275 ;
        RECT 96.620 120.605 97.285 120.775 ;
        RECT 96.620 119.615 96.850 120.605 ;
        RECT 97.020 119.785 97.370 120.435 ;
        RECT 97.585 120.305 97.815 121.445 ;
        RECT 97.985 120.295 98.315 121.275 ;
        RECT 98.485 120.305 98.695 121.445 ;
        RECT 98.925 120.370 99.195 121.275 ;
        RECT 99.365 120.685 99.695 121.445 ;
        RECT 99.875 120.515 100.045 121.275 ;
        RECT 97.565 119.885 97.895 120.135 ;
        RECT 96.620 119.445 97.285 119.615 ;
        RECT 96.615 118.895 96.945 119.275 ;
        RECT 97.115 119.155 97.285 119.445 ;
        RECT 97.585 118.895 97.815 119.715 ;
        RECT 98.065 119.695 98.315 120.295 ;
        RECT 97.985 119.065 98.315 119.695 ;
        RECT 98.485 118.895 98.695 119.715 ;
        RECT 98.925 119.570 99.095 120.370 ;
        RECT 99.380 120.345 100.045 120.515 ;
        RECT 100.305 120.370 100.575 121.275 ;
        RECT 100.745 120.685 101.075 121.445 ;
        RECT 101.255 120.515 101.425 121.275 ;
        RECT 99.380 120.200 99.550 120.345 ;
        RECT 99.265 119.870 99.550 120.200 ;
        RECT 99.380 119.615 99.550 119.870 ;
        RECT 99.785 119.795 100.115 120.165 ;
        RECT 98.925 119.065 99.185 119.570 ;
        RECT 99.380 119.445 100.045 119.615 ;
        RECT 99.365 118.895 99.695 119.275 ;
        RECT 99.875 119.065 100.045 119.445 ;
        RECT 100.305 119.570 100.475 120.370 ;
        RECT 100.760 120.345 101.425 120.515 ;
        RECT 100.760 120.200 100.930 120.345 ;
        RECT 101.685 120.280 101.975 121.445 ;
        RECT 102.155 120.635 102.450 121.445 ;
        RECT 100.645 119.870 100.930 120.200 ;
        RECT 100.760 119.615 100.930 119.870 ;
        RECT 101.165 119.795 101.495 120.165 ;
        RECT 102.630 120.135 102.875 121.275 ;
        RECT 103.050 120.635 103.310 121.445 ;
        RECT 103.910 121.440 110.185 121.445 ;
        RECT 103.490 120.135 103.740 121.270 ;
        RECT 103.910 120.645 104.170 121.440 ;
        RECT 104.340 120.545 104.600 121.270 ;
        RECT 104.770 120.715 105.030 121.440 ;
        RECT 105.200 120.545 105.460 121.270 ;
        RECT 105.630 120.715 105.890 121.440 ;
        RECT 106.060 120.545 106.320 121.270 ;
        RECT 106.490 120.715 106.750 121.440 ;
        RECT 106.920 120.545 107.180 121.270 ;
        RECT 107.350 120.715 107.595 121.440 ;
        RECT 107.765 120.545 108.025 121.270 ;
        RECT 108.210 120.715 108.455 121.440 ;
        RECT 108.625 120.545 108.885 121.270 ;
        RECT 109.070 120.715 109.315 121.440 ;
        RECT 109.485 120.545 109.745 121.270 ;
        RECT 109.930 120.715 110.185 121.440 ;
        RECT 104.340 120.530 109.745 120.545 ;
        RECT 110.355 120.530 110.645 121.270 ;
        RECT 110.815 120.700 111.085 121.445 ;
        RECT 111.400 120.575 111.685 121.445 ;
        RECT 111.855 120.815 112.115 121.275 ;
        RECT 112.290 120.985 112.545 121.445 ;
        RECT 112.715 120.815 112.975 121.275 ;
        RECT 111.855 120.645 112.975 120.815 ;
        RECT 113.145 120.645 113.455 121.445 ;
        RECT 104.340 120.305 111.085 120.530 ;
        RECT 111.855 120.395 112.115 120.645 ;
        RECT 113.625 120.475 113.935 121.275 ;
        RECT 100.305 119.065 100.565 119.570 ;
        RECT 100.760 119.445 101.425 119.615 ;
        RECT 100.745 118.895 101.075 119.275 ;
        RECT 101.255 119.065 101.425 119.445 ;
        RECT 101.685 118.895 101.975 119.620 ;
        RECT 102.145 119.575 102.460 120.135 ;
        RECT 102.630 119.885 109.750 120.135 ;
        RECT 102.145 118.895 102.450 119.405 ;
        RECT 102.630 119.075 102.880 119.885 ;
        RECT 103.050 118.895 103.310 119.420 ;
        RECT 103.490 119.075 103.740 119.885 ;
        RECT 109.920 119.745 111.085 120.305 ;
        RECT 111.360 120.225 112.115 120.395 ;
        RECT 112.905 120.305 113.935 120.475 ;
        RECT 109.920 119.715 111.115 119.745 ;
        RECT 104.340 119.575 111.115 119.715 ;
        RECT 111.360 119.715 111.765 120.225 ;
        RECT 112.905 120.055 113.075 120.305 ;
        RECT 111.935 119.885 113.075 120.055 ;
        RECT 104.340 119.545 111.085 119.575 ;
        RECT 111.360 119.545 113.010 119.715 ;
        RECT 113.245 119.565 113.595 120.135 ;
        RECT 103.910 118.895 104.170 119.455 ;
        RECT 104.340 119.090 104.600 119.545 ;
        RECT 104.770 118.895 105.030 119.375 ;
        RECT 105.200 119.090 105.460 119.545 ;
        RECT 105.630 118.895 105.890 119.375 ;
        RECT 106.060 119.090 106.320 119.545 ;
        RECT 106.490 118.895 106.735 119.375 ;
        RECT 106.905 119.090 107.180 119.545 ;
        RECT 107.350 118.895 107.595 119.375 ;
        RECT 107.765 119.090 108.025 119.545 ;
        RECT 108.205 118.895 108.455 119.375 ;
        RECT 108.625 119.090 108.885 119.545 ;
        RECT 109.065 118.895 109.315 119.375 ;
        RECT 109.485 119.090 109.745 119.545 ;
        RECT 109.925 118.895 110.185 119.375 ;
        RECT 110.355 119.090 110.615 119.545 ;
        RECT 110.785 118.895 111.085 119.375 ;
        RECT 111.405 118.895 111.685 119.375 ;
        RECT 111.855 119.155 112.115 119.545 ;
        RECT 112.290 118.895 112.545 119.375 ;
        RECT 112.715 119.155 113.010 119.545 ;
        RECT 113.765 119.395 113.935 120.305 ;
        RECT 114.105 120.355 115.315 121.445 ;
        RECT 115.485 120.685 116.000 121.095 ;
        RECT 116.235 120.685 116.405 121.445 ;
        RECT 116.575 121.105 118.605 121.275 ;
        RECT 114.105 119.815 114.625 120.355 ;
        RECT 114.795 119.645 115.315 120.185 ;
        RECT 115.485 119.875 115.825 120.685 ;
        RECT 116.575 120.440 116.745 121.105 ;
        RECT 117.140 120.765 118.265 120.935 ;
        RECT 115.995 120.250 116.745 120.440 ;
        RECT 116.915 120.425 117.925 120.595 ;
        RECT 115.485 119.705 116.715 119.875 ;
        RECT 113.190 118.895 113.465 119.375 ;
        RECT 113.635 119.065 113.935 119.395 ;
        RECT 114.105 118.895 115.315 119.645 ;
        RECT 115.760 119.100 116.005 119.705 ;
        RECT 116.225 118.895 116.735 119.430 ;
        RECT 116.915 119.065 117.105 120.425 ;
        RECT 117.275 120.085 117.550 120.225 ;
        RECT 117.275 119.915 117.555 120.085 ;
        RECT 117.275 119.065 117.550 119.915 ;
        RECT 117.755 119.625 117.925 120.425 ;
        RECT 118.095 119.635 118.265 120.765 ;
        RECT 118.435 120.135 118.605 121.105 ;
        RECT 118.775 120.305 118.945 121.445 ;
        RECT 119.115 120.305 119.450 121.275 ;
        RECT 119.715 120.515 119.885 121.275 ;
        RECT 120.065 120.685 120.395 121.445 ;
        RECT 119.715 120.345 120.380 120.515 ;
        RECT 120.565 120.370 120.835 121.275 ;
        RECT 118.435 119.805 118.630 120.135 ;
        RECT 118.855 119.805 119.110 120.135 ;
        RECT 118.855 119.635 119.025 119.805 ;
        RECT 119.280 119.635 119.450 120.305 ;
        RECT 120.210 120.200 120.380 120.345 ;
        RECT 119.645 119.795 119.975 120.165 ;
        RECT 120.210 119.870 120.495 120.200 ;
        RECT 118.095 119.465 119.025 119.635 ;
        RECT 118.095 119.430 118.270 119.465 ;
        RECT 117.740 119.065 118.270 119.430 ;
        RECT 118.695 118.895 119.025 119.295 ;
        RECT 119.195 119.065 119.450 119.635 ;
        RECT 120.210 119.615 120.380 119.870 ;
        RECT 119.715 119.445 120.380 119.615 ;
        RECT 120.665 119.570 120.835 120.370 ;
        RECT 121.095 120.515 121.265 121.275 ;
        RECT 121.445 120.685 121.775 121.445 ;
        RECT 121.095 120.345 121.760 120.515 ;
        RECT 121.945 120.370 122.215 121.275 ;
        RECT 121.590 120.200 121.760 120.345 ;
        RECT 121.025 119.795 121.355 120.165 ;
        RECT 121.590 119.870 121.875 120.200 ;
        RECT 121.590 119.615 121.760 119.870 ;
        RECT 119.715 119.065 119.885 119.445 ;
        RECT 120.065 118.895 120.395 119.275 ;
        RECT 120.575 119.065 120.835 119.570 ;
        RECT 121.095 119.445 121.760 119.615 ;
        RECT 122.045 119.570 122.215 120.370 ;
        RECT 122.845 120.355 126.355 121.445 ;
        RECT 126.525 120.355 127.735 121.445 ;
        RECT 122.845 119.835 124.535 120.355 ;
        RECT 124.705 119.665 126.355 120.185 ;
        RECT 126.525 119.815 127.045 120.355 ;
        RECT 121.095 119.065 121.265 119.445 ;
        RECT 121.445 118.895 121.775 119.275 ;
        RECT 121.955 119.065 122.215 119.570 ;
        RECT 122.845 118.895 126.355 119.665 ;
        RECT 127.215 119.645 127.735 120.185 ;
        RECT 126.525 118.895 127.735 119.645 ;
        RECT 14.660 118.725 127.820 118.895 ;
        RECT 14.745 117.975 15.955 118.725 ;
        RECT 14.745 117.435 15.265 117.975 ;
        RECT 16.125 117.955 17.795 118.725 ;
        RECT 18.340 118.385 18.595 118.545 ;
        RECT 18.255 118.215 18.595 118.385 ;
        RECT 18.775 118.265 19.060 118.725 ;
        RECT 15.435 117.265 15.955 117.805 ;
        RECT 14.745 116.175 15.955 117.265 ;
        RECT 16.125 117.265 16.875 117.785 ;
        RECT 17.045 117.435 17.795 117.955 ;
        RECT 18.340 118.015 18.595 118.215 ;
        RECT 16.125 116.175 17.795 117.265 ;
        RECT 18.340 117.155 18.520 118.015 ;
        RECT 19.240 117.815 19.490 118.465 ;
        RECT 18.690 117.485 19.490 117.815 ;
        RECT 18.340 116.485 18.595 117.155 ;
        RECT 18.775 116.175 19.060 116.975 ;
        RECT 19.240 116.895 19.490 117.485 ;
        RECT 19.690 118.130 20.010 118.460 ;
        RECT 20.190 118.245 20.850 118.725 ;
        RECT 21.050 118.335 21.900 118.505 ;
        RECT 19.690 117.235 19.880 118.130 ;
        RECT 20.200 117.805 20.860 118.075 ;
        RECT 20.530 117.745 20.860 117.805 ;
        RECT 20.050 117.575 20.380 117.635 ;
        RECT 21.050 117.575 21.220 118.335 ;
        RECT 22.460 118.265 22.780 118.725 ;
        RECT 22.980 118.085 23.230 118.515 ;
        RECT 23.520 118.285 23.930 118.725 ;
        RECT 24.100 118.345 25.115 118.545 ;
        RECT 21.390 117.915 22.640 118.085 ;
        RECT 21.390 117.795 21.720 117.915 ;
        RECT 20.050 117.405 21.950 117.575 ;
        RECT 19.690 117.065 21.610 117.235 ;
        RECT 19.690 117.045 20.010 117.065 ;
        RECT 19.240 116.385 19.570 116.895 ;
        RECT 19.840 116.435 20.010 117.045 ;
        RECT 21.780 116.895 21.950 117.405 ;
        RECT 22.120 117.335 22.300 117.745 ;
        RECT 22.470 117.155 22.640 117.915 ;
        RECT 20.180 116.175 20.510 116.865 ;
        RECT 20.740 116.725 21.950 116.895 ;
        RECT 22.120 116.845 22.640 117.155 ;
        RECT 22.810 117.745 23.230 118.085 ;
        RECT 23.520 117.745 23.930 118.075 ;
        RECT 22.810 116.975 23.000 117.745 ;
        RECT 24.100 117.615 24.270 118.345 ;
        RECT 25.415 118.175 25.585 118.505 ;
        RECT 25.755 118.345 26.085 118.725 ;
        RECT 24.440 117.795 24.790 118.165 ;
        RECT 24.100 117.575 24.520 117.615 ;
        RECT 23.170 117.405 24.520 117.575 ;
        RECT 23.170 117.245 23.420 117.405 ;
        RECT 23.930 116.975 24.180 117.235 ;
        RECT 22.810 116.725 24.180 116.975 ;
        RECT 20.740 116.435 20.980 116.725 ;
        RECT 21.780 116.645 21.950 116.725 ;
        RECT 21.180 116.175 21.600 116.555 ;
        RECT 21.780 116.395 22.410 116.645 ;
        RECT 22.880 116.175 23.210 116.555 ;
        RECT 23.380 116.435 23.550 116.725 ;
        RECT 24.350 116.560 24.520 117.405 ;
        RECT 24.970 117.235 25.190 118.105 ;
        RECT 25.415 117.985 26.110 118.175 ;
        RECT 24.690 116.855 25.190 117.235 ;
        RECT 25.360 117.185 25.770 117.805 ;
        RECT 25.940 117.015 26.110 117.985 ;
        RECT 25.415 116.845 26.110 117.015 ;
        RECT 23.730 116.175 24.110 116.555 ;
        RECT 24.350 116.390 25.180 116.560 ;
        RECT 25.415 116.345 25.585 116.845 ;
        RECT 25.755 116.175 26.085 116.675 ;
        RECT 26.300 116.345 26.525 118.465 ;
        RECT 26.695 118.345 27.025 118.725 ;
        RECT 27.195 118.175 27.365 118.465 ;
        RECT 27.715 118.245 28.015 118.725 ;
        RECT 26.700 118.005 27.365 118.175 ;
        RECT 28.185 118.075 28.445 118.530 ;
        RECT 28.615 118.245 28.875 118.725 ;
        RECT 29.055 118.075 29.315 118.530 ;
        RECT 29.485 118.245 29.735 118.725 ;
        RECT 29.915 118.075 30.175 118.530 ;
        RECT 30.345 118.245 30.595 118.725 ;
        RECT 30.775 118.075 31.035 118.530 ;
        RECT 31.205 118.245 31.450 118.725 ;
        RECT 31.620 118.075 31.895 118.530 ;
        RECT 32.065 118.245 32.310 118.725 ;
        RECT 32.480 118.075 32.740 118.530 ;
        RECT 32.910 118.245 33.170 118.725 ;
        RECT 33.340 118.075 33.600 118.530 ;
        RECT 33.770 118.245 34.030 118.725 ;
        RECT 34.200 118.075 34.460 118.530 ;
        RECT 34.630 118.165 34.890 118.725 ;
        RECT 26.700 117.015 26.930 118.005 ;
        RECT 27.715 117.905 34.460 118.075 ;
        RECT 27.100 117.185 27.450 117.835 ;
        RECT 27.715 117.315 28.880 117.905 ;
        RECT 35.060 117.735 35.310 118.545 ;
        RECT 35.490 118.200 35.750 118.725 ;
        RECT 35.920 117.735 36.170 118.545 ;
        RECT 36.350 118.215 36.655 118.725 ;
        RECT 29.050 117.485 36.170 117.735 ;
        RECT 36.340 117.485 36.655 118.045 ;
        RECT 37.285 118.000 37.575 118.725 ;
        RECT 38.120 118.385 38.375 118.545 ;
        RECT 38.035 118.215 38.375 118.385 ;
        RECT 38.555 118.265 38.840 118.725 ;
        RECT 38.120 118.015 38.375 118.215 ;
        RECT 27.715 117.090 34.460 117.315 ;
        RECT 26.700 116.845 27.365 117.015 ;
        RECT 26.695 116.175 27.025 116.675 ;
        RECT 27.195 116.345 27.365 116.845 ;
        RECT 27.715 116.175 27.985 116.920 ;
        RECT 28.155 116.350 28.445 117.090 ;
        RECT 29.055 117.075 34.460 117.090 ;
        RECT 28.615 116.180 28.870 116.905 ;
        RECT 29.055 116.350 29.315 117.075 ;
        RECT 29.485 116.180 29.730 116.905 ;
        RECT 29.915 116.350 30.175 117.075 ;
        RECT 30.345 116.180 30.590 116.905 ;
        RECT 30.775 116.350 31.035 117.075 ;
        RECT 31.205 116.180 31.450 116.905 ;
        RECT 31.620 116.350 31.880 117.075 ;
        RECT 32.050 116.180 32.310 116.905 ;
        RECT 32.480 116.350 32.740 117.075 ;
        RECT 32.910 116.180 33.170 116.905 ;
        RECT 33.340 116.350 33.600 117.075 ;
        RECT 33.770 116.180 34.030 116.905 ;
        RECT 34.200 116.350 34.460 117.075 ;
        RECT 34.630 116.180 34.890 116.975 ;
        RECT 35.060 116.350 35.310 117.485 ;
        RECT 28.615 116.175 34.890 116.180 ;
        RECT 35.490 116.175 35.750 116.985 ;
        RECT 35.925 116.345 36.170 117.485 ;
        RECT 36.350 116.175 36.645 116.985 ;
        RECT 37.285 116.175 37.575 117.340 ;
        RECT 38.120 117.155 38.300 118.015 ;
        RECT 39.020 117.815 39.270 118.465 ;
        RECT 38.470 117.485 39.270 117.815 ;
        RECT 38.120 116.485 38.375 117.155 ;
        RECT 38.555 116.175 38.840 116.975 ;
        RECT 39.020 116.895 39.270 117.485 ;
        RECT 39.470 118.130 39.790 118.460 ;
        RECT 39.970 118.245 40.630 118.725 ;
        RECT 40.830 118.335 41.680 118.505 ;
        RECT 39.470 117.235 39.660 118.130 ;
        RECT 39.980 117.805 40.640 118.075 ;
        RECT 40.310 117.745 40.640 117.805 ;
        RECT 39.830 117.575 40.160 117.635 ;
        RECT 40.830 117.575 41.000 118.335 ;
        RECT 42.240 118.265 42.560 118.725 ;
        RECT 42.760 118.085 43.010 118.515 ;
        RECT 43.300 118.285 43.710 118.725 ;
        RECT 43.880 118.345 44.895 118.545 ;
        RECT 41.170 117.915 42.420 118.085 ;
        RECT 41.170 117.795 41.500 117.915 ;
        RECT 39.830 117.405 41.730 117.575 ;
        RECT 39.470 117.065 41.390 117.235 ;
        RECT 39.470 117.045 39.790 117.065 ;
        RECT 39.020 116.385 39.350 116.895 ;
        RECT 39.620 116.435 39.790 117.045 ;
        RECT 41.560 116.895 41.730 117.405 ;
        RECT 41.900 117.335 42.080 117.745 ;
        RECT 42.250 117.155 42.420 117.915 ;
        RECT 39.960 116.175 40.290 116.865 ;
        RECT 40.520 116.725 41.730 116.895 ;
        RECT 41.900 116.845 42.420 117.155 ;
        RECT 42.590 117.745 43.010 118.085 ;
        RECT 43.300 117.745 43.710 118.075 ;
        RECT 42.590 116.975 42.780 117.745 ;
        RECT 43.880 117.615 44.050 118.345 ;
        RECT 45.195 118.175 45.365 118.505 ;
        RECT 45.535 118.345 45.865 118.725 ;
        RECT 44.220 117.795 44.570 118.165 ;
        RECT 43.880 117.575 44.300 117.615 ;
        RECT 42.950 117.405 44.300 117.575 ;
        RECT 42.950 117.245 43.200 117.405 ;
        RECT 43.710 116.975 43.960 117.235 ;
        RECT 42.590 116.725 43.960 116.975 ;
        RECT 40.520 116.435 40.760 116.725 ;
        RECT 41.560 116.645 41.730 116.725 ;
        RECT 40.960 116.175 41.380 116.555 ;
        RECT 41.560 116.395 42.190 116.645 ;
        RECT 42.660 116.175 42.990 116.555 ;
        RECT 43.160 116.435 43.330 116.725 ;
        RECT 44.130 116.560 44.300 117.405 ;
        RECT 44.750 117.235 44.970 118.105 ;
        RECT 45.195 117.985 45.890 118.175 ;
        RECT 44.470 116.855 44.970 117.235 ;
        RECT 45.140 117.185 45.550 117.805 ;
        RECT 45.720 117.015 45.890 117.985 ;
        RECT 45.195 116.845 45.890 117.015 ;
        RECT 43.510 116.175 43.890 116.555 ;
        RECT 44.130 116.390 44.960 116.560 ;
        RECT 45.195 116.345 45.365 116.845 ;
        RECT 45.535 116.175 45.865 116.675 ;
        RECT 46.080 116.345 46.305 118.465 ;
        RECT 46.475 118.345 46.805 118.725 ;
        RECT 46.975 118.175 47.145 118.465 ;
        RECT 46.480 118.005 47.145 118.175 ;
        RECT 46.480 117.015 46.710 118.005 ;
        RECT 47.555 117.925 47.885 118.725 ;
        RECT 48.055 118.075 48.225 118.555 ;
        RECT 48.395 118.245 48.725 118.725 ;
        RECT 48.895 118.075 49.065 118.555 ;
        RECT 49.315 118.245 49.555 118.725 ;
        RECT 49.735 118.075 49.905 118.555 ;
        RECT 48.055 117.905 49.065 118.075 ;
        RECT 49.270 117.905 49.905 118.075 ;
        RECT 50.165 117.975 51.375 118.725 ;
        RECT 51.920 118.385 52.175 118.545 ;
        RECT 51.835 118.215 52.175 118.385 ;
        RECT 52.355 118.265 52.640 118.725 ;
        RECT 46.880 117.185 47.230 117.835 ;
        RECT 48.055 117.365 48.550 117.905 ;
        RECT 49.270 117.735 49.440 117.905 ;
        RECT 48.940 117.565 49.440 117.735 ;
        RECT 46.480 116.845 47.145 117.015 ;
        RECT 46.475 116.175 46.805 116.675 ;
        RECT 46.975 116.345 47.145 116.845 ;
        RECT 47.555 116.175 47.885 117.325 ;
        RECT 48.055 117.195 49.065 117.365 ;
        RECT 48.055 116.345 48.225 117.195 ;
        RECT 48.395 116.175 48.725 116.975 ;
        RECT 48.895 116.345 49.065 117.195 ;
        RECT 49.270 117.325 49.440 117.565 ;
        RECT 49.610 117.495 49.990 117.735 ;
        RECT 49.270 117.155 49.985 117.325 ;
        RECT 49.245 116.175 49.485 116.975 ;
        RECT 49.655 116.345 49.985 117.155 ;
        RECT 50.165 117.265 50.685 117.805 ;
        RECT 50.855 117.435 51.375 117.975 ;
        RECT 51.920 118.015 52.175 118.215 ;
        RECT 50.165 116.175 51.375 117.265 ;
        RECT 51.920 117.155 52.100 118.015 ;
        RECT 52.820 117.815 53.070 118.465 ;
        RECT 52.270 117.485 53.070 117.815 ;
        RECT 51.920 116.485 52.175 117.155 ;
        RECT 52.355 116.175 52.640 116.975 ;
        RECT 52.820 116.895 53.070 117.485 ;
        RECT 53.270 118.130 53.590 118.460 ;
        RECT 53.770 118.245 54.430 118.725 ;
        RECT 54.630 118.335 55.480 118.505 ;
        RECT 53.270 117.235 53.460 118.130 ;
        RECT 53.780 117.805 54.440 118.075 ;
        RECT 54.110 117.745 54.440 117.805 ;
        RECT 53.630 117.575 53.960 117.635 ;
        RECT 54.630 117.575 54.800 118.335 ;
        RECT 56.040 118.265 56.360 118.725 ;
        RECT 56.560 118.085 56.810 118.515 ;
        RECT 57.100 118.285 57.510 118.725 ;
        RECT 57.680 118.345 58.695 118.545 ;
        RECT 54.970 117.915 56.220 118.085 ;
        RECT 54.970 117.795 55.300 117.915 ;
        RECT 53.630 117.405 55.530 117.575 ;
        RECT 53.270 117.065 55.190 117.235 ;
        RECT 53.270 117.045 53.590 117.065 ;
        RECT 52.820 116.385 53.150 116.895 ;
        RECT 53.420 116.435 53.590 117.045 ;
        RECT 55.360 116.895 55.530 117.405 ;
        RECT 55.700 117.335 55.880 117.745 ;
        RECT 56.050 117.155 56.220 117.915 ;
        RECT 53.760 116.175 54.090 116.865 ;
        RECT 54.320 116.725 55.530 116.895 ;
        RECT 55.700 116.845 56.220 117.155 ;
        RECT 56.390 117.745 56.810 118.085 ;
        RECT 57.100 117.745 57.510 118.075 ;
        RECT 56.390 116.975 56.580 117.745 ;
        RECT 57.680 117.615 57.850 118.345 ;
        RECT 58.995 118.175 59.165 118.505 ;
        RECT 59.335 118.345 59.665 118.725 ;
        RECT 58.020 117.795 58.370 118.165 ;
        RECT 57.680 117.575 58.100 117.615 ;
        RECT 56.750 117.405 58.100 117.575 ;
        RECT 56.750 117.245 57.000 117.405 ;
        RECT 57.510 116.975 57.760 117.235 ;
        RECT 56.390 116.725 57.760 116.975 ;
        RECT 54.320 116.435 54.560 116.725 ;
        RECT 55.360 116.645 55.530 116.725 ;
        RECT 54.760 116.175 55.180 116.555 ;
        RECT 55.360 116.395 55.990 116.645 ;
        RECT 56.460 116.175 56.790 116.555 ;
        RECT 56.960 116.435 57.130 116.725 ;
        RECT 57.930 116.560 58.100 117.405 ;
        RECT 58.550 117.235 58.770 118.105 ;
        RECT 58.995 117.985 59.690 118.175 ;
        RECT 58.270 116.855 58.770 117.235 ;
        RECT 58.940 117.185 59.350 117.805 ;
        RECT 59.520 117.015 59.690 117.985 ;
        RECT 58.995 116.845 59.690 117.015 ;
        RECT 57.310 116.175 57.690 116.555 ;
        RECT 57.930 116.390 58.760 116.560 ;
        RECT 58.995 116.345 59.165 116.845 ;
        RECT 59.335 116.175 59.665 116.675 ;
        RECT 59.880 116.345 60.105 118.465 ;
        RECT 60.275 118.345 60.605 118.725 ;
        RECT 60.775 118.175 60.945 118.465 ;
        RECT 60.280 118.005 60.945 118.175 ;
        RECT 61.205 118.050 61.465 118.555 ;
        RECT 61.645 118.345 61.975 118.725 ;
        RECT 62.155 118.175 62.325 118.555 ;
        RECT 60.280 117.015 60.510 118.005 ;
        RECT 60.680 117.185 61.030 117.835 ;
        RECT 61.205 117.250 61.375 118.050 ;
        RECT 61.660 118.005 62.325 118.175 ;
        RECT 61.660 117.750 61.830 118.005 ;
        RECT 63.045 118.000 63.335 118.725 ;
        RECT 63.965 117.955 65.635 118.725 ;
        RECT 61.545 117.420 61.830 117.750 ;
        RECT 62.065 117.455 62.395 117.825 ;
        RECT 61.660 117.275 61.830 117.420 ;
        RECT 60.280 116.845 60.945 117.015 ;
        RECT 60.275 116.175 60.605 116.675 ;
        RECT 60.775 116.345 60.945 116.845 ;
        RECT 61.205 116.345 61.475 117.250 ;
        RECT 61.660 117.105 62.325 117.275 ;
        RECT 61.645 116.175 61.975 116.935 ;
        RECT 62.155 116.345 62.325 117.105 ;
        RECT 63.045 116.175 63.335 117.340 ;
        RECT 63.965 117.265 64.715 117.785 ;
        RECT 64.885 117.435 65.635 117.955 ;
        RECT 66.080 117.915 66.325 118.520 ;
        RECT 66.545 118.190 67.055 118.725 ;
        RECT 65.805 117.745 67.035 117.915 ;
        RECT 63.965 116.175 65.635 117.265 ;
        RECT 65.805 116.935 66.145 117.745 ;
        RECT 66.315 117.180 67.065 117.370 ;
        RECT 65.805 116.525 66.320 116.935 ;
        RECT 66.555 116.175 66.725 116.935 ;
        RECT 66.895 116.515 67.065 117.180 ;
        RECT 67.235 117.195 67.425 118.555 ;
        RECT 67.595 117.705 67.870 118.555 ;
        RECT 68.060 118.190 68.590 118.555 ;
        RECT 69.015 118.325 69.345 118.725 ;
        RECT 68.415 118.155 68.590 118.190 ;
        RECT 67.595 117.535 67.875 117.705 ;
        RECT 67.595 117.395 67.870 117.535 ;
        RECT 68.075 117.195 68.245 117.995 ;
        RECT 67.235 117.025 68.245 117.195 ;
        RECT 68.415 117.985 69.345 118.155 ;
        RECT 69.515 117.985 69.770 118.555 ;
        RECT 70.495 118.175 70.665 118.555 ;
        RECT 70.845 118.345 71.175 118.725 ;
        RECT 70.495 118.005 71.160 118.175 ;
        RECT 71.355 118.050 71.615 118.555 ;
        RECT 68.415 116.855 68.585 117.985 ;
        RECT 69.175 117.815 69.345 117.985 ;
        RECT 67.460 116.685 68.585 116.855 ;
        RECT 68.755 117.485 68.950 117.815 ;
        RECT 69.175 117.485 69.430 117.815 ;
        RECT 68.755 116.515 68.925 117.485 ;
        RECT 69.600 117.315 69.770 117.985 ;
        RECT 70.425 117.455 70.755 117.825 ;
        RECT 70.990 117.750 71.160 118.005 ;
        RECT 66.895 116.345 68.925 116.515 ;
        RECT 69.095 116.175 69.265 117.315 ;
        RECT 69.435 116.345 69.770 117.315 ;
        RECT 70.990 117.420 71.275 117.750 ;
        RECT 70.990 117.275 71.160 117.420 ;
        RECT 70.495 117.105 71.160 117.275 ;
        RECT 71.445 117.250 71.615 118.050 ;
        RECT 72.705 117.955 76.215 118.725 ;
        RECT 70.495 116.345 70.665 117.105 ;
        RECT 70.845 116.175 71.175 116.935 ;
        RECT 71.345 116.345 71.615 117.250 ;
        RECT 72.705 117.265 74.395 117.785 ;
        RECT 74.565 117.435 76.215 117.955 ;
        RECT 76.425 117.905 76.655 118.725 ;
        RECT 76.825 117.925 77.155 118.555 ;
        RECT 76.405 117.485 76.735 117.735 ;
        RECT 76.905 117.325 77.155 117.925 ;
        RECT 77.325 117.905 77.535 118.725 ;
        RECT 77.765 118.050 78.025 118.555 ;
        RECT 78.205 118.345 78.535 118.725 ;
        RECT 78.715 118.175 78.885 118.555 ;
        RECT 72.705 116.175 76.215 117.265 ;
        RECT 76.425 116.175 76.655 117.315 ;
        RECT 76.825 116.345 77.155 117.325 ;
        RECT 77.325 116.175 77.535 117.315 ;
        RECT 77.765 117.250 77.935 118.050 ;
        RECT 78.220 118.005 78.885 118.175 ;
        RECT 79.235 118.175 79.405 118.465 ;
        RECT 79.575 118.345 79.905 118.725 ;
        RECT 79.235 118.005 79.900 118.175 ;
        RECT 78.220 117.750 78.390 118.005 ;
        RECT 78.105 117.420 78.390 117.750 ;
        RECT 78.625 117.455 78.955 117.825 ;
        RECT 78.220 117.275 78.390 117.420 ;
        RECT 77.765 116.345 78.035 117.250 ;
        RECT 78.220 117.105 78.885 117.275 ;
        RECT 79.150 117.185 79.500 117.835 ;
        RECT 78.205 116.175 78.535 116.935 ;
        RECT 78.715 116.345 78.885 117.105 ;
        RECT 79.670 117.015 79.900 118.005 ;
        RECT 79.235 116.845 79.900 117.015 ;
        RECT 79.235 116.345 79.405 116.845 ;
        RECT 79.575 116.175 79.905 116.675 ;
        RECT 80.075 116.345 80.300 118.465 ;
        RECT 80.515 118.345 80.845 118.725 ;
        RECT 81.015 118.175 81.185 118.505 ;
        RECT 81.485 118.345 82.500 118.545 ;
        RECT 80.490 117.985 81.185 118.175 ;
        RECT 80.490 117.015 80.660 117.985 ;
        RECT 80.830 117.185 81.240 117.805 ;
        RECT 81.410 117.235 81.630 118.105 ;
        RECT 81.810 117.795 82.160 118.165 ;
        RECT 82.330 117.615 82.500 118.345 ;
        RECT 82.670 118.285 83.080 118.725 ;
        RECT 83.370 118.085 83.620 118.515 ;
        RECT 83.820 118.265 84.140 118.725 ;
        RECT 84.700 118.335 85.550 118.505 ;
        RECT 82.670 117.745 83.080 118.075 ;
        RECT 83.370 117.745 83.790 118.085 ;
        RECT 82.080 117.575 82.500 117.615 ;
        RECT 82.080 117.405 83.430 117.575 ;
        RECT 80.490 116.845 81.185 117.015 ;
        RECT 81.410 116.855 81.910 117.235 ;
        RECT 80.515 116.175 80.845 116.675 ;
        RECT 81.015 116.345 81.185 116.845 ;
        RECT 82.080 116.560 82.250 117.405 ;
        RECT 83.180 117.245 83.430 117.405 ;
        RECT 82.420 116.975 82.670 117.235 ;
        RECT 83.600 116.975 83.790 117.745 ;
        RECT 82.420 116.725 83.790 116.975 ;
        RECT 83.960 117.915 85.210 118.085 ;
        RECT 83.960 117.155 84.130 117.915 ;
        RECT 84.880 117.795 85.210 117.915 ;
        RECT 84.300 117.335 84.480 117.745 ;
        RECT 85.380 117.575 85.550 118.335 ;
        RECT 85.750 118.245 86.410 118.725 ;
        RECT 86.590 118.130 86.910 118.460 ;
        RECT 85.740 117.805 86.400 118.075 ;
        RECT 85.740 117.745 86.070 117.805 ;
        RECT 86.220 117.575 86.550 117.635 ;
        RECT 84.650 117.405 86.550 117.575 ;
        RECT 83.960 116.845 84.480 117.155 ;
        RECT 84.650 116.895 84.820 117.405 ;
        RECT 86.720 117.235 86.910 118.130 ;
        RECT 84.990 117.065 86.910 117.235 ;
        RECT 86.590 117.045 86.910 117.065 ;
        RECT 87.110 117.815 87.360 118.465 ;
        RECT 87.540 118.265 87.825 118.725 ;
        RECT 88.005 118.015 88.260 118.545 ;
        RECT 87.110 117.485 87.910 117.815 ;
        RECT 84.650 116.725 85.860 116.895 ;
        RECT 81.420 116.390 82.250 116.560 ;
        RECT 82.490 116.175 82.870 116.555 ;
        RECT 83.050 116.435 83.220 116.725 ;
        RECT 84.650 116.645 84.820 116.725 ;
        RECT 83.390 116.175 83.720 116.555 ;
        RECT 84.190 116.395 84.820 116.645 ;
        RECT 85.000 116.175 85.420 116.555 ;
        RECT 85.620 116.435 85.860 116.725 ;
        RECT 86.090 116.175 86.420 116.865 ;
        RECT 86.590 116.435 86.760 117.045 ;
        RECT 87.110 116.895 87.360 117.485 ;
        RECT 88.080 117.365 88.260 118.015 ;
        RECT 88.805 118.000 89.095 118.725 ;
        RECT 89.325 117.905 89.535 118.725 ;
        RECT 89.705 117.925 90.035 118.555 ;
        RECT 88.080 117.195 88.345 117.365 ;
        RECT 88.080 117.155 88.260 117.195 ;
        RECT 87.030 116.385 87.360 116.895 ;
        RECT 87.540 116.175 87.825 116.975 ;
        RECT 88.005 116.485 88.260 117.155 ;
        RECT 88.805 116.175 89.095 117.340 ;
        RECT 89.705 117.325 89.955 117.925 ;
        RECT 90.205 117.905 90.435 118.725 ;
        RECT 91.840 117.915 92.085 118.520 ;
        RECT 92.305 118.190 92.815 118.725 ;
        RECT 91.565 117.745 92.795 117.915 ;
        RECT 90.125 117.485 90.455 117.735 ;
        RECT 89.325 116.175 89.535 117.315 ;
        RECT 89.705 116.345 90.035 117.325 ;
        RECT 90.205 116.175 90.435 117.315 ;
        RECT 91.565 116.935 91.905 117.745 ;
        RECT 92.075 117.180 92.825 117.370 ;
        RECT 91.565 116.525 92.080 116.935 ;
        RECT 92.315 116.175 92.485 116.935 ;
        RECT 92.655 116.515 92.825 117.180 ;
        RECT 92.995 117.195 93.185 118.555 ;
        RECT 93.355 118.385 93.630 118.555 ;
        RECT 93.355 118.215 93.635 118.385 ;
        RECT 93.355 117.395 93.630 118.215 ;
        RECT 93.820 118.190 94.350 118.555 ;
        RECT 94.775 118.325 95.105 118.725 ;
        RECT 94.175 118.155 94.350 118.190 ;
        RECT 93.835 117.195 94.005 117.995 ;
        RECT 92.995 117.025 94.005 117.195 ;
        RECT 94.175 117.985 95.105 118.155 ;
        RECT 95.275 117.985 95.530 118.555 ;
        RECT 94.175 116.855 94.345 117.985 ;
        RECT 94.935 117.815 95.105 117.985 ;
        RECT 93.220 116.685 94.345 116.855 ;
        RECT 94.515 117.485 94.710 117.815 ;
        RECT 94.935 117.485 95.190 117.815 ;
        RECT 94.515 116.515 94.685 117.485 ;
        RECT 95.360 117.315 95.530 117.985 ;
        RECT 96.165 117.955 97.835 118.725 ;
        RECT 98.010 118.180 103.355 118.725 ;
        RECT 92.655 116.345 94.685 116.515 ;
        RECT 94.855 116.175 95.025 117.315 ;
        RECT 95.195 116.345 95.530 117.315 ;
        RECT 96.165 117.265 96.915 117.785 ;
        RECT 97.085 117.435 97.835 117.955 ;
        RECT 96.165 116.175 97.835 117.265 ;
        RECT 99.600 116.610 99.950 117.860 ;
        RECT 101.430 117.350 101.770 118.180 ;
        RECT 103.565 117.905 103.795 118.725 ;
        RECT 103.965 117.925 104.295 118.555 ;
        RECT 103.545 117.485 103.875 117.735 ;
        RECT 104.045 117.325 104.295 117.925 ;
        RECT 104.465 117.905 104.675 118.725 ;
        RECT 105.180 117.915 105.425 118.520 ;
        RECT 105.645 118.190 106.155 118.725 ;
        RECT 98.010 116.175 103.355 116.610 ;
        RECT 103.565 116.175 103.795 117.315 ;
        RECT 103.965 116.345 104.295 117.325 ;
        RECT 104.905 117.745 106.135 117.915 ;
        RECT 104.465 116.175 104.675 117.315 ;
        RECT 104.905 116.935 105.245 117.745 ;
        RECT 105.415 117.180 106.165 117.370 ;
        RECT 104.905 116.525 105.420 116.935 ;
        RECT 105.655 116.175 105.825 116.935 ;
        RECT 105.995 116.515 106.165 117.180 ;
        RECT 106.335 117.195 106.525 118.555 ;
        RECT 106.695 117.705 106.970 118.555 ;
        RECT 107.160 118.190 107.690 118.555 ;
        RECT 108.115 118.325 108.445 118.725 ;
        RECT 107.515 118.155 107.690 118.190 ;
        RECT 106.695 117.535 106.975 117.705 ;
        RECT 106.695 117.395 106.970 117.535 ;
        RECT 107.175 117.195 107.345 117.995 ;
        RECT 106.335 117.025 107.345 117.195 ;
        RECT 107.515 117.985 108.445 118.155 ;
        RECT 108.615 117.985 108.870 118.555 ;
        RECT 109.135 118.175 109.305 118.555 ;
        RECT 109.485 118.345 109.815 118.725 ;
        RECT 109.135 118.005 109.800 118.175 ;
        RECT 109.995 118.050 110.255 118.555 ;
        RECT 107.515 116.855 107.685 117.985 ;
        RECT 108.275 117.815 108.445 117.985 ;
        RECT 106.560 116.685 107.685 116.855 ;
        RECT 107.855 117.485 108.050 117.815 ;
        RECT 108.275 117.485 108.530 117.815 ;
        RECT 107.855 116.515 108.025 117.485 ;
        RECT 108.700 117.315 108.870 117.985 ;
        RECT 109.065 117.455 109.395 117.825 ;
        RECT 109.630 117.750 109.800 118.005 ;
        RECT 105.995 116.345 108.025 116.515 ;
        RECT 108.195 116.175 108.365 117.315 ;
        RECT 108.535 116.345 108.870 117.315 ;
        RECT 109.630 117.420 109.915 117.750 ;
        RECT 109.630 117.275 109.800 117.420 ;
        RECT 109.135 117.105 109.800 117.275 ;
        RECT 110.085 117.250 110.255 118.050 ;
        RECT 110.700 117.915 110.945 118.520 ;
        RECT 111.165 118.190 111.675 118.725 ;
        RECT 109.135 116.345 109.305 117.105 ;
        RECT 109.485 116.175 109.815 116.935 ;
        RECT 109.985 116.345 110.255 117.250 ;
        RECT 110.425 117.745 111.655 117.915 ;
        RECT 110.425 116.935 110.765 117.745 ;
        RECT 110.935 117.180 111.685 117.370 ;
        RECT 110.425 116.525 110.940 116.935 ;
        RECT 111.175 116.175 111.345 116.935 ;
        RECT 111.515 116.515 111.685 117.180 ;
        RECT 111.855 117.195 112.045 118.555 ;
        RECT 112.215 118.385 112.490 118.555 ;
        RECT 112.215 118.215 112.495 118.385 ;
        RECT 112.215 117.395 112.490 118.215 ;
        RECT 112.680 118.190 113.210 118.555 ;
        RECT 113.635 118.325 113.965 118.725 ;
        RECT 113.035 118.155 113.210 118.190 ;
        RECT 112.695 117.195 112.865 117.995 ;
        RECT 111.855 117.025 112.865 117.195 ;
        RECT 113.035 117.985 113.965 118.155 ;
        RECT 114.135 117.985 114.390 118.555 ;
        RECT 114.565 118.000 114.855 118.725 ;
        RECT 113.035 116.855 113.205 117.985 ;
        RECT 113.795 117.815 113.965 117.985 ;
        RECT 112.080 116.685 113.205 116.855 ;
        RECT 113.375 117.485 113.570 117.815 ;
        RECT 113.795 117.485 114.050 117.815 ;
        RECT 113.375 116.515 113.545 117.485 ;
        RECT 114.220 117.315 114.390 117.985 ;
        RECT 115.025 117.975 116.235 118.725 ;
        RECT 111.515 116.345 113.545 116.515 ;
        RECT 113.715 116.175 113.885 117.315 ;
        RECT 114.055 116.345 114.390 117.315 ;
        RECT 114.565 116.175 114.855 117.340 ;
        RECT 115.025 117.265 115.545 117.805 ;
        RECT 115.715 117.435 116.235 117.975 ;
        RECT 116.465 117.905 116.675 118.725 ;
        RECT 116.845 117.925 117.175 118.555 ;
        RECT 116.845 117.325 117.095 117.925 ;
        RECT 117.345 117.905 117.575 118.725 ;
        RECT 118.795 118.175 118.965 118.555 ;
        RECT 119.145 118.345 119.475 118.725 ;
        RECT 118.795 118.005 119.460 118.175 ;
        RECT 119.655 118.050 119.915 118.555 ;
        RECT 121.010 118.180 126.355 118.725 ;
        RECT 117.265 117.485 117.595 117.735 ;
        RECT 118.725 117.455 119.055 117.825 ;
        RECT 119.290 117.750 119.460 118.005 ;
        RECT 119.290 117.420 119.575 117.750 ;
        RECT 115.025 116.175 116.235 117.265 ;
        RECT 116.465 116.175 116.675 117.315 ;
        RECT 116.845 116.345 117.175 117.325 ;
        RECT 117.345 116.175 117.575 117.315 ;
        RECT 119.290 117.275 119.460 117.420 ;
        RECT 118.795 117.105 119.460 117.275 ;
        RECT 119.745 117.250 119.915 118.050 ;
        RECT 118.795 116.345 118.965 117.105 ;
        RECT 119.145 116.175 119.475 116.935 ;
        RECT 119.645 116.345 119.915 117.250 ;
        RECT 122.600 116.610 122.950 117.860 ;
        RECT 124.430 117.350 124.770 118.180 ;
        RECT 126.525 117.975 127.735 118.725 ;
        RECT 126.525 117.265 127.045 117.805 ;
        RECT 127.215 117.435 127.735 117.975 ;
        RECT 121.010 116.175 126.355 116.610 ;
        RECT 126.525 116.175 127.735 117.265 ;
        RECT 14.660 116.005 127.820 116.175 ;
        RECT 14.745 114.915 15.955 116.005 ;
        RECT 14.745 114.205 15.265 114.745 ;
        RECT 15.435 114.375 15.955 114.915 ;
        RECT 16.125 114.915 17.335 116.005 ;
        RECT 17.510 115.570 22.855 116.005 ;
        RECT 16.125 114.375 16.645 114.915 ;
        RECT 16.815 114.205 17.335 114.745 ;
        RECT 19.100 114.320 19.450 115.570 ;
        RECT 23.115 115.075 23.285 115.835 ;
        RECT 23.465 115.245 23.795 116.005 ;
        RECT 23.115 114.905 23.780 115.075 ;
        RECT 23.965 114.930 24.235 115.835 ;
        RECT 14.745 113.455 15.955 114.205 ;
        RECT 16.125 113.455 17.335 114.205 ;
        RECT 20.930 114.000 21.270 114.830 ;
        RECT 23.610 114.760 23.780 114.905 ;
        RECT 23.045 114.355 23.375 114.725 ;
        RECT 23.610 114.430 23.895 114.760 ;
        RECT 23.610 114.175 23.780 114.430 ;
        RECT 23.115 114.005 23.780 114.175 ;
        RECT 24.065 114.130 24.235 114.930 ;
        RECT 24.405 114.840 24.695 116.005 ;
        RECT 25.325 114.915 27.915 116.005 ;
        RECT 25.325 114.395 26.535 114.915 ;
        RECT 28.125 114.865 28.355 116.005 ;
        RECT 28.525 114.855 28.855 115.835 ;
        RECT 29.025 114.865 29.235 116.005 ;
        RECT 29.470 114.865 29.805 115.835 ;
        RECT 29.975 114.865 30.145 116.005 ;
        RECT 30.315 115.665 32.345 115.835 ;
        RECT 26.705 114.225 27.915 114.745 ;
        RECT 28.105 114.445 28.435 114.695 ;
        RECT 17.510 113.455 22.855 114.000 ;
        RECT 23.115 113.625 23.285 114.005 ;
        RECT 23.465 113.455 23.795 113.835 ;
        RECT 23.975 113.625 24.235 114.130 ;
        RECT 24.405 113.455 24.695 114.180 ;
        RECT 25.325 113.455 27.915 114.225 ;
        RECT 28.125 113.455 28.355 114.275 ;
        RECT 28.605 114.255 28.855 114.855 ;
        RECT 28.525 113.625 28.855 114.255 ;
        RECT 29.025 113.455 29.235 114.275 ;
        RECT 29.470 114.195 29.640 114.865 ;
        RECT 30.315 114.695 30.485 115.665 ;
        RECT 29.810 114.365 30.065 114.695 ;
        RECT 30.290 114.365 30.485 114.695 ;
        RECT 30.655 115.325 31.780 115.495 ;
        RECT 29.895 114.195 30.065 114.365 ;
        RECT 30.655 114.195 30.825 115.325 ;
        RECT 29.470 113.625 29.725 114.195 ;
        RECT 29.895 114.025 30.825 114.195 ;
        RECT 30.995 114.985 32.005 115.155 ;
        RECT 30.995 114.185 31.165 114.985 ;
        RECT 31.370 114.645 31.645 114.785 ;
        RECT 31.365 114.475 31.645 114.645 ;
        RECT 30.650 113.990 30.825 114.025 ;
        RECT 29.895 113.455 30.225 113.855 ;
        RECT 30.650 113.625 31.180 113.990 ;
        RECT 31.370 113.625 31.645 114.475 ;
        RECT 31.815 113.625 32.005 114.985 ;
        RECT 32.175 115.000 32.345 115.665 ;
        RECT 32.515 115.245 32.685 116.005 ;
        RECT 32.920 115.245 33.435 115.655 ;
        RECT 32.175 114.810 32.925 115.000 ;
        RECT 33.095 114.435 33.435 115.245 ;
        RECT 34.615 115.075 34.785 115.835 ;
        RECT 34.965 115.245 35.295 116.005 ;
        RECT 34.615 114.905 35.280 115.075 ;
        RECT 35.465 114.930 35.735 115.835 ;
        RECT 35.110 114.760 35.280 114.905 ;
        RECT 32.205 114.265 33.435 114.435 ;
        RECT 34.545 114.355 34.875 114.725 ;
        RECT 35.110 114.430 35.395 114.760 ;
        RECT 32.185 113.455 32.695 113.990 ;
        RECT 32.915 113.660 33.160 114.265 ;
        RECT 35.110 114.175 35.280 114.430 ;
        RECT 34.615 114.005 35.280 114.175 ;
        RECT 35.565 114.130 35.735 114.930 ;
        RECT 35.945 114.865 36.175 116.005 ;
        RECT 36.345 114.855 36.675 115.835 ;
        RECT 36.845 114.865 37.055 116.005 ;
        RECT 37.285 114.915 38.955 116.005 ;
        RECT 39.130 115.570 44.475 116.005 ;
        RECT 35.925 114.445 36.255 114.695 ;
        RECT 34.615 113.625 34.785 114.005 ;
        RECT 34.965 113.455 35.295 113.835 ;
        RECT 35.475 113.625 35.735 114.130 ;
        RECT 35.945 113.455 36.175 114.275 ;
        RECT 36.425 114.255 36.675 114.855 ;
        RECT 37.285 114.395 38.035 114.915 ;
        RECT 36.345 113.625 36.675 114.255 ;
        RECT 36.845 113.455 37.055 114.275 ;
        RECT 38.205 114.225 38.955 114.745 ;
        RECT 40.720 114.320 41.070 115.570 ;
        RECT 44.735 115.075 44.905 115.835 ;
        RECT 45.085 115.245 45.415 116.005 ;
        RECT 44.735 114.905 45.400 115.075 ;
        RECT 45.585 114.930 45.855 115.835 ;
        RECT 37.285 113.455 38.955 114.225 ;
        RECT 42.550 114.000 42.890 114.830 ;
        RECT 45.230 114.760 45.400 114.905 ;
        RECT 44.665 114.355 44.995 114.725 ;
        RECT 45.230 114.430 45.515 114.760 ;
        RECT 45.230 114.175 45.400 114.430 ;
        RECT 44.735 114.005 45.400 114.175 ;
        RECT 45.685 114.130 45.855 114.930 ;
        RECT 46.485 114.915 49.995 116.005 ;
        RECT 46.485 114.395 48.175 114.915 ;
        RECT 50.165 114.840 50.455 116.005 ;
        RECT 50.625 114.915 51.835 116.005 ;
        RECT 52.005 114.915 55.515 116.005 ;
        RECT 55.685 115.245 56.200 115.655 ;
        RECT 56.435 115.245 56.605 116.005 ;
        RECT 56.775 115.665 58.805 115.835 ;
        RECT 48.345 114.225 49.995 114.745 ;
        RECT 50.625 114.375 51.145 114.915 ;
        RECT 39.130 113.455 44.475 114.000 ;
        RECT 44.735 113.625 44.905 114.005 ;
        RECT 45.085 113.455 45.415 113.835 ;
        RECT 45.595 113.625 45.855 114.130 ;
        RECT 46.485 113.455 49.995 114.225 ;
        RECT 51.315 114.205 51.835 114.745 ;
        RECT 52.005 114.395 53.695 114.915 ;
        RECT 53.865 114.225 55.515 114.745 ;
        RECT 55.685 114.435 56.025 115.245 ;
        RECT 56.775 115.000 56.945 115.665 ;
        RECT 57.340 115.325 58.465 115.495 ;
        RECT 56.195 114.810 56.945 115.000 ;
        RECT 57.115 114.985 58.125 115.155 ;
        RECT 55.685 114.265 56.915 114.435 ;
        RECT 50.165 113.455 50.455 114.180 ;
        RECT 50.625 113.455 51.835 114.205 ;
        RECT 52.005 113.455 55.515 114.225 ;
        RECT 55.960 113.660 56.205 114.265 ;
        RECT 56.425 113.455 56.935 113.990 ;
        RECT 57.115 113.625 57.305 114.985 ;
        RECT 57.475 114.645 57.750 114.785 ;
        RECT 57.475 114.475 57.755 114.645 ;
        RECT 57.475 113.625 57.750 114.475 ;
        RECT 57.955 114.185 58.125 114.985 ;
        RECT 58.295 114.195 58.465 115.325 ;
        RECT 58.635 114.695 58.805 115.665 ;
        RECT 58.975 114.865 59.145 116.005 ;
        RECT 59.315 114.865 59.650 115.835 ;
        RECT 59.830 115.570 65.175 116.005 ;
        RECT 65.720 115.665 65.975 115.695 ;
        RECT 58.635 114.365 58.830 114.695 ;
        RECT 59.055 114.365 59.310 114.695 ;
        RECT 59.055 114.195 59.225 114.365 ;
        RECT 59.480 114.195 59.650 114.865 ;
        RECT 61.420 114.320 61.770 115.570 ;
        RECT 65.635 115.495 65.975 115.665 ;
        RECT 65.720 115.025 65.975 115.495 ;
        RECT 66.155 115.205 66.440 116.005 ;
        RECT 66.620 115.285 66.950 115.795 ;
        RECT 58.295 114.025 59.225 114.195 ;
        RECT 58.295 113.990 58.470 114.025 ;
        RECT 57.940 113.625 58.470 113.990 ;
        RECT 58.895 113.455 59.225 113.855 ;
        RECT 59.395 113.625 59.650 114.195 ;
        RECT 63.250 114.000 63.590 114.830 ;
        RECT 65.720 114.165 65.900 115.025 ;
        RECT 66.620 114.695 66.870 115.285 ;
        RECT 67.220 115.135 67.390 115.745 ;
        RECT 67.560 115.315 67.890 116.005 ;
        RECT 68.120 115.455 68.360 115.745 ;
        RECT 68.560 115.625 68.980 116.005 ;
        RECT 69.160 115.535 69.790 115.785 ;
        RECT 70.260 115.625 70.590 116.005 ;
        RECT 69.160 115.455 69.330 115.535 ;
        RECT 70.760 115.455 70.930 115.745 ;
        RECT 71.110 115.625 71.490 116.005 ;
        RECT 71.730 115.620 72.560 115.790 ;
        RECT 68.120 115.285 69.330 115.455 ;
        RECT 66.070 114.365 66.870 114.695 ;
        RECT 59.830 113.455 65.175 114.000 ;
        RECT 65.720 113.635 65.975 114.165 ;
        RECT 66.155 113.455 66.440 113.915 ;
        RECT 66.620 113.715 66.870 114.365 ;
        RECT 67.070 115.115 67.390 115.135 ;
        RECT 67.070 114.945 68.990 115.115 ;
        RECT 67.070 114.050 67.260 114.945 ;
        RECT 69.160 114.775 69.330 115.285 ;
        RECT 69.500 115.025 70.020 115.335 ;
        RECT 67.430 114.605 69.330 114.775 ;
        RECT 67.430 114.545 67.760 114.605 ;
        RECT 67.910 114.375 68.240 114.435 ;
        RECT 67.580 114.105 68.240 114.375 ;
        RECT 67.070 113.720 67.390 114.050 ;
        RECT 67.570 113.455 68.230 113.935 ;
        RECT 68.430 113.845 68.600 114.605 ;
        RECT 69.500 114.435 69.680 114.845 ;
        RECT 68.770 114.265 69.100 114.385 ;
        RECT 69.850 114.265 70.020 115.025 ;
        RECT 68.770 114.095 70.020 114.265 ;
        RECT 70.190 115.205 71.560 115.455 ;
        RECT 70.190 114.435 70.380 115.205 ;
        RECT 71.310 114.945 71.560 115.205 ;
        RECT 70.550 114.775 70.800 114.935 ;
        RECT 71.730 114.775 71.900 115.620 ;
        RECT 72.795 115.335 72.965 115.835 ;
        RECT 73.135 115.505 73.465 116.005 ;
        RECT 72.070 114.945 72.570 115.325 ;
        RECT 72.795 115.165 73.490 115.335 ;
        RECT 70.550 114.605 71.900 114.775 ;
        RECT 71.480 114.565 71.900 114.605 ;
        RECT 70.190 114.095 70.610 114.435 ;
        RECT 70.900 114.105 71.310 114.435 ;
        RECT 68.430 113.675 69.280 113.845 ;
        RECT 69.840 113.455 70.160 113.915 ;
        RECT 70.360 113.665 70.610 114.095 ;
        RECT 70.900 113.455 71.310 113.895 ;
        RECT 71.480 113.835 71.650 114.565 ;
        RECT 71.820 114.015 72.170 114.385 ;
        RECT 72.350 114.075 72.570 114.945 ;
        RECT 72.740 114.375 73.150 114.995 ;
        RECT 73.320 114.195 73.490 115.165 ;
        RECT 72.795 114.005 73.490 114.195 ;
        RECT 71.480 113.635 72.495 113.835 ;
        RECT 72.795 113.675 72.965 114.005 ;
        RECT 73.135 113.455 73.465 113.835 ;
        RECT 73.680 113.715 73.905 115.835 ;
        RECT 74.075 115.505 74.405 116.005 ;
        RECT 74.575 115.335 74.745 115.835 ;
        RECT 74.080 115.165 74.745 115.335 ;
        RECT 74.080 114.175 74.310 115.165 ;
        RECT 74.480 114.345 74.830 114.995 ;
        RECT 75.925 114.840 76.215 116.005 ;
        RECT 76.845 114.915 79.435 116.005 ;
        RECT 79.610 115.570 84.955 116.005 ;
        RECT 76.845 114.395 78.055 114.915 ;
        RECT 78.225 114.225 79.435 114.745 ;
        RECT 81.200 114.320 81.550 115.570 ;
        RECT 85.125 115.245 85.640 115.655 ;
        RECT 85.875 115.245 86.045 116.005 ;
        RECT 86.215 115.665 88.245 115.835 ;
        RECT 74.080 114.005 74.745 114.175 ;
        RECT 74.075 113.455 74.405 113.835 ;
        RECT 74.575 113.715 74.745 114.005 ;
        RECT 75.925 113.455 76.215 114.180 ;
        RECT 76.845 113.455 79.435 114.225 ;
        RECT 83.030 114.000 83.370 114.830 ;
        RECT 85.125 114.435 85.465 115.245 ;
        RECT 86.215 115.000 86.385 115.665 ;
        RECT 86.780 115.325 87.905 115.495 ;
        RECT 85.635 114.810 86.385 115.000 ;
        RECT 86.555 114.985 87.565 115.155 ;
        RECT 85.125 114.265 86.355 114.435 ;
        RECT 79.610 113.455 84.955 114.000 ;
        RECT 85.400 113.660 85.645 114.265 ;
        RECT 85.865 113.455 86.375 113.990 ;
        RECT 86.555 113.625 86.745 114.985 ;
        RECT 86.915 114.645 87.190 114.785 ;
        RECT 86.915 114.475 87.195 114.645 ;
        RECT 86.915 113.625 87.190 114.475 ;
        RECT 87.395 114.185 87.565 114.985 ;
        RECT 87.735 114.195 87.905 115.325 ;
        RECT 88.075 114.695 88.245 115.665 ;
        RECT 88.415 114.865 88.585 116.005 ;
        RECT 88.755 114.865 89.090 115.835 ;
        RECT 88.075 114.365 88.270 114.695 ;
        RECT 88.495 114.365 88.750 114.695 ;
        RECT 88.495 114.195 88.665 114.365 ;
        RECT 88.920 114.195 89.090 114.865 ;
        RECT 87.735 114.025 88.665 114.195 ;
        RECT 87.735 113.990 87.910 114.025 ;
        RECT 87.380 113.625 87.910 113.990 ;
        RECT 88.335 113.455 88.665 113.855 ;
        RECT 88.835 113.625 89.090 114.195 ;
        RECT 89.265 114.930 89.535 115.835 ;
        RECT 89.705 115.245 90.035 116.005 ;
        RECT 90.215 115.075 90.385 115.835 ;
        RECT 90.650 115.570 95.995 116.005 ;
        RECT 96.170 115.570 101.515 116.005 ;
        RECT 89.265 114.130 89.435 114.930 ;
        RECT 89.720 114.905 90.385 115.075 ;
        RECT 89.720 114.760 89.890 114.905 ;
        RECT 89.605 114.430 89.890 114.760 ;
        RECT 89.720 114.175 89.890 114.430 ;
        RECT 90.125 114.355 90.455 114.725 ;
        RECT 92.240 114.320 92.590 115.570 ;
        RECT 89.265 113.625 89.525 114.130 ;
        RECT 89.720 114.005 90.385 114.175 ;
        RECT 89.705 113.455 90.035 113.835 ;
        RECT 90.215 113.625 90.385 114.005 ;
        RECT 94.070 114.000 94.410 114.830 ;
        RECT 97.760 114.320 98.110 115.570 ;
        RECT 101.685 114.840 101.975 116.005 ;
        RECT 102.980 115.665 103.235 115.695 ;
        RECT 102.895 115.495 103.235 115.665 ;
        RECT 102.980 115.025 103.235 115.495 ;
        RECT 103.415 115.205 103.700 116.005 ;
        RECT 103.880 115.285 104.210 115.795 ;
        RECT 99.590 114.000 99.930 114.830 ;
        RECT 90.650 113.455 95.995 114.000 ;
        RECT 96.170 113.455 101.515 114.000 ;
        RECT 101.685 113.455 101.975 114.180 ;
        RECT 102.980 114.165 103.160 115.025 ;
        RECT 103.880 114.695 104.130 115.285 ;
        RECT 104.480 115.135 104.650 115.745 ;
        RECT 104.820 115.315 105.150 116.005 ;
        RECT 105.380 115.455 105.620 115.745 ;
        RECT 105.820 115.625 106.240 116.005 ;
        RECT 106.420 115.535 107.050 115.785 ;
        RECT 107.520 115.625 107.850 116.005 ;
        RECT 106.420 115.455 106.590 115.535 ;
        RECT 108.020 115.455 108.190 115.745 ;
        RECT 108.370 115.625 108.750 116.005 ;
        RECT 108.990 115.620 109.820 115.790 ;
        RECT 105.380 115.285 106.590 115.455 ;
        RECT 103.330 114.365 104.130 114.695 ;
        RECT 102.980 113.635 103.235 114.165 ;
        RECT 103.415 113.455 103.700 113.915 ;
        RECT 103.880 113.715 104.130 114.365 ;
        RECT 104.330 115.115 104.650 115.135 ;
        RECT 104.330 114.945 106.250 115.115 ;
        RECT 104.330 114.050 104.520 114.945 ;
        RECT 106.420 114.775 106.590 115.285 ;
        RECT 106.760 115.025 107.280 115.335 ;
        RECT 104.690 114.605 106.590 114.775 ;
        RECT 104.690 114.545 105.020 114.605 ;
        RECT 105.170 114.375 105.500 114.435 ;
        RECT 104.840 114.105 105.500 114.375 ;
        RECT 104.330 113.720 104.650 114.050 ;
        RECT 104.830 113.455 105.490 113.935 ;
        RECT 105.690 113.845 105.860 114.605 ;
        RECT 106.760 114.435 106.940 114.845 ;
        RECT 106.030 114.265 106.360 114.385 ;
        RECT 107.110 114.265 107.280 115.025 ;
        RECT 106.030 114.095 107.280 114.265 ;
        RECT 107.450 115.205 108.820 115.455 ;
        RECT 107.450 114.435 107.640 115.205 ;
        RECT 108.570 114.945 108.820 115.205 ;
        RECT 107.810 114.775 108.060 114.935 ;
        RECT 108.990 114.775 109.160 115.620 ;
        RECT 110.055 115.335 110.225 115.835 ;
        RECT 110.395 115.505 110.725 116.005 ;
        RECT 109.330 114.945 109.830 115.325 ;
        RECT 110.055 115.165 110.750 115.335 ;
        RECT 107.810 114.605 109.160 114.775 ;
        RECT 108.740 114.565 109.160 114.605 ;
        RECT 107.450 114.095 107.870 114.435 ;
        RECT 108.160 114.105 108.570 114.435 ;
        RECT 105.690 113.675 106.540 113.845 ;
        RECT 107.100 113.455 107.420 113.915 ;
        RECT 107.620 113.665 107.870 114.095 ;
        RECT 108.160 113.455 108.570 113.895 ;
        RECT 108.740 113.835 108.910 114.565 ;
        RECT 109.080 114.015 109.430 114.385 ;
        RECT 109.610 114.075 109.830 114.945 ;
        RECT 110.000 114.375 110.410 114.995 ;
        RECT 110.580 114.195 110.750 115.165 ;
        RECT 110.055 114.005 110.750 114.195 ;
        RECT 108.740 113.635 109.755 113.835 ;
        RECT 110.055 113.675 110.225 114.005 ;
        RECT 110.395 113.455 110.725 113.835 ;
        RECT 110.940 113.715 111.165 115.835 ;
        RECT 111.335 115.505 111.665 116.005 ;
        RECT 111.835 115.335 112.005 115.835 ;
        RECT 113.100 115.665 113.355 115.695 ;
        RECT 113.015 115.495 113.355 115.665 ;
        RECT 111.340 115.165 112.005 115.335 ;
        RECT 111.340 114.175 111.570 115.165 ;
        RECT 113.100 115.025 113.355 115.495 ;
        RECT 113.535 115.205 113.820 116.005 ;
        RECT 114.000 115.285 114.330 115.795 ;
        RECT 111.740 114.345 112.090 114.995 ;
        RECT 111.340 114.005 112.005 114.175 ;
        RECT 111.335 113.455 111.665 113.835 ;
        RECT 111.835 113.715 112.005 114.005 ;
        RECT 113.100 114.165 113.280 115.025 ;
        RECT 114.000 114.695 114.250 115.285 ;
        RECT 114.600 115.135 114.770 115.745 ;
        RECT 114.940 115.315 115.270 116.005 ;
        RECT 115.500 115.455 115.740 115.745 ;
        RECT 115.940 115.625 116.360 116.005 ;
        RECT 116.540 115.535 117.170 115.785 ;
        RECT 117.640 115.625 117.970 116.005 ;
        RECT 116.540 115.455 116.710 115.535 ;
        RECT 118.140 115.455 118.310 115.745 ;
        RECT 118.490 115.625 118.870 116.005 ;
        RECT 119.110 115.620 119.940 115.790 ;
        RECT 115.500 115.285 116.710 115.455 ;
        RECT 113.450 114.365 114.250 114.695 ;
        RECT 113.100 113.635 113.355 114.165 ;
        RECT 113.535 113.455 113.820 113.915 ;
        RECT 114.000 113.715 114.250 114.365 ;
        RECT 114.450 115.115 114.770 115.135 ;
        RECT 114.450 114.945 116.370 115.115 ;
        RECT 114.450 114.050 114.640 114.945 ;
        RECT 116.540 114.775 116.710 115.285 ;
        RECT 116.880 115.025 117.400 115.335 ;
        RECT 114.810 114.605 116.710 114.775 ;
        RECT 114.810 114.545 115.140 114.605 ;
        RECT 115.290 114.375 115.620 114.435 ;
        RECT 114.960 114.105 115.620 114.375 ;
        RECT 114.450 113.720 114.770 114.050 ;
        RECT 114.950 113.455 115.610 113.935 ;
        RECT 115.810 113.845 115.980 114.605 ;
        RECT 116.880 114.435 117.060 114.845 ;
        RECT 116.150 114.265 116.480 114.385 ;
        RECT 117.230 114.265 117.400 115.025 ;
        RECT 116.150 114.095 117.400 114.265 ;
        RECT 117.570 115.205 118.940 115.455 ;
        RECT 117.570 114.435 117.760 115.205 ;
        RECT 118.690 114.945 118.940 115.205 ;
        RECT 117.930 114.775 118.180 114.935 ;
        RECT 119.110 114.775 119.280 115.620 ;
        RECT 120.175 115.335 120.345 115.835 ;
        RECT 120.515 115.505 120.845 116.005 ;
        RECT 119.450 114.945 119.950 115.325 ;
        RECT 120.175 115.165 120.870 115.335 ;
        RECT 117.930 114.605 119.280 114.775 ;
        RECT 118.860 114.565 119.280 114.605 ;
        RECT 117.570 114.095 117.990 114.435 ;
        RECT 118.280 114.105 118.690 114.435 ;
        RECT 115.810 113.675 116.660 113.845 ;
        RECT 117.220 113.455 117.540 113.915 ;
        RECT 117.740 113.665 117.990 114.095 ;
        RECT 118.280 113.455 118.690 113.895 ;
        RECT 118.860 113.835 119.030 114.565 ;
        RECT 119.200 114.015 119.550 114.385 ;
        RECT 119.730 114.075 119.950 114.945 ;
        RECT 120.120 114.375 120.530 114.995 ;
        RECT 120.700 114.195 120.870 115.165 ;
        RECT 120.175 114.005 120.870 114.195 ;
        RECT 118.860 113.635 119.875 113.835 ;
        RECT 120.175 113.675 120.345 114.005 ;
        RECT 120.515 113.455 120.845 113.835 ;
        RECT 121.060 113.715 121.285 115.835 ;
        RECT 121.455 115.505 121.785 116.005 ;
        RECT 121.955 115.335 122.125 115.835 ;
        RECT 121.460 115.165 122.125 115.335 ;
        RECT 121.460 114.175 121.690 115.165 ;
        RECT 121.860 114.345 122.210 114.995 ;
        RECT 122.845 114.915 126.355 116.005 ;
        RECT 126.525 114.915 127.735 116.005 ;
        RECT 122.845 114.395 124.535 114.915 ;
        RECT 124.705 114.225 126.355 114.745 ;
        RECT 126.525 114.375 127.045 114.915 ;
        RECT 121.460 114.005 122.125 114.175 ;
        RECT 121.455 113.455 121.785 113.835 ;
        RECT 121.955 113.715 122.125 114.005 ;
        RECT 122.845 113.455 126.355 114.225 ;
        RECT 127.215 114.205 127.735 114.745 ;
        RECT 126.525 113.455 127.735 114.205 ;
        RECT 14.660 113.285 127.820 113.455 ;
        RECT 14.745 112.535 15.955 113.285 ;
        RECT 14.745 111.995 15.265 112.535 ;
        RECT 17.045 112.515 20.555 113.285 ;
        RECT 15.435 111.825 15.955 112.365 ;
        RECT 14.745 110.735 15.955 111.825 ;
        RECT 17.045 111.825 18.735 112.345 ;
        RECT 18.905 111.995 20.555 112.515 ;
        RECT 20.730 112.575 20.985 113.105 ;
        RECT 21.155 112.825 21.460 113.285 ;
        RECT 21.705 112.905 22.775 113.075 ;
        RECT 20.730 111.925 20.940 112.575 ;
        RECT 21.705 112.550 22.025 112.905 ;
        RECT 21.700 112.375 22.025 112.550 ;
        RECT 21.110 112.075 22.025 112.375 ;
        RECT 22.195 112.335 22.435 112.735 ;
        RECT 22.605 112.675 22.775 112.905 ;
        RECT 22.945 112.845 23.135 113.285 ;
        RECT 23.305 112.835 24.255 113.115 ;
        RECT 24.475 112.925 24.825 113.095 ;
        RECT 22.605 112.505 23.135 112.675 ;
        RECT 21.110 112.045 21.850 112.075 ;
        RECT 17.045 110.735 20.555 111.825 ;
        RECT 20.730 111.045 20.985 111.925 ;
        RECT 21.155 110.735 21.460 111.875 ;
        RECT 21.680 111.455 21.850 112.045 ;
        RECT 22.195 111.965 22.735 112.335 ;
        RECT 22.915 112.225 23.135 112.505 ;
        RECT 23.305 112.055 23.475 112.835 ;
        RECT 23.070 111.885 23.475 112.055 ;
        RECT 23.645 112.045 23.995 112.665 ;
        RECT 23.070 111.795 23.240 111.885 ;
        RECT 24.165 111.875 24.375 112.665 ;
        RECT 22.020 111.625 23.240 111.795 ;
        RECT 23.700 111.715 24.375 111.875 ;
        RECT 21.680 111.285 22.480 111.455 ;
        RECT 21.800 110.735 22.130 111.115 ;
        RECT 22.310 110.995 22.480 111.285 ;
        RECT 23.070 111.245 23.240 111.625 ;
        RECT 23.410 111.705 24.375 111.715 ;
        RECT 24.565 112.535 24.825 112.925 ;
        RECT 25.035 112.825 25.365 113.285 ;
        RECT 26.240 112.895 27.095 113.065 ;
        RECT 27.300 112.895 27.795 113.065 ;
        RECT 27.965 112.925 28.295 113.285 ;
        RECT 24.565 111.845 24.735 112.535 ;
        RECT 24.905 112.185 25.075 112.365 ;
        RECT 25.245 112.355 26.035 112.605 ;
        RECT 26.240 112.185 26.410 112.895 ;
        RECT 26.580 112.385 26.935 112.605 ;
        RECT 24.905 112.015 26.595 112.185 ;
        RECT 23.410 111.415 23.870 111.705 ;
        RECT 24.565 111.675 26.065 111.845 ;
        RECT 24.565 111.535 24.735 111.675 ;
        RECT 24.175 111.365 24.735 111.535 ;
        RECT 22.650 110.735 22.900 111.195 ;
        RECT 23.070 110.905 23.940 111.245 ;
        RECT 24.175 110.905 24.345 111.365 ;
        RECT 25.180 111.335 26.255 111.505 ;
        RECT 24.515 110.735 24.885 111.195 ;
        RECT 25.180 110.995 25.350 111.335 ;
        RECT 25.520 110.735 25.850 111.165 ;
        RECT 26.085 110.995 26.255 111.335 ;
        RECT 26.425 111.235 26.595 112.015 ;
        RECT 26.765 111.795 26.935 112.385 ;
        RECT 27.105 111.985 27.455 112.605 ;
        RECT 26.765 111.405 27.230 111.795 ;
        RECT 27.625 111.535 27.795 112.895 ;
        RECT 27.965 111.705 28.425 112.755 ;
        RECT 27.400 111.365 27.795 111.535 ;
        RECT 27.400 111.235 27.570 111.365 ;
        RECT 26.425 110.905 27.105 111.235 ;
        RECT 27.320 110.905 27.570 111.235 ;
        RECT 27.740 110.735 27.990 111.195 ;
        RECT 28.160 110.920 28.485 111.705 ;
        RECT 28.655 110.905 28.825 113.025 ;
        RECT 28.995 112.905 29.325 113.285 ;
        RECT 29.495 112.735 29.750 113.025 ;
        RECT 29.000 112.565 29.750 112.735 ;
        RECT 29.000 111.575 29.230 112.565 ;
        RECT 29.925 112.515 31.595 113.285 ;
        RECT 31.770 112.740 37.115 113.285 ;
        RECT 29.400 111.745 29.750 112.395 ;
        RECT 29.925 111.825 30.675 112.345 ;
        RECT 30.845 111.995 31.595 112.515 ;
        RECT 29.000 111.405 29.750 111.575 ;
        RECT 28.995 110.735 29.325 111.235 ;
        RECT 29.495 110.905 29.750 111.405 ;
        RECT 29.925 110.735 31.595 111.825 ;
        RECT 33.360 111.170 33.710 112.420 ;
        RECT 35.190 111.910 35.530 112.740 ;
        RECT 37.285 112.560 37.575 113.285 ;
        RECT 38.205 112.515 41.715 113.285 ;
        RECT 41.975 112.735 42.145 113.115 ;
        RECT 42.325 112.905 42.655 113.285 ;
        RECT 41.975 112.565 42.640 112.735 ;
        RECT 42.835 112.610 43.095 113.115 ;
        RECT 31.770 110.735 37.115 111.170 ;
        RECT 37.285 110.735 37.575 111.900 ;
        RECT 38.205 111.825 39.895 112.345 ;
        RECT 40.065 111.995 41.715 112.515 ;
        RECT 41.905 112.015 42.235 112.385 ;
        RECT 42.470 112.310 42.640 112.565 ;
        RECT 42.470 111.980 42.755 112.310 ;
        RECT 42.470 111.835 42.640 111.980 ;
        RECT 38.205 110.735 41.715 111.825 ;
        RECT 41.975 111.665 42.640 111.835 ;
        RECT 42.925 111.810 43.095 112.610 ;
        RECT 43.725 112.515 47.235 113.285 ;
        RECT 47.410 112.740 52.755 113.285 ;
        RECT 53.300 112.945 53.555 113.105 ;
        RECT 53.215 112.775 53.555 112.945 ;
        RECT 53.735 112.825 54.020 113.285 ;
        RECT 41.975 110.905 42.145 111.665 ;
        RECT 42.325 110.735 42.655 111.495 ;
        RECT 42.825 110.905 43.095 111.810 ;
        RECT 43.725 111.825 45.415 112.345 ;
        RECT 45.585 111.995 47.235 112.515 ;
        RECT 43.725 110.735 47.235 111.825 ;
        RECT 49.000 111.170 49.350 112.420 ;
        RECT 50.830 111.910 51.170 112.740 ;
        RECT 53.300 112.575 53.555 112.775 ;
        RECT 53.300 111.715 53.480 112.575 ;
        RECT 54.200 112.375 54.450 113.025 ;
        RECT 53.650 112.045 54.450 112.375 ;
        RECT 47.410 110.735 52.755 111.170 ;
        RECT 53.300 111.045 53.555 111.715 ;
        RECT 53.735 110.735 54.020 111.535 ;
        RECT 54.200 111.455 54.450 112.045 ;
        RECT 54.650 112.690 54.970 113.020 ;
        RECT 55.150 112.805 55.810 113.285 ;
        RECT 56.010 112.895 56.860 113.065 ;
        RECT 54.650 111.795 54.840 112.690 ;
        RECT 55.160 112.365 55.820 112.635 ;
        RECT 55.490 112.305 55.820 112.365 ;
        RECT 55.010 112.135 55.340 112.195 ;
        RECT 56.010 112.135 56.180 112.895 ;
        RECT 57.420 112.825 57.740 113.285 ;
        RECT 57.940 112.645 58.190 113.075 ;
        RECT 58.480 112.845 58.890 113.285 ;
        RECT 59.060 112.905 60.075 113.105 ;
        RECT 56.350 112.475 57.600 112.645 ;
        RECT 56.350 112.355 56.680 112.475 ;
        RECT 55.010 111.965 56.910 112.135 ;
        RECT 54.650 111.625 56.570 111.795 ;
        RECT 54.650 111.605 54.970 111.625 ;
        RECT 54.200 110.945 54.530 111.455 ;
        RECT 54.800 110.995 54.970 111.605 ;
        RECT 56.740 111.455 56.910 111.965 ;
        RECT 57.080 111.895 57.260 112.305 ;
        RECT 57.430 111.715 57.600 112.475 ;
        RECT 55.140 110.735 55.470 111.425 ;
        RECT 55.700 111.285 56.910 111.455 ;
        RECT 57.080 111.405 57.600 111.715 ;
        RECT 57.770 112.305 58.190 112.645 ;
        RECT 58.480 112.305 58.890 112.635 ;
        RECT 57.770 111.535 57.960 112.305 ;
        RECT 59.060 112.175 59.230 112.905 ;
        RECT 60.375 112.735 60.545 113.065 ;
        RECT 60.715 112.905 61.045 113.285 ;
        RECT 59.400 112.355 59.750 112.725 ;
        RECT 59.060 112.135 59.480 112.175 ;
        RECT 58.130 111.965 59.480 112.135 ;
        RECT 58.130 111.805 58.380 111.965 ;
        RECT 58.890 111.535 59.140 111.795 ;
        RECT 57.770 111.285 59.140 111.535 ;
        RECT 55.700 110.995 55.940 111.285 ;
        RECT 56.740 111.205 56.910 111.285 ;
        RECT 56.140 110.735 56.560 111.115 ;
        RECT 56.740 110.955 57.370 111.205 ;
        RECT 57.840 110.735 58.170 111.115 ;
        RECT 58.340 110.995 58.510 111.285 ;
        RECT 59.310 111.120 59.480 111.965 ;
        RECT 59.930 111.795 60.150 112.665 ;
        RECT 60.375 112.545 61.070 112.735 ;
        RECT 59.650 111.415 60.150 111.795 ;
        RECT 60.320 111.745 60.730 112.365 ;
        RECT 60.900 111.575 61.070 112.545 ;
        RECT 60.375 111.405 61.070 111.575 ;
        RECT 58.690 110.735 59.070 111.115 ;
        RECT 59.310 110.950 60.140 111.120 ;
        RECT 60.375 110.905 60.545 111.405 ;
        RECT 60.715 110.735 61.045 111.235 ;
        RECT 61.260 110.905 61.485 113.025 ;
        RECT 61.655 112.905 61.985 113.285 ;
        RECT 62.155 112.735 62.325 113.025 ;
        RECT 61.660 112.565 62.325 112.735 ;
        RECT 61.660 111.575 61.890 112.565 ;
        RECT 63.045 112.560 63.335 113.285 ;
        RECT 63.510 112.740 68.855 113.285 ;
        RECT 62.060 111.745 62.410 112.395 ;
        RECT 61.660 111.405 62.325 111.575 ;
        RECT 61.655 110.735 61.985 111.235 ;
        RECT 62.155 110.905 62.325 111.405 ;
        RECT 63.045 110.735 63.335 111.900 ;
        RECT 65.100 111.170 65.450 112.420 ;
        RECT 66.930 111.910 67.270 112.740 ;
        RECT 69.085 112.465 69.295 113.285 ;
        RECT 69.465 112.485 69.795 113.115 ;
        RECT 69.465 111.885 69.715 112.485 ;
        RECT 69.965 112.465 70.195 113.285 ;
        RECT 70.405 112.515 72.075 113.285 ;
        RECT 72.250 112.740 77.595 113.285 ;
        RECT 77.770 112.740 83.115 113.285 ;
        RECT 83.290 112.740 88.635 113.285 ;
        RECT 69.885 112.045 70.215 112.295 ;
        RECT 63.510 110.735 68.855 111.170 ;
        RECT 69.085 110.735 69.295 111.875 ;
        RECT 69.465 110.905 69.795 111.885 ;
        RECT 69.965 110.735 70.195 111.875 ;
        RECT 70.405 111.825 71.155 112.345 ;
        RECT 71.325 111.995 72.075 112.515 ;
        RECT 70.405 110.735 72.075 111.825 ;
        RECT 73.840 111.170 74.190 112.420 ;
        RECT 75.670 111.910 76.010 112.740 ;
        RECT 79.360 111.170 79.710 112.420 ;
        RECT 81.190 111.910 81.530 112.740 ;
        RECT 84.880 111.170 85.230 112.420 ;
        RECT 86.710 111.910 87.050 112.740 ;
        RECT 88.805 112.560 89.095 113.285 ;
        RECT 89.725 112.515 93.235 113.285 ;
        RECT 93.410 112.740 98.755 113.285 ;
        RECT 72.250 110.735 77.595 111.170 ;
        RECT 77.770 110.735 83.115 111.170 ;
        RECT 83.290 110.735 88.635 111.170 ;
        RECT 88.805 110.735 89.095 111.900 ;
        RECT 89.725 111.825 91.415 112.345 ;
        RECT 91.585 111.995 93.235 112.515 ;
        RECT 89.725 110.735 93.235 111.825 ;
        RECT 95.000 111.170 95.350 112.420 ;
        RECT 96.830 111.910 97.170 112.740 ;
        RECT 99.015 112.735 99.185 113.115 ;
        RECT 99.365 112.905 99.695 113.285 ;
        RECT 99.015 112.565 99.680 112.735 ;
        RECT 99.875 112.610 100.135 113.115 ;
        RECT 98.945 112.015 99.275 112.385 ;
        RECT 99.510 112.310 99.680 112.565 ;
        RECT 99.510 111.980 99.795 112.310 ;
        RECT 99.510 111.835 99.680 111.980 ;
        RECT 99.015 111.665 99.680 111.835 ;
        RECT 99.965 111.810 100.135 112.610 ;
        RECT 100.305 112.515 102.895 113.285 ;
        RECT 103.070 112.740 108.415 113.285 ;
        RECT 93.410 110.735 98.755 111.170 ;
        RECT 99.015 110.905 99.185 111.665 ;
        RECT 99.365 110.735 99.695 111.495 ;
        RECT 99.865 110.905 100.135 111.810 ;
        RECT 100.305 111.825 101.515 112.345 ;
        RECT 101.685 111.995 102.895 112.515 ;
        RECT 100.305 110.735 102.895 111.825 ;
        RECT 104.660 111.170 105.010 112.420 ;
        RECT 106.490 111.910 106.830 112.740 ;
        RECT 108.675 112.735 108.845 113.115 ;
        RECT 109.025 112.905 109.355 113.285 ;
        RECT 108.675 112.565 109.340 112.735 ;
        RECT 109.535 112.610 109.795 113.115 ;
        RECT 108.605 112.015 108.935 112.385 ;
        RECT 109.170 112.310 109.340 112.565 ;
        RECT 109.170 111.980 109.455 112.310 ;
        RECT 109.170 111.835 109.340 111.980 ;
        RECT 108.675 111.665 109.340 111.835 ;
        RECT 109.625 111.810 109.795 112.610 ;
        RECT 110.885 112.515 114.395 113.285 ;
        RECT 114.565 112.560 114.855 113.285 ;
        RECT 115.490 112.740 120.835 113.285 ;
        RECT 103.070 110.735 108.415 111.170 ;
        RECT 108.675 110.905 108.845 111.665 ;
        RECT 109.025 110.735 109.355 111.495 ;
        RECT 109.525 110.905 109.795 111.810 ;
        RECT 110.885 111.825 112.575 112.345 ;
        RECT 112.745 111.995 114.395 112.515 ;
        RECT 110.885 110.735 114.395 111.825 ;
        RECT 114.565 110.735 114.855 111.900 ;
        RECT 117.080 111.170 117.430 112.420 ;
        RECT 118.910 111.910 119.250 112.740 ;
        RECT 121.095 112.735 121.265 113.115 ;
        RECT 121.445 112.905 121.775 113.285 ;
        RECT 121.095 112.565 121.760 112.735 ;
        RECT 121.955 112.610 122.215 113.115 ;
        RECT 121.025 112.015 121.355 112.385 ;
        RECT 121.590 112.310 121.760 112.565 ;
        RECT 121.590 111.980 121.875 112.310 ;
        RECT 121.590 111.835 121.760 111.980 ;
        RECT 121.095 111.665 121.760 111.835 ;
        RECT 122.045 111.810 122.215 112.610 ;
        RECT 115.490 110.735 120.835 111.170 ;
        RECT 121.095 110.905 121.265 111.665 ;
        RECT 121.445 110.735 121.775 111.495 ;
        RECT 121.945 110.905 122.215 111.810 ;
        RECT 122.385 112.610 122.645 113.115 ;
        RECT 122.825 112.905 123.155 113.285 ;
        RECT 123.335 112.735 123.505 113.115 ;
        RECT 122.385 111.810 122.555 112.610 ;
        RECT 122.840 112.565 123.505 112.735 ;
        RECT 122.840 112.310 123.010 112.565 ;
        RECT 123.765 112.515 126.355 113.285 ;
        RECT 126.525 112.535 127.735 113.285 ;
        RECT 122.725 111.980 123.010 112.310 ;
        RECT 123.245 112.015 123.575 112.385 ;
        RECT 122.840 111.835 123.010 111.980 ;
        RECT 122.385 110.905 122.655 111.810 ;
        RECT 122.840 111.665 123.505 111.835 ;
        RECT 122.825 110.735 123.155 111.495 ;
        RECT 123.335 110.905 123.505 111.665 ;
        RECT 123.765 111.825 124.975 112.345 ;
        RECT 125.145 111.995 126.355 112.515 ;
        RECT 126.525 111.825 127.045 112.365 ;
        RECT 127.215 111.995 127.735 112.535 ;
        RECT 123.765 110.735 126.355 111.825 ;
        RECT 126.525 110.735 127.735 111.825 ;
        RECT 14.660 110.565 127.820 110.735 ;
        RECT 14.745 109.475 15.955 110.565 ;
        RECT 14.745 108.765 15.265 109.305 ;
        RECT 15.435 108.935 15.955 109.475 ;
        RECT 16.125 109.475 17.335 110.565 ;
        RECT 17.510 110.130 22.855 110.565 ;
        RECT 16.125 108.935 16.645 109.475 ;
        RECT 16.815 108.765 17.335 109.305 ;
        RECT 19.100 108.880 19.450 110.130 ;
        RECT 23.065 109.425 23.295 110.565 ;
        RECT 23.465 109.415 23.795 110.395 ;
        RECT 23.965 109.425 24.175 110.565 ;
        RECT 14.745 108.015 15.955 108.765 ;
        RECT 16.125 108.015 17.335 108.765 ;
        RECT 20.930 108.560 21.270 109.390 ;
        RECT 23.045 109.005 23.375 109.255 ;
        RECT 17.510 108.015 22.855 108.560 ;
        RECT 23.065 108.015 23.295 108.835 ;
        RECT 23.545 108.815 23.795 109.415 ;
        RECT 24.405 109.400 24.695 110.565 ;
        RECT 25.385 109.425 25.595 110.565 ;
        RECT 25.765 109.415 26.095 110.395 ;
        RECT 26.265 109.425 26.495 110.565 ;
        RECT 26.795 109.635 26.965 110.395 ;
        RECT 27.145 109.805 27.475 110.565 ;
        RECT 26.795 109.465 27.460 109.635 ;
        RECT 27.645 109.490 27.915 110.395 ;
        RECT 23.465 108.185 23.795 108.815 ;
        RECT 23.965 108.015 24.175 108.835 ;
        RECT 24.405 108.015 24.695 108.740 ;
        RECT 25.385 108.015 25.595 108.835 ;
        RECT 25.765 108.815 26.015 109.415 ;
        RECT 27.290 109.320 27.460 109.465 ;
        RECT 26.185 109.005 26.515 109.255 ;
        RECT 26.725 108.915 27.055 109.285 ;
        RECT 27.290 108.990 27.575 109.320 ;
        RECT 25.765 108.185 26.095 108.815 ;
        RECT 26.265 108.015 26.495 108.835 ;
        RECT 27.290 108.735 27.460 108.990 ;
        RECT 26.795 108.565 27.460 108.735 ;
        RECT 27.745 108.690 27.915 109.490 ;
        RECT 28.085 109.475 29.755 110.565 ;
        RECT 28.085 108.955 28.835 109.475 ;
        RECT 29.965 109.425 30.195 110.565 ;
        RECT 30.365 109.415 30.695 110.395 ;
        RECT 30.865 109.425 31.075 110.565 ;
        RECT 31.305 109.490 31.575 110.395 ;
        RECT 31.745 109.805 32.075 110.565 ;
        RECT 32.255 109.635 32.425 110.395 ;
        RECT 29.005 108.785 29.755 109.305 ;
        RECT 29.945 109.005 30.275 109.255 ;
        RECT 26.795 108.185 26.965 108.565 ;
        RECT 27.145 108.015 27.475 108.395 ;
        RECT 27.655 108.185 27.915 108.690 ;
        RECT 28.085 108.015 29.755 108.785 ;
        RECT 29.965 108.015 30.195 108.835 ;
        RECT 30.445 108.815 30.695 109.415 ;
        RECT 30.365 108.185 30.695 108.815 ;
        RECT 30.865 108.015 31.075 108.835 ;
        RECT 31.305 108.690 31.475 109.490 ;
        RECT 31.760 109.465 32.425 109.635 ;
        RECT 32.685 109.490 32.955 110.395 ;
        RECT 33.125 109.805 33.455 110.565 ;
        RECT 33.635 109.635 33.805 110.395 ;
        RECT 31.760 109.320 31.930 109.465 ;
        RECT 31.645 108.990 31.930 109.320 ;
        RECT 31.760 108.735 31.930 108.990 ;
        RECT 32.165 108.915 32.495 109.285 ;
        RECT 31.305 108.185 31.565 108.690 ;
        RECT 31.760 108.565 32.425 108.735 ;
        RECT 31.745 108.015 32.075 108.395 ;
        RECT 32.255 108.185 32.425 108.565 ;
        RECT 32.685 108.690 32.855 109.490 ;
        RECT 33.140 109.465 33.805 109.635 ;
        RECT 34.155 109.635 34.325 110.395 ;
        RECT 34.505 109.805 34.835 110.565 ;
        RECT 34.155 109.465 34.820 109.635 ;
        RECT 35.005 109.490 35.275 110.395 ;
        RECT 33.140 109.320 33.310 109.465 ;
        RECT 33.025 108.990 33.310 109.320 ;
        RECT 34.650 109.320 34.820 109.465 ;
        RECT 33.140 108.735 33.310 108.990 ;
        RECT 33.545 108.915 33.875 109.285 ;
        RECT 34.085 108.915 34.415 109.285 ;
        RECT 34.650 108.990 34.935 109.320 ;
        RECT 34.650 108.735 34.820 108.990 ;
        RECT 32.685 108.185 32.945 108.690 ;
        RECT 33.140 108.565 33.805 108.735 ;
        RECT 33.125 108.015 33.455 108.395 ;
        RECT 33.635 108.185 33.805 108.565 ;
        RECT 34.155 108.565 34.820 108.735 ;
        RECT 35.105 108.690 35.275 109.490 ;
        RECT 34.155 108.185 34.325 108.565 ;
        RECT 34.505 108.015 34.835 108.395 ;
        RECT 35.015 108.185 35.275 108.690 ;
        RECT 35.450 109.375 35.705 110.255 ;
        RECT 35.875 109.425 36.180 110.565 ;
        RECT 36.520 110.185 36.850 110.565 ;
        RECT 37.030 110.015 37.200 110.305 ;
        RECT 37.370 110.105 37.620 110.565 ;
        RECT 36.400 109.845 37.200 110.015 ;
        RECT 37.790 110.055 38.660 110.395 ;
        RECT 35.450 108.725 35.660 109.375 ;
        RECT 36.400 109.255 36.570 109.845 ;
        RECT 37.790 109.675 37.960 110.055 ;
        RECT 38.895 109.935 39.065 110.395 ;
        RECT 39.235 110.105 39.605 110.565 ;
        RECT 39.900 109.965 40.070 110.305 ;
        RECT 40.240 110.135 40.570 110.565 ;
        RECT 40.805 109.965 40.975 110.305 ;
        RECT 36.740 109.505 37.960 109.675 ;
        RECT 38.130 109.595 38.590 109.885 ;
        RECT 38.895 109.765 39.455 109.935 ;
        RECT 39.900 109.795 40.975 109.965 ;
        RECT 41.145 110.065 41.825 110.395 ;
        RECT 42.040 110.065 42.290 110.395 ;
        RECT 42.460 110.105 42.710 110.565 ;
        RECT 39.285 109.625 39.455 109.765 ;
        RECT 38.130 109.585 39.095 109.595 ;
        RECT 37.790 109.415 37.960 109.505 ;
        RECT 38.420 109.425 39.095 109.585 ;
        RECT 35.830 109.225 36.570 109.255 ;
        RECT 35.830 108.925 36.745 109.225 ;
        RECT 36.420 108.750 36.745 108.925 ;
        RECT 35.450 108.195 35.705 108.725 ;
        RECT 35.875 108.015 36.180 108.475 ;
        RECT 36.425 108.395 36.745 108.750 ;
        RECT 36.915 108.965 37.455 109.335 ;
        RECT 37.790 109.245 38.195 109.415 ;
        RECT 36.915 108.565 37.155 108.965 ;
        RECT 37.635 108.795 37.855 109.075 ;
        RECT 37.325 108.625 37.855 108.795 ;
        RECT 37.325 108.395 37.495 108.625 ;
        RECT 38.025 108.465 38.195 109.245 ;
        RECT 38.365 108.635 38.715 109.255 ;
        RECT 38.885 108.635 39.095 109.425 ;
        RECT 39.285 109.455 40.785 109.625 ;
        RECT 39.285 108.765 39.455 109.455 ;
        RECT 41.145 109.285 41.315 110.065 ;
        RECT 42.120 109.935 42.290 110.065 ;
        RECT 39.625 109.115 41.315 109.285 ;
        RECT 41.485 109.505 41.950 109.895 ;
        RECT 42.120 109.765 42.515 109.935 ;
        RECT 39.625 108.935 39.795 109.115 ;
        RECT 36.425 108.225 37.495 108.395 ;
        RECT 37.665 108.015 37.855 108.455 ;
        RECT 38.025 108.185 38.975 108.465 ;
        RECT 39.285 108.375 39.545 108.765 ;
        RECT 39.965 108.695 40.755 108.945 ;
        RECT 39.195 108.205 39.545 108.375 ;
        RECT 39.755 108.015 40.085 108.475 ;
        RECT 40.960 108.405 41.130 109.115 ;
        RECT 41.485 108.915 41.655 109.505 ;
        RECT 41.300 108.695 41.655 108.915 ;
        RECT 41.825 108.695 42.175 109.315 ;
        RECT 42.345 108.405 42.515 109.765 ;
        RECT 42.880 109.595 43.205 110.380 ;
        RECT 42.685 108.545 43.145 109.595 ;
        RECT 40.960 108.235 41.815 108.405 ;
        RECT 42.020 108.235 42.515 108.405 ;
        RECT 42.685 108.015 43.015 108.375 ;
        RECT 43.375 108.275 43.545 110.395 ;
        RECT 43.715 110.065 44.045 110.565 ;
        RECT 44.215 109.895 44.470 110.395 ;
        RECT 43.720 109.725 44.470 109.895 ;
        RECT 43.720 108.735 43.950 109.725 ;
        RECT 45.195 109.635 45.365 110.395 ;
        RECT 45.545 109.805 45.875 110.565 ;
        RECT 44.120 108.905 44.470 109.555 ;
        RECT 45.195 109.465 45.860 109.635 ;
        RECT 46.045 109.490 46.315 110.395 ;
        RECT 45.690 109.320 45.860 109.465 ;
        RECT 45.125 108.915 45.455 109.285 ;
        RECT 45.690 108.990 45.975 109.320 ;
        RECT 45.690 108.735 45.860 108.990 ;
        RECT 43.720 108.565 44.470 108.735 ;
        RECT 43.715 108.015 44.045 108.395 ;
        RECT 44.215 108.275 44.470 108.565 ;
        RECT 45.195 108.565 45.860 108.735 ;
        RECT 46.145 108.690 46.315 109.490 ;
        RECT 47.555 109.415 47.885 110.565 ;
        RECT 48.055 109.545 48.225 110.395 ;
        RECT 48.395 109.765 48.725 110.565 ;
        RECT 48.895 109.545 49.065 110.395 ;
        RECT 49.245 109.765 49.485 110.565 ;
        RECT 49.655 109.585 49.985 110.395 ;
        RECT 48.055 109.375 49.065 109.545 ;
        RECT 49.270 109.415 49.985 109.585 ;
        RECT 48.055 108.865 48.550 109.375 ;
        RECT 49.270 109.175 49.440 109.415 ;
        RECT 50.165 109.400 50.455 110.565 ;
        RECT 50.630 110.130 55.975 110.565 ;
        RECT 48.940 109.005 49.440 109.175 ;
        RECT 49.610 109.005 49.990 109.245 ;
        RECT 48.055 108.835 48.555 108.865 ;
        RECT 49.270 108.835 49.440 109.005 ;
        RECT 52.220 108.880 52.570 110.130 ;
        RECT 56.185 109.425 56.415 110.565 ;
        RECT 56.585 109.415 56.915 110.395 ;
        RECT 57.085 109.425 57.295 110.565 ;
        RECT 57.525 109.475 59.195 110.565 ;
        RECT 59.455 109.635 59.625 110.395 ;
        RECT 59.805 109.805 60.135 110.565 ;
        RECT 45.195 108.185 45.365 108.565 ;
        RECT 45.545 108.015 45.875 108.395 ;
        RECT 46.055 108.185 46.315 108.690 ;
        RECT 47.555 108.015 47.885 108.815 ;
        RECT 48.055 108.665 49.065 108.835 ;
        RECT 49.270 108.665 49.905 108.835 ;
        RECT 48.055 108.185 48.225 108.665 ;
        RECT 48.395 108.015 48.725 108.495 ;
        RECT 48.895 108.185 49.065 108.665 ;
        RECT 49.315 108.015 49.555 108.495 ;
        RECT 49.735 108.185 49.905 108.665 ;
        RECT 50.165 108.015 50.455 108.740 ;
        RECT 54.050 108.560 54.390 109.390 ;
        RECT 56.165 109.005 56.495 109.255 ;
        RECT 50.630 108.015 55.975 108.560 ;
        RECT 56.185 108.015 56.415 108.835 ;
        RECT 56.665 108.815 56.915 109.415 ;
        RECT 57.525 108.955 58.275 109.475 ;
        RECT 59.455 109.465 60.120 109.635 ;
        RECT 60.305 109.490 60.575 110.395 ;
        RECT 59.950 109.320 60.120 109.465 ;
        RECT 56.585 108.185 56.915 108.815 ;
        RECT 57.085 108.015 57.295 108.835 ;
        RECT 58.445 108.785 59.195 109.305 ;
        RECT 59.385 108.915 59.715 109.285 ;
        RECT 59.950 108.990 60.235 109.320 ;
        RECT 57.525 108.015 59.195 108.785 ;
        RECT 59.950 108.735 60.120 108.990 ;
        RECT 59.455 108.565 60.120 108.735 ;
        RECT 60.405 108.690 60.575 109.490 ;
        RECT 60.745 109.475 61.955 110.565 ;
        RECT 62.130 110.130 67.475 110.565 ;
        RECT 60.745 108.935 61.265 109.475 ;
        RECT 61.435 108.765 61.955 109.305 ;
        RECT 63.720 108.880 64.070 110.130 ;
        RECT 67.735 109.635 67.905 110.395 ;
        RECT 68.085 109.805 68.415 110.565 ;
        RECT 67.735 109.465 68.400 109.635 ;
        RECT 68.585 109.490 68.855 110.395 ;
        RECT 69.030 110.130 74.375 110.565 ;
        RECT 59.455 108.185 59.625 108.565 ;
        RECT 59.805 108.015 60.135 108.395 ;
        RECT 60.315 108.185 60.575 108.690 ;
        RECT 60.745 108.015 61.955 108.765 ;
        RECT 65.550 108.560 65.890 109.390 ;
        RECT 68.230 109.320 68.400 109.465 ;
        RECT 67.665 108.915 67.995 109.285 ;
        RECT 68.230 108.990 68.515 109.320 ;
        RECT 68.230 108.735 68.400 108.990 ;
        RECT 67.735 108.565 68.400 108.735 ;
        RECT 68.685 108.690 68.855 109.490 ;
        RECT 70.620 108.880 70.970 110.130 ;
        RECT 74.605 109.425 74.815 110.565 ;
        RECT 74.985 109.415 75.315 110.395 ;
        RECT 75.485 109.425 75.715 110.565 ;
        RECT 62.130 108.015 67.475 108.560 ;
        RECT 67.735 108.185 67.905 108.565 ;
        RECT 68.085 108.015 68.415 108.395 ;
        RECT 68.595 108.185 68.855 108.690 ;
        RECT 72.450 108.560 72.790 109.390 ;
        RECT 69.030 108.015 74.375 108.560 ;
        RECT 74.605 108.015 74.815 108.835 ;
        RECT 74.985 108.815 75.235 109.415 ;
        RECT 75.925 109.400 76.215 110.565 ;
        RECT 76.385 109.475 78.055 110.565 ;
        RECT 75.405 109.005 75.735 109.255 ;
        RECT 76.385 108.955 77.135 109.475 ;
        RECT 78.285 109.425 78.495 110.565 ;
        RECT 78.665 109.415 78.995 110.395 ;
        RECT 79.165 109.425 79.395 110.565 ;
        RECT 79.695 109.635 79.865 110.395 ;
        RECT 80.045 109.805 80.375 110.565 ;
        RECT 79.695 109.465 80.360 109.635 ;
        RECT 80.545 109.490 80.815 110.395 ;
        RECT 74.985 108.185 75.315 108.815 ;
        RECT 75.485 108.015 75.715 108.835 ;
        RECT 77.305 108.785 78.055 109.305 ;
        RECT 75.925 108.015 76.215 108.740 ;
        RECT 76.385 108.015 78.055 108.785 ;
        RECT 78.285 108.015 78.495 108.835 ;
        RECT 78.665 108.815 78.915 109.415 ;
        RECT 80.190 109.320 80.360 109.465 ;
        RECT 79.085 109.005 79.415 109.255 ;
        RECT 79.625 108.915 79.955 109.285 ;
        RECT 80.190 108.990 80.475 109.320 ;
        RECT 78.665 108.185 78.995 108.815 ;
        RECT 79.165 108.015 79.395 108.835 ;
        RECT 80.190 108.735 80.360 108.990 ;
        RECT 79.695 108.565 80.360 108.735 ;
        RECT 80.645 108.690 80.815 109.490 ;
        RECT 80.995 109.585 81.325 110.395 ;
        RECT 81.495 109.765 81.735 110.565 ;
        RECT 80.995 109.415 81.710 109.585 ;
        RECT 80.990 109.005 81.370 109.245 ;
        RECT 81.540 109.175 81.710 109.415 ;
        RECT 81.915 109.545 82.085 110.395 ;
        RECT 82.255 109.765 82.585 110.565 ;
        RECT 82.755 109.545 82.925 110.395 ;
        RECT 81.915 109.375 82.925 109.545 ;
        RECT 83.095 109.415 83.425 110.565 ;
        RECT 84.205 109.475 86.795 110.565 ;
        RECT 82.430 109.205 82.925 109.375 ;
        RECT 81.540 109.005 82.040 109.175 ;
        RECT 82.425 109.035 82.925 109.205 ;
        RECT 81.540 108.835 81.710 109.005 ;
        RECT 82.430 108.835 82.925 109.035 ;
        RECT 84.205 108.955 85.415 109.475 ;
        RECT 87.005 109.425 87.235 110.565 ;
        RECT 87.405 109.415 87.735 110.395 ;
        RECT 87.905 109.425 88.115 110.565 ;
        RECT 88.345 109.475 89.555 110.565 ;
        RECT 79.695 108.185 79.865 108.565 ;
        RECT 80.045 108.015 80.375 108.395 ;
        RECT 80.555 108.185 80.815 108.690 ;
        RECT 81.075 108.665 81.710 108.835 ;
        RECT 81.915 108.665 82.925 108.835 ;
        RECT 81.075 108.185 81.245 108.665 ;
        RECT 81.425 108.015 81.665 108.495 ;
        RECT 81.915 108.185 82.085 108.665 ;
        RECT 82.255 108.015 82.585 108.495 ;
        RECT 82.755 108.185 82.925 108.665 ;
        RECT 83.095 108.015 83.425 108.815 ;
        RECT 85.585 108.785 86.795 109.305 ;
        RECT 86.985 109.005 87.315 109.255 ;
        RECT 84.205 108.015 86.795 108.785 ;
        RECT 87.005 108.015 87.235 108.835 ;
        RECT 87.485 108.815 87.735 109.415 ;
        RECT 88.345 108.935 88.865 109.475 ;
        RECT 89.765 109.425 89.995 110.565 ;
        RECT 90.165 109.415 90.495 110.395 ;
        RECT 90.665 109.425 90.875 110.565 ;
        RECT 91.195 109.635 91.365 110.395 ;
        RECT 91.545 109.805 91.875 110.565 ;
        RECT 91.195 109.465 91.860 109.635 ;
        RECT 92.045 109.490 92.315 110.395 ;
        RECT 87.405 108.185 87.735 108.815 ;
        RECT 87.905 108.015 88.115 108.835 ;
        RECT 89.035 108.765 89.555 109.305 ;
        RECT 89.745 109.005 90.075 109.255 ;
        RECT 88.345 108.015 89.555 108.765 ;
        RECT 89.765 108.015 89.995 108.835 ;
        RECT 90.245 108.815 90.495 109.415 ;
        RECT 91.690 109.320 91.860 109.465 ;
        RECT 91.125 108.915 91.455 109.285 ;
        RECT 91.690 108.990 91.975 109.320 ;
        RECT 90.165 108.185 90.495 108.815 ;
        RECT 90.665 108.015 90.875 108.835 ;
        RECT 91.690 108.735 91.860 108.990 ;
        RECT 91.195 108.565 91.860 108.735 ;
        RECT 92.145 108.690 92.315 109.490 ;
        RECT 91.195 108.185 91.365 108.565 ;
        RECT 91.545 108.015 91.875 108.395 ;
        RECT 92.055 108.185 92.315 108.690 ;
        RECT 92.490 109.375 92.745 110.255 ;
        RECT 92.915 109.425 93.220 110.565 ;
        RECT 93.560 110.185 93.890 110.565 ;
        RECT 94.070 110.015 94.240 110.305 ;
        RECT 94.410 110.105 94.660 110.565 ;
        RECT 93.440 109.845 94.240 110.015 ;
        RECT 94.830 110.055 95.700 110.395 ;
        RECT 92.490 108.725 92.700 109.375 ;
        RECT 93.440 109.255 93.610 109.845 ;
        RECT 94.830 109.675 95.000 110.055 ;
        RECT 95.935 109.935 96.105 110.395 ;
        RECT 96.275 110.105 96.645 110.565 ;
        RECT 96.940 109.965 97.110 110.305 ;
        RECT 97.280 110.135 97.610 110.565 ;
        RECT 97.845 109.965 98.015 110.305 ;
        RECT 93.780 109.505 95.000 109.675 ;
        RECT 95.170 109.595 95.630 109.885 ;
        RECT 95.935 109.765 96.495 109.935 ;
        RECT 96.940 109.795 98.015 109.965 ;
        RECT 98.185 110.065 98.865 110.395 ;
        RECT 99.080 110.065 99.330 110.395 ;
        RECT 99.500 110.105 99.750 110.565 ;
        RECT 96.325 109.625 96.495 109.765 ;
        RECT 95.170 109.585 96.135 109.595 ;
        RECT 94.830 109.415 95.000 109.505 ;
        RECT 95.460 109.425 96.135 109.585 ;
        RECT 92.870 109.225 93.610 109.255 ;
        RECT 92.870 108.925 93.785 109.225 ;
        RECT 93.460 108.750 93.785 108.925 ;
        RECT 92.490 108.195 92.745 108.725 ;
        RECT 92.915 108.015 93.220 108.475 ;
        RECT 93.465 108.395 93.785 108.750 ;
        RECT 93.955 108.965 94.495 109.335 ;
        RECT 94.830 109.245 95.235 109.415 ;
        RECT 93.955 108.565 94.195 108.965 ;
        RECT 94.675 108.795 94.895 109.075 ;
        RECT 94.365 108.625 94.895 108.795 ;
        RECT 94.365 108.395 94.535 108.625 ;
        RECT 95.065 108.465 95.235 109.245 ;
        RECT 95.405 108.635 95.755 109.255 ;
        RECT 95.925 108.635 96.135 109.425 ;
        RECT 96.325 109.455 97.825 109.625 ;
        RECT 96.325 108.765 96.495 109.455 ;
        RECT 98.185 109.285 98.355 110.065 ;
        RECT 99.160 109.935 99.330 110.065 ;
        RECT 96.665 109.115 98.355 109.285 ;
        RECT 98.525 109.505 98.990 109.895 ;
        RECT 99.160 109.765 99.555 109.935 ;
        RECT 96.665 108.935 96.835 109.115 ;
        RECT 93.465 108.225 94.535 108.395 ;
        RECT 94.705 108.015 94.895 108.455 ;
        RECT 95.065 108.185 96.015 108.465 ;
        RECT 96.325 108.375 96.585 108.765 ;
        RECT 97.005 108.695 97.795 108.945 ;
        RECT 96.235 108.205 96.585 108.375 ;
        RECT 96.795 108.015 97.125 108.475 ;
        RECT 98.000 108.405 98.170 109.115 ;
        RECT 98.525 108.915 98.695 109.505 ;
        RECT 98.340 108.695 98.695 108.915 ;
        RECT 98.865 108.695 99.215 109.315 ;
        RECT 99.385 108.405 99.555 109.765 ;
        RECT 99.920 109.595 100.245 110.380 ;
        RECT 99.725 108.545 100.185 109.595 ;
        RECT 98.000 108.235 98.855 108.405 ;
        RECT 99.060 108.235 99.555 108.405 ;
        RECT 99.725 108.015 100.055 108.375 ;
        RECT 100.415 108.275 100.585 110.395 ;
        RECT 100.755 110.065 101.085 110.565 ;
        RECT 101.255 109.895 101.510 110.395 ;
        RECT 100.760 109.725 101.510 109.895 ;
        RECT 100.760 108.735 100.990 109.725 ;
        RECT 101.160 108.905 101.510 109.555 ;
        RECT 101.685 109.400 101.975 110.565 ;
        RECT 102.665 109.425 102.875 110.565 ;
        RECT 103.045 109.415 103.375 110.395 ;
        RECT 103.545 109.425 103.775 110.565 ;
        RECT 104.535 109.635 104.705 110.395 ;
        RECT 104.885 109.805 105.215 110.565 ;
        RECT 104.535 109.465 105.200 109.635 ;
        RECT 105.385 109.490 105.655 110.395 ;
        RECT 100.760 108.565 101.510 108.735 ;
        RECT 100.755 108.015 101.085 108.395 ;
        RECT 101.255 108.275 101.510 108.565 ;
        RECT 101.685 108.015 101.975 108.740 ;
        RECT 102.665 108.015 102.875 108.835 ;
        RECT 103.045 108.815 103.295 109.415 ;
        RECT 105.030 109.320 105.200 109.465 ;
        RECT 103.465 109.005 103.795 109.255 ;
        RECT 104.465 108.915 104.795 109.285 ;
        RECT 105.030 108.990 105.315 109.320 ;
        RECT 103.045 108.185 103.375 108.815 ;
        RECT 103.545 108.015 103.775 108.835 ;
        RECT 105.030 108.735 105.200 108.990 ;
        RECT 104.535 108.565 105.200 108.735 ;
        RECT 105.485 108.690 105.655 109.490 ;
        RECT 105.825 109.475 107.035 110.565 ;
        RECT 105.825 108.935 106.345 109.475 ;
        RECT 107.265 109.425 107.475 110.565 ;
        RECT 107.645 109.415 107.975 110.395 ;
        RECT 108.145 109.425 108.375 110.565 ;
        RECT 108.585 109.475 110.255 110.565 ;
        RECT 110.430 110.130 115.775 110.565 ;
        RECT 106.515 108.765 107.035 109.305 ;
        RECT 104.535 108.185 104.705 108.565 ;
        RECT 104.885 108.015 105.215 108.395 ;
        RECT 105.395 108.185 105.655 108.690 ;
        RECT 105.825 108.015 107.035 108.765 ;
        RECT 107.265 108.015 107.475 108.835 ;
        RECT 107.645 108.815 107.895 109.415 ;
        RECT 108.065 109.005 108.395 109.255 ;
        RECT 108.585 108.955 109.335 109.475 ;
        RECT 107.645 108.185 107.975 108.815 ;
        RECT 108.145 108.015 108.375 108.835 ;
        RECT 109.505 108.785 110.255 109.305 ;
        RECT 112.020 108.880 112.370 110.130 ;
        RECT 115.985 109.425 116.215 110.565 ;
        RECT 116.385 109.415 116.715 110.395 ;
        RECT 116.885 109.425 117.095 110.565 ;
        RECT 108.585 108.015 110.255 108.785 ;
        RECT 113.850 108.560 114.190 109.390 ;
        RECT 115.965 109.005 116.295 109.255 ;
        RECT 110.430 108.015 115.775 108.560 ;
        RECT 115.985 108.015 116.215 108.835 ;
        RECT 116.465 108.815 116.715 109.415 ;
        RECT 117.330 109.375 117.585 110.255 ;
        RECT 117.755 109.425 118.060 110.565 ;
        RECT 118.400 110.185 118.730 110.565 ;
        RECT 118.910 110.015 119.080 110.305 ;
        RECT 119.250 110.105 119.500 110.565 ;
        RECT 118.280 109.845 119.080 110.015 ;
        RECT 119.670 110.055 120.540 110.395 ;
        RECT 116.385 108.185 116.715 108.815 ;
        RECT 116.885 108.015 117.095 108.835 ;
        RECT 117.330 108.725 117.540 109.375 ;
        RECT 118.280 109.255 118.450 109.845 ;
        RECT 119.670 109.675 119.840 110.055 ;
        RECT 120.775 109.935 120.945 110.395 ;
        RECT 121.115 110.105 121.485 110.565 ;
        RECT 121.780 109.965 121.950 110.305 ;
        RECT 122.120 110.135 122.450 110.565 ;
        RECT 122.685 109.965 122.855 110.305 ;
        RECT 118.620 109.505 119.840 109.675 ;
        RECT 120.010 109.595 120.470 109.885 ;
        RECT 120.775 109.765 121.335 109.935 ;
        RECT 121.780 109.795 122.855 109.965 ;
        RECT 123.025 110.065 123.705 110.395 ;
        RECT 123.920 110.065 124.170 110.395 ;
        RECT 124.340 110.105 124.590 110.565 ;
        RECT 121.165 109.625 121.335 109.765 ;
        RECT 120.010 109.585 120.975 109.595 ;
        RECT 119.670 109.415 119.840 109.505 ;
        RECT 120.300 109.425 120.975 109.585 ;
        RECT 117.710 109.225 118.450 109.255 ;
        RECT 117.710 108.925 118.625 109.225 ;
        RECT 118.300 108.750 118.625 108.925 ;
        RECT 117.330 108.195 117.585 108.725 ;
        RECT 117.755 108.015 118.060 108.475 ;
        RECT 118.305 108.395 118.625 108.750 ;
        RECT 118.795 108.965 119.335 109.335 ;
        RECT 119.670 109.245 120.075 109.415 ;
        RECT 118.795 108.565 119.035 108.965 ;
        RECT 119.515 108.795 119.735 109.075 ;
        RECT 119.205 108.625 119.735 108.795 ;
        RECT 119.205 108.395 119.375 108.625 ;
        RECT 119.905 108.465 120.075 109.245 ;
        RECT 120.245 108.635 120.595 109.255 ;
        RECT 120.765 108.635 120.975 109.425 ;
        RECT 121.165 109.455 122.665 109.625 ;
        RECT 121.165 108.765 121.335 109.455 ;
        RECT 123.025 109.285 123.195 110.065 ;
        RECT 124.000 109.935 124.170 110.065 ;
        RECT 121.505 109.115 123.195 109.285 ;
        RECT 123.365 109.505 123.830 109.895 ;
        RECT 124.000 109.765 124.395 109.935 ;
        RECT 121.505 108.935 121.675 109.115 ;
        RECT 118.305 108.225 119.375 108.395 ;
        RECT 119.545 108.015 119.735 108.455 ;
        RECT 119.905 108.185 120.855 108.465 ;
        RECT 121.165 108.375 121.425 108.765 ;
        RECT 121.845 108.695 122.635 108.945 ;
        RECT 121.075 108.205 121.425 108.375 ;
        RECT 121.635 108.015 121.965 108.475 ;
        RECT 122.840 108.405 123.010 109.115 ;
        RECT 123.365 108.915 123.535 109.505 ;
        RECT 123.180 108.695 123.535 108.915 ;
        RECT 123.705 108.695 124.055 109.315 ;
        RECT 124.225 108.405 124.395 109.765 ;
        RECT 124.760 109.595 125.085 110.380 ;
        RECT 124.565 108.545 125.025 109.595 ;
        RECT 122.840 108.235 123.695 108.405 ;
        RECT 123.900 108.235 124.395 108.405 ;
        RECT 124.565 108.015 124.895 108.375 ;
        RECT 125.255 108.275 125.425 110.395 ;
        RECT 125.595 110.065 125.925 110.565 ;
        RECT 126.095 109.895 126.350 110.395 ;
        RECT 125.600 109.725 126.350 109.895 ;
        RECT 125.600 108.735 125.830 109.725 ;
        RECT 126.000 108.905 126.350 109.555 ;
        RECT 126.525 109.475 127.735 110.565 ;
        RECT 126.525 108.935 127.045 109.475 ;
        RECT 127.215 108.765 127.735 109.305 ;
        RECT 125.600 108.565 126.350 108.735 ;
        RECT 125.595 108.015 125.925 108.395 ;
        RECT 126.095 108.275 126.350 108.565 ;
        RECT 126.525 108.015 127.735 108.765 ;
        RECT 14.660 107.845 127.820 108.015 ;
        RECT 14.745 107.095 15.955 107.845 ;
        RECT 16.125 107.095 17.335 107.845 ;
        RECT 14.745 106.555 15.265 107.095 ;
        RECT 15.435 106.385 15.955 106.925 ;
        RECT 14.745 105.295 15.955 106.385 ;
        RECT 16.125 106.385 16.645 106.925 ;
        RECT 16.815 106.555 17.335 107.095 ;
        RECT 17.565 107.025 17.775 107.845 ;
        RECT 17.945 107.045 18.275 107.675 ;
        RECT 17.945 106.445 18.195 107.045 ;
        RECT 18.445 107.025 18.675 107.845 ;
        RECT 18.890 107.135 19.145 107.665 ;
        RECT 19.315 107.385 19.620 107.845 ;
        RECT 19.865 107.465 20.935 107.635 ;
        RECT 18.365 106.605 18.695 106.855 ;
        RECT 18.890 106.485 19.100 107.135 ;
        RECT 19.865 107.110 20.185 107.465 ;
        RECT 19.860 106.935 20.185 107.110 ;
        RECT 19.270 106.635 20.185 106.935 ;
        RECT 20.355 106.895 20.595 107.295 ;
        RECT 20.765 107.235 20.935 107.465 ;
        RECT 21.105 107.405 21.295 107.845 ;
        RECT 21.465 107.395 22.415 107.675 ;
        RECT 22.635 107.485 22.985 107.655 ;
        RECT 20.765 107.065 21.295 107.235 ;
        RECT 19.270 106.605 20.010 106.635 ;
        RECT 16.125 105.295 17.335 106.385 ;
        RECT 17.565 105.295 17.775 106.435 ;
        RECT 17.945 105.465 18.275 106.445 ;
        RECT 18.445 105.295 18.675 106.435 ;
        RECT 18.890 105.605 19.145 106.485 ;
        RECT 19.315 105.295 19.620 106.435 ;
        RECT 19.840 106.015 20.010 106.605 ;
        RECT 20.355 106.525 20.895 106.895 ;
        RECT 21.075 106.785 21.295 107.065 ;
        RECT 21.465 106.615 21.635 107.395 ;
        RECT 21.230 106.445 21.635 106.615 ;
        RECT 21.805 106.605 22.155 107.225 ;
        RECT 21.230 106.355 21.400 106.445 ;
        RECT 22.325 106.435 22.535 107.225 ;
        RECT 20.180 106.185 21.400 106.355 ;
        RECT 21.860 106.275 22.535 106.435 ;
        RECT 19.840 105.845 20.640 106.015 ;
        RECT 19.960 105.295 20.290 105.675 ;
        RECT 20.470 105.555 20.640 105.845 ;
        RECT 21.230 105.805 21.400 106.185 ;
        RECT 21.570 106.265 22.535 106.275 ;
        RECT 22.725 107.095 22.985 107.485 ;
        RECT 23.195 107.385 23.525 107.845 ;
        RECT 24.400 107.455 25.255 107.625 ;
        RECT 25.460 107.455 25.955 107.625 ;
        RECT 26.125 107.485 26.455 107.845 ;
        RECT 22.725 106.405 22.895 107.095 ;
        RECT 23.065 106.745 23.235 106.925 ;
        RECT 23.405 106.915 24.195 107.165 ;
        RECT 24.400 106.745 24.570 107.455 ;
        RECT 24.740 106.945 25.095 107.165 ;
        RECT 23.065 106.575 24.755 106.745 ;
        RECT 21.570 105.975 22.030 106.265 ;
        RECT 22.725 106.235 24.225 106.405 ;
        RECT 22.725 106.095 22.895 106.235 ;
        RECT 22.335 105.925 22.895 106.095 ;
        RECT 20.810 105.295 21.060 105.755 ;
        RECT 21.230 105.465 22.100 105.805 ;
        RECT 22.335 105.465 22.505 105.925 ;
        RECT 23.340 105.895 24.415 106.065 ;
        RECT 22.675 105.295 23.045 105.755 ;
        RECT 23.340 105.555 23.510 105.895 ;
        RECT 23.680 105.295 24.010 105.725 ;
        RECT 24.245 105.555 24.415 105.895 ;
        RECT 24.585 105.795 24.755 106.575 ;
        RECT 24.925 106.355 25.095 106.945 ;
        RECT 25.265 106.545 25.615 107.165 ;
        RECT 24.925 105.965 25.390 106.355 ;
        RECT 25.785 106.095 25.955 107.455 ;
        RECT 26.125 106.265 26.585 107.315 ;
        RECT 25.560 105.925 25.955 106.095 ;
        RECT 25.560 105.795 25.730 105.925 ;
        RECT 24.585 105.465 25.265 105.795 ;
        RECT 25.480 105.465 25.730 105.795 ;
        RECT 25.900 105.295 26.150 105.755 ;
        RECT 26.320 105.480 26.645 106.265 ;
        RECT 26.815 105.465 26.985 107.585 ;
        RECT 27.155 107.465 27.485 107.845 ;
        RECT 27.655 107.295 27.910 107.585 ;
        RECT 27.160 107.125 27.910 107.295 ;
        RECT 28.090 107.135 28.345 107.665 ;
        RECT 28.515 107.385 28.820 107.845 ;
        RECT 29.065 107.465 30.135 107.635 ;
        RECT 27.160 106.135 27.390 107.125 ;
        RECT 27.560 106.305 27.910 106.955 ;
        RECT 28.090 106.485 28.300 107.135 ;
        RECT 29.065 107.110 29.385 107.465 ;
        RECT 29.060 106.935 29.385 107.110 ;
        RECT 28.470 106.635 29.385 106.935 ;
        RECT 29.555 106.895 29.795 107.295 ;
        RECT 29.965 107.235 30.135 107.465 ;
        RECT 30.305 107.405 30.495 107.845 ;
        RECT 30.665 107.395 31.615 107.675 ;
        RECT 31.835 107.485 32.185 107.655 ;
        RECT 29.965 107.065 30.495 107.235 ;
        RECT 28.470 106.605 29.210 106.635 ;
        RECT 27.160 105.965 27.910 106.135 ;
        RECT 27.155 105.295 27.485 105.795 ;
        RECT 27.655 105.465 27.910 105.965 ;
        RECT 28.090 105.605 28.345 106.485 ;
        RECT 28.515 105.295 28.820 106.435 ;
        RECT 29.040 106.015 29.210 106.605 ;
        RECT 29.555 106.525 30.095 106.895 ;
        RECT 30.275 106.785 30.495 107.065 ;
        RECT 30.665 106.615 30.835 107.395 ;
        RECT 30.430 106.445 30.835 106.615 ;
        RECT 31.005 106.605 31.355 107.225 ;
        RECT 30.430 106.355 30.600 106.445 ;
        RECT 31.525 106.435 31.735 107.225 ;
        RECT 29.380 106.185 30.600 106.355 ;
        RECT 31.060 106.275 31.735 106.435 ;
        RECT 29.040 105.845 29.840 106.015 ;
        RECT 29.160 105.295 29.490 105.675 ;
        RECT 29.670 105.555 29.840 105.845 ;
        RECT 30.430 105.805 30.600 106.185 ;
        RECT 30.770 106.265 31.735 106.275 ;
        RECT 31.925 107.095 32.185 107.485 ;
        RECT 32.395 107.385 32.725 107.845 ;
        RECT 33.600 107.455 34.455 107.625 ;
        RECT 34.660 107.455 35.155 107.625 ;
        RECT 35.325 107.485 35.655 107.845 ;
        RECT 31.925 106.405 32.095 107.095 ;
        RECT 32.265 106.745 32.435 106.925 ;
        RECT 32.605 106.915 33.395 107.165 ;
        RECT 33.600 106.745 33.770 107.455 ;
        RECT 33.940 106.945 34.295 107.165 ;
        RECT 32.265 106.575 33.955 106.745 ;
        RECT 30.770 105.975 31.230 106.265 ;
        RECT 31.925 106.235 33.425 106.405 ;
        RECT 31.925 106.095 32.095 106.235 ;
        RECT 31.535 105.925 32.095 106.095 ;
        RECT 30.010 105.295 30.260 105.755 ;
        RECT 30.430 105.465 31.300 105.805 ;
        RECT 31.535 105.465 31.705 105.925 ;
        RECT 32.540 105.895 33.615 106.065 ;
        RECT 31.875 105.295 32.245 105.755 ;
        RECT 32.540 105.555 32.710 105.895 ;
        RECT 32.880 105.295 33.210 105.725 ;
        RECT 33.445 105.555 33.615 105.895 ;
        RECT 33.785 105.795 33.955 106.575 ;
        RECT 34.125 106.355 34.295 106.945 ;
        RECT 34.465 106.545 34.815 107.165 ;
        RECT 34.125 105.965 34.590 106.355 ;
        RECT 34.985 106.095 35.155 107.455 ;
        RECT 35.325 106.265 35.785 107.315 ;
        RECT 34.760 105.925 35.155 106.095 ;
        RECT 34.760 105.795 34.930 105.925 ;
        RECT 33.785 105.465 34.465 105.795 ;
        RECT 34.680 105.465 34.930 105.795 ;
        RECT 35.100 105.295 35.350 105.755 ;
        RECT 35.520 105.480 35.845 106.265 ;
        RECT 36.015 105.465 36.185 107.585 ;
        RECT 36.355 107.465 36.685 107.845 ;
        RECT 36.855 107.295 37.110 107.585 ;
        RECT 36.360 107.125 37.110 107.295 ;
        RECT 36.360 106.135 36.590 107.125 ;
        RECT 37.285 107.120 37.575 107.845 ;
        RECT 38.245 107.025 38.475 107.845 ;
        RECT 38.645 107.045 38.975 107.675 ;
        RECT 36.760 106.305 37.110 106.955 ;
        RECT 38.225 106.605 38.555 106.855 ;
        RECT 36.360 105.965 37.110 106.135 ;
        RECT 36.355 105.295 36.685 105.795 ;
        RECT 36.855 105.465 37.110 105.965 ;
        RECT 37.285 105.295 37.575 106.460 ;
        RECT 38.725 106.445 38.975 107.045 ;
        RECT 39.145 107.025 39.355 107.845 ;
        RECT 39.590 107.135 39.845 107.665 ;
        RECT 40.015 107.385 40.320 107.845 ;
        RECT 40.565 107.465 41.635 107.635 ;
        RECT 38.245 105.295 38.475 106.435 ;
        RECT 38.645 105.465 38.975 106.445 ;
        RECT 39.590 106.485 39.800 107.135 ;
        RECT 40.565 107.110 40.885 107.465 ;
        RECT 40.560 106.935 40.885 107.110 ;
        RECT 39.970 106.635 40.885 106.935 ;
        RECT 41.055 106.895 41.295 107.295 ;
        RECT 41.465 107.235 41.635 107.465 ;
        RECT 41.805 107.405 41.995 107.845 ;
        RECT 42.165 107.395 43.115 107.675 ;
        RECT 43.335 107.485 43.685 107.655 ;
        RECT 41.465 107.065 41.995 107.235 ;
        RECT 39.970 106.605 40.710 106.635 ;
        RECT 39.145 105.295 39.355 106.435 ;
        RECT 39.590 105.605 39.845 106.485 ;
        RECT 40.015 105.295 40.320 106.435 ;
        RECT 40.540 106.015 40.710 106.605 ;
        RECT 41.055 106.525 41.595 106.895 ;
        RECT 41.775 106.785 41.995 107.065 ;
        RECT 42.165 106.615 42.335 107.395 ;
        RECT 41.930 106.445 42.335 106.615 ;
        RECT 42.505 106.605 42.855 107.225 ;
        RECT 41.930 106.355 42.100 106.445 ;
        RECT 43.025 106.435 43.235 107.225 ;
        RECT 40.880 106.185 42.100 106.355 ;
        RECT 42.560 106.275 43.235 106.435 ;
        RECT 40.540 105.845 41.340 106.015 ;
        RECT 40.660 105.295 40.990 105.675 ;
        RECT 41.170 105.555 41.340 105.845 ;
        RECT 41.930 105.805 42.100 106.185 ;
        RECT 42.270 106.265 43.235 106.275 ;
        RECT 43.425 107.095 43.685 107.485 ;
        RECT 43.895 107.385 44.225 107.845 ;
        RECT 45.100 107.455 45.955 107.625 ;
        RECT 46.160 107.455 46.655 107.625 ;
        RECT 46.825 107.485 47.155 107.845 ;
        RECT 43.425 106.405 43.595 107.095 ;
        RECT 43.765 106.745 43.935 106.925 ;
        RECT 44.105 106.915 44.895 107.165 ;
        RECT 45.100 106.745 45.270 107.455 ;
        RECT 45.440 106.945 45.795 107.165 ;
        RECT 43.765 106.575 45.455 106.745 ;
        RECT 42.270 105.975 42.730 106.265 ;
        RECT 43.425 106.235 44.925 106.405 ;
        RECT 43.425 106.095 43.595 106.235 ;
        RECT 43.035 105.925 43.595 106.095 ;
        RECT 41.510 105.295 41.760 105.755 ;
        RECT 41.930 105.465 42.800 105.805 ;
        RECT 43.035 105.465 43.205 105.925 ;
        RECT 44.040 105.895 45.115 106.065 ;
        RECT 43.375 105.295 43.745 105.755 ;
        RECT 44.040 105.555 44.210 105.895 ;
        RECT 44.380 105.295 44.710 105.725 ;
        RECT 44.945 105.555 45.115 105.895 ;
        RECT 45.285 105.795 45.455 106.575 ;
        RECT 45.625 106.355 45.795 106.945 ;
        RECT 45.965 106.545 46.315 107.165 ;
        RECT 45.625 105.965 46.090 106.355 ;
        RECT 46.485 106.095 46.655 107.455 ;
        RECT 46.825 106.265 47.285 107.315 ;
        RECT 46.260 105.925 46.655 106.095 ;
        RECT 46.260 105.795 46.430 105.925 ;
        RECT 45.285 105.465 45.965 105.795 ;
        RECT 46.180 105.465 46.430 105.795 ;
        RECT 46.600 105.295 46.850 105.755 ;
        RECT 47.020 105.480 47.345 106.265 ;
        RECT 47.515 105.465 47.685 107.585 ;
        RECT 47.855 107.465 48.185 107.845 ;
        RECT 48.355 107.295 48.610 107.585 ;
        RECT 47.860 107.125 48.610 107.295 ;
        RECT 48.785 107.170 49.045 107.675 ;
        RECT 49.225 107.465 49.555 107.845 ;
        RECT 49.735 107.295 49.905 107.675 ;
        RECT 47.860 106.135 48.090 107.125 ;
        RECT 48.260 106.305 48.610 106.955 ;
        RECT 48.785 106.370 48.955 107.170 ;
        RECT 49.240 107.125 49.905 107.295 ;
        RECT 49.240 106.870 49.410 107.125 ;
        RECT 50.165 107.095 51.375 107.845 ;
        RECT 51.635 107.295 51.805 107.675 ;
        RECT 51.985 107.465 52.315 107.845 ;
        RECT 51.635 107.125 52.300 107.295 ;
        RECT 52.495 107.170 52.755 107.675 ;
        RECT 49.125 106.540 49.410 106.870 ;
        RECT 49.645 106.575 49.975 106.945 ;
        RECT 49.240 106.395 49.410 106.540 ;
        RECT 47.860 105.965 48.610 106.135 ;
        RECT 47.855 105.295 48.185 105.795 ;
        RECT 48.355 105.465 48.610 105.965 ;
        RECT 48.785 105.465 49.055 106.370 ;
        RECT 49.240 106.225 49.905 106.395 ;
        RECT 49.225 105.295 49.555 106.055 ;
        RECT 49.735 105.465 49.905 106.225 ;
        RECT 50.165 106.385 50.685 106.925 ;
        RECT 50.855 106.555 51.375 107.095 ;
        RECT 51.565 106.575 51.895 106.945 ;
        RECT 52.130 106.870 52.300 107.125 ;
        RECT 52.130 106.540 52.415 106.870 ;
        RECT 52.130 106.395 52.300 106.540 ;
        RECT 50.165 105.295 51.375 106.385 ;
        RECT 51.635 106.225 52.300 106.395 ;
        RECT 52.585 106.370 52.755 107.170 ;
        RECT 51.635 105.465 51.805 106.225 ;
        RECT 51.985 105.295 52.315 106.055 ;
        RECT 52.485 105.465 52.755 106.370 ;
        RECT 53.845 107.170 54.105 107.675 ;
        RECT 54.285 107.465 54.615 107.845 ;
        RECT 54.795 107.295 54.965 107.675 ;
        RECT 53.845 106.370 54.015 107.170 ;
        RECT 54.300 107.125 54.965 107.295 ;
        RECT 54.300 106.870 54.470 107.125 ;
        RECT 55.725 107.025 55.955 107.845 ;
        RECT 56.125 107.045 56.455 107.675 ;
        RECT 54.185 106.540 54.470 106.870 ;
        RECT 54.705 106.575 55.035 106.945 ;
        RECT 55.705 106.605 56.035 106.855 ;
        RECT 54.300 106.395 54.470 106.540 ;
        RECT 56.205 106.445 56.455 107.045 ;
        RECT 56.625 107.025 56.835 107.845 ;
        RECT 57.985 107.075 61.495 107.845 ;
        RECT 53.845 105.465 54.115 106.370 ;
        RECT 54.300 106.225 54.965 106.395 ;
        RECT 54.285 105.295 54.615 106.055 ;
        RECT 54.795 105.465 54.965 106.225 ;
        RECT 55.725 105.295 55.955 106.435 ;
        RECT 56.125 105.465 56.455 106.445 ;
        RECT 56.625 105.295 56.835 106.435 ;
        RECT 57.985 106.385 59.675 106.905 ;
        RECT 59.845 106.555 61.495 107.075 ;
        RECT 61.705 107.025 61.935 107.845 ;
        RECT 62.105 107.045 62.435 107.675 ;
        RECT 61.685 106.605 62.015 106.855 ;
        RECT 62.185 106.445 62.435 107.045 ;
        RECT 62.605 107.025 62.815 107.845 ;
        RECT 63.045 107.120 63.335 107.845 ;
        RECT 63.510 107.135 63.765 107.665 ;
        RECT 63.935 107.385 64.240 107.845 ;
        RECT 64.485 107.465 65.555 107.635 ;
        RECT 63.510 106.485 63.720 107.135 ;
        RECT 64.485 107.110 64.805 107.465 ;
        RECT 64.480 106.935 64.805 107.110 ;
        RECT 63.890 106.635 64.805 106.935 ;
        RECT 64.975 106.895 65.215 107.295 ;
        RECT 65.385 107.235 65.555 107.465 ;
        RECT 65.725 107.405 65.915 107.845 ;
        RECT 66.085 107.395 67.035 107.675 ;
        RECT 67.255 107.485 67.605 107.655 ;
        RECT 65.385 107.065 65.915 107.235 ;
        RECT 63.890 106.605 64.630 106.635 ;
        RECT 57.985 105.295 61.495 106.385 ;
        RECT 61.705 105.295 61.935 106.435 ;
        RECT 62.105 105.465 62.435 106.445 ;
        RECT 62.605 105.295 62.815 106.435 ;
        RECT 63.045 105.295 63.335 106.460 ;
        RECT 63.510 105.605 63.765 106.485 ;
        RECT 63.935 105.295 64.240 106.435 ;
        RECT 64.460 106.015 64.630 106.605 ;
        RECT 64.975 106.525 65.515 106.895 ;
        RECT 65.695 106.785 65.915 107.065 ;
        RECT 66.085 106.615 66.255 107.395 ;
        RECT 65.850 106.445 66.255 106.615 ;
        RECT 66.425 106.605 66.775 107.225 ;
        RECT 65.850 106.355 66.020 106.445 ;
        RECT 66.945 106.435 67.155 107.225 ;
        RECT 64.800 106.185 66.020 106.355 ;
        RECT 66.480 106.275 67.155 106.435 ;
        RECT 64.460 105.845 65.260 106.015 ;
        RECT 64.580 105.295 64.910 105.675 ;
        RECT 65.090 105.555 65.260 105.845 ;
        RECT 65.850 105.805 66.020 106.185 ;
        RECT 66.190 106.265 67.155 106.275 ;
        RECT 67.345 107.095 67.605 107.485 ;
        RECT 67.815 107.385 68.145 107.845 ;
        RECT 69.020 107.455 69.875 107.625 ;
        RECT 70.080 107.455 70.575 107.625 ;
        RECT 70.745 107.485 71.075 107.845 ;
        RECT 67.345 106.405 67.515 107.095 ;
        RECT 67.685 106.745 67.855 106.925 ;
        RECT 68.025 106.915 68.815 107.165 ;
        RECT 69.020 106.745 69.190 107.455 ;
        RECT 69.360 106.945 69.715 107.165 ;
        RECT 67.685 106.575 69.375 106.745 ;
        RECT 66.190 105.975 66.650 106.265 ;
        RECT 67.345 106.235 68.845 106.405 ;
        RECT 67.345 106.095 67.515 106.235 ;
        RECT 66.955 105.925 67.515 106.095 ;
        RECT 65.430 105.295 65.680 105.755 ;
        RECT 65.850 105.465 66.720 105.805 ;
        RECT 66.955 105.465 67.125 105.925 ;
        RECT 67.960 105.895 69.035 106.065 ;
        RECT 67.295 105.295 67.665 105.755 ;
        RECT 67.960 105.555 68.130 105.895 ;
        RECT 68.300 105.295 68.630 105.725 ;
        RECT 68.865 105.555 69.035 105.895 ;
        RECT 69.205 105.795 69.375 106.575 ;
        RECT 69.545 106.355 69.715 106.945 ;
        RECT 69.885 106.545 70.235 107.165 ;
        RECT 69.545 105.965 70.010 106.355 ;
        RECT 70.405 106.095 70.575 107.455 ;
        RECT 70.745 106.265 71.205 107.315 ;
        RECT 70.180 105.925 70.575 106.095 ;
        RECT 70.180 105.795 70.350 105.925 ;
        RECT 69.205 105.465 69.885 105.795 ;
        RECT 70.100 105.465 70.350 105.795 ;
        RECT 70.520 105.295 70.770 105.755 ;
        RECT 70.940 105.480 71.265 106.265 ;
        RECT 71.435 105.465 71.605 107.585 ;
        RECT 71.775 107.465 72.105 107.845 ;
        RECT 72.275 107.295 72.530 107.585 ;
        RECT 71.780 107.125 72.530 107.295 ;
        RECT 73.630 107.135 73.885 107.665 ;
        RECT 74.055 107.385 74.360 107.845 ;
        RECT 74.605 107.465 75.675 107.635 ;
        RECT 71.780 106.135 72.010 107.125 ;
        RECT 72.180 106.305 72.530 106.955 ;
        RECT 73.630 106.485 73.840 107.135 ;
        RECT 74.605 107.110 74.925 107.465 ;
        RECT 74.600 106.935 74.925 107.110 ;
        RECT 74.010 106.635 74.925 106.935 ;
        RECT 75.095 106.895 75.335 107.295 ;
        RECT 75.505 107.235 75.675 107.465 ;
        RECT 75.845 107.405 76.035 107.845 ;
        RECT 76.205 107.395 77.155 107.675 ;
        RECT 77.375 107.485 77.725 107.655 ;
        RECT 75.505 107.065 76.035 107.235 ;
        RECT 74.010 106.605 74.750 106.635 ;
        RECT 71.780 105.965 72.530 106.135 ;
        RECT 71.775 105.295 72.105 105.795 ;
        RECT 72.275 105.465 72.530 105.965 ;
        RECT 73.630 105.605 73.885 106.485 ;
        RECT 74.055 105.295 74.360 106.435 ;
        RECT 74.580 106.015 74.750 106.605 ;
        RECT 75.095 106.525 75.635 106.895 ;
        RECT 75.815 106.785 76.035 107.065 ;
        RECT 76.205 106.615 76.375 107.395 ;
        RECT 75.970 106.445 76.375 106.615 ;
        RECT 76.545 106.605 76.895 107.225 ;
        RECT 75.970 106.355 76.140 106.445 ;
        RECT 77.065 106.435 77.275 107.225 ;
        RECT 74.920 106.185 76.140 106.355 ;
        RECT 76.600 106.275 77.275 106.435 ;
        RECT 74.580 105.845 75.380 106.015 ;
        RECT 74.700 105.295 75.030 105.675 ;
        RECT 75.210 105.555 75.380 105.845 ;
        RECT 75.970 105.805 76.140 106.185 ;
        RECT 76.310 106.265 77.275 106.275 ;
        RECT 77.465 107.095 77.725 107.485 ;
        RECT 77.935 107.385 78.265 107.845 ;
        RECT 79.140 107.455 79.995 107.625 ;
        RECT 80.200 107.455 80.695 107.625 ;
        RECT 80.865 107.485 81.195 107.845 ;
        RECT 77.465 106.405 77.635 107.095 ;
        RECT 77.805 106.745 77.975 106.925 ;
        RECT 78.145 106.915 78.935 107.165 ;
        RECT 79.140 106.745 79.310 107.455 ;
        RECT 79.480 106.945 79.835 107.165 ;
        RECT 77.805 106.575 79.495 106.745 ;
        RECT 76.310 105.975 76.770 106.265 ;
        RECT 77.465 106.235 78.965 106.405 ;
        RECT 77.465 106.095 77.635 106.235 ;
        RECT 77.075 105.925 77.635 106.095 ;
        RECT 75.550 105.295 75.800 105.755 ;
        RECT 75.970 105.465 76.840 105.805 ;
        RECT 77.075 105.465 77.245 105.925 ;
        RECT 78.080 105.895 79.155 106.065 ;
        RECT 77.415 105.295 77.785 105.755 ;
        RECT 78.080 105.555 78.250 105.895 ;
        RECT 78.420 105.295 78.750 105.725 ;
        RECT 78.985 105.555 79.155 105.895 ;
        RECT 79.325 105.795 79.495 106.575 ;
        RECT 79.665 106.355 79.835 106.945 ;
        RECT 80.005 106.545 80.355 107.165 ;
        RECT 79.665 105.965 80.130 106.355 ;
        RECT 80.525 106.095 80.695 107.455 ;
        RECT 80.865 106.265 81.325 107.315 ;
        RECT 80.300 105.925 80.695 106.095 ;
        RECT 80.300 105.795 80.470 105.925 ;
        RECT 79.325 105.465 80.005 105.795 ;
        RECT 80.220 105.465 80.470 105.795 ;
        RECT 80.640 105.295 80.890 105.755 ;
        RECT 81.060 105.480 81.385 106.265 ;
        RECT 81.555 105.465 81.725 107.585 ;
        RECT 81.895 107.465 82.225 107.845 ;
        RECT 82.395 107.295 82.650 107.585 ;
        RECT 81.900 107.125 82.650 107.295 ;
        RECT 82.915 107.295 83.085 107.675 ;
        RECT 83.265 107.465 83.595 107.845 ;
        RECT 82.915 107.125 83.580 107.295 ;
        RECT 83.775 107.170 84.035 107.675 ;
        RECT 81.900 106.135 82.130 107.125 ;
        RECT 82.300 106.305 82.650 106.955 ;
        RECT 82.845 106.575 83.175 106.945 ;
        RECT 83.410 106.870 83.580 107.125 ;
        RECT 83.410 106.540 83.695 106.870 ;
        RECT 83.410 106.395 83.580 106.540 ;
        RECT 82.915 106.225 83.580 106.395 ;
        RECT 83.865 106.370 84.035 107.170 ;
        RECT 84.265 107.025 84.475 107.845 ;
        RECT 84.645 107.045 84.975 107.675 ;
        RECT 84.645 106.445 84.895 107.045 ;
        RECT 85.145 107.025 85.375 107.845 ;
        RECT 86.595 107.295 86.765 107.675 ;
        RECT 86.945 107.465 87.275 107.845 ;
        RECT 86.595 107.125 87.260 107.295 ;
        RECT 87.455 107.170 87.715 107.675 ;
        RECT 85.065 106.605 85.395 106.855 ;
        RECT 86.525 106.575 86.855 106.945 ;
        RECT 87.090 106.870 87.260 107.125 ;
        RECT 87.090 106.540 87.375 106.870 ;
        RECT 81.900 105.965 82.650 106.135 ;
        RECT 81.895 105.295 82.225 105.795 ;
        RECT 82.395 105.465 82.650 105.965 ;
        RECT 82.915 105.465 83.085 106.225 ;
        RECT 83.265 105.295 83.595 106.055 ;
        RECT 83.765 105.465 84.035 106.370 ;
        RECT 84.265 105.295 84.475 106.435 ;
        RECT 84.645 105.465 84.975 106.445 ;
        RECT 85.145 105.295 85.375 106.435 ;
        RECT 87.090 106.395 87.260 106.540 ;
        RECT 86.595 106.225 87.260 106.395 ;
        RECT 87.545 106.370 87.715 107.170 ;
        RECT 88.805 107.120 89.095 107.845 ;
        RECT 89.270 107.135 89.525 107.665 ;
        RECT 89.695 107.385 90.000 107.845 ;
        RECT 90.245 107.465 91.315 107.635 ;
        RECT 89.270 106.485 89.480 107.135 ;
        RECT 90.245 107.110 90.565 107.465 ;
        RECT 90.240 106.935 90.565 107.110 ;
        RECT 89.650 106.635 90.565 106.935 ;
        RECT 90.735 106.895 90.975 107.295 ;
        RECT 91.145 107.235 91.315 107.465 ;
        RECT 91.485 107.405 91.675 107.845 ;
        RECT 91.845 107.395 92.795 107.675 ;
        RECT 93.015 107.485 93.365 107.655 ;
        RECT 91.145 107.065 91.675 107.235 ;
        RECT 89.650 106.605 90.390 106.635 ;
        RECT 86.595 105.465 86.765 106.225 ;
        RECT 86.945 105.295 87.275 106.055 ;
        RECT 87.445 105.465 87.715 106.370 ;
        RECT 88.805 105.295 89.095 106.460 ;
        RECT 89.270 105.605 89.525 106.485 ;
        RECT 89.695 105.295 90.000 106.435 ;
        RECT 90.220 106.015 90.390 106.605 ;
        RECT 90.735 106.525 91.275 106.895 ;
        RECT 91.455 106.785 91.675 107.065 ;
        RECT 91.845 106.615 92.015 107.395 ;
        RECT 91.610 106.445 92.015 106.615 ;
        RECT 92.185 106.605 92.535 107.225 ;
        RECT 91.610 106.355 91.780 106.445 ;
        RECT 92.705 106.435 92.915 107.225 ;
        RECT 90.560 106.185 91.780 106.355 ;
        RECT 92.240 106.275 92.915 106.435 ;
        RECT 90.220 105.845 91.020 106.015 ;
        RECT 90.340 105.295 90.670 105.675 ;
        RECT 90.850 105.555 91.020 105.845 ;
        RECT 91.610 105.805 91.780 106.185 ;
        RECT 91.950 106.265 92.915 106.275 ;
        RECT 93.105 107.095 93.365 107.485 ;
        RECT 93.575 107.385 93.905 107.845 ;
        RECT 94.780 107.455 95.635 107.625 ;
        RECT 95.840 107.455 96.335 107.625 ;
        RECT 96.505 107.485 96.835 107.845 ;
        RECT 93.105 106.405 93.275 107.095 ;
        RECT 93.445 106.745 93.615 106.925 ;
        RECT 93.785 106.915 94.575 107.165 ;
        RECT 94.780 106.745 94.950 107.455 ;
        RECT 95.120 106.945 95.475 107.165 ;
        RECT 93.445 106.575 95.135 106.745 ;
        RECT 91.950 105.975 92.410 106.265 ;
        RECT 93.105 106.235 94.605 106.405 ;
        RECT 93.105 106.095 93.275 106.235 ;
        RECT 92.715 105.925 93.275 106.095 ;
        RECT 91.190 105.295 91.440 105.755 ;
        RECT 91.610 105.465 92.480 105.805 ;
        RECT 92.715 105.465 92.885 105.925 ;
        RECT 93.720 105.895 94.795 106.065 ;
        RECT 93.055 105.295 93.425 105.755 ;
        RECT 93.720 105.555 93.890 105.895 ;
        RECT 94.060 105.295 94.390 105.725 ;
        RECT 94.625 105.555 94.795 105.895 ;
        RECT 94.965 105.795 95.135 106.575 ;
        RECT 95.305 106.355 95.475 106.945 ;
        RECT 95.645 106.545 95.995 107.165 ;
        RECT 95.305 105.965 95.770 106.355 ;
        RECT 96.165 106.095 96.335 107.455 ;
        RECT 96.505 106.265 96.965 107.315 ;
        RECT 95.940 105.925 96.335 106.095 ;
        RECT 95.940 105.795 96.110 105.925 ;
        RECT 94.965 105.465 95.645 105.795 ;
        RECT 95.860 105.465 96.110 105.795 ;
        RECT 96.280 105.295 96.530 105.755 ;
        RECT 96.700 105.480 97.025 106.265 ;
        RECT 97.195 105.465 97.365 107.585 ;
        RECT 97.535 107.465 97.865 107.845 ;
        RECT 98.035 107.295 98.290 107.585 ;
        RECT 97.540 107.125 98.290 107.295 ;
        RECT 97.540 106.135 97.770 107.125 ;
        RECT 98.525 107.025 98.735 107.845 ;
        RECT 98.905 107.045 99.235 107.675 ;
        RECT 97.940 106.305 98.290 106.955 ;
        RECT 98.905 106.445 99.155 107.045 ;
        RECT 99.405 107.025 99.635 107.845 ;
        RECT 99.850 107.135 100.105 107.665 ;
        RECT 100.275 107.385 100.580 107.845 ;
        RECT 100.825 107.465 101.895 107.635 ;
        RECT 99.325 106.605 99.655 106.855 ;
        RECT 99.850 106.485 100.060 107.135 ;
        RECT 100.825 107.110 101.145 107.465 ;
        RECT 100.820 106.935 101.145 107.110 ;
        RECT 100.230 106.635 101.145 106.935 ;
        RECT 101.315 106.895 101.555 107.295 ;
        RECT 101.725 107.235 101.895 107.465 ;
        RECT 102.065 107.405 102.255 107.845 ;
        RECT 102.425 107.395 103.375 107.675 ;
        RECT 103.595 107.485 103.945 107.655 ;
        RECT 101.725 107.065 102.255 107.235 ;
        RECT 100.230 106.605 100.970 106.635 ;
        RECT 97.540 105.965 98.290 106.135 ;
        RECT 97.535 105.295 97.865 105.795 ;
        RECT 98.035 105.465 98.290 105.965 ;
        RECT 98.525 105.295 98.735 106.435 ;
        RECT 98.905 105.465 99.235 106.445 ;
        RECT 99.405 105.295 99.635 106.435 ;
        RECT 99.850 105.605 100.105 106.485 ;
        RECT 100.275 105.295 100.580 106.435 ;
        RECT 100.800 106.015 100.970 106.605 ;
        RECT 101.315 106.525 101.855 106.895 ;
        RECT 102.035 106.785 102.255 107.065 ;
        RECT 102.425 106.615 102.595 107.395 ;
        RECT 102.190 106.445 102.595 106.615 ;
        RECT 102.765 106.605 103.115 107.225 ;
        RECT 102.190 106.355 102.360 106.445 ;
        RECT 103.285 106.435 103.495 107.225 ;
        RECT 101.140 106.185 102.360 106.355 ;
        RECT 102.820 106.275 103.495 106.435 ;
        RECT 100.800 105.845 101.600 106.015 ;
        RECT 100.920 105.295 101.250 105.675 ;
        RECT 101.430 105.555 101.600 105.845 ;
        RECT 102.190 105.805 102.360 106.185 ;
        RECT 102.530 106.265 103.495 106.275 ;
        RECT 103.685 107.095 103.945 107.485 ;
        RECT 104.155 107.385 104.485 107.845 ;
        RECT 105.360 107.455 106.215 107.625 ;
        RECT 106.420 107.455 106.915 107.625 ;
        RECT 107.085 107.485 107.415 107.845 ;
        RECT 103.685 106.405 103.855 107.095 ;
        RECT 104.025 106.745 104.195 106.925 ;
        RECT 104.365 106.915 105.155 107.165 ;
        RECT 105.360 106.745 105.530 107.455 ;
        RECT 105.700 106.945 106.055 107.165 ;
        RECT 104.025 106.575 105.715 106.745 ;
        RECT 102.530 105.975 102.990 106.265 ;
        RECT 103.685 106.235 105.185 106.405 ;
        RECT 103.685 106.095 103.855 106.235 ;
        RECT 103.295 105.925 103.855 106.095 ;
        RECT 101.770 105.295 102.020 105.755 ;
        RECT 102.190 105.465 103.060 105.805 ;
        RECT 103.295 105.465 103.465 105.925 ;
        RECT 104.300 105.895 105.375 106.065 ;
        RECT 103.635 105.295 104.005 105.755 ;
        RECT 104.300 105.555 104.470 105.895 ;
        RECT 104.640 105.295 104.970 105.725 ;
        RECT 105.205 105.555 105.375 105.895 ;
        RECT 105.545 105.795 105.715 106.575 ;
        RECT 105.885 106.355 106.055 106.945 ;
        RECT 106.225 106.545 106.575 107.165 ;
        RECT 105.885 105.965 106.350 106.355 ;
        RECT 106.745 106.095 106.915 107.455 ;
        RECT 107.085 106.265 107.545 107.315 ;
        RECT 106.520 105.925 106.915 106.095 ;
        RECT 106.520 105.795 106.690 105.925 ;
        RECT 105.545 105.465 106.225 105.795 ;
        RECT 106.440 105.465 106.690 105.795 ;
        RECT 106.860 105.295 107.110 105.755 ;
        RECT 107.280 105.480 107.605 106.265 ;
        RECT 107.775 105.465 107.945 107.585 ;
        RECT 108.115 107.465 108.445 107.845 ;
        RECT 108.615 107.295 108.870 107.585 ;
        RECT 108.120 107.125 108.870 107.295 ;
        RECT 109.135 107.295 109.305 107.675 ;
        RECT 109.485 107.465 109.815 107.845 ;
        RECT 109.135 107.125 109.800 107.295 ;
        RECT 109.995 107.170 110.255 107.675 ;
        RECT 108.120 106.135 108.350 107.125 ;
        RECT 108.520 106.305 108.870 106.955 ;
        RECT 109.065 106.575 109.395 106.945 ;
        RECT 109.630 106.870 109.800 107.125 ;
        RECT 109.630 106.540 109.915 106.870 ;
        RECT 109.630 106.395 109.800 106.540 ;
        RECT 109.135 106.225 109.800 106.395 ;
        RECT 110.085 106.370 110.255 107.170 ;
        RECT 110.425 107.095 111.635 107.845 ;
        RECT 108.120 105.965 108.870 106.135 ;
        RECT 108.115 105.295 108.445 105.795 ;
        RECT 108.615 105.465 108.870 105.965 ;
        RECT 109.135 105.465 109.305 106.225 ;
        RECT 109.485 105.295 109.815 106.055 ;
        RECT 109.985 105.465 110.255 106.370 ;
        RECT 110.425 106.385 110.945 106.925 ;
        RECT 111.115 106.555 111.635 107.095 ;
        RECT 111.845 107.025 112.075 107.845 ;
        RECT 112.245 107.045 112.575 107.675 ;
        RECT 111.825 106.605 112.155 106.855 ;
        RECT 112.325 106.445 112.575 107.045 ;
        RECT 112.745 107.025 112.955 107.845 ;
        RECT 113.275 107.295 113.445 107.675 ;
        RECT 113.625 107.465 113.955 107.845 ;
        RECT 113.275 107.125 113.940 107.295 ;
        RECT 114.135 107.170 114.395 107.675 ;
        RECT 113.205 106.575 113.535 106.945 ;
        RECT 113.770 106.870 113.940 107.125 ;
        RECT 110.425 105.295 111.635 106.385 ;
        RECT 111.845 105.295 112.075 106.435 ;
        RECT 112.245 105.465 112.575 106.445 ;
        RECT 113.770 106.540 114.055 106.870 ;
        RECT 112.745 105.295 112.955 106.435 ;
        RECT 113.770 106.395 113.940 106.540 ;
        RECT 113.275 106.225 113.940 106.395 ;
        RECT 114.225 106.370 114.395 107.170 ;
        RECT 114.565 107.120 114.855 107.845 ;
        RECT 115.065 107.025 115.295 107.845 ;
        RECT 115.465 107.045 115.795 107.675 ;
        RECT 115.045 106.605 115.375 106.855 ;
        RECT 113.275 105.465 113.445 106.225 ;
        RECT 113.625 105.295 113.955 106.055 ;
        RECT 114.125 105.465 114.395 106.370 ;
        RECT 114.565 105.295 114.855 106.460 ;
        RECT 115.545 106.445 115.795 107.045 ;
        RECT 115.965 107.025 116.175 107.845 ;
        RECT 117.330 107.295 117.585 107.585 ;
        RECT 117.755 107.465 118.085 107.845 ;
        RECT 117.330 107.125 118.080 107.295 ;
        RECT 115.065 105.295 115.295 106.435 ;
        RECT 115.465 105.465 115.795 106.445 ;
        RECT 115.965 105.295 116.175 106.435 ;
        RECT 117.330 106.305 117.680 106.955 ;
        RECT 117.850 106.135 118.080 107.125 ;
        RECT 117.330 105.965 118.080 106.135 ;
        RECT 117.330 105.465 117.585 105.965 ;
        RECT 117.755 105.295 118.085 105.795 ;
        RECT 118.255 105.465 118.425 107.585 ;
        RECT 118.785 107.485 119.115 107.845 ;
        RECT 119.285 107.455 119.780 107.625 ;
        RECT 119.985 107.455 120.840 107.625 ;
        RECT 118.655 106.265 119.115 107.315 ;
        RECT 118.595 105.480 118.920 106.265 ;
        RECT 119.285 106.095 119.455 107.455 ;
        RECT 119.625 106.545 119.975 107.165 ;
        RECT 120.145 106.945 120.500 107.165 ;
        RECT 120.145 106.355 120.315 106.945 ;
        RECT 120.670 106.745 120.840 107.455 ;
        RECT 121.715 107.385 122.045 107.845 ;
        RECT 122.255 107.485 122.605 107.655 ;
        RECT 121.045 106.915 121.835 107.165 ;
        RECT 122.255 107.095 122.515 107.485 ;
        RECT 122.825 107.395 123.775 107.675 ;
        RECT 123.945 107.405 124.135 107.845 ;
        RECT 124.305 107.465 125.375 107.635 ;
        RECT 122.005 106.745 122.175 106.925 ;
        RECT 119.285 105.925 119.680 106.095 ;
        RECT 119.850 105.965 120.315 106.355 ;
        RECT 120.485 106.575 122.175 106.745 ;
        RECT 119.510 105.795 119.680 105.925 ;
        RECT 120.485 105.795 120.655 106.575 ;
        RECT 122.345 106.405 122.515 107.095 ;
        RECT 121.015 106.235 122.515 106.405 ;
        RECT 122.705 106.435 122.915 107.225 ;
        RECT 123.085 106.605 123.435 107.225 ;
        RECT 123.605 106.615 123.775 107.395 ;
        RECT 124.305 107.235 124.475 107.465 ;
        RECT 123.945 107.065 124.475 107.235 ;
        RECT 123.945 106.785 124.165 107.065 ;
        RECT 124.645 106.895 124.885 107.295 ;
        RECT 123.605 106.445 124.010 106.615 ;
        RECT 124.345 106.525 124.885 106.895 ;
        RECT 125.055 107.110 125.375 107.465 ;
        RECT 125.620 107.385 125.925 107.845 ;
        RECT 126.095 107.135 126.350 107.665 ;
        RECT 125.055 106.935 125.380 107.110 ;
        RECT 125.055 106.635 125.970 106.935 ;
        RECT 125.230 106.605 125.970 106.635 ;
        RECT 122.705 106.275 123.380 106.435 ;
        RECT 123.840 106.355 124.010 106.445 ;
        RECT 122.705 106.265 123.670 106.275 ;
        RECT 122.345 106.095 122.515 106.235 ;
        RECT 119.090 105.295 119.340 105.755 ;
        RECT 119.510 105.465 119.760 105.795 ;
        RECT 119.975 105.465 120.655 105.795 ;
        RECT 120.825 105.895 121.900 106.065 ;
        RECT 122.345 105.925 122.905 106.095 ;
        RECT 123.210 105.975 123.670 106.265 ;
        RECT 123.840 106.185 125.060 106.355 ;
        RECT 120.825 105.555 120.995 105.895 ;
        RECT 121.230 105.295 121.560 105.725 ;
        RECT 121.730 105.555 121.900 105.895 ;
        RECT 122.195 105.295 122.565 105.755 ;
        RECT 122.735 105.465 122.905 105.925 ;
        RECT 123.840 105.805 124.010 106.185 ;
        RECT 125.230 106.015 125.400 106.605 ;
        RECT 126.140 106.485 126.350 107.135 ;
        RECT 126.525 107.095 127.735 107.845 ;
        RECT 123.140 105.465 124.010 105.805 ;
        RECT 124.600 105.845 125.400 106.015 ;
        RECT 124.180 105.295 124.430 105.755 ;
        RECT 124.600 105.555 124.770 105.845 ;
        RECT 124.950 105.295 125.280 105.675 ;
        RECT 125.620 105.295 125.925 106.435 ;
        RECT 126.095 105.605 126.350 106.485 ;
        RECT 126.525 106.385 127.045 106.925 ;
        RECT 127.215 106.555 127.735 107.095 ;
        RECT 126.525 105.295 127.735 106.385 ;
        RECT 14.660 105.125 127.820 105.295 ;
        RECT 14.745 104.035 15.955 105.125 ;
        RECT 14.745 103.325 15.265 103.865 ;
        RECT 15.435 103.495 15.955 104.035 ;
        RECT 16.125 104.035 18.715 105.125 ;
        RECT 18.890 104.690 24.235 105.125 ;
        RECT 16.125 103.515 17.335 104.035 ;
        RECT 17.505 103.345 18.715 103.865 ;
        RECT 20.480 103.440 20.830 104.690 ;
        RECT 24.405 103.960 24.695 105.125 ;
        RECT 14.745 102.575 15.955 103.325 ;
        RECT 16.125 102.575 18.715 103.345 ;
        RECT 22.310 103.120 22.650 103.950 ;
        RECT 24.870 103.935 25.125 104.815 ;
        RECT 25.295 103.985 25.600 105.125 ;
        RECT 25.940 104.745 26.270 105.125 ;
        RECT 26.450 104.575 26.620 104.865 ;
        RECT 26.790 104.665 27.040 105.125 ;
        RECT 25.820 104.405 26.620 104.575 ;
        RECT 27.210 104.615 28.080 104.955 ;
        RECT 18.890 102.575 24.235 103.120 ;
        RECT 24.405 102.575 24.695 103.300 ;
        RECT 24.870 103.285 25.080 103.935 ;
        RECT 25.820 103.815 25.990 104.405 ;
        RECT 27.210 104.235 27.380 104.615 ;
        RECT 28.315 104.495 28.485 104.955 ;
        RECT 28.655 104.665 29.025 105.125 ;
        RECT 29.320 104.525 29.490 104.865 ;
        RECT 29.660 104.695 29.990 105.125 ;
        RECT 30.225 104.525 30.395 104.865 ;
        RECT 26.160 104.065 27.380 104.235 ;
        RECT 27.550 104.155 28.010 104.445 ;
        RECT 28.315 104.325 28.875 104.495 ;
        RECT 29.320 104.355 30.395 104.525 ;
        RECT 30.565 104.625 31.245 104.955 ;
        RECT 31.460 104.625 31.710 104.955 ;
        RECT 31.880 104.665 32.130 105.125 ;
        RECT 28.705 104.185 28.875 104.325 ;
        RECT 27.550 104.145 28.515 104.155 ;
        RECT 27.210 103.975 27.380 104.065 ;
        RECT 27.840 103.985 28.515 104.145 ;
        RECT 25.250 103.785 25.990 103.815 ;
        RECT 25.250 103.485 26.165 103.785 ;
        RECT 25.840 103.310 26.165 103.485 ;
        RECT 24.870 102.755 25.125 103.285 ;
        RECT 25.295 102.575 25.600 103.035 ;
        RECT 25.845 102.955 26.165 103.310 ;
        RECT 26.335 103.525 26.875 103.895 ;
        RECT 27.210 103.805 27.615 103.975 ;
        RECT 26.335 103.125 26.575 103.525 ;
        RECT 27.055 103.355 27.275 103.635 ;
        RECT 26.745 103.185 27.275 103.355 ;
        RECT 26.745 102.955 26.915 103.185 ;
        RECT 27.445 103.025 27.615 103.805 ;
        RECT 27.785 103.195 28.135 103.815 ;
        RECT 28.305 103.195 28.515 103.985 ;
        RECT 28.705 104.015 30.205 104.185 ;
        RECT 28.705 103.325 28.875 104.015 ;
        RECT 30.565 103.845 30.735 104.625 ;
        RECT 31.540 104.495 31.710 104.625 ;
        RECT 29.045 103.675 30.735 103.845 ;
        RECT 30.905 104.065 31.370 104.455 ;
        RECT 31.540 104.325 31.935 104.495 ;
        RECT 29.045 103.495 29.215 103.675 ;
        RECT 25.845 102.785 26.915 102.955 ;
        RECT 27.085 102.575 27.275 103.015 ;
        RECT 27.445 102.745 28.395 103.025 ;
        RECT 28.705 102.935 28.965 103.325 ;
        RECT 29.385 103.255 30.175 103.505 ;
        RECT 28.615 102.765 28.965 102.935 ;
        RECT 29.175 102.575 29.505 103.035 ;
        RECT 30.380 102.965 30.550 103.675 ;
        RECT 30.905 103.475 31.075 104.065 ;
        RECT 30.720 103.255 31.075 103.475 ;
        RECT 31.245 103.255 31.595 103.875 ;
        RECT 31.765 102.965 31.935 104.325 ;
        RECT 32.300 104.155 32.625 104.940 ;
        RECT 32.105 103.105 32.565 104.155 ;
        RECT 30.380 102.795 31.235 102.965 ;
        RECT 31.440 102.795 31.935 102.965 ;
        RECT 32.105 102.575 32.435 102.935 ;
        RECT 32.795 102.835 32.965 104.955 ;
        RECT 33.135 104.625 33.465 105.125 ;
        RECT 33.635 104.455 33.890 104.955 ;
        RECT 33.140 104.285 33.890 104.455 ;
        RECT 33.140 103.295 33.370 104.285 ;
        RECT 33.540 103.465 33.890 104.115 ;
        RECT 34.525 104.035 38.035 105.125 ;
        RECT 34.525 103.515 36.215 104.035 ;
        RECT 38.265 103.985 38.475 105.125 ;
        RECT 38.645 103.975 38.975 104.955 ;
        RECT 39.145 103.985 39.375 105.125 ;
        RECT 39.585 104.035 40.795 105.125 ;
        RECT 40.970 104.455 41.225 104.955 ;
        RECT 41.395 104.625 41.725 105.125 ;
        RECT 40.970 104.285 41.720 104.455 ;
        RECT 36.385 103.345 38.035 103.865 ;
        RECT 33.140 103.125 33.890 103.295 ;
        RECT 33.135 102.575 33.465 102.955 ;
        RECT 33.635 102.835 33.890 103.125 ;
        RECT 34.525 102.575 38.035 103.345 ;
        RECT 38.265 102.575 38.475 103.395 ;
        RECT 38.645 103.375 38.895 103.975 ;
        RECT 39.065 103.565 39.395 103.815 ;
        RECT 39.585 103.495 40.105 104.035 ;
        RECT 38.645 102.745 38.975 103.375 ;
        RECT 39.145 102.575 39.375 103.395 ;
        RECT 40.275 103.325 40.795 103.865 ;
        RECT 40.970 103.465 41.320 104.115 ;
        RECT 39.585 102.575 40.795 103.325 ;
        RECT 41.490 103.295 41.720 104.285 ;
        RECT 40.970 103.125 41.720 103.295 ;
        RECT 40.970 102.835 41.225 103.125 ;
        RECT 41.395 102.575 41.725 102.955 ;
        RECT 41.895 102.835 42.065 104.955 ;
        RECT 42.235 104.155 42.560 104.940 ;
        RECT 42.730 104.665 42.980 105.125 ;
        RECT 43.150 104.625 43.400 104.955 ;
        RECT 43.615 104.625 44.295 104.955 ;
        RECT 43.150 104.495 43.320 104.625 ;
        RECT 42.925 104.325 43.320 104.495 ;
        RECT 42.295 103.105 42.755 104.155 ;
        RECT 42.925 102.965 43.095 104.325 ;
        RECT 43.490 104.065 43.955 104.455 ;
        RECT 43.265 103.255 43.615 103.875 ;
        RECT 43.785 103.475 43.955 104.065 ;
        RECT 44.125 103.845 44.295 104.625 ;
        RECT 44.465 104.525 44.635 104.865 ;
        RECT 44.870 104.695 45.200 105.125 ;
        RECT 45.370 104.525 45.540 104.865 ;
        RECT 45.835 104.665 46.205 105.125 ;
        RECT 44.465 104.355 45.540 104.525 ;
        RECT 46.375 104.495 46.545 104.955 ;
        RECT 46.780 104.615 47.650 104.955 ;
        RECT 47.820 104.665 48.070 105.125 ;
        RECT 45.985 104.325 46.545 104.495 ;
        RECT 45.985 104.185 46.155 104.325 ;
        RECT 44.655 104.015 46.155 104.185 ;
        RECT 46.850 104.155 47.310 104.445 ;
        RECT 44.125 103.675 45.815 103.845 ;
        RECT 43.785 103.255 44.140 103.475 ;
        RECT 44.310 102.965 44.480 103.675 ;
        RECT 44.685 103.255 45.475 103.505 ;
        RECT 45.645 103.495 45.815 103.675 ;
        RECT 45.985 103.325 46.155 104.015 ;
        RECT 42.425 102.575 42.755 102.935 ;
        RECT 42.925 102.795 43.420 102.965 ;
        RECT 43.625 102.795 44.480 102.965 ;
        RECT 45.355 102.575 45.685 103.035 ;
        RECT 45.895 102.935 46.155 103.325 ;
        RECT 46.345 104.145 47.310 104.155 ;
        RECT 47.480 104.235 47.650 104.615 ;
        RECT 48.240 104.575 48.410 104.865 ;
        RECT 48.590 104.745 48.920 105.125 ;
        RECT 48.240 104.405 49.040 104.575 ;
        RECT 46.345 103.985 47.020 104.145 ;
        RECT 47.480 104.065 48.700 104.235 ;
        RECT 46.345 103.195 46.555 103.985 ;
        RECT 47.480 103.975 47.650 104.065 ;
        RECT 46.725 103.195 47.075 103.815 ;
        RECT 47.245 103.805 47.650 103.975 ;
        RECT 47.245 103.025 47.415 103.805 ;
        RECT 47.585 103.355 47.805 103.635 ;
        RECT 47.985 103.525 48.525 103.895 ;
        RECT 48.870 103.815 49.040 104.405 ;
        RECT 49.260 103.985 49.565 105.125 ;
        RECT 49.735 103.935 49.990 104.815 ;
        RECT 50.165 103.960 50.455 105.125 ;
        RECT 51.090 104.455 51.345 104.955 ;
        RECT 51.515 104.625 51.845 105.125 ;
        RECT 51.090 104.285 51.840 104.455 ;
        RECT 48.870 103.785 49.610 103.815 ;
        RECT 47.585 103.185 48.115 103.355 ;
        RECT 45.895 102.765 46.245 102.935 ;
        RECT 46.465 102.745 47.415 103.025 ;
        RECT 47.585 102.575 47.775 103.015 ;
        RECT 47.945 102.955 48.115 103.185 ;
        RECT 48.285 103.125 48.525 103.525 ;
        RECT 48.695 103.485 49.610 103.785 ;
        RECT 48.695 103.310 49.020 103.485 ;
        RECT 48.695 102.955 49.015 103.310 ;
        RECT 49.780 103.285 49.990 103.935 ;
        RECT 51.090 103.465 51.440 104.115 ;
        RECT 47.945 102.785 49.015 102.955 ;
        RECT 49.260 102.575 49.565 103.035 ;
        RECT 49.735 102.755 49.990 103.285 ;
        RECT 50.165 102.575 50.455 103.300 ;
        RECT 51.610 103.295 51.840 104.285 ;
        RECT 51.090 103.125 51.840 103.295 ;
        RECT 51.090 102.835 51.345 103.125 ;
        RECT 51.515 102.575 51.845 102.955 ;
        RECT 52.015 102.835 52.185 104.955 ;
        RECT 52.355 104.155 52.680 104.940 ;
        RECT 52.850 104.665 53.100 105.125 ;
        RECT 53.270 104.625 53.520 104.955 ;
        RECT 53.735 104.625 54.415 104.955 ;
        RECT 53.270 104.495 53.440 104.625 ;
        RECT 53.045 104.325 53.440 104.495 ;
        RECT 52.415 103.105 52.875 104.155 ;
        RECT 53.045 102.965 53.215 104.325 ;
        RECT 53.610 104.065 54.075 104.455 ;
        RECT 53.385 103.255 53.735 103.875 ;
        RECT 53.905 103.475 54.075 104.065 ;
        RECT 54.245 103.845 54.415 104.625 ;
        RECT 54.585 104.525 54.755 104.865 ;
        RECT 54.990 104.695 55.320 105.125 ;
        RECT 55.490 104.525 55.660 104.865 ;
        RECT 55.955 104.665 56.325 105.125 ;
        RECT 54.585 104.355 55.660 104.525 ;
        RECT 56.495 104.495 56.665 104.955 ;
        RECT 56.900 104.615 57.770 104.955 ;
        RECT 57.940 104.665 58.190 105.125 ;
        RECT 56.105 104.325 56.665 104.495 ;
        RECT 56.105 104.185 56.275 104.325 ;
        RECT 54.775 104.015 56.275 104.185 ;
        RECT 56.970 104.155 57.430 104.445 ;
        RECT 54.245 103.675 55.935 103.845 ;
        RECT 53.905 103.255 54.260 103.475 ;
        RECT 54.430 102.965 54.600 103.675 ;
        RECT 54.805 103.255 55.595 103.505 ;
        RECT 55.765 103.495 55.935 103.675 ;
        RECT 56.105 103.325 56.275 104.015 ;
        RECT 52.545 102.575 52.875 102.935 ;
        RECT 53.045 102.795 53.540 102.965 ;
        RECT 53.745 102.795 54.600 102.965 ;
        RECT 55.475 102.575 55.805 103.035 ;
        RECT 56.015 102.935 56.275 103.325 ;
        RECT 56.465 104.145 57.430 104.155 ;
        RECT 57.600 104.235 57.770 104.615 ;
        RECT 58.360 104.575 58.530 104.865 ;
        RECT 58.710 104.745 59.040 105.125 ;
        RECT 58.360 104.405 59.160 104.575 ;
        RECT 56.465 103.985 57.140 104.145 ;
        RECT 57.600 104.065 58.820 104.235 ;
        RECT 56.465 103.195 56.675 103.985 ;
        RECT 57.600 103.975 57.770 104.065 ;
        RECT 56.845 103.195 57.195 103.815 ;
        RECT 57.365 103.805 57.770 103.975 ;
        RECT 57.365 103.025 57.535 103.805 ;
        RECT 57.705 103.355 57.925 103.635 ;
        RECT 58.105 103.525 58.645 103.895 ;
        RECT 58.990 103.815 59.160 104.405 ;
        RECT 59.380 103.985 59.685 105.125 ;
        RECT 59.855 103.935 60.110 104.815 ;
        RECT 58.990 103.785 59.730 103.815 ;
        RECT 57.705 103.185 58.235 103.355 ;
        RECT 56.015 102.765 56.365 102.935 ;
        RECT 56.585 102.745 57.535 103.025 ;
        RECT 57.705 102.575 57.895 103.015 ;
        RECT 58.065 102.955 58.235 103.185 ;
        RECT 58.405 103.125 58.645 103.525 ;
        RECT 58.815 103.485 59.730 103.785 ;
        RECT 58.815 103.310 59.140 103.485 ;
        RECT 58.815 102.955 59.135 103.310 ;
        RECT 59.900 103.285 60.110 103.935 ;
        RECT 58.065 102.785 59.135 102.955 ;
        RECT 59.380 102.575 59.685 103.035 ;
        RECT 59.855 102.755 60.110 103.285 ;
        RECT 60.290 103.935 60.545 104.815 ;
        RECT 60.715 103.985 61.020 105.125 ;
        RECT 61.360 104.745 61.690 105.125 ;
        RECT 61.870 104.575 62.040 104.865 ;
        RECT 62.210 104.665 62.460 105.125 ;
        RECT 61.240 104.405 62.040 104.575 ;
        RECT 62.630 104.615 63.500 104.955 ;
        RECT 60.290 103.285 60.500 103.935 ;
        RECT 61.240 103.815 61.410 104.405 ;
        RECT 62.630 104.235 62.800 104.615 ;
        RECT 63.735 104.495 63.905 104.955 ;
        RECT 64.075 104.665 64.445 105.125 ;
        RECT 64.740 104.525 64.910 104.865 ;
        RECT 65.080 104.695 65.410 105.125 ;
        RECT 65.645 104.525 65.815 104.865 ;
        RECT 61.580 104.065 62.800 104.235 ;
        RECT 62.970 104.155 63.430 104.445 ;
        RECT 63.735 104.325 64.295 104.495 ;
        RECT 64.740 104.355 65.815 104.525 ;
        RECT 65.985 104.625 66.665 104.955 ;
        RECT 66.880 104.625 67.130 104.955 ;
        RECT 67.300 104.665 67.550 105.125 ;
        RECT 64.125 104.185 64.295 104.325 ;
        RECT 62.970 104.145 63.935 104.155 ;
        RECT 62.630 103.975 62.800 104.065 ;
        RECT 63.260 103.985 63.935 104.145 ;
        RECT 60.670 103.785 61.410 103.815 ;
        RECT 60.670 103.485 61.585 103.785 ;
        RECT 61.260 103.310 61.585 103.485 ;
        RECT 60.290 102.755 60.545 103.285 ;
        RECT 60.715 102.575 61.020 103.035 ;
        RECT 61.265 102.955 61.585 103.310 ;
        RECT 61.755 103.525 62.295 103.895 ;
        RECT 62.630 103.805 63.035 103.975 ;
        RECT 61.755 103.125 61.995 103.525 ;
        RECT 62.475 103.355 62.695 103.635 ;
        RECT 62.165 103.185 62.695 103.355 ;
        RECT 62.165 102.955 62.335 103.185 ;
        RECT 62.865 103.025 63.035 103.805 ;
        RECT 63.205 103.195 63.555 103.815 ;
        RECT 63.725 103.195 63.935 103.985 ;
        RECT 64.125 104.015 65.625 104.185 ;
        RECT 64.125 103.325 64.295 104.015 ;
        RECT 65.985 103.845 66.155 104.625 ;
        RECT 66.960 104.495 67.130 104.625 ;
        RECT 64.465 103.675 66.155 103.845 ;
        RECT 66.325 104.065 66.790 104.455 ;
        RECT 66.960 104.325 67.355 104.495 ;
        RECT 64.465 103.495 64.635 103.675 ;
        RECT 61.265 102.785 62.335 102.955 ;
        RECT 62.505 102.575 62.695 103.015 ;
        RECT 62.865 102.745 63.815 103.025 ;
        RECT 64.125 102.935 64.385 103.325 ;
        RECT 64.805 103.255 65.595 103.505 ;
        RECT 64.035 102.765 64.385 102.935 ;
        RECT 64.595 102.575 64.925 103.035 ;
        RECT 65.800 102.965 65.970 103.675 ;
        RECT 66.325 103.475 66.495 104.065 ;
        RECT 66.140 103.255 66.495 103.475 ;
        RECT 66.665 103.255 67.015 103.875 ;
        RECT 67.185 102.965 67.355 104.325 ;
        RECT 67.720 104.155 68.045 104.940 ;
        RECT 67.525 103.105 67.985 104.155 ;
        RECT 65.800 102.795 66.655 102.965 ;
        RECT 66.860 102.795 67.355 102.965 ;
        RECT 67.525 102.575 67.855 102.935 ;
        RECT 68.215 102.835 68.385 104.955 ;
        RECT 68.555 104.625 68.885 105.125 ;
        RECT 69.055 104.455 69.310 104.955 ;
        RECT 70.410 104.690 75.755 105.125 ;
        RECT 68.560 104.285 69.310 104.455 ;
        RECT 68.560 103.295 68.790 104.285 ;
        RECT 68.960 103.465 69.310 104.115 ;
        RECT 72.000 103.440 72.350 104.690 ;
        RECT 75.925 103.960 76.215 105.125 ;
        RECT 68.560 103.125 69.310 103.295 ;
        RECT 68.555 102.575 68.885 102.955 ;
        RECT 69.055 102.835 69.310 103.125 ;
        RECT 73.830 103.120 74.170 103.950 ;
        RECT 76.390 103.935 76.645 104.815 ;
        RECT 76.815 103.985 77.120 105.125 ;
        RECT 77.460 104.745 77.790 105.125 ;
        RECT 77.970 104.575 78.140 104.865 ;
        RECT 78.310 104.665 78.560 105.125 ;
        RECT 77.340 104.405 78.140 104.575 ;
        RECT 78.730 104.615 79.600 104.955 ;
        RECT 70.410 102.575 75.755 103.120 ;
        RECT 75.925 102.575 76.215 103.300 ;
        RECT 76.390 103.285 76.600 103.935 ;
        RECT 77.340 103.815 77.510 104.405 ;
        RECT 78.730 104.235 78.900 104.615 ;
        RECT 79.835 104.495 80.005 104.955 ;
        RECT 80.175 104.665 80.545 105.125 ;
        RECT 80.840 104.525 81.010 104.865 ;
        RECT 81.180 104.695 81.510 105.125 ;
        RECT 81.745 104.525 81.915 104.865 ;
        RECT 77.680 104.065 78.900 104.235 ;
        RECT 79.070 104.155 79.530 104.445 ;
        RECT 79.835 104.325 80.395 104.495 ;
        RECT 80.840 104.355 81.915 104.525 ;
        RECT 82.085 104.625 82.765 104.955 ;
        RECT 82.980 104.625 83.230 104.955 ;
        RECT 83.400 104.665 83.650 105.125 ;
        RECT 80.225 104.185 80.395 104.325 ;
        RECT 79.070 104.145 80.035 104.155 ;
        RECT 78.730 103.975 78.900 104.065 ;
        RECT 79.360 103.985 80.035 104.145 ;
        RECT 76.770 103.785 77.510 103.815 ;
        RECT 76.770 103.485 77.685 103.785 ;
        RECT 77.360 103.310 77.685 103.485 ;
        RECT 76.390 102.755 76.645 103.285 ;
        RECT 76.815 102.575 77.120 103.035 ;
        RECT 77.365 102.955 77.685 103.310 ;
        RECT 77.855 103.525 78.395 103.895 ;
        RECT 78.730 103.805 79.135 103.975 ;
        RECT 77.855 103.125 78.095 103.525 ;
        RECT 78.575 103.355 78.795 103.635 ;
        RECT 78.265 103.185 78.795 103.355 ;
        RECT 78.265 102.955 78.435 103.185 ;
        RECT 78.965 103.025 79.135 103.805 ;
        RECT 79.305 103.195 79.655 103.815 ;
        RECT 79.825 103.195 80.035 103.985 ;
        RECT 80.225 104.015 81.725 104.185 ;
        RECT 80.225 103.325 80.395 104.015 ;
        RECT 82.085 103.845 82.255 104.625 ;
        RECT 83.060 104.495 83.230 104.625 ;
        RECT 80.565 103.675 82.255 103.845 ;
        RECT 82.425 104.065 82.890 104.455 ;
        RECT 83.060 104.325 83.455 104.495 ;
        RECT 80.565 103.495 80.735 103.675 ;
        RECT 77.365 102.785 78.435 102.955 ;
        RECT 78.605 102.575 78.795 103.015 ;
        RECT 78.965 102.745 79.915 103.025 ;
        RECT 80.225 102.935 80.485 103.325 ;
        RECT 80.905 103.255 81.695 103.505 ;
        RECT 80.135 102.765 80.485 102.935 ;
        RECT 80.695 102.575 81.025 103.035 ;
        RECT 81.900 102.965 82.070 103.675 ;
        RECT 82.425 103.475 82.595 104.065 ;
        RECT 82.240 103.255 82.595 103.475 ;
        RECT 82.765 103.255 83.115 103.875 ;
        RECT 83.285 102.965 83.455 104.325 ;
        RECT 83.820 104.155 84.145 104.940 ;
        RECT 83.625 103.105 84.085 104.155 ;
        RECT 81.900 102.795 82.755 102.965 ;
        RECT 82.960 102.795 83.455 102.965 ;
        RECT 83.625 102.575 83.955 102.935 ;
        RECT 84.315 102.835 84.485 104.955 ;
        RECT 84.655 104.625 84.985 105.125 ;
        RECT 85.155 104.455 85.410 104.955 ;
        RECT 84.660 104.285 85.410 104.455 ;
        RECT 84.660 103.295 84.890 104.285 ;
        RECT 85.060 103.465 85.410 104.115 ;
        RECT 85.590 103.935 85.845 104.815 ;
        RECT 86.015 103.985 86.320 105.125 ;
        RECT 86.660 104.745 86.990 105.125 ;
        RECT 87.170 104.575 87.340 104.865 ;
        RECT 87.510 104.665 87.760 105.125 ;
        RECT 86.540 104.405 87.340 104.575 ;
        RECT 87.930 104.615 88.800 104.955 ;
        RECT 84.660 103.125 85.410 103.295 ;
        RECT 84.655 102.575 84.985 102.955 ;
        RECT 85.155 102.835 85.410 103.125 ;
        RECT 85.590 103.285 85.800 103.935 ;
        RECT 86.540 103.815 86.710 104.405 ;
        RECT 87.930 104.235 88.100 104.615 ;
        RECT 89.035 104.495 89.205 104.955 ;
        RECT 89.375 104.665 89.745 105.125 ;
        RECT 90.040 104.525 90.210 104.865 ;
        RECT 90.380 104.695 90.710 105.125 ;
        RECT 90.945 104.525 91.115 104.865 ;
        RECT 86.880 104.065 88.100 104.235 ;
        RECT 88.270 104.155 88.730 104.445 ;
        RECT 89.035 104.325 89.595 104.495 ;
        RECT 90.040 104.355 91.115 104.525 ;
        RECT 91.285 104.625 91.965 104.955 ;
        RECT 92.180 104.625 92.430 104.955 ;
        RECT 92.600 104.665 92.850 105.125 ;
        RECT 89.425 104.185 89.595 104.325 ;
        RECT 88.270 104.145 89.235 104.155 ;
        RECT 87.930 103.975 88.100 104.065 ;
        RECT 88.560 103.985 89.235 104.145 ;
        RECT 85.970 103.785 86.710 103.815 ;
        RECT 85.970 103.485 86.885 103.785 ;
        RECT 86.560 103.310 86.885 103.485 ;
        RECT 85.590 102.755 85.845 103.285 ;
        RECT 86.015 102.575 86.320 103.035 ;
        RECT 86.565 102.955 86.885 103.310 ;
        RECT 87.055 103.525 87.595 103.895 ;
        RECT 87.930 103.805 88.335 103.975 ;
        RECT 87.055 103.125 87.295 103.525 ;
        RECT 87.775 103.355 87.995 103.635 ;
        RECT 87.465 103.185 87.995 103.355 ;
        RECT 87.465 102.955 87.635 103.185 ;
        RECT 88.165 103.025 88.335 103.805 ;
        RECT 88.505 103.195 88.855 103.815 ;
        RECT 89.025 103.195 89.235 103.985 ;
        RECT 89.425 104.015 90.925 104.185 ;
        RECT 89.425 103.325 89.595 104.015 ;
        RECT 91.285 103.845 91.455 104.625 ;
        RECT 92.260 104.495 92.430 104.625 ;
        RECT 89.765 103.675 91.455 103.845 ;
        RECT 91.625 104.065 92.090 104.455 ;
        RECT 92.260 104.325 92.655 104.495 ;
        RECT 89.765 103.495 89.935 103.675 ;
        RECT 86.565 102.785 87.635 102.955 ;
        RECT 87.805 102.575 87.995 103.015 ;
        RECT 88.165 102.745 89.115 103.025 ;
        RECT 89.425 102.935 89.685 103.325 ;
        RECT 90.105 103.255 90.895 103.505 ;
        RECT 89.335 102.765 89.685 102.935 ;
        RECT 89.895 102.575 90.225 103.035 ;
        RECT 91.100 102.965 91.270 103.675 ;
        RECT 91.625 103.475 91.795 104.065 ;
        RECT 91.440 103.255 91.795 103.475 ;
        RECT 91.965 103.255 92.315 103.875 ;
        RECT 92.485 102.965 92.655 104.325 ;
        RECT 93.020 104.155 93.345 104.940 ;
        RECT 92.825 103.105 93.285 104.155 ;
        RECT 91.100 102.795 91.955 102.965 ;
        RECT 92.160 102.795 92.655 102.965 ;
        RECT 92.825 102.575 93.155 102.935 ;
        RECT 93.515 102.835 93.685 104.955 ;
        RECT 93.855 104.625 94.185 105.125 ;
        RECT 94.355 104.455 94.610 104.955 ;
        RECT 93.860 104.285 94.610 104.455 ;
        RECT 93.860 103.295 94.090 104.285 ;
        RECT 94.260 103.465 94.610 104.115 ;
        RECT 94.785 104.035 95.995 105.125 ;
        RECT 96.170 104.690 101.515 105.125 ;
        RECT 94.785 103.495 95.305 104.035 ;
        RECT 95.475 103.325 95.995 103.865 ;
        RECT 97.760 103.440 98.110 104.690 ;
        RECT 101.685 103.960 101.975 105.125 ;
        RECT 102.605 104.035 104.275 105.125 ;
        RECT 93.860 103.125 94.610 103.295 ;
        RECT 93.855 102.575 94.185 102.955 ;
        RECT 94.355 102.835 94.610 103.125 ;
        RECT 94.785 102.575 95.995 103.325 ;
        RECT 99.590 103.120 99.930 103.950 ;
        RECT 102.605 103.515 103.355 104.035 ;
        RECT 104.450 103.935 104.705 104.815 ;
        RECT 104.875 103.985 105.180 105.125 ;
        RECT 105.520 104.745 105.850 105.125 ;
        RECT 106.030 104.575 106.200 104.865 ;
        RECT 106.370 104.665 106.620 105.125 ;
        RECT 105.400 104.405 106.200 104.575 ;
        RECT 106.790 104.615 107.660 104.955 ;
        RECT 103.525 103.345 104.275 103.865 ;
        RECT 96.170 102.575 101.515 103.120 ;
        RECT 101.685 102.575 101.975 103.300 ;
        RECT 102.605 102.575 104.275 103.345 ;
        RECT 104.450 103.285 104.660 103.935 ;
        RECT 105.400 103.815 105.570 104.405 ;
        RECT 106.790 104.235 106.960 104.615 ;
        RECT 107.895 104.495 108.065 104.955 ;
        RECT 108.235 104.665 108.605 105.125 ;
        RECT 108.900 104.525 109.070 104.865 ;
        RECT 109.240 104.695 109.570 105.125 ;
        RECT 109.805 104.525 109.975 104.865 ;
        RECT 105.740 104.065 106.960 104.235 ;
        RECT 107.130 104.155 107.590 104.445 ;
        RECT 107.895 104.325 108.455 104.495 ;
        RECT 108.900 104.355 109.975 104.525 ;
        RECT 110.145 104.625 110.825 104.955 ;
        RECT 111.040 104.625 111.290 104.955 ;
        RECT 111.460 104.665 111.710 105.125 ;
        RECT 108.285 104.185 108.455 104.325 ;
        RECT 107.130 104.145 108.095 104.155 ;
        RECT 106.790 103.975 106.960 104.065 ;
        RECT 107.420 103.985 108.095 104.145 ;
        RECT 104.830 103.785 105.570 103.815 ;
        RECT 104.830 103.485 105.745 103.785 ;
        RECT 105.420 103.310 105.745 103.485 ;
        RECT 104.450 102.755 104.705 103.285 ;
        RECT 104.875 102.575 105.180 103.035 ;
        RECT 105.425 102.955 105.745 103.310 ;
        RECT 105.915 103.525 106.455 103.895 ;
        RECT 106.790 103.805 107.195 103.975 ;
        RECT 105.915 103.125 106.155 103.525 ;
        RECT 106.635 103.355 106.855 103.635 ;
        RECT 106.325 103.185 106.855 103.355 ;
        RECT 106.325 102.955 106.495 103.185 ;
        RECT 107.025 103.025 107.195 103.805 ;
        RECT 107.365 103.195 107.715 103.815 ;
        RECT 107.885 103.195 108.095 103.985 ;
        RECT 108.285 104.015 109.785 104.185 ;
        RECT 108.285 103.325 108.455 104.015 ;
        RECT 110.145 103.845 110.315 104.625 ;
        RECT 111.120 104.495 111.290 104.625 ;
        RECT 108.625 103.675 110.315 103.845 ;
        RECT 110.485 104.065 110.950 104.455 ;
        RECT 111.120 104.325 111.515 104.495 ;
        RECT 108.625 103.495 108.795 103.675 ;
        RECT 105.425 102.785 106.495 102.955 ;
        RECT 106.665 102.575 106.855 103.015 ;
        RECT 107.025 102.745 107.975 103.025 ;
        RECT 108.285 102.935 108.545 103.325 ;
        RECT 108.965 103.255 109.755 103.505 ;
        RECT 108.195 102.765 108.545 102.935 ;
        RECT 108.755 102.575 109.085 103.035 ;
        RECT 109.960 102.965 110.130 103.675 ;
        RECT 110.485 103.475 110.655 104.065 ;
        RECT 110.300 103.255 110.655 103.475 ;
        RECT 110.825 103.255 111.175 103.875 ;
        RECT 111.345 102.965 111.515 104.325 ;
        RECT 111.880 104.155 112.205 104.940 ;
        RECT 111.685 103.105 112.145 104.155 ;
        RECT 109.960 102.795 110.815 102.965 ;
        RECT 111.020 102.795 111.515 102.965 ;
        RECT 111.685 102.575 112.015 102.935 ;
        RECT 112.375 102.835 112.545 104.955 ;
        RECT 112.715 104.625 113.045 105.125 ;
        RECT 113.215 104.455 113.470 104.955 ;
        RECT 112.720 104.285 113.470 104.455 ;
        RECT 112.720 103.295 112.950 104.285 ;
        RECT 113.120 103.465 113.470 104.115 ;
        RECT 113.650 103.935 113.905 104.815 ;
        RECT 114.075 103.985 114.380 105.125 ;
        RECT 114.720 104.745 115.050 105.125 ;
        RECT 115.230 104.575 115.400 104.865 ;
        RECT 115.570 104.665 115.820 105.125 ;
        RECT 114.600 104.405 115.400 104.575 ;
        RECT 115.990 104.615 116.860 104.955 ;
        RECT 112.720 103.125 113.470 103.295 ;
        RECT 112.715 102.575 113.045 102.955 ;
        RECT 113.215 102.835 113.470 103.125 ;
        RECT 113.650 103.285 113.860 103.935 ;
        RECT 114.600 103.815 114.770 104.405 ;
        RECT 115.990 104.235 116.160 104.615 ;
        RECT 117.095 104.495 117.265 104.955 ;
        RECT 117.435 104.665 117.805 105.125 ;
        RECT 118.100 104.525 118.270 104.865 ;
        RECT 118.440 104.695 118.770 105.125 ;
        RECT 119.005 104.525 119.175 104.865 ;
        RECT 114.940 104.065 116.160 104.235 ;
        RECT 116.330 104.155 116.790 104.445 ;
        RECT 117.095 104.325 117.655 104.495 ;
        RECT 118.100 104.355 119.175 104.525 ;
        RECT 119.345 104.625 120.025 104.955 ;
        RECT 120.240 104.625 120.490 104.955 ;
        RECT 120.660 104.665 120.910 105.125 ;
        RECT 117.485 104.185 117.655 104.325 ;
        RECT 116.330 104.145 117.295 104.155 ;
        RECT 115.990 103.975 116.160 104.065 ;
        RECT 116.620 103.985 117.295 104.145 ;
        RECT 114.030 103.785 114.770 103.815 ;
        RECT 114.030 103.485 114.945 103.785 ;
        RECT 114.620 103.310 114.945 103.485 ;
        RECT 113.650 102.755 113.905 103.285 ;
        RECT 114.075 102.575 114.380 103.035 ;
        RECT 114.625 102.955 114.945 103.310 ;
        RECT 115.115 103.525 115.655 103.895 ;
        RECT 115.990 103.805 116.395 103.975 ;
        RECT 115.115 103.125 115.355 103.525 ;
        RECT 115.835 103.355 116.055 103.635 ;
        RECT 115.525 103.185 116.055 103.355 ;
        RECT 115.525 102.955 115.695 103.185 ;
        RECT 116.225 103.025 116.395 103.805 ;
        RECT 116.565 103.195 116.915 103.815 ;
        RECT 117.085 103.195 117.295 103.985 ;
        RECT 117.485 104.015 118.985 104.185 ;
        RECT 117.485 103.325 117.655 104.015 ;
        RECT 119.345 103.845 119.515 104.625 ;
        RECT 120.320 104.495 120.490 104.625 ;
        RECT 117.825 103.675 119.515 103.845 ;
        RECT 119.685 104.065 120.150 104.455 ;
        RECT 120.320 104.325 120.715 104.495 ;
        RECT 117.825 103.495 117.995 103.675 ;
        RECT 114.625 102.785 115.695 102.955 ;
        RECT 115.865 102.575 116.055 103.015 ;
        RECT 116.225 102.745 117.175 103.025 ;
        RECT 117.485 102.935 117.745 103.325 ;
        RECT 118.165 103.255 118.955 103.505 ;
        RECT 117.395 102.765 117.745 102.935 ;
        RECT 117.955 102.575 118.285 103.035 ;
        RECT 119.160 102.965 119.330 103.675 ;
        RECT 119.685 103.475 119.855 104.065 ;
        RECT 119.500 103.255 119.855 103.475 ;
        RECT 120.025 103.255 120.375 103.875 ;
        RECT 120.545 102.965 120.715 104.325 ;
        RECT 121.080 104.155 121.405 104.940 ;
        RECT 120.885 103.105 121.345 104.155 ;
        RECT 119.160 102.795 120.015 102.965 ;
        RECT 120.220 102.795 120.715 102.965 ;
        RECT 120.885 102.575 121.215 102.935 ;
        RECT 121.575 102.835 121.745 104.955 ;
        RECT 121.915 104.625 122.245 105.125 ;
        RECT 122.415 104.455 122.670 104.955 ;
        RECT 121.920 104.285 122.670 104.455 ;
        RECT 121.920 103.295 122.150 104.285 ;
        RECT 122.320 103.465 122.670 104.115 ;
        RECT 123.305 104.035 124.975 105.125 ;
        RECT 125.145 104.050 125.415 104.955 ;
        RECT 125.585 104.365 125.915 105.125 ;
        RECT 126.095 104.195 126.275 104.955 ;
        RECT 123.305 103.515 124.055 104.035 ;
        RECT 124.225 103.345 124.975 103.865 ;
        RECT 121.920 103.125 122.670 103.295 ;
        RECT 121.915 102.575 122.245 102.955 ;
        RECT 122.415 102.835 122.670 103.125 ;
        RECT 123.305 102.575 124.975 103.345 ;
        RECT 125.145 103.250 125.325 104.050 ;
        RECT 125.600 104.025 126.275 104.195 ;
        RECT 126.525 104.035 127.735 105.125 ;
        RECT 125.600 103.880 125.770 104.025 ;
        RECT 125.495 103.550 125.770 103.880 ;
        RECT 125.600 103.295 125.770 103.550 ;
        RECT 125.995 103.475 126.335 103.845 ;
        RECT 126.525 103.495 127.045 104.035 ;
        RECT 127.215 103.325 127.735 103.865 ;
        RECT 125.145 102.745 125.405 103.250 ;
        RECT 125.600 103.125 126.265 103.295 ;
        RECT 125.585 102.575 125.915 102.955 ;
        RECT 126.095 102.745 126.265 103.125 ;
        RECT 126.525 102.575 127.735 103.325 ;
        RECT 14.660 102.405 127.820 102.575 ;
        RECT 14.745 101.655 15.955 102.405 ;
        RECT 14.745 101.115 15.265 101.655 ;
        RECT 16.125 101.635 18.715 102.405 ;
        RECT 18.890 101.860 24.235 102.405 ;
        RECT 15.435 100.945 15.955 101.485 ;
        RECT 14.745 99.855 15.955 100.945 ;
        RECT 16.125 100.945 17.335 101.465 ;
        RECT 17.505 101.115 18.715 101.635 ;
        RECT 16.125 99.855 18.715 100.945 ;
        RECT 20.480 100.290 20.830 101.540 ;
        RECT 22.310 101.030 22.650 101.860 ;
        RECT 24.405 101.680 24.695 102.405 ;
        RECT 24.865 101.655 26.075 102.405 ;
        RECT 26.250 101.860 31.595 102.405 ;
        RECT 31.770 101.860 37.115 102.405 ;
        RECT 18.890 99.855 24.235 100.290 ;
        RECT 24.405 99.855 24.695 101.020 ;
        RECT 24.865 100.945 25.385 101.485 ;
        RECT 25.555 101.115 26.075 101.655 ;
        RECT 24.865 99.855 26.075 100.945 ;
        RECT 27.840 100.290 28.190 101.540 ;
        RECT 29.670 101.030 30.010 101.860 ;
        RECT 33.360 100.290 33.710 101.540 ;
        RECT 35.190 101.030 35.530 101.860 ;
        RECT 37.285 101.680 37.575 102.405 ;
        RECT 37.745 101.635 41.255 102.405 ;
        RECT 41.430 101.860 46.775 102.405 ;
        RECT 26.250 99.855 31.595 100.290 ;
        RECT 31.770 99.855 37.115 100.290 ;
        RECT 37.285 99.855 37.575 101.020 ;
        RECT 37.745 100.945 39.435 101.465 ;
        RECT 39.605 101.115 41.255 101.635 ;
        RECT 37.745 99.855 41.255 100.945 ;
        RECT 43.020 100.290 43.370 101.540 ;
        RECT 44.850 101.030 45.190 101.860 ;
        RECT 47.005 101.585 47.215 102.405 ;
        RECT 47.385 101.605 47.715 102.235 ;
        RECT 47.385 101.005 47.635 101.605 ;
        RECT 47.885 101.585 48.115 102.405 ;
        RECT 48.325 101.635 49.995 102.405 ;
        RECT 50.165 101.680 50.455 102.405 ;
        RECT 50.625 101.655 51.835 102.405 ;
        RECT 52.010 101.860 57.355 102.405 ;
        RECT 57.530 101.860 62.875 102.405 ;
        RECT 47.805 101.165 48.135 101.415 ;
        RECT 41.430 99.855 46.775 100.290 ;
        RECT 47.005 99.855 47.215 100.995 ;
        RECT 47.385 100.025 47.715 101.005 ;
        RECT 47.885 99.855 48.115 100.995 ;
        RECT 48.325 100.945 49.075 101.465 ;
        RECT 49.245 101.115 49.995 101.635 ;
        RECT 48.325 99.855 49.995 100.945 ;
        RECT 50.165 99.855 50.455 101.020 ;
        RECT 50.625 100.945 51.145 101.485 ;
        RECT 51.315 101.115 51.835 101.655 ;
        RECT 50.625 99.855 51.835 100.945 ;
        RECT 53.600 100.290 53.950 101.540 ;
        RECT 55.430 101.030 55.770 101.860 ;
        RECT 59.120 100.290 59.470 101.540 ;
        RECT 60.950 101.030 61.290 101.860 ;
        RECT 63.045 101.680 63.335 102.405 ;
        RECT 64.465 101.585 64.695 102.405 ;
        RECT 64.865 101.605 65.195 102.235 ;
        RECT 64.445 101.165 64.775 101.415 ;
        RECT 52.010 99.855 57.355 100.290 ;
        RECT 57.530 99.855 62.875 100.290 ;
        RECT 63.045 99.855 63.335 101.020 ;
        RECT 64.945 101.005 65.195 101.605 ;
        RECT 65.365 101.585 65.575 102.405 ;
        RECT 66.725 101.635 70.235 102.405 ;
        RECT 70.410 101.860 75.755 102.405 ;
        RECT 64.465 99.855 64.695 100.995 ;
        RECT 64.865 100.025 65.195 101.005 ;
        RECT 65.365 99.855 65.575 100.995 ;
        RECT 66.725 100.945 68.415 101.465 ;
        RECT 68.585 101.115 70.235 101.635 ;
        RECT 66.725 99.855 70.235 100.945 ;
        RECT 72.000 100.290 72.350 101.540 ;
        RECT 73.830 101.030 74.170 101.860 ;
        RECT 75.925 101.680 76.215 102.405 ;
        RECT 76.385 101.655 77.595 102.405 ;
        RECT 77.770 101.860 83.115 102.405 ;
        RECT 83.290 101.860 88.635 102.405 ;
        RECT 70.410 99.855 75.755 100.290 ;
        RECT 75.925 99.855 76.215 101.020 ;
        RECT 76.385 100.945 76.905 101.485 ;
        RECT 77.075 101.115 77.595 101.655 ;
        RECT 76.385 99.855 77.595 100.945 ;
        RECT 79.360 100.290 79.710 101.540 ;
        RECT 81.190 101.030 81.530 101.860 ;
        RECT 84.880 100.290 85.230 101.540 ;
        RECT 86.710 101.030 87.050 101.860 ;
        RECT 88.805 101.680 89.095 102.405 ;
        RECT 89.265 101.655 90.475 102.405 ;
        RECT 90.650 101.860 95.995 102.405 ;
        RECT 96.170 101.860 101.515 102.405 ;
        RECT 77.770 99.855 83.115 100.290 ;
        RECT 83.290 99.855 88.635 100.290 ;
        RECT 88.805 99.855 89.095 101.020 ;
        RECT 89.265 100.945 89.785 101.485 ;
        RECT 89.955 101.115 90.475 101.655 ;
        RECT 89.265 99.855 90.475 100.945 ;
        RECT 92.240 100.290 92.590 101.540 ;
        RECT 94.070 101.030 94.410 101.860 ;
        RECT 97.760 100.290 98.110 101.540 ;
        RECT 99.590 101.030 99.930 101.860 ;
        RECT 101.685 101.680 101.975 102.405 ;
        RECT 102.145 101.655 103.355 102.405 ;
        RECT 103.530 101.860 108.875 102.405 ;
        RECT 109.050 101.860 114.395 102.405 ;
        RECT 90.650 99.855 95.995 100.290 ;
        RECT 96.170 99.855 101.515 100.290 ;
        RECT 101.685 99.855 101.975 101.020 ;
        RECT 102.145 100.945 102.665 101.485 ;
        RECT 102.835 101.115 103.355 101.655 ;
        RECT 102.145 99.855 103.355 100.945 ;
        RECT 105.120 100.290 105.470 101.540 ;
        RECT 106.950 101.030 107.290 101.860 ;
        RECT 110.640 100.290 110.990 101.540 ;
        RECT 112.470 101.030 112.810 101.860 ;
        RECT 114.565 101.680 114.855 102.405 ;
        RECT 115.490 101.860 120.835 102.405 ;
        RECT 121.010 101.860 126.355 102.405 ;
        RECT 103.530 99.855 108.875 100.290 ;
        RECT 109.050 99.855 114.395 100.290 ;
        RECT 114.565 99.855 114.855 101.020 ;
        RECT 117.080 100.290 117.430 101.540 ;
        RECT 118.910 101.030 119.250 101.860 ;
        RECT 122.600 100.290 122.950 101.540 ;
        RECT 124.430 101.030 124.770 101.860 ;
        RECT 126.525 101.655 127.735 102.405 ;
        RECT 126.525 100.945 127.045 101.485 ;
        RECT 127.215 101.115 127.735 101.655 ;
        RECT 115.490 99.855 120.835 100.290 ;
        RECT 121.010 99.855 126.355 100.290 ;
        RECT 126.525 99.855 127.735 100.945 ;
        RECT 14.660 99.685 127.820 99.855 ;
        RECT 19.165 66.070 30.165 66.940 ;
        RECT 19.165 54.930 20.835 66.070 ;
        RECT 21.465 65.555 26.465 65.725 ;
        RECT 21.235 55.300 21.405 65.340 ;
        RECT 26.525 55.300 26.695 65.340 ;
        RECT 27.095 54.930 27.265 66.070 ;
        RECT 27.895 65.555 28.895 65.725 ;
        RECT 27.665 55.300 27.835 65.340 ;
        RECT 28.955 55.300 29.125 65.340 ;
        RECT 29.525 54.930 30.165 66.070 ;
        RECT 19.165 52.860 30.165 54.930 ;
        RECT 19.165 49.370 21.005 52.860 ;
        RECT 22.765 52.780 30.165 52.860 ;
        RECT 21.635 52.350 22.135 52.520 ;
        RECT 21.405 50.095 21.575 52.135 ;
        RECT 22.195 50.095 22.365 52.135 ;
        RECT 21.635 49.710 22.135 49.880 ;
        RECT 22.765 49.370 25.085 52.780 ;
        RECT 25.715 52.270 26.215 52.440 ;
        RECT 19.165 48.650 25.085 49.370 ;
        RECT 19.135 48.040 23.045 48.260 ;
        RECT 19.135 45.640 20.855 48.040 ;
        RECT 21.485 47.530 21.985 47.700 ;
        RECT 21.255 46.320 21.425 47.360 ;
        RECT 22.045 46.320 22.215 47.360 ;
        RECT 21.485 45.980 21.985 46.150 ;
        RECT 22.615 45.640 23.045 48.040 ;
        RECT 24.025 46.290 25.085 48.650 ;
        RECT 25.485 47.015 25.655 52.055 ;
        RECT 26.275 47.015 26.445 52.055 ;
        RECT 25.715 46.630 26.215 46.800 ;
        RECT 26.845 46.290 27.015 52.780 ;
        RECT 27.645 52.270 28.145 52.440 ;
        RECT 27.415 47.015 27.585 52.055 ;
        RECT 28.205 47.015 28.375 52.055 ;
        RECT 27.645 46.630 28.145 46.800 ;
        RECT 28.775 46.290 30.165 52.780 ;
        RECT 30.365 66.080 41.365 66.950 ;
        RECT 30.365 54.940 32.035 66.080 ;
        RECT 32.665 65.565 37.665 65.735 ;
        RECT 32.435 55.310 32.605 65.350 ;
        RECT 37.725 55.310 37.895 65.350 ;
        RECT 38.295 54.940 38.465 66.080 ;
        RECT 39.095 65.565 40.095 65.735 ;
        RECT 38.865 55.310 39.035 65.350 ;
        RECT 40.155 55.310 40.325 65.350 ;
        RECT 40.725 54.940 41.365 66.080 ;
        RECT 30.365 52.870 41.365 54.940 ;
        RECT 30.365 49.380 32.205 52.870 ;
        RECT 33.965 52.790 41.365 52.870 ;
        RECT 32.835 52.360 33.335 52.530 ;
        RECT 32.605 50.105 32.775 52.145 ;
        RECT 33.395 50.105 33.565 52.145 ;
        RECT 32.835 49.720 33.335 49.890 ;
        RECT 33.965 49.380 36.285 52.790 ;
        RECT 36.915 52.280 37.415 52.450 ;
        RECT 30.365 48.660 36.285 49.380 ;
        RECT 24.025 45.800 30.165 46.290 ;
        RECT 30.335 48.050 34.245 48.270 ;
        RECT 19.135 45.370 23.045 45.640 ;
        RECT 30.335 45.650 32.055 48.050 ;
        RECT 32.685 47.540 33.185 47.710 ;
        RECT 32.455 46.330 32.625 47.370 ;
        RECT 33.245 46.330 33.415 47.370 ;
        RECT 32.685 45.990 33.185 46.160 ;
        RECT 33.815 45.650 34.245 48.050 ;
        RECT 35.225 46.300 36.285 48.660 ;
        RECT 36.685 47.025 36.855 52.065 ;
        RECT 37.475 47.025 37.645 52.065 ;
        RECT 36.915 46.640 37.415 46.810 ;
        RECT 38.045 46.300 38.215 52.790 ;
        RECT 38.845 52.280 39.345 52.450 ;
        RECT 38.615 47.025 38.785 52.065 ;
        RECT 39.405 47.025 39.575 52.065 ;
        RECT 38.845 46.640 39.345 46.810 ;
        RECT 39.975 46.300 41.365 52.790 ;
        RECT 41.585 66.050 52.585 66.920 ;
        RECT 41.585 54.910 43.255 66.050 ;
        RECT 43.885 65.535 48.885 65.705 ;
        RECT 43.655 55.280 43.825 65.320 ;
        RECT 48.945 55.280 49.115 65.320 ;
        RECT 49.515 54.910 49.685 66.050 ;
        RECT 50.315 65.535 51.315 65.705 ;
        RECT 50.085 55.280 50.255 65.320 ;
        RECT 51.375 55.280 51.545 65.320 ;
        RECT 51.945 54.910 52.585 66.050 ;
        RECT 41.585 52.840 52.585 54.910 ;
        RECT 41.585 49.350 43.425 52.840 ;
        RECT 45.185 52.760 52.585 52.840 ;
        RECT 44.055 52.330 44.555 52.500 ;
        RECT 43.825 50.075 43.995 52.115 ;
        RECT 44.615 50.075 44.785 52.115 ;
        RECT 44.055 49.690 44.555 49.860 ;
        RECT 45.185 49.350 47.505 52.760 ;
        RECT 48.135 52.250 48.635 52.420 ;
        RECT 41.585 48.630 47.505 49.350 ;
        RECT 35.225 45.810 41.365 46.300 ;
        RECT 41.555 48.020 45.465 48.240 ;
        RECT 30.335 45.380 34.245 45.650 ;
        RECT 41.555 45.620 43.275 48.020 ;
        RECT 43.905 47.510 44.405 47.680 ;
        RECT 43.675 46.300 43.845 47.340 ;
        RECT 44.465 46.300 44.635 47.340 ;
        RECT 43.905 45.960 44.405 46.130 ;
        RECT 45.035 45.620 45.465 48.020 ;
        RECT 46.445 46.270 47.505 48.630 ;
        RECT 47.905 46.995 48.075 52.035 ;
        RECT 48.695 46.995 48.865 52.035 ;
        RECT 48.135 46.610 48.635 46.780 ;
        RECT 49.265 46.270 49.435 52.760 ;
        RECT 50.065 52.250 50.565 52.420 ;
        RECT 49.835 46.995 50.005 52.035 ;
        RECT 50.625 46.995 50.795 52.035 ;
        RECT 50.065 46.610 50.565 46.780 ;
        RECT 51.195 46.270 52.585 52.760 ;
        RECT 52.835 66.030 63.835 66.900 ;
        RECT 52.835 54.890 54.505 66.030 ;
        RECT 55.135 65.515 60.135 65.685 ;
        RECT 54.905 55.260 55.075 65.300 ;
        RECT 60.195 55.260 60.365 65.300 ;
        RECT 60.765 54.890 60.935 66.030 ;
        RECT 61.565 65.515 62.565 65.685 ;
        RECT 61.335 55.260 61.505 65.300 ;
        RECT 62.625 55.260 62.795 65.300 ;
        RECT 63.195 54.890 63.835 66.030 ;
        RECT 52.835 52.820 63.835 54.890 ;
        RECT 52.835 49.330 54.675 52.820 ;
        RECT 56.435 52.740 63.835 52.820 ;
        RECT 55.305 52.310 55.805 52.480 ;
        RECT 55.075 50.055 55.245 52.095 ;
        RECT 55.865 50.055 56.035 52.095 ;
        RECT 55.305 49.670 55.805 49.840 ;
        RECT 56.435 49.330 58.755 52.740 ;
        RECT 59.385 52.230 59.885 52.400 ;
        RECT 52.835 48.610 58.755 49.330 ;
        RECT 46.445 45.780 52.585 46.270 ;
        RECT 52.805 48.000 56.715 48.220 ;
        RECT 41.555 45.350 45.465 45.620 ;
        RECT 52.805 45.600 54.525 48.000 ;
        RECT 55.155 47.490 55.655 47.660 ;
        RECT 54.925 46.280 55.095 47.320 ;
        RECT 55.715 46.280 55.885 47.320 ;
        RECT 55.155 45.940 55.655 46.110 ;
        RECT 56.285 45.600 56.715 48.000 ;
        RECT 57.695 46.250 58.755 48.610 ;
        RECT 59.155 46.975 59.325 52.015 ;
        RECT 59.945 46.975 60.115 52.015 ;
        RECT 59.385 46.590 59.885 46.760 ;
        RECT 60.515 46.250 60.685 52.740 ;
        RECT 61.315 52.230 61.815 52.400 ;
        RECT 61.085 46.975 61.255 52.015 ;
        RECT 61.875 46.975 62.045 52.015 ;
        RECT 61.315 46.590 61.815 46.760 ;
        RECT 62.445 46.250 63.835 52.740 ;
        RECT 64.055 66.020 75.055 66.890 ;
        RECT 64.055 54.880 65.725 66.020 ;
        RECT 66.355 65.505 71.355 65.675 ;
        RECT 66.125 55.250 66.295 65.290 ;
        RECT 71.415 55.250 71.585 65.290 ;
        RECT 71.985 54.880 72.155 66.020 ;
        RECT 72.785 65.505 73.785 65.675 ;
        RECT 72.555 55.250 72.725 65.290 ;
        RECT 73.845 55.250 74.015 65.290 ;
        RECT 74.415 54.880 75.055 66.020 ;
        RECT 64.055 52.810 75.055 54.880 ;
        RECT 64.055 49.320 65.895 52.810 ;
        RECT 67.655 52.730 75.055 52.810 ;
        RECT 66.525 52.300 67.025 52.470 ;
        RECT 66.295 50.045 66.465 52.085 ;
        RECT 67.085 50.045 67.255 52.085 ;
        RECT 66.525 49.660 67.025 49.830 ;
        RECT 67.655 49.320 69.975 52.730 ;
        RECT 70.605 52.220 71.105 52.390 ;
        RECT 64.055 48.600 69.975 49.320 ;
        RECT 57.695 45.760 63.835 46.250 ;
        RECT 64.025 47.990 67.935 48.210 ;
        RECT 52.805 45.330 56.715 45.600 ;
        RECT 64.025 45.590 65.745 47.990 ;
        RECT 66.375 47.480 66.875 47.650 ;
        RECT 66.145 46.270 66.315 47.310 ;
        RECT 66.935 46.270 67.105 47.310 ;
        RECT 66.375 45.930 66.875 46.100 ;
        RECT 67.505 45.590 67.935 47.990 ;
        RECT 68.915 46.240 69.975 48.600 ;
        RECT 70.375 46.965 70.545 52.005 ;
        RECT 71.165 46.965 71.335 52.005 ;
        RECT 70.605 46.580 71.105 46.750 ;
        RECT 71.735 46.240 71.905 52.730 ;
        RECT 72.535 52.220 73.035 52.390 ;
        RECT 72.305 46.965 72.475 52.005 ;
        RECT 73.095 46.965 73.265 52.005 ;
        RECT 72.535 46.580 73.035 46.750 ;
        RECT 73.665 46.240 75.055 52.730 ;
        RECT 75.295 66.010 86.295 66.880 ;
        RECT 75.295 54.870 76.965 66.010 ;
        RECT 77.595 65.495 82.595 65.665 ;
        RECT 77.365 55.240 77.535 65.280 ;
        RECT 82.655 55.240 82.825 65.280 ;
        RECT 83.225 54.870 83.395 66.010 ;
        RECT 84.025 65.495 85.025 65.665 ;
        RECT 83.795 55.240 83.965 65.280 ;
        RECT 85.085 55.240 85.255 65.280 ;
        RECT 85.655 54.870 86.295 66.010 ;
        RECT 75.295 52.800 86.295 54.870 ;
        RECT 75.295 49.310 77.135 52.800 ;
        RECT 78.895 52.720 86.295 52.800 ;
        RECT 77.765 52.290 78.265 52.460 ;
        RECT 77.535 50.035 77.705 52.075 ;
        RECT 78.325 50.035 78.495 52.075 ;
        RECT 77.765 49.650 78.265 49.820 ;
        RECT 78.895 49.310 81.215 52.720 ;
        RECT 81.845 52.210 82.345 52.380 ;
        RECT 75.295 48.590 81.215 49.310 ;
        RECT 68.915 45.750 75.055 46.240 ;
        RECT 75.265 47.980 79.175 48.200 ;
        RECT 64.025 45.320 67.935 45.590 ;
        RECT 75.265 45.580 76.985 47.980 ;
        RECT 77.615 47.470 78.115 47.640 ;
        RECT 77.385 46.260 77.555 47.300 ;
        RECT 78.175 46.260 78.345 47.300 ;
        RECT 77.615 45.920 78.115 46.090 ;
        RECT 78.745 45.580 79.175 47.980 ;
        RECT 80.155 46.230 81.215 48.590 ;
        RECT 81.615 46.955 81.785 51.995 ;
        RECT 82.405 46.955 82.575 51.995 ;
        RECT 81.845 46.570 82.345 46.740 ;
        RECT 82.975 46.230 83.145 52.720 ;
        RECT 83.775 52.210 84.275 52.380 ;
        RECT 83.545 46.955 83.715 51.995 ;
        RECT 84.335 46.955 84.505 51.995 ;
        RECT 83.775 46.570 84.275 46.740 ;
        RECT 84.905 46.230 86.295 52.720 ;
        RECT 86.545 66.020 97.545 66.890 ;
        RECT 131.125 66.880 140.025 66.890 ;
        RECT 86.545 54.880 88.215 66.020 ;
        RECT 88.845 65.505 93.845 65.675 ;
        RECT 88.615 55.250 88.785 65.290 ;
        RECT 93.905 55.250 94.075 65.290 ;
        RECT 94.475 54.880 94.645 66.020 ;
        RECT 95.275 65.505 96.275 65.675 ;
        RECT 95.045 55.250 95.215 65.290 ;
        RECT 96.335 55.250 96.505 65.290 ;
        RECT 96.905 54.880 97.545 66.020 ;
        RECT 86.545 52.810 97.545 54.880 ;
        RECT 86.545 49.320 88.385 52.810 ;
        RECT 90.145 52.730 97.545 52.810 ;
        RECT 89.015 52.300 89.515 52.470 ;
        RECT 88.785 50.045 88.955 52.085 ;
        RECT 89.575 50.045 89.745 52.085 ;
        RECT 89.015 49.660 89.515 49.830 ;
        RECT 90.145 49.320 92.465 52.730 ;
        RECT 93.095 52.220 93.595 52.390 ;
        RECT 86.545 48.600 92.465 49.320 ;
        RECT 80.155 45.740 86.295 46.230 ;
        RECT 86.515 47.990 90.425 48.210 ;
        RECT 75.265 45.310 79.175 45.580 ;
        RECT 86.515 45.590 88.235 47.990 ;
        RECT 88.865 47.480 89.365 47.650 ;
        RECT 88.635 46.270 88.805 47.310 ;
        RECT 89.425 46.270 89.595 47.310 ;
        RECT 88.865 45.930 89.365 46.100 ;
        RECT 89.995 45.590 90.425 47.990 ;
        RECT 91.405 46.240 92.465 48.600 ;
        RECT 92.865 46.965 93.035 52.005 ;
        RECT 93.655 46.965 93.825 52.005 ;
        RECT 93.095 46.580 93.595 46.750 ;
        RECT 94.225 46.240 94.395 52.730 ;
        RECT 95.025 52.220 95.525 52.390 ;
        RECT 94.795 46.965 94.965 52.005 ;
        RECT 95.585 46.965 95.755 52.005 ;
        RECT 95.025 46.580 95.525 46.750 ;
        RECT 96.155 46.240 97.545 52.730 ;
        RECT 97.825 66.010 108.825 66.880 ;
        RECT 97.825 54.870 99.495 66.010 ;
        RECT 100.125 65.495 105.125 65.665 ;
        RECT 99.895 55.240 100.065 65.280 ;
        RECT 105.185 55.240 105.355 65.280 ;
        RECT 105.755 54.870 105.925 66.010 ;
        RECT 106.555 65.495 107.555 65.665 ;
        RECT 106.325 55.240 106.495 65.280 ;
        RECT 107.615 55.240 107.785 65.280 ;
        RECT 108.185 54.870 108.825 66.010 ;
        RECT 97.825 52.800 108.825 54.870 ;
        RECT 97.825 49.310 99.665 52.800 ;
        RECT 101.425 52.720 108.825 52.800 ;
        RECT 100.295 52.290 100.795 52.460 ;
        RECT 100.065 50.035 100.235 52.075 ;
        RECT 100.855 50.035 101.025 52.075 ;
        RECT 100.295 49.650 100.795 49.820 ;
        RECT 101.425 49.310 103.745 52.720 ;
        RECT 104.375 52.210 104.875 52.380 ;
        RECT 97.825 48.590 103.745 49.310 ;
        RECT 91.405 45.750 97.545 46.240 ;
        RECT 97.795 47.980 101.705 48.200 ;
        RECT 86.515 45.320 90.425 45.590 ;
        RECT 97.795 45.580 99.515 47.980 ;
        RECT 100.145 47.470 100.645 47.640 ;
        RECT 99.915 46.260 100.085 47.300 ;
        RECT 100.705 46.260 100.875 47.300 ;
        RECT 100.145 45.920 100.645 46.090 ;
        RECT 101.275 45.580 101.705 47.980 ;
        RECT 102.685 46.230 103.745 48.590 ;
        RECT 104.145 46.955 104.315 51.995 ;
        RECT 104.935 46.955 105.105 51.995 ;
        RECT 104.375 46.570 104.875 46.740 ;
        RECT 105.505 46.230 105.675 52.720 ;
        RECT 106.305 52.210 106.805 52.380 ;
        RECT 106.075 46.955 106.245 51.995 ;
        RECT 106.865 46.955 107.035 51.995 ;
        RECT 106.305 46.570 106.805 46.740 ;
        RECT 107.435 46.230 108.825 52.720 ;
        RECT 109.095 66.010 120.095 66.880 ;
        RECT 109.095 54.870 110.765 66.010 ;
        RECT 111.395 65.495 116.395 65.665 ;
        RECT 111.165 55.240 111.335 65.280 ;
        RECT 116.455 55.240 116.625 65.280 ;
        RECT 117.025 54.870 117.195 66.010 ;
        RECT 117.825 65.495 118.825 65.665 ;
        RECT 117.595 55.240 117.765 65.280 ;
        RECT 118.885 55.240 119.055 65.280 ;
        RECT 119.455 54.870 120.095 66.010 ;
        RECT 109.095 52.800 120.095 54.870 ;
        RECT 109.095 49.310 110.935 52.800 ;
        RECT 112.695 52.720 120.095 52.800 ;
        RECT 111.565 52.290 112.065 52.460 ;
        RECT 111.335 50.035 111.505 52.075 ;
        RECT 112.125 50.035 112.295 52.075 ;
        RECT 111.565 49.650 112.065 49.820 ;
        RECT 112.695 49.310 115.015 52.720 ;
        RECT 115.645 52.210 116.145 52.380 ;
        RECT 109.095 48.590 115.015 49.310 ;
        RECT 102.685 45.740 108.825 46.230 ;
        RECT 109.065 47.980 112.975 48.200 ;
        RECT 97.795 45.310 101.705 45.580 ;
        RECT 109.065 45.580 110.785 47.980 ;
        RECT 111.415 47.470 111.915 47.640 ;
        RECT 111.185 46.260 111.355 47.300 ;
        RECT 111.975 46.260 112.145 47.300 ;
        RECT 111.415 45.920 111.915 46.090 ;
        RECT 112.545 45.580 112.975 47.980 ;
        RECT 113.955 46.230 115.015 48.590 ;
        RECT 115.415 46.955 115.585 51.995 ;
        RECT 116.205 46.955 116.375 51.995 ;
        RECT 115.645 46.570 116.145 46.740 ;
        RECT 116.775 46.230 116.945 52.720 ;
        RECT 117.575 52.210 118.075 52.380 ;
        RECT 117.345 46.955 117.515 51.995 ;
        RECT 118.135 46.955 118.305 51.995 ;
        RECT 117.575 46.570 118.075 46.740 ;
        RECT 118.705 46.230 120.095 52.720 ;
        RECT 120.345 66.010 140.025 66.880 ;
        RECT 120.345 54.870 122.015 66.010 ;
        RECT 122.645 65.495 127.645 65.665 ;
        RECT 122.415 55.240 122.585 65.280 ;
        RECT 127.705 55.240 127.875 65.280 ;
        RECT 128.275 54.870 128.445 66.010 ;
        RECT 130.705 65.980 140.025 66.010 ;
        RECT 129.075 65.495 130.075 65.665 ;
        RECT 128.845 55.240 129.015 65.280 ;
        RECT 130.135 55.240 130.305 65.280 ;
        RECT 130.705 54.870 132.765 65.980 ;
        RECT 133.395 65.465 138.395 65.635 ;
        RECT 133.165 55.210 133.335 65.250 ;
        RECT 138.455 55.210 138.625 65.250 ;
        RECT 120.345 54.840 132.765 54.870 ;
        RECT 139.025 54.840 140.025 65.980 ;
        RECT 120.345 54.720 140.025 54.840 ;
        RECT 120.345 53.550 140.035 54.720 ;
        RECT 120.345 52.800 131.345 53.550 ;
        RECT 120.345 49.310 122.185 52.800 ;
        RECT 123.945 52.720 131.345 52.800 ;
        RECT 122.815 52.290 123.315 52.460 ;
        RECT 122.585 50.035 122.755 52.075 ;
        RECT 123.375 50.035 123.545 52.075 ;
        RECT 122.815 49.650 123.315 49.820 ;
        RECT 123.945 49.310 126.265 52.720 ;
        RECT 126.895 52.210 127.395 52.380 ;
        RECT 120.345 48.590 126.265 49.310 ;
        RECT 113.955 45.740 120.095 46.230 ;
        RECT 120.315 47.980 124.225 48.200 ;
        RECT 109.065 45.310 112.975 45.580 ;
        RECT 120.315 45.580 122.035 47.980 ;
        RECT 122.665 47.470 123.165 47.640 ;
        RECT 122.435 46.260 122.605 47.300 ;
        RECT 123.225 46.260 123.395 47.300 ;
        RECT 122.665 45.920 123.165 46.090 ;
        RECT 123.795 45.580 124.225 47.980 ;
        RECT 125.205 46.230 126.265 48.590 ;
        RECT 126.665 46.955 126.835 51.995 ;
        RECT 127.455 46.955 127.625 51.995 ;
        RECT 126.895 46.570 127.395 46.740 ;
        RECT 128.025 46.230 128.195 52.720 ;
        RECT 128.825 52.210 129.325 52.380 ;
        RECT 128.595 46.955 128.765 51.995 ;
        RECT 129.385 46.955 129.555 51.995 ;
        RECT 128.825 46.570 129.325 46.740 ;
        RECT 129.955 46.230 131.345 52.720 ;
        RECT 125.205 45.740 131.345 46.230 ;
        RECT 120.315 45.310 124.225 45.580 ;
        RECT 25.695 39.770 29.605 40.040 ;
        RECT 18.575 39.120 24.715 39.610 ;
        RECT 18.575 32.630 19.965 39.120 ;
        RECT 20.595 38.610 21.095 38.780 ;
        RECT 20.365 33.355 20.535 38.395 ;
        RECT 21.155 33.355 21.325 38.395 ;
        RECT 20.595 32.970 21.095 33.140 ;
        RECT 21.725 32.630 21.895 39.120 ;
        RECT 22.525 38.610 23.025 38.780 ;
        RECT 22.295 33.355 22.465 38.395 ;
        RECT 23.085 33.355 23.255 38.395 ;
        RECT 23.655 36.760 24.715 39.120 ;
        RECT 25.695 37.370 26.125 39.770 ;
        RECT 26.755 39.260 27.255 39.430 ;
        RECT 26.525 38.050 26.695 39.090 ;
        RECT 27.315 38.050 27.485 39.090 ;
        RECT 26.755 37.710 27.255 37.880 ;
        RECT 27.885 37.370 29.605 39.770 ;
        RECT 36.975 39.770 40.885 40.040 ;
        RECT 25.695 37.150 29.605 37.370 ;
        RECT 29.855 39.120 35.995 39.610 ;
        RECT 23.655 36.040 29.575 36.760 ;
        RECT 22.525 32.970 23.025 33.140 ;
        RECT 23.655 32.630 25.975 36.040 ;
        RECT 26.605 35.530 27.105 35.700 ;
        RECT 26.375 33.275 26.545 35.315 ;
        RECT 27.165 33.275 27.335 35.315 ;
        RECT 26.605 32.890 27.105 33.060 ;
        RECT 18.575 32.550 25.975 32.630 ;
        RECT 27.735 32.550 29.575 36.040 ;
        RECT 18.575 30.480 29.575 32.550 ;
        RECT 18.575 19.340 19.215 30.480 ;
        RECT 19.615 20.070 19.785 30.110 ;
        RECT 20.905 20.070 21.075 30.110 ;
        RECT 19.845 19.685 20.845 19.855 ;
        RECT 21.475 19.340 21.645 30.480 ;
        RECT 22.045 20.070 22.215 30.110 ;
        RECT 27.335 20.070 27.505 30.110 ;
        RECT 22.275 19.685 27.275 19.855 ;
        RECT 27.905 19.340 29.575 30.480 ;
        RECT 18.575 18.470 29.575 19.340 ;
        RECT 29.855 32.630 31.245 39.120 ;
        RECT 31.875 38.610 32.375 38.780 ;
        RECT 31.645 33.355 31.815 38.395 ;
        RECT 32.435 33.355 32.605 38.395 ;
        RECT 31.875 32.970 32.375 33.140 ;
        RECT 33.005 32.630 33.175 39.120 ;
        RECT 33.805 38.610 34.305 38.780 ;
        RECT 33.575 33.355 33.745 38.395 ;
        RECT 34.365 33.355 34.535 38.395 ;
        RECT 34.935 36.760 35.995 39.120 ;
        RECT 36.975 37.370 37.405 39.770 ;
        RECT 38.035 39.260 38.535 39.430 ;
        RECT 37.805 38.050 37.975 39.090 ;
        RECT 38.595 38.050 38.765 39.090 ;
        RECT 38.035 37.710 38.535 37.880 ;
        RECT 39.165 37.370 40.885 39.770 ;
        RECT 48.265 39.750 52.175 40.020 ;
        RECT 36.975 37.150 40.885 37.370 ;
        RECT 41.145 39.100 47.285 39.590 ;
        RECT 34.935 36.040 40.855 36.760 ;
        RECT 33.805 32.970 34.305 33.140 ;
        RECT 34.935 32.630 37.255 36.040 ;
        RECT 37.885 35.530 38.385 35.700 ;
        RECT 37.655 33.275 37.825 35.315 ;
        RECT 38.445 33.275 38.615 35.315 ;
        RECT 37.885 32.890 38.385 33.060 ;
        RECT 29.855 32.550 37.255 32.630 ;
        RECT 39.015 32.550 40.855 36.040 ;
        RECT 29.855 30.480 40.855 32.550 ;
        RECT 29.855 19.340 30.495 30.480 ;
        RECT 30.895 20.070 31.065 30.110 ;
        RECT 32.185 20.070 32.355 30.110 ;
        RECT 31.125 19.685 32.125 19.855 ;
        RECT 32.755 19.340 32.925 30.480 ;
        RECT 33.325 20.070 33.495 30.110 ;
        RECT 38.615 20.070 38.785 30.110 ;
        RECT 33.555 19.685 38.555 19.855 ;
        RECT 39.185 19.340 40.855 30.480 ;
        RECT 29.855 18.470 40.855 19.340 ;
        RECT 41.145 32.610 42.535 39.100 ;
        RECT 43.165 38.590 43.665 38.760 ;
        RECT 42.935 33.335 43.105 38.375 ;
        RECT 43.725 33.335 43.895 38.375 ;
        RECT 43.165 32.950 43.665 33.120 ;
        RECT 44.295 32.610 44.465 39.100 ;
        RECT 45.095 38.590 45.595 38.760 ;
        RECT 44.865 33.335 45.035 38.375 ;
        RECT 45.655 33.335 45.825 38.375 ;
        RECT 46.225 36.740 47.285 39.100 ;
        RECT 48.265 37.350 48.695 39.750 ;
        RECT 49.325 39.240 49.825 39.410 ;
        RECT 49.095 38.030 49.265 39.070 ;
        RECT 49.885 38.030 50.055 39.070 ;
        RECT 49.325 37.690 49.825 37.860 ;
        RECT 50.455 37.350 52.175 39.750 ;
        RECT 59.485 39.750 63.395 40.020 ;
        RECT 48.265 37.130 52.175 37.350 ;
        RECT 52.365 39.100 58.505 39.590 ;
        RECT 46.225 36.020 52.145 36.740 ;
        RECT 45.095 32.950 45.595 33.120 ;
        RECT 46.225 32.610 48.545 36.020 ;
        RECT 49.175 35.510 49.675 35.680 ;
        RECT 48.945 33.255 49.115 35.295 ;
        RECT 49.735 33.255 49.905 35.295 ;
        RECT 49.175 32.870 49.675 33.040 ;
        RECT 41.145 32.530 48.545 32.610 ;
        RECT 50.305 32.530 52.145 36.020 ;
        RECT 41.145 30.460 52.145 32.530 ;
        RECT 41.145 19.320 41.785 30.460 ;
        RECT 42.185 20.050 42.355 30.090 ;
        RECT 43.475 20.050 43.645 30.090 ;
        RECT 42.415 19.665 43.415 19.835 ;
        RECT 44.045 19.320 44.215 30.460 ;
        RECT 44.615 20.050 44.785 30.090 ;
        RECT 49.905 20.050 50.075 30.090 ;
        RECT 44.845 19.665 49.845 19.835 ;
        RECT 50.475 19.320 52.145 30.460 ;
        RECT 41.145 18.450 52.145 19.320 ;
        RECT 52.365 32.610 53.755 39.100 ;
        RECT 54.385 38.590 54.885 38.760 ;
        RECT 54.155 33.335 54.325 38.375 ;
        RECT 54.945 33.335 55.115 38.375 ;
        RECT 54.385 32.950 54.885 33.120 ;
        RECT 55.515 32.610 55.685 39.100 ;
        RECT 56.315 38.590 56.815 38.760 ;
        RECT 56.085 33.335 56.255 38.375 ;
        RECT 56.875 33.335 57.045 38.375 ;
        RECT 57.445 36.740 58.505 39.100 ;
        RECT 59.485 37.350 59.915 39.750 ;
        RECT 60.545 39.240 61.045 39.410 ;
        RECT 60.315 38.030 60.485 39.070 ;
        RECT 61.105 38.030 61.275 39.070 ;
        RECT 60.545 37.690 61.045 37.860 ;
        RECT 61.675 37.350 63.395 39.750 ;
        RECT 70.685 39.750 74.595 40.020 ;
        RECT 59.485 37.130 63.395 37.350 ;
        RECT 63.565 39.100 69.705 39.590 ;
        RECT 57.445 36.020 63.365 36.740 ;
        RECT 56.315 32.950 56.815 33.120 ;
        RECT 57.445 32.610 59.765 36.020 ;
        RECT 60.395 35.510 60.895 35.680 ;
        RECT 60.165 33.255 60.335 35.295 ;
        RECT 60.955 33.255 61.125 35.295 ;
        RECT 60.395 32.870 60.895 33.040 ;
        RECT 52.365 32.530 59.765 32.610 ;
        RECT 61.525 32.530 63.365 36.020 ;
        RECT 52.365 30.460 63.365 32.530 ;
        RECT 52.365 19.320 53.005 30.460 ;
        RECT 53.405 20.050 53.575 30.090 ;
        RECT 54.695 20.050 54.865 30.090 ;
        RECT 53.635 19.665 54.635 19.835 ;
        RECT 55.265 19.320 55.435 30.460 ;
        RECT 55.835 20.050 56.005 30.090 ;
        RECT 61.125 20.050 61.295 30.090 ;
        RECT 56.065 19.665 61.065 19.835 ;
        RECT 61.695 19.320 63.365 30.460 ;
        RECT 52.365 18.450 63.365 19.320 ;
        RECT 63.565 32.610 64.955 39.100 ;
        RECT 65.585 38.590 66.085 38.760 ;
        RECT 65.355 33.335 65.525 38.375 ;
        RECT 66.145 33.335 66.315 38.375 ;
        RECT 65.585 32.950 66.085 33.120 ;
        RECT 66.715 32.610 66.885 39.100 ;
        RECT 67.515 38.590 68.015 38.760 ;
        RECT 67.285 33.335 67.455 38.375 ;
        RECT 68.075 33.335 68.245 38.375 ;
        RECT 68.645 36.740 69.705 39.100 ;
        RECT 70.685 37.350 71.115 39.750 ;
        RECT 71.745 39.240 72.245 39.410 ;
        RECT 71.515 38.030 71.685 39.070 ;
        RECT 72.305 38.030 72.475 39.070 ;
        RECT 71.745 37.690 72.245 37.860 ;
        RECT 72.875 37.350 74.595 39.750 ;
        RECT 81.975 39.740 85.885 40.010 ;
        RECT 70.685 37.130 74.595 37.350 ;
        RECT 74.855 39.090 80.995 39.580 ;
        RECT 68.645 36.020 74.565 36.740 ;
        RECT 67.515 32.950 68.015 33.120 ;
        RECT 68.645 32.610 70.965 36.020 ;
        RECT 71.595 35.510 72.095 35.680 ;
        RECT 71.365 33.255 71.535 35.295 ;
        RECT 72.155 33.255 72.325 35.295 ;
        RECT 71.595 32.870 72.095 33.040 ;
        RECT 63.565 32.530 70.965 32.610 ;
        RECT 72.725 32.530 74.565 36.020 ;
        RECT 63.565 30.460 74.565 32.530 ;
        RECT 63.565 19.320 64.205 30.460 ;
        RECT 64.605 20.050 64.775 30.090 ;
        RECT 65.895 20.050 66.065 30.090 ;
        RECT 64.835 19.665 65.835 19.835 ;
        RECT 66.465 19.320 66.635 30.460 ;
        RECT 67.035 20.050 67.205 30.090 ;
        RECT 72.325 20.050 72.495 30.090 ;
        RECT 67.265 19.665 72.265 19.835 ;
        RECT 72.895 19.320 74.565 30.460 ;
        RECT 63.565 18.450 74.565 19.320 ;
        RECT 74.855 32.600 76.245 39.090 ;
        RECT 76.875 38.580 77.375 38.750 ;
        RECT 76.645 33.325 76.815 38.365 ;
        RECT 77.435 33.325 77.605 38.365 ;
        RECT 76.875 32.940 77.375 33.110 ;
        RECT 78.005 32.600 78.175 39.090 ;
        RECT 78.805 38.580 79.305 38.750 ;
        RECT 78.575 33.325 78.745 38.365 ;
        RECT 79.365 33.325 79.535 38.365 ;
        RECT 79.935 36.730 80.995 39.090 ;
        RECT 81.975 37.340 82.405 39.740 ;
        RECT 83.035 39.230 83.535 39.400 ;
        RECT 82.805 38.020 82.975 39.060 ;
        RECT 83.595 38.020 83.765 39.060 ;
        RECT 83.035 37.680 83.535 37.850 ;
        RECT 84.165 37.340 85.885 39.740 ;
        RECT 93.215 39.760 97.125 40.030 ;
        RECT 81.975 37.120 85.885 37.340 ;
        RECT 86.095 39.110 92.235 39.600 ;
        RECT 79.935 36.010 85.855 36.730 ;
        RECT 78.805 32.940 79.305 33.110 ;
        RECT 79.935 32.600 82.255 36.010 ;
        RECT 82.885 35.500 83.385 35.670 ;
        RECT 82.655 33.245 82.825 35.285 ;
        RECT 83.445 33.245 83.615 35.285 ;
        RECT 82.885 32.860 83.385 33.030 ;
        RECT 74.855 32.520 82.255 32.600 ;
        RECT 84.015 32.520 85.855 36.010 ;
        RECT 74.855 30.450 85.855 32.520 ;
        RECT 74.855 19.310 75.495 30.450 ;
        RECT 75.895 20.040 76.065 30.080 ;
        RECT 77.185 20.040 77.355 30.080 ;
        RECT 76.125 19.655 77.125 19.825 ;
        RECT 77.755 19.310 77.925 30.450 ;
        RECT 78.325 20.040 78.495 30.080 ;
        RECT 83.615 20.040 83.785 30.080 ;
        RECT 78.555 19.655 83.555 19.825 ;
        RECT 84.185 19.310 85.855 30.450 ;
        RECT 74.855 18.440 85.855 19.310 ;
        RECT 86.095 32.620 87.485 39.110 ;
        RECT 88.115 38.600 88.615 38.770 ;
        RECT 87.885 33.345 88.055 38.385 ;
        RECT 88.675 33.345 88.845 38.385 ;
        RECT 88.115 32.960 88.615 33.130 ;
        RECT 89.245 32.620 89.415 39.110 ;
        RECT 90.045 38.600 90.545 38.770 ;
        RECT 89.815 33.345 89.985 38.385 ;
        RECT 90.605 33.345 90.775 38.385 ;
        RECT 91.175 36.750 92.235 39.110 ;
        RECT 93.215 37.360 93.645 39.760 ;
        RECT 94.275 39.250 94.775 39.420 ;
        RECT 94.045 38.040 94.215 39.080 ;
        RECT 94.835 38.040 95.005 39.080 ;
        RECT 94.275 37.700 94.775 37.870 ;
        RECT 95.405 37.360 97.125 39.760 ;
        RECT 104.425 39.780 108.335 40.050 ;
        RECT 93.215 37.140 97.125 37.360 ;
        RECT 97.305 39.130 103.445 39.620 ;
        RECT 91.175 36.030 97.095 36.750 ;
        RECT 90.045 32.960 90.545 33.130 ;
        RECT 91.175 32.620 93.495 36.030 ;
        RECT 94.125 35.520 94.625 35.690 ;
        RECT 93.895 33.265 94.065 35.305 ;
        RECT 94.685 33.265 94.855 35.305 ;
        RECT 94.125 32.880 94.625 33.050 ;
        RECT 86.095 32.540 93.495 32.620 ;
        RECT 95.255 32.540 97.095 36.030 ;
        RECT 86.095 30.470 97.095 32.540 ;
        RECT 86.095 19.330 86.735 30.470 ;
        RECT 87.135 20.060 87.305 30.100 ;
        RECT 88.425 20.060 88.595 30.100 ;
        RECT 87.365 19.675 88.365 19.845 ;
        RECT 88.995 19.330 89.165 30.470 ;
        RECT 89.565 20.060 89.735 30.100 ;
        RECT 94.855 20.060 95.025 30.100 ;
        RECT 89.795 19.675 94.795 19.845 ;
        RECT 95.425 19.330 97.095 30.470 ;
        RECT 86.095 18.460 97.095 19.330 ;
        RECT 97.305 32.640 98.695 39.130 ;
        RECT 99.325 38.620 99.825 38.790 ;
        RECT 99.095 33.365 99.265 38.405 ;
        RECT 99.885 33.365 100.055 38.405 ;
        RECT 99.325 32.980 99.825 33.150 ;
        RECT 100.455 32.640 100.625 39.130 ;
        RECT 101.255 38.620 101.755 38.790 ;
        RECT 101.025 33.365 101.195 38.405 ;
        RECT 101.815 33.365 101.985 38.405 ;
        RECT 102.385 36.770 103.445 39.130 ;
        RECT 104.425 37.380 104.855 39.780 ;
        RECT 105.485 39.270 105.985 39.440 ;
        RECT 105.255 38.060 105.425 39.100 ;
        RECT 106.045 38.060 106.215 39.100 ;
        RECT 105.485 37.720 105.985 37.890 ;
        RECT 106.615 37.380 108.335 39.780 ;
        RECT 115.625 39.820 119.535 40.090 ;
        RECT 104.425 37.160 108.335 37.380 ;
        RECT 108.505 39.170 114.645 39.660 ;
        RECT 102.385 36.050 108.305 36.770 ;
        RECT 101.255 32.980 101.755 33.150 ;
        RECT 102.385 32.640 104.705 36.050 ;
        RECT 105.335 35.540 105.835 35.710 ;
        RECT 105.105 33.285 105.275 35.325 ;
        RECT 105.895 33.285 106.065 35.325 ;
        RECT 105.335 32.900 105.835 33.070 ;
        RECT 97.305 32.560 104.705 32.640 ;
        RECT 106.465 32.560 108.305 36.050 ;
        RECT 97.305 30.490 108.305 32.560 ;
        RECT 97.305 19.350 97.945 30.490 ;
        RECT 98.345 20.080 98.515 30.120 ;
        RECT 99.635 20.080 99.805 30.120 ;
        RECT 98.575 19.695 99.575 19.865 ;
        RECT 100.205 19.350 100.375 30.490 ;
        RECT 100.775 20.080 100.945 30.120 ;
        RECT 106.065 20.080 106.235 30.120 ;
        RECT 101.005 19.695 106.005 19.865 ;
        RECT 106.635 19.350 108.305 30.490 ;
        RECT 97.305 18.480 108.305 19.350 ;
        RECT 108.505 32.680 109.895 39.170 ;
        RECT 110.525 38.660 111.025 38.830 ;
        RECT 110.295 33.405 110.465 38.445 ;
        RECT 111.085 33.405 111.255 38.445 ;
        RECT 110.525 33.020 111.025 33.190 ;
        RECT 111.655 32.680 111.825 39.170 ;
        RECT 112.455 38.660 112.955 38.830 ;
        RECT 112.225 33.405 112.395 38.445 ;
        RECT 113.015 33.405 113.185 38.445 ;
        RECT 113.585 36.810 114.645 39.170 ;
        RECT 115.625 37.420 116.055 39.820 ;
        RECT 116.685 39.310 117.185 39.480 ;
        RECT 116.455 38.100 116.625 39.140 ;
        RECT 117.245 38.100 117.415 39.140 ;
        RECT 116.685 37.760 117.185 37.930 ;
        RECT 117.815 37.420 119.535 39.820 ;
        RECT 126.835 39.840 130.745 40.110 ;
        RECT 115.625 37.200 119.535 37.420 ;
        RECT 119.715 39.190 125.855 39.680 ;
        RECT 113.585 36.090 119.505 36.810 ;
        RECT 112.455 33.020 112.955 33.190 ;
        RECT 113.585 32.680 115.905 36.090 ;
        RECT 116.535 35.580 117.035 35.750 ;
        RECT 116.305 33.325 116.475 35.365 ;
        RECT 117.095 33.325 117.265 35.365 ;
        RECT 116.535 32.940 117.035 33.110 ;
        RECT 108.505 32.600 115.905 32.680 ;
        RECT 117.665 32.600 119.505 36.090 ;
        RECT 108.505 30.530 119.505 32.600 ;
        RECT 108.505 19.390 109.145 30.530 ;
        RECT 109.545 20.120 109.715 30.160 ;
        RECT 110.835 20.120 111.005 30.160 ;
        RECT 109.775 19.735 110.775 19.905 ;
        RECT 111.405 19.390 111.575 30.530 ;
        RECT 111.975 20.120 112.145 30.160 ;
        RECT 117.265 20.120 117.435 30.160 ;
        RECT 112.205 19.735 117.205 19.905 ;
        RECT 117.835 19.390 119.505 30.530 ;
        RECT 108.505 18.520 119.505 19.390 ;
        RECT 119.715 32.700 121.105 39.190 ;
        RECT 121.735 38.680 122.235 38.850 ;
        RECT 121.505 33.425 121.675 38.465 ;
        RECT 122.295 33.425 122.465 38.465 ;
        RECT 121.735 33.040 122.235 33.210 ;
        RECT 122.865 32.700 123.035 39.190 ;
        RECT 123.665 38.680 124.165 38.850 ;
        RECT 123.435 33.425 123.605 38.465 ;
        RECT 124.225 33.425 124.395 38.465 ;
        RECT 124.795 36.830 125.855 39.190 ;
        RECT 126.835 37.440 127.265 39.840 ;
        RECT 127.895 39.330 128.395 39.500 ;
        RECT 127.665 38.120 127.835 39.160 ;
        RECT 128.455 38.120 128.625 39.160 ;
        RECT 127.895 37.780 128.395 37.950 ;
        RECT 129.025 37.440 130.745 39.840 ;
        RECT 126.835 37.220 130.745 37.440 ;
        RECT 124.795 36.110 130.715 36.830 ;
        RECT 123.665 33.040 124.165 33.210 ;
        RECT 124.795 32.700 127.115 36.110 ;
        RECT 127.745 35.600 128.245 35.770 ;
        RECT 127.515 33.345 127.685 35.385 ;
        RECT 128.305 33.345 128.475 35.385 ;
        RECT 127.745 32.960 128.245 33.130 ;
        RECT 119.715 32.620 127.115 32.700 ;
        RECT 128.875 32.620 130.715 36.110 ;
        RECT 119.715 31.140 130.715 32.620 ;
        RECT 119.715 30.550 139.465 31.140 ;
        RECT 119.715 19.410 120.355 30.550 ;
        RECT 120.755 20.140 120.925 30.180 ;
        RECT 122.045 20.140 122.215 30.180 ;
        RECT 120.985 19.755 121.985 19.925 ;
        RECT 122.615 19.410 122.785 30.550 ;
        RECT 129.045 30.520 139.465 30.550 ;
        RECT 123.185 20.140 123.355 30.180 ;
        RECT 128.475 20.140 128.645 30.180 ;
        RECT 123.415 19.755 128.415 19.925 ;
        RECT 129.045 19.410 132.075 30.520 ;
        RECT 132.475 20.110 132.645 30.150 ;
        RECT 137.765 20.110 137.935 30.150 ;
        RECT 132.705 19.725 137.705 19.895 ;
        RECT 119.715 19.380 132.075 19.410 ;
        RECT 138.335 19.380 139.465 30.520 ;
        RECT 119.715 18.540 139.465 19.380 ;
        RECT 131.925 18.520 139.465 18.540 ;
      LAYER met1 ;
        RECT 135.340 223.880 136.790 225.180 ;
        RECT 14.660 211.050 127.820 211.530 ;
        RECT 14.660 208.330 127.820 208.810 ;
        RECT 14.660 205.610 127.820 206.090 ;
        RECT 14.660 202.890 127.820 203.370 ;
        RECT 61.765 202.350 62.055 202.395 ;
        RECT 64.885 202.350 65.175 202.395 ;
        RECT 66.775 202.350 67.065 202.395 ;
        RECT 61.765 202.210 67.065 202.350 ;
        RECT 61.765 202.165 62.055 202.210 ;
        RECT 64.885 202.165 65.175 202.210 ;
        RECT 66.775 202.165 67.065 202.210 ;
        RECT 58.905 202.010 59.195 202.055 ;
        RECT 64.410 202.010 64.730 202.070 ;
        RECT 58.905 201.870 64.730 202.010 ;
        RECT 58.905 201.825 59.195 201.870 ;
        RECT 64.410 201.810 64.730 201.870 ;
        RECT 60.685 201.375 60.975 201.690 ;
        RECT 61.765 201.670 62.055 201.715 ;
        RECT 65.345 201.670 65.635 201.715 ;
        RECT 67.180 201.670 67.470 201.715 ;
        RECT 61.765 201.530 67.470 201.670 ;
        RECT 61.765 201.485 62.055 201.530 ;
        RECT 65.345 201.485 65.635 201.530 ;
        RECT 67.180 201.485 67.470 201.530 ;
        RECT 67.645 201.670 67.935 201.715 ;
        RECT 68.550 201.670 68.870 201.730 ;
        RECT 67.645 201.530 68.870 201.670 ;
        RECT 67.645 201.485 67.935 201.530 ;
        RECT 68.550 201.470 68.870 201.530 ;
        RECT 60.385 201.330 60.975 201.375 ;
        RECT 62.570 201.330 62.890 201.390 ;
        RECT 63.625 201.330 64.275 201.375 ;
        RECT 60.385 201.190 64.275 201.330 ;
        RECT 60.385 201.145 60.675 201.190 ;
        RECT 62.570 201.130 62.890 201.190 ;
        RECT 63.625 201.145 64.275 201.190 ;
        RECT 66.265 201.330 66.555 201.375 ;
        RECT 69.010 201.330 69.330 201.390 ;
        RECT 66.265 201.190 69.330 201.330 ;
        RECT 66.265 201.145 66.555 201.190 ;
        RECT 69.010 201.130 69.330 201.190 ;
        RECT 14.660 200.170 127.820 200.650 ;
        RECT 62.125 199.970 62.415 200.015 ;
        RECT 62.570 199.970 62.890 200.030 ;
        RECT 62.125 199.830 62.890 199.970 ;
        RECT 62.125 199.785 62.415 199.830 ;
        RECT 62.570 199.770 62.890 199.830 ;
        RECT 70.325 199.630 70.615 199.675 ;
        RECT 70.850 199.630 71.170 199.690 ;
        RECT 64.500 199.490 70.160 199.630 ;
        RECT 64.500 199.335 64.640 199.490 ;
        RECT 62.585 199.290 62.875 199.335 ;
        RECT 64.425 199.290 64.715 199.335 ;
        RECT 62.585 199.150 64.715 199.290 ;
        RECT 62.585 199.105 62.875 199.150 ;
        RECT 64.425 199.105 64.715 199.150 ;
        RECT 68.565 199.290 68.855 199.335 ;
        RECT 70.020 199.290 70.160 199.490 ;
        RECT 70.325 199.490 71.170 199.630 ;
        RECT 70.325 199.445 70.615 199.490 ;
        RECT 70.850 199.430 71.170 199.490 ;
        RECT 71.310 199.430 71.630 199.690 ;
        RECT 76.485 199.630 76.775 199.675 ;
        RECT 77.290 199.630 77.610 199.690 ;
        RECT 79.725 199.630 80.375 199.675 ;
        RECT 76.485 199.490 80.375 199.630 ;
        RECT 76.485 199.445 77.075 199.490 ;
        RECT 75.910 199.290 76.230 199.350 ;
        RECT 68.565 199.150 69.700 199.290 ;
        RECT 70.020 199.150 76.230 199.290 ;
        RECT 68.565 199.105 68.855 199.150 ;
        RECT 69.560 198.655 69.700 199.150 ;
        RECT 75.910 199.090 76.230 199.150 ;
        RECT 76.785 199.130 77.075 199.445 ;
        RECT 77.290 199.430 77.610 199.490 ;
        RECT 79.725 199.445 80.375 199.490 ;
        RECT 77.865 199.290 78.155 199.335 ;
        RECT 81.445 199.290 81.735 199.335 ;
        RECT 83.280 199.290 83.570 199.335 ;
        RECT 77.865 199.150 83.570 199.290 ;
        RECT 77.865 199.105 78.155 199.150 ;
        RECT 81.445 199.105 81.735 199.150 ;
        RECT 83.280 199.105 83.570 199.150 ;
        RECT 110.425 199.290 110.715 199.335 ;
        RECT 111.790 199.290 112.110 199.350 ;
        RECT 113.185 199.290 113.475 199.335 ;
        RECT 110.425 199.150 113.475 199.290 ;
        RECT 110.425 199.105 110.715 199.150 ;
        RECT 111.790 199.090 112.110 199.150 ;
        RECT 113.185 199.105 113.475 199.150 ;
        RECT 82.350 198.750 82.670 199.010 ;
        RECT 83.745 198.950 84.035 198.995 ;
        RECT 93.850 198.950 94.170 199.010 ;
        RECT 83.745 198.810 94.170 198.950 ;
        RECT 83.745 198.765 84.035 198.810 ;
        RECT 93.850 198.750 94.170 198.810 ;
        RECT 69.485 198.425 69.775 198.655 ;
        RECT 77.865 198.610 78.155 198.655 ;
        RECT 80.985 198.610 81.275 198.655 ;
        RECT 82.875 198.610 83.165 198.655 ;
        RECT 77.865 198.470 83.165 198.610 ;
        RECT 77.865 198.425 78.155 198.470 ;
        RECT 80.985 198.425 81.275 198.470 ;
        RECT 82.875 198.425 83.165 198.470 ;
        RECT 63.950 198.070 64.270 198.330 ;
        RECT 67.170 198.270 67.490 198.330 ;
        RECT 67.645 198.270 67.935 198.315 ;
        RECT 67.170 198.130 67.935 198.270 ;
        RECT 67.170 198.070 67.490 198.130 ;
        RECT 67.645 198.085 67.935 198.130 ;
        RECT 70.390 198.070 70.710 198.330 ;
        RECT 71.770 198.270 72.090 198.330 ;
        RECT 75.005 198.270 75.295 198.315 ;
        RECT 71.770 198.130 75.295 198.270 ;
        RECT 71.770 198.070 72.090 198.130 ;
        RECT 75.005 198.085 75.295 198.130 ;
        RECT 109.950 198.070 110.270 198.330 ;
        RECT 113.645 198.270 113.935 198.315 ;
        RECT 115.470 198.270 115.790 198.330 ;
        RECT 113.645 198.130 115.790 198.270 ;
        RECT 113.645 198.085 113.935 198.130 ;
        RECT 115.470 198.070 115.790 198.130 ;
        RECT 14.660 197.450 127.820 197.930 ;
        RECT 64.410 197.250 64.730 197.310 ;
        RECT 64.410 197.110 71.080 197.250 ;
        RECT 64.410 197.050 64.730 197.110 ;
        RECT 62.685 196.910 62.975 196.955 ;
        RECT 65.805 196.910 66.095 196.955 ;
        RECT 67.695 196.910 67.985 196.955 ;
        RECT 62.685 196.770 67.985 196.910 ;
        RECT 62.685 196.725 62.975 196.770 ;
        RECT 65.805 196.725 66.095 196.770 ;
        RECT 67.695 196.725 67.985 196.770 ;
        RECT 69.010 196.710 69.330 196.970 ;
        RECT 67.170 196.370 67.490 196.630 ;
        RECT 68.550 196.370 68.870 196.630 ;
        RECT 70.390 196.370 70.710 196.630 ;
        RECT 43.250 196.030 43.570 196.290 ;
        RECT 70.940 196.275 71.080 197.110 ;
        RECT 77.290 197.050 77.610 197.310 ;
        RECT 80.525 197.250 80.815 197.295 ;
        RECT 82.350 197.250 82.670 197.310 ;
        RECT 80.525 197.110 82.670 197.250 ;
        RECT 80.525 197.065 80.815 197.110 ;
        RECT 82.350 197.050 82.670 197.110 ;
        RECT 89.220 196.910 89.510 196.955 ;
        RECT 92.000 196.910 92.290 196.955 ;
        RECT 93.860 196.910 94.150 196.955 ;
        RECT 89.220 196.770 94.150 196.910 ;
        RECT 89.220 196.725 89.510 196.770 ;
        RECT 92.000 196.725 92.290 196.770 ;
        RECT 93.860 196.725 94.150 196.770 ;
        RECT 109.145 196.910 109.435 196.955 ;
        RECT 112.265 196.910 112.555 196.955 ;
        RECT 114.155 196.910 114.445 196.955 ;
        RECT 109.145 196.770 114.445 196.910 ;
        RECT 109.145 196.725 109.435 196.770 ;
        RECT 112.265 196.725 112.555 196.770 ;
        RECT 114.155 196.725 114.445 196.770 ;
        RECT 118.345 196.910 118.635 196.955 ;
        RECT 121.465 196.910 121.755 196.955 ;
        RECT 123.355 196.910 123.645 196.955 ;
        RECT 118.345 196.770 123.645 196.910 ;
        RECT 118.345 196.725 118.635 196.770 ;
        RECT 121.465 196.725 121.755 196.770 ;
        RECT 123.355 196.725 123.645 196.770 ;
        RECT 76.370 196.570 76.690 196.630 ;
        RECT 78.685 196.570 78.975 196.615 ;
        RECT 76.370 196.430 78.975 196.570 ;
        RECT 76.370 196.370 76.690 196.430 ;
        RECT 78.685 196.385 78.975 196.430 ;
        RECT 91.550 196.570 91.870 196.630 ;
        RECT 92.485 196.570 92.775 196.615 ;
        RECT 91.550 196.430 92.775 196.570 ;
        RECT 91.550 196.370 91.870 196.430 ;
        RECT 92.485 196.385 92.775 196.430 ;
        RECT 111.330 196.570 111.650 196.630 ;
        RECT 115.485 196.570 115.775 196.615 ;
        RECT 111.330 196.430 115.775 196.570 ;
        RECT 111.330 196.370 111.650 196.430 ;
        RECT 115.485 196.385 115.775 196.430 ;
        RECT 116.390 196.570 116.710 196.630 ;
        RECT 122.845 196.570 123.135 196.615 ;
        RECT 116.390 196.430 123.135 196.570 ;
        RECT 116.390 196.370 116.710 196.430 ;
        RECT 122.845 196.385 123.135 196.430 ;
        RECT 61.605 195.935 61.895 196.250 ;
        RECT 62.685 196.230 62.975 196.275 ;
        RECT 66.265 196.230 66.555 196.275 ;
        RECT 68.100 196.230 68.390 196.275 ;
        RECT 62.685 196.090 68.390 196.230 ;
        RECT 62.685 196.045 62.975 196.090 ;
        RECT 66.265 196.045 66.555 196.090 ;
        RECT 68.100 196.045 68.390 196.090 ;
        RECT 70.865 196.045 71.155 196.275 ;
        RECT 75.910 196.230 76.230 196.290 ;
        RECT 76.845 196.230 77.135 196.275 ;
        RECT 75.910 196.090 77.135 196.230 ;
        RECT 75.910 196.030 76.230 196.090 ;
        RECT 76.845 196.045 77.135 196.090 ;
        RECT 79.145 196.045 79.435 196.275 ;
        RECT 89.220 196.230 89.510 196.275 ;
        RECT 93.850 196.230 94.170 196.290 ;
        RECT 94.325 196.230 94.615 196.275 ;
        RECT 89.220 196.090 91.755 196.230 ;
        RECT 89.220 196.045 89.510 196.090 ;
        RECT 58.445 195.705 58.735 195.935 ;
        RECT 61.305 195.890 61.895 195.935 ;
        RECT 63.950 195.890 64.270 195.950 ;
        RECT 64.545 195.890 65.195 195.935 ;
        RECT 61.305 195.750 65.195 195.890 ;
        RECT 61.305 195.705 61.595 195.750 ;
        RECT 42.805 195.550 43.095 195.595 ;
        RECT 44.170 195.550 44.490 195.610 ;
        RECT 42.805 195.410 44.490 195.550 ;
        RECT 58.520 195.550 58.660 195.705 ;
        RECT 63.950 195.690 64.270 195.750 ;
        RECT 64.545 195.705 65.195 195.750 ;
        RECT 73.610 195.890 73.930 195.950 ;
        RECT 79.220 195.890 79.360 196.045 ;
        RECT 73.610 195.750 79.360 195.890 ;
        RECT 86.490 195.890 86.810 195.950 ;
        RECT 91.540 195.935 91.755 196.090 ;
        RECT 93.850 196.090 94.615 196.230 ;
        RECT 93.850 196.030 94.170 196.090 ;
        RECT 94.325 196.045 94.615 196.090 ;
        RECT 100.290 196.030 100.610 196.290 ;
        RECT 108.065 195.935 108.355 196.250 ;
        RECT 109.145 196.230 109.435 196.275 ;
        RECT 112.725 196.230 113.015 196.275 ;
        RECT 114.560 196.230 114.850 196.275 ;
        RECT 109.145 196.090 114.850 196.230 ;
        RECT 109.145 196.045 109.435 196.090 ;
        RECT 112.725 196.045 113.015 196.090 ;
        RECT 114.560 196.045 114.850 196.090 ;
        RECT 115.025 196.045 115.315 196.275 ;
        RECT 87.360 195.890 87.650 195.935 ;
        RECT 90.620 195.890 90.910 195.935 ;
        RECT 86.490 195.750 90.910 195.890 ;
        RECT 73.610 195.690 73.930 195.750 ;
        RECT 86.490 195.690 86.810 195.750 ;
        RECT 87.360 195.705 87.650 195.750 ;
        RECT 90.620 195.705 90.910 195.750 ;
        RECT 91.540 195.890 91.830 195.935 ;
        RECT 93.400 195.890 93.690 195.935 ;
        RECT 91.540 195.750 93.690 195.890 ;
        RECT 91.540 195.705 91.830 195.750 ;
        RECT 93.400 195.705 93.690 195.750 ;
        RECT 107.765 195.890 108.355 195.935 ;
        RECT 109.950 195.890 110.270 195.950 ;
        RECT 111.005 195.890 111.655 195.935 ;
        RECT 107.765 195.750 111.655 195.890 ;
        RECT 107.765 195.705 108.055 195.750 ;
        RECT 109.950 195.690 110.270 195.750 ;
        RECT 111.005 195.705 111.655 195.750 ;
        RECT 112.250 195.890 112.570 195.950 ;
        RECT 113.645 195.890 113.935 195.935 ;
        RECT 112.250 195.750 113.935 195.890 ;
        RECT 112.250 195.690 112.570 195.750 ;
        RECT 113.645 195.705 113.935 195.750 ;
        RECT 67.630 195.550 67.950 195.610 ;
        RECT 58.520 195.410 67.950 195.550 ;
        RECT 42.805 195.365 43.095 195.410 ;
        RECT 44.170 195.350 44.490 195.410 ;
        RECT 67.630 195.350 67.950 195.410 ;
        RECT 71.310 195.550 71.630 195.610 ;
        RECT 74.990 195.550 75.310 195.610 ;
        RECT 71.310 195.410 75.310 195.550 ;
        RECT 71.310 195.350 71.630 195.410 ;
        RECT 74.990 195.350 75.310 195.410 ;
        RECT 85.355 195.550 85.645 195.595 ;
        RECT 86.030 195.550 86.350 195.610 ;
        RECT 85.355 195.410 86.350 195.550 ;
        RECT 85.355 195.365 85.645 195.410 ;
        RECT 86.030 195.350 86.350 195.410 ;
        RECT 101.225 195.550 101.515 195.595 ;
        RECT 102.590 195.550 102.910 195.610 ;
        RECT 101.225 195.410 102.910 195.550 ;
        RECT 101.225 195.365 101.515 195.410 ;
        RECT 102.590 195.350 102.910 195.410 ;
        RECT 106.270 195.350 106.590 195.610 ;
        RECT 115.100 195.550 115.240 196.045 ;
        RECT 115.470 195.890 115.790 195.950 ;
        RECT 117.265 195.935 117.555 196.250 ;
        RECT 118.345 196.230 118.635 196.275 ;
        RECT 121.925 196.230 122.215 196.275 ;
        RECT 123.760 196.230 124.050 196.275 ;
        RECT 118.345 196.090 124.050 196.230 ;
        RECT 118.345 196.045 118.635 196.090 ;
        RECT 121.925 196.045 122.215 196.090 ;
        RECT 123.760 196.045 124.050 196.090 ;
        RECT 124.225 196.045 124.515 196.275 ;
        RECT 116.965 195.890 117.555 195.935 ;
        RECT 120.205 195.890 120.855 195.935 ;
        RECT 115.470 195.750 120.855 195.890 ;
        RECT 115.470 195.690 115.790 195.750 ;
        RECT 116.965 195.705 117.255 195.750 ;
        RECT 120.205 195.705 120.855 195.750 ;
        RECT 124.300 195.610 124.440 196.045 ;
        RECT 124.210 195.550 124.530 195.610 ;
        RECT 115.100 195.410 124.530 195.550 ;
        RECT 124.210 195.350 124.530 195.410 ;
        RECT 14.660 194.730 127.820 195.210 ;
        RECT 43.250 194.530 43.570 194.590 ;
        RECT 43.250 194.390 45.780 194.530 ;
        RECT 43.250 194.330 43.570 194.390 ;
        RECT 41.405 194.190 42.055 194.235 ;
        RECT 44.170 194.190 44.490 194.250 ;
        RECT 45.005 194.190 45.295 194.235 ;
        RECT 41.405 194.050 45.295 194.190 ;
        RECT 41.405 194.005 42.055 194.050 ;
        RECT 44.170 193.990 44.490 194.050 ;
        RECT 44.705 194.005 45.295 194.050 ;
        RECT 38.210 193.850 38.500 193.895 ;
        RECT 40.045 193.850 40.335 193.895 ;
        RECT 43.625 193.850 43.915 193.895 ;
        RECT 38.210 193.710 43.915 193.850 ;
        RECT 38.210 193.665 38.500 193.710 ;
        RECT 40.045 193.665 40.335 193.710 ;
        RECT 43.625 193.665 43.915 193.710 ;
        RECT 44.705 193.690 44.995 194.005 ;
        RECT 45.640 193.910 45.780 194.390 ;
        RECT 64.960 194.390 69.700 194.530 ;
        RECT 48.325 194.190 48.615 194.235 ;
        RECT 50.725 194.190 51.015 194.235 ;
        RECT 53.965 194.190 54.615 194.235 ;
        RECT 48.325 194.050 54.615 194.190 ;
        RECT 48.325 194.005 48.615 194.050 ;
        RECT 50.725 194.005 51.315 194.050 ;
        RECT 53.965 194.005 54.615 194.050 ;
        RECT 56.130 194.190 56.450 194.250 ;
        RECT 56.605 194.190 56.895 194.235 ;
        RECT 56.130 194.050 56.895 194.190 ;
        RECT 45.550 193.850 45.870 193.910 ;
        RECT 47.865 193.850 48.155 193.895 ;
        RECT 45.550 193.710 48.155 193.850 ;
        RECT 45.550 193.650 45.870 193.710 ;
        RECT 47.865 193.665 48.155 193.710 ;
        RECT 51.025 193.690 51.315 194.005 ;
        RECT 56.130 193.990 56.450 194.050 ;
        RECT 56.605 194.005 56.895 194.050 ;
        RECT 64.960 193.895 65.100 194.390 ;
        RECT 66.800 194.050 69.240 194.190 ;
        RECT 66.800 193.895 66.940 194.050 ;
        RECT 52.105 193.850 52.395 193.895 ;
        RECT 55.685 193.850 55.975 193.895 ;
        RECT 57.520 193.850 57.810 193.895 ;
        RECT 52.105 193.710 57.810 193.850 ;
        RECT 52.105 193.665 52.395 193.710 ;
        RECT 55.685 193.665 55.975 193.710 ;
        RECT 57.520 193.665 57.810 193.710 ;
        RECT 64.885 193.665 65.175 193.895 ;
        RECT 66.725 193.665 67.015 193.895 ;
        RECT 67.630 193.850 67.950 193.910 ;
        RECT 68.565 193.850 68.855 193.895 ;
        RECT 67.630 193.710 68.855 193.850 ;
        RECT 67.630 193.650 67.950 193.710 ;
        RECT 68.565 193.665 68.855 193.710 ;
        RECT 69.100 193.570 69.240 194.050 ;
        RECT 69.560 193.895 69.700 194.390 ;
        RECT 70.850 194.330 71.170 194.590 ;
        RECT 71.310 194.330 71.630 194.590 ;
        RECT 73.610 194.530 73.930 194.590 ;
        RECT 71.860 194.390 73.930 194.530 ;
        RECT 69.485 193.665 69.775 193.895 ;
        RECT 69.930 193.850 70.250 193.910 ;
        RECT 71.860 193.850 72.000 194.390 ;
        RECT 73.610 194.330 73.930 194.390 ;
        RECT 77.305 194.345 77.595 194.575 ;
        RECT 74.990 194.235 75.310 194.250 ;
        RECT 74.990 194.005 75.595 194.235 ;
        RECT 76.370 194.190 76.690 194.250 ;
        RECT 77.380 194.190 77.520 194.345 ;
        RECT 91.550 194.330 91.870 194.590 ;
        RECT 95.245 194.530 95.535 194.575 ;
        RECT 95.245 194.390 106.960 194.530 ;
        RECT 95.245 194.345 95.535 194.390 ;
        RECT 106.820 194.250 106.960 194.390 ;
        RECT 112.250 194.330 112.570 194.590 ;
        RECT 116.390 194.330 116.710 194.590 ;
        RECT 76.370 194.050 77.520 194.190 ;
        RECT 86.505 194.190 86.795 194.235 ;
        RECT 86.950 194.190 87.270 194.250 ;
        RECT 86.505 194.050 87.270 194.190 ;
        RECT 74.990 193.990 75.310 194.005 ;
        RECT 76.370 193.990 76.690 194.050 ;
        RECT 86.505 194.005 86.795 194.050 ;
        RECT 86.950 193.990 87.270 194.050 ;
        RECT 94.325 194.190 94.615 194.235 ;
        RECT 96.725 194.190 97.015 194.235 ;
        RECT 99.965 194.190 100.615 194.235 ;
        RECT 94.325 194.050 100.615 194.190 ;
        RECT 94.325 194.005 94.615 194.050 ;
        RECT 96.725 194.005 97.315 194.050 ;
        RECT 99.965 194.005 100.615 194.050 ;
        RECT 74.085 193.850 74.375 193.895 ;
        RECT 69.930 193.710 72.000 193.850 ;
        RECT 73.240 193.710 74.375 193.850 ;
        RECT 24.850 193.510 25.170 193.570 ;
        RECT 37.745 193.510 38.035 193.555 ;
        RECT 24.850 193.370 38.035 193.510 ;
        RECT 24.850 193.310 25.170 193.370 ;
        RECT 37.745 193.325 38.035 193.370 ;
        RECT 39.110 193.310 39.430 193.570 ;
        RECT 57.970 193.510 58.290 193.570 ;
        RECT 68.090 193.510 68.410 193.570 ;
        RECT 57.970 193.370 68.410 193.510 ;
        RECT 57.970 193.310 58.290 193.370 ;
        RECT 68.090 193.310 68.410 193.370 ;
        RECT 69.010 193.310 69.330 193.570 ;
        RECT 69.560 193.510 69.700 193.665 ;
        RECT 69.930 193.650 70.250 193.710 ;
        RECT 72.230 193.510 72.550 193.570 ;
        RECT 69.560 193.370 72.550 193.510 ;
        RECT 72.230 193.310 72.550 193.370 ;
        RECT 72.705 193.325 72.995 193.555 ;
        RECT 38.615 193.170 38.905 193.215 ;
        RECT 40.505 193.170 40.795 193.215 ;
        RECT 43.625 193.170 43.915 193.215 ;
        RECT 38.615 193.030 43.915 193.170 ;
        RECT 38.615 192.985 38.905 193.030 ;
        RECT 40.505 192.985 40.795 193.030 ;
        RECT 43.625 192.985 43.915 193.030 ;
        RECT 52.105 193.170 52.395 193.215 ;
        RECT 55.225 193.170 55.515 193.215 ;
        RECT 57.115 193.170 57.405 193.215 ;
        RECT 52.105 193.030 57.405 193.170 ;
        RECT 52.105 192.985 52.395 193.030 ;
        RECT 55.225 192.985 55.515 193.030 ;
        RECT 57.115 192.985 57.405 193.030 ;
        RECT 67.645 193.170 67.935 193.215 ;
        RECT 72.780 193.170 72.920 193.325 ;
        RECT 67.645 193.030 72.920 193.170 ;
        RECT 67.645 192.985 67.935 193.030 ;
        RECT 42.790 192.830 43.110 192.890 ;
        RECT 46.485 192.830 46.775 192.875 ;
        RECT 42.790 192.690 46.775 192.830 ;
        RECT 42.790 192.630 43.110 192.690 ;
        RECT 46.485 192.645 46.775 192.690 ;
        RECT 49.245 192.830 49.535 192.875 ;
        RECT 50.150 192.830 50.470 192.890 ;
        RECT 49.245 192.690 50.470 192.830 ;
        RECT 49.245 192.645 49.535 192.690 ;
        RECT 50.150 192.630 50.470 192.690 ;
        RECT 64.410 192.830 64.730 192.890 ;
        RECT 65.345 192.830 65.635 192.875 ;
        RECT 67.170 192.830 67.490 192.890 ;
        RECT 64.410 192.690 67.490 192.830 ;
        RECT 64.410 192.630 64.730 192.690 ;
        RECT 65.345 192.645 65.635 192.690 ;
        RECT 67.170 192.630 67.490 192.690 ;
        RECT 68.090 192.830 68.410 192.890 ;
        RECT 70.850 192.830 71.170 192.890 ;
        RECT 73.240 192.830 73.380 193.710 ;
        RECT 74.085 193.665 74.375 193.710 ;
        RECT 76.830 193.650 77.150 193.910 ;
        RECT 77.750 193.650 78.070 193.910 ;
        RECT 90.645 193.850 90.935 193.895 ;
        RECT 88.420 193.710 90.935 193.850 ;
        RECT 85.110 193.310 85.430 193.570 ;
        RECT 86.030 193.310 86.350 193.570 ;
        RECT 88.420 193.215 88.560 193.710 ;
        RECT 90.645 193.665 90.935 193.710 ;
        RECT 93.865 193.665 94.155 193.895 ;
        RECT 97.025 193.690 97.315 194.005 ;
        RECT 102.590 193.990 102.910 194.250 ;
        RECT 106.730 194.190 107.050 194.250 ;
        RECT 108.585 194.190 108.875 194.235 ;
        RECT 106.730 194.050 108.875 194.190 ;
        RECT 106.730 193.990 107.050 194.050 ;
        RECT 108.585 194.005 108.875 194.050 ;
        RECT 98.105 193.850 98.395 193.895 ;
        RECT 101.685 193.850 101.975 193.895 ;
        RECT 103.520 193.850 103.810 193.895 ;
        RECT 98.105 193.710 103.810 193.850 ;
        RECT 98.105 193.665 98.395 193.710 ;
        RECT 101.685 193.665 101.975 193.710 ;
        RECT 103.520 193.665 103.810 193.710 ;
        RECT 106.270 193.850 106.590 193.910 ;
        RECT 111.345 193.850 111.635 193.895 ;
        RECT 106.270 193.710 108.340 193.850 ;
        RECT 88.345 192.985 88.635 193.215 ;
        RECT 68.090 192.690 73.380 192.830 ;
        RECT 68.090 192.630 68.410 192.690 ;
        RECT 70.850 192.630 71.170 192.690 ;
        RECT 73.610 192.630 73.930 192.890 ;
        RECT 74.530 192.630 74.850 192.890 ;
        RECT 75.450 192.630 75.770 192.890 ;
        RECT 76.370 192.830 76.690 192.890 ;
        RECT 93.940 192.830 94.080 193.665 ;
        RECT 106.270 193.650 106.590 193.710 ;
        RECT 103.985 193.510 104.275 193.555 ;
        RECT 105.810 193.510 106.130 193.570 ;
        RECT 108.200 193.555 108.340 193.710 ;
        RECT 110.500 193.710 111.635 193.850 ;
        RECT 103.985 193.370 106.130 193.510 ;
        RECT 103.985 193.325 104.275 193.370 ;
        RECT 105.810 193.310 106.130 193.370 ;
        RECT 107.205 193.325 107.495 193.555 ;
        RECT 108.125 193.510 108.415 193.555 ;
        RECT 109.950 193.510 110.270 193.570 ;
        RECT 108.125 193.370 110.270 193.510 ;
        RECT 108.125 193.325 108.415 193.370 ;
        RECT 98.105 193.170 98.395 193.215 ;
        RECT 101.225 193.170 101.515 193.215 ;
        RECT 103.115 193.170 103.405 193.215 ;
        RECT 98.105 193.030 103.405 193.170 ;
        RECT 98.105 192.985 98.395 193.030 ;
        RECT 101.225 192.985 101.515 193.030 ;
        RECT 103.115 192.985 103.405 193.030 ;
        RECT 105.350 193.170 105.670 193.230 ;
        RECT 107.280 193.170 107.420 193.325 ;
        RECT 109.950 193.310 110.270 193.370 ;
        RECT 110.500 193.215 110.640 193.710 ;
        RECT 111.345 193.665 111.635 193.710 ;
        RECT 115.470 193.650 115.790 193.910 ;
        RECT 105.350 193.030 107.420 193.170 ;
        RECT 105.350 192.970 105.670 193.030 ;
        RECT 110.425 192.985 110.715 193.215 ;
        RECT 111.790 192.830 112.110 192.890 ;
        RECT 76.370 192.690 112.110 192.830 ;
        RECT 76.370 192.630 76.690 192.690 ;
        RECT 111.790 192.630 112.110 192.690 ;
        RECT 14.660 192.010 127.820 192.490 ;
        RECT 39.110 191.810 39.430 191.870 ;
        RECT 42.345 191.810 42.635 191.855 ;
        RECT 39.110 191.670 42.635 191.810 ;
        RECT 39.110 191.610 39.430 191.670 ;
        RECT 42.345 191.625 42.635 191.670 ;
        RECT 55.685 191.810 55.975 191.855 ;
        RECT 56.130 191.810 56.450 191.870 ;
        RECT 55.685 191.670 56.450 191.810 ;
        RECT 55.685 191.625 55.975 191.670 ;
        RECT 56.130 191.610 56.450 191.670 ;
        RECT 68.565 191.810 68.855 191.855 ;
        RECT 69.930 191.810 70.250 191.870 ;
        RECT 68.565 191.670 70.250 191.810 ;
        RECT 68.565 191.625 68.855 191.670 ;
        RECT 69.930 191.610 70.250 191.670 ;
        RECT 70.390 191.610 70.710 191.870 ;
        RECT 70.850 191.810 71.170 191.870 ;
        RECT 74.545 191.810 74.835 191.855 ;
        RECT 75.450 191.810 75.770 191.870 ;
        RECT 70.850 191.670 72.000 191.810 ;
        RECT 70.850 191.610 71.170 191.670 ;
        RECT 36.350 191.470 36.670 191.530 ;
        RECT 33.220 191.330 38.420 191.470 ;
        RECT 33.220 191.175 33.360 191.330 ;
        RECT 36.350 191.270 36.670 191.330 ;
        RECT 38.280 191.175 38.420 191.330 ;
        RECT 54.305 191.285 54.595 191.515 ;
        RECT 70.020 191.470 70.160 191.610 ;
        RECT 70.020 191.330 71.080 191.470 ;
        RECT 33.145 190.945 33.435 191.175 ;
        RECT 38.205 190.945 38.495 191.175 ;
        RECT 39.125 191.130 39.415 191.175 ;
        RECT 42.790 191.130 43.110 191.190 ;
        RECT 39.125 190.990 43.110 191.130 ;
        RECT 39.125 190.945 39.415 190.990 ;
        RECT 42.790 190.930 43.110 190.990 ;
        RECT 50.610 191.130 50.930 191.190 ;
        RECT 51.085 191.130 51.375 191.175 ;
        RECT 50.610 190.990 51.375 191.130 ;
        RECT 50.610 190.930 50.930 190.990 ;
        RECT 51.085 190.945 51.375 190.990 ;
        RECT 26.230 190.790 26.550 190.850 ;
        RECT 30.845 190.790 31.135 190.835 ;
        RECT 43.265 190.790 43.555 190.835 ;
        RECT 26.230 190.650 31.135 190.790 ;
        RECT 26.230 190.590 26.550 190.650 ;
        RECT 30.845 190.605 31.135 190.650 ;
        RECT 41.500 190.650 43.555 190.790 ;
        RECT 38.190 190.450 38.510 190.510 ;
        RECT 39.585 190.450 39.875 190.495 ;
        RECT 33.680 190.310 39.875 190.450 ;
        RECT 33.680 190.170 33.820 190.310 ;
        RECT 38.190 190.250 38.510 190.310 ;
        RECT 39.585 190.265 39.875 190.310 ;
        RECT 31.290 189.910 31.610 190.170 ;
        RECT 33.590 189.910 33.910 190.170 ;
        RECT 34.065 190.110 34.355 190.155 ;
        RECT 35.430 190.110 35.750 190.170 ;
        RECT 34.065 189.970 35.750 190.110 ;
        RECT 34.065 189.925 34.355 189.970 ;
        RECT 35.430 189.910 35.750 189.970 ;
        RECT 35.890 189.910 36.210 190.170 ;
        RECT 41.500 190.155 41.640 190.650 ;
        RECT 43.265 190.605 43.555 190.650 ;
        RECT 45.105 190.790 45.395 190.835 ;
        RECT 45.550 190.790 45.870 190.850 ;
        RECT 45.105 190.650 45.870 190.790 ;
        RECT 45.105 190.605 45.395 190.650 ;
        RECT 45.550 190.590 45.870 190.650 ;
        RECT 49.230 190.590 49.550 190.850 ;
        RECT 54.380 190.790 54.520 191.285 ;
        RECT 69.010 191.130 69.330 191.190 ;
        RECT 69.945 191.130 70.235 191.175 ;
        RECT 69.010 190.990 70.235 191.130 ;
        RECT 69.010 190.930 69.330 190.990 ;
        RECT 69.945 190.945 70.235 190.990 ;
        RECT 54.765 190.790 55.055 190.835 ;
        RECT 54.380 190.650 55.055 190.790 ;
        RECT 54.765 190.605 55.055 190.650 ;
        RECT 42.790 190.450 43.110 190.510 ;
        RECT 52.465 190.450 52.755 190.495 ;
        RECT 42.790 190.310 52.755 190.450 ;
        RECT 69.100 190.450 69.240 190.930 ;
        RECT 69.485 190.790 69.775 190.835 ;
        RECT 70.390 190.790 70.710 190.850 ;
        RECT 69.485 190.650 70.710 190.790 ;
        RECT 70.940 190.790 71.080 191.330 ;
        RECT 71.860 190.835 72.000 191.670 ;
        RECT 74.545 191.670 75.770 191.810 ;
        RECT 74.545 191.625 74.835 191.670 ;
        RECT 75.450 191.610 75.770 191.670 ;
        RECT 85.110 191.810 85.430 191.870 ;
        RECT 99.385 191.810 99.675 191.855 ;
        RECT 100.290 191.810 100.610 191.870 ;
        RECT 85.110 191.670 95.920 191.810 ;
        RECT 85.110 191.610 85.430 191.670 ;
        RECT 88.300 191.470 88.590 191.515 ;
        RECT 91.080 191.470 91.370 191.515 ;
        RECT 92.940 191.470 93.230 191.515 ;
        RECT 88.300 191.330 93.230 191.470 ;
        RECT 88.300 191.285 88.590 191.330 ;
        RECT 91.080 191.285 91.370 191.330 ;
        RECT 92.940 191.285 93.230 191.330 ;
        RECT 72.230 191.130 72.550 191.190 ;
        RECT 74.990 191.130 75.310 191.190 ;
        RECT 76.830 191.130 77.150 191.190 ;
        RECT 72.230 190.990 77.150 191.130 ;
        RECT 72.230 190.930 72.550 190.990 ;
        RECT 72.780 190.835 72.920 190.990 ;
        RECT 74.990 190.930 75.310 190.990 ;
        RECT 76.830 190.930 77.150 190.990 ;
        RECT 86.030 191.130 86.350 191.190 ;
        RECT 95.780 191.130 95.920 191.670 ;
        RECT 99.385 191.670 100.610 191.810 ;
        RECT 99.385 191.625 99.675 191.670 ;
        RECT 100.290 191.610 100.610 191.670 ;
        RECT 113.645 191.810 113.935 191.855 ;
        RECT 115.470 191.810 115.790 191.870 ;
        RECT 113.645 191.670 115.790 191.810 ;
        RECT 113.645 191.625 113.935 191.670 ;
        RECT 115.470 191.610 115.790 191.670 ;
        RECT 96.165 191.130 96.455 191.175 ;
        RECT 103.050 191.130 103.370 191.190 ;
        RECT 105.350 191.130 105.670 191.190 ;
        RECT 110.425 191.130 110.715 191.175 ;
        RECT 86.030 190.990 94.540 191.130 ;
        RECT 95.780 190.990 110.715 191.130 ;
        RECT 86.030 190.930 86.350 190.990 ;
        RECT 71.325 190.790 71.615 190.835 ;
        RECT 70.940 190.650 71.615 190.790 ;
        RECT 69.485 190.605 69.775 190.650 ;
        RECT 70.390 190.590 70.710 190.650 ;
        RECT 71.325 190.605 71.615 190.650 ;
        RECT 71.785 190.605 72.075 190.835 ;
        RECT 72.705 190.605 72.995 190.835 ;
        RECT 73.625 190.790 73.915 190.835 ;
        RECT 77.750 190.790 78.070 190.850 ;
        RECT 73.625 190.650 78.070 190.790 ;
        RECT 73.625 190.605 73.915 190.650 ;
        RECT 73.700 190.450 73.840 190.605 ;
        RECT 77.750 190.590 78.070 190.650 ;
        RECT 88.300 190.790 88.590 190.835 ;
        RECT 88.300 190.650 90.835 190.790 ;
        RECT 88.300 190.605 88.590 190.650 ;
        RECT 69.100 190.310 73.840 190.450 ;
        RECT 86.440 190.450 86.730 190.495 ;
        RECT 87.870 190.450 88.190 190.510 ;
        RECT 90.620 190.495 90.835 190.650 ;
        RECT 91.550 190.590 91.870 190.850 ;
        RECT 93.405 190.790 93.695 190.835 ;
        RECT 93.850 190.790 94.170 190.850 ;
        RECT 93.405 190.650 94.170 190.790 ;
        RECT 94.400 190.790 94.540 190.990 ;
        RECT 96.165 190.945 96.455 190.990 ;
        RECT 103.050 190.930 103.370 190.990 ;
        RECT 105.350 190.930 105.670 190.990 ;
        RECT 110.425 190.945 110.715 190.990 ;
        RECT 111.330 190.930 111.650 191.190 ;
        RECT 97.545 190.790 97.835 190.835 ;
        RECT 94.400 190.650 97.835 190.790 ;
        RECT 93.405 190.605 93.695 190.650 ;
        RECT 93.850 190.590 94.170 190.650 ;
        RECT 97.545 190.605 97.835 190.650 ;
        RECT 89.700 190.450 89.990 190.495 ;
        RECT 86.440 190.310 89.990 190.450 ;
        RECT 42.790 190.250 43.110 190.310 ;
        RECT 52.465 190.265 52.755 190.310 ;
        RECT 86.440 190.265 86.730 190.310 ;
        RECT 87.870 190.250 88.190 190.310 ;
        RECT 89.700 190.265 89.990 190.310 ;
        RECT 90.620 190.450 90.910 190.495 ;
        RECT 92.480 190.450 92.770 190.495 ;
        RECT 90.620 190.310 92.770 190.450 ;
        RECT 90.620 190.265 90.910 190.310 ;
        RECT 92.480 190.265 92.770 190.310 ;
        RECT 41.425 189.925 41.715 190.155 ;
        RECT 44.630 189.910 44.950 190.170 ;
        RECT 46.470 190.110 46.790 190.170 ;
        RECT 48.325 190.110 48.615 190.155 ;
        RECT 46.470 189.970 48.615 190.110 ;
        RECT 46.470 189.910 46.790 189.970 ;
        RECT 48.325 189.925 48.615 189.970 ;
        RECT 50.150 190.110 50.470 190.170 ;
        RECT 52.005 190.110 52.295 190.155 ;
        RECT 50.150 189.970 52.295 190.110 ;
        RECT 50.150 189.910 50.470 189.970 ;
        RECT 52.005 189.925 52.295 189.970 ;
        RECT 70.865 190.110 71.155 190.155 ;
        RECT 72.230 190.110 72.550 190.170 ;
        RECT 70.865 189.970 72.550 190.110 ;
        RECT 70.865 189.925 71.155 189.970 ;
        RECT 72.230 189.910 72.550 189.970 ;
        RECT 84.435 190.110 84.725 190.155 ;
        RECT 86.950 190.110 87.270 190.170 ;
        RECT 84.435 189.970 87.270 190.110 ;
        RECT 84.435 189.925 84.725 189.970 ;
        RECT 86.950 189.910 87.270 189.970 ;
        RECT 97.085 190.110 97.375 190.155 ;
        RECT 106.270 190.110 106.590 190.170 ;
        RECT 97.085 189.970 106.590 190.110 ;
        RECT 97.085 189.925 97.375 189.970 ;
        RECT 106.270 189.910 106.590 189.970 ;
        RECT 109.950 190.110 110.270 190.170 ;
        RECT 111.805 190.110 112.095 190.155 ;
        RECT 109.950 189.970 112.095 190.110 ;
        RECT 109.950 189.910 110.270 189.970 ;
        RECT 111.805 189.925 112.095 189.970 ;
        RECT 14.660 189.290 127.820 189.770 ;
        RECT 27.855 189.090 28.145 189.135 ;
        RECT 33.590 189.090 33.910 189.150 ;
        RECT 37.745 189.090 38.035 189.135 ;
        RECT 27.855 188.950 33.910 189.090 ;
        RECT 27.855 188.905 28.145 188.950 ;
        RECT 33.590 188.890 33.910 188.950 ;
        RECT 36.440 188.950 38.035 189.090 ;
        RECT 29.860 188.750 30.150 188.795 ;
        RECT 31.290 188.750 31.610 188.810 ;
        RECT 33.120 188.750 33.410 188.795 ;
        RECT 29.860 188.610 33.410 188.750 ;
        RECT 29.860 188.565 30.150 188.610 ;
        RECT 31.290 188.550 31.610 188.610 ;
        RECT 33.120 188.565 33.410 188.610 ;
        RECT 34.040 188.750 34.330 188.795 ;
        RECT 35.900 188.750 36.190 188.795 ;
        RECT 34.040 188.610 36.190 188.750 ;
        RECT 34.040 188.565 34.330 188.610 ;
        RECT 35.900 188.565 36.190 188.610 ;
        RECT 26.230 188.210 26.550 188.470 ;
        RECT 26.705 188.410 26.995 188.455 ;
        RECT 30.370 188.410 30.690 188.470 ;
        RECT 26.705 188.270 30.690 188.410 ;
        RECT 26.705 188.225 26.995 188.270 ;
        RECT 30.370 188.210 30.690 188.270 ;
        RECT 31.720 188.410 32.010 188.455 ;
        RECT 34.040 188.410 34.255 188.565 ;
        RECT 31.720 188.270 34.255 188.410 ;
        RECT 34.985 188.410 35.275 188.455 ;
        RECT 36.440 188.410 36.580 188.950 ;
        RECT 37.745 188.905 38.035 188.950 ;
        RECT 46.470 189.090 46.790 189.150 ;
        RECT 46.470 188.950 47.620 189.090 ;
        RECT 46.470 188.890 46.790 188.950 ;
        RECT 44.630 188.795 44.950 188.810 ;
        RECT 47.480 188.795 47.620 188.950 ;
        RECT 86.490 188.890 86.810 189.150 ;
        RECT 87.870 188.890 88.190 189.150 ;
        RECT 90.645 189.090 90.935 189.135 ;
        RECT 91.550 189.090 91.870 189.150 ;
        RECT 90.645 188.950 91.870 189.090 ;
        RECT 90.645 188.905 90.935 188.950 ;
        RECT 91.550 188.890 91.870 188.950 ;
        RECT 41.525 188.750 41.815 188.795 ;
        RECT 44.630 188.750 45.415 188.795 ;
        RECT 41.525 188.610 45.415 188.750 ;
        RECT 41.525 188.565 42.115 188.610 ;
        RECT 38.665 188.410 38.955 188.455 ;
        RECT 34.985 188.270 36.580 188.410 ;
        RECT 37.360 188.270 38.955 188.410 ;
        RECT 31.720 188.225 32.010 188.270 ;
        RECT 34.985 188.225 35.275 188.270 ;
        RECT 24.850 188.070 25.170 188.130 ;
        RECT 36.790 188.070 37.080 188.115 ;
        RECT 24.850 187.930 37.080 188.070 ;
        RECT 24.850 187.870 25.170 187.930 ;
        RECT 36.790 187.885 37.080 187.930 ;
        RECT 31.720 187.730 32.010 187.775 ;
        RECT 34.500 187.730 34.790 187.775 ;
        RECT 36.360 187.730 36.650 187.775 ;
        RECT 31.720 187.590 36.650 187.730 ;
        RECT 31.720 187.545 32.010 187.590 ;
        RECT 34.500 187.545 34.790 187.590 ;
        RECT 36.360 187.545 36.650 187.590 ;
        RECT 35.890 187.390 36.210 187.450 ;
        RECT 37.360 187.390 37.500 188.270 ;
        RECT 38.665 188.225 38.955 188.270 ;
        RECT 41.825 188.250 42.115 188.565 ;
        RECT 44.630 188.565 45.415 188.610 ;
        RECT 47.405 188.565 47.695 188.795 ;
        RECT 50.725 188.750 51.015 188.795 ;
        RECT 51.530 188.750 51.850 188.810 ;
        RECT 53.965 188.750 54.615 188.795 ;
        RECT 97.545 188.750 97.835 188.795 ;
        RECT 99.945 188.750 100.235 188.795 ;
        RECT 103.185 188.750 103.835 188.795 ;
        RECT 50.725 188.610 54.615 188.750 ;
        RECT 50.725 188.565 51.315 188.610 ;
        RECT 44.630 188.550 44.950 188.565 ;
        RECT 42.905 188.410 43.195 188.455 ;
        RECT 46.485 188.410 46.775 188.455 ;
        RECT 48.320 188.410 48.610 188.455 ;
        RECT 42.905 188.270 48.610 188.410 ;
        RECT 42.905 188.225 43.195 188.270 ;
        RECT 46.485 188.225 46.775 188.270 ;
        RECT 48.320 188.225 48.610 188.270 ;
        RECT 51.025 188.250 51.315 188.565 ;
        RECT 51.530 188.550 51.850 188.610 ;
        RECT 53.965 188.565 54.615 188.610 ;
        RECT 87.500 188.610 90.860 188.750 ;
        RECT 52.105 188.410 52.395 188.455 ;
        RECT 55.685 188.410 55.975 188.455 ;
        RECT 57.520 188.410 57.810 188.455 ;
        RECT 52.105 188.270 57.810 188.410 ;
        RECT 52.105 188.225 52.395 188.270 ;
        RECT 55.685 188.225 55.975 188.270 ;
        RECT 57.520 188.225 57.810 188.270 ;
        RECT 57.970 188.210 58.290 188.470 ;
        RECT 73.625 188.225 73.915 188.455 ;
        RECT 74.530 188.410 74.850 188.470 ;
        RECT 87.500 188.455 87.640 188.610 ;
        RECT 90.720 188.470 90.860 188.610 ;
        RECT 97.545 188.610 103.835 188.750 ;
        RECT 97.545 188.565 97.835 188.610 ;
        RECT 99.945 188.565 100.535 188.610 ;
        RECT 103.185 188.565 103.835 188.610 ;
        RECT 116.965 188.750 117.255 188.795 ;
        RECT 119.150 188.750 119.470 188.810 ;
        RECT 120.205 188.750 120.855 188.795 ;
        RECT 116.965 188.610 120.855 188.750 ;
        RECT 116.965 188.565 117.555 188.610 ;
        RECT 76.845 188.410 77.135 188.455 ;
        RECT 74.530 188.270 77.135 188.410 ;
        RECT 48.785 188.070 49.075 188.115 ;
        RECT 58.060 188.070 58.200 188.210 ;
        RECT 48.785 187.930 58.200 188.070 ;
        RECT 72.230 188.070 72.550 188.130 ;
        RECT 73.165 188.070 73.455 188.115 ;
        RECT 72.230 187.930 73.455 188.070 ;
        RECT 73.700 188.070 73.840 188.225 ;
        RECT 74.530 188.210 74.850 188.270 ;
        RECT 76.845 188.225 77.135 188.270 ;
        RECT 86.045 188.410 86.335 188.455 ;
        RECT 87.425 188.410 87.715 188.455 ;
        RECT 86.045 188.270 87.715 188.410 ;
        RECT 86.045 188.225 86.335 188.270 ;
        RECT 87.425 188.225 87.715 188.270 ;
        RECT 89.710 188.210 90.030 188.470 ;
        RECT 90.630 188.410 90.950 188.470 ;
        RECT 97.085 188.410 97.375 188.455 ;
        RECT 90.630 188.270 97.375 188.410 ;
        RECT 90.630 188.210 90.950 188.270 ;
        RECT 97.085 188.225 97.375 188.270 ;
        RECT 100.245 188.250 100.535 188.565 ;
        RECT 101.325 188.410 101.615 188.455 ;
        RECT 104.905 188.410 105.195 188.455 ;
        RECT 106.740 188.410 107.030 188.455 ;
        RECT 101.325 188.270 107.030 188.410 ;
        RECT 101.325 188.225 101.615 188.270 ;
        RECT 104.905 188.225 105.195 188.270 ;
        RECT 106.740 188.225 107.030 188.270 ;
        RECT 117.265 188.250 117.555 188.565 ;
        RECT 119.150 188.550 119.470 188.610 ;
        RECT 120.205 188.565 120.855 188.610 ;
        RECT 118.345 188.410 118.635 188.455 ;
        RECT 121.925 188.410 122.215 188.455 ;
        RECT 123.760 188.410 124.050 188.455 ;
        RECT 118.345 188.270 124.050 188.410 ;
        RECT 118.345 188.225 118.635 188.270 ;
        RECT 121.925 188.225 122.215 188.270 ;
        RECT 123.760 188.225 124.050 188.270 ;
        RECT 124.210 188.210 124.530 188.470 ;
        RECT 76.370 188.070 76.690 188.130 ;
        RECT 73.700 187.930 76.690 188.070 ;
        RECT 48.785 187.885 49.075 187.930 ;
        RECT 72.230 187.870 72.550 187.930 ;
        RECT 73.165 187.885 73.455 187.930 ;
        RECT 76.370 187.870 76.690 187.930 ;
        RECT 105.810 188.070 106.130 188.130 ;
        RECT 107.205 188.070 107.495 188.115 ;
        RECT 105.810 187.930 107.495 188.070 ;
        RECT 105.810 187.870 106.130 187.930 ;
        RECT 107.205 187.885 107.495 187.930 ;
        RECT 112.250 188.070 112.570 188.130 ;
        RECT 115.485 188.070 115.775 188.115 ;
        RECT 112.250 187.930 115.775 188.070 ;
        RECT 112.250 187.870 112.570 187.930 ;
        RECT 115.485 187.885 115.775 187.930 ;
        RECT 42.905 187.730 43.195 187.775 ;
        RECT 46.025 187.730 46.315 187.775 ;
        RECT 47.915 187.730 48.205 187.775 ;
        RECT 42.905 187.590 48.205 187.730 ;
        RECT 42.905 187.545 43.195 187.590 ;
        RECT 46.025 187.545 46.315 187.590 ;
        RECT 47.915 187.545 48.205 187.590 ;
        RECT 52.105 187.730 52.395 187.775 ;
        RECT 55.225 187.730 55.515 187.775 ;
        RECT 57.115 187.730 57.405 187.775 ;
        RECT 52.105 187.590 57.405 187.730 ;
        RECT 52.105 187.545 52.395 187.590 ;
        RECT 55.225 187.545 55.515 187.590 ;
        RECT 57.115 187.545 57.405 187.590 ;
        RECT 101.325 187.730 101.615 187.775 ;
        RECT 104.445 187.730 104.735 187.775 ;
        RECT 106.335 187.730 106.625 187.775 ;
        RECT 101.325 187.590 106.625 187.730 ;
        RECT 101.325 187.545 101.615 187.590 ;
        RECT 104.445 187.545 104.735 187.590 ;
        RECT 106.335 187.545 106.625 187.590 ;
        RECT 118.345 187.730 118.635 187.775 ;
        RECT 121.465 187.730 121.755 187.775 ;
        RECT 123.355 187.730 123.645 187.775 ;
        RECT 118.345 187.590 123.645 187.730 ;
        RECT 118.345 187.545 118.635 187.590 ;
        RECT 121.465 187.545 121.755 187.590 ;
        RECT 123.355 187.545 123.645 187.590 ;
        RECT 35.890 187.250 37.500 187.390 ;
        RECT 35.890 187.190 36.210 187.250 ;
        RECT 40.030 187.190 40.350 187.450 ;
        RECT 48.770 187.390 49.090 187.450 ;
        RECT 49.245 187.390 49.535 187.435 ;
        RECT 48.770 187.250 49.535 187.390 ;
        RECT 48.770 187.190 49.090 187.250 ;
        RECT 49.245 187.205 49.535 187.250 ;
        RECT 55.670 187.390 55.990 187.450 ;
        RECT 56.670 187.390 56.960 187.435 ;
        RECT 55.670 187.250 56.960 187.390 ;
        RECT 55.670 187.190 55.990 187.250 ;
        RECT 56.670 187.205 56.960 187.250 ;
        RECT 74.070 187.390 74.390 187.450 ;
        RECT 75.925 187.390 76.215 187.435 ;
        RECT 74.070 187.250 76.215 187.390 ;
        RECT 74.070 187.190 74.390 187.250 ;
        RECT 75.925 187.205 76.215 187.250 ;
        RECT 98.450 187.190 98.770 187.450 ;
        RECT 105.920 187.390 106.210 187.435 ;
        RECT 106.730 187.390 107.050 187.450 ;
        RECT 105.920 187.250 107.050 187.390 ;
        RECT 105.920 187.205 106.210 187.250 ;
        RECT 106.730 187.190 107.050 187.250 ;
        RECT 120.990 187.390 121.310 187.450 ;
        RECT 122.910 187.390 123.200 187.435 ;
        RECT 120.990 187.250 123.200 187.390 ;
        RECT 120.990 187.190 121.310 187.250 ;
        RECT 122.910 187.205 123.200 187.250 ;
        RECT 14.660 186.570 127.820 187.050 ;
        RECT 49.230 186.370 49.550 186.430 ;
        RECT 49.705 186.370 49.995 186.415 ;
        RECT 49.230 186.230 49.995 186.370 ;
        RECT 49.230 186.170 49.550 186.230 ;
        RECT 49.705 186.185 49.995 186.230 ;
        RECT 51.530 186.370 51.850 186.430 ;
        RECT 52.005 186.370 52.295 186.415 ;
        RECT 51.530 186.230 52.295 186.370 ;
        RECT 51.530 186.170 51.850 186.230 ;
        RECT 52.005 186.185 52.295 186.230 ;
        RECT 55.670 186.370 55.990 186.430 ;
        RECT 56.605 186.370 56.895 186.415 ;
        RECT 55.670 186.230 56.895 186.370 ;
        RECT 55.670 186.170 55.990 186.230 ;
        RECT 56.605 186.185 56.895 186.230 ;
        RECT 89.265 186.370 89.555 186.415 ;
        RECT 89.710 186.370 90.030 186.430 ;
        RECT 89.265 186.230 90.030 186.370 ;
        RECT 89.265 186.185 89.555 186.230 ;
        RECT 89.710 186.170 90.030 186.230 ;
        RECT 106.730 186.170 107.050 186.430 ;
        RECT 119.150 186.370 119.470 186.430 ;
        RECT 120.545 186.370 120.835 186.415 ;
        RECT 119.150 186.230 120.835 186.370 ;
        RECT 119.150 186.170 119.470 186.230 ;
        RECT 120.545 186.185 120.835 186.230 ;
        RECT 120.990 186.370 121.310 186.430 ;
        RECT 122.385 186.370 122.675 186.415 ;
        RECT 120.990 186.230 122.675 186.370 ;
        RECT 120.990 186.170 121.310 186.230 ;
        RECT 122.385 186.185 122.675 186.230 ;
        RECT 25.735 186.030 26.025 186.075 ;
        RECT 27.625 186.030 27.915 186.075 ;
        RECT 30.745 186.030 31.035 186.075 ;
        RECT 69.585 186.030 69.875 186.075 ;
        RECT 72.705 186.030 72.995 186.075 ;
        RECT 74.595 186.030 74.885 186.075 ;
        RECT 25.735 185.890 31.035 186.030 ;
        RECT 25.735 185.845 26.025 185.890 ;
        RECT 27.625 185.845 27.915 185.890 ;
        RECT 30.745 185.845 31.035 185.890 ;
        RECT 47.020 185.890 50.380 186.030 ;
        RECT 24.850 185.490 25.170 185.750 ;
        RECT 47.020 185.735 47.160 185.890 ;
        RECT 46.945 185.505 47.235 185.735 ;
        RECT 50.240 185.690 50.380 185.890 ;
        RECT 69.585 185.890 74.885 186.030 ;
        RECT 69.585 185.845 69.875 185.890 ;
        RECT 72.705 185.845 72.995 185.890 ;
        RECT 74.595 185.845 74.885 185.890 ;
        RECT 106.285 185.845 106.575 186.075 ;
        RECT 113.745 186.030 114.035 186.075 ;
        RECT 116.865 186.030 117.155 186.075 ;
        RECT 118.755 186.030 119.045 186.075 ;
        RECT 113.745 185.890 119.045 186.030 ;
        RECT 113.745 185.845 114.035 185.890 ;
        RECT 116.865 185.845 117.155 185.890 ;
        RECT 118.755 185.845 119.045 185.890 ;
        RECT 50.610 185.690 50.930 185.750 ;
        RECT 50.240 185.550 50.930 185.690 ;
        RECT 50.610 185.490 50.930 185.550 ;
        RECT 51.620 185.550 58.200 185.690 ;
        RECT 25.330 185.350 25.620 185.395 ;
        RECT 27.165 185.350 27.455 185.395 ;
        RECT 30.745 185.350 31.035 185.395 ;
        RECT 25.330 185.210 31.035 185.350 ;
        RECT 25.330 185.165 25.620 185.210 ;
        RECT 27.165 185.165 27.455 185.210 ;
        RECT 30.745 185.165 31.035 185.210 ;
        RECT 26.230 184.810 26.550 185.070 ;
        RECT 28.525 185.010 29.175 185.055 ;
        RECT 29.910 185.010 30.230 185.070 ;
        RECT 31.825 185.055 32.115 185.370 ;
        RECT 46.010 185.350 46.330 185.410 ;
        RECT 47.865 185.350 48.155 185.395 ;
        RECT 49.230 185.350 49.550 185.410 ;
        RECT 51.620 185.395 51.760 185.550 ;
        RECT 51.545 185.350 51.835 185.395 ;
        RECT 46.010 185.210 49.550 185.350 ;
        RECT 46.010 185.150 46.330 185.210 ;
        RECT 47.865 185.165 48.155 185.210 ;
        RECT 49.230 185.150 49.550 185.210 ;
        RECT 50.470 185.210 51.835 185.350 ;
        RECT 31.825 185.010 32.415 185.055 ;
        RECT 28.525 184.870 32.415 185.010 ;
        RECT 28.525 184.825 29.175 184.870 ;
        RECT 29.910 184.810 30.230 184.870 ;
        RECT 32.125 184.825 32.415 184.870 ;
        RECT 45.550 185.010 45.870 185.070 ;
        RECT 50.470 185.010 50.610 185.210 ;
        RECT 51.545 185.165 51.835 185.210 ;
        RECT 53.370 185.350 53.690 185.410 ;
        RECT 58.060 185.395 58.200 185.550 ;
        RECT 74.070 185.490 74.390 185.750 ;
        RECT 85.110 185.690 85.430 185.750 ;
        RECT 86.045 185.690 86.335 185.735 ;
        RECT 85.110 185.550 86.335 185.690 ;
        RECT 85.110 185.490 85.430 185.550 ;
        RECT 86.045 185.505 86.335 185.550 ;
        RECT 103.050 185.490 103.370 185.750 ;
        RECT 55.685 185.350 55.975 185.395 ;
        RECT 53.370 185.210 55.975 185.350 ;
        RECT 53.370 185.150 53.690 185.210 ;
        RECT 55.685 185.165 55.975 185.210 ;
        RECT 57.985 185.350 58.275 185.395 ;
        RECT 63.950 185.350 64.270 185.410 ;
        RECT 57.985 185.210 64.270 185.350 ;
        RECT 57.985 185.165 58.275 185.210 ;
        RECT 63.950 185.150 64.270 185.210 ;
        RECT 68.505 185.055 68.795 185.370 ;
        RECT 69.585 185.350 69.875 185.395 ;
        RECT 73.165 185.350 73.455 185.395 ;
        RECT 75.000 185.350 75.290 185.395 ;
        RECT 69.585 185.210 75.290 185.350 ;
        RECT 69.585 185.165 69.875 185.210 ;
        RECT 73.165 185.165 73.455 185.210 ;
        RECT 75.000 185.165 75.290 185.210 ;
        RECT 75.450 185.150 75.770 185.410 ;
        RECT 76.370 185.350 76.690 185.410 ;
        RECT 77.305 185.350 77.595 185.395 ;
        RECT 76.370 185.210 77.595 185.350 ;
        RECT 76.370 185.150 76.690 185.210 ;
        RECT 77.305 185.165 77.595 185.210 ;
        RECT 98.450 185.350 98.770 185.410 ;
        RECT 103.985 185.350 104.275 185.395 ;
        RECT 98.450 185.210 104.275 185.350 ;
        RECT 106.360 185.350 106.500 185.845 ;
        RECT 111.790 185.690 112.110 185.750 ;
        RECT 113.170 185.690 113.490 185.750 ;
        RECT 109.580 185.550 113.490 185.690 ;
        RECT 109.580 185.395 109.720 185.550 ;
        RECT 111.790 185.490 112.110 185.550 ;
        RECT 113.170 185.490 113.490 185.550 ;
        RECT 119.625 185.690 119.915 185.735 ;
        RECT 124.210 185.690 124.530 185.750 ;
        RECT 119.625 185.550 124.530 185.690 ;
        RECT 119.625 185.505 119.915 185.550 ;
        RECT 124.210 185.490 124.530 185.550 ;
        RECT 107.665 185.350 107.955 185.395 ;
        RECT 106.360 185.210 107.955 185.350 ;
        RECT 98.450 185.150 98.770 185.210 ;
        RECT 103.985 185.165 104.275 185.210 ;
        RECT 107.665 185.165 107.955 185.210 ;
        RECT 109.505 185.165 109.795 185.395 ;
        RECT 45.550 184.870 50.610 185.010 ;
        RECT 68.205 185.010 68.795 185.055 ;
        RECT 71.445 185.010 72.095 185.055 ;
        RECT 76.845 185.010 77.135 185.055 ;
        RECT 68.205 184.870 77.135 185.010 ;
        RECT 45.550 184.810 45.870 184.870 ;
        RECT 68.205 184.825 68.495 184.870 ;
        RECT 71.445 184.825 72.095 184.870 ;
        RECT 76.845 184.825 77.135 184.870 ;
        RECT 84.650 185.010 84.970 185.070 ;
        RECT 112.665 185.055 112.955 185.370 ;
        RECT 113.745 185.350 114.035 185.395 ;
        RECT 117.325 185.350 117.615 185.395 ;
        RECT 119.160 185.350 119.450 185.395 ;
        RECT 113.745 185.210 119.450 185.350 ;
        RECT 113.745 185.165 114.035 185.210 ;
        RECT 117.325 185.165 117.615 185.210 ;
        RECT 119.160 185.165 119.450 185.210 ;
        RECT 120.085 185.165 120.375 185.395 ;
        RECT 120.530 185.350 120.850 185.410 ;
        RECT 121.465 185.350 121.755 185.395 ;
        RECT 120.530 185.210 121.755 185.350 ;
        RECT 87.425 185.010 87.715 185.055 ;
        RECT 84.650 184.870 87.715 185.010 ;
        RECT 84.650 184.810 84.970 184.870 ;
        RECT 87.425 184.825 87.715 184.870 ;
        RECT 109.965 185.010 110.255 185.055 ;
        RECT 112.365 185.010 112.955 185.055 ;
        RECT 115.605 185.010 116.255 185.055 ;
        RECT 109.965 184.870 116.255 185.010 ;
        RECT 109.965 184.825 110.255 184.870 ;
        RECT 112.365 184.825 112.655 184.870 ;
        RECT 115.605 184.825 116.255 184.870 ;
        RECT 118.230 184.810 118.550 185.070 ;
        RECT 33.605 184.670 33.895 184.715 ;
        RECT 34.050 184.670 34.370 184.730 ;
        RECT 35.430 184.670 35.750 184.730 ;
        RECT 33.605 184.530 35.750 184.670 ;
        RECT 33.605 184.485 33.895 184.530 ;
        RECT 34.050 184.470 34.370 184.530 ;
        RECT 35.430 184.470 35.750 184.530 ;
        RECT 46.470 184.670 46.790 184.730 ;
        RECT 47.405 184.670 47.695 184.715 ;
        RECT 46.470 184.530 47.695 184.670 ;
        RECT 46.470 184.470 46.790 184.530 ;
        RECT 47.405 184.485 47.695 184.530 ;
        RECT 57.510 184.470 57.830 184.730 ;
        RECT 66.725 184.670 67.015 184.715 ;
        RECT 67.630 184.670 67.950 184.730 ;
        RECT 66.725 184.530 67.950 184.670 ;
        RECT 66.725 184.485 67.015 184.530 ;
        RECT 67.630 184.470 67.950 184.530 ;
        RECT 86.950 184.470 87.270 184.730 ;
        RECT 101.210 184.670 101.530 184.730 ;
        RECT 104.445 184.670 104.735 184.715 ;
        RECT 110.885 184.670 111.175 184.715 ;
        RECT 111.790 184.670 112.110 184.730 ;
        RECT 101.210 184.530 112.110 184.670 ;
        RECT 101.210 184.470 101.530 184.530 ;
        RECT 104.445 184.485 104.735 184.530 ;
        RECT 110.885 184.485 111.175 184.530 ;
        RECT 111.790 184.470 112.110 184.530 ;
        RECT 113.170 184.670 113.490 184.730 ;
        RECT 120.160 184.670 120.300 185.165 ;
        RECT 120.530 185.150 120.850 185.210 ;
        RECT 121.465 185.165 121.755 185.210 ;
        RECT 113.170 184.530 120.300 184.670 ;
        RECT 113.170 184.470 113.490 184.530 ;
        RECT 14.660 183.850 127.820 184.330 ;
        RECT 26.230 183.650 26.550 183.710 ;
        RECT 27.625 183.650 27.915 183.695 ;
        RECT 26.230 183.510 27.915 183.650 ;
        RECT 26.230 183.450 26.550 183.510 ;
        RECT 27.625 183.465 27.915 183.510 ;
        RECT 46.930 183.650 47.250 183.710 ;
        RECT 49.230 183.650 49.550 183.710 ;
        RECT 51.085 183.650 51.375 183.695 ;
        RECT 46.930 183.510 49.000 183.650 ;
        RECT 46.930 183.450 47.250 183.510 ;
        RECT 40.030 183.310 40.350 183.370 ;
        RECT 43.725 183.310 44.015 183.355 ;
        RECT 46.470 183.310 46.790 183.370 ;
        RECT 40.030 183.170 48.540 183.310 ;
        RECT 40.030 183.110 40.350 183.170 ;
        RECT 43.725 183.125 44.015 183.170 ;
        RECT 46.470 183.110 46.790 183.170 ;
        RECT 28.545 182.970 28.835 183.015 ;
        RECT 28.545 182.830 29.220 182.970 ;
        RECT 28.545 182.785 28.835 182.830 ;
        RECT 29.080 182.335 29.220 182.830 ;
        RECT 30.830 182.770 31.150 183.030 ;
        RECT 31.305 182.970 31.595 183.015 ;
        RECT 34.050 182.970 34.370 183.030 ;
        RECT 45.090 182.970 45.410 183.030 ;
        RECT 48.400 183.015 48.540 183.170 ;
        RECT 47.405 182.970 47.695 183.015 ;
        RECT 31.305 182.830 34.370 182.970 ;
        RECT 31.305 182.785 31.595 182.830 ;
        RECT 34.050 182.770 34.370 182.830 ;
        RECT 42.420 182.830 44.400 182.970 ;
        RECT 32.225 182.630 32.515 182.675 ;
        RECT 35.430 182.630 35.750 182.690 ;
        RECT 36.350 182.630 36.670 182.690 ;
        RECT 42.420 182.675 42.560 182.830 ;
        RECT 42.345 182.630 42.635 182.675 ;
        RECT 32.225 182.490 42.635 182.630 ;
        RECT 32.225 182.445 32.515 182.490 ;
        RECT 35.430 182.430 35.750 182.490 ;
        RECT 36.350 182.430 36.670 182.490 ;
        RECT 42.345 182.445 42.635 182.490 ;
        RECT 43.265 182.630 43.555 182.675 ;
        RECT 43.710 182.630 44.030 182.690 ;
        RECT 43.265 182.490 44.030 182.630 ;
        RECT 44.260 182.630 44.400 182.830 ;
        RECT 45.090 182.830 47.695 182.970 ;
        RECT 45.090 182.770 45.410 182.830 ;
        RECT 47.405 182.785 47.695 182.830 ;
        RECT 47.865 182.785 48.155 183.015 ;
        RECT 48.325 182.785 48.615 183.015 ;
        RECT 48.860 182.970 49.000 183.510 ;
        RECT 49.230 183.510 51.375 183.650 ;
        RECT 49.230 183.450 49.550 183.510 ;
        RECT 51.085 183.465 51.375 183.510 ;
        RECT 53.370 183.450 53.690 183.710 ;
        RECT 64.425 183.650 64.715 183.695 ;
        RECT 69.010 183.650 69.330 183.710 ;
        RECT 64.425 183.510 69.330 183.650 ;
        RECT 64.425 183.465 64.715 183.510 ;
        RECT 69.010 183.450 69.330 183.510 ;
        RECT 88.345 183.465 88.635 183.695 ;
        RECT 55.325 183.310 55.615 183.355 ;
        RECT 57.510 183.310 57.830 183.370 ;
        RECT 58.565 183.310 59.215 183.355 ;
        RECT 55.325 183.170 59.215 183.310 ;
        RECT 55.325 183.125 55.915 183.170 ;
        RECT 49.245 182.970 49.535 183.015 ;
        RECT 48.860 182.830 49.535 182.970 ;
        RECT 49.245 182.785 49.535 182.830 ;
        RECT 51.545 182.970 51.835 183.015 ;
        RECT 53.830 182.970 54.150 183.030 ;
        RECT 51.545 182.830 54.150 182.970 ;
        RECT 51.545 182.785 51.835 182.830 ;
        RECT 47.940 182.630 48.080 182.785 ;
        RECT 53.830 182.770 54.150 182.830 ;
        RECT 55.625 182.810 55.915 183.125 ;
        RECT 57.510 183.110 57.830 183.170 ;
        RECT 58.565 183.125 59.215 183.170 ;
        RECT 61.190 183.110 61.510 183.370 ;
        RECT 65.805 183.310 66.095 183.355 ;
        RECT 66.710 183.310 67.030 183.370 ;
        RECT 65.805 183.170 67.030 183.310 ;
        RECT 65.805 183.125 66.095 183.170 ;
        RECT 66.710 183.110 67.030 183.170 ;
        RECT 71.425 183.310 71.715 183.355 ;
        RECT 72.230 183.310 72.550 183.370 ;
        RECT 74.665 183.310 75.315 183.355 ;
        RECT 71.425 183.170 75.315 183.310 ;
        RECT 71.425 183.125 72.015 183.170 ;
        RECT 56.705 182.970 56.995 183.015 ;
        RECT 60.285 182.970 60.575 183.015 ;
        RECT 62.120 182.970 62.410 183.015 ;
        RECT 56.705 182.830 62.410 182.970 ;
        RECT 56.705 182.785 56.995 182.830 ;
        RECT 60.285 182.785 60.575 182.830 ;
        RECT 62.120 182.785 62.410 182.830 ;
        RECT 63.965 182.785 64.255 183.015 ;
        RECT 69.485 182.970 69.775 183.015 ;
        RECT 70.390 182.970 70.710 183.030 ;
        RECT 69.485 182.830 70.710 182.970 ;
        RECT 69.485 182.785 69.775 182.830 ;
        RECT 49.690 182.630 50.010 182.690 ;
        RECT 44.260 182.490 47.620 182.630 ;
        RECT 47.940 182.490 50.010 182.630 ;
        RECT 43.265 182.445 43.555 182.490 ;
        RECT 43.710 182.430 44.030 182.490 ;
        RECT 29.005 182.105 29.295 182.335 ;
        RECT 41.410 182.290 41.730 182.350 ;
        RECT 46.025 182.290 46.315 182.335 ;
        RECT 41.410 182.150 46.315 182.290 ;
        RECT 47.480 182.290 47.620 182.490 ;
        RECT 49.690 182.430 50.010 182.490 ;
        RECT 50.610 182.430 50.930 182.690 ;
        RECT 57.970 182.630 58.290 182.690 ;
        RECT 62.585 182.630 62.875 182.675 ;
        RECT 57.970 182.490 62.875 182.630 ;
        RECT 64.040 182.630 64.180 182.785 ;
        RECT 70.390 182.770 70.710 182.830 ;
        RECT 71.725 182.810 72.015 183.125 ;
        RECT 72.230 183.110 72.550 183.170 ;
        RECT 74.665 183.125 75.315 183.170 ;
        RECT 77.290 183.110 77.610 183.370 ;
        RECT 72.805 182.970 73.095 183.015 ;
        RECT 76.385 182.970 76.675 183.015 ;
        RECT 78.220 182.970 78.510 183.015 ;
        RECT 72.805 182.830 78.510 182.970 ;
        RECT 72.805 182.785 73.095 182.830 ;
        RECT 76.385 182.785 76.675 182.830 ;
        RECT 78.220 182.785 78.510 182.830 ;
        RECT 84.650 182.970 84.970 183.030 ;
        RECT 86.045 182.970 86.335 183.015 ;
        RECT 84.650 182.830 86.335 182.970 ;
        RECT 84.650 182.770 84.970 182.830 ;
        RECT 86.045 182.785 86.335 182.830 ;
        RECT 86.490 182.770 86.810 183.030 ;
        RECT 88.420 182.970 88.560 183.465 ;
        RECT 111.790 183.450 112.110 183.710 ;
        RECT 114.105 183.465 114.395 183.695 ;
        RECT 116.865 183.650 117.155 183.695 ;
        RECT 118.230 183.650 118.550 183.710 ;
        RECT 116.865 183.510 118.550 183.650 ;
        RECT 116.865 183.465 117.155 183.510 ;
        RECT 94.885 183.310 95.175 183.355 ;
        RECT 98.125 183.310 98.775 183.355 ;
        RECT 94.885 183.170 98.775 183.310 ;
        RECT 94.885 183.125 95.475 183.170 ;
        RECT 98.125 183.125 98.775 183.170 ;
        RECT 95.185 183.030 95.475 183.125 ;
        RECT 90.645 182.970 90.935 183.015 ;
        RECT 88.420 182.830 90.935 182.970 ;
        RECT 90.645 182.785 90.935 182.830 ;
        RECT 95.185 182.810 95.550 183.030 ;
        RECT 95.230 182.770 95.550 182.810 ;
        RECT 96.265 182.970 96.555 183.015 ;
        RECT 99.845 182.970 100.135 183.015 ;
        RECT 101.680 182.970 101.970 183.015 ;
        RECT 96.265 182.830 101.970 182.970 ;
        RECT 96.265 182.785 96.555 182.830 ;
        RECT 99.845 182.785 100.135 182.830 ;
        RECT 101.680 182.785 101.970 182.830 ;
        RECT 102.145 182.970 102.435 183.015 ;
        RECT 105.810 182.970 106.130 183.030 ;
        RECT 102.145 182.830 106.130 182.970 ;
        RECT 102.145 182.785 102.435 182.830 ;
        RECT 105.810 182.770 106.130 182.830 ;
        RECT 112.250 182.770 112.570 183.030 ;
        RECT 114.180 182.970 114.320 183.465 ;
        RECT 118.230 183.450 118.550 183.510 ;
        RECT 115.945 182.970 116.235 183.015 ;
        RECT 114.180 182.830 116.235 182.970 ;
        RECT 115.945 182.785 116.235 182.830 ;
        RECT 68.090 182.630 68.410 182.690 ;
        RECT 64.040 182.490 68.410 182.630 ;
        RECT 57.970 182.430 58.290 182.490 ;
        RECT 62.585 182.445 62.875 182.490 ;
        RECT 68.090 182.430 68.410 182.490 ;
        RECT 68.550 182.430 68.870 182.690 ;
        RECT 73.610 182.630 73.930 182.690 ;
        RECT 70.020 182.490 73.930 182.630 ;
        RECT 50.700 182.290 50.840 182.430 ;
        RECT 54.750 182.290 55.070 182.350 ;
        RECT 47.480 182.150 55.070 182.290 ;
        RECT 41.410 182.090 41.730 182.150 ;
        RECT 46.025 182.105 46.315 182.150 ;
        RECT 54.750 182.090 55.070 182.150 ;
        RECT 56.705 182.290 56.995 182.335 ;
        RECT 59.825 182.290 60.115 182.335 ;
        RECT 61.715 182.290 62.005 182.335 ;
        RECT 56.705 182.150 62.005 182.290 ;
        RECT 56.705 182.105 56.995 182.150 ;
        RECT 59.825 182.105 60.115 182.150 ;
        RECT 61.715 182.105 62.005 182.150 ;
        RECT 65.805 182.290 66.095 182.335 ;
        RECT 70.020 182.290 70.160 182.490 ;
        RECT 73.610 182.430 73.930 182.490 ;
        RECT 75.450 182.630 75.770 182.690 ;
        RECT 78.685 182.630 78.975 182.675 ;
        RECT 75.450 182.490 78.975 182.630 ;
        RECT 75.450 182.430 75.770 182.490 ;
        RECT 78.685 182.445 78.975 182.490 ;
        RECT 65.805 182.150 70.160 182.290 ;
        RECT 72.805 182.290 73.095 182.335 ;
        RECT 75.925 182.290 76.215 182.335 ;
        RECT 77.815 182.290 78.105 182.335 ;
        RECT 72.805 182.150 78.105 182.290 ;
        RECT 78.760 182.290 78.900 182.445 ;
        RECT 85.110 182.430 85.430 182.690 ;
        RECT 86.580 182.630 86.720 182.770 ;
        RECT 93.405 182.630 93.695 182.675 ;
        RECT 97.530 182.630 97.850 182.690 ;
        RECT 86.580 182.490 97.850 182.630 ;
        RECT 93.405 182.445 93.695 182.490 ;
        RECT 97.530 182.430 97.850 182.490 ;
        RECT 100.750 182.430 101.070 182.690 ;
        RECT 103.050 182.630 103.370 182.690 ;
        RECT 110.885 182.630 111.175 182.675 ;
        RECT 111.790 182.630 112.110 182.690 ;
        RECT 103.050 182.490 112.110 182.630 ;
        RECT 103.050 182.430 103.370 182.490 ;
        RECT 110.885 182.445 111.175 182.490 ;
        RECT 111.790 182.430 112.110 182.490 ;
        RECT 93.850 182.290 94.170 182.350 ;
        RECT 78.760 182.150 94.170 182.290 ;
        RECT 65.805 182.105 66.095 182.150 ;
        RECT 72.805 182.105 73.095 182.150 ;
        RECT 75.925 182.105 76.215 182.150 ;
        RECT 77.815 182.105 78.105 182.150 ;
        RECT 93.850 182.090 94.170 182.150 ;
        RECT 96.265 182.290 96.555 182.335 ;
        RECT 99.385 182.290 99.675 182.335 ;
        RECT 101.275 182.290 101.565 182.335 ;
        RECT 96.265 182.150 101.565 182.290 ;
        RECT 96.265 182.105 96.555 182.150 ;
        RECT 99.385 182.105 99.675 182.150 ;
        RECT 101.275 182.105 101.565 182.150 ;
        RECT 45.565 181.950 45.855 181.995 ;
        RECT 47.850 181.950 48.170 182.010 ;
        RECT 45.565 181.810 48.170 181.950 ;
        RECT 45.565 181.765 45.855 181.810 ;
        RECT 47.850 181.750 48.170 181.810 ;
        RECT 53.830 181.750 54.150 182.010 ;
        RECT 68.550 181.950 68.870 182.010 ;
        RECT 69.470 181.950 69.790 182.010 ;
        RECT 69.945 181.950 70.235 181.995 ;
        RECT 68.550 181.810 70.235 181.950 ;
        RECT 68.550 181.750 68.870 181.810 ;
        RECT 69.470 181.750 69.790 181.810 ;
        RECT 69.945 181.765 70.235 181.810 ;
        RECT 91.090 181.950 91.410 182.010 ;
        RECT 91.565 181.950 91.855 181.995 ;
        RECT 91.090 181.810 91.855 181.950 ;
        RECT 91.090 181.750 91.410 181.810 ;
        RECT 91.565 181.765 91.855 181.810 ;
        RECT 14.660 181.130 127.820 181.610 ;
        RECT 59.825 180.930 60.115 180.975 ;
        RECT 61.190 180.930 61.510 180.990 ;
        RECT 59.825 180.790 61.510 180.930 ;
        RECT 59.825 180.745 60.115 180.790 ;
        RECT 61.190 180.730 61.510 180.790 ;
        RECT 75.005 180.930 75.295 180.975 ;
        RECT 77.290 180.930 77.610 180.990 ;
        RECT 75.005 180.790 77.610 180.930 ;
        RECT 75.005 180.745 75.295 180.790 ;
        RECT 77.290 180.730 77.610 180.790 ;
        RECT 85.110 180.930 85.430 180.990 ;
        RECT 85.110 180.790 94.080 180.930 ;
        RECT 85.110 180.730 85.430 180.790 ;
        RECT 40.605 180.590 40.895 180.635 ;
        RECT 43.725 180.590 44.015 180.635 ;
        RECT 45.615 180.590 45.905 180.635 ;
        RECT 40.605 180.450 45.905 180.590 ;
        RECT 40.605 180.405 40.895 180.450 ;
        RECT 43.725 180.405 44.015 180.450 ;
        RECT 45.615 180.405 45.905 180.450 ;
        RECT 57.525 180.405 57.815 180.635 ;
        RECT 64.410 180.590 64.730 180.650 ;
        RECT 66.710 180.590 67.030 180.650 ;
        RECT 70.850 180.590 71.170 180.650 ;
        RECT 81.430 180.590 81.750 180.650 ;
        RECT 84.650 180.590 84.970 180.650 ;
        RECT 64.410 180.450 72.920 180.590 ;
        RECT 46.485 180.250 46.775 180.295 ;
        RECT 54.290 180.250 54.610 180.310 ;
        RECT 46.485 180.110 54.610 180.250 ;
        RECT 46.485 180.065 46.775 180.110 ;
        RECT 54.290 180.050 54.610 180.110 ;
        RECT 54.750 180.250 55.070 180.310 ;
        RECT 57.050 180.250 57.370 180.310 ;
        RECT 54.750 180.110 57.370 180.250 ;
        RECT 54.750 180.050 55.070 180.110 ;
        RECT 57.050 180.050 57.370 180.110 ;
        RECT 25.770 179.910 26.090 179.970 ;
        RECT 36.365 179.910 36.655 179.955 ;
        RECT 25.770 179.770 36.655 179.910 ;
        RECT 25.770 179.710 26.090 179.770 ;
        RECT 36.365 179.725 36.655 179.770 ;
        RECT 39.525 179.615 39.815 179.930 ;
        RECT 40.605 179.910 40.895 179.955 ;
        RECT 44.185 179.910 44.475 179.955 ;
        RECT 46.020 179.910 46.310 179.955 ;
        RECT 40.605 179.770 46.310 179.910 ;
        RECT 40.605 179.725 40.895 179.770 ;
        RECT 44.185 179.725 44.475 179.770 ;
        RECT 46.020 179.725 46.310 179.770 ;
        RECT 47.850 179.710 48.170 179.970 ;
        RECT 57.600 179.910 57.740 180.405 ;
        RECT 64.410 180.390 64.730 180.450 ;
        RECT 66.710 180.390 67.030 180.450 ;
        RECT 70.850 180.390 71.170 180.450 ;
        RECT 68.090 180.250 68.410 180.310 ;
        RECT 70.280 180.250 70.570 180.295 ;
        RECT 68.090 180.110 70.570 180.250 ;
        RECT 68.090 180.050 68.410 180.110 ;
        RECT 70.280 180.065 70.570 180.110 ;
        RECT 71.310 180.050 71.630 180.310 ;
        RECT 72.780 180.295 72.920 180.450 ;
        RECT 81.430 180.450 84.970 180.590 ;
        RECT 81.430 180.390 81.750 180.450 ;
        RECT 84.650 180.390 84.970 180.450 ;
        RECT 87.525 180.590 87.815 180.635 ;
        RECT 90.645 180.590 90.935 180.635 ;
        RECT 92.535 180.590 92.825 180.635 ;
        RECT 87.525 180.450 92.825 180.590 ;
        RECT 87.525 180.405 87.815 180.450 ;
        RECT 90.645 180.405 90.935 180.450 ;
        RECT 92.535 180.405 92.825 180.450 ;
        RECT 72.705 180.065 72.995 180.295 ;
        RECT 76.370 180.250 76.690 180.310 ;
        RECT 85.110 180.250 85.430 180.310 ;
        RECT 76.370 180.110 85.430 180.250 ;
        RECT 76.370 180.050 76.690 180.110 ;
        RECT 85.110 180.050 85.430 180.110 ;
        RECT 91.550 180.250 91.870 180.310 ;
        RECT 92.025 180.250 92.315 180.295 ;
        RECT 91.550 180.110 92.315 180.250 ;
        RECT 93.940 180.250 94.080 180.790 ;
        RECT 95.230 180.730 95.550 180.990 ;
        RECT 100.750 180.930 101.070 180.990 ;
        RECT 101.225 180.930 101.515 180.975 ;
        RECT 100.750 180.790 101.515 180.930 ;
        RECT 100.750 180.730 101.070 180.790 ;
        RECT 101.225 180.745 101.515 180.790 ;
        RECT 115.945 180.930 116.235 180.975 ;
        RECT 119.150 180.930 119.470 180.990 ;
        RECT 115.945 180.790 119.470 180.930 ;
        RECT 115.945 180.745 116.235 180.790 ;
        RECT 119.150 180.730 119.470 180.790 ;
        RECT 99.845 180.405 100.135 180.635 ;
        RECT 100.840 180.450 118.920 180.590 ;
        RECT 96.625 180.250 96.915 180.295 ;
        RECT 93.940 180.110 96.915 180.250 ;
        RECT 91.550 180.050 91.870 180.110 ;
        RECT 92.025 180.065 92.315 180.110 ;
        RECT 96.625 180.065 96.915 180.110 ;
        RECT 97.530 180.050 97.850 180.310 ;
        RECT 58.905 179.910 59.195 179.955 ;
        RECT 57.600 179.770 59.195 179.910 ;
        RECT 58.905 179.725 59.195 179.770 ;
        RECT 69.025 179.910 69.315 179.955 ;
        RECT 69.470 179.910 69.790 179.970 ;
        RECT 70.865 179.910 71.155 179.955 ;
        RECT 69.025 179.770 71.155 179.910 ;
        RECT 69.025 179.725 69.315 179.770 ;
        RECT 69.470 179.710 69.790 179.770 ;
        RECT 70.865 179.725 71.155 179.770 ;
        RECT 74.545 179.910 74.835 179.955 ;
        RECT 74.990 179.910 75.310 179.970 ;
        RECT 80.985 179.910 81.275 179.955 ;
        RECT 84.650 179.910 84.970 179.970 ;
        RECT 74.545 179.770 75.310 179.910 ;
        RECT 74.545 179.725 74.835 179.770 ;
        RECT 36.825 179.570 37.115 179.615 ;
        RECT 39.225 179.570 39.815 179.615 ;
        RECT 42.465 179.570 43.115 179.615 ;
        RECT 36.825 179.430 43.115 179.570 ;
        RECT 36.825 179.385 37.115 179.430 ;
        RECT 39.225 179.385 39.515 179.430 ;
        RECT 42.465 179.385 43.115 179.430 ;
        RECT 45.105 179.385 45.395 179.615 ;
        RECT 49.230 179.570 49.550 179.630 ;
        RECT 50.150 179.570 50.470 179.630 ;
        RECT 55.685 179.570 55.975 179.615 ;
        RECT 72.230 179.570 72.550 179.630 ;
        RECT 74.620 179.570 74.760 179.725 ;
        RECT 74.990 179.710 75.310 179.770 ;
        RECT 76.460 179.770 84.970 179.910 ;
        RECT 49.230 179.430 55.975 179.570 ;
        RECT 37.745 179.230 38.035 179.275 ;
        RECT 43.710 179.230 44.030 179.290 ;
        RECT 37.745 179.090 44.030 179.230 ;
        RECT 45.180 179.230 45.320 179.385 ;
        RECT 49.230 179.370 49.550 179.430 ;
        RECT 50.150 179.370 50.470 179.430 ;
        RECT 55.685 179.385 55.975 179.430 ;
        RECT 68.180 179.430 74.760 179.570 ;
        RECT 46.945 179.230 47.235 179.275 ;
        RECT 45.180 179.090 47.235 179.230 ;
        RECT 37.745 179.045 38.035 179.090 ;
        RECT 43.710 179.030 44.030 179.090 ;
        RECT 46.945 179.045 47.235 179.090 ;
        RECT 53.830 179.230 54.150 179.290 ;
        RECT 68.180 179.275 68.320 179.430 ;
        RECT 72.230 179.370 72.550 179.430 ;
        RECT 55.225 179.230 55.515 179.275 ;
        RECT 53.830 179.090 55.515 179.230 ;
        RECT 53.830 179.030 54.150 179.090 ;
        RECT 55.225 179.045 55.515 179.090 ;
        RECT 68.105 179.045 68.395 179.275 ;
        RECT 69.470 179.030 69.790 179.290 ;
        RECT 69.930 179.230 70.250 179.290 ;
        RECT 76.460 179.230 76.600 179.770 ;
        RECT 80.985 179.725 81.275 179.770 ;
        RECT 84.650 179.710 84.970 179.770 ;
        RECT 76.830 179.570 77.150 179.630 ;
        RECT 86.445 179.615 86.735 179.930 ;
        RECT 87.525 179.910 87.815 179.955 ;
        RECT 91.105 179.910 91.395 179.955 ;
        RECT 92.940 179.910 93.230 179.955 ;
        RECT 87.525 179.770 93.230 179.910 ;
        RECT 87.525 179.725 87.815 179.770 ;
        RECT 91.105 179.725 91.395 179.770 ;
        RECT 92.940 179.725 93.230 179.770 ;
        RECT 93.405 179.910 93.695 179.955 ;
        RECT 93.850 179.910 94.170 179.970 ;
        RECT 93.405 179.770 94.170 179.910 ;
        RECT 93.405 179.725 93.695 179.770 ;
        RECT 93.850 179.710 94.170 179.770 ;
        RECT 94.785 179.725 95.075 179.955 ;
        RECT 98.005 179.910 98.295 179.955 ;
        RECT 98.450 179.910 98.770 179.970 ;
        RECT 98.005 179.770 98.770 179.910 ;
        RECT 99.920 179.910 100.060 180.405 ;
        RECT 100.305 179.910 100.595 179.955 ;
        RECT 99.920 179.770 100.595 179.910 ;
        RECT 98.005 179.725 98.295 179.770 ;
        RECT 82.365 179.570 82.655 179.615 ;
        RECT 76.830 179.430 82.655 179.570 ;
        RECT 76.830 179.370 77.150 179.430 ;
        RECT 82.365 179.385 82.655 179.430 ;
        RECT 86.145 179.570 86.735 179.615 ;
        RECT 88.330 179.570 88.650 179.630 ;
        RECT 89.385 179.570 90.035 179.615 ;
        RECT 86.145 179.430 90.035 179.570 ;
        RECT 86.145 179.385 86.435 179.430 ;
        RECT 88.330 179.370 88.650 179.430 ;
        RECT 89.385 179.385 90.035 179.430 ;
        RECT 90.630 179.570 90.950 179.630 ;
        RECT 94.860 179.570 95.000 179.725 ;
        RECT 98.450 179.710 98.770 179.770 ;
        RECT 100.305 179.725 100.595 179.770 ;
        RECT 100.840 179.570 100.980 180.450 ;
        RECT 111.790 180.250 112.110 180.310 ;
        RECT 112.725 180.250 113.015 180.295 ;
        RECT 109.580 180.110 111.560 180.250 ;
        RECT 105.350 179.910 105.670 179.970 ;
        RECT 109.580 179.955 109.720 180.110 ;
        RECT 111.420 179.970 111.560 180.110 ;
        RECT 111.790 180.110 113.015 180.250 ;
        RECT 111.790 180.050 112.110 180.110 ;
        RECT 112.725 180.065 113.015 180.110 ;
        RECT 118.780 179.970 118.920 180.450 ;
        RECT 108.585 179.910 108.875 179.955 ;
        RECT 105.350 179.770 108.875 179.910 ;
        RECT 105.350 179.710 105.670 179.770 ;
        RECT 108.585 179.725 108.875 179.770 ;
        RECT 109.045 179.725 109.335 179.955 ;
        RECT 109.505 179.725 109.795 179.955 ;
        RECT 90.630 179.430 100.980 179.570 ;
        RECT 109.120 179.570 109.260 179.725 ;
        RECT 110.410 179.710 110.730 179.970 ;
        RECT 111.330 179.910 111.650 179.970 ;
        RECT 114.105 179.910 114.395 179.955 ;
        RECT 111.330 179.770 114.395 179.910 ;
        RECT 111.330 179.710 111.650 179.770 ;
        RECT 114.105 179.725 114.395 179.770 ;
        RECT 118.690 179.910 119.010 179.970 ;
        RECT 119.165 179.910 119.455 179.955 ;
        RECT 118.690 179.770 119.455 179.910 ;
        RECT 118.690 179.710 119.010 179.770 ;
        RECT 119.165 179.725 119.455 179.770 ;
        RECT 110.870 179.570 111.190 179.630 ;
        RECT 109.120 179.430 111.190 179.570 ;
        RECT 90.630 179.370 90.950 179.430 ;
        RECT 110.870 179.370 111.190 179.430 ;
        RECT 69.930 179.090 76.600 179.230 ;
        RECT 107.205 179.230 107.495 179.275 ;
        RECT 109.030 179.230 109.350 179.290 ;
        RECT 107.205 179.090 109.350 179.230 ;
        RECT 69.930 179.030 70.250 179.090 ;
        RECT 107.205 179.045 107.495 179.090 ;
        RECT 109.030 179.030 109.350 179.090 ;
        RECT 109.490 179.230 109.810 179.290 ;
        RECT 112.250 179.230 112.570 179.290 ;
        RECT 113.645 179.230 113.935 179.275 ;
        RECT 109.490 179.090 113.935 179.230 ;
        RECT 109.490 179.030 109.810 179.090 ;
        RECT 112.250 179.030 112.570 179.090 ;
        RECT 113.645 179.045 113.935 179.090 ;
        RECT 118.705 179.230 118.995 179.275 ;
        RECT 119.150 179.230 119.470 179.290 ;
        RECT 118.705 179.090 119.470 179.230 ;
        RECT 118.705 179.045 118.995 179.090 ;
        RECT 119.150 179.030 119.470 179.090 ;
        RECT 14.660 178.410 127.820 178.890 ;
        RECT 30.830 178.210 31.150 178.270 ;
        RECT 31.305 178.210 31.595 178.255 ;
        RECT 43.250 178.210 43.570 178.270 ;
        RECT 66.710 178.210 67.030 178.270 ;
        RECT 69.930 178.210 70.250 178.270 ;
        RECT 30.830 178.070 34.740 178.210 ;
        RECT 30.830 178.010 31.150 178.070 ;
        RECT 31.305 178.025 31.595 178.070 ;
        RECT 23.930 177.670 24.250 177.930 ;
        RECT 26.230 177.915 26.550 177.930 ;
        RECT 26.225 177.870 26.875 177.915 ;
        RECT 29.825 177.870 30.115 177.915 ;
        RECT 26.225 177.730 30.115 177.870 ;
        RECT 26.225 177.685 26.875 177.730 ;
        RECT 29.525 177.685 30.115 177.730 ;
        RECT 30.370 177.870 30.690 177.930 ;
        RECT 30.370 177.730 33.820 177.870 ;
        RECT 26.230 177.670 26.550 177.685 ;
        RECT 23.030 177.530 23.320 177.575 ;
        RECT 24.865 177.530 25.155 177.575 ;
        RECT 28.445 177.530 28.735 177.575 ;
        RECT 23.030 177.390 28.735 177.530 ;
        RECT 23.030 177.345 23.320 177.390 ;
        RECT 24.865 177.345 25.155 177.390 ;
        RECT 28.445 177.345 28.735 177.390 ;
        RECT 29.525 177.370 29.815 177.685 ;
        RECT 30.370 177.670 30.690 177.730 ;
        RECT 33.680 177.575 33.820 177.730 ;
        RECT 34.600 177.590 34.740 178.070 ;
        RECT 36.670 178.070 64.640 178.210 ;
        RECT 35.890 177.870 36.210 177.930 ;
        RECT 35.060 177.730 36.210 177.870 ;
        RECT 33.145 177.345 33.435 177.575 ;
        RECT 33.605 177.345 33.895 177.575 ;
        RECT 22.565 177.190 22.855 177.235 ;
        RECT 24.390 177.190 24.710 177.250 ;
        RECT 22.565 177.050 24.710 177.190 ;
        RECT 33.220 177.190 33.360 177.345 ;
        RECT 34.510 177.330 34.830 177.590 ;
        RECT 35.060 177.575 35.200 177.730 ;
        RECT 35.890 177.670 36.210 177.730 ;
        RECT 34.985 177.345 35.275 177.575 ;
        RECT 35.445 177.530 35.735 177.575 ;
        RECT 36.670 177.530 36.810 178.070 ;
        RECT 43.250 178.010 43.570 178.070 ;
        RECT 54.290 177.870 54.610 177.930 ;
        RECT 57.970 177.870 58.290 177.930 ;
        RECT 54.290 177.730 58.290 177.870 ;
        RECT 54.290 177.670 54.610 177.730 ;
        RECT 57.970 177.670 58.290 177.730 ;
        RECT 35.445 177.390 36.810 177.530 ;
        RECT 35.445 177.345 35.735 177.390 ;
        RECT 41.885 177.345 42.175 177.575 ;
        RECT 36.350 177.190 36.670 177.250 ;
        RECT 33.220 177.050 36.670 177.190 ;
        RECT 22.565 177.005 22.855 177.050 ;
        RECT 24.390 176.990 24.710 177.050 ;
        RECT 36.350 176.990 36.670 177.050 ;
        RECT 23.435 176.850 23.725 176.895 ;
        RECT 25.325 176.850 25.615 176.895 ;
        RECT 28.445 176.850 28.735 176.895 ;
        RECT 23.435 176.710 28.735 176.850 ;
        RECT 23.435 176.665 23.725 176.710 ;
        RECT 25.325 176.665 25.615 176.710 ;
        RECT 28.445 176.665 28.735 176.710 ;
        RECT 30.830 176.850 31.150 176.910 ;
        RECT 36.825 176.850 37.115 176.895 ;
        RECT 30.830 176.710 37.115 176.850 ;
        RECT 41.960 176.850 42.100 177.345 ;
        RECT 42.790 177.330 43.110 177.590 ;
        RECT 43.265 177.345 43.555 177.575 ;
        RECT 43.725 177.530 44.015 177.575 ;
        RECT 44.170 177.530 44.490 177.590 ;
        RECT 45.090 177.530 45.410 177.590 ;
        RECT 43.725 177.390 45.410 177.530 ;
        RECT 43.725 177.345 44.015 177.390 ;
        RECT 43.340 177.190 43.480 177.345 ;
        RECT 44.170 177.330 44.490 177.390 ;
        RECT 45.090 177.330 45.410 177.390 ;
        RECT 45.550 177.330 45.870 177.590 ;
        RECT 50.470 177.390 64.180 177.530 ;
        RECT 44.630 177.190 44.950 177.250 ;
        RECT 43.340 177.050 44.950 177.190 ;
        RECT 44.630 176.990 44.950 177.050 ;
        RECT 48.310 177.190 48.630 177.250 ;
        RECT 50.470 177.190 50.610 177.390 ;
        RECT 48.310 177.050 50.610 177.190 ;
        RECT 48.310 176.990 48.630 177.050 ;
        RECT 41.960 176.710 46.700 176.850 ;
        RECT 30.830 176.650 31.150 176.710 ;
        RECT 36.825 176.665 37.115 176.710 ;
        RECT 46.560 176.570 46.700 176.710 ;
        RECT 31.290 176.510 31.610 176.570 ;
        RECT 32.225 176.510 32.515 176.555 ;
        RECT 31.290 176.370 32.515 176.510 ;
        RECT 31.290 176.310 31.610 176.370 ;
        RECT 32.225 176.325 32.515 176.370 ;
        RECT 45.090 176.310 45.410 176.570 ;
        RECT 46.470 176.510 46.790 176.570 ;
        RECT 54.750 176.510 55.070 176.570 ;
        RECT 64.040 176.555 64.180 177.390 ;
        RECT 64.500 176.850 64.640 178.070 ;
        RECT 66.710 178.070 70.250 178.210 ;
        RECT 66.710 178.010 67.030 178.070 ;
        RECT 69.930 178.010 70.250 178.070 ;
        RECT 76.370 178.010 76.690 178.270 ;
        RECT 77.290 178.210 77.610 178.270 ;
        RECT 87.885 178.210 88.175 178.255 ;
        RECT 88.330 178.210 88.650 178.270 ;
        RECT 110.870 178.210 111.190 178.270 ;
        RECT 77.290 178.070 84.420 178.210 ;
        RECT 77.290 178.010 77.610 178.070 ;
        RECT 81.430 177.870 81.750 177.930 ;
        RECT 78.300 177.730 81.750 177.870 ;
        RECT 64.870 177.330 65.190 177.590 ;
        RECT 65.345 177.530 65.635 177.575 ;
        RECT 66.250 177.530 66.570 177.590 ;
        RECT 65.345 177.390 66.570 177.530 ;
        RECT 65.345 177.345 65.635 177.390 ;
        RECT 66.250 177.330 66.570 177.390 ;
        RECT 69.930 177.530 70.250 177.590 ;
        RECT 75.005 177.530 75.295 177.575 ;
        RECT 69.930 177.390 75.295 177.530 ;
        RECT 69.930 177.330 70.250 177.390 ;
        RECT 75.005 177.345 75.295 177.390 ;
        RECT 76.370 177.530 76.690 177.590 ;
        RECT 77.290 177.530 77.610 177.590 ;
        RECT 78.300 177.575 78.440 177.730 ;
        RECT 81.430 177.670 81.750 177.730 ;
        RECT 76.370 177.390 77.610 177.530 ;
        RECT 76.370 177.330 76.690 177.390 ;
        RECT 77.290 177.330 77.610 177.390 ;
        RECT 78.225 177.345 78.515 177.575 ;
        RECT 78.670 177.330 78.990 177.590 ;
        RECT 79.130 177.530 79.450 177.590 ;
        RECT 84.280 177.575 84.420 178.070 ;
        RECT 87.885 178.070 88.650 178.210 ;
        RECT 87.885 178.025 88.175 178.070 ;
        RECT 88.330 178.010 88.650 178.070 ;
        RECT 109.580 178.070 111.190 178.210 ;
        RECT 99.830 177.870 100.150 177.930 ;
        RECT 109.580 177.870 109.720 178.070 ;
        RECT 110.870 178.010 111.190 178.070 ;
        RECT 99.830 177.730 109.720 177.870 ;
        RECT 99.830 177.670 100.150 177.730 ;
        RECT 82.365 177.530 82.655 177.575 ;
        RECT 79.130 177.390 82.655 177.530 ;
        RECT 79.130 177.330 79.450 177.390 ;
        RECT 82.365 177.345 82.655 177.390 ;
        RECT 82.825 177.345 83.115 177.575 ;
        RECT 83.285 177.345 83.575 177.575 ;
        RECT 84.205 177.345 84.495 177.575 ;
        RECT 65.790 177.190 66.110 177.250 ;
        RECT 69.010 177.190 69.330 177.250 ;
        RECT 72.690 177.190 73.010 177.250 ;
        RECT 80.970 177.190 81.290 177.250 ;
        RECT 82.900 177.190 83.040 177.345 ;
        RECT 65.790 177.050 73.010 177.190 ;
        RECT 65.790 176.990 66.110 177.050 ;
        RECT 69.010 176.990 69.330 177.050 ;
        RECT 72.690 176.990 73.010 177.050 ;
        RECT 73.240 177.050 81.290 177.190 ;
        RECT 66.265 176.850 66.555 176.895 ;
        RECT 73.240 176.850 73.380 177.050 ;
        RECT 80.970 176.990 81.290 177.050 ;
        RECT 82.440 177.050 83.040 177.190 ;
        RECT 83.360 177.190 83.500 177.345 ;
        RECT 84.650 177.330 84.970 177.590 ;
        RECT 86.045 177.530 86.335 177.575 ;
        RECT 88.345 177.530 88.635 177.575 ;
        RECT 90.630 177.530 90.950 177.590 ;
        RECT 86.045 177.390 90.950 177.530 ;
        RECT 86.045 177.345 86.335 177.390 ;
        RECT 88.345 177.345 88.635 177.390 ;
        RECT 90.630 177.330 90.950 177.390 ;
        RECT 100.305 177.530 100.595 177.575 ;
        RECT 100.750 177.530 101.070 177.590 ;
        RECT 100.305 177.390 101.070 177.530 ;
        RECT 100.305 177.345 100.595 177.390 ;
        RECT 100.750 177.330 101.070 177.390 ;
        RECT 101.210 177.330 101.530 177.590 ;
        RECT 101.760 177.575 101.900 177.730 ;
        RECT 101.685 177.345 101.975 177.575 ;
        RECT 102.145 177.530 102.435 177.575 ;
        RECT 105.350 177.530 105.670 177.590 ;
        RECT 105.900 177.575 106.040 177.730 ;
        RECT 102.145 177.390 105.670 177.530 ;
        RECT 102.145 177.345 102.435 177.390 ;
        RECT 86.950 177.190 87.270 177.250 ;
        RECT 83.360 177.050 87.270 177.190 ;
        RECT 64.500 176.710 73.380 176.850 ;
        RECT 78.670 176.850 78.990 176.910 ;
        RECT 82.440 176.850 82.580 177.050 ;
        RECT 86.950 176.990 87.270 177.050 ;
        RECT 99.370 177.190 99.690 177.250 ;
        RECT 102.220 177.190 102.360 177.345 ;
        RECT 105.350 177.330 105.670 177.390 ;
        RECT 105.825 177.345 106.115 177.575 ;
        RECT 106.270 177.330 106.590 177.590 ;
        RECT 107.205 177.530 107.495 177.575 ;
        RECT 108.570 177.530 108.890 177.590 ;
        RECT 109.580 177.575 109.720 177.730 ;
        RECT 116.965 177.870 117.255 177.915 ;
        RECT 119.150 177.870 119.470 177.930 ;
        RECT 120.205 177.870 120.855 177.915 ;
        RECT 116.965 177.730 120.855 177.870 ;
        RECT 116.965 177.685 117.555 177.730 ;
        RECT 109.045 177.530 109.335 177.575 ;
        RECT 107.205 177.390 107.880 177.530 ;
        RECT 107.205 177.345 107.495 177.390 ;
        RECT 99.370 177.050 102.360 177.190 ;
        RECT 105.440 177.190 105.580 177.330 ;
        RECT 106.730 177.190 107.050 177.250 ;
        RECT 105.440 177.050 107.050 177.190 ;
        RECT 99.370 176.990 99.690 177.050 ;
        RECT 106.730 176.990 107.050 177.050 ;
        RECT 107.740 177.190 107.880 177.390 ;
        RECT 108.570 177.390 109.335 177.530 ;
        RECT 108.570 177.330 108.890 177.390 ;
        RECT 109.045 177.345 109.335 177.390 ;
        RECT 109.505 177.345 109.795 177.575 ;
        RECT 109.950 177.330 110.270 177.590 ;
        RECT 110.885 177.345 111.175 177.575 ;
        RECT 117.265 177.370 117.555 177.685 ;
        RECT 119.150 177.670 119.470 177.730 ;
        RECT 120.205 177.685 120.855 177.730 ;
        RECT 118.345 177.530 118.635 177.575 ;
        RECT 121.925 177.530 122.215 177.575 ;
        RECT 123.760 177.530 124.050 177.575 ;
        RECT 118.345 177.390 124.050 177.530 ;
        RECT 118.345 177.345 118.635 177.390 ;
        RECT 121.925 177.345 122.215 177.390 ;
        RECT 123.760 177.345 124.050 177.390 ;
        RECT 110.410 177.190 110.730 177.250 ;
        RECT 110.960 177.190 111.100 177.345 ;
        RECT 107.740 177.050 111.100 177.190 ;
        RECT 120.990 177.190 121.310 177.250 ;
        RECT 122.845 177.190 123.135 177.235 ;
        RECT 120.990 177.050 123.135 177.190 ;
        RECT 78.670 176.710 82.580 176.850 ;
        RECT 100.750 176.850 101.070 176.910 ;
        RECT 107.740 176.850 107.880 177.050 ;
        RECT 110.410 176.990 110.730 177.050 ;
        RECT 120.990 176.990 121.310 177.050 ;
        RECT 122.845 177.005 123.135 177.050 ;
        RECT 124.210 177.190 124.530 177.250 ;
        RECT 125.590 177.190 125.910 177.250 ;
        RECT 124.210 177.050 125.910 177.190 ;
        RECT 124.210 176.990 124.530 177.050 ;
        RECT 125.590 176.990 125.910 177.050 ;
        RECT 100.750 176.710 107.880 176.850 ;
        RECT 118.345 176.850 118.635 176.895 ;
        RECT 121.465 176.850 121.755 176.895 ;
        RECT 123.355 176.850 123.645 176.895 ;
        RECT 118.345 176.710 123.645 176.850 ;
        RECT 66.265 176.665 66.555 176.710 ;
        RECT 78.670 176.650 78.990 176.710 ;
        RECT 100.750 176.650 101.070 176.710 ;
        RECT 118.345 176.665 118.635 176.710 ;
        RECT 121.465 176.665 121.755 176.710 ;
        RECT 123.355 176.665 123.645 176.710 ;
        RECT 46.470 176.370 55.070 176.510 ;
        RECT 46.470 176.310 46.790 176.370 ;
        RECT 54.750 176.310 55.070 176.370 ;
        RECT 63.965 176.510 64.255 176.555 ;
        RECT 80.050 176.510 80.370 176.570 ;
        RECT 63.965 176.370 80.370 176.510 ;
        RECT 63.965 176.325 64.255 176.370 ;
        RECT 80.050 176.310 80.370 176.370 ;
        RECT 80.510 176.310 80.830 176.570 ;
        RECT 80.985 176.510 81.275 176.555 ;
        RECT 82.810 176.510 83.130 176.570 ;
        RECT 80.985 176.370 83.130 176.510 ;
        RECT 80.985 176.325 81.275 176.370 ;
        RECT 82.810 176.310 83.130 176.370 ;
        RECT 101.670 176.510 101.990 176.570 ;
        RECT 103.525 176.510 103.815 176.555 ;
        RECT 101.670 176.370 103.815 176.510 ;
        RECT 101.670 176.310 101.990 176.370 ;
        RECT 103.525 176.325 103.815 176.370 ;
        RECT 103.970 176.310 104.290 176.570 ;
        RECT 104.890 176.510 105.210 176.570 ;
        RECT 107.665 176.510 107.955 176.555 ;
        RECT 104.890 176.370 107.955 176.510 ;
        RECT 104.890 176.310 105.210 176.370 ;
        RECT 107.665 176.325 107.955 176.370 ;
        RECT 109.950 176.510 110.270 176.570 ;
        RECT 115.485 176.510 115.775 176.555 ;
        RECT 109.950 176.370 115.775 176.510 ;
        RECT 109.950 176.310 110.270 176.370 ;
        RECT 115.485 176.325 115.775 176.370 ;
        RECT 14.660 175.690 127.820 176.170 ;
        RECT 23.930 175.490 24.250 175.550 ;
        RECT 25.785 175.490 26.075 175.535 ;
        RECT 23.930 175.350 26.075 175.490 ;
        RECT 23.930 175.290 24.250 175.350 ;
        RECT 25.785 175.305 26.075 175.350 ;
        RECT 36.350 175.290 36.670 175.550 ;
        RECT 44.630 175.490 44.950 175.550 ;
        RECT 47.850 175.490 48.170 175.550 ;
        RECT 49.690 175.490 50.010 175.550 ;
        RECT 44.630 175.350 53.600 175.490 ;
        RECT 44.630 175.290 44.950 175.350 ;
        RECT 47.850 175.290 48.170 175.350 ;
        RECT 49.690 175.290 50.010 175.350 ;
        RECT 22.105 175.150 22.395 175.195 ;
        RECT 26.230 175.150 26.550 175.210 ;
        RECT 22.105 175.010 26.550 175.150 ;
        RECT 22.105 174.965 22.395 175.010 ;
        RECT 26.230 174.950 26.550 175.010 ;
        RECT 28.035 175.150 28.325 175.195 ;
        RECT 29.925 175.150 30.215 175.195 ;
        RECT 33.045 175.150 33.335 175.195 ;
        RECT 28.035 175.010 33.335 175.150 ;
        RECT 28.035 174.965 28.325 175.010 ;
        RECT 29.925 174.965 30.215 175.010 ;
        RECT 33.045 174.965 33.335 175.010 ;
        RECT 24.390 174.810 24.710 174.870 ;
        RECT 27.165 174.810 27.455 174.855 ;
        RECT 24.390 174.670 27.455 174.810 ;
        RECT 24.390 174.610 24.710 174.670 ;
        RECT 27.165 174.625 27.455 174.670 ;
        RECT 28.545 174.810 28.835 174.855 ;
        RECT 31.290 174.810 31.610 174.870 ;
        RECT 28.545 174.670 31.610 174.810 ;
        RECT 28.545 174.625 28.835 174.670 ;
        RECT 31.290 174.610 31.610 174.670 ;
        RECT 35.430 174.810 35.750 174.870 ;
        RECT 39.125 174.810 39.415 174.855 ;
        RECT 35.430 174.670 39.415 174.810 ;
        RECT 35.430 174.610 35.750 174.670 ;
        RECT 39.125 174.625 39.415 174.670 ;
        RECT 22.565 174.470 22.855 174.515 ;
        RECT 23.025 174.470 23.315 174.515 ;
        RECT 23.930 174.470 24.250 174.530 ;
        RECT 25.770 174.470 26.090 174.530 ;
        RECT 22.565 174.330 26.090 174.470 ;
        RECT 22.565 174.285 22.855 174.330 ;
        RECT 23.025 174.285 23.315 174.330 ;
        RECT 23.930 174.270 24.250 174.330 ;
        RECT 25.770 174.270 26.090 174.330 ;
        RECT 26.690 174.270 27.010 174.530 ;
        RECT 27.630 174.470 27.920 174.515 ;
        RECT 29.465 174.470 29.755 174.515 ;
        RECT 33.045 174.470 33.335 174.515 ;
        RECT 27.630 174.330 33.335 174.470 ;
        RECT 27.630 174.285 27.920 174.330 ;
        RECT 29.465 174.285 29.755 174.330 ;
        RECT 33.045 174.285 33.335 174.330 ;
        RECT 34.125 174.175 34.415 174.490 ;
        RECT 38.205 174.470 38.495 174.515 ;
        RECT 43.710 174.470 44.030 174.530 ;
        RECT 44.720 174.515 44.860 175.290 ;
        RECT 46.010 175.150 46.330 175.210 ;
        RECT 45.180 175.010 46.330 175.150 ;
        RECT 45.180 174.515 45.320 175.010 ;
        RECT 46.010 174.950 46.330 175.010 ;
        RECT 49.230 174.810 49.550 174.870 ;
        RECT 47.480 174.670 49.550 174.810 ;
        RECT 38.205 174.330 44.030 174.470 ;
        RECT 38.205 174.285 38.495 174.330 ;
        RECT 43.710 174.270 44.030 174.330 ;
        RECT 44.185 174.285 44.475 174.515 ;
        RECT 44.645 174.285 44.935 174.515 ;
        RECT 45.105 174.285 45.395 174.515 ;
        RECT 46.025 174.470 46.315 174.515 ;
        RECT 46.470 174.470 46.790 174.530 ;
        RECT 47.480 174.515 47.620 174.670 ;
        RECT 49.230 174.610 49.550 174.670 ;
        RECT 53.460 174.530 53.600 175.350 ;
        RECT 57.050 175.290 57.370 175.550 ;
        RECT 64.870 175.490 65.190 175.550 ;
        RECT 67.185 175.490 67.475 175.535 ;
        RECT 64.870 175.350 67.475 175.490 ;
        RECT 64.870 175.290 65.190 175.350 ;
        RECT 67.185 175.305 67.475 175.350 ;
        RECT 68.550 175.490 68.870 175.550 ;
        RECT 70.405 175.490 70.695 175.535 ;
        RECT 68.550 175.350 70.695 175.490 ;
        RECT 68.550 175.290 68.870 175.350 ;
        RECT 70.405 175.305 70.695 175.350 ;
        RECT 70.850 175.490 71.170 175.550 ;
        RECT 71.310 175.490 71.630 175.550 ;
        RECT 70.850 175.350 71.630 175.490 ;
        RECT 70.850 175.290 71.170 175.350 ;
        RECT 71.310 175.290 71.630 175.350 ;
        RECT 80.050 175.490 80.370 175.550 ;
        RECT 99.830 175.490 100.150 175.550 ;
        RECT 80.050 175.350 100.150 175.490 ;
        RECT 80.050 175.290 80.370 175.350 ;
        RECT 99.830 175.290 100.150 175.350 ;
        RECT 120.990 175.290 121.310 175.550 ;
        RECT 62.585 174.965 62.875 175.195 ;
        RECT 73.610 175.150 73.930 175.210 ;
        RECT 86.030 175.150 86.350 175.210 ;
        RECT 65.420 175.010 73.930 175.150 ;
        RECT 62.660 174.810 62.800 174.965 ;
        RECT 54.380 174.670 62.800 174.810 ;
        RECT 64.410 174.810 64.730 174.870 ;
        RECT 65.420 174.855 65.560 175.010 ;
        RECT 64.885 174.810 65.175 174.855 ;
        RECT 64.410 174.670 65.175 174.810 ;
        RECT 46.025 174.330 46.790 174.470 ;
        RECT 46.025 174.285 46.315 174.330 ;
        RECT 23.485 174.130 23.775 174.175 ;
        RECT 30.825 174.130 31.475 174.175 ;
        RECT 34.125 174.130 34.715 174.175 ;
        RECT 38.665 174.130 38.955 174.175 ;
        RECT 23.485 173.990 34.715 174.130 ;
        RECT 23.485 173.945 23.775 173.990 ;
        RECT 30.825 173.945 31.475 173.990 ;
        RECT 34.425 173.945 34.715 173.990 ;
        RECT 35.980 173.990 38.955 174.130 ;
        RECT 34.970 173.790 35.290 173.850 ;
        RECT 35.980 173.835 36.120 173.990 ;
        RECT 38.665 173.945 38.955 173.990 ;
        RECT 42.790 173.930 43.110 174.190 ;
        RECT 44.260 174.130 44.400 174.285 ;
        RECT 46.470 174.270 46.790 174.330 ;
        RECT 47.405 174.285 47.695 174.515 ;
        RECT 47.850 174.270 48.170 174.530 ;
        RECT 48.325 174.470 48.615 174.515 ;
        RECT 50.150 174.470 50.470 174.530 ;
        RECT 52.925 174.470 53.215 174.515 ;
        RECT 48.325 174.330 53.215 174.470 ;
        RECT 48.325 174.285 48.615 174.330 ;
        RECT 50.150 174.270 50.470 174.330 ;
        RECT 52.925 174.285 53.215 174.330 ;
        RECT 49.705 174.130 49.995 174.175 ;
        RECT 51.545 174.130 51.835 174.175 ;
        RECT 44.260 173.990 44.860 174.130 ;
        RECT 44.720 173.850 44.860 173.990 ;
        RECT 45.640 173.990 49.995 174.130 ;
        RECT 45.640 173.850 45.780 173.990 ;
        RECT 49.705 173.945 49.995 173.990 ;
        RECT 50.240 173.990 51.835 174.130 ;
        RECT 53.000 174.130 53.140 174.285 ;
        RECT 53.370 174.270 53.690 174.530 ;
        RECT 53.830 174.270 54.150 174.530 ;
        RECT 54.380 174.130 54.520 174.670 ;
        RECT 64.410 174.610 64.730 174.670 ;
        RECT 64.885 174.625 65.175 174.670 ;
        RECT 65.345 174.625 65.635 174.855 ;
        RECT 65.790 174.610 66.110 174.870 ;
        RECT 68.180 174.855 68.320 175.010 ;
        RECT 66.265 174.625 66.555 174.855 ;
        RECT 68.105 174.625 68.395 174.855 ;
        RECT 54.750 174.270 55.070 174.530 ;
        RECT 63.505 174.470 63.795 174.515 ;
        RECT 66.340 174.470 66.480 174.625 ;
        RECT 69.010 174.610 69.330 174.870 ;
        RECT 69.485 174.810 69.775 174.855 ;
        RECT 70.850 174.810 71.170 174.870 ;
        RECT 71.860 174.855 72.000 175.010 ;
        RECT 73.610 174.950 73.930 175.010 ;
        RECT 78.300 175.010 86.350 175.150 ;
        RECT 71.325 174.810 71.615 174.855 ;
        RECT 69.485 174.670 71.615 174.810 ;
        RECT 69.485 174.625 69.775 174.670 ;
        RECT 70.850 174.610 71.170 174.670 ;
        RECT 71.325 174.625 71.615 174.670 ;
        RECT 71.785 174.625 72.075 174.855 ;
        RECT 72.230 174.610 72.550 174.870 ;
        RECT 72.690 174.610 73.010 174.870 ;
        RECT 68.565 174.470 68.855 174.515 ;
        RECT 72.320 174.470 72.460 174.610 ;
        RECT 63.505 174.330 64.180 174.470 ;
        RECT 66.340 174.330 72.460 174.470 ;
        RECT 76.370 174.470 76.690 174.530 ;
        RECT 78.300 174.515 78.440 175.010 ;
        RECT 86.030 174.950 86.350 175.010 ;
        RECT 86.505 175.150 86.795 175.195 ;
        RECT 92.010 175.150 92.330 175.210 ;
        RECT 93.850 175.150 94.170 175.210 ;
        RECT 86.505 175.010 94.170 175.150 ;
        RECT 99.920 175.150 100.060 175.290 ;
        RECT 99.920 175.010 109.260 175.150 ;
        RECT 86.505 174.965 86.795 175.010 ;
        RECT 92.010 174.950 92.330 175.010 ;
        RECT 93.850 174.950 94.170 175.010 ;
        RECT 80.970 174.810 81.290 174.870 ;
        RECT 98.450 174.810 98.770 174.870 ;
        RECT 80.970 174.670 98.220 174.810 ;
        RECT 80.970 174.610 81.290 174.670 ;
        RECT 77.305 174.470 77.595 174.515 ;
        RECT 76.370 174.330 77.595 174.470 ;
        RECT 63.505 174.285 63.795 174.330 ;
        RECT 64.040 174.175 64.180 174.330 ;
        RECT 68.565 174.285 68.855 174.330 ;
        RECT 76.370 174.270 76.690 174.330 ;
        RECT 77.305 174.285 77.595 174.330 ;
        RECT 78.225 174.285 78.515 174.515 ;
        RECT 78.670 174.270 78.990 174.530 ;
        RECT 79.130 174.270 79.450 174.530 ;
        RECT 98.080 174.470 98.220 174.670 ;
        RECT 98.450 174.670 100.520 174.810 ;
        RECT 98.450 174.610 98.770 174.670 ;
        RECT 99.370 174.470 99.690 174.530 ;
        RECT 80.140 174.330 97.300 174.470 ;
        RECT 98.080 174.330 99.690 174.470 ;
        RECT 53.000 173.990 54.520 174.130 ;
        RECT 58.445 174.130 58.735 174.175 ;
        RECT 63.965 174.130 64.255 174.175 ;
        RECT 66.250 174.130 66.570 174.190 ;
        RECT 58.445 173.990 63.720 174.130 ;
        RECT 35.905 173.790 36.195 173.835 ;
        RECT 34.970 173.650 36.195 173.790 ;
        RECT 34.970 173.590 35.290 173.650 ;
        RECT 35.905 173.605 36.195 173.650 ;
        RECT 44.630 173.590 44.950 173.850 ;
        RECT 45.550 173.590 45.870 173.850 ;
        RECT 46.010 173.790 46.330 173.850 ;
        RECT 48.310 173.790 48.630 173.850 ;
        RECT 46.010 173.650 48.630 173.790 ;
        RECT 50.240 173.790 50.380 173.990 ;
        RECT 51.545 173.945 51.835 173.990 ;
        RECT 58.445 173.945 58.735 173.990 ;
        RECT 51.070 173.790 51.390 173.850 ;
        RECT 50.240 173.650 51.390 173.790 ;
        RECT 63.580 173.790 63.720 173.990 ;
        RECT 63.965 173.990 66.570 174.130 ;
        RECT 63.965 173.945 64.255 173.990 ;
        RECT 66.250 173.930 66.570 173.990 ;
        RECT 69.010 174.130 69.330 174.190 ;
        RECT 78.760 174.130 78.900 174.270 ;
        RECT 79.590 174.130 79.910 174.190 ;
        RECT 69.010 173.990 78.440 174.130 ;
        RECT 78.760 173.990 79.910 174.130 ;
        RECT 69.010 173.930 69.330 173.990 ;
        RECT 69.930 173.790 70.250 173.850 ;
        RECT 63.580 173.650 70.250 173.790 ;
        RECT 78.300 173.790 78.440 173.990 ;
        RECT 79.590 173.930 79.910 173.990 ;
        RECT 80.140 173.790 80.280 174.330 ;
        RECT 80.510 173.930 80.830 174.190 ;
        RECT 92.930 173.930 93.250 174.190 ;
        RECT 78.300 173.650 80.280 173.790 ;
        RECT 97.160 173.790 97.300 174.330 ;
        RECT 99.370 174.270 99.690 174.330 ;
        RECT 99.830 174.270 100.150 174.530 ;
        RECT 100.380 174.515 100.520 174.670 ;
        RECT 100.305 174.285 100.595 174.515 ;
        RECT 100.750 174.470 101.070 174.530 ;
        RECT 101.225 174.470 101.515 174.515 ;
        RECT 100.750 174.330 101.515 174.470 ;
        RECT 100.750 174.270 101.070 174.330 ;
        RECT 101.225 174.285 101.515 174.330 ;
        RECT 97.530 174.130 97.850 174.190 ;
        RECT 98.005 174.130 98.295 174.175 ;
        RECT 101.300 174.130 101.440 174.285 ;
        RECT 106.270 174.270 106.590 174.530 ;
        RECT 106.730 174.470 107.050 174.530 ;
        RECT 106.730 174.455 108.340 174.470 ;
        RECT 108.570 174.455 108.890 174.530 ;
        RECT 109.120 174.515 109.260 175.010 ;
        RECT 114.090 174.810 114.410 174.870 ;
        RECT 114.090 174.670 120.300 174.810 ;
        RECT 114.090 174.610 114.410 174.670 ;
        RECT 106.730 174.330 108.890 174.455 ;
        RECT 106.730 174.270 107.050 174.330 ;
        RECT 108.200 174.315 108.890 174.330 ;
        RECT 108.570 174.270 108.890 174.315 ;
        RECT 109.045 174.285 109.335 174.515 ;
        RECT 109.490 174.270 109.810 174.530 ;
        RECT 110.410 174.270 110.730 174.530 ;
        RECT 118.245 174.470 118.535 174.515 ;
        RECT 119.150 174.470 119.470 174.530 ;
        RECT 120.160 174.515 120.300 174.670 ;
        RECT 135.635 174.550 136.775 223.880 ;
        RECT 138.130 223.810 139.580 225.110 ;
        RECT 143.180 223.840 144.630 225.140 ;
        RECT 118.245 174.330 119.470 174.470 ;
        RECT 118.245 174.285 118.535 174.330 ;
        RECT 119.150 174.270 119.470 174.330 ;
        RECT 120.085 174.285 120.375 174.515 ;
        RECT 97.530 173.990 98.295 174.130 ;
        RECT 97.530 173.930 97.850 173.990 ;
        RECT 98.005 173.945 98.295 173.990 ;
        RECT 98.540 173.990 101.440 174.130 ;
        RECT 105.350 174.130 105.670 174.190 ;
        RECT 107.205 174.130 107.495 174.175 ;
        RECT 105.350 173.990 107.495 174.130 ;
        RECT 98.540 173.790 98.680 173.990 ;
        RECT 105.350 173.930 105.670 173.990 ;
        RECT 107.205 173.945 107.495 173.990 ;
        RECT 118.705 173.945 118.995 174.175 ;
        RECT 97.160 173.650 98.680 173.790 ;
        RECT 118.230 173.790 118.550 173.850 ;
        RECT 118.780 173.790 118.920 173.945 ;
        RECT 118.230 173.650 118.920 173.790 ;
        RECT 46.010 173.590 46.330 173.650 ;
        RECT 48.310 173.590 48.630 173.650 ;
        RECT 51.070 173.590 51.390 173.650 ;
        RECT 69.930 173.590 70.250 173.650 ;
        RECT 118.230 173.590 118.550 173.650 ;
        RECT 14.660 172.970 127.820 173.450 ;
        RECT 135.580 173.430 136.830 174.550 ;
        RECT 135.635 173.420 136.775 173.430 ;
        RECT 26.690 172.770 27.010 172.830 ;
        RECT 32.225 172.770 32.515 172.815 ;
        RECT 26.690 172.630 32.515 172.770 ;
        RECT 26.690 172.570 27.010 172.630 ;
        RECT 32.225 172.585 32.515 172.630 ;
        RECT 34.510 172.570 34.830 172.830 ;
        RECT 39.110 172.770 39.430 172.830 ;
        RECT 43.250 172.770 43.570 172.830 ;
        RECT 39.110 172.630 43.570 172.770 ;
        RECT 39.110 172.570 39.430 172.630 ;
        RECT 43.250 172.570 43.570 172.630 ;
        RECT 44.630 172.770 44.950 172.830 ;
        RECT 47.390 172.770 47.710 172.830 ;
        RECT 49.690 172.770 50.010 172.830 ;
        RECT 64.885 172.770 65.175 172.815 ;
        RECT 44.630 172.630 47.160 172.770 ;
        RECT 44.630 172.570 44.950 172.630 ;
        RECT 38.190 172.430 38.510 172.490 ;
        RECT 46.010 172.430 46.330 172.490 ;
        RECT 38.190 172.290 40.260 172.430 ;
        RECT 38.190 172.230 38.510 172.290 ;
        RECT 24.390 172.090 24.710 172.150 ;
        RECT 30.845 172.090 31.135 172.135 ;
        RECT 24.390 171.950 31.135 172.090 ;
        RECT 24.390 171.890 24.710 171.950 ;
        RECT 30.845 171.905 31.135 171.950 ;
        RECT 34.065 172.090 34.355 172.135 ;
        RECT 34.970 172.090 35.290 172.150 ;
        RECT 34.065 171.950 35.290 172.090 ;
        RECT 34.065 171.905 34.355 171.950 ;
        RECT 34.970 171.890 35.290 171.950 ;
        RECT 39.110 171.890 39.430 172.150 ;
        RECT 40.120 172.135 40.260 172.290 ;
        RECT 43.800 172.290 46.330 172.430 ;
        RECT 39.585 171.905 39.875 172.135 ;
        RECT 40.045 171.905 40.335 172.135 ;
        RECT 35.430 171.550 35.750 171.810 ;
        RECT 35.890 171.750 36.210 171.810 ;
        RECT 39.660 171.750 39.800 171.905 ;
        RECT 40.950 171.890 41.270 172.150 ;
        RECT 43.250 171.890 43.570 172.150 ;
        RECT 43.800 172.135 43.940 172.290 ;
        RECT 46.010 172.230 46.330 172.290 ;
        RECT 47.020 172.430 47.160 172.630 ;
        RECT 47.390 172.630 65.175 172.770 ;
        RECT 47.390 172.570 47.710 172.630 ;
        RECT 49.690 172.570 50.010 172.630 ;
        RECT 64.885 172.585 65.175 172.630 ;
        RECT 72.245 172.770 72.535 172.815 ;
        RECT 73.610 172.770 73.930 172.830 ;
        RECT 72.245 172.630 73.930 172.770 ;
        RECT 72.245 172.585 72.535 172.630 ;
        RECT 73.610 172.570 73.930 172.630 ;
        RECT 103.065 172.770 103.355 172.815 ;
        RECT 106.270 172.770 106.590 172.830 ;
        RECT 103.065 172.630 106.590 172.770 ;
        RECT 103.065 172.585 103.355 172.630 ;
        RECT 106.270 172.570 106.590 172.630 ;
        RECT 114.090 172.570 114.410 172.830 ;
        RECT 50.150 172.430 50.470 172.490 ;
        RECT 47.020 172.290 50.470 172.430 ;
        RECT 43.725 171.905 44.015 172.135 ;
        RECT 43.800 171.750 43.940 171.905 ;
        RECT 44.170 171.890 44.490 172.150 ;
        RECT 45.105 172.090 45.395 172.135 ;
        RECT 46.470 172.090 46.790 172.150 ;
        RECT 47.020 172.135 47.160 172.290 ;
        RECT 50.150 172.230 50.470 172.290 ;
        RECT 66.250 172.230 66.570 172.490 ;
        RECT 69.930 172.230 70.250 172.490 ;
        RECT 71.310 172.430 71.630 172.490 ;
        RECT 74.545 172.430 74.835 172.475 ;
        RECT 71.310 172.290 74.835 172.430 ;
        RECT 71.310 172.230 71.630 172.290 ;
        RECT 74.545 172.245 74.835 172.290 ;
        RECT 79.590 172.430 79.910 172.490 ;
        RECT 86.490 172.430 86.810 172.490 ;
        RECT 79.590 172.290 83.960 172.430 ;
        RECT 79.590 172.230 79.910 172.290 ;
        RECT 45.105 171.950 46.790 172.090 ;
        RECT 45.105 171.905 45.395 171.950 ;
        RECT 46.470 171.890 46.790 171.950 ;
        RECT 46.945 171.905 47.235 172.135 ;
        RECT 47.390 171.890 47.710 172.150 ;
        RECT 47.865 171.905 48.155 172.135 ;
        RECT 48.785 172.090 49.075 172.135 ;
        RECT 52.910 172.090 53.230 172.150 ;
        RECT 48.785 171.950 53.230 172.090 ;
        RECT 48.785 171.905 49.075 171.950 ;
        RECT 35.890 171.610 43.940 171.750 ;
        RECT 35.890 171.550 36.210 171.610 ;
        RECT 34.050 171.410 34.370 171.470 ;
        RECT 47.940 171.410 48.080 171.905 ;
        RECT 52.910 171.890 53.230 171.950 ;
        RECT 54.290 171.890 54.610 172.150 ;
        RECT 64.870 172.090 65.190 172.150 ;
        RECT 65.805 172.090 66.095 172.135 ;
        RECT 67.645 172.090 67.935 172.135 ;
        RECT 64.870 171.950 67.935 172.090 ;
        RECT 64.870 171.890 65.190 171.950 ;
        RECT 65.805 171.905 66.095 171.950 ;
        RECT 67.645 171.905 67.935 171.950 ;
        RECT 69.485 171.905 69.775 172.135 ;
        RECT 69.560 171.750 69.700 171.905 ;
        RECT 70.850 171.890 71.170 172.150 ;
        RECT 71.785 172.090 72.075 172.135 ;
        RECT 72.690 172.090 73.010 172.150 ;
        RECT 71.785 171.950 73.010 172.090 ;
        RECT 71.785 171.905 72.075 171.950 ;
        RECT 72.690 171.890 73.010 171.950 ;
        RECT 75.465 171.905 75.755 172.135 ;
        RECT 79.130 172.090 79.450 172.150 ;
        RECT 83.820 172.135 83.960 172.290 ;
        RECT 84.280 172.290 86.810 172.430 ;
        RECT 84.280 172.135 84.420 172.290 ;
        RECT 86.490 172.230 86.810 172.290 ;
        RECT 105.810 172.430 106.130 172.490 ;
        RECT 109.505 172.430 109.795 172.475 ;
        RECT 105.810 172.290 109.795 172.430 ;
        RECT 105.810 172.230 106.130 172.290 ;
        RECT 109.505 172.245 109.795 172.290 ;
        RECT 117.425 172.430 117.715 172.475 ;
        RECT 118.230 172.430 118.550 172.490 ;
        RECT 120.665 172.430 121.315 172.475 ;
        RECT 117.425 172.290 121.315 172.430 ;
        RECT 117.425 172.245 118.015 172.290 ;
        RECT 83.285 172.090 83.575 172.135 ;
        RECT 79.130 171.950 83.575 172.090 ;
        RECT 69.930 171.750 70.250 171.810 ;
        RECT 69.560 171.610 70.250 171.750 ;
        RECT 69.930 171.550 70.250 171.610 ;
        RECT 70.405 171.750 70.695 171.795 ;
        RECT 75.540 171.750 75.680 171.905 ;
        RECT 79.130 171.890 79.450 171.950 ;
        RECT 83.285 171.905 83.575 171.950 ;
        RECT 83.745 171.905 84.035 172.135 ;
        RECT 84.205 171.905 84.495 172.135 ;
        RECT 85.125 171.905 85.415 172.135 ;
        RECT 92.010 172.090 92.330 172.150 ;
        RECT 92.945 172.090 93.235 172.135 ;
        RECT 92.010 171.950 93.235 172.090 ;
        RECT 85.200 171.750 85.340 171.905 ;
        RECT 92.010 171.890 92.330 171.950 ;
        RECT 92.945 171.905 93.235 171.950 ;
        RECT 70.405 171.610 75.680 171.750 ;
        RECT 76.460 171.610 85.340 171.750 ;
        RECT 93.020 171.750 93.160 171.905 ;
        RECT 96.150 171.890 96.470 172.150 ;
        RECT 109.950 172.090 110.270 172.150 ;
        RECT 111.805 172.090 112.095 172.135 ;
        RECT 109.950 171.950 112.095 172.090 ;
        RECT 109.950 171.890 110.270 171.950 ;
        RECT 111.805 171.905 112.095 171.950 ;
        RECT 112.265 172.090 112.555 172.135 ;
        RECT 115.470 172.090 115.790 172.150 ;
        RECT 112.265 171.950 115.790 172.090 ;
        RECT 112.265 171.905 112.555 171.950 ;
        RECT 115.470 171.890 115.790 171.950 ;
        RECT 117.725 171.930 118.015 172.245 ;
        RECT 118.230 172.230 118.550 172.290 ;
        RECT 120.665 172.245 121.315 172.290 ;
        RECT 133.700 172.190 134.930 172.680 ;
        RECT 118.805 172.090 119.095 172.135 ;
        RECT 122.385 172.090 122.675 172.135 ;
        RECT 124.220 172.090 124.510 172.135 ;
        RECT 118.805 171.950 124.510 172.090 ;
        RECT 118.805 171.905 119.095 171.950 ;
        RECT 122.385 171.905 122.675 171.950 ;
        RECT 124.220 171.905 124.510 171.950 ;
        RECT 133.700 171.930 136.690 172.190 ;
        RECT 138.330 171.930 139.470 223.810 ;
        RECT 99.830 171.750 100.150 171.810 ;
        RECT 93.020 171.610 100.150 171.750 ;
        RECT 70.405 171.565 70.695 171.610 ;
        RECT 71.860 171.470 72.000 171.610 ;
        RECT 76.460 171.470 76.600 171.610 ;
        RECT 99.830 171.550 100.150 171.610 ;
        RECT 110.410 171.750 110.730 171.810 ;
        RECT 110.885 171.750 111.175 171.795 ;
        RECT 110.410 171.610 111.175 171.750 ;
        RECT 110.410 171.550 110.730 171.610 ;
        RECT 110.885 171.565 111.175 171.610 ;
        RECT 121.450 171.750 121.770 171.810 ;
        RECT 123.305 171.750 123.595 171.795 ;
        RECT 121.450 171.610 123.595 171.750 ;
        RECT 121.450 171.550 121.770 171.610 ;
        RECT 123.305 171.565 123.595 171.610 ;
        RECT 124.685 171.750 124.975 171.795 ;
        RECT 125.590 171.750 125.910 171.810 ;
        RECT 124.685 171.610 125.910 171.750 ;
        RECT 124.685 171.565 124.975 171.610 ;
        RECT 125.590 171.550 125.910 171.610 ;
        RECT 34.050 171.270 48.080 171.410 ;
        RECT 34.050 171.210 34.370 171.270 ;
        RECT 71.770 171.210 72.090 171.470 ;
        RECT 72.230 171.410 72.550 171.470 ;
        RECT 74.545 171.410 74.835 171.455 ;
        RECT 72.230 171.270 74.835 171.410 ;
        RECT 72.230 171.210 72.550 171.270 ;
        RECT 74.545 171.225 74.835 171.270 ;
        RECT 76.370 171.210 76.690 171.470 ;
        RECT 118.805 171.410 119.095 171.455 ;
        RECT 121.925 171.410 122.215 171.455 ;
        RECT 123.815 171.410 124.105 171.455 ;
        RECT 118.805 171.270 124.105 171.410 ;
        RECT 118.805 171.225 119.095 171.270 ;
        RECT 121.925 171.225 122.215 171.270 ;
        RECT 123.815 171.225 124.105 171.270 ;
        RECT 37.270 171.070 37.590 171.130 ;
        RECT 37.745 171.070 38.035 171.115 ;
        RECT 37.270 170.930 38.035 171.070 ;
        RECT 37.270 170.870 37.590 170.930 ;
        RECT 37.745 170.885 38.035 170.930 ;
        RECT 41.870 170.870 42.190 171.130 ;
        RECT 45.565 171.070 45.855 171.115 ;
        RECT 46.010 171.070 46.330 171.130 ;
        RECT 45.565 170.930 46.330 171.070 ;
        RECT 45.565 170.885 45.855 170.930 ;
        RECT 46.010 170.870 46.330 170.930 ;
        RECT 50.150 171.070 50.470 171.130 ;
        RECT 50.610 171.070 50.930 171.130 ;
        RECT 50.150 170.930 50.930 171.070 ;
        RECT 50.150 170.870 50.470 170.930 ;
        RECT 50.610 170.870 50.930 170.930 ;
        RECT 53.370 171.070 53.690 171.130 ;
        RECT 79.590 171.070 79.910 171.130 ;
        RECT 53.370 170.930 79.910 171.070 ;
        RECT 53.370 170.870 53.690 170.930 ;
        RECT 79.590 170.870 79.910 170.930 ;
        RECT 80.050 171.070 80.370 171.130 ;
        RECT 81.905 171.070 82.195 171.115 ;
        RECT 80.050 170.930 82.195 171.070 ;
        RECT 80.050 170.870 80.370 170.930 ;
        RECT 81.905 170.885 82.195 170.930 ;
        RECT 97.070 170.870 97.390 171.130 ;
        RECT 115.470 171.070 115.790 171.130 ;
        RECT 115.945 171.070 116.235 171.115 ;
        RECT 115.470 170.930 116.235 171.070 ;
        RECT 115.470 170.870 115.790 170.930 ;
        RECT 115.945 170.885 116.235 170.930 ;
        RECT 133.700 170.790 139.470 171.930 ;
        RECT 14.660 170.250 127.820 170.730 ;
        RECT 133.700 170.600 136.690 170.790 ;
        RECT 133.700 170.120 134.930 170.600 ;
        RECT 69.025 170.050 69.315 170.095 ;
        RECT 71.770 170.050 72.090 170.110 ;
        RECT 69.025 169.910 72.090 170.050 ;
        RECT 69.025 169.865 69.315 169.910 ;
        RECT 71.770 169.850 72.090 169.910 ;
        RECT 93.020 169.910 102.820 170.050 ;
        RECT 86.045 169.710 86.335 169.755 ;
        RECT 90.170 169.710 90.490 169.770 ;
        RECT 86.045 169.570 90.490 169.710 ;
        RECT 86.045 169.525 86.335 169.570 ;
        RECT 90.170 169.510 90.490 169.570 ;
        RECT 24.390 169.370 24.710 169.430 ;
        RECT 24.865 169.370 25.155 169.415 ;
        RECT 40.950 169.370 41.270 169.430 ;
        RECT 43.250 169.370 43.570 169.430 ;
        RECT 59.825 169.370 60.115 169.415 ;
        RECT 24.390 169.230 25.155 169.370 ;
        RECT 24.390 169.170 24.710 169.230 ;
        RECT 24.865 169.185 25.155 169.230 ;
        RECT 34.140 169.230 43.570 169.370 ;
        RECT 30.370 169.030 30.690 169.090 ;
        RECT 34.140 169.075 34.280 169.230 ;
        RECT 40.950 169.170 41.270 169.230 ;
        RECT 43.250 169.170 43.570 169.230 ;
        RECT 56.220 169.230 60.115 169.370 ;
        RECT 34.065 169.030 34.355 169.075 ;
        RECT 30.370 168.890 34.355 169.030 ;
        RECT 30.370 168.830 30.690 168.890 ;
        RECT 34.065 168.845 34.355 168.890 ;
        RECT 34.970 168.830 35.290 169.090 ;
        RECT 35.430 168.830 35.750 169.090 ;
        RECT 35.905 169.030 36.195 169.075 ;
        RECT 39.110 169.030 39.430 169.090 ;
        RECT 35.905 168.890 39.430 169.030 ;
        RECT 35.905 168.845 36.195 168.890 ;
        RECT 39.110 168.830 39.430 168.890 ;
        RECT 52.450 169.030 52.770 169.090 ;
        RECT 56.220 169.075 56.360 169.230 ;
        RECT 59.825 169.185 60.115 169.230 ;
        RECT 71.310 169.170 71.630 169.430 ;
        RECT 72.245 169.370 72.535 169.415 ;
        RECT 73.610 169.370 73.930 169.430 ;
        RECT 72.245 169.230 73.930 169.370 ;
        RECT 72.245 169.185 72.535 169.230 ;
        RECT 73.610 169.170 73.930 169.230 ;
        RECT 83.270 169.170 83.590 169.430 ;
        RECT 56.145 169.030 56.435 169.075 ;
        RECT 52.450 168.890 56.435 169.030 ;
        RECT 52.450 168.830 52.770 168.890 ;
        RECT 56.145 168.845 56.435 168.890 ;
        RECT 57.525 168.845 57.815 169.075 ;
        RECT 33.605 168.690 33.895 168.735 ;
        RECT 36.350 168.690 36.670 168.750 ;
        RECT 33.605 168.550 36.670 168.690 ;
        RECT 33.605 168.505 33.895 168.550 ;
        RECT 36.350 168.490 36.670 168.550 ;
        RECT 53.830 168.690 54.150 168.750 ;
        RECT 57.600 168.690 57.740 168.845 ;
        RECT 61.190 168.830 61.510 169.090 ;
        RECT 67.170 169.030 67.490 169.090 ;
        RECT 68.565 169.030 68.855 169.075 ;
        RECT 70.865 169.030 71.155 169.075 ;
        RECT 67.170 168.890 71.155 169.030 ;
        RECT 67.170 168.830 67.490 168.890 ;
        RECT 68.565 168.845 68.855 168.890 ;
        RECT 70.865 168.845 71.155 168.890 ;
        RECT 71.785 169.030 72.075 169.075 ;
        RECT 72.690 169.030 73.010 169.090 ;
        RECT 71.785 168.890 73.010 169.030 ;
        RECT 71.785 168.845 72.075 168.890 ;
        RECT 72.690 168.830 73.010 168.890 ;
        RECT 87.425 169.030 87.715 169.075 ;
        RECT 88.790 169.030 89.110 169.090 ;
        RECT 87.425 168.890 89.110 169.030 ;
        RECT 87.425 168.845 87.715 168.890 ;
        RECT 88.790 168.830 89.110 168.890 ;
        RECT 90.185 169.030 90.475 169.075 ;
        RECT 93.020 169.030 93.160 169.910 ;
        RECT 94.425 169.710 94.715 169.755 ;
        RECT 97.545 169.710 97.835 169.755 ;
        RECT 99.435 169.710 99.725 169.755 ;
        RECT 94.425 169.570 99.725 169.710 ;
        RECT 94.425 169.525 94.715 169.570 ;
        RECT 97.545 169.525 97.835 169.570 ;
        RECT 99.435 169.525 99.725 169.570 ;
        RECT 97.070 169.370 97.390 169.430 ;
        RECT 98.925 169.370 99.215 169.415 ;
        RECT 97.070 169.230 99.215 169.370 ;
        RECT 97.070 169.170 97.390 169.230 ;
        RECT 98.925 169.185 99.215 169.230 ;
        RECT 102.680 169.090 102.820 169.910 ;
        RECT 106.270 169.850 106.590 170.110 ;
        RECT 121.450 169.850 121.770 170.110 ;
        RECT 106.360 169.370 106.500 169.850 ;
        RECT 106.845 169.710 107.135 169.755 ;
        RECT 109.965 169.710 110.255 169.755 ;
        RECT 111.855 169.710 112.145 169.755 ;
        RECT 106.845 169.570 112.145 169.710 ;
        RECT 106.845 169.525 107.135 169.570 ;
        RECT 109.965 169.525 110.255 169.570 ;
        RECT 111.855 169.525 112.145 169.570 ;
        RECT 111.330 169.370 111.650 169.430 ;
        RECT 112.725 169.370 113.015 169.415 ;
        RECT 125.590 169.370 125.910 169.430 ;
        RECT 106.360 169.230 125.910 169.370 ;
        RECT 111.330 169.170 111.650 169.230 ;
        RECT 112.725 169.185 113.015 169.230 ;
        RECT 125.590 169.170 125.910 169.230 ;
        RECT 90.185 168.890 93.160 169.030 ;
        RECT 90.185 168.845 90.475 168.890 ;
        RECT 53.830 168.550 57.740 168.690 ;
        RECT 68.090 168.690 68.410 168.750 ;
        RECT 69.945 168.690 70.235 168.735 ;
        RECT 68.090 168.550 70.235 168.690 ;
        RECT 53.830 168.490 54.150 168.550 ;
        RECT 68.090 168.490 68.410 168.550 ;
        RECT 69.945 168.505 70.235 168.550 ;
        RECT 83.730 168.490 84.050 168.750 ;
        RECT 93.345 168.735 93.635 169.050 ;
        RECT 94.425 169.030 94.715 169.075 ;
        RECT 98.005 169.030 98.295 169.075 ;
        RECT 99.840 169.030 100.130 169.075 ;
        RECT 94.425 168.890 100.130 169.030 ;
        RECT 94.425 168.845 94.715 168.890 ;
        RECT 98.005 168.845 98.295 168.890 ;
        RECT 99.840 168.845 100.130 168.890 ;
        RECT 100.290 168.830 100.610 169.090 ;
        RECT 102.590 168.830 102.910 169.090 ;
        RECT 105.765 168.735 106.055 169.050 ;
        RECT 106.845 169.030 107.135 169.075 ;
        RECT 110.425 169.030 110.715 169.075 ;
        RECT 112.260 169.030 112.550 169.075 ;
        RECT 106.845 168.890 112.550 169.030 ;
        RECT 106.845 168.845 107.135 168.890 ;
        RECT 110.425 168.845 110.715 168.890 ;
        RECT 112.260 168.845 112.550 168.890 ;
        RECT 118.690 169.030 119.010 169.090 ;
        RECT 120.545 169.030 120.835 169.075 ;
        RECT 118.690 168.890 120.835 169.030 ;
        RECT 118.690 168.830 119.010 168.890 ;
        RECT 120.545 168.845 120.835 168.890 ;
        RECT 122.845 169.030 123.135 169.075 ;
        RECT 130.190 169.030 130.510 169.090 ;
        RECT 122.845 168.890 130.510 169.030 ;
        RECT 122.845 168.845 123.135 168.890 ;
        RECT 130.190 168.830 130.510 168.890 ;
        RECT 90.645 168.690 90.935 168.735 ;
        RECT 93.045 168.690 93.635 168.735 ;
        RECT 96.285 168.690 96.935 168.735 ;
        RECT 90.645 168.550 96.935 168.690 ;
        RECT 90.645 168.505 90.935 168.550 ;
        RECT 93.045 168.505 93.335 168.550 ;
        RECT 96.285 168.505 96.935 168.550 ;
        RECT 103.065 168.690 103.355 168.735 ;
        RECT 105.465 168.690 106.055 168.735 ;
        RECT 108.705 168.690 109.355 168.735 ;
        RECT 103.065 168.550 109.355 168.690 ;
        RECT 103.065 168.505 103.355 168.550 ;
        RECT 105.465 168.505 105.755 168.550 ;
        RECT 108.705 168.505 109.355 168.550 ;
        RECT 111.345 168.690 111.635 168.735 ;
        RECT 111.790 168.690 112.110 168.750 ;
        RECT 111.345 168.550 112.110 168.690 ;
        RECT 111.345 168.505 111.635 168.550 ;
        RECT 111.790 168.490 112.110 168.550 ;
        RECT 119.610 168.690 119.930 168.750 ;
        RECT 121.925 168.690 122.215 168.735 ;
        RECT 119.610 168.550 122.215 168.690 ;
        RECT 119.610 168.490 119.930 168.550 ;
        RECT 121.925 168.505 122.215 168.550 ;
        RECT 36.810 168.350 37.130 168.410 ;
        RECT 37.285 168.350 37.575 168.395 ;
        RECT 36.810 168.210 37.575 168.350 ;
        RECT 36.810 168.150 37.130 168.210 ;
        RECT 37.285 168.165 37.575 168.210 ;
        RECT 55.670 168.150 55.990 168.410 ;
        RECT 58.445 168.350 58.735 168.395 ;
        RECT 59.350 168.350 59.670 168.410 ;
        RECT 58.445 168.210 59.670 168.350 ;
        RECT 58.445 168.165 58.735 168.210 ;
        RECT 59.350 168.150 59.670 168.210 ;
        RECT 81.430 168.350 81.750 168.410 ;
        RECT 84.205 168.350 84.495 168.395 ;
        RECT 81.430 168.210 84.495 168.350 ;
        RECT 81.430 168.150 81.750 168.210 ;
        RECT 84.205 168.165 84.495 168.210 ;
        RECT 84.650 168.350 84.970 168.410 ;
        RECT 86.965 168.350 87.255 168.395 ;
        RECT 84.650 168.210 87.255 168.350 ;
        RECT 84.650 168.150 84.970 168.210 ;
        RECT 86.965 168.165 87.255 168.210 ;
        RECT 91.565 168.350 91.855 168.395 ;
        RECT 94.310 168.350 94.630 168.410 ;
        RECT 91.565 168.210 94.630 168.350 ;
        RECT 91.565 168.165 91.855 168.210 ;
        RECT 94.310 168.150 94.630 168.210 ;
        RECT 103.985 168.350 104.275 168.395 ;
        RECT 104.430 168.350 104.750 168.410 ;
        RECT 103.985 168.210 104.750 168.350 ;
        RECT 103.985 168.165 104.275 168.210 ;
        RECT 104.430 168.150 104.750 168.210 ;
        RECT 14.660 167.530 127.820 168.010 ;
        RECT 46.470 167.330 46.790 167.390 ;
        RECT 76.370 167.330 76.690 167.390 ;
        RECT 46.470 167.190 70.620 167.330 ;
        RECT 46.470 167.130 46.790 167.190 ;
        RECT 18.360 166.990 18.650 167.035 ;
        RECT 19.330 166.990 19.650 167.050 ;
        RECT 21.620 166.990 21.910 167.035 ;
        RECT 18.360 166.850 21.910 166.990 ;
        RECT 18.360 166.805 18.650 166.850 ;
        RECT 19.330 166.790 19.650 166.850 ;
        RECT 21.620 166.805 21.910 166.850 ;
        RECT 22.540 166.990 22.830 167.035 ;
        RECT 24.400 166.990 24.690 167.035 ;
        RECT 22.540 166.850 24.690 166.990 ;
        RECT 22.540 166.805 22.830 166.850 ;
        RECT 24.400 166.805 24.690 166.850 ;
        RECT 53.485 166.990 53.775 167.035 ;
        RECT 55.670 166.990 55.990 167.050 ;
        RECT 56.725 166.990 57.375 167.035 ;
        RECT 53.485 166.850 57.375 166.990 ;
        RECT 53.485 166.805 54.075 166.850 ;
        RECT 20.220 166.650 20.510 166.695 ;
        RECT 22.540 166.650 22.755 166.805 ;
        RECT 20.220 166.510 22.755 166.650 ;
        RECT 20.220 166.465 20.510 166.510 ;
        RECT 53.785 166.490 54.075 166.805 ;
        RECT 55.670 166.790 55.990 166.850 ;
        RECT 56.725 166.805 57.375 166.850 ;
        RECT 59.350 166.790 59.670 167.050 ;
        RECT 70.480 166.990 70.620 167.190 ;
        RECT 71.170 167.190 76.690 167.330 ;
        RECT 71.170 166.990 71.310 167.190 ;
        RECT 76.370 167.130 76.690 167.190 ;
        RECT 83.730 167.330 84.050 167.390 ;
        RECT 95.245 167.330 95.535 167.375 ;
        RECT 96.150 167.330 96.470 167.390 ;
        RECT 83.730 167.190 86.720 167.330 ;
        RECT 83.730 167.130 84.050 167.190 ;
        RECT 70.480 166.850 71.310 166.990 ;
        RECT 80.070 166.990 80.360 167.035 ;
        RECT 81.930 166.990 82.220 167.035 ;
        RECT 80.070 166.850 82.220 166.990 ;
        RECT 80.070 166.805 80.360 166.850 ;
        RECT 81.930 166.805 82.220 166.850 ;
        RECT 82.850 166.990 83.140 167.035 ;
        RECT 84.650 166.990 84.970 167.050 ;
        RECT 86.110 166.990 86.400 167.035 ;
        RECT 82.850 166.850 86.400 166.990 ;
        RECT 86.580 166.990 86.720 167.190 ;
        RECT 95.245 167.190 96.470 167.330 ;
        RECT 95.245 167.145 95.535 167.190 ;
        RECT 96.150 167.130 96.470 167.190 ;
        RECT 102.590 167.330 102.910 167.390 ;
        RECT 111.345 167.330 111.635 167.375 ;
        RECT 111.790 167.330 112.110 167.390 ;
        RECT 102.590 167.190 106.040 167.330 ;
        RECT 102.590 167.130 102.910 167.190 ;
        RECT 88.115 166.990 88.405 167.035 ;
        RECT 93.405 166.990 93.695 167.035 ;
        RECT 86.580 166.850 93.695 166.990 ;
        RECT 105.900 166.990 106.040 167.190 ;
        RECT 111.345 167.190 112.110 167.330 ;
        RECT 111.345 167.145 111.635 167.190 ;
        RECT 111.790 167.130 112.110 167.190 ;
        RECT 118.690 167.130 119.010 167.390 ;
        RECT 105.900 166.850 119.380 166.990 ;
        RECT 82.850 166.805 83.140 166.850 ;
        RECT 54.865 166.650 55.155 166.695 ;
        RECT 58.445 166.650 58.735 166.695 ;
        RECT 60.280 166.650 60.570 166.695 ;
        RECT 54.865 166.510 60.570 166.650 ;
        RECT 54.865 166.465 55.155 166.510 ;
        RECT 58.445 166.465 58.735 166.510 ;
        RECT 60.280 166.465 60.570 166.510 ;
        RECT 71.770 166.450 72.090 166.710 ;
        RECT 80.970 166.450 81.290 166.710 ;
        RECT 82.005 166.650 82.220 166.805 ;
        RECT 84.650 166.790 84.970 166.850 ;
        RECT 86.110 166.805 86.400 166.850 ;
        RECT 88.115 166.805 88.405 166.850 ;
        RECT 93.405 166.805 93.695 166.850 ;
        RECT 119.240 166.710 119.380 166.850 ;
        RECT 84.250 166.650 84.540 166.695 ;
        RECT 82.005 166.510 84.540 166.650 ;
        RECT 84.250 166.465 84.540 166.510 ;
        RECT 90.170 166.450 90.490 166.710 ;
        RECT 100.750 166.650 101.070 166.710 ;
        RECT 103.985 166.650 104.275 166.695 ;
        RECT 100.750 166.510 104.275 166.650 ;
        RECT 100.750 166.450 101.070 166.510 ;
        RECT 103.985 166.465 104.275 166.510 ;
        RECT 104.430 166.650 104.750 166.710 ;
        RECT 108.585 166.650 108.875 166.695 ;
        RECT 104.430 166.510 108.875 166.650 ;
        RECT 104.430 166.450 104.750 166.510 ;
        RECT 108.585 166.465 108.875 166.510 ;
        RECT 109.045 166.650 109.335 166.695 ;
        RECT 109.950 166.650 110.270 166.710 ;
        RECT 112.265 166.650 112.555 166.695 ;
        RECT 109.045 166.510 110.270 166.650 ;
        RECT 109.045 166.465 109.335 166.510 ;
        RECT 109.950 166.450 110.270 166.510 ;
        RECT 110.960 166.510 112.555 166.650 ;
        RECT 19.790 166.310 20.110 166.370 ;
        RECT 23.485 166.310 23.775 166.355 ;
        RECT 19.790 166.170 23.775 166.310 ;
        RECT 19.790 166.110 20.110 166.170 ;
        RECT 23.485 166.125 23.775 166.170 ;
        RECT 24.390 166.310 24.710 166.370 ;
        RECT 25.325 166.310 25.615 166.355 ;
        RECT 24.390 166.170 25.615 166.310 ;
        RECT 24.390 166.110 24.710 166.170 ;
        RECT 25.325 166.125 25.615 166.170 ;
        RECT 60.730 166.110 61.050 166.370 ;
        RECT 79.145 166.310 79.435 166.355 ;
        RECT 86.030 166.310 86.350 166.370 ;
        RECT 79.145 166.170 86.350 166.310 ;
        RECT 79.145 166.125 79.435 166.170 ;
        RECT 86.030 166.110 86.350 166.170 ;
        RECT 92.025 166.125 92.315 166.355 ;
        RECT 92.945 166.310 93.235 166.355 ;
        RECT 94.310 166.310 94.630 166.370 ;
        RECT 92.945 166.170 94.630 166.310 ;
        RECT 92.945 166.125 93.235 166.170 ;
        RECT 20.220 165.970 20.510 166.015 ;
        RECT 23.000 165.970 23.290 166.015 ;
        RECT 24.860 165.970 25.150 166.015 ;
        RECT 20.220 165.830 25.150 165.970 ;
        RECT 20.220 165.785 20.510 165.830 ;
        RECT 23.000 165.785 23.290 165.830 ;
        RECT 24.860 165.785 25.150 165.830 ;
        RECT 54.865 165.970 55.155 166.015 ;
        RECT 57.985 165.970 58.275 166.015 ;
        RECT 59.875 165.970 60.165 166.015 ;
        RECT 54.865 165.830 60.165 165.970 ;
        RECT 54.865 165.785 55.155 165.830 ;
        RECT 57.985 165.785 58.275 165.830 ;
        RECT 59.875 165.785 60.165 165.830 ;
        RECT 69.930 165.970 70.250 166.030 ;
        RECT 71.310 165.970 71.630 166.030 ;
        RECT 69.930 165.830 71.630 165.970 ;
        RECT 69.930 165.770 70.250 165.830 ;
        RECT 71.310 165.770 71.630 165.830 ;
        RECT 79.610 165.970 79.900 166.015 ;
        RECT 81.470 165.970 81.760 166.015 ;
        RECT 84.250 165.970 84.540 166.015 ;
        RECT 79.610 165.830 84.540 165.970 ;
        RECT 79.610 165.785 79.900 165.830 ;
        RECT 81.470 165.785 81.760 165.830 ;
        RECT 84.250 165.785 84.540 165.830 ;
        RECT 85.110 165.970 85.430 166.030 ;
        RECT 92.100 165.970 92.240 166.125 ;
        RECT 94.310 166.110 94.630 166.170 ;
        RECT 103.065 166.310 103.355 166.355 ;
        RECT 107.650 166.310 107.970 166.370 ;
        RECT 103.065 166.170 107.970 166.310 ;
        RECT 103.065 166.125 103.355 166.170 ;
        RECT 95.690 165.970 96.010 166.030 ;
        RECT 103.140 165.970 103.280 166.125 ;
        RECT 107.650 166.110 107.970 166.170 ;
        RECT 110.960 166.015 111.100 166.510 ;
        RECT 112.265 166.465 112.555 166.510 ;
        RECT 115.470 166.650 115.790 166.710 ;
        RECT 116.405 166.650 116.695 166.695 ;
        RECT 115.470 166.510 116.695 166.650 ;
        RECT 115.470 166.450 115.790 166.510 ;
        RECT 116.405 166.465 116.695 166.510 ;
        RECT 116.850 166.450 117.170 166.710 ;
        RECT 119.150 166.450 119.470 166.710 ;
        RECT 120.990 166.450 121.310 166.710 ;
        RECT 115.945 166.125 116.235 166.355 ;
        RECT 85.110 165.830 103.280 165.970 ;
        RECT 85.110 165.770 85.430 165.830 ;
        RECT 95.690 165.770 96.010 165.830 ;
        RECT 110.885 165.785 111.175 166.015 ;
        RECT 16.355 165.630 16.645 165.675 ;
        RECT 22.550 165.630 22.870 165.690 ;
        RECT 16.355 165.490 22.870 165.630 ;
        RECT 16.355 165.445 16.645 165.490 ;
        RECT 22.550 165.430 22.870 165.490 ;
        RECT 23.930 165.630 24.250 165.690 ;
        RECT 28.530 165.630 28.850 165.690 ;
        RECT 44.170 165.630 44.490 165.690 ;
        RECT 23.930 165.490 44.490 165.630 ;
        RECT 23.930 165.430 24.250 165.490 ;
        RECT 28.530 165.430 28.850 165.490 ;
        RECT 44.170 165.430 44.490 165.490 ;
        RECT 49.230 165.630 49.550 165.690 ;
        RECT 52.005 165.630 52.295 165.675 ;
        RECT 49.230 165.490 52.295 165.630 ;
        RECT 49.230 165.430 49.550 165.490 ;
        RECT 52.005 165.445 52.295 165.490 ;
        RECT 52.910 165.630 53.230 165.690 ;
        RECT 64.870 165.630 65.190 165.690 ;
        RECT 70.865 165.630 71.155 165.675 ;
        RECT 52.910 165.490 71.155 165.630 ;
        RECT 52.910 165.430 53.230 165.490 ;
        RECT 64.870 165.430 65.190 165.490 ;
        RECT 70.865 165.445 71.155 165.490 ;
        RECT 80.970 165.630 81.290 165.690 ;
        RECT 89.265 165.630 89.555 165.675 ;
        RECT 80.970 165.490 89.555 165.630 ;
        RECT 80.970 165.430 81.290 165.490 ;
        RECT 89.265 165.445 89.555 165.490 ;
        RECT 106.270 165.430 106.590 165.690 ;
        RECT 110.410 165.630 110.730 165.690 ;
        RECT 116.020 165.630 116.160 166.125 ;
        RECT 110.410 165.490 116.160 165.630 ;
        RECT 119.625 165.630 119.915 165.675 ;
        RECT 120.070 165.630 120.390 165.690 ;
        RECT 119.625 165.490 120.390 165.630 ;
        RECT 110.410 165.430 110.730 165.490 ;
        RECT 119.625 165.445 119.915 165.490 ;
        RECT 120.070 165.430 120.390 165.490 ;
        RECT 121.450 165.630 121.770 165.690 ;
        RECT 121.925 165.630 122.215 165.675 ;
        RECT 121.450 165.490 122.215 165.630 ;
        RECT 121.450 165.430 121.770 165.490 ;
        RECT 121.925 165.445 122.215 165.490 ;
        RECT 135.580 165.470 136.830 166.590 ;
        RECT 14.660 164.810 127.820 165.290 ;
        RECT 19.330 164.410 19.650 164.670 ;
        RECT 29.925 164.610 30.215 164.655 ;
        RECT 35.430 164.610 35.750 164.670 ;
        RECT 29.925 164.470 35.750 164.610 ;
        RECT 29.925 164.425 30.215 164.470 ;
        RECT 35.430 164.410 35.750 164.470 ;
        RECT 43.250 164.610 43.570 164.670 ;
        RECT 49.705 164.610 49.995 164.655 ;
        RECT 53.830 164.610 54.150 164.670 ;
        RECT 69.010 164.610 69.330 164.670 ;
        RECT 43.250 164.470 48.540 164.610 ;
        RECT 43.250 164.410 43.570 164.470 ;
        RECT 23.945 164.085 24.235 164.315 ;
        RECT 25.310 164.270 25.630 164.330 ;
        RECT 26.245 164.270 26.535 164.315 ;
        RECT 25.310 164.130 26.535 164.270 ;
        RECT 21.185 163.930 21.475 163.975 ;
        RECT 22.090 163.930 22.410 163.990 ;
        RECT 21.185 163.790 22.410 163.930 ;
        RECT 21.185 163.745 21.475 163.790 ;
        RECT 22.090 163.730 22.410 163.790 ;
        RECT 18.870 163.390 19.190 163.650 ;
        RECT 24.020 163.590 24.160 164.085 ;
        RECT 25.310 164.070 25.630 164.130 ;
        RECT 26.245 164.085 26.535 164.130 ;
        RECT 32.785 164.270 33.075 164.315 ;
        RECT 35.905 164.270 36.195 164.315 ;
        RECT 37.795 164.270 38.085 164.315 ;
        RECT 32.785 164.130 38.085 164.270 ;
        RECT 48.400 164.270 48.540 164.470 ;
        RECT 49.705 164.470 54.150 164.610 ;
        RECT 49.705 164.425 49.995 164.470 ;
        RECT 53.830 164.410 54.150 164.470 ;
        RECT 56.220 164.470 69.330 164.610 ;
        RECT 56.220 164.270 56.360 164.470 ;
        RECT 69.010 164.410 69.330 164.470 ;
        RECT 69.470 164.610 69.790 164.670 ;
        RECT 70.865 164.610 71.155 164.655 ;
        RECT 88.345 164.610 88.635 164.655 ;
        RECT 69.470 164.470 71.155 164.610 ;
        RECT 69.470 164.410 69.790 164.470 ;
        RECT 70.865 164.425 71.155 164.470 ;
        RECT 80.600 164.470 88.635 164.610 ;
        RECT 48.400 164.130 56.360 164.270 ;
        RECT 56.705 164.270 56.995 164.315 ;
        RECT 59.825 164.270 60.115 164.315 ;
        RECT 61.715 164.270 62.005 164.315 ;
        RECT 56.705 164.130 62.005 164.270 ;
        RECT 32.785 164.085 33.075 164.130 ;
        RECT 35.905 164.085 36.195 164.130 ;
        RECT 37.795 164.085 38.085 164.130 ;
        RECT 56.705 164.085 56.995 164.130 ;
        RECT 59.825 164.085 60.115 164.130 ;
        RECT 61.715 164.085 62.005 164.130 ;
        RECT 63.950 164.270 64.270 164.330 ;
        RECT 74.070 164.270 74.390 164.330 ;
        RECT 63.950 164.130 74.390 164.270 ;
        RECT 63.950 164.070 64.270 164.130 ;
        RECT 34.970 163.930 35.290 163.990 ;
        RECT 28.160 163.790 35.290 163.930 ;
        RECT 25.325 163.590 25.615 163.635 ;
        RECT 24.020 163.450 25.615 163.590 ;
        RECT 25.325 163.405 25.615 163.450 ;
        RECT 21.630 163.250 21.950 163.310 ;
        RECT 28.160 163.250 28.300 163.790 ;
        RECT 34.970 163.730 35.290 163.790 ;
        RECT 35.430 163.930 35.750 163.990 ;
        RECT 41.425 163.930 41.715 163.975 ;
        RECT 35.430 163.790 41.715 163.930 ;
        RECT 35.430 163.730 35.750 163.790 ;
        RECT 41.425 163.745 41.715 163.790 ;
        RECT 42.345 163.930 42.635 163.975 ;
        RECT 46.485 163.930 46.775 163.975 ;
        RECT 54.750 163.930 55.070 163.990 ;
        RECT 42.345 163.790 55.070 163.930 ;
        RECT 42.345 163.745 42.635 163.790 ;
        RECT 46.485 163.745 46.775 163.790 ;
        RECT 54.750 163.730 55.070 163.790 ;
        RECT 59.350 163.930 59.670 163.990 ;
        RECT 61.205 163.930 61.495 163.975 ;
        RECT 59.350 163.790 61.495 163.930 ;
        RECT 59.350 163.730 59.670 163.790 ;
        RECT 61.205 163.745 61.495 163.790 ;
        RECT 65.805 163.930 66.095 163.975 ;
        RECT 66.250 163.930 66.570 163.990 ;
        RECT 68.640 163.975 68.780 164.130 ;
        RECT 74.070 164.070 74.390 164.130 ;
        RECT 65.805 163.790 66.570 163.930 ;
        RECT 65.805 163.745 66.095 163.790 ;
        RECT 28.530 163.390 28.850 163.650 ;
        RECT 31.705 163.295 31.995 163.610 ;
        RECT 32.785 163.590 33.075 163.635 ;
        RECT 36.365 163.590 36.655 163.635 ;
        RECT 38.200 163.590 38.490 163.635 ;
        RECT 32.785 163.450 38.490 163.590 ;
        RECT 32.785 163.405 33.075 163.450 ;
        RECT 36.365 163.405 36.655 163.450 ;
        RECT 38.200 163.405 38.490 163.450 ;
        RECT 38.665 163.405 38.955 163.635 ;
        RECT 40.965 163.590 41.255 163.635 ;
        RECT 43.710 163.590 44.030 163.650 ;
        RECT 40.965 163.450 44.030 163.590 ;
        RECT 40.965 163.405 41.255 163.450 ;
        RECT 21.630 163.110 28.300 163.250 ;
        RECT 29.005 163.250 29.295 163.295 ;
        RECT 31.405 163.250 31.995 163.295 ;
        RECT 34.645 163.250 35.295 163.295 ;
        RECT 29.005 163.110 35.295 163.250 ;
        RECT 21.630 163.050 21.950 163.110 ;
        RECT 29.005 163.065 29.295 163.110 ;
        RECT 31.405 163.065 31.695 163.110 ;
        RECT 34.645 163.065 35.295 163.110 ;
        RECT 37.285 163.250 37.575 163.295 ;
        RECT 37.730 163.250 38.050 163.310 ;
        RECT 37.285 163.110 38.050 163.250 ;
        RECT 37.285 163.065 37.575 163.110 ;
        RECT 37.730 163.050 38.050 163.110 ;
        RECT 22.105 162.910 22.395 162.955 ;
        RECT 22.550 162.910 22.870 162.970 ;
        RECT 22.105 162.770 22.870 162.910 ;
        RECT 22.105 162.725 22.395 162.770 ;
        RECT 22.550 162.710 22.870 162.770 ;
        RECT 24.390 162.910 24.710 162.970 ;
        RECT 38.740 162.910 38.880 163.405 ;
        RECT 43.710 163.390 44.030 163.450 ;
        RECT 44.170 163.590 44.490 163.650 ;
        RECT 52.450 163.590 52.770 163.650 ;
        RECT 44.170 163.450 52.770 163.590 ;
        RECT 44.170 163.390 44.490 163.450 ;
        RECT 52.450 163.390 52.770 163.450 ;
        RECT 47.405 163.250 47.695 163.295 ;
        RECT 49.230 163.250 49.550 163.310 ;
        RECT 55.625 163.295 55.915 163.610 ;
        RECT 56.705 163.590 56.995 163.635 ;
        RECT 60.285 163.590 60.575 163.635 ;
        RECT 62.120 163.590 62.410 163.635 ;
        RECT 56.705 163.450 62.410 163.590 ;
        RECT 56.705 163.405 56.995 163.450 ;
        RECT 60.285 163.405 60.575 163.450 ;
        RECT 62.120 163.405 62.410 163.450 ;
        RECT 62.585 163.405 62.875 163.635 ;
        RECT 63.950 163.590 64.270 163.650 ;
        RECT 65.880 163.590 66.020 163.745 ;
        RECT 66.250 163.730 66.570 163.790 ;
        RECT 68.565 163.745 68.855 163.975 ;
        RECT 71.310 163.930 71.630 163.990 ;
        RECT 71.785 163.930 72.075 163.975 ;
        RECT 71.310 163.790 72.075 163.930 ;
        RECT 71.310 163.730 71.630 163.790 ;
        RECT 71.785 163.745 72.075 163.790 ;
        RECT 63.950 163.450 66.020 163.590 ;
        RECT 66.710 163.590 67.030 163.650 ;
        RECT 69.485 163.590 69.775 163.635 ;
        RECT 69.930 163.590 70.250 163.650 ;
        RECT 66.710 163.450 70.250 163.590 ;
        RECT 47.405 163.110 49.550 163.250 ;
        RECT 47.405 163.065 47.695 163.110 ;
        RECT 49.230 163.050 49.550 163.110 ;
        RECT 52.925 163.250 53.215 163.295 ;
        RECT 55.325 163.250 55.915 163.295 ;
        RECT 58.565 163.250 59.215 163.295 ;
        RECT 52.925 163.110 59.215 163.250 ;
        RECT 52.925 163.065 53.215 163.110 ;
        RECT 55.325 163.065 55.615 163.110 ;
        RECT 58.565 163.065 59.215 163.110 ;
        RECT 60.730 163.250 61.050 163.310 ;
        RECT 62.660 163.250 62.800 163.405 ;
        RECT 63.950 163.390 64.270 163.450 ;
        RECT 66.710 163.390 67.030 163.450 ;
        RECT 69.485 163.405 69.775 163.450 ;
        RECT 69.930 163.390 70.250 163.450 ;
        RECT 70.405 163.405 70.695 163.635 ;
        RECT 71.860 163.590 72.000 163.745 ;
        RECT 72.230 163.730 72.550 163.990 ;
        RECT 73.150 163.590 73.470 163.650 ;
        RECT 71.860 163.450 73.470 163.590 ;
        RECT 60.730 163.110 62.800 163.250 ;
        RECT 68.550 163.250 68.870 163.310 ;
        RECT 70.480 163.250 70.620 163.405 ;
        RECT 73.150 163.390 73.470 163.450 ;
        RECT 75.465 163.590 75.755 163.635 ;
        RECT 79.590 163.590 79.910 163.650 ;
        RECT 75.465 163.450 79.910 163.590 ;
        RECT 75.465 163.405 75.755 163.450 ;
        RECT 79.590 163.390 79.910 163.450 ;
        RECT 68.550 163.110 70.620 163.250 ;
        RECT 60.730 163.050 61.050 163.110 ;
        RECT 68.550 163.050 68.870 163.110 ;
        RECT 73.625 163.065 73.915 163.295 ;
        RECT 79.080 163.250 79.370 163.295 ;
        RECT 80.600 163.250 80.740 164.470 ;
        RECT 88.345 164.425 88.635 164.470 ;
        RECT 107.650 164.610 107.970 164.670 ;
        RECT 110.410 164.610 110.730 164.670 ;
        RECT 120.990 164.610 121.310 164.670 ;
        RECT 107.650 164.470 112.940 164.610 ;
        RECT 107.650 164.410 107.970 164.470 ;
        RECT 110.410 164.410 110.730 164.470 ;
        RECT 80.940 164.270 81.230 164.315 ;
        RECT 83.720 164.270 84.010 164.315 ;
        RECT 85.580 164.270 85.870 164.315 ;
        RECT 99.830 164.270 100.150 164.330 ;
        RECT 80.940 164.130 85.870 164.270 ;
        RECT 80.940 164.085 81.230 164.130 ;
        RECT 83.720 164.085 84.010 164.130 ;
        RECT 85.580 164.085 85.870 164.130 ;
        RECT 86.120 164.130 100.150 164.270 ;
        RECT 86.120 163.990 86.260 164.130 ;
        RECT 99.830 164.070 100.150 164.130 ;
        RECT 106.240 164.270 106.530 164.315 ;
        RECT 109.020 164.270 109.310 164.315 ;
        RECT 110.880 164.270 111.170 164.315 ;
        RECT 106.240 164.130 111.170 164.270 ;
        RECT 106.240 164.085 106.530 164.130 ;
        RECT 109.020 164.085 109.310 164.130 ;
        RECT 110.880 164.085 111.170 164.130 ;
        RECT 83.270 163.930 83.590 163.990 ;
        RECT 84.650 163.930 84.970 163.990 ;
        RECT 83.270 163.790 84.970 163.930 ;
        RECT 83.270 163.730 83.590 163.790 ;
        RECT 84.650 163.730 84.970 163.790 ;
        RECT 86.030 163.730 86.350 163.990 ;
        RECT 95.690 163.730 96.010 163.990 ;
        RECT 100.750 163.930 101.070 163.990 ;
        RECT 102.375 163.930 102.665 163.975 ;
        RECT 97.160 163.790 102.665 163.930 ;
        RECT 80.940 163.590 81.230 163.635 ;
        RECT 84.205 163.590 84.495 163.635 ;
        RECT 80.940 163.450 83.475 163.590 ;
        RECT 80.940 163.405 81.230 163.450 ;
        RECT 83.260 163.295 83.475 163.450 ;
        RECT 84.205 163.450 86.720 163.590 ;
        RECT 84.205 163.405 84.495 163.450 ;
        RECT 82.340 163.250 82.630 163.295 ;
        RECT 79.080 163.110 82.630 163.250 ;
        RECT 79.080 163.065 79.370 163.110 ;
        RECT 82.340 163.065 82.630 163.110 ;
        RECT 83.260 163.250 83.550 163.295 ;
        RECT 85.120 163.250 85.410 163.295 ;
        RECT 83.260 163.110 85.410 163.250 ;
        RECT 83.260 163.065 83.550 163.110 ;
        RECT 85.120 163.065 85.410 163.110 ;
        RECT 24.390 162.770 38.880 162.910 ;
        RECT 24.390 162.710 24.710 162.770 ;
        RECT 39.110 162.710 39.430 162.970 ;
        RECT 43.725 162.910 44.015 162.955 ;
        RECT 44.170 162.910 44.490 162.970 ;
        RECT 43.725 162.770 44.490 162.910 ;
        RECT 43.725 162.725 44.015 162.770 ;
        RECT 44.170 162.710 44.490 162.770 ;
        RECT 46.470 162.910 46.790 162.970 ;
        RECT 47.865 162.910 48.155 162.955 ;
        RECT 53.830 162.910 54.150 162.970 ;
        RECT 46.470 162.770 54.150 162.910 ;
        RECT 46.470 162.710 46.790 162.770 ;
        RECT 47.865 162.725 48.155 162.770 ;
        RECT 53.830 162.710 54.150 162.770 ;
        RECT 72.230 162.910 72.550 162.970 ;
        RECT 73.700 162.910 73.840 163.065 ;
        RECT 72.230 162.770 73.840 162.910 ;
        RECT 77.075 162.910 77.365 162.955 ;
        RECT 81.430 162.910 81.750 162.970 ;
        RECT 86.580 162.955 86.720 163.450 ;
        RECT 87.410 163.390 87.730 163.650 ;
        RECT 88.790 163.590 89.110 163.650 ;
        RECT 97.160 163.635 97.300 163.790 ;
        RECT 100.750 163.730 101.070 163.790 ;
        RECT 102.375 163.745 102.665 163.790 ;
        RECT 103.140 163.790 110.180 163.930 ;
        RECT 88.790 163.450 95.920 163.590 ;
        RECT 88.790 163.390 89.110 163.450 ;
        RECT 95.780 163.310 95.920 163.450 ;
        RECT 97.085 163.405 97.375 163.635 ;
        RECT 100.305 163.590 100.595 163.635 ;
        RECT 103.140 163.590 103.280 163.790 ;
        RECT 100.305 163.450 103.280 163.590 ;
        RECT 106.240 163.590 106.530 163.635 ;
        RECT 106.240 163.450 108.775 163.590 ;
        RECT 100.305 163.405 100.595 163.450 ;
        RECT 106.240 163.405 106.530 163.450 ;
        RECT 95.690 163.250 96.010 163.310 ;
        RECT 100.380 163.250 100.520 163.405 ;
        RECT 108.560 163.295 108.775 163.450 ;
        RECT 109.490 163.390 109.810 163.650 ;
        RECT 110.040 163.590 110.180 163.790 ;
        RECT 111.330 163.730 111.650 163.990 ;
        RECT 112.800 163.975 112.940 164.470 ;
        RECT 117.860 164.470 121.310 164.610 ;
        RECT 115.945 164.270 116.235 164.315 ;
        RECT 117.860 164.270 118.000 164.470 ;
        RECT 120.990 164.410 121.310 164.470 ;
        RECT 115.945 164.130 118.000 164.270 ;
        RECT 119.265 164.270 119.555 164.315 ;
        RECT 122.385 164.270 122.675 164.315 ;
        RECT 124.275 164.270 124.565 164.315 ;
        RECT 119.265 164.130 124.565 164.270 ;
        RECT 115.945 164.085 116.235 164.130 ;
        RECT 119.265 164.085 119.555 164.130 ;
        RECT 122.385 164.085 122.675 164.130 ;
        RECT 124.275 164.085 124.565 164.130 ;
        RECT 112.725 163.745 113.015 163.975 ;
        RECT 121.450 163.930 121.770 163.990 ;
        RECT 123.765 163.930 124.055 163.975 ;
        RECT 121.450 163.790 124.055 163.930 ;
        RECT 121.450 163.730 121.770 163.790 ;
        RECT 123.765 163.745 124.055 163.790 ;
        RECT 117.310 163.590 117.630 163.650 ;
        RECT 110.040 163.450 117.630 163.590 ;
        RECT 117.310 163.390 117.630 163.450 ;
        RECT 95.690 163.110 100.520 163.250 ;
        RECT 100.765 163.250 101.055 163.295 ;
        RECT 104.380 163.250 104.670 163.295 ;
        RECT 107.640 163.250 107.930 163.295 ;
        RECT 100.765 163.110 107.930 163.250 ;
        RECT 95.690 163.050 96.010 163.110 ;
        RECT 100.765 163.065 101.055 163.110 ;
        RECT 104.380 163.065 104.670 163.110 ;
        RECT 107.640 163.065 107.930 163.110 ;
        RECT 108.560 163.250 108.850 163.295 ;
        RECT 110.420 163.250 110.710 163.295 ;
        RECT 108.560 163.110 110.710 163.250 ;
        RECT 108.560 163.065 108.850 163.110 ;
        RECT 110.420 163.065 110.710 163.110 ;
        RECT 113.170 163.250 113.490 163.310 ;
        RECT 113.645 163.250 113.935 163.295 ;
        RECT 116.850 163.250 117.170 163.310 ;
        RECT 118.185 163.295 118.475 163.610 ;
        RECT 119.265 163.590 119.555 163.635 ;
        RECT 122.845 163.590 123.135 163.635 ;
        RECT 124.680 163.590 124.970 163.635 ;
        RECT 119.265 163.450 124.970 163.590 ;
        RECT 119.265 163.405 119.555 163.450 ;
        RECT 122.845 163.405 123.135 163.450 ;
        RECT 124.680 163.405 124.970 163.450 ;
        RECT 125.145 163.590 125.435 163.635 ;
        RECT 125.590 163.590 125.910 163.650 ;
        RECT 125.145 163.450 125.910 163.590 ;
        RECT 125.145 163.405 125.435 163.450 ;
        RECT 125.590 163.390 125.910 163.450 ;
        RECT 113.170 163.110 117.170 163.250 ;
        RECT 113.170 163.050 113.490 163.110 ;
        RECT 113.645 163.065 113.935 163.110 ;
        RECT 77.075 162.770 81.750 162.910 ;
        RECT 72.230 162.710 72.550 162.770 ;
        RECT 77.075 162.725 77.365 162.770 ;
        RECT 81.430 162.710 81.750 162.770 ;
        RECT 86.505 162.725 86.795 162.955 ;
        RECT 93.850 162.910 94.170 162.970 ;
        RECT 96.625 162.910 96.915 162.955 ;
        RECT 93.850 162.770 96.915 162.910 ;
        RECT 93.850 162.710 94.170 162.770 ;
        RECT 96.625 162.725 96.915 162.770 ;
        RECT 98.925 162.910 99.215 162.955 ;
        RECT 101.210 162.910 101.530 162.970 ;
        RECT 98.925 162.770 101.530 162.910 ;
        RECT 98.925 162.725 99.215 162.770 ;
        RECT 101.210 162.710 101.530 162.770 ;
        RECT 110.870 162.910 111.190 162.970 ;
        RECT 116.480 162.955 116.620 163.110 ;
        RECT 116.850 163.050 117.170 163.110 ;
        RECT 117.885 163.250 118.475 163.295 ;
        RECT 120.070 163.250 120.390 163.310 ;
        RECT 121.125 163.250 121.775 163.295 ;
        RECT 117.885 163.110 121.775 163.250 ;
        RECT 117.885 163.065 118.175 163.110 ;
        RECT 120.070 163.050 120.390 163.110 ;
        RECT 121.125 163.065 121.775 163.110 ;
        RECT 114.105 162.910 114.395 162.955 ;
        RECT 110.870 162.770 114.395 162.910 ;
        RECT 110.870 162.710 111.190 162.770 ;
        RECT 114.105 162.725 114.395 162.770 ;
        RECT 116.405 162.725 116.695 162.955 ;
        RECT 14.660 162.090 127.820 162.570 ;
        RECT 18.195 161.890 18.485 161.935 ;
        RECT 21.630 161.890 21.950 161.950 ;
        RECT 18.195 161.750 21.950 161.890 ;
        RECT 18.195 161.705 18.485 161.750 ;
        RECT 21.630 161.690 21.950 161.750 ;
        RECT 38.190 161.890 38.510 161.950 ;
        RECT 39.125 161.890 39.415 161.935 ;
        RECT 38.190 161.750 39.415 161.890 ;
        RECT 38.190 161.690 38.510 161.750 ;
        RECT 39.125 161.705 39.415 161.750 ;
        RECT 40.505 161.890 40.795 161.935 ;
        RECT 43.710 161.890 44.030 161.950 ;
        RECT 49.705 161.890 49.995 161.935 ;
        RECT 40.505 161.750 44.030 161.890 ;
        RECT 40.505 161.705 40.795 161.750 ;
        RECT 43.710 161.690 44.030 161.750 ;
        RECT 47.940 161.750 49.995 161.890 ;
        RECT 31.290 161.595 31.610 161.610 ;
        RECT 17.045 161.550 17.335 161.595 ;
        RECT 20.200 161.550 20.490 161.595 ;
        RECT 23.460 161.550 23.750 161.595 ;
        RECT 17.045 161.410 23.750 161.550 ;
        RECT 17.045 161.365 17.335 161.410 ;
        RECT 20.200 161.365 20.490 161.410 ;
        RECT 23.460 161.365 23.750 161.410 ;
        RECT 24.380 161.550 24.670 161.595 ;
        RECT 26.240 161.550 26.530 161.595 ;
        RECT 24.380 161.410 26.530 161.550 ;
        RECT 24.380 161.365 24.670 161.410 ;
        RECT 26.240 161.365 26.530 161.410 ;
        RECT 28.550 161.550 28.840 161.595 ;
        RECT 30.410 161.550 30.700 161.595 ;
        RECT 28.550 161.410 30.700 161.550 ;
        RECT 28.550 161.365 28.840 161.410 ;
        RECT 30.410 161.365 30.700 161.410 ;
        RECT 17.505 161.210 17.795 161.255 ;
        RECT 18.870 161.210 19.190 161.270 ;
        RECT 20.710 161.210 21.030 161.270 ;
        RECT 17.505 161.070 21.030 161.210 ;
        RECT 17.505 161.025 17.795 161.070 ;
        RECT 18.870 161.010 19.190 161.070 ;
        RECT 20.710 161.010 21.030 161.070 ;
        RECT 22.060 161.210 22.350 161.255 ;
        RECT 24.380 161.210 24.595 161.365 ;
        RECT 22.060 161.070 24.595 161.210 ;
        RECT 22.060 161.025 22.350 161.070 ;
        RECT 25.310 161.010 25.630 161.270 ;
        RECT 30.485 161.210 30.700 161.365 ;
        RECT 31.290 161.550 31.620 161.595 ;
        RECT 34.590 161.550 34.880 161.595 ;
        RECT 31.290 161.410 34.880 161.550 ;
        RECT 31.290 161.365 31.620 161.410 ;
        RECT 34.590 161.365 34.880 161.410 ;
        RECT 41.985 161.550 42.275 161.595 ;
        RECT 44.170 161.550 44.490 161.610 ;
        RECT 47.940 161.595 48.080 161.750 ;
        RECT 49.705 161.705 49.995 161.750 ;
        RECT 53.830 161.890 54.150 161.950 ;
        RECT 54.765 161.890 55.055 161.935 ;
        RECT 53.830 161.750 55.055 161.890 ;
        RECT 53.830 161.690 54.150 161.750 ;
        RECT 54.765 161.705 55.055 161.750 ;
        RECT 59.350 161.890 59.670 161.950 ;
        RECT 59.825 161.890 60.115 161.935 ;
        RECT 59.350 161.750 60.115 161.890 ;
        RECT 59.350 161.690 59.670 161.750 ;
        RECT 59.825 161.705 60.115 161.750 ;
        RECT 69.010 161.890 69.330 161.950 ;
        RECT 70.405 161.890 70.695 161.935 ;
        RECT 69.010 161.750 70.695 161.890 ;
        RECT 69.010 161.690 69.330 161.750 ;
        RECT 70.405 161.705 70.695 161.750 ;
        RECT 80.985 161.890 81.275 161.935 ;
        RECT 81.430 161.890 81.750 161.950 ;
        RECT 80.985 161.750 81.750 161.890 ;
        RECT 80.985 161.705 81.275 161.750 ;
        RECT 81.430 161.690 81.750 161.750 ;
        RECT 83.285 161.890 83.575 161.935 ;
        RECT 87.410 161.890 87.730 161.950 ;
        RECT 83.285 161.750 87.730 161.890 ;
        RECT 83.285 161.705 83.575 161.750 ;
        RECT 87.410 161.690 87.730 161.750 ;
        RECT 100.305 161.705 100.595 161.935 ;
        RECT 107.205 161.890 107.495 161.935 ;
        RECT 109.490 161.890 109.810 161.950 ;
        RECT 107.205 161.750 109.810 161.890 ;
        RECT 107.205 161.705 107.495 161.750 ;
        RECT 45.225 161.550 45.875 161.595 ;
        RECT 41.985 161.410 45.875 161.550 ;
        RECT 41.985 161.365 42.575 161.410 ;
        RECT 31.290 161.350 31.610 161.365 ;
        RECT 32.730 161.210 33.020 161.255 ;
        RECT 30.485 161.070 33.020 161.210 ;
        RECT 32.730 161.025 33.020 161.070 ;
        RECT 38.650 161.010 38.970 161.270 ;
        RECT 39.110 161.210 39.430 161.270 ;
        RECT 40.045 161.210 40.335 161.255 ;
        RECT 39.110 161.070 40.335 161.210 ;
        RECT 39.110 161.010 39.430 161.070 ;
        RECT 40.045 161.025 40.335 161.070 ;
        RECT 42.285 161.050 42.575 161.365 ;
        RECT 44.170 161.350 44.490 161.410 ;
        RECT 45.225 161.365 45.875 161.410 ;
        RECT 47.865 161.365 48.155 161.595 ;
        RECT 54.290 161.550 54.610 161.610 ;
        RECT 60.730 161.550 61.050 161.610 ;
        RECT 49.320 161.410 61.050 161.550 ;
        RECT 49.320 161.255 49.460 161.410 ;
        RECT 54.290 161.350 54.610 161.410 ;
        RECT 60.730 161.350 61.050 161.410 ;
        RECT 67.645 161.550 67.935 161.595 ;
        RECT 72.230 161.550 72.550 161.610 ;
        RECT 88.790 161.550 89.110 161.610 ;
        RECT 67.645 161.410 72.550 161.550 ;
        RECT 67.645 161.365 67.935 161.410 ;
        RECT 72.230 161.350 72.550 161.410 ;
        RECT 85.660 161.410 89.110 161.550 ;
        RECT 43.365 161.210 43.655 161.255 ;
        RECT 46.945 161.210 47.235 161.255 ;
        RECT 48.780 161.210 49.070 161.255 ;
        RECT 43.365 161.070 49.070 161.210 ;
        RECT 43.365 161.025 43.655 161.070 ;
        RECT 46.945 161.025 47.235 161.070 ;
        RECT 48.780 161.025 49.070 161.070 ;
        RECT 49.245 161.025 49.535 161.255 ;
        RECT 49.690 161.210 50.010 161.270 ;
        RECT 50.625 161.210 50.915 161.255 ;
        RECT 49.690 161.070 50.915 161.210 ;
        RECT 49.690 161.010 50.010 161.070 ;
        RECT 50.625 161.025 50.915 161.070 ;
        RECT 52.005 161.210 52.295 161.255 ;
        RECT 52.450 161.210 52.770 161.270 ;
        RECT 52.005 161.070 52.770 161.210 ;
        RECT 52.005 161.025 52.295 161.070 ;
        RECT 52.450 161.010 52.770 161.070 ;
        RECT 52.910 161.210 53.230 161.270 ;
        RECT 55.225 161.210 55.515 161.255 ;
        RECT 58.905 161.210 59.195 161.255 ;
        RECT 52.910 161.070 55.515 161.210 ;
        RECT 52.910 161.010 53.230 161.070 ;
        RECT 55.225 161.025 55.515 161.070 ;
        RECT 57.140 161.070 59.195 161.210 ;
        RECT 24.390 160.870 24.710 160.930 ;
        RECT 26.230 160.870 26.550 160.930 ;
        RECT 27.165 160.870 27.455 160.915 ;
        RECT 27.625 160.870 27.915 160.915 ;
        RECT 24.390 160.730 27.915 160.870 ;
        RECT 24.390 160.670 24.710 160.730 ;
        RECT 26.230 160.670 26.550 160.730 ;
        RECT 27.165 160.685 27.455 160.730 ;
        RECT 27.625 160.685 27.915 160.730 ;
        RECT 29.465 160.870 29.755 160.915 ;
        RECT 29.465 160.730 37.960 160.870 ;
        RECT 29.465 160.685 29.755 160.730 ;
        RECT 37.820 160.575 37.960 160.730 ;
        RECT 54.305 160.685 54.595 160.915 ;
        RECT 22.060 160.530 22.350 160.575 ;
        RECT 24.840 160.530 25.130 160.575 ;
        RECT 26.700 160.530 26.990 160.575 ;
        RECT 22.060 160.390 26.990 160.530 ;
        RECT 22.060 160.345 22.350 160.390 ;
        RECT 24.840 160.345 25.130 160.390 ;
        RECT 26.700 160.345 26.990 160.390 ;
        RECT 28.090 160.530 28.380 160.575 ;
        RECT 29.950 160.530 30.240 160.575 ;
        RECT 32.730 160.530 33.020 160.575 ;
        RECT 28.090 160.390 33.020 160.530 ;
        RECT 28.090 160.345 28.380 160.390 ;
        RECT 29.950 160.345 30.240 160.390 ;
        RECT 32.730 160.345 33.020 160.390 ;
        RECT 37.745 160.345 38.035 160.575 ;
        RECT 43.365 160.530 43.655 160.575 ;
        RECT 46.485 160.530 46.775 160.575 ;
        RECT 48.375 160.530 48.665 160.575 ;
        RECT 43.365 160.390 48.665 160.530 ;
        RECT 43.365 160.345 43.655 160.390 ;
        RECT 46.485 160.345 46.775 160.390 ;
        RECT 48.375 160.345 48.665 160.390 ;
        RECT 54.380 160.250 54.520 160.685 ;
        RECT 57.140 160.575 57.280 161.070 ;
        RECT 58.905 161.025 59.195 161.070 ;
        RECT 61.650 161.210 61.970 161.270 ;
        RECT 62.585 161.210 62.875 161.255 ;
        RECT 66.710 161.210 67.030 161.270 ;
        RECT 61.650 161.070 67.030 161.210 ;
        RECT 61.650 161.010 61.970 161.070 ;
        RECT 62.585 161.025 62.875 161.070 ;
        RECT 66.710 161.010 67.030 161.070 ;
        RECT 71.325 161.210 71.615 161.255 ;
        RECT 71.770 161.210 72.090 161.270 ;
        RECT 71.325 161.070 72.090 161.210 ;
        RECT 71.325 161.025 71.615 161.070 ;
        RECT 71.770 161.010 72.090 161.070 ;
        RECT 81.430 161.010 81.750 161.270 ;
        RECT 85.660 161.255 85.800 161.410 ;
        RECT 88.790 161.350 89.110 161.410 ;
        RECT 92.880 161.550 93.170 161.595 ;
        RECT 95.230 161.550 95.550 161.610 ;
        RECT 96.140 161.550 96.430 161.595 ;
        RECT 92.880 161.410 96.430 161.550 ;
        RECT 92.880 161.365 93.170 161.410 ;
        RECT 95.230 161.350 95.550 161.410 ;
        RECT 96.140 161.365 96.430 161.410 ;
        RECT 97.060 161.550 97.350 161.595 ;
        RECT 98.920 161.550 99.210 161.595 ;
        RECT 97.060 161.410 99.210 161.550 ;
        RECT 97.060 161.365 97.350 161.410 ;
        RECT 98.920 161.365 99.210 161.410 ;
        RECT 85.585 161.025 85.875 161.255 ;
        RECT 86.950 161.010 87.270 161.270 ;
        RECT 94.740 161.210 95.030 161.255 ;
        RECT 97.060 161.210 97.275 161.365 ;
        RECT 94.740 161.070 97.275 161.210 ;
        RECT 98.005 161.210 98.295 161.255 ;
        RECT 100.380 161.210 100.520 161.705 ;
        RECT 109.490 161.690 109.810 161.750 ;
        RECT 98.005 161.070 100.520 161.210 ;
        RECT 94.740 161.025 95.030 161.070 ;
        RECT 98.005 161.025 98.295 161.070 ;
        RECT 101.210 161.010 101.530 161.270 ;
        RECT 106.270 161.010 106.590 161.270 ;
        RECT 115.930 161.210 116.250 161.270 ;
        RECT 119.610 161.210 119.930 161.270 ;
        RECT 115.930 161.070 119.930 161.210 ;
        RECT 115.930 161.010 116.250 161.070 ;
        RECT 119.610 161.010 119.930 161.070 ;
        RECT 57.510 160.870 57.830 160.930 ;
        RECT 61.205 160.870 61.495 160.915 ;
        RECT 57.510 160.730 61.495 160.870 ;
        RECT 57.510 160.670 57.830 160.730 ;
        RECT 61.205 160.685 61.495 160.730 ;
        RECT 79.590 160.870 79.910 160.930 ;
        RECT 80.065 160.870 80.355 160.915 ;
        RECT 83.270 160.870 83.590 160.930 ;
        RECT 79.590 160.730 83.590 160.870 ;
        RECT 79.590 160.670 79.910 160.730 ;
        RECT 80.065 160.685 80.355 160.730 ;
        RECT 83.270 160.670 83.590 160.730 ;
        RECT 99.830 160.670 100.150 160.930 ;
        RECT 117.310 160.870 117.630 160.930 ;
        RECT 118.245 160.870 118.535 160.915 ;
        RECT 117.310 160.730 118.535 160.870 ;
        RECT 117.310 160.670 117.630 160.730 ;
        RECT 118.245 160.685 118.535 160.730 ;
        RECT 57.065 160.345 57.355 160.575 ;
        RECT 84.190 160.530 84.510 160.590 ;
        RECT 90.875 160.530 91.165 160.575 ;
        RECT 93.850 160.530 94.170 160.590 ;
        RECT 84.190 160.390 94.170 160.530 ;
        RECT 84.190 160.330 84.510 160.390 ;
        RECT 90.875 160.345 91.165 160.390 ;
        RECT 93.850 160.330 94.170 160.390 ;
        RECT 94.740 160.530 95.030 160.575 ;
        RECT 97.520 160.530 97.810 160.575 ;
        RECT 99.380 160.530 99.670 160.575 ;
        RECT 94.740 160.390 99.670 160.530 ;
        RECT 94.740 160.345 95.030 160.390 ;
        RECT 97.520 160.345 97.810 160.390 ;
        RECT 99.380 160.345 99.670 160.390 ;
        RECT 104.430 160.530 104.750 160.590 ;
        RECT 106.270 160.530 106.590 160.590 ;
        RECT 104.430 160.390 106.590 160.530 ;
        RECT 104.430 160.330 104.750 160.390 ;
        RECT 106.270 160.330 106.590 160.390 ;
        RECT 35.890 160.190 36.210 160.250 ;
        RECT 36.595 160.190 36.885 160.235 ;
        RECT 35.890 160.050 36.885 160.190 ;
        RECT 35.890 159.990 36.210 160.050 ;
        RECT 36.595 160.005 36.885 160.050 ;
        RECT 52.450 159.990 52.770 160.250 ;
        RECT 54.290 160.190 54.610 160.250 ;
        RECT 66.265 160.190 66.555 160.235 ;
        RECT 54.290 160.050 66.555 160.190 ;
        RECT 54.290 159.990 54.610 160.050 ;
        RECT 66.265 160.005 66.555 160.050 ;
        RECT 84.650 160.190 84.970 160.250 ;
        RECT 85.125 160.190 85.415 160.235 ;
        RECT 84.650 160.050 85.415 160.190 ;
        RECT 84.650 159.990 84.970 160.050 ;
        RECT 85.125 160.005 85.415 160.050 ;
        RECT 87.885 160.190 88.175 160.235 ;
        RECT 88.330 160.190 88.650 160.250 ;
        RECT 87.885 160.050 88.650 160.190 ;
        RECT 87.885 160.005 88.175 160.050 ;
        RECT 88.330 159.990 88.650 160.050 ;
        RECT 94.310 160.190 94.630 160.250 ;
        RECT 106.730 160.190 107.050 160.250 ;
        RECT 94.310 160.050 107.050 160.190 ;
        RECT 94.310 159.990 94.630 160.050 ;
        RECT 106.730 159.990 107.050 160.050 ;
        RECT 14.660 159.370 127.820 159.850 ;
        RECT 19.790 158.970 20.110 159.230 ;
        RECT 31.290 159.170 31.610 159.230 ;
        RECT 32.225 159.170 32.515 159.215 ;
        RECT 31.290 159.030 32.515 159.170 ;
        RECT 31.290 158.970 31.610 159.030 ;
        RECT 32.225 158.985 32.515 159.030 ;
        RECT 36.825 159.170 37.115 159.215 ;
        RECT 38.650 159.170 38.970 159.230 ;
        RECT 36.825 159.030 38.970 159.170 ;
        RECT 36.825 158.985 37.115 159.030 ;
        RECT 38.650 158.970 38.970 159.030 ;
        RECT 49.690 158.970 50.010 159.230 ;
        RECT 52.005 159.170 52.295 159.215 ;
        RECT 52.910 159.170 53.230 159.230 ;
        RECT 70.865 159.170 71.155 159.215 ;
        RECT 79.130 159.170 79.450 159.230 ;
        RECT 94.310 159.170 94.630 159.230 ;
        RECT 52.005 159.030 53.230 159.170 ;
        RECT 52.005 158.985 52.295 159.030 ;
        RECT 52.910 158.970 53.230 159.030 ;
        RECT 54.380 159.030 79.450 159.170 ;
        RECT 20.265 158.645 20.555 158.875 ;
        RECT 53.830 158.830 54.150 158.890 ;
        RECT 34.140 158.690 54.150 158.830 ;
        RECT 18.885 158.150 19.175 158.195 ;
        RECT 20.340 158.150 20.480 158.645 ;
        RECT 22.090 158.490 22.410 158.550 ;
        RECT 34.140 158.535 34.280 158.690 ;
        RECT 23.485 158.490 23.775 158.535 ;
        RECT 34.065 158.490 34.355 158.535 ;
        RECT 44.170 158.490 44.490 158.550 ;
        RECT 47.020 158.535 47.160 158.690 ;
        RECT 53.830 158.630 54.150 158.690 ;
        RECT 22.090 158.350 34.355 158.490 ;
        RECT 22.090 158.290 22.410 158.350 ;
        RECT 23.485 158.305 23.775 158.350 ;
        RECT 34.065 158.305 34.355 158.350 ;
        RECT 41.960 158.350 44.490 158.490 ;
        RECT 18.885 158.010 20.480 158.150 ;
        RECT 20.710 158.150 21.030 158.210 ;
        RECT 31.750 158.150 32.070 158.210 ;
        RECT 20.710 158.010 32.070 158.150 ;
        RECT 18.885 157.965 19.175 158.010 ;
        RECT 20.710 157.950 21.030 158.010 ;
        RECT 31.750 157.950 32.070 158.010 ;
        RECT 40.950 158.150 41.270 158.210 ;
        RECT 41.960 158.195 42.100 158.350 ;
        RECT 44.170 158.290 44.490 158.350 ;
        RECT 46.945 158.305 47.235 158.535 ;
        RECT 51.070 158.490 51.390 158.550 ;
        RECT 54.380 158.490 54.520 159.030 ;
        RECT 70.865 158.985 71.155 159.030 ;
        RECT 79.130 158.970 79.450 159.030 ;
        RECT 79.680 159.030 94.630 159.170 ;
        RECT 54.865 158.830 55.155 158.875 ;
        RECT 57.985 158.830 58.275 158.875 ;
        RECT 59.875 158.830 60.165 158.875 ;
        RECT 54.865 158.690 60.165 158.830 ;
        RECT 54.865 158.645 55.155 158.690 ;
        RECT 57.985 158.645 58.275 158.690 ;
        RECT 59.875 158.645 60.165 158.690 ;
        RECT 61.190 158.830 61.510 158.890 ;
        RECT 69.025 158.830 69.315 158.875 ;
        RECT 79.680 158.830 79.820 159.030 ;
        RECT 94.310 158.970 94.630 159.030 ;
        RECT 94.785 159.170 95.075 159.215 ;
        RECT 95.230 159.170 95.550 159.230 ;
        RECT 94.785 159.030 95.550 159.170 ;
        RECT 94.785 158.985 95.075 159.030 ;
        RECT 95.230 158.970 95.550 159.030 ;
        RECT 61.190 158.690 79.820 158.830 ;
        RECT 85.080 158.830 85.370 158.875 ;
        RECT 87.860 158.830 88.150 158.875 ;
        RECT 89.720 158.830 90.010 158.875 ;
        RECT 85.080 158.690 90.010 158.830 ;
        RECT 61.190 158.630 61.510 158.690 ;
        RECT 69.025 158.645 69.315 158.690 ;
        RECT 85.080 158.645 85.370 158.690 ;
        RECT 87.860 158.645 88.150 158.690 ;
        RECT 89.720 158.645 90.010 158.690 ;
        RECT 102.130 158.830 102.450 158.890 ;
        RECT 102.130 158.690 117.080 158.830 ;
        RECT 102.130 158.630 102.450 158.690 ;
        RECT 68.550 158.490 68.870 158.550 ;
        RECT 86.030 158.490 86.350 158.550 ;
        RECT 51.070 158.350 54.520 158.490 ;
        RECT 65.880 158.350 70.160 158.490 ;
        RECT 51.070 158.290 51.390 158.350 ;
        RECT 41.425 158.150 41.715 158.195 ;
        RECT 40.950 158.010 41.715 158.150 ;
        RECT 40.950 157.950 41.270 158.010 ;
        RECT 41.425 157.965 41.715 158.010 ;
        RECT 41.885 157.965 42.175 158.195 ;
        RECT 42.345 157.965 42.635 158.195 ;
        RECT 34.970 157.810 35.290 157.870 ;
        RECT 42.420 157.810 42.560 157.965 ;
        RECT 43.250 157.950 43.570 158.210 ;
        RECT 34.970 157.670 42.560 157.810 ;
        RECT 52.450 157.810 52.770 157.870 ;
        RECT 53.785 157.855 54.075 158.170 ;
        RECT 54.865 158.150 55.155 158.195 ;
        RECT 58.445 158.150 58.735 158.195 ;
        RECT 60.280 158.150 60.570 158.195 ;
        RECT 54.865 158.010 60.570 158.150 ;
        RECT 54.865 157.965 55.155 158.010 ;
        RECT 58.445 157.965 58.735 158.010 ;
        RECT 60.280 157.965 60.570 158.010 ;
        RECT 60.730 157.950 61.050 158.210 ;
        RECT 65.880 158.195 66.020 158.350 ;
        RECT 68.550 158.290 68.870 158.350 ;
        RECT 65.805 157.965 66.095 158.195 ;
        RECT 67.645 158.150 67.935 158.195 ;
        RECT 68.105 158.150 68.395 158.195 ;
        RECT 69.470 158.150 69.790 158.210 ;
        RECT 70.020 158.195 70.160 158.350 ;
        RECT 86.030 158.350 88.100 158.490 ;
        RECT 86.030 158.290 86.350 158.350 ;
        RECT 67.645 158.010 69.790 158.150 ;
        RECT 67.645 157.965 67.935 158.010 ;
        RECT 68.105 157.965 68.395 158.010 ;
        RECT 69.470 157.950 69.790 158.010 ;
        RECT 69.945 157.965 70.235 158.195 ;
        RECT 85.080 158.150 85.370 158.195 ;
        RECT 87.960 158.150 88.100 158.350 ;
        RECT 88.330 158.290 88.650 158.550 ;
        RECT 104.430 158.490 104.750 158.550 ;
        RECT 110.870 158.490 111.190 158.550 ;
        RECT 116.940 158.535 117.080 158.690 ;
        RECT 104.430 158.350 106.500 158.490 ;
        RECT 104.430 158.290 104.750 158.350 ;
        RECT 90.185 158.150 90.475 158.195 ;
        RECT 85.080 158.010 87.615 158.150 ;
        RECT 87.960 158.010 90.475 158.150 ;
        RECT 85.080 157.965 85.370 158.010 ;
        RECT 53.485 157.810 54.075 157.855 ;
        RECT 56.725 157.810 57.375 157.855 ;
        RECT 52.450 157.670 57.375 157.810 ;
        RECT 34.970 157.610 35.290 157.670 ;
        RECT 52.450 157.610 52.770 157.670 ;
        RECT 53.485 157.625 53.775 157.670 ;
        RECT 56.725 157.625 57.375 157.670 ;
        RECT 59.350 157.610 59.670 157.870 ;
        RECT 81.430 157.855 81.750 157.870 ;
        RECT 64.960 157.670 67.400 157.810 ;
        RECT 21.630 157.470 21.950 157.530 ;
        RECT 22.105 157.470 22.395 157.515 ;
        RECT 21.630 157.330 22.395 157.470 ;
        RECT 21.630 157.270 21.950 157.330 ;
        RECT 22.105 157.285 22.395 157.330 ;
        RECT 22.550 157.470 22.870 157.530 ;
        RECT 31.290 157.470 31.610 157.530 ;
        RECT 22.550 157.330 31.610 157.470 ;
        RECT 22.550 157.270 22.870 157.330 ;
        RECT 31.290 157.270 31.610 157.330 ;
        RECT 34.525 157.470 34.815 157.515 ;
        RECT 35.890 157.470 36.210 157.530 ;
        RECT 36.810 157.470 37.130 157.530 ;
        RECT 34.525 157.330 37.130 157.470 ;
        RECT 34.525 157.285 34.815 157.330 ;
        RECT 35.890 157.270 36.210 157.330 ;
        RECT 36.810 157.270 37.130 157.330 ;
        RECT 40.030 157.270 40.350 157.530 ;
        RECT 43.710 157.470 44.030 157.530 ;
        RECT 47.405 157.470 47.695 157.515 ;
        RECT 43.710 157.330 47.695 157.470 ;
        RECT 43.710 157.270 44.030 157.330 ;
        RECT 47.405 157.285 47.695 157.330 ;
        RECT 47.865 157.470 48.155 157.515 ;
        RECT 49.230 157.470 49.550 157.530 ;
        RECT 47.865 157.330 49.550 157.470 ;
        RECT 47.865 157.285 48.155 157.330 ;
        RECT 49.230 157.270 49.550 157.330 ;
        RECT 50.150 157.470 50.470 157.530 ;
        RECT 64.960 157.515 65.100 157.670 ;
        RECT 64.885 157.470 65.175 157.515 ;
        RECT 50.150 157.330 65.175 157.470 ;
        RECT 50.150 157.270 50.470 157.330 ;
        RECT 64.885 157.285 65.175 157.330 ;
        RECT 66.710 157.270 67.030 157.530 ;
        RECT 67.260 157.470 67.400 157.670 ;
        RECT 81.215 157.625 81.750 157.855 ;
        RECT 83.220 157.810 83.510 157.855 ;
        RECT 84.650 157.810 84.970 157.870 ;
        RECT 87.400 157.855 87.615 158.010 ;
        RECT 90.185 157.965 90.475 158.010 ;
        RECT 95.230 157.950 95.550 158.210 ;
        RECT 106.360 158.195 106.500 158.350 ;
        RECT 106.820 158.350 111.190 158.490 ;
        RECT 106.820 158.210 106.960 158.350 ;
        RECT 110.870 158.290 111.190 158.350 ;
        RECT 116.865 158.305 117.155 158.535 ;
        RECT 105.825 157.965 106.115 158.195 ;
        RECT 106.285 157.965 106.575 158.195 ;
        RECT 86.480 157.810 86.770 157.855 ;
        RECT 83.220 157.670 86.770 157.810 ;
        RECT 83.220 157.625 83.510 157.670 ;
        RECT 81.430 157.610 81.750 157.625 ;
        RECT 84.650 157.610 84.970 157.670 ;
        RECT 86.480 157.625 86.770 157.670 ;
        RECT 87.400 157.810 87.690 157.855 ;
        RECT 89.260 157.810 89.550 157.855 ;
        RECT 103.050 157.810 103.370 157.870 ;
        RECT 105.900 157.810 106.040 157.965 ;
        RECT 106.730 157.950 107.050 158.210 ;
        RECT 107.665 158.150 107.955 158.195 ;
        RECT 109.490 158.150 109.810 158.210 ;
        RECT 107.665 158.010 109.810 158.150 ;
        RECT 107.665 157.965 107.955 158.010 ;
        RECT 109.490 157.950 109.810 158.010 ;
        RECT 115.930 157.950 116.250 158.210 ;
        RECT 111.790 157.810 112.110 157.870 ;
        RECT 87.400 157.670 89.550 157.810 ;
        RECT 87.400 157.625 87.690 157.670 ;
        RECT 89.260 157.625 89.550 157.670 ;
        RECT 99.460 157.670 112.110 157.810 ;
        RECT 99.460 157.530 99.600 157.670 ;
        RECT 103.050 157.610 103.370 157.670 ;
        RECT 111.790 157.610 112.110 157.670 ;
        RECT 99.370 157.470 99.690 157.530 ;
        RECT 67.260 157.330 99.690 157.470 ;
        RECT 99.370 157.270 99.690 157.330 ;
        RECT 103.510 157.470 103.830 157.530 ;
        RECT 104.445 157.470 104.735 157.515 ;
        RECT 103.510 157.330 104.735 157.470 ;
        RECT 103.510 157.270 103.830 157.330 ;
        RECT 104.445 157.285 104.735 157.330 ;
        RECT 14.660 156.650 127.820 157.130 ;
        RECT 36.810 156.450 37.130 156.510 ;
        RECT 37.730 156.450 38.050 156.510 ;
        RECT 52.925 156.450 53.215 156.495 ;
        RECT 36.810 156.310 53.215 156.450 ;
        RECT 36.810 156.250 37.130 156.310 ;
        RECT 37.730 156.250 38.050 156.310 ;
        RECT 52.925 156.265 53.215 156.310 ;
        RECT 57.525 156.450 57.815 156.495 ;
        RECT 59.350 156.450 59.670 156.510 ;
        RECT 57.525 156.310 59.670 156.450 ;
        RECT 57.525 156.265 57.815 156.310 ;
        RECT 59.350 156.250 59.670 156.310 ;
        RECT 86.505 156.450 86.795 156.495 ;
        RECT 86.950 156.450 87.270 156.510 ;
        RECT 86.505 156.310 87.270 156.450 ;
        RECT 86.505 156.265 86.795 156.310 ;
        RECT 86.950 156.250 87.270 156.310 ;
        RECT 94.310 156.450 94.630 156.510 ;
        RECT 104.430 156.450 104.750 156.510 ;
        RECT 109.030 156.450 109.350 156.510 ;
        RECT 94.310 156.310 112.940 156.450 ;
        RECT 94.310 156.250 94.630 156.310 ;
        RECT 19.330 156.155 19.650 156.170 ;
        RECT 19.280 156.110 19.650 156.155 ;
        RECT 22.540 156.110 22.830 156.155 ;
        RECT 19.280 155.970 22.830 156.110 ;
        RECT 19.280 155.925 19.650 155.970 ;
        RECT 22.540 155.925 22.830 155.970 ;
        RECT 23.460 156.110 23.750 156.155 ;
        RECT 25.320 156.110 25.610 156.155 ;
        RECT 23.460 155.970 25.610 156.110 ;
        RECT 23.460 155.925 23.750 155.970 ;
        RECT 25.320 155.925 25.610 155.970 ;
        RECT 42.330 156.110 42.650 156.170 ;
        RECT 61.190 156.110 61.510 156.170 ;
        RECT 42.330 155.970 61.510 156.110 ;
        RECT 19.330 155.910 19.650 155.925 ;
        RECT 21.140 155.770 21.430 155.815 ;
        RECT 23.460 155.770 23.675 155.925 ;
        RECT 42.330 155.910 42.650 155.970 ;
        RECT 61.190 155.910 61.510 155.970 ;
        RECT 66.710 156.110 67.030 156.170 ;
        RECT 79.590 156.110 79.910 156.170 ;
        RECT 81.430 156.110 81.750 156.170 ;
        RECT 84.205 156.110 84.495 156.155 ;
        RECT 66.710 155.970 80.740 156.110 ;
        RECT 66.710 155.910 67.030 155.970 ;
        RECT 79.590 155.910 79.910 155.970 ;
        RECT 21.140 155.630 23.675 155.770 ;
        RECT 52.465 155.770 52.755 155.815 ;
        RECT 52.910 155.770 53.230 155.830 ;
        RECT 56.605 155.770 56.895 155.815 ;
        RECT 52.465 155.630 53.230 155.770 ;
        RECT 21.140 155.585 21.430 155.630 ;
        RECT 52.465 155.585 52.755 155.630 ;
        RECT 52.910 155.570 53.230 155.630 ;
        RECT 54.840 155.630 56.895 155.770 ;
        RECT 24.390 155.230 24.710 155.490 ;
        RECT 26.230 155.430 26.550 155.490 ;
        RECT 28.990 155.430 29.310 155.490 ;
        RECT 26.230 155.290 29.310 155.430 ;
        RECT 26.230 155.230 26.550 155.290 ;
        RECT 28.990 155.230 29.310 155.290 ;
        RECT 31.750 155.430 32.070 155.490 ;
        RECT 51.530 155.430 51.850 155.490 ;
        RECT 31.750 155.290 51.850 155.430 ;
        RECT 31.750 155.230 32.070 155.290 ;
        RECT 51.530 155.230 51.850 155.290 ;
        RECT 52.005 155.430 52.295 155.475 ;
        RECT 53.830 155.430 54.150 155.490 ;
        RECT 52.005 155.290 54.150 155.430 ;
        RECT 52.005 155.245 52.295 155.290 ;
        RECT 53.830 155.230 54.150 155.290 ;
        RECT 21.140 155.090 21.430 155.135 ;
        RECT 23.920 155.090 24.210 155.135 ;
        RECT 25.780 155.090 26.070 155.135 ;
        RECT 21.140 154.950 26.070 155.090 ;
        RECT 21.140 154.905 21.430 154.950 ;
        RECT 23.920 154.905 24.210 154.950 ;
        RECT 25.780 154.905 26.070 154.950 ;
        RECT 39.570 155.090 39.890 155.150 ;
        RECT 50.150 155.090 50.470 155.150 ;
        RECT 54.840 155.135 54.980 155.630 ;
        RECT 56.605 155.585 56.895 155.630 ;
        RECT 67.645 155.770 67.935 155.815 ;
        RECT 68.105 155.770 68.395 155.815 ;
        RECT 67.645 155.630 68.395 155.770 ;
        RECT 67.645 155.585 67.935 155.630 ;
        RECT 68.105 155.585 68.395 155.630 ;
        RECT 69.945 155.770 70.235 155.815 ;
        RECT 70.390 155.770 70.710 155.830 ;
        RECT 69.945 155.630 70.710 155.770 ;
        RECT 69.945 155.585 70.235 155.630 ;
        RECT 68.180 155.430 68.320 155.585 ;
        RECT 70.390 155.570 70.710 155.630 ;
        RECT 71.770 155.770 72.090 155.830 ;
        RECT 73.165 155.770 73.455 155.815 ;
        RECT 74.530 155.770 74.850 155.830 ;
        RECT 71.770 155.630 74.850 155.770 ;
        RECT 71.770 155.570 72.090 155.630 ;
        RECT 73.165 155.585 73.455 155.630 ;
        RECT 74.530 155.570 74.850 155.630 ;
        RECT 79.130 155.770 79.450 155.830 ;
        RECT 80.600 155.815 80.740 155.970 ;
        RECT 81.060 155.970 84.495 156.110 ;
        RECT 81.060 155.815 81.200 155.970 ;
        RECT 81.430 155.910 81.750 155.970 ;
        RECT 84.205 155.925 84.495 155.970 ;
        RECT 80.065 155.770 80.355 155.815 ;
        RECT 79.130 155.630 80.355 155.770 ;
        RECT 79.130 155.570 79.450 155.630 ;
        RECT 80.065 155.585 80.355 155.630 ;
        RECT 80.525 155.585 80.815 155.815 ;
        RECT 80.985 155.585 81.275 155.815 ;
        RECT 81.905 155.585 82.195 155.815 ;
        RECT 82.350 155.770 82.670 155.830 ;
        RECT 84.665 155.770 84.955 155.815 ;
        RECT 82.350 155.630 84.955 155.770 ;
        RECT 71.860 155.430 72.000 155.570 ;
        RECT 68.180 155.290 72.000 155.430 ;
        RECT 72.230 155.430 72.550 155.490 ;
        RECT 81.980 155.430 82.120 155.585 ;
        RECT 82.350 155.570 82.670 155.630 ;
        RECT 84.280 155.490 84.420 155.630 ;
        RECT 84.665 155.585 84.955 155.630 ;
        RECT 99.370 155.570 99.690 155.830 ;
        RECT 99.920 155.815 100.060 156.310 ;
        RECT 104.430 156.250 104.750 156.310 ;
        RECT 103.050 156.110 103.370 156.170 ;
        RECT 105.900 156.110 106.040 156.310 ;
        RECT 109.030 156.250 109.350 156.310 ;
        RECT 111.790 156.110 112.110 156.170 ;
        RECT 103.050 155.970 104.660 156.110 ;
        RECT 103.050 155.910 103.370 155.970 ;
        RECT 99.845 155.585 100.135 155.815 ;
        RECT 100.305 155.770 100.595 155.815 ;
        RECT 100.750 155.770 101.070 155.830 ;
        RECT 100.305 155.630 101.070 155.770 ;
        RECT 100.305 155.585 100.595 155.630 ;
        RECT 100.750 155.570 101.070 155.630 ;
        RECT 101.225 155.770 101.515 155.815 ;
        RECT 102.590 155.770 102.910 155.830 ;
        RECT 101.225 155.630 102.910 155.770 ;
        RECT 104.520 155.785 104.660 155.970 ;
        RECT 105.440 155.970 106.040 156.110 ;
        RECT 108.660 155.970 112.110 156.110 ;
        RECT 105.440 155.815 105.580 155.970 ;
        RECT 108.660 155.830 108.800 155.970 ;
        RECT 111.790 155.910 112.110 155.970 ;
        RECT 104.905 155.785 105.195 155.815 ;
        RECT 104.520 155.645 105.195 155.785 ;
        RECT 101.225 155.585 101.515 155.630 ;
        RECT 72.230 155.290 82.120 155.430 ;
        RECT 72.230 155.230 72.550 155.290 ;
        RECT 39.570 154.950 50.470 155.090 ;
        RECT 39.570 154.890 39.890 154.950 ;
        RECT 50.150 154.890 50.470 154.950 ;
        RECT 54.765 154.905 55.055 155.135 ;
        RECT 66.725 155.090 67.015 155.135 ;
        RECT 68.550 155.090 68.870 155.150 ;
        RECT 81.980 155.090 82.120 155.290 ;
        RECT 83.270 155.230 83.590 155.490 ;
        RECT 84.190 155.230 84.510 155.490 ;
        RECT 101.300 155.430 101.440 155.585 ;
        RECT 102.590 155.570 102.910 155.630 ;
        RECT 104.905 155.585 105.195 155.645 ;
        RECT 105.350 155.585 105.640 155.815 ;
        RECT 105.825 155.785 106.115 155.815 ;
        RECT 106.270 155.785 106.590 155.830 ;
        RECT 105.825 155.645 106.590 155.785 ;
        RECT 105.825 155.585 106.115 155.645 ;
        RECT 106.270 155.570 106.590 155.645 ;
        RECT 106.730 155.570 107.050 155.830 ;
        RECT 108.570 155.570 108.890 155.830 ;
        RECT 109.030 155.570 109.350 155.830 ;
        RECT 109.505 155.770 109.795 155.815 ;
        RECT 109.950 155.770 110.270 155.830 ;
        RECT 109.505 155.630 110.270 155.770 ;
        RECT 109.505 155.585 109.795 155.630 ;
        RECT 109.950 155.570 110.270 155.630 ;
        RECT 110.425 155.585 110.715 155.815 ;
        RECT 111.880 155.770 112.020 155.910 ;
        RECT 112.800 155.815 112.940 156.310 ;
        RECT 115.485 156.110 115.775 156.155 ;
        RECT 117.885 156.110 118.175 156.155 ;
        RECT 121.125 156.110 121.775 156.155 ;
        RECT 115.485 155.970 121.775 156.110 ;
        RECT 115.485 155.925 115.775 155.970 ;
        RECT 117.885 155.925 118.475 155.970 ;
        RECT 121.125 155.925 121.775 155.970 ;
        RECT 123.765 156.110 124.055 156.155 ;
        RECT 124.210 156.110 124.530 156.170 ;
        RECT 123.765 155.970 124.530 156.110 ;
        RECT 123.765 155.925 124.055 155.970 ;
        RECT 112.265 155.770 112.555 155.815 ;
        RECT 111.880 155.630 112.555 155.770 ;
        RECT 112.265 155.585 112.555 155.630 ;
        RECT 112.725 155.585 113.015 155.815 ;
        RECT 97.620 155.290 101.440 155.430 ;
        RECT 84.650 155.090 84.970 155.150 ;
        RECT 66.725 154.950 81.660 155.090 ;
        RECT 81.980 154.950 84.970 155.090 ;
        RECT 66.725 154.905 67.015 154.950 ;
        RECT 68.550 154.890 68.870 154.950 ;
        RECT 17.275 154.750 17.565 154.795 ;
        RECT 21.630 154.750 21.950 154.810 ;
        RECT 17.275 154.610 21.950 154.750 ;
        RECT 17.275 154.565 17.565 154.610 ;
        RECT 21.630 154.550 21.950 154.610 ;
        RECT 45.550 154.750 45.870 154.810 ;
        RECT 47.390 154.750 47.710 154.810 ;
        RECT 45.550 154.610 47.710 154.750 ;
        RECT 45.550 154.550 45.870 154.610 ;
        RECT 47.390 154.550 47.710 154.610 ;
        RECT 51.530 154.750 51.850 154.810 ;
        RECT 53.370 154.750 53.690 154.810 ;
        RECT 57.050 154.750 57.370 154.810 ;
        RECT 51.530 154.610 57.370 154.750 ;
        RECT 51.530 154.550 51.850 154.610 ;
        RECT 53.370 154.550 53.690 154.610 ;
        RECT 57.050 154.550 57.370 154.610 ;
        RECT 67.630 154.750 67.950 154.810 ;
        RECT 69.025 154.750 69.315 154.795 ;
        RECT 67.630 154.610 69.315 154.750 ;
        RECT 67.630 154.550 67.950 154.610 ;
        RECT 69.025 154.565 69.315 154.610 ;
        RECT 69.470 154.750 69.790 154.810 ;
        RECT 70.865 154.750 71.155 154.795 ;
        RECT 69.470 154.610 71.155 154.750 ;
        RECT 69.470 154.550 69.790 154.610 ;
        RECT 70.865 154.565 71.155 154.610 ;
        RECT 72.230 154.550 72.550 154.810 ;
        RECT 78.685 154.750 78.975 154.795 ;
        RECT 80.970 154.750 81.290 154.810 ;
        RECT 78.685 154.610 81.290 154.750 ;
        RECT 81.520 154.750 81.660 154.950 ;
        RECT 84.650 154.890 84.970 154.950 ;
        RECT 97.620 154.750 97.760 155.290 ;
        RECT 109.950 155.090 110.270 155.150 ;
        RECT 110.500 155.090 110.640 155.585 ;
        RECT 113.170 155.570 113.490 155.830 ;
        RECT 114.105 155.585 114.395 155.815 ;
        RECT 115.025 155.770 115.315 155.815 ;
        RECT 117.310 155.770 117.630 155.830 ;
        RECT 115.025 155.630 117.630 155.770 ;
        RECT 115.025 155.585 115.315 155.630 ;
        RECT 114.180 155.090 114.320 155.585 ;
        RECT 117.310 155.570 117.630 155.630 ;
        RECT 118.185 155.610 118.475 155.925 ;
        RECT 124.210 155.910 124.530 155.970 ;
        RECT 119.265 155.770 119.555 155.815 ;
        RECT 122.845 155.770 123.135 155.815 ;
        RECT 124.680 155.770 124.970 155.815 ;
        RECT 119.265 155.630 124.970 155.770 ;
        RECT 119.265 155.585 119.555 155.630 ;
        RECT 122.845 155.585 123.135 155.630 ;
        RECT 124.680 155.585 124.970 155.630 ;
        RECT 125.145 155.430 125.435 155.475 ;
        RECT 125.590 155.430 125.910 155.490 ;
        RECT 125.145 155.290 125.910 155.430 ;
        RECT 125.145 155.245 125.435 155.290 ;
        RECT 125.590 155.230 125.910 155.290 ;
        RECT 109.950 154.950 114.320 155.090 ;
        RECT 119.265 155.090 119.555 155.135 ;
        RECT 122.385 155.090 122.675 155.135 ;
        RECT 124.275 155.090 124.565 155.135 ;
        RECT 119.265 154.950 124.565 155.090 ;
        RECT 109.950 154.890 110.270 154.950 ;
        RECT 119.265 154.905 119.555 154.950 ;
        RECT 122.385 154.905 122.675 154.950 ;
        RECT 124.275 154.905 124.565 154.950 ;
        RECT 81.520 154.610 97.760 154.750 ;
        RECT 78.685 154.565 78.975 154.610 ;
        RECT 80.970 154.550 81.290 154.610 ;
        RECT 97.990 154.550 98.310 154.810 ;
        RECT 103.050 154.750 103.370 154.810 ;
        RECT 103.525 154.750 103.815 154.795 ;
        RECT 103.050 154.610 103.815 154.750 ;
        RECT 103.050 154.550 103.370 154.610 ;
        RECT 103.525 154.565 103.815 154.610 ;
        RECT 107.205 154.750 107.495 154.795 ;
        RECT 109.490 154.750 109.810 154.810 ;
        RECT 107.205 154.610 109.810 154.750 ;
        RECT 107.205 154.565 107.495 154.610 ;
        RECT 109.490 154.550 109.810 154.610 ;
        RECT 110.870 154.550 111.190 154.810 ;
        RECT 116.390 154.550 116.710 154.810 ;
        RECT 14.660 153.930 127.820 154.410 ;
        RECT 44.170 153.730 44.490 153.790 ;
        RECT 47.850 153.730 48.170 153.790 ;
        RECT 50.610 153.730 50.930 153.790 ;
        RECT 52.450 153.730 52.770 153.790 ;
        RECT 66.710 153.730 67.030 153.790 ;
        RECT 44.170 153.590 67.030 153.730 ;
        RECT 44.170 153.530 44.490 153.590 ;
        RECT 47.850 153.530 48.170 153.590 ;
        RECT 50.610 153.530 50.930 153.590 ;
        RECT 52.450 153.530 52.770 153.590 ;
        RECT 66.710 153.530 67.030 153.590 ;
        RECT 70.850 153.730 71.170 153.790 ;
        RECT 73.150 153.730 73.470 153.790 ;
        RECT 70.850 153.590 73.470 153.730 ;
        RECT 70.850 153.530 71.170 153.590 ;
        RECT 73.150 153.530 73.470 153.590 ;
        RECT 79.590 153.730 79.910 153.790 ;
        RECT 104.430 153.730 104.750 153.790 ;
        RECT 110.870 153.730 111.190 153.790 ;
        RECT 79.590 153.590 83.500 153.730 ;
        RECT 79.590 153.530 79.910 153.590 ;
        RECT 22.090 153.390 22.410 153.450 ;
        RECT 39.570 153.390 39.890 153.450 ;
        RECT 48.310 153.390 48.630 153.450 ;
        RECT 21.260 153.250 27.380 153.390 ;
        RECT 21.260 153.095 21.400 153.250 ;
        RECT 22.090 153.190 22.410 153.250 ;
        RECT 27.240 153.095 27.380 153.250 ;
        RECT 36.440 153.250 39.890 153.390 ;
        RECT 21.185 152.865 21.475 153.095 ;
        RECT 27.165 152.865 27.455 153.095 ;
        RECT 35.430 153.050 35.750 153.110 ;
        RECT 28.620 152.910 35.750 153.050 ;
        RECT 28.620 152.755 28.760 152.910 ;
        RECT 35.430 152.850 35.750 152.910 ;
        RECT 28.545 152.525 28.835 152.755 ;
        RECT 31.305 152.525 31.595 152.755 ;
        RECT 22.090 152.370 22.410 152.430 ;
        RECT 31.380 152.370 31.520 152.525 ;
        RECT 32.210 152.510 32.530 152.770 ;
        RECT 32.670 152.510 32.990 152.770 ;
        RECT 36.440 152.755 36.580 153.250 ;
        RECT 39.570 153.190 39.890 153.250 ;
        RECT 44.720 153.250 48.630 153.390 ;
        RECT 40.950 153.050 41.270 153.110 ;
        RECT 43.250 153.050 43.570 153.110 ;
        RECT 44.720 153.050 44.860 153.250 ;
        RECT 48.310 153.190 48.630 153.250 ;
        RECT 63.965 153.205 64.255 153.435 ;
        RECT 40.950 152.910 44.860 153.050 ;
        RECT 40.950 152.850 41.270 152.910 ;
        RECT 43.250 152.850 43.570 152.910 ;
        RECT 33.145 152.710 33.435 152.755 ;
        RECT 36.365 152.710 36.655 152.755 ;
        RECT 33.145 152.570 36.655 152.710 ;
        RECT 33.145 152.525 33.435 152.570 ;
        RECT 36.365 152.525 36.655 152.570 ;
        RECT 36.810 152.510 37.130 152.770 ;
        RECT 37.285 152.695 37.575 152.740 ;
        RECT 37.730 152.695 38.050 152.770 ;
        RECT 37.285 152.555 38.050 152.695 ;
        RECT 37.285 152.510 37.575 152.555 ;
        RECT 37.730 152.510 38.050 152.555 ;
        RECT 38.190 152.510 38.510 152.770 ;
        RECT 42.790 152.510 43.110 152.770 ;
        RECT 43.710 152.510 44.030 152.770 ;
        RECT 44.170 152.510 44.490 152.770 ;
        RECT 44.720 152.755 44.860 152.910 ;
        RECT 46.010 153.050 46.330 153.110 ;
        RECT 50.625 153.050 50.915 153.095 ;
        RECT 46.010 152.910 50.915 153.050 ;
        RECT 64.040 153.050 64.180 153.205 ;
        RECT 64.410 153.050 64.730 153.110 ;
        RECT 70.940 153.050 71.080 153.530 ;
        RECT 79.130 153.390 79.450 153.450 ;
        RECT 81.430 153.390 81.750 153.450 ;
        RECT 79.130 153.250 82.580 153.390 ;
        RECT 79.130 153.190 79.450 153.250 ;
        RECT 81.430 153.190 81.750 153.250 ;
        RECT 73.610 153.050 73.930 153.110 ;
        RECT 74.085 153.050 74.375 153.095 ;
        RECT 64.040 152.910 64.730 153.050 ;
        RECT 46.010 152.850 46.330 152.910 ;
        RECT 50.625 152.865 50.915 152.910 ;
        RECT 64.410 152.850 64.730 152.910 ;
        RECT 65.420 152.910 71.080 153.050 ;
        RECT 71.860 152.910 73.380 153.050 ;
        RECT 44.645 152.525 44.935 152.755 ;
        RECT 46.485 152.525 46.775 152.755 ;
        RECT 46.930 152.710 47.250 152.770 ;
        RECT 47.405 152.710 47.695 152.755 ;
        RECT 46.930 152.570 47.695 152.710 ;
        RECT 33.590 152.370 33.910 152.430 ;
        RECT 22.090 152.230 27.380 152.370 ;
        RECT 31.380 152.230 36.810 152.370 ;
        RECT 22.090 152.170 22.410 152.230 ;
        RECT 21.630 151.830 21.950 152.090 ;
        RECT 23.930 151.830 24.250 152.090 ;
        RECT 27.240 152.030 27.380 152.230 ;
        RECT 33.590 152.170 33.910 152.230 ;
        RECT 28.085 152.030 28.375 152.075 ;
        RECT 28.530 152.030 28.850 152.090 ;
        RECT 27.240 151.890 28.850 152.030 ;
        RECT 28.085 151.845 28.375 151.890 ;
        RECT 28.530 151.830 28.850 151.890 ;
        RECT 30.370 151.830 30.690 152.090 ;
        RECT 34.050 152.030 34.370 152.090 ;
        RECT 34.525 152.030 34.815 152.075 ;
        RECT 34.050 151.890 34.815 152.030 ;
        RECT 34.050 151.830 34.370 151.890 ;
        RECT 34.525 151.845 34.815 151.890 ;
        RECT 34.970 151.830 35.290 152.090 ;
        RECT 36.670 152.030 36.810 152.230 ;
        RECT 37.730 152.030 38.050 152.090 ;
        RECT 36.670 151.890 38.050 152.030 ;
        RECT 37.730 151.830 38.050 151.890 ;
        RECT 43.710 152.030 44.030 152.090 ;
        RECT 44.260 152.030 44.400 152.510 ;
        RECT 46.560 152.370 46.700 152.525 ;
        RECT 46.930 152.510 47.250 152.570 ;
        RECT 47.405 152.525 47.695 152.570 ;
        RECT 47.850 152.510 48.170 152.770 ;
        RECT 48.310 152.710 48.630 152.770 ;
        RECT 51.070 152.710 51.390 152.770 ;
        RECT 52.005 152.710 52.295 152.755 ;
        RECT 48.310 152.570 52.295 152.710 ;
        RECT 48.310 152.510 48.630 152.570 ;
        RECT 51.070 152.510 51.390 152.570 ;
        RECT 52.005 152.525 52.295 152.570 ;
        RECT 52.450 152.510 52.770 152.770 ;
        RECT 52.910 152.510 53.230 152.770 ;
        RECT 53.830 152.510 54.150 152.770 ;
        RECT 62.125 152.710 62.415 152.755 ;
        RECT 63.950 152.710 64.270 152.770 ;
        RECT 62.125 152.570 64.270 152.710 ;
        RECT 62.125 152.525 62.415 152.570 ;
        RECT 63.950 152.510 64.270 152.570 ;
        RECT 64.885 152.720 65.175 152.755 ;
        RECT 65.420 152.720 65.560 152.910 ;
        RECT 64.885 152.580 65.560 152.720 ;
        RECT 64.885 152.525 65.175 152.580 ;
        RECT 66.710 152.510 67.030 152.770 ;
        RECT 67.185 152.525 67.475 152.755 ;
        RECT 67.645 152.525 67.935 152.755 ;
        RECT 53.920 152.370 54.060 152.510 ;
        RECT 46.560 152.230 54.060 152.370 ;
        RECT 64.410 152.370 64.730 152.430 ;
        RECT 67.260 152.370 67.400 152.525 ;
        RECT 64.410 152.230 67.400 152.370 ;
        RECT 67.720 152.370 67.860 152.525 ;
        RECT 68.550 152.510 68.870 152.770 ;
        RECT 70.390 152.710 70.710 152.770 ;
        RECT 71.860 152.755 72.000 152.910 ;
        RECT 70.390 152.570 71.310 152.710 ;
        RECT 70.390 152.510 70.710 152.570 ;
        RECT 69.930 152.370 70.250 152.430 ;
        RECT 67.720 152.230 70.250 152.370 ;
        RECT 71.170 152.370 71.310 152.570 ;
        RECT 71.785 152.525 72.075 152.755 ;
        RECT 72.705 152.525 72.995 152.755 ;
        RECT 73.240 152.710 73.380 152.910 ;
        RECT 73.610 152.910 74.375 153.050 ;
        RECT 73.610 152.850 73.930 152.910 ;
        RECT 74.085 152.865 74.375 152.910 ;
        RECT 74.530 152.850 74.850 153.110 ;
        RECT 81.890 153.050 82.210 153.110 ;
        RECT 80.140 152.910 82.210 153.050 ;
        RECT 73.240 152.570 75.220 152.710 ;
        RECT 72.780 152.370 72.920 152.525 ;
        RECT 71.170 152.230 72.920 152.370 ;
        RECT 64.410 152.170 64.730 152.230 ;
        RECT 69.930 152.170 70.250 152.230 ;
        RECT 75.080 152.090 75.220 152.570 ;
        RECT 79.130 152.510 79.450 152.770 ;
        RECT 79.590 152.510 79.910 152.770 ;
        RECT 80.140 152.755 80.280 152.910 ;
        RECT 81.890 152.850 82.210 152.910 ;
        RECT 80.065 152.525 80.355 152.755 ;
        RECT 80.985 152.710 81.275 152.755 ;
        RECT 82.440 152.710 82.580 153.250 ;
        RECT 83.360 152.755 83.500 153.590 ;
        RECT 104.430 153.590 111.190 153.730 ;
        RECT 104.430 153.530 104.750 153.590 ;
        RECT 110.870 153.530 111.190 153.590 ;
        RECT 123.765 153.730 124.055 153.775 ;
        RECT 124.210 153.730 124.530 153.790 ;
        RECT 123.765 153.590 124.530 153.730 ;
        RECT 123.765 153.545 124.055 153.590 ;
        RECT 124.210 153.530 124.530 153.590 ;
        RECT 102.130 153.390 102.450 153.450 ;
        RECT 92.100 153.250 102.450 153.390 ;
        RECT 90.630 153.050 90.950 153.110 ;
        RECT 92.100 153.050 92.240 153.250 ;
        RECT 102.130 153.190 102.450 153.250 ;
        RECT 109.030 153.190 109.350 153.450 ;
        RECT 117.310 153.390 117.630 153.450 ;
        RECT 117.310 153.250 119.840 153.390 ;
        RECT 117.310 153.190 117.630 153.250 ;
        RECT 90.630 152.910 92.240 153.050 ;
        RECT 109.120 153.050 109.260 153.190 ;
        RECT 115.470 153.050 115.790 153.110 ;
        RECT 109.120 152.910 109.720 153.050 ;
        RECT 90.630 152.850 90.950 152.910 ;
        RECT 82.825 152.710 83.115 152.755 ;
        RECT 80.985 152.570 82.120 152.710 ;
        RECT 82.440 152.570 83.115 152.710 ;
        RECT 80.985 152.525 81.275 152.570 ;
        RECT 43.710 151.890 44.400 152.030 ;
        RECT 45.550 152.030 45.870 152.090 ;
        RECT 46.025 152.030 46.315 152.075 ;
        RECT 45.550 151.890 46.315 152.030 ;
        RECT 43.710 151.830 44.030 151.890 ;
        RECT 45.550 151.830 45.870 151.890 ;
        RECT 46.025 151.845 46.315 151.890 ;
        RECT 49.705 152.030 49.995 152.075 ;
        RECT 50.150 152.030 50.470 152.090 ;
        RECT 49.705 151.890 50.470 152.030 ;
        RECT 49.705 151.845 49.995 151.890 ;
        RECT 50.150 151.830 50.470 151.890 ;
        RECT 62.585 152.030 62.875 152.075 ;
        RECT 63.950 152.030 64.270 152.090 ;
        RECT 62.585 151.890 64.270 152.030 ;
        RECT 62.585 151.845 62.875 151.890 ;
        RECT 63.950 151.830 64.270 151.890 ;
        RECT 65.330 151.830 65.650 152.090 ;
        RECT 69.010 152.030 69.330 152.090 ;
        RECT 70.405 152.030 70.695 152.075 ;
        RECT 69.010 151.890 70.695 152.030 ;
        RECT 69.010 151.830 69.330 151.890 ;
        RECT 70.405 151.845 70.695 151.890 ;
        RECT 74.990 151.830 75.310 152.090 ;
        RECT 76.370 152.030 76.690 152.090 ;
        RECT 77.765 152.030 78.055 152.075 ;
        RECT 76.370 151.890 78.055 152.030 ;
        RECT 76.370 151.830 76.690 151.890 ;
        RECT 77.765 151.845 78.055 151.890 ;
        RECT 79.130 152.030 79.450 152.090 ;
        RECT 81.445 152.030 81.735 152.075 ;
        RECT 79.130 151.890 81.735 152.030 ;
        RECT 81.980 152.030 82.120 152.570 ;
        RECT 82.825 152.525 83.115 152.570 ;
        RECT 83.285 152.525 83.575 152.755 ;
        RECT 83.730 152.510 84.050 152.770 ;
        RECT 84.650 152.510 84.970 152.770 ;
        RECT 95.230 152.710 95.550 152.770 ;
        RECT 96.165 152.710 96.455 152.755 ;
        RECT 95.230 152.570 96.455 152.710 ;
        RECT 95.230 152.510 95.550 152.570 ;
        RECT 96.165 152.525 96.455 152.570 ;
        RECT 96.610 152.710 96.930 152.770 ;
        RECT 97.545 152.710 97.835 152.755 ;
        RECT 96.610 152.570 97.835 152.710 ;
        RECT 96.610 152.510 96.930 152.570 ;
        RECT 97.545 152.525 97.835 152.570 ;
        RECT 108.570 152.710 108.890 152.770 ;
        RECT 109.580 152.755 109.720 152.910 ;
        RECT 110.040 152.910 115.790 153.050 ;
        RECT 110.040 152.755 110.180 152.910 ;
        RECT 115.470 152.850 115.790 152.910 ;
        RECT 115.945 152.865 116.235 153.095 ;
        RECT 109.045 152.710 109.335 152.755 ;
        RECT 108.570 152.570 109.335 152.710 ;
        RECT 108.570 152.510 108.890 152.570 ;
        RECT 109.045 152.525 109.335 152.570 ;
        RECT 109.505 152.525 109.795 152.755 ;
        RECT 109.965 152.525 110.255 152.755 ;
        RECT 110.410 152.710 110.730 152.770 ;
        RECT 110.885 152.710 111.175 152.755 ;
        RECT 110.410 152.570 111.175 152.710 ;
        RECT 116.020 152.710 116.160 152.865 ;
        RECT 117.310 152.710 117.630 152.770 ;
        RECT 119.700 152.755 119.840 153.250 ;
        RECT 116.020 152.570 117.630 152.710 ;
        RECT 110.410 152.510 110.730 152.570 ;
        RECT 110.885 152.525 111.175 152.570 ;
        RECT 117.310 152.510 117.630 152.570 ;
        RECT 119.625 152.710 119.915 152.755 ;
        RECT 120.990 152.710 121.310 152.770 ;
        RECT 119.625 152.570 121.310 152.710 ;
        RECT 119.625 152.525 119.915 152.570 ;
        RECT 120.990 152.510 121.310 152.570 ;
        RECT 121.450 152.510 121.770 152.770 ;
        RECT 122.845 152.525 123.135 152.755 ;
        RECT 122.920 152.370 123.060 152.525 ;
        RECT 119.470 152.230 123.060 152.370 ;
        RECT 84.650 152.030 84.970 152.090 ;
        RECT 81.980 151.890 84.970 152.030 ;
        RECT 79.130 151.830 79.450 151.890 ;
        RECT 81.445 151.845 81.735 151.890 ;
        RECT 84.650 151.830 84.970 151.890 ;
        RECT 95.705 152.030 95.995 152.075 ;
        RECT 96.150 152.030 96.470 152.090 ;
        RECT 95.705 151.890 96.470 152.030 ;
        RECT 95.705 151.845 95.995 151.890 ;
        RECT 96.150 151.830 96.470 151.890 ;
        RECT 98.450 151.830 98.770 152.090 ;
        RECT 107.665 152.030 107.955 152.075 ;
        RECT 109.030 152.030 109.350 152.090 ;
        RECT 107.665 151.890 109.350 152.030 ;
        RECT 107.665 151.845 107.955 151.890 ;
        RECT 109.030 151.830 109.350 151.890 ;
        RECT 116.390 151.830 116.710 152.090 ;
        RECT 116.850 151.830 117.170 152.090 ;
        RECT 118.705 152.030 118.995 152.075 ;
        RECT 119.470 152.030 119.610 152.230 ;
        RECT 118.705 151.890 119.610 152.030 ;
        RECT 118.705 151.845 118.995 151.890 ;
        RECT 120.070 151.830 120.390 152.090 ;
        RECT 122.385 152.030 122.675 152.075 ;
        RECT 123.750 152.030 124.070 152.090 ;
        RECT 122.385 151.890 124.070 152.030 ;
        RECT 122.385 151.845 122.675 151.890 ;
        RECT 123.750 151.830 124.070 151.890 ;
        RECT 14.660 151.210 127.820 151.690 ;
        RECT 17.505 151.010 17.795 151.055 ;
        RECT 19.330 151.010 19.650 151.070 ;
        RECT 17.505 150.870 19.650 151.010 ;
        RECT 17.505 150.825 17.795 150.870 ;
        RECT 19.330 150.810 19.650 150.870 ;
        RECT 32.670 151.010 32.990 151.070 ;
        RECT 36.810 151.010 37.130 151.070 ;
        RECT 32.670 150.870 37.130 151.010 ;
        RECT 32.670 150.810 32.990 150.870 ;
        RECT 36.810 150.810 37.130 150.870 ;
        RECT 40.490 151.010 40.810 151.070 ;
        RECT 41.870 151.010 42.190 151.070 ;
        RECT 53.830 151.010 54.150 151.070 ;
        RECT 72.230 151.010 72.550 151.070 ;
        RECT 40.490 150.870 42.190 151.010 ;
        RECT 40.490 150.810 40.810 150.870 ;
        RECT 41.870 150.810 42.190 150.870 ;
        RECT 45.640 150.870 72.550 151.010 ;
        RECT 18.885 150.670 19.175 150.715 ;
        RECT 22.040 150.670 22.330 150.715 ;
        RECT 25.300 150.670 25.590 150.715 ;
        RECT 18.885 150.530 25.590 150.670 ;
        RECT 18.885 150.485 19.175 150.530 ;
        RECT 22.040 150.485 22.330 150.530 ;
        RECT 25.300 150.485 25.590 150.530 ;
        RECT 26.220 150.670 26.510 150.715 ;
        RECT 28.080 150.670 28.370 150.715 ;
        RECT 26.220 150.530 28.370 150.670 ;
        RECT 26.220 150.485 26.510 150.530 ;
        RECT 28.080 150.485 28.370 150.530 ;
        RECT 28.530 150.670 28.850 150.730 ;
        RECT 42.790 150.670 43.110 150.730 ;
        RECT 45.640 150.670 45.780 150.870 ;
        RECT 28.530 150.530 41.180 150.670 ;
        RECT 17.965 150.330 18.255 150.375 ;
        RECT 18.425 150.330 18.715 150.375 ;
        RECT 20.710 150.330 21.030 150.390 ;
        RECT 17.965 150.190 21.030 150.330 ;
        RECT 17.965 150.145 18.255 150.190 ;
        RECT 18.425 150.145 18.715 150.190 ;
        RECT 20.710 150.130 21.030 150.190 ;
        RECT 23.900 150.330 24.190 150.375 ;
        RECT 26.220 150.330 26.435 150.485 ;
        RECT 28.530 150.470 28.850 150.530 ;
        RECT 23.900 150.190 26.435 150.330 ;
        RECT 23.900 150.145 24.190 150.190 ;
        RECT 28.990 150.130 29.310 150.390 ;
        RECT 30.370 150.130 30.690 150.390 ;
        RECT 33.590 150.130 33.910 150.390 ;
        RECT 34.525 150.145 34.815 150.375 ;
        RECT 34.985 150.145 35.275 150.375 ;
        RECT 35.445 150.330 35.735 150.375 ;
        RECT 39.570 150.330 39.890 150.390 ;
        RECT 41.040 150.375 41.180 150.530 ;
        RECT 41.960 150.530 45.780 150.670 ;
        RECT 41.960 150.375 42.100 150.530 ;
        RECT 42.790 150.470 43.110 150.530 ;
        RECT 40.045 150.330 40.335 150.375 ;
        RECT 35.445 150.190 40.335 150.330 ;
        RECT 35.445 150.145 35.735 150.190 ;
        RECT 20.035 149.990 20.325 150.035 ;
        RECT 22.090 149.990 22.410 150.050 ;
        RECT 20.035 149.850 22.410 149.990 ;
        RECT 20.035 149.805 20.325 149.850 ;
        RECT 22.090 149.790 22.410 149.850 ;
        RECT 27.165 149.990 27.455 150.035 ;
        RECT 27.165 149.850 29.680 149.990 ;
        RECT 27.165 149.805 27.455 149.850 ;
        RECT 29.540 149.695 29.680 149.850 ;
        RECT 23.900 149.650 24.190 149.695 ;
        RECT 26.680 149.650 26.970 149.695 ;
        RECT 28.540 149.650 28.830 149.695 ;
        RECT 23.900 149.510 28.830 149.650 ;
        RECT 23.900 149.465 24.190 149.510 ;
        RECT 26.680 149.465 26.970 149.510 ;
        RECT 28.540 149.465 28.830 149.510 ;
        RECT 29.465 149.465 29.755 149.695 ;
        RECT 21.630 149.310 21.950 149.370 ;
        RECT 34.600 149.310 34.740 150.145 ;
        RECT 35.060 149.990 35.200 150.145 ;
        RECT 39.570 150.130 39.890 150.190 ;
        RECT 40.045 150.145 40.335 150.190 ;
        RECT 40.505 150.145 40.795 150.375 ;
        RECT 40.965 150.145 41.255 150.375 ;
        RECT 41.885 150.145 42.175 150.375 ;
        RECT 36.810 149.990 37.130 150.050 ;
        RECT 40.580 149.990 40.720 150.145 ;
        RECT 42.330 150.130 42.650 150.390 ;
        RECT 43.250 150.330 43.570 150.390 ;
        RECT 45.640 150.375 45.780 150.530 ;
        RECT 49.230 150.670 49.550 150.730 ;
        RECT 49.230 150.530 51.300 150.670 ;
        RECT 49.230 150.470 49.550 150.530 ;
        RECT 43.725 150.330 44.015 150.375 ;
        RECT 43.250 150.190 44.015 150.330 ;
        RECT 43.250 150.130 43.570 150.190 ;
        RECT 43.725 150.145 44.015 150.190 ;
        RECT 44.185 150.145 44.475 150.375 ;
        RECT 44.645 150.330 44.935 150.375 ;
        RECT 44.645 150.190 45.320 150.330 ;
        RECT 44.645 150.145 44.935 150.190 ;
        RECT 42.420 149.990 42.560 150.130 ;
        RECT 44.260 149.990 44.400 150.145 ;
        RECT 35.060 149.850 42.560 149.990 ;
        RECT 43.800 149.850 44.400 149.990 ;
        RECT 36.810 149.790 37.130 149.850 ;
        RECT 43.800 149.710 43.940 149.850 ;
        RECT 35.430 149.650 35.750 149.710 ;
        RECT 35.430 149.510 43.020 149.650 ;
        RECT 35.430 149.450 35.750 149.510 ;
        RECT 21.630 149.170 34.740 149.310 ;
        RECT 35.890 149.310 36.210 149.370 ;
        RECT 36.825 149.310 37.115 149.355 ;
        RECT 35.890 149.170 37.115 149.310 ;
        RECT 21.630 149.110 21.950 149.170 ;
        RECT 35.890 149.110 36.210 149.170 ;
        RECT 36.825 149.125 37.115 149.170 ;
        RECT 38.650 149.110 38.970 149.370 ;
        RECT 41.870 149.310 42.190 149.370 ;
        RECT 42.345 149.310 42.635 149.355 ;
        RECT 41.870 149.170 42.635 149.310 ;
        RECT 42.880 149.310 43.020 149.510 ;
        RECT 43.710 149.450 44.030 149.710 ;
        RECT 45.180 149.310 45.320 150.190 ;
        RECT 45.565 150.145 45.855 150.375 ;
        RECT 50.165 150.145 50.455 150.375 ;
        RECT 50.240 149.650 50.380 150.145 ;
        RECT 50.610 150.130 50.930 150.390 ;
        RECT 51.160 150.375 51.300 150.530 ;
        RECT 51.085 150.145 51.375 150.375 ;
        RECT 52.005 150.330 52.295 150.375 ;
        RECT 52.540 150.330 52.680 150.870 ;
        RECT 53.830 150.810 54.150 150.870 ;
        RECT 72.230 150.810 72.550 150.870 ;
        RECT 78.225 151.010 78.515 151.055 ;
        RECT 85.110 151.010 85.430 151.070 ;
        RECT 78.225 150.870 85.430 151.010 ;
        RECT 78.225 150.825 78.515 150.870 ;
        RECT 85.110 150.810 85.430 150.870 ;
        RECT 92.485 151.010 92.775 151.055 ;
        RECT 95.690 151.010 96.010 151.070 ;
        RECT 92.485 150.870 96.010 151.010 ;
        RECT 92.485 150.825 92.775 150.870 ;
        RECT 95.690 150.810 96.010 150.870 ;
        RECT 103.525 151.010 103.815 151.055 ;
        RECT 120.530 151.010 120.850 151.070 ;
        RECT 103.525 150.870 108.340 151.010 ;
        RECT 103.525 150.825 103.815 150.870 ;
        RECT 66.710 150.670 67.030 150.730 ;
        RECT 60.820 150.530 67.030 150.670 ;
        RECT 60.820 150.375 60.960 150.530 ;
        RECT 66.710 150.470 67.030 150.530 ;
        RECT 70.390 150.670 70.710 150.730 ;
        RECT 74.990 150.670 75.310 150.730 ;
        RECT 76.845 150.670 77.135 150.715 ;
        RECT 70.390 150.530 72.920 150.670 ;
        RECT 70.390 150.470 70.710 150.530 ;
        RECT 52.005 150.190 52.680 150.330 ;
        RECT 52.005 150.145 52.295 150.190 ;
        RECT 60.745 150.145 61.035 150.375 ;
        RECT 61.205 150.145 61.495 150.375 ;
        RECT 51.070 149.650 51.390 149.710 ;
        RECT 50.240 149.510 51.390 149.650 ;
        RECT 61.280 149.650 61.420 150.145 ;
        RECT 61.650 150.130 61.970 150.390 ;
        RECT 62.585 150.330 62.875 150.375 ;
        RECT 64.870 150.330 65.190 150.390 ;
        RECT 65.790 150.330 66.110 150.390 ;
        RECT 62.585 150.190 66.110 150.330 ;
        RECT 62.585 150.145 62.875 150.190 ;
        RECT 64.870 150.130 65.190 150.190 ;
        RECT 65.790 150.130 66.110 150.190 ;
        RECT 72.230 150.130 72.550 150.390 ;
        RECT 72.780 150.375 72.920 150.530 ;
        RECT 74.990 150.530 77.135 150.670 ;
        RECT 74.990 150.470 75.310 150.530 ;
        RECT 76.845 150.485 77.135 150.530 ;
        RECT 79.590 150.670 79.910 150.730 ;
        RECT 93.965 150.670 94.255 150.715 ;
        RECT 96.150 150.670 96.470 150.730 ;
        RECT 97.205 150.670 97.855 150.715 ;
        RECT 79.590 150.530 81.660 150.670 ;
        RECT 79.590 150.470 79.910 150.530 ;
        RECT 72.705 150.145 72.995 150.375 ;
        RECT 73.150 150.330 73.470 150.390 ;
        RECT 81.520 150.375 81.660 150.530 ;
        RECT 93.965 150.530 97.855 150.670 ;
        RECT 93.965 150.485 94.555 150.530 ;
        RECT 74.545 150.330 74.835 150.375 ;
        RECT 73.150 150.190 74.835 150.330 ;
        RECT 73.150 150.130 73.470 150.190 ;
        RECT 74.545 150.145 74.835 150.190 ;
        RECT 80.985 150.145 81.275 150.375 ;
        RECT 81.445 150.145 81.735 150.375 ;
        RECT 81.905 150.330 82.195 150.375 ;
        RECT 82.350 150.330 82.670 150.390 ;
        RECT 81.905 150.190 82.670 150.330 ;
        RECT 81.905 150.145 82.195 150.190 ;
        RECT 81.060 149.990 81.200 150.145 ;
        RECT 82.350 150.130 82.670 150.190 ;
        RECT 82.825 150.330 83.115 150.375 ;
        RECT 84.650 150.330 84.970 150.390 ;
        RECT 82.825 150.190 84.970 150.330 ;
        RECT 82.825 150.145 83.115 150.190 ;
        RECT 84.650 150.130 84.970 150.190 ;
        RECT 90.630 150.130 90.950 150.390 ;
        RECT 91.090 150.130 91.410 150.390 ;
        RECT 94.265 150.170 94.555 150.485 ;
        RECT 96.150 150.470 96.470 150.530 ;
        RECT 97.205 150.485 97.855 150.530 ;
        RECT 98.450 150.670 98.770 150.730 ;
        RECT 99.845 150.670 100.135 150.715 ;
        RECT 98.450 150.530 100.135 150.670 ;
        RECT 108.200 150.670 108.340 150.870 ;
        RECT 117.400 150.870 120.850 151.010 ;
        RECT 117.400 150.670 117.540 150.870 ;
        RECT 120.530 150.810 120.850 150.870 ;
        RECT 108.200 150.530 117.540 150.670 ;
        RECT 118.640 150.670 118.930 150.715 ;
        RECT 120.070 150.670 120.390 150.730 ;
        RECT 121.900 150.670 122.190 150.715 ;
        RECT 118.640 150.530 122.190 150.670 ;
        RECT 98.450 150.470 98.770 150.530 ;
        RECT 99.845 150.485 100.135 150.530 ;
        RECT 118.640 150.485 118.930 150.530 ;
        RECT 120.070 150.470 120.390 150.530 ;
        RECT 121.900 150.485 122.190 150.530 ;
        RECT 122.820 150.670 123.110 150.715 ;
        RECT 124.680 150.670 124.970 150.715 ;
        RECT 122.820 150.530 124.970 150.670 ;
        RECT 122.820 150.485 123.110 150.530 ;
        RECT 124.680 150.485 124.970 150.530 ;
        RECT 95.345 150.330 95.635 150.375 ;
        RECT 98.925 150.330 99.215 150.375 ;
        RECT 100.760 150.330 101.050 150.375 ;
        RECT 95.345 150.190 101.050 150.330 ;
        RECT 95.345 150.145 95.635 150.190 ;
        RECT 98.925 150.145 99.215 150.190 ;
        RECT 100.760 150.145 101.050 150.190 ;
        RECT 104.430 150.130 104.750 150.390 ;
        RECT 104.890 150.130 105.210 150.390 ;
        RECT 105.825 150.145 106.115 150.375 ;
        RECT 106.285 150.330 106.575 150.375 ;
        RECT 106.730 150.330 107.050 150.390 ;
        RECT 106.285 150.190 107.050 150.330 ;
        RECT 106.285 150.145 106.575 150.190 ;
        RECT 99.830 149.990 100.150 150.050 ;
        RECT 101.225 149.990 101.515 150.035 ;
        RECT 81.060 149.850 81.660 149.990 ;
        RECT 81.520 149.710 81.660 149.850 ;
        RECT 99.830 149.850 101.515 149.990 ;
        RECT 105.900 149.990 106.040 150.145 ;
        RECT 106.730 150.130 107.050 150.190 ;
        RECT 107.190 150.130 107.510 150.390 ;
        RECT 107.665 150.330 107.955 150.375 ;
        RECT 109.030 150.330 109.350 150.390 ;
        RECT 107.665 150.190 109.350 150.330 ;
        RECT 107.665 150.145 107.955 150.190 ;
        RECT 109.030 150.130 109.350 150.190 ;
        RECT 109.950 150.330 110.270 150.390 ;
        RECT 110.425 150.330 110.715 150.375 ;
        RECT 109.950 150.190 110.715 150.330 ;
        RECT 109.950 150.130 110.270 150.190 ;
        RECT 110.425 150.145 110.715 150.190 ;
        RECT 110.870 150.130 111.190 150.390 ;
        RECT 111.345 150.145 111.635 150.375 ;
        RECT 111.420 149.990 111.560 150.145 ;
        RECT 112.250 150.130 112.570 150.390 ;
        RECT 120.500 150.330 120.790 150.375 ;
        RECT 122.820 150.330 123.035 150.485 ;
        RECT 120.500 150.190 123.035 150.330 ;
        RECT 120.500 150.145 120.790 150.190 ;
        RECT 123.750 150.130 124.070 150.390 ;
        RECT 125.590 150.130 125.910 150.390 ;
        RECT 116.390 149.990 116.710 150.050 ;
        RECT 105.900 149.850 109.260 149.990 ;
        RECT 111.420 149.850 116.710 149.990 ;
        RECT 99.830 149.790 100.150 149.850 ;
        RECT 101.225 149.805 101.515 149.850 ;
        RECT 64.410 149.650 64.730 149.710 ;
        RECT 61.280 149.510 64.730 149.650 ;
        RECT 51.070 149.450 51.390 149.510 ;
        RECT 64.410 149.450 64.730 149.510 ;
        RECT 68.550 149.650 68.870 149.710 ;
        RECT 69.470 149.650 69.790 149.710 ;
        RECT 73.625 149.650 73.915 149.695 ;
        RECT 68.550 149.510 69.790 149.650 ;
        RECT 68.550 149.450 68.870 149.510 ;
        RECT 69.470 149.450 69.790 149.510 ;
        RECT 71.170 149.510 81.200 149.650 ;
        RECT 42.880 149.170 45.320 149.310 ;
        RECT 48.785 149.310 49.075 149.355 ;
        RECT 49.230 149.310 49.550 149.370 ;
        RECT 48.785 149.170 49.550 149.310 ;
        RECT 41.870 149.110 42.190 149.170 ;
        RECT 42.345 149.125 42.635 149.170 ;
        RECT 48.785 149.125 49.075 149.170 ;
        RECT 49.230 149.110 49.550 149.170 ;
        RECT 59.350 149.110 59.670 149.370 ;
        RECT 60.270 149.310 60.590 149.370 ;
        RECT 61.650 149.310 61.970 149.370 ;
        RECT 60.270 149.170 61.970 149.310 ;
        RECT 60.270 149.110 60.590 149.170 ;
        RECT 61.650 149.110 61.970 149.170 ;
        RECT 64.870 149.110 65.190 149.370 ;
        RECT 66.710 149.310 67.030 149.370 ;
        RECT 71.170 149.310 71.310 149.510 ;
        RECT 73.625 149.465 73.915 149.510 ;
        RECT 66.710 149.170 71.310 149.310 ;
        RECT 71.770 149.310 72.090 149.370 ;
        RECT 75.465 149.310 75.755 149.355 ;
        RECT 71.770 149.170 75.755 149.310 ;
        RECT 66.710 149.110 67.030 149.170 ;
        RECT 71.770 149.110 72.090 149.170 ;
        RECT 75.465 149.125 75.755 149.170 ;
        RECT 79.590 149.110 79.910 149.370 ;
        RECT 81.060 149.310 81.200 149.510 ;
        RECT 81.430 149.450 81.750 149.710 ;
        RECT 95.345 149.650 95.635 149.695 ;
        RECT 98.465 149.650 98.755 149.695 ;
        RECT 100.355 149.650 100.645 149.695 ;
        RECT 105.810 149.650 106.130 149.710 ;
        RECT 109.120 149.695 109.260 149.850 ;
        RECT 116.390 149.790 116.710 149.850 ;
        RECT 89.800 149.510 95.000 149.650 ;
        RECT 89.800 149.310 89.940 149.510 ;
        RECT 81.060 149.170 89.940 149.310 ;
        RECT 90.185 149.310 90.475 149.355 ;
        RECT 90.630 149.310 90.950 149.370 ;
        RECT 90.185 149.170 90.950 149.310 ;
        RECT 90.185 149.125 90.475 149.170 ;
        RECT 90.630 149.110 90.950 149.170 ;
        RECT 92.025 149.310 92.315 149.355 ;
        RECT 93.850 149.310 94.170 149.370 ;
        RECT 92.025 149.170 94.170 149.310 ;
        RECT 94.860 149.310 95.000 149.510 ;
        RECT 95.345 149.510 100.645 149.650 ;
        RECT 95.345 149.465 95.635 149.510 ;
        RECT 98.465 149.465 98.755 149.510 ;
        RECT 100.355 149.465 100.645 149.510 ;
        RECT 102.220 149.510 106.130 149.650 ;
        RECT 100.750 149.310 101.070 149.370 ;
        RECT 102.220 149.310 102.360 149.510 ;
        RECT 105.810 149.450 106.130 149.510 ;
        RECT 109.045 149.465 109.335 149.695 ;
        RECT 110.870 149.650 111.190 149.710 ;
        RECT 119.610 149.650 119.930 149.710 ;
        RECT 110.870 149.510 119.930 149.650 ;
        RECT 110.870 149.450 111.190 149.510 ;
        RECT 119.610 149.450 119.930 149.510 ;
        RECT 120.500 149.650 120.790 149.695 ;
        RECT 123.280 149.650 123.570 149.695 ;
        RECT 125.140 149.650 125.430 149.695 ;
        RECT 120.500 149.510 125.430 149.650 ;
        RECT 120.500 149.465 120.790 149.510 ;
        RECT 123.280 149.465 123.570 149.510 ;
        RECT 125.140 149.465 125.430 149.510 ;
        RECT 94.860 149.170 102.360 149.310 ;
        RECT 102.590 149.310 102.910 149.370 ;
        RECT 104.445 149.310 104.735 149.355 ;
        RECT 102.590 149.170 104.735 149.310 ;
        RECT 92.025 149.125 92.315 149.170 ;
        RECT 93.850 149.110 94.170 149.170 ;
        RECT 100.750 149.110 101.070 149.170 ;
        RECT 102.590 149.110 102.910 149.170 ;
        RECT 104.445 149.125 104.735 149.170 ;
        RECT 106.270 149.110 106.590 149.370 ;
        RECT 108.585 149.310 108.875 149.355 ;
        RECT 112.710 149.310 113.030 149.370 ;
        RECT 108.585 149.170 113.030 149.310 ;
        RECT 108.585 149.125 108.875 149.170 ;
        RECT 112.710 149.110 113.030 149.170 ;
        RECT 116.635 149.310 116.925 149.355 ;
        RECT 118.230 149.310 118.550 149.370 ;
        RECT 116.635 149.170 118.550 149.310 ;
        RECT 116.635 149.125 116.925 149.170 ;
        RECT 118.230 149.110 118.550 149.170 ;
        RECT 14.660 148.490 127.820 148.970 ;
        RECT 23.945 148.290 24.235 148.335 ;
        RECT 24.390 148.290 24.710 148.350 ;
        RECT 23.945 148.150 24.710 148.290 ;
        RECT 23.945 148.105 24.235 148.150 ;
        RECT 24.390 148.090 24.710 148.150 ;
        RECT 35.430 148.090 35.750 148.350 ;
        RECT 39.110 148.090 39.430 148.350 ;
        RECT 65.330 148.290 65.650 148.350 ;
        RECT 63.120 148.150 70.160 148.290 ;
        RECT 63.120 147.950 63.260 148.150 ;
        RECT 65.330 148.090 65.650 148.150 ;
        RECT 39.200 147.810 63.260 147.950 ;
        RECT 63.460 147.950 63.750 147.995 ;
        RECT 66.240 147.950 66.530 147.995 ;
        RECT 68.100 147.950 68.390 147.995 ;
        RECT 63.460 147.810 68.390 147.950 ;
        RECT 35.445 147.610 35.735 147.655 ;
        RECT 37.270 147.610 37.590 147.670 ;
        RECT 35.445 147.470 37.590 147.610 ;
        RECT 35.445 147.425 35.735 147.470 ;
        RECT 37.270 147.410 37.590 147.470 ;
        RECT 23.025 147.270 23.315 147.315 ;
        RECT 23.930 147.270 24.250 147.330 ;
        RECT 23.025 147.130 24.250 147.270 ;
        RECT 23.025 147.085 23.315 147.130 ;
        RECT 23.930 147.070 24.250 147.130 ;
        RECT 34.525 147.270 34.815 147.315 ;
        RECT 34.970 147.270 35.290 147.330 ;
        RECT 39.200 147.315 39.340 147.810 ;
        RECT 63.460 147.765 63.750 147.810 ;
        RECT 66.240 147.765 66.530 147.810 ;
        RECT 68.100 147.765 68.390 147.810 ;
        RECT 69.025 147.765 69.315 147.995 ;
        RECT 40.030 147.410 40.350 147.670 ;
        RECT 58.430 147.610 58.750 147.670 ;
        RECT 59.595 147.610 59.885 147.655 ;
        RECT 60.270 147.610 60.590 147.670 ;
        RECT 58.430 147.470 60.590 147.610 ;
        RECT 58.430 147.410 58.750 147.470 ;
        RECT 59.595 147.425 59.885 147.470 ;
        RECT 60.270 147.410 60.590 147.470 ;
        RECT 60.730 147.610 61.050 147.670 ;
        RECT 66.725 147.610 67.015 147.655 ;
        RECT 69.100 147.610 69.240 147.765 ;
        RECT 60.730 147.470 66.480 147.610 ;
        RECT 60.730 147.410 61.050 147.470 ;
        RECT 34.525 147.130 35.290 147.270 ;
        RECT 34.525 147.085 34.815 147.130 ;
        RECT 34.970 147.070 35.290 147.130 ;
        RECT 39.125 147.085 39.415 147.315 ;
        RECT 40.505 147.270 40.795 147.315 ;
        RECT 44.170 147.270 44.490 147.330 ;
        RECT 40.505 147.130 44.490 147.270 ;
        RECT 40.505 147.085 40.795 147.130 ;
        RECT 44.170 147.070 44.490 147.130 ;
        RECT 53.370 147.070 53.690 147.330 ;
        RECT 63.460 147.270 63.750 147.315 ;
        RECT 66.340 147.270 66.480 147.470 ;
        RECT 66.725 147.470 69.240 147.610 ;
        RECT 66.725 147.425 67.015 147.470 ;
        RECT 70.020 147.315 70.160 148.150 ;
        RECT 104.430 148.090 104.750 148.350 ;
        RECT 106.730 148.290 107.050 148.350 ;
        RECT 109.045 148.290 109.335 148.335 ;
        RECT 106.730 148.150 109.335 148.290 ;
        RECT 106.730 148.090 107.050 148.150 ;
        RECT 109.045 148.105 109.335 148.150 ;
        RECT 120.085 148.290 120.375 148.335 ;
        RECT 121.450 148.290 121.770 148.350 ;
        RECT 120.085 148.150 121.770 148.290 ;
        RECT 120.085 148.105 120.375 148.150 ;
        RECT 121.450 148.090 121.770 148.150 ;
        RECT 90.140 147.950 90.430 147.995 ;
        RECT 92.920 147.950 93.210 147.995 ;
        RECT 94.780 147.950 95.070 147.995 ;
        RECT 90.140 147.810 95.070 147.950 ;
        RECT 90.140 147.765 90.430 147.810 ;
        RECT 92.920 147.765 93.210 147.810 ;
        RECT 94.780 147.765 95.070 147.810 ;
        RECT 102.605 147.950 102.895 147.995 ;
        RECT 110.870 147.950 111.190 148.010 ;
        RECT 102.605 147.810 111.190 147.950 ;
        RECT 102.605 147.765 102.895 147.810 ;
        RECT 110.870 147.750 111.190 147.810 ;
        RECT 70.850 147.610 71.170 147.670 ;
        RECT 73.610 147.610 73.930 147.670 ;
        RECT 70.480 147.470 73.930 147.610 ;
        RECT 70.480 147.315 70.620 147.470 ;
        RECT 70.850 147.410 71.170 147.470 ;
        RECT 73.610 147.410 73.930 147.470 ;
        RECT 93.405 147.610 93.695 147.655 ;
        RECT 93.850 147.610 94.170 147.670 ;
        RECT 93.405 147.470 94.170 147.610 ;
        RECT 93.405 147.425 93.695 147.470 ;
        RECT 93.850 147.410 94.170 147.470 ;
        RECT 103.970 147.410 104.290 147.670 ;
        RECT 105.810 147.410 106.130 147.670 ;
        RECT 116.850 147.610 117.170 147.670 ;
        RECT 107.740 147.470 117.170 147.610 ;
        RECT 68.565 147.270 68.855 147.315 ;
        RECT 63.460 147.130 65.995 147.270 ;
        RECT 66.340 147.130 68.855 147.270 ;
        RECT 63.460 147.085 63.750 147.130 ;
        RECT 35.905 146.930 36.195 146.975 ;
        RECT 59.350 146.930 59.670 146.990 ;
        RECT 35.905 146.790 59.670 146.930 ;
        RECT 35.905 146.745 36.195 146.790 ;
        RECT 59.350 146.730 59.670 146.790 ;
        RECT 61.600 146.930 61.890 146.975 ;
        RECT 63.950 146.930 64.270 146.990 ;
        RECT 65.780 146.975 65.995 147.130 ;
        RECT 68.565 147.085 68.855 147.130 ;
        RECT 69.945 147.085 70.235 147.315 ;
        RECT 70.405 147.085 70.695 147.315 ;
        RECT 71.785 147.270 72.075 147.315 ;
        RECT 71.400 147.130 72.075 147.270 ;
        RECT 64.860 146.930 65.150 146.975 ;
        RECT 61.600 146.790 65.150 146.930 ;
        RECT 61.600 146.745 61.890 146.790 ;
        RECT 63.950 146.730 64.270 146.790 ;
        RECT 64.860 146.745 65.150 146.790 ;
        RECT 65.780 146.930 66.070 146.975 ;
        RECT 67.640 146.930 67.930 146.975 ;
        RECT 65.780 146.790 67.930 146.930 ;
        RECT 65.780 146.745 66.070 146.790 ;
        RECT 67.640 146.745 67.930 146.790 ;
        RECT 69.010 146.930 69.330 146.990 ;
        RECT 70.865 146.930 71.155 146.975 ;
        RECT 69.010 146.790 71.155 146.930 ;
        RECT 69.010 146.730 69.330 146.790 ;
        RECT 70.865 146.745 71.155 146.790 ;
        RECT 27.610 146.590 27.930 146.650 ;
        RECT 33.605 146.590 33.895 146.635 ;
        RECT 27.610 146.450 33.895 146.590 ;
        RECT 27.610 146.390 27.930 146.450 ;
        RECT 33.605 146.405 33.895 146.450 ;
        RECT 34.970 146.590 35.290 146.650 ;
        RECT 38.205 146.590 38.495 146.635 ;
        RECT 34.970 146.450 38.495 146.590 ;
        RECT 34.970 146.390 35.290 146.450 ;
        RECT 38.205 146.405 38.495 146.450 ;
        RECT 53.370 146.590 53.690 146.650 ;
        RECT 53.845 146.590 54.135 146.635 ;
        RECT 53.370 146.450 54.135 146.590 ;
        RECT 53.370 146.390 53.690 146.450 ;
        RECT 53.845 146.405 54.135 146.450 ;
        RECT 60.270 146.590 60.590 146.650 ;
        RECT 71.400 146.590 71.540 147.130 ;
        RECT 71.785 147.085 72.075 147.130 ;
        RECT 90.140 147.270 90.430 147.315 ;
        RECT 90.140 147.130 92.675 147.270 ;
        RECT 90.140 147.085 90.430 147.130 ;
        RECT 88.280 146.930 88.570 146.975 ;
        RECT 90.630 146.930 90.950 146.990 ;
        RECT 92.460 146.975 92.675 147.130 ;
        RECT 95.230 147.070 95.550 147.330 ;
        RECT 103.510 147.070 103.830 147.330 ;
        RECT 105.900 147.270 106.040 147.410 ;
        RECT 106.730 147.270 107.050 147.330 ;
        RECT 107.740 147.315 107.880 147.470 ;
        RECT 116.850 147.410 117.170 147.470 ;
        RECT 117.310 147.410 117.630 147.670 ;
        RECT 105.900 147.130 107.050 147.270 ;
        RECT 106.730 147.070 107.050 147.130 ;
        RECT 107.205 147.085 107.495 147.315 ;
        RECT 107.665 147.085 107.955 147.315 ;
        RECT 108.585 147.270 108.875 147.315 ;
        RECT 109.030 147.270 109.350 147.330 ;
        RECT 108.585 147.130 109.350 147.270 ;
        RECT 108.585 147.085 108.875 147.130 ;
        RECT 91.540 146.930 91.830 146.975 ;
        RECT 88.280 146.790 91.830 146.930 ;
        RECT 88.280 146.745 88.570 146.790 ;
        RECT 90.630 146.730 90.950 146.790 ;
        RECT 91.540 146.745 91.830 146.790 ;
        RECT 92.460 146.930 92.750 146.975 ;
        RECT 94.320 146.930 94.610 146.975 ;
        RECT 92.460 146.790 94.610 146.930 ;
        RECT 92.460 146.745 92.750 146.790 ;
        RECT 94.320 146.745 94.610 146.790 ;
        RECT 104.905 146.930 105.195 146.975 ;
        RECT 105.365 146.930 105.655 146.975 ;
        RECT 104.905 146.790 105.655 146.930 ;
        RECT 104.905 146.745 105.195 146.790 ;
        RECT 105.365 146.745 105.655 146.790 ;
        RECT 105.810 146.930 106.130 146.990 ;
        RECT 107.280 146.930 107.420 147.085 ;
        RECT 105.810 146.790 107.420 146.930 ;
        RECT 105.810 146.730 106.130 146.790 ;
        RECT 60.270 146.450 71.540 146.590 ;
        RECT 86.030 146.635 86.350 146.650 ;
        RECT 60.270 146.390 60.590 146.450 ;
        RECT 86.030 146.405 86.565 146.635 ;
        RECT 95.690 146.590 96.010 146.650 ;
        RECT 107.740 146.590 107.880 147.085 ;
        RECT 109.030 147.070 109.350 147.130 ;
        RECT 110.425 147.085 110.715 147.315 ;
        RECT 108.110 146.930 108.430 146.990 ;
        RECT 109.950 146.930 110.270 146.990 ;
        RECT 110.500 146.930 110.640 147.085 ;
        RECT 110.870 147.070 111.190 147.330 ;
        RECT 111.345 147.085 111.635 147.315 ;
        RECT 108.110 146.790 110.640 146.930 ;
        RECT 111.420 146.930 111.560 147.085 ;
        RECT 112.250 147.070 112.570 147.330 ;
        RECT 116.390 147.270 116.710 147.330 ;
        RECT 118.245 147.270 118.535 147.315 ;
        RECT 116.390 147.130 118.535 147.270 ;
        RECT 116.390 147.070 116.710 147.130 ;
        RECT 118.245 147.085 118.535 147.130 ;
        RECT 111.420 146.790 118.000 146.930 ;
        RECT 108.110 146.730 108.430 146.790 ;
        RECT 109.950 146.730 110.270 146.790 ;
        RECT 117.860 146.635 118.000 146.790 ;
        RECT 95.690 146.450 107.880 146.590 ;
        RECT 117.785 146.590 118.075 146.635 ;
        RECT 118.230 146.590 118.550 146.650 ;
        RECT 117.785 146.450 118.550 146.590 ;
        RECT 86.030 146.390 86.350 146.405 ;
        RECT 95.690 146.390 96.010 146.450 ;
        RECT 117.785 146.405 118.075 146.450 ;
        RECT 118.230 146.390 118.550 146.450 ;
        RECT 14.660 145.770 127.820 146.250 ;
        RECT 54.750 145.570 55.070 145.630 ;
        RECT 68.550 145.570 68.870 145.630 ;
        RECT 71.770 145.570 72.090 145.630 ;
        RECT 81.430 145.570 81.750 145.630 ;
        RECT 82.810 145.570 83.130 145.630 ;
        RECT 86.505 145.570 86.795 145.615 ;
        RECT 49.320 145.430 67.860 145.570 ;
        RECT 18.360 145.230 18.650 145.275 ;
        RECT 18.870 145.230 19.190 145.290 ;
        RECT 21.620 145.230 21.910 145.275 ;
        RECT 18.360 145.090 21.910 145.230 ;
        RECT 18.360 145.045 18.650 145.090 ;
        RECT 18.870 145.030 19.190 145.090 ;
        RECT 21.620 145.045 21.910 145.090 ;
        RECT 22.540 145.230 22.830 145.275 ;
        RECT 24.400 145.230 24.690 145.275 ;
        RECT 22.540 145.090 24.690 145.230 ;
        RECT 22.540 145.045 22.830 145.090 ;
        RECT 24.400 145.045 24.690 145.090 ;
        RECT 44.645 145.230 44.935 145.275 ;
        RECT 47.405 145.230 47.695 145.275 ;
        RECT 44.645 145.090 47.695 145.230 ;
        RECT 44.645 145.045 44.935 145.090 ;
        RECT 47.405 145.045 47.695 145.090 ;
        RECT 20.220 144.890 20.510 144.935 ;
        RECT 22.540 144.890 22.755 145.045 ;
        RECT 20.220 144.750 22.755 144.890 ;
        RECT 20.220 144.705 20.510 144.750 ;
        RECT 34.050 144.690 34.370 144.950 ;
        RECT 35.445 144.890 35.735 144.935 ;
        RECT 36.810 144.890 37.130 144.950 ;
        RECT 35.445 144.750 37.130 144.890 ;
        RECT 35.445 144.705 35.735 144.750 ;
        RECT 36.810 144.690 37.130 144.750 ;
        RECT 46.010 144.690 46.330 144.950 ;
        RECT 49.320 144.935 49.460 145.430 ;
        RECT 54.750 145.370 55.070 145.430 ;
        RECT 52.565 145.230 52.855 145.275 ;
        RECT 53.370 145.230 53.690 145.290 ;
        RECT 55.805 145.230 56.455 145.275 ;
        RECT 52.565 145.090 56.455 145.230 ;
        RECT 52.565 145.045 53.155 145.090 ;
        RECT 48.785 144.705 49.075 144.935 ;
        RECT 49.245 144.705 49.535 144.935 ;
        RECT 49.705 144.705 49.995 144.935 ;
        RECT 50.625 144.890 50.915 144.935 ;
        RECT 50.625 144.750 52.680 144.890 ;
        RECT 50.625 144.705 50.915 144.750 ;
        RECT 21.170 144.550 21.490 144.610 ;
        RECT 23.485 144.550 23.775 144.595 ;
        RECT 21.170 144.410 23.775 144.550 ;
        RECT 21.170 144.350 21.490 144.410 ;
        RECT 23.485 144.365 23.775 144.410 ;
        RECT 25.310 144.350 25.630 144.610 ;
        RECT 30.830 144.550 31.150 144.610 ;
        RECT 34.525 144.550 34.815 144.595 ;
        RECT 30.830 144.410 34.815 144.550 ;
        RECT 30.830 144.350 31.150 144.410 ;
        RECT 34.525 144.365 34.815 144.410 ;
        RECT 45.090 144.350 45.410 144.610 ;
        RECT 48.860 144.550 49.000 144.705 ;
        RECT 49.780 144.550 49.920 144.705 ;
        RECT 52.540 144.550 52.680 144.750 ;
        RECT 52.865 144.730 53.155 145.045 ;
        RECT 53.370 145.030 53.690 145.090 ;
        RECT 55.805 145.045 56.455 145.090 ;
        RECT 53.945 144.890 54.235 144.935 ;
        RECT 57.525 144.890 57.815 144.935 ;
        RECT 59.360 144.890 59.650 144.935 ;
        RECT 53.945 144.750 59.650 144.890 ;
        RECT 53.945 144.705 54.235 144.750 ;
        RECT 57.525 144.705 57.815 144.750 ;
        RECT 59.360 144.705 59.650 144.750 ;
        RECT 61.190 144.690 61.510 144.950 ;
        RECT 65.345 144.705 65.635 144.935 ;
        RECT 55.210 144.550 55.530 144.610 ;
        RECT 48.860 144.410 49.460 144.550 ;
        RECT 49.780 144.410 51.300 144.550 ;
        RECT 52.540 144.410 55.530 144.550 ;
        RECT 20.220 144.210 20.510 144.255 ;
        RECT 23.000 144.210 23.290 144.255 ;
        RECT 24.860 144.210 25.150 144.255 ;
        RECT 20.220 144.070 25.150 144.210 ;
        RECT 49.320 144.210 49.460 144.410 ;
        RECT 50.610 144.210 50.930 144.270 ;
        RECT 49.320 144.070 50.930 144.210 ;
        RECT 20.220 144.025 20.510 144.070 ;
        RECT 23.000 144.025 23.290 144.070 ;
        RECT 24.860 144.025 25.150 144.070 ;
        RECT 50.610 144.010 50.930 144.070 ;
        RECT 16.355 143.870 16.645 143.915 ;
        RECT 21.630 143.870 21.950 143.930 ;
        RECT 16.355 143.730 21.950 143.870 ;
        RECT 16.355 143.685 16.645 143.730 ;
        RECT 21.630 143.670 21.950 143.730 ;
        RECT 30.370 143.870 30.690 143.930 ;
        RECT 33.145 143.870 33.435 143.915 ;
        RECT 30.370 143.730 33.435 143.870 ;
        RECT 30.370 143.670 30.690 143.730 ;
        RECT 33.145 143.685 33.435 143.730 ;
        RECT 34.050 143.670 34.370 143.930 ;
        RECT 46.010 143.670 46.330 143.930 ;
        RECT 46.930 143.670 47.250 143.930 ;
        RECT 51.160 143.915 51.300 144.410 ;
        RECT 55.210 144.350 55.530 144.410 ;
        RECT 58.445 144.550 58.735 144.595 ;
        RECT 58.445 144.410 59.580 144.550 ;
        RECT 58.445 144.365 58.735 144.410 ;
        RECT 53.945 144.210 54.235 144.255 ;
        RECT 57.065 144.210 57.355 144.255 ;
        RECT 58.955 144.210 59.245 144.255 ;
        RECT 53.945 144.070 59.245 144.210 ;
        RECT 59.440 144.210 59.580 144.410 ;
        RECT 59.810 144.350 60.130 144.610 ;
        RECT 65.420 144.550 65.560 144.705 ;
        RECT 65.790 144.690 66.110 144.950 ;
        RECT 66.250 144.690 66.570 144.950 ;
        RECT 67.185 144.705 67.475 144.935 ;
        RECT 66.710 144.550 67.030 144.610 ;
        RECT 65.420 144.410 67.030 144.550 ;
        RECT 66.710 144.350 67.030 144.410 ;
        RECT 60.285 144.210 60.575 144.255 ;
        RECT 59.440 144.070 60.575 144.210 ;
        RECT 53.945 144.025 54.235 144.070 ;
        RECT 57.065 144.025 57.355 144.070 ;
        RECT 58.955 144.025 59.245 144.070 ;
        RECT 60.285 144.025 60.575 144.070 ;
        RECT 65.330 144.210 65.650 144.270 ;
        RECT 67.260 144.210 67.400 144.705 ;
        RECT 65.330 144.070 67.400 144.210 ;
        RECT 67.720 144.210 67.860 145.430 ;
        RECT 68.550 145.430 71.080 145.570 ;
        RECT 68.550 145.370 68.870 145.430 ;
        RECT 70.390 145.030 70.710 145.290 ;
        RECT 70.940 145.230 71.080 145.430 ;
        RECT 71.770 145.430 82.580 145.570 ;
        RECT 71.770 145.370 72.090 145.430 ;
        RECT 81.430 145.370 81.750 145.430 ;
        RECT 80.525 145.230 80.815 145.275 ;
        RECT 80.985 145.230 81.275 145.275 ;
        RECT 70.940 145.090 80.280 145.230 ;
        RECT 73.625 144.890 73.915 144.935 ;
        RECT 72.320 144.750 73.915 144.890 ;
        RECT 69.010 144.350 69.330 144.610 ;
        RECT 69.930 144.350 70.250 144.610 ;
        RECT 71.770 144.210 72.090 144.270 ;
        RECT 72.320 144.255 72.460 144.750 ;
        RECT 73.625 144.705 73.915 144.750 ;
        RECT 79.130 144.690 79.450 144.950 ;
        RECT 80.140 144.890 80.280 145.090 ;
        RECT 80.525 145.090 81.275 145.230 ;
        RECT 82.440 145.230 82.580 145.430 ;
        RECT 82.810 145.430 86.795 145.570 ;
        RECT 82.810 145.370 83.130 145.430 ;
        RECT 86.505 145.385 86.795 145.430 ;
        RECT 88.345 145.570 88.635 145.615 ;
        RECT 91.090 145.570 91.410 145.630 ;
        RECT 88.345 145.430 91.410 145.570 ;
        RECT 88.345 145.385 88.635 145.430 ;
        RECT 91.090 145.370 91.410 145.430 ;
        RECT 94.325 145.570 94.615 145.615 ;
        RECT 95.690 145.570 96.010 145.630 ;
        RECT 94.325 145.430 96.010 145.570 ;
        RECT 94.325 145.385 94.615 145.430 ;
        RECT 95.690 145.370 96.010 145.430 ;
        RECT 96.610 145.370 96.930 145.630 ;
        RECT 86.030 145.230 86.350 145.290 ;
        RECT 94.785 145.230 95.075 145.275 ;
        RECT 82.440 145.090 83.040 145.230 ;
        RECT 80.525 145.045 80.815 145.090 ;
        RECT 80.985 145.045 81.275 145.090 ;
        RECT 81.890 144.890 82.210 144.950 ;
        RECT 82.900 144.935 83.040 145.090 ;
        RECT 83.360 145.090 95.075 145.230 ;
        RECT 83.360 144.935 83.500 145.090 ;
        RECT 86.030 145.030 86.350 145.090 ;
        RECT 94.785 145.045 95.075 145.090 ;
        RECT 109.030 145.230 109.350 145.290 ;
        RECT 112.250 145.230 112.570 145.290 ;
        RECT 109.030 145.090 112.570 145.230 ;
        RECT 109.030 145.030 109.350 145.090 ;
        RECT 82.365 144.890 82.655 144.935 ;
        RECT 80.140 144.750 82.655 144.890 ;
        RECT 81.890 144.690 82.210 144.750 ;
        RECT 82.365 144.705 82.655 144.750 ;
        RECT 82.825 144.705 83.115 144.935 ;
        RECT 83.285 144.705 83.575 144.935 ;
        RECT 83.730 144.890 84.050 144.950 ;
        RECT 84.205 144.890 84.495 144.935 ;
        RECT 83.730 144.750 84.495 144.890 ;
        RECT 83.730 144.690 84.050 144.750 ;
        RECT 84.205 144.705 84.495 144.750 ;
        RECT 109.950 144.690 110.270 144.950 ;
        RECT 110.410 144.690 110.730 144.950 ;
        RECT 111.880 144.935 112.020 145.090 ;
        RECT 112.250 145.030 112.570 145.090 ;
        RECT 110.885 144.705 111.175 144.935 ;
        RECT 111.805 144.705 112.095 144.935 ;
        RECT 80.065 144.550 80.355 144.595 ;
        RECT 80.510 144.550 80.830 144.610 ;
        RECT 80.065 144.410 80.830 144.550 ;
        RECT 80.065 144.365 80.355 144.410 ;
        RECT 80.510 144.350 80.830 144.410 ;
        RECT 85.110 144.550 85.430 144.610 ;
        RECT 93.405 144.550 93.695 144.595 ;
        RECT 110.500 144.550 110.640 144.690 ;
        RECT 85.110 144.410 93.695 144.550 ;
        RECT 85.110 144.350 85.430 144.410 ;
        RECT 93.405 144.365 93.695 144.410 ;
        RECT 108.200 144.410 110.640 144.550 ;
        RECT 110.960 144.550 111.100 144.705 ;
        RECT 114.090 144.550 114.410 144.610 ;
        RECT 110.960 144.410 114.410 144.550 ;
        RECT 108.200 144.270 108.340 144.410 ;
        RECT 114.090 144.350 114.410 144.410 ;
        RECT 67.720 144.070 72.090 144.210 ;
        RECT 65.330 144.010 65.650 144.070 ;
        RECT 71.770 144.010 72.090 144.070 ;
        RECT 72.245 144.025 72.535 144.255 ;
        RECT 100.290 144.210 100.610 144.270 ;
        RECT 105.810 144.210 106.130 144.270 ;
        RECT 108.110 144.210 108.430 144.270 ;
        RECT 74.160 144.070 108.430 144.210 ;
        RECT 51.085 143.870 51.375 143.915 ;
        RECT 57.970 143.870 58.290 143.930 ;
        RECT 51.085 143.730 58.290 143.870 ;
        RECT 51.085 143.685 51.375 143.730 ;
        RECT 57.970 143.670 58.290 143.730 ;
        RECT 60.730 143.870 61.050 143.930 ;
        RECT 63.965 143.870 64.255 143.915 ;
        RECT 60.730 143.730 64.255 143.870 ;
        RECT 60.730 143.670 61.050 143.730 ;
        RECT 63.965 143.685 64.255 143.730 ;
        RECT 64.410 143.870 64.730 143.930 ;
        RECT 65.790 143.870 66.110 143.930 ;
        RECT 74.160 143.870 74.300 144.070 ;
        RECT 100.290 144.010 100.610 144.070 ;
        RECT 105.810 144.010 106.130 144.070 ;
        RECT 108.110 144.010 108.430 144.070 ;
        RECT 64.410 143.730 74.300 143.870 ;
        RECT 64.410 143.670 64.730 143.730 ;
        RECT 65.790 143.670 66.110 143.730 ;
        RECT 74.530 143.670 74.850 143.930 ;
        RECT 78.210 143.670 78.530 143.930 ;
        RECT 80.525 143.870 80.815 143.915 ;
        RECT 84.190 143.870 84.510 143.930 ;
        RECT 80.525 143.730 84.510 143.870 ;
        RECT 80.525 143.685 80.815 143.730 ;
        RECT 84.190 143.670 84.510 143.730 ;
        RECT 102.130 143.870 102.450 143.930 ;
        RECT 103.970 143.870 104.290 143.930 ;
        RECT 102.130 143.730 104.290 143.870 ;
        RECT 102.130 143.670 102.450 143.730 ;
        RECT 103.970 143.670 104.290 143.730 ;
        RECT 107.190 143.870 107.510 143.930 ;
        RECT 108.585 143.870 108.875 143.915 ;
        RECT 107.190 143.730 108.875 143.870 ;
        RECT 107.190 143.670 107.510 143.730 ;
        RECT 108.585 143.685 108.875 143.730 ;
        RECT 14.660 143.050 127.820 143.530 ;
        RECT 35.445 142.665 35.735 142.895 ;
        RECT 46.930 142.850 47.250 142.910 ;
        RECT 58.890 142.850 59.210 142.910 ;
        RECT 46.930 142.710 59.210 142.850 ;
        RECT 34.065 142.510 34.355 142.555 ;
        RECT 35.520 142.510 35.660 142.665 ;
        RECT 46.930 142.650 47.250 142.710 ;
        RECT 58.890 142.650 59.210 142.710 ;
        RECT 60.285 142.850 60.575 142.895 ;
        RECT 61.190 142.850 61.510 142.910 ;
        RECT 60.285 142.710 61.510 142.850 ;
        RECT 60.285 142.665 60.575 142.710 ;
        RECT 61.190 142.650 61.510 142.710 ;
        RECT 66.495 142.850 66.785 142.895 ;
        RECT 69.930 142.850 70.250 142.910 ;
        RECT 66.495 142.710 70.250 142.850 ;
        RECT 66.495 142.665 66.785 142.710 ;
        RECT 69.930 142.650 70.250 142.710 ;
        RECT 79.130 142.650 79.450 142.910 ;
        RECT 80.510 142.850 80.830 142.910 ;
        RECT 83.730 142.850 84.050 142.910 ;
        RECT 80.510 142.710 84.050 142.850 ;
        RECT 80.510 142.650 80.830 142.710 ;
        RECT 83.730 142.650 84.050 142.710 ;
        RECT 104.890 142.650 105.210 142.910 ;
        RECT 117.310 142.850 117.630 142.910 ;
        RECT 112.800 142.710 117.630 142.850 ;
        RECT 34.065 142.370 35.660 142.510 ;
        RECT 36.810 142.510 37.130 142.570 ;
        RECT 62.585 142.510 62.875 142.555 ;
        RECT 36.810 142.370 62.875 142.510 ;
        RECT 34.065 142.325 34.355 142.370 ;
        RECT 36.810 142.310 37.130 142.370 ;
        RECT 62.585 142.325 62.875 142.370 ;
        RECT 67.630 142.510 67.950 142.570 ;
        RECT 68.550 142.510 68.870 142.570 ;
        RECT 67.630 142.370 68.870 142.510 ;
        RECT 67.630 142.310 67.950 142.370 ;
        RECT 68.550 142.310 68.870 142.370 ;
        RECT 70.360 142.510 70.650 142.555 ;
        RECT 73.140 142.510 73.430 142.555 ;
        RECT 75.000 142.510 75.290 142.555 ;
        RECT 102.130 142.510 102.450 142.570 ;
        RECT 109.490 142.510 109.810 142.570 ;
        RECT 70.360 142.370 75.290 142.510 ;
        RECT 70.360 142.325 70.650 142.370 ;
        RECT 73.140 142.325 73.430 142.370 ;
        RECT 75.000 142.325 75.290 142.370 ;
        RECT 75.540 142.370 102.450 142.510 ;
        RECT 36.350 141.970 36.670 142.230 ;
        RECT 57.510 141.970 57.830 142.230 ;
        RECT 60.730 142.170 61.050 142.230 ;
        RECT 66.710 142.170 67.030 142.230 ;
        RECT 73.625 142.170 73.915 142.215 ;
        RECT 74.530 142.170 74.850 142.230 ;
        RECT 75.540 142.170 75.680 142.370 ;
        RECT 102.130 142.310 102.450 142.370 ;
        RECT 104.520 142.370 109.810 142.510 ;
        RECT 58.060 142.030 61.050 142.170 ;
        RECT 20.710 141.830 21.030 141.890 ;
        RECT 32.225 141.830 32.515 141.875 ;
        RECT 20.710 141.690 32.515 141.830 ;
        RECT 20.710 141.630 21.030 141.690 ;
        RECT 32.225 141.645 32.515 141.690 ;
        RECT 33.130 141.630 33.450 141.890 ;
        RECT 35.445 141.830 35.735 141.875 ;
        RECT 35.890 141.830 36.210 141.890 ;
        RECT 35.445 141.690 36.210 141.830 ;
        RECT 35.445 141.645 35.735 141.690 ;
        RECT 35.890 141.630 36.210 141.690 ;
        RECT 36.825 141.830 37.115 141.875 ;
        RECT 58.060 141.830 58.200 142.030 ;
        RECT 60.730 141.970 61.050 142.030 ;
        RECT 64.040 142.030 67.030 142.170 ;
        RECT 36.825 141.690 58.200 141.830 ;
        RECT 36.825 141.645 37.115 141.690 ;
        RECT 58.430 141.630 58.750 141.890 ;
        RECT 64.040 141.875 64.180 142.030 ;
        RECT 66.710 141.970 67.030 142.030 ;
        RECT 70.020 142.030 73.380 142.170 ;
        RECT 63.965 141.645 64.255 141.875 ;
        RECT 64.410 141.630 64.730 141.890 ;
        RECT 64.870 141.630 65.190 141.890 ;
        RECT 65.330 141.830 65.650 141.890 ;
        RECT 65.805 141.830 66.095 141.875 ;
        RECT 70.020 141.830 70.160 142.030 ;
        RECT 65.330 141.690 70.160 141.830 ;
        RECT 70.360 141.830 70.650 141.875 ;
        RECT 73.240 141.830 73.380 142.030 ;
        RECT 73.625 142.030 74.850 142.170 ;
        RECT 73.625 141.985 73.915 142.030 ;
        RECT 74.530 141.970 74.850 142.030 ;
        RECT 75.080 142.030 75.680 142.170 ;
        RECT 78.685 142.170 78.975 142.215 ;
        RECT 83.270 142.170 83.590 142.230 ;
        RECT 78.685 142.030 83.590 142.170 ;
        RECT 75.080 141.830 75.220 142.030 ;
        RECT 78.685 141.985 78.975 142.030 ;
        RECT 83.270 141.970 83.590 142.030 ;
        RECT 85.110 141.970 85.430 142.230 ;
        RECT 70.360 141.690 72.895 141.830 ;
        RECT 73.240 141.690 75.220 141.830 ;
        RECT 65.330 141.630 65.650 141.690 ;
        RECT 65.805 141.645 66.095 141.690 ;
        RECT 70.360 141.645 70.650 141.690 ;
        RECT 57.510 141.490 57.830 141.550 ;
        RECT 58.890 141.490 59.210 141.550 ;
        RECT 67.630 141.490 67.950 141.550 ;
        RECT 71.770 141.535 72.090 141.550 ;
        RECT 57.510 141.350 58.660 141.490 ;
        RECT 57.510 141.290 57.830 141.350 ;
        RECT 34.510 140.950 34.830 141.210 ;
        RECT 57.970 140.950 58.290 141.210 ;
        RECT 58.520 141.150 58.660 141.350 ;
        RECT 58.890 141.350 67.950 141.490 ;
        RECT 58.890 141.290 59.210 141.350 ;
        RECT 67.630 141.290 67.950 141.350 ;
        RECT 68.500 141.490 68.790 141.535 ;
        RECT 71.760 141.490 72.090 141.535 ;
        RECT 68.500 141.350 72.090 141.490 ;
        RECT 68.500 141.305 68.790 141.350 ;
        RECT 71.760 141.305 72.090 141.350 ;
        RECT 72.680 141.535 72.895 141.690 ;
        RECT 75.450 141.630 75.770 141.890 ;
        RECT 76.370 141.830 76.690 141.890 ;
        RECT 79.145 141.830 79.435 141.875 ;
        RECT 76.370 141.690 79.435 141.830 ;
        RECT 76.370 141.630 76.690 141.690 ;
        RECT 79.145 141.645 79.435 141.690 ;
        RECT 81.890 141.630 82.210 141.890 ;
        RECT 82.365 141.645 82.655 141.875 ;
        RECT 72.680 141.490 72.970 141.535 ;
        RECT 74.540 141.490 74.830 141.535 ;
        RECT 72.680 141.350 74.830 141.490 ;
        RECT 72.680 141.305 72.970 141.350 ;
        RECT 74.540 141.305 74.830 141.350 ;
        RECT 77.765 141.490 78.055 141.535 ;
        RECT 80.525 141.490 80.815 141.535 ;
        RECT 77.765 141.350 80.815 141.490 ;
        RECT 77.765 141.305 78.055 141.350 ;
        RECT 80.525 141.305 80.815 141.350 ;
        RECT 81.430 141.490 81.750 141.550 ;
        RECT 82.440 141.490 82.580 141.645 ;
        RECT 82.810 141.630 83.130 141.890 ;
        RECT 83.730 141.630 84.050 141.890 ;
        RECT 86.045 141.830 86.335 141.875 ;
        RECT 84.280 141.690 86.335 141.830 ;
        RECT 81.430 141.350 82.580 141.490 ;
        RECT 82.900 141.490 83.040 141.630 ;
        RECT 84.280 141.490 84.420 141.690 ;
        RECT 86.045 141.645 86.335 141.690 ;
        RECT 89.710 141.630 90.030 141.890 ;
        RECT 104.520 141.875 104.660 142.370 ;
        RECT 109.490 142.310 109.810 142.370 ;
        RECT 105.350 141.970 105.670 142.230 ;
        RECT 109.950 142.170 110.270 142.230 ;
        RECT 107.740 142.030 110.270 142.170 ;
        RECT 104.445 141.645 104.735 141.875 ;
        RECT 105.825 141.830 106.115 141.875 ;
        RECT 107.190 141.830 107.510 141.890 ;
        RECT 107.740 141.875 107.880 142.030 ;
        RECT 109.950 141.970 110.270 142.030 ;
        RECT 112.250 142.170 112.570 142.230 ;
        RECT 112.800 142.215 112.940 142.710 ;
        RECT 117.310 142.650 117.630 142.710 ;
        RECT 115.930 142.310 116.250 142.570 ;
        RECT 117.400 142.510 117.540 142.650 ;
        RECT 117.400 142.370 119.380 142.510 ;
        RECT 119.240 142.215 119.380 142.370 ;
        RECT 112.725 142.170 113.015 142.215 ;
        RECT 118.705 142.170 118.995 142.215 ;
        RECT 112.250 142.030 113.015 142.170 ;
        RECT 112.250 141.970 112.570 142.030 ;
        RECT 112.725 141.985 113.015 142.030 ;
        RECT 114.180 142.030 118.995 142.170 ;
        RECT 114.180 141.890 114.320 142.030 ;
        RECT 118.705 141.985 118.995 142.030 ;
        RECT 119.165 141.985 119.455 142.215 ;
        RECT 105.825 141.690 107.510 141.830 ;
        RECT 105.825 141.645 106.115 141.690 ;
        RECT 107.190 141.630 107.510 141.690 ;
        RECT 107.665 141.645 107.955 141.875 ;
        RECT 108.110 141.630 108.430 141.890 ;
        RECT 108.585 141.645 108.875 141.875 ;
        RECT 109.030 141.830 109.350 141.890 ;
        RECT 109.505 141.830 109.795 141.875 ;
        RECT 109.030 141.690 109.795 141.830 ;
        RECT 82.900 141.350 84.420 141.490 ;
        RECT 84.650 141.490 84.970 141.550 ;
        RECT 89.265 141.490 89.555 141.535 ;
        RECT 108.660 141.490 108.800 141.645 ;
        RECT 109.030 141.630 109.350 141.690 ;
        RECT 109.505 141.645 109.795 141.690 ;
        RECT 114.090 141.630 114.410 141.890 ;
        RECT 118.230 141.630 118.550 141.890 ;
        RECT 120.070 141.830 120.390 141.890 ;
        RECT 120.545 141.830 120.835 141.875 ;
        RECT 120.990 141.830 121.310 141.890 ;
        RECT 120.070 141.690 121.310 141.830 ;
        RECT 120.070 141.630 120.390 141.690 ;
        RECT 120.545 141.645 120.835 141.690 ;
        RECT 120.990 141.630 121.310 141.690 ;
        RECT 113.645 141.490 113.935 141.535 ;
        RECT 114.550 141.490 114.870 141.550 ;
        RECT 84.650 141.350 89.555 141.490 ;
        RECT 71.770 141.290 72.090 141.305 ;
        RECT 81.430 141.290 81.750 141.350 ;
        RECT 84.650 141.290 84.970 141.350 ;
        RECT 89.265 141.305 89.555 141.350 ;
        RECT 103.600 141.350 106.960 141.490 ;
        RECT 108.660 141.350 114.870 141.490 ;
        RECT 69.010 141.150 69.330 141.210 ;
        RECT 58.520 141.010 69.330 141.150 ;
        RECT 69.010 140.950 69.330 141.010 ;
        RECT 80.065 141.150 80.355 141.195 ;
        RECT 82.350 141.150 82.670 141.210 ;
        RECT 80.065 141.010 82.670 141.150 ;
        RECT 80.065 140.965 80.355 141.010 ;
        RECT 82.350 140.950 82.670 141.010 ;
        RECT 86.030 141.150 86.350 141.210 ;
        RECT 86.505 141.150 86.795 141.195 ;
        RECT 86.030 141.010 86.795 141.150 ;
        RECT 86.030 140.950 86.350 141.010 ;
        RECT 86.505 140.965 86.795 141.010 ;
        RECT 88.345 141.150 88.635 141.195 ;
        RECT 90.170 141.150 90.490 141.210 ;
        RECT 103.600 141.195 103.740 141.350 ;
        RECT 88.345 141.010 90.490 141.150 ;
        RECT 88.345 140.965 88.635 141.010 ;
        RECT 90.170 140.950 90.490 141.010 ;
        RECT 103.525 140.965 103.815 141.195 ;
        RECT 106.270 140.950 106.590 141.210 ;
        RECT 106.820 141.150 106.960 141.350 ;
        RECT 113.645 141.305 113.935 141.350 ;
        RECT 114.550 141.290 114.870 141.350 ;
        RECT 135.635 141.220 136.775 165.470 ;
        RECT 110.410 141.150 110.730 141.210 ;
        RECT 106.820 141.010 110.730 141.150 ;
        RECT 110.410 140.950 110.730 141.010 ;
        RECT 113.170 141.150 113.490 141.210 ;
        RECT 116.405 141.150 116.695 141.195 ;
        RECT 113.170 141.010 116.695 141.150 ;
        RECT 113.170 140.950 113.490 141.010 ;
        RECT 116.405 140.965 116.695 141.010 ;
        RECT 120.990 140.950 121.310 141.210 ;
        RECT 14.660 140.330 127.820 140.810 ;
        RECT 135.580 140.230 136.830 141.220 ;
        RECT 21.630 140.130 21.950 140.190 ;
        RECT 32.225 140.130 32.515 140.175 ;
        RECT 34.050 140.130 34.370 140.190 ;
        RECT 21.630 139.990 26.460 140.130 ;
        RECT 21.630 139.930 21.950 139.990 ;
        RECT 18.820 139.790 19.110 139.835 ;
        RECT 19.330 139.790 19.650 139.850 ;
        RECT 22.080 139.790 22.370 139.835 ;
        RECT 18.820 139.650 22.370 139.790 ;
        RECT 18.820 139.605 19.110 139.650 ;
        RECT 19.330 139.590 19.650 139.650 ;
        RECT 22.080 139.605 22.370 139.650 ;
        RECT 23.000 139.790 23.290 139.835 ;
        RECT 24.860 139.790 25.150 139.835 ;
        RECT 23.000 139.650 25.150 139.790 ;
        RECT 23.000 139.605 23.290 139.650 ;
        RECT 24.860 139.605 25.150 139.650 ;
        RECT 20.680 139.450 20.970 139.495 ;
        RECT 23.000 139.450 23.215 139.605 ;
        RECT 20.680 139.310 23.215 139.450 ;
        RECT 25.310 139.450 25.630 139.510 ;
        RECT 25.785 139.450 26.075 139.495 ;
        RECT 25.310 139.310 26.075 139.450 ;
        RECT 20.680 139.265 20.970 139.310 ;
        RECT 25.310 139.250 25.630 139.310 ;
        RECT 25.785 139.265 26.075 139.310 ;
        RECT 23.945 139.110 24.235 139.155 ;
        RECT 24.850 139.110 25.170 139.170 ;
        RECT 23.945 138.970 25.170 139.110 ;
        RECT 26.320 139.110 26.460 139.990 ;
        RECT 32.225 139.990 34.370 140.130 ;
        RECT 32.225 139.945 32.515 139.990 ;
        RECT 34.050 139.930 34.370 139.990 ;
        RECT 34.525 140.130 34.815 140.175 ;
        RECT 36.350 140.130 36.670 140.190 ;
        RECT 34.525 139.990 36.670 140.130 ;
        RECT 34.525 139.945 34.815 139.990 ;
        RECT 36.350 139.930 36.670 139.990 ;
        RECT 51.070 140.130 51.390 140.190 ;
        RECT 51.545 140.130 51.835 140.175 ;
        RECT 51.070 139.990 51.835 140.130 ;
        RECT 51.070 139.930 51.390 139.990 ;
        RECT 51.545 139.945 51.835 139.990 ;
        RECT 57.970 139.930 58.290 140.190 ;
        RECT 59.825 139.945 60.115 140.175 ;
        RECT 64.870 140.130 65.190 140.190 ;
        RECT 69.470 140.130 69.790 140.190 ;
        RECT 70.390 140.130 70.710 140.190 ;
        RECT 64.870 139.990 70.710 140.130 ;
        RECT 49.245 139.790 49.535 139.835 ;
        RECT 52.005 139.790 52.295 139.835 ;
        RECT 54.750 139.790 55.070 139.850 ;
        RECT 33.680 139.650 36.120 139.790 ;
        RECT 31.305 139.450 31.595 139.495 ;
        RECT 33.130 139.450 33.450 139.510 ;
        RECT 33.680 139.495 33.820 139.650 ;
        RECT 33.605 139.450 33.895 139.495 ;
        RECT 31.305 139.310 33.895 139.450 ;
        RECT 31.305 139.265 31.595 139.310 ;
        RECT 33.130 139.250 33.450 139.310 ;
        RECT 33.605 139.265 33.895 139.310 ;
        RECT 34.970 139.250 35.290 139.510 ;
        RECT 35.980 139.495 36.120 139.650 ;
        RECT 49.245 139.650 52.295 139.790 ;
        RECT 49.245 139.605 49.535 139.650 ;
        RECT 52.005 139.605 52.295 139.650 ;
        RECT 52.540 139.650 55.070 139.790 ;
        RECT 35.905 139.450 36.195 139.495 ;
        RECT 36.350 139.450 36.670 139.510 ;
        RECT 35.905 139.310 36.670 139.450 ;
        RECT 35.905 139.265 36.195 139.310 ;
        RECT 36.350 139.250 36.670 139.310 ;
        RECT 46.470 139.450 46.790 139.510 ;
        RECT 46.470 139.310 46.985 139.450 ;
        RECT 46.470 139.250 46.790 139.310 ;
        RECT 50.610 139.250 50.930 139.510 ;
        RECT 51.530 139.450 51.850 139.510 ;
        RECT 52.540 139.450 52.680 139.650 ;
        RECT 51.530 139.310 52.680 139.450 ;
        RECT 51.530 139.250 51.850 139.310 ;
        RECT 53.370 139.250 53.690 139.510 ;
        RECT 53.920 139.495 54.060 139.650 ;
        RECT 54.750 139.590 55.070 139.650 ;
        RECT 57.510 139.590 57.830 139.850 ;
        RECT 53.845 139.265 54.135 139.495 ;
        RECT 54.305 139.265 54.595 139.495 ;
        RECT 30.385 139.110 30.675 139.155 ;
        RECT 26.320 138.970 30.675 139.110 ;
        RECT 23.945 138.925 24.235 138.970 ;
        RECT 24.850 138.910 25.170 138.970 ;
        RECT 30.385 138.925 30.675 138.970 ;
        RECT 32.685 138.925 32.975 139.155 ;
        RECT 36.825 139.110 37.115 139.155 ;
        RECT 39.110 139.110 39.430 139.170 ;
        RECT 36.825 138.970 39.430 139.110 ;
        RECT 36.825 138.925 37.115 138.970 ;
        RECT 20.680 138.770 20.970 138.815 ;
        RECT 23.460 138.770 23.750 138.815 ;
        RECT 25.320 138.770 25.610 138.815 ;
        RECT 20.680 138.630 25.610 138.770 ;
        RECT 20.680 138.585 20.970 138.630 ;
        RECT 23.460 138.585 23.750 138.630 ;
        RECT 25.320 138.585 25.610 138.630 ;
        RECT 29.910 138.770 30.230 138.830 ;
        RECT 32.760 138.770 32.900 138.925 ;
        RECT 39.110 138.910 39.430 138.970 ;
        RECT 42.330 139.110 42.650 139.170 ;
        RECT 45.565 139.110 45.855 139.155 ;
        RECT 42.330 138.970 45.855 139.110 ;
        RECT 42.330 138.910 42.650 138.970 ;
        RECT 45.565 138.925 45.855 138.970 ;
        RECT 46.930 139.110 47.250 139.170 ;
        RECT 49.705 139.110 49.995 139.155 ;
        RECT 46.930 138.970 49.995 139.110 ;
        RECT 46.930 138.910 47.250 138.970 ;
        RECT 49.705 138.925 49.995 138.970 ;
        RECT 29.910 138.630 32.900 138.770 ;
        RECT 54.380 138.770 54.520 139.265 ;
        RECT 55.210 139.250 55.530 139.510 ;
        RECT 57.600 139.450 57.740 139.590 ;
        RECT 57.140 139.310 57.740 139.450 ;
        RECT 59.900 139.450 60.040 139.945 ;
        RECT 64.870 139.930 65.190 139.990 ;
        RECT 69.470 139.930 69.790 139.990 ;
        RECT 70.390 139.930 70.710 139.990 ;
        RECT 71.770 140.130 72.090 140.190 ;
        RECT 72.705 140.130 72.995 140.175 ;
        RECT 71.770 139.990 72.995 140.130 ;
        RECT 71.770 139.930 72.090 139.990 ;
        RECT 72.705 139.945 72.995 139.990 ;
        RECT 79.375 140.130 79.665 140.175 ;
        RECT 82.810 140.130 83.130 140.190 ;
        RECT 79.375 139.990 83.130 140.130 ;
        RECT 79.375 139.945 79.665 139.990 ;
        RECT 82.810 139.930 83.130 139.990 ;
        RECT 89.265 139.945 89.555 140.175 ;
        RECT 68.550 139.790 68.870 139.850 ;
        RECT 80.510 139.790 80.830 139.850 ;
        RECT 84.650 139.835 84.970 139.850 ;
        RECT 68.550 139.650 80.830 139.790 ;
        RECT 68.550 139.590 68.870 139.650 ;
        RECT 80.510 139.590 80.830 139.650 ;
        RECT 81.380 139.790 81.670 139.835 ;
        RECT 84.640 139.790 84.970 139.835 ;
        RECT 81.380 139.650 84.970 139.790 ;
        RECT 81.380 139.605 81.670 139.650 ;
        RECT 84.640 139.605 84.970 139.650 ;
        RECT 84.650 139.590 84.970 139.605 ;
        RECT 85.560 139.790 85.850 139.835 ;
        RECT 87.420 139.790 87.710 139.835 ;
        RECT 85.560 139.650 87.710 139.790 ;
        RECT 85.560 139.605 85.850 139.650 ;
        RECT 87.420 139.605 87.710 139.650 ;
        RECT 60.285 139.450 60.575 139.495 ;
        RECT 68.640 139.450 68.780 139.590 ;
        RECT 59.900 139.310 60.575 139.450 ;
        RECT 57.140 139.155 57.280 139.310 ;
        RECT 60.285 139.265 60.575 139.310 ;
        RECT 60.820 139.310 68.780 139.450 ;
        RECT 72.690 139.450 73.010 139.510 ;
        RECT 73.165 139.450 73.455 139.495 ;
        RECT 72.690 139.310 73.455 139.450 ;
        RECT 57.065 138.925 57.355 139.155 ;
        RECT 57.525 139.110 57.815 139.155 ;
        RECT 58.890 139.110 59.210 139.170 ;
        RECT 57.525 138.970 59.210 139.110 ;
        RECT 57.525 138.925 57.815 138.970 ;
        RECT 57.600 138.770 57.740 138.925 ;
        RECT 58.890 138.910 59.210 138.970 ;
        RECT 54.380 138.630 57.740 138.770 ;
        RECT 29.910 138.570 30.230 138.630 ;
        RECT 16.815 138.430 17.105 138.475 ;
        RECT 22.090 138.430 22.410 138.490 ;
        RECT 34.970 138.430 35.290 138.490 ;
        RECT 16.815 138.290 35.290 138.430 ;
        RECT 16.815 138.245 17.105 138.290 ;
        RECT 22.090 138.230 22.410 138.290 ;
        RECT 34.970 138.230 35.290 138.290 ;
        RECT 47.405 138.430 47.695 138.475 ;
        RECT 49.245 138.430 49.535 138.475 ;
        RECT 47.405 138.290 49.535 138.430 ;
        RECT 47.405 138.245 47.695 138.290 ;
        RECT 49.245 138.245 49.535 138.290 ;
        RECT 55.210 138.430 55.530 138.490 ;
        RECT 60.820 138.430 60.960 139.310 ;
        RECT 72.690 139.250 73.010 139.310 ;
        RECT 73.165 139.265 73.455 139.310 ;
        RECT 75.450 139.450 75.770 139.510 ;
        RECT 83.240 139.450 83.530 139.495 ;
        RECT 85.560 139.450 85.775 139.605 ;
        RECT 75.450 139.310 78.440 139.450 ;
        RECT 75.450 139.250 75.770 139.310 ;
        RECT 78.300 139.110 78.440 139.310 ;
        RECT 83.240 139.310 85.775 139.450 ;
        RECT 86.505 139.450 86.795 139.495 ;
        RECT 89.340 139.450 89.480 139.945 ;
        RECT 98.910 139.930 99.230 140.190 ;
        RECT 103.510 139.930 103.830 140.190 ;
        RECT 109.030 140.130 109.350 140.190 ;
        RECT 105.440 139.990 109.350 140.130 ;
        RECT 96.625 139.790 96.915 139.835 ;
        RECT 99.385 139.790 99.675 139.835 ;
        RECT 96.625 139.650 99.675 139.790 ;
        RECT 96.625 139.605 96.915 139.650 ;
        RECT 99.385 139.605 99.675 139.650 ;
        RECT 100.290 139.790 100.610 139.850 ;
        RECT 105.440 139.790 105.580 139.990 ;
        RECT 109.030 139.930 109.350 139.990 ;
        RECT 114.090 140.130 114.410 140.190 ;
        RECT 116.635 140.130 116.925 140.175 ;
        RECT 120.070 140.130 120.390 140.190 ;
        RECT 135.635 140.155 136.775 140.230 ;
        RECT 114.090 139.990 116.925 140.130 ;
        RECT 114.090 139.930 114.410 139.990 ;
        RECT 116.635 139.945 116.925 139.990 ;
        RECT 118.320 139.990 120.390 140.130 ;
        RECT 100.290 139.650 101.440 139.790 ;
        RECT 100.290 139.590 100.610 139.650 ;
        RECT 86.505 139.310 89.480 139.450 ;
        RECT 83.240 139.265 83.530 139.310 ;
        RECT 86.505 139.265 86.795 139.310 ;
        RECT 90.170 139.250 90.490 139.510 ;
        RECT 97.990 139.250 98.310 139.510 ;
        RECT 100.750 139.250 101.070 139.510 ;
        RECT 101.300 139.495 101.440 139.650 ;
        RECT 102.680 139.650 105.580 139.790 ;
        RECT 105.825 139.790 106.115 139.835 ;
        RECT 106.270 139.790 106.590 139.850 ;
        RECT 105.825 139.650 106.590 139.790 ;
        RECT 101.225 139.265 101.515 139.495 ;
        RECT 101.670 139.250 101.990 139.510 ;
        RECT 102.130 139.450 102.450 139.510 ;
        RECT 102.680 139.495 102.820 139.650 ;
        RECT 105.825 139.605 106.115 139.650 ;
        RECT 106.270 139.590 106.590 139.650 ;
        RECT 109.505 139.790 109.795 139.835 ;
        RECT 114.550 139.790 114.870 139.850 ;
        RECT 109.505 139.650 114.870 139.790 ;
        RECT 109.505 139.605 109.795 139.650 ;
        RECT 114.550 139.590 114.870 139.650 ;
        RECT 102.605 139.450 102.895 139.495 ;
        RECT 102.130 139.310 102.895 139.450 ;
        RECT 102.130 139.250 102.450 139.310 ;
        RECT 102.605 139.265 102.895 139.310 ;
        RECT 103.050 139.450 103.370 139.510 ;
        RECT 104.445 139.450 104.735 139.495 ;
        RECT 112.250 139.450 112.570 139.510 ;
        RECT 103.050 139.310 104.735 139.450 ;
        RECT 103.050 139.250 103.370 139.310 ;
        RECT 104.445 139.265 104.735 139.310 ;
        RECT 108.200 139.310 112.570 139.450 ;
        RECT 108.200 139.170 108.340 139.310 ;
        RECT 112.250 139.250 112.570 139.310 ;
        RECT 113.170 139.250 113.490 139.510 ;
        RECT 115.025 139.265 115.315 139.495 ;
        RECT 88.345 139.110 88.635 139.155 ;
        RECT 95.230 139.110 95.550 139.170 ;
        RECT 78.300 138.970 95.550 139.110 ;
        RECT 88.345 138.925 88.635 138.970 ;
        RECT 95.230 138.910 95.550 138.970 ;
        RECT 97.070 138.910 97.390 139.170 ;
        RECT 104.905 139.110 105.195 139.155 ;
        RECT 101.300 138.970 105.195 139.110 ;
        RECT 101.300 138.830 101.440 138.970 ;
        RECT 104.905 138.925 105.195 138.970 ;
        RECT 108.110 138.910 108.430 139.170 ;
        RECT 109.045 138.925 109.335 139.155 ;
        RECT 115.100 139.110 115.240 139.265 ;
        RECT 115.470 139.250 115.790 139.510 ;
        RECT 118.320 139.110 118.460 139.990 ;
        RECT 120.070 139.930 120.390 139.990 ;
        RECT 118.640 139.790 118.930 139.835 ;
        RECT 120.990 139.790 121.310 139.850 ;
        RECT 121.900 139.790 122.190 139.835 ;
        RECT 118.640 139.650 122.190 139.790 ;
        RECT 118.640 139.605 118.930 139.650 ;
        RECT 120.990 139.590 121.310 139.650 ;
        RECT 121.900 139.605 122.190 139.650 ;
        RECT 122.820 139.790 123.110 139.835 ;
        RECT 124.680 139.790 124.970 139.835 ;
        RECT 122.820 139.650 124.970 139.790 ;
        RECT 122.820 139.605 123.110 139.650 ;
        RECT 124.680 139.605 124.970 139.650 ;
        RECT 120.500 139.450 120.790 139.495 ;
        RECT 122.820 139.450 123.035 139.605 ;
        RECT 120.500 139.310 123.035 139.450 ;
        RECT 120.500 139.265 120.790 139.310 ;
        RECT 129.090 139.190 134.150 139.405 ;
        RECT 143.370 139.390 144.510 223.840 ;
        RECT 137.240 139.380 144.510 139.390 ;
        RECT 136.210 139.190 144.510 139.380 ;
        RECT 123.765 139.110 124.055 139.155 ;
        RECT 115.100 138.970 118.460 139.110 ;
        RECT 119.470 138.970 124.055 139.110 ;
        RECT 83.240 138.770 83.530 138.815 ;
        RECT 86.020 138.770 86.310 138.815 ;
        RECT 87.880 138.770 88.170 138.815 ;
        RECT 83.240 138.630 88.170 138.770 ;
        RECT 83.240 138.585 83.530 138.630 ;
        RECT 86.020 138.585 86.310 138.630 ;
        RECT 87.880 138.585 88.170 138.630 ;
        RECT 101.210 138.570 101.530 138.830 ;
        RECT 101.670 138.770 101.990 138.830 ;
        RECT 109.120 138.770 109.260 138.925 ;
        RECT 101.670 138.630 109.260 138.770 ;
        RECT 114.105 138.770 114.395 138.815 ;
        RECT 119.470 138.770 119.610 138.970 ;
        RECT 123.765 138.925 124.055 138.970 ;
        RECT 125.590 138.910 125.910 139.170 ;
        RECT 114.105 138.630 119.610 138.770 ;
        RECT 120.500 138.770 120.790 138.815 ;
        RECT 123.280 138.770 123.570 138.815 ;
        RECT 125.140 138.770 125.430 138.815 ;
        RECT 120.500 138.630 125.430 138.770 ;
        RECT 101.670 138.570 101.990 138.630 ;
        RECT 114.105 138.585 114.395 138.630 ;
        RECT 120.500 138.585 120.790 138.630 ;
        RECT 123.280 138.585 123.570 138.630 ;
        RECT 125.140 138.585 125.430 138.630 ;
        RECT 129.090 138.530 144.510 139.190 ;
        RECT 55.210 138.290 60.960 138.430 ;
        RECT 55.210 138.230 55.530 138.290 ;
        RECT 61.190 138.230 61.510 138.490 ;
        RECT 97.530 138.230 97.850 138.490 ;
        RECT 105.350 138.230 105.670 138.490 ;
        RECT 111.330 138.230 111.650 138.490 ;
        RECT 129.090 138.225 134.150 138.530 ;
        RECT 136.210 138.250 144.510 138.530 ;
        RECT 136.210 138.240 138.350 138.250 ;
        RECT 14.660 137.610 127.820 138.090 ;
        RECT 17.965 137.410 18.255 137.455 ;
        RECT 18.870 137.410 19.190 137.470 ;
        RECT 17.965 137.270 19.190 137.410 ;
        RECT 17.965 137.225 18.255 137.270 ;
        RECT 18.870 137.210 19.190 137.270 ;
        RECT 19.330 137.210 19.650 137.470 ;
        RECT 24.850 137.210 25.170 137.470 ;
        RECT 26.230 137.410 26.550 137.470 ;
        RECT 46.010 137.410 46.330 137.470 ;
        RECT 46.945 137.410 47.235 137.455 ;
        RECT 26.230 137.270 29.220 137.410 ;
        RECT 26.230 137.210 26.550 137.270 ;
        RECT 29.080 137.070 29.220 137.270 ;
        RECT 46.010 137.270 47.235 137.410 ;
        RECT 46.010 137.210 46.330 137.270 ;
        RECT 46.945 137.225 47.235 137.270 ;
        RECT 114.550 137.410 114.870 137.470 ;
        RECT 116.175 137.410 116.465 137.455 ;
        RECT 114.550 137.270 116.465 137.410 ;
        RECT 114.550 137.210 114.870 137.270 ;
        RECT 116.175 137.225 116.465 137.270 ;
        RECT 36.320 137.070 36.610 137.115 ;
        RECT 39.100 137.070 39.390 137.115 ;
        RECT 40.960 137.070 41.250 137.115 ;
        RECT 21.260 136.930 22.320 137.070 ;
        RECT 21.260 136.775 21.400 136.930 ;
        RECT 21.185 136.545 21.475 136.775 ;
        RECT 21.630 136.530 21.950 136.790 ;
        RECT 22.180 136.730 22.320 136.930 ;
        RECT 29.080 136.930 35.660 137.070 ;
        RECT 23.010 136.730 23.330 136.790 ;
        RECT 26.230 136.730 26.550 136.790 ;
        RECT 29.080 136.775 29.220 136.930 ;
        RECT 22.180 136.590 26.550 136.730 ;
        RECT 23.010 136.530 23.330 136.590 ;
        RECT 26.230 136.530 26.550 136.590 ;
        RECT 29.005 136.545 29.295 136.775 ;
        RECT 29.465 136.730 29.755 136.775 ;
        RECT 34.970 136.730 35.290 136.790 ;
        RECT 29.465 136.590 35.290 136.730 ;
        RECT 35.520 136.730 35.660 136.930 ;
        RECT 36.320 136.930 41.250 137.070 ;
        RECT 36.320 136.885 36.610 136.930 ;
        RECT 39.100 136.885 39.390 136.930 ;
        RECT 40.960 136.885 41.250 136.930 ;
        RECT 58.400 137.070 58.690 137.115 ;
        RECT 61.180 137.070 61.470 137.115 ;
        RECT 63.040 137.070 63.330 137.115 ;
        RECT 58.400 136.930 63.330 137.070 ;
        RECT 58.400 136.885 58.690 136.930 ;
        RECT 61.180 136.885 61.470 136.930 ;
        RECT 63.040 136.885 63.330 136.930 ;
        RECT 83.730 136.870 84.050 137.130 ;
        RECT 85.110 137.070 85.430 137.130 ;
        RECT 108.110 137.070 108.430 137.130 ;
        RECT 85.110 136.930 108.430 137.070 ;
        RECT 85.110 136.870 85.430 136.930 ;
        RECT 37.270 136.730 37.590 136.790 ;
        RECT 43.725 136.730 44.015 136.775 ;
        RECT 35.520 136.590 44.015 136.730 ;
        RECT 29.465 136.545 29.755 136.590 ;
        RECT 34.970 136.530 35.290 136.590 ;
        RECT 37.270 136.530 37.590 136.590 ;
        RECT 43.725 136.545 44.015 136.590 ;
        RECT 59.810 136.730 60.130 136.790 ;
        RECT 63.505 136.730 63.795 136.775 ;
        RECT 59.810 136.590 63.795 136.730 ;
        RECT 83.820 136.730 83.960 136.870 ;
        RECT 97.160 136.775 97.300 136.930 ;
        RECT 108.110 136.870 108.430 136.930 ;
        RECT 109.000 137.070 109.290 137.115 ;
        RECT 111.780 137.070 112.070 137.115 ;
        RECT 113.640 137.070 113.930 137.115 ;
        RECT 109.000 136.930 113.930 137.070 ;
        RECT 109.000 136.885 109.290 136.930 ;
        RECT 111.780 136.885 112.070 136.930 ;
        RECT 113.640 136.885 113.930 136.930 ;
        RECT 120.040 137.070 120.330 137.115 ;
        RECT 122.820 137.070 123.110 137.115 ;
        RECT 124.680 137.070 124.970 137.115 ;
        RECT 120.040 136.930 124.970 137.070 ;
        RECT 120.040 136.885 120.330 136.930 ;
        RECT 122.820 136.885 123.110 136.930 ;
        RECT 124.680 136.885 124.970 136.930 ;
        RECT 83.820 136.590 85.340 136.730 ;
        RECT 59.810 136.530 60.130 136.590 ;
        RECT 63.505 136.545 63.795 136.590 ;
        RECT 17.505 136.390 17.795 136.435 ;
        RECT 18.885 136.390 19.175 136.435 ;
        RECT 17.505 136.250 19.175 136.390 ;
        RECT 17.505 136.205 17.795 136.250 ;
        RECT 18.885 136.205 19.175 136.250 ;
        RECT 18.960 136.050 19.100 136.205 ;
        RECT 22.090 136.190 22.410 136.450 ;
        RECT 25.770 136.190 26.090 136.450 ;
        RECT 26.705 136.390 26.995 136.435 ;
        RECT 31.750 136.390 32.070 136.450 ;
        RECT 26.705 136.250 32.070 136.390 ;
        RECT 26.705 136.205 26.995 136.250 ;
        RECT 26.780 136.050 26.920 136.205 ;
        RECT 31.750 136.190 32.070 136.250 ;
        RECT 36.320 136.390 36.610 136.435 ;
        RECT 39.110 136.390 39.430 136.450 ;
        RECT 39.585 136.390 39.875 136.435 ;
        RECT 36.320 136.250 38.855 136.390 ;
        RECT 36.320 136.205 36.610 136.250 ;
        RECT 18.960 135.910 26.920 136.050 ;
        RECT 34.460 136.050 34.750 136.095 ;
        RECT 35.890 136.050 36.210 136.110 ;
        RECT 38.640 136.095 38.855 136.250 ;
        RECT 39.110 136.250 39.875 136.390 ;
        RECT 39.110 136.190 39.430 136.250 ;
        RECT 39.585 136.205 39.875 136.250 ;
        RECT 41.410 136.190 41.730 136.450 ;
        RECT 42.330 136.390 42.650 136.450 ;
        RECT 44.645 136.390 44.935 136.435 ;
        RECT 42.330 136.250 44.935 136.390 ;
        RECT 42.330 136.190 42.650 136.250 ;
        RECT 44.645 136.205 44.935 136.250 ;
        RECT 46.010 136.390 46.330 136.450 ;
        RECT 47.865 136.390 48.155 136.435 ;
        RECT 46.010 136.250 48.155 136.390 ;
        RECT 46.010 136.190 46.330 136.250 ;
        RECT 47.865 136.205 48.155 136.250 ;
        RECT 48.325 136.205 48.615 136.435 ;
        RECT 58.400 136.390 58.690 136.435 ;
        RECT 61.190 136.390 61.510 136.450 ;
        RECT 61.665 136.390 61.955 136.435 ;
        RECT 58.400 136.250 60.935 136.390 ;
        RECT 58.400 136.205 58.690 136.250 ;
        RECT 37.720 136.050 38.010 136.095 ;
        RECT 34.460 135.910 38.010 136.050 ;
        RECT 34.460 135.865 34.750 135.910 ;
        RECT 35.890 135.850 36.210 135.910 ;
        RECT 37.720 135.865 38.010 135.910 ;
        RECT 38.640 136.050 38.930 136.095 ;
        RECT 40.500 136.050 40.790 136.095 ;
        RECT 48.400 136.050 48.540 136.205 ;
        RECT 38.640 135.910 40.790 136.050 ;
        RECT 38.640 135.865 38.930 135.910 ;
        RECT 40.500 135.865 40.790 135.910 ;
        RECT 44.260 135.910 48.540 136.050 ;
        RECT 56.540 136.050 56.830 136.095 ;
        RECT 57.970 136.050 58.290 136.110 ;
        RECT 60.720 136.095 60.935 136.250 ;
        RECT 61.190 136.250 61.955 136.390 ;
        RECT 61.190 136.190 61.510 136.250 ;
        RECT 61.665 136.205 61.955 136.250 ;
        RECT 81.890 136.390 82.210 136.450 ;
        RECT 83.285 136.390 83.575 136.435 ;
        RECT 81.890 136.250 83.575 136.390 ;
        RECT 81.890 136.190 82.210 136.250 ;
        RECT 83.285 136.205 83.575 136.250 ;
        RECT 83.745 136.205 84.035 136.435 ;
        RECT 84.205 136.390 84.495 136.435 ;
        RECT 84.650 136.390 84.970 136.450 ;
        RECT 85.200 136.435 85.340 136.590 ;
        RECT 97.085 136.545 97.375 136.775 ;
        RECT 112.250 136.530 112.570 136.790 ;
        RECT 119.470 136.590 123.060 136.730 ;
        RECT 84.205 136.250 84.970 136.390 ;
        RECT 84.205 136.205 84.495 136.250 ;
        RECT 59.800 136.050 60.090 136.095 ;
        RECT 56.540 135.910 60.090 136.050 ;
        RECT 23.945 135.710 24.235 135.755 ;
        RECT 25.770 135.710 26.090 135.770 ;
        RECT 23.945 135.570 26.090 135.710 ;
        RECT 23.945 135.525 24.235 135.570 ;
        RECT 25.770 135.510 26.090 135.570 ;
        RECT 27.150 135.510 27.470 135.770 ;
        RECT 29.910 135.510 30.230 135.770 ;
        RECT 31.290 135.710 31.610 135.770 ;
        RECT 31.765 135.710 32.055 135.755 ;
        RECT 31.290 135.570 32.055 135.710 ;
        RECT 31.290 135.510 31.610 135.570 ;
        RECT 31.765 135.525 32.055 135.570 ;
        RECT 32.455 135.710 32.745 135.755 ;
        RECT 36.810 135.710 37.130 135.770 ;
        RECT 44.260 135.755 44.400 135.910 ;
        RECT 56.540 135.865 56.830 135.910 ;
        RECT 57.970 135.850 58.290 135.910 ;
        RECT 59.800 135.865 60.090 135.910 ;
        RECT 60.720 136.050 61.010 136.095 ;
        RECT 62.580 136.050 62.870 136.095 ;
        RECT 60.720 135.910 62.870 136.050 ;
        RECT 60.720 135.865 61.010 135.910 ;
        RECT 62.580 135.865 62.870 135.910 ;
        RECT 81.430 136.050 81.750 136.110 ;
        RECT 83.820 136.050 83.960 136.205 ;
        RECT 84.650 136.190 84.970 136.250 ;
        RECT 85.125 136.205 85.415 136.435 ;
        RECT 98.465 136.390 98.755 136.435 ;
        RECT 101.670 136.390 101.990 136.450 ;
        RECT 105.135 136.390 105.425 136.435 ;
        RECT 98.465 136.250 105.425 136.390 ;
        RECT 98.465 136.205 98.755 136.250 ;
        RECT 101.670 136.190 101.990 136.250 ;
        RECT 105.135 136.205 105.425 136.250 ;
        RECT 109.000 136.390 109.290 136.435 ;
        RECT 111.790 136.390 112.110 136.450 ;
        RECT 114.105 136.390 114.395 136.435 ;
        RECT 119.470 136.390 119.610 136.590 ;
        RECT 109.000 136.250 111.535 136.390 ;
        RECT 109.000 136.205 109.290 136.250 ;
        RECT 81.430 135.910 83.960 136.050 ;
        RECT 107.140 136.050 107.430 136.095 ;
        RECT 109.490 136.050 109.810 136.110 ;
        RECT 111.320 136.095 111.535 136.250 ;
        RECT 111.790 136.250 119.610 136.390 ;
        RECT 120.040 136.390 120.330 136.435 ;
        RECT 122.920 136.390 123.060 136.590 ;
        RECT 123.290 136.530 123.610 136.790 ;
        RECT 125.145 136.730 125.435 136.775 ;
        RECT 125.590 136.730 125.910 136.790 ;
        RECT 125.145 136.590 125.910 136.730 ;
        RECT 125.145 136.545 125.435 136.590 ;
        RECT 125.220 136.390 125.360 136.545 ;
        RECT 125.590 136.530 125.910 136.590 ;
        RECT 120.040 136.250 122.575 136.390 ;
        RECT 122.920 136.250 125.360 136.390 ;
        RECT 111.790 136.190 112.110 136.250 ;
        RECT 114.105 136.205 114.395 136.250 ;
        RECT 120.040 136.205 120.330 136.250 ;
        RECT 110.400 136.050 110.690 136.095 ;
        RECT 107.140 135.910 110.690 136.050 ;
        RECT 81.430 135.850 81.750 135.910 ;
        RECT 107.140 135.865 107.430 135.910 ;
        RECT 109.490 135.850 109.810 135.910 ;
        RECT 110.400 135.865 110.690 135.910 ;
        RECT 111.320 136.050 111.610 136.095 ;
        RECT 113.180 136.050 113.470 136.095 ;
        RECT 111.320 135.910 113.470 136.050 ;
        RECT 111.320 135.865 111.610 135.910 ;
        RECT 113.180 135.865 113.470 135.910 ;
        RECT 115.470 136.050 115.790 136.110 ;
        RECT 122.360 136.095 122.575 136.250 ;
        RECT 118.180 136.050 118.470 136.095 ;
        RECT 121.440 136.050 121.730 136.095 ;
        RECT 115.470 135.910 121.730 136.050 ;
        RECT 115.470 135.850 115.790 135.910 ;
        RECT 118.180 135.865 118.470 135.910 ;
        RECT 121.440 135.865 121.730 135.910 ;
        RECT 122.360 136.050 122.650 136.095 ;
        RECT 124.220 136.050 124.510 136.095 ;
        RECT 122.360 135.910 124.510 136.050 ;
        RECT 122.360 135.865 122.650 135.910 ;
        RECT 124.220 135.865 124.510 135.910 ;
        RECT 44.185 135.710 44.475 135.755 ;
        RECT 32.455 135.570 44.475 135.710 ;
        RECT 32.455 135.525 32.745 135.570 ;
        RECT 36.810 135.510 37.130 135.570 ;
        RECT 44.185 135.525 44.475 135.570 ;
        RECT 45.550 135.710 45.870 135.770 ;
        RECT 46.485 135.710 46.775 135.755 ;
        RECT 45.550 135.570 46.775 135.710 ;
        RECT 45.550 135.510 45.870 135.570 ;
        RECT 46.485 135.525 46.775 135.570 ;
        RECT 54.535 135.710 54.825 135.755 ;
        RECT 58.890 135.710 59.210 135.770 ;
        RECT 54.535 135.570 59.210 135.710 ;
        RECT 54.535 135.525 54.825 135.570 ;
        RECT 58.890 135.510 59.210 135.570 ;
        RECT 81.890 135.510 82.210 135.770 ;
        RECT 97.990 135.510 98.310 135.770 ;
        RECT 100.305 135.710 100.595 135.755 ;
        RECT 103.050 135.710 103.370 135.770 ;
        RECT 100.305 135.570 103.370 135.710 ;
        RECT 100.305 135.525 100.595 135.570 ;
        RECT 103.050 135.510 103.370 135.570 ;
        RECT 14.660 134.890 127.820 135.370 ;
        RECT 19.345 134.690 19.635 134.735 ;
        RECT 21.170 134.690 21.490 134.750 ;
        RECT 19.345 134.550 21.490 134.690 ;
        RECT 19.345 134.505 19.635 134.550 ;
        RECT 21.170 134.490 21.490 134.550 ;
        RECT 21.630 134.490 21.950 134.750 ;
        RECT 24.175 134.690 24.465 134.735 ;
        RECT 29.910 134.690 30.230 134.750 ;
        RECT 24.175 134.550 30.230 134.690 ;
        RECT 24.175 134.505 24.465 134.550 ;
        RECT 29.910 134.490 30.230 134.550 ;
        RECT 35.890 134.490 36.210 134.750 ;
        RECT 39.110 134.490 39.430 134.750 ;
        RECT 57.970 134.490 58.290 134.750 ;
        RECT 69.470 134.490 69.790 134.750 ;
        RECT 78.225 134.690 78.515 134.735 ;
        RECT 81.430 134.690 81.750 134.750 ;
        RECT 86.030 134.690 86.350 134.750 ;
        RECT 78.225 134.550 80.280 134.690 ;
        RECT 78.225 134.505 78.515 134.550 ;
        RECT 26.180 134.350 26.470 134.395 ;
        RECT 27.150 134.350 27.470 134.410 ;
        RECT 29.440 134.350 29.730 134.395 ;
        RECT 26.180 134.210 29.730 134.350 ;
        RECT 26.180 134.165 26.470 134.210 ;
        RECT 27.150 134.150 27.470 134.210 ;
        RECT 29.440 134.165 29.730 134.210 ;
        RECT 30.360 134.350 30.650 134.395 ;
        RECT 32.220 134.350 32.510 134.395 ;
        RECT 30.360 134.210 32.510 134.350 ;
        RECT 30.360 134.165 30.650 134.210 ;
        RECT 32.220 134.165 32.510 134.210 ;
        RECT 41.820 134.350 42.110 134.395 ;
        RECT 43.250 134.350 43.570 134.410 ;
        RECT 45.080 134.350 45.370 134.395 ;
        RECT 41.820 134.210 45.370 134.350 ;
        RECT 41.820 134.165 42.110 134.210 ;
        RECT 18.425 134.010 18.715 134.055 ;
        RECT 28.040 134.010 28.330 134.055 ;
        RECT 30.360 134.010 30.575 134.165 ;
        RECT 43.250 134.150 43.570 134.210 ;
        RECT 45.080 134.165 45.370 134.210 ;
        RECT 46.000 134.350 46.290 134.395 ;
        RECT 47.860 134.350 48.150 134.395 ;
        RECT 46.000 134.210 48.150 134.350 ;
        RECT 46.000 134.165 46.290 134.210 ;
        RECT 47.860 134.165 48.150 134.210 ;
        RECT 67.185 134.350 67.475 134.395 ;
        RECT 68.090 134.350 68.410 134.410 ;
        RECT 70.390 134.350 70.710 134.410 ;
        RECT 72.705 134.350 72.995 134.395 ;
        RECT 67.185 134.210 72.995 134.350 ;
        RECT 67.185 134.165 67.475 134.210 ;
        RECT 18.425 133.870 20.020 134.010 ;
        RECT 18.425 133.825 18.715 133.870 ;
        RECT 19.880 133.375 20.020 133.870 ;
        RECT 28.040 133.870 30.575 134.010 ;
        RECT 30.830 134.010 31.150 134.070 ;
        RECT 31.305 134.010 31.595 134.055 ;
        RECT 30.830 133.870 31.595 134.010 ;
        RECT 28.040 133.825 28.330 133.870 ;
        RECT 30.830 133.810 31.150 133.870 ;
        RECT 31.305 133.825 31.595 133.870 ;
        RECT 31.750 134.010 32.070 134.070 ;
        RECT 35.445 134.010 35.735 134.055 ;
        RECT 37.730 134.010 38.050 134.070 ;
        RECT 31.750 133.870 38.050 134.010 ;
        RECT 31.750 133.810 32.070 133.870 ;
        RECT 35.445 133.825 35.735 133.870 ;
        RECT 37.730 133.810 38.050 133.870 ;
        RECT 38.190 133.810 38.510 134.070 ;
        RECT 43.680 134.010 43.970 134.055 ;
        RECT 46.000 134.010 46.215 134.165 ;
        RECT 68.090 134.150 68.410 134.210 ;
        RECT 70.390 134.150 70.710 134.210 ;
        RECT 72.705 134.165 72.995 134.210 ;
        RECT 43.680 133.870 46.215 134.010 ;
        RECT 53.830 134.010 54.150 134.070 ;
        RECT 55.670 134.010 55.990 134.070 ;
        RECT 57.525 134.010 57.815 134.055 ;
        RECT 53.830 133.870 57.815 134.010 ;
        RECT 43.680 133.825 43.970 133.870 ;
        RECT 53.830 133.810 54.150 133.870 ;
        RECT 55.670 133.810 55.990 133.870 ;
        RECT 57.525 133.825 57.815 133.870 ;
        RECT 66.250 134.010 66.570 134.070 ;
        RECT 69.945 134.010 70.235 134.055 ;
        RECT 66.250 133.870 70.235 134.010 ;
        RECT 66.250 133.810 66.570 133.870 ;
        RECT 69.945 133.825 70.235 133.870 ;
        RECT 79.145 134.010 79.435 134.055 ;
        RECT 79.590 134.010 79.910 134.070 ;
        RECT 79.145 133.870 79.910 134.010 ;
        RECT 80.140 134.010 80.280 134.550 ;
        RECT 81.430 134.550 82.580 134.690 ;
        RECT 81.430 134.490 81.750 134.550 ;
        RECT 80.525 134.350 80.815 134.395 ;
        RECT 81.890 134.350 82.210 134.410 ;
        RECT 80.525 134.210 82.210 134.350 ;
        RECT 82.440 134.350 82.580 134.550 ;
        RECT 83.360 134.550 86.350 134.690 ;
        RECT 82.440 134.210 83.040 134.350 ;
        RECT 80.525 134.165 80.815 134.210 ;
        RECT 81.890 134.150 82.210 134.210 ;
        RECT 80.140 133.870 81.660 134.010 ;
        RECT 79.145 133.825 79.435 133.870 ;
        RECT 79.590 133.810 79.910 133.870 ;
        RECT 20.710 133.670 21.030 133.730 ;
        RECT 22.090 133.670 22.410 133.730 ;
        RECT 20.710 133.530 22.410 133.670 ;
        RECT 20.710 133.470 21.030 133.530 ;
        RECT 22.090 133.470 22.410 133.530 ;
        RECT 23.010 133.470 23.330 133.730 ;
        RECT 25.310 133.670 25.630 133.730 ;
        RECT 33.145 133.670 33.435 133.715 ;
        RECT 41.410 133.670 41.730 133.730 ;
        RECT 25.310 133.530 41.730 133.670 ;
        RECT 25.310 133.470 25.630 133.530 ;
        RECT 33.145 133.485 33.435 133.530 ;
        RECT 41.410 133.470 41.730 133.530 ;
        RECT 46.930 133.470 47.250 133.730 ;
        RECT 48.785 133.670 49.075 133.715 ;
        RECT 60.270 133.670 60.590 133.730 ;
        RECT 48.785 133.530 60.590 133.670 ;
        RECT 48.785 133.485 49.075 133.530 ;
        RECT 60.270 133.470 60.590 133.530 ;
        RECT 69.010 133.470 69.330 133.730 ;
        RECT 80.050 133.470 80.370 133.730 ;
        RECT 81.520 133.670 81.660 133.870 ;
        RECT 82.350 133.810 82.670 134.070 ;
        RECT 82.900 134.055 83.040 134.210 ;
        RECT 83.360 134.055 83.500 134.550 ;
        RECT 86.030 134.490 86.350 134.550 ;
        RECT 102.145 134.505 102.435 134.735 ;
        RECT 109.045 134.690 109.335 134.735 ;
        RECT 109.490 134.690 109.810 134.750 ;
        RECT 109.045 134.550 109.810 134.690 ;
        RECT 109.045 134.505 109.335 134.550 ;
        RECT 84.650 134.350 84.970 134.410 ;
        RECT 86.505 134.350 86.795 134.395 ;
        RECT 94.720 134.350 95.010 134.395 ;
        RECT 96.150 134.350 96.470 134.410 ;
        RECT 97.980 134.350 98.270 134.395 ;
        RECT 84.650 134.210 91.320 134.350 ;
        RECT 84.650 134.150 84.970 134.210 ;
        RECT 86.505 134.165 86.795 134.210 ;
        RECT 82.825 133.825 83.115 134.055 ;
        RECT 83.285 133.825 83.575 134.055 ;
        RECT 83.730 134.010 84.050 134.070 ;
        RECT 84.205 134.010 84.495 134.055 ;
        RECT 83.730 133.870 84.495 134.010 ;
        RECT 83.730 133.810 84.050 133.870 ;
        RECT 84.205 133.825 84.495 133.870 ;
        RECT 90.170 133.810 90.490 134.070 ;
        RECT 90.645 133.825 90.935 134.055 ;
        RECT 84.650 133.670 84.970 133.730 ;
        RECT 81.520 133.530 84.970 133.670 ;
        RECT 84.650 133.470 84.970 133.530 ;
        RECT 85.110 133.470 85.430 133.730 ;
        RECT 90.720 133.670 90.860 133.825 ;
        RECT 88.420 133.530 90.860 133.670 ;
        RECT 91.180 133.670 91.320 134.210 ;
        RECT 94.720 134.210 98.270 134.350 ;
        RECT 94.720 134.165 95.010 134.210 ;
        RECT 96.150 134.150 96.470 134.210 ;
        RECT 97.980 134.165 98.270 134.210 ;
        RECT 98.900 134.350 99.190 134.395 ;
        RECT 100.760 134.350 101.050 134.395 ;
        RECT 98.900 134.210 101.050 134.350 ;
        RECT 98.900 134.165 99.190 134.210 ;
        RECT 100.760 134.165 101.050 134.210 ;
        RECT 96.580 134.010 96.870 134.055 ;
        RECT 98.900 134.010 99.115 134.165 ;
        RECT 96.580 133.870 99.115 134.010 ;
        RECT 99.845 134.010 100.135 134.055 ;
        RECT 102.220 134.010 102.360 134.505 ;
        RECT 109.490 134.490 109.810 134.550 ;
        RECT 112.250 134.490 112.570 134.750 ;
        RECT 121.925 134.690 122.215 134.735 ;
        RECT 123.290 134.690 123.610 134.750 ;
        RECT 121.925 134.550 123.610 134.690 ;
        RECT 121.925 134.505 122.215 134.550 ;
        RECT 123.290 134.490 123.610 134.550 ;
        RECT 135.660 134.480 136.800 134.510 ;
        RECT 99.845 133.870 102.360 134.010 ;
        RECT 96.580 133.825 96.870 133.870 ;
        RECT 99.845 133.825 100.135 133.870 ;
        RECT 103.050 133.810 103.370 134.070 ;
        RECT 103.970 134.010 104.290 134.070 ;
        RECT 109.505 134.010 109.795 134.055 ;
        RECT 103.970 133.870 109.795 134.010 ;
        RECT 103.970 133.810 104.290 133.870 ;
        RECT 109.505 133.825 109.795 133.870 ;
        RECT 111.330 133.810 111.650 134.070 ;
        RECT 115.930 134.010 116.250 134.070 ;
        RECT 121.005 134.010 121.295 134.055 ;
        RECT 115.930 133.870 121.295 134.010 ;
        RECT 115.930 133.810 116.250 133.870 ;
        RECT 121.005 133.825 121.295 133.870 ;
        RECT 92.715 133.670 93.005 133.715 ;
        RECT 97.990 133.670 98.310 133.730 ;
        RECT 91.180 133.530 98.310 133.670 ;
        RECT 19.805 133.145 20.095 133.375 ;
        RECT 28.040 133.330 28.330 133.375 ;
        RECT 30.820 133.330 31.110 133.375 ;
        RECT 32.680 133.330 32.970 133.375 ;
        RECT 28.040 133.190 32.970 133.330 ;
        RECT 28.040 133.145 28.330 133.190 ;
        RECT 30.820 133.145 31.110 133.190 ;
        RECT 32.680 133.145 32.970 133.190 ;
        RECT 36.350 133.330 36.670 133.390 ;
        RECT 43.680 133.330 43.970 133.375 ;
        RECT 46.460 133.330 46.750 133.375 ;
        RECT 48.320 133.330 48.610 133.375 ;
        RECT 36.350 133.190 43.020 133.330 ;
        RECT 36.350 133.130 36.670 133.190 ;
        RECT 39.815 132.990 40.105 133.035 ;
        RECT 41.410 132.990 41.730 133.050 ;
        RECT 42.330 132.990 42.650 133.050 ;
        RECT 39.815 132.850 42.650 132.990 ;
        RECT 42.880 132.990 43.020 133.190 ;
        RECT 43.680 133.190 48.610 133.330 ;
        RECT 43.680 133.145 43.970 133.190 ;
        RECT 46.460 133.145 46.750 133.190 ;
        RECT 48.320 133.145 48.610 133.190 ;
        RECT 73.610 133.130 73.930 133.390 ;
        RECT 88.420 133.375 88.560 133.530 ;
        RECT 92.715 133.485 93.005 133.530 ;
        RECT 97.990 133.470 98.310 133.530 ;
        RECT 101.685 133.670 101.975 133.715 ;
        RECT 111.790 133.670 112.110 133.730 ;
        RECT 101.685 133.530 112.110 133.670 ;
        RECT 101.685 133.485 101.975 133.530 ;
        RECT 111.790 133.470 112.110 133.530 ;
        RECT 135.590 133.400 136.850 134.480 ;
        RECT 80.985 133.330 81.275 133.375 ;
        RECT 80.140 133.190 81.275 133.330 ;
        RECT 80.140 133.050 80.280 133.190 ;
        RECT 80.985 133.145 81.275 133.190 ;
        RECT 88.345 133.145 88.635 133.375 ;
        RECT 96.580 133.330 96.870 133.375 ;
        RECT 99.360 133.330 99.650 133.375 ;
        RECT 101.220 133.330 101.510 133.375 ;
        RECT 96.580 133.190 101.510 133.330 ;
        RECT 96.580 133.145 96.870 133.190 ;
        RECT 99.360 133.145 99.650 133.190 ;
        RECT 101.220 133.145 101.510 133.190 ;
        RECT 66.725 132.990 67.015 133.035 ;
        RECT 69.930 132.990 70.250 133.050 ;
        RECT 42.880 132.850 70.250 132.990 ;
        RECT 39.815 132.805 40.105 132.850 ;
        RECT 41.410 132.790 41.730 132.850 ;
        RECT 42.330 132.790 42.650 132.850 ;
        RECT 66.725 132.805 67.015 132.850 ;
        RECT 69.930 132.790 70.250 132.850 ;
        RECT 71.785 132.990 72.075 133.035 ;
        RECT 77.290 132.990 77.610 133.050 ;
        RECT 71.785 132.850 77.610 132.990 ;
        RECT 71.785 132.805 72.075 132.850 ;
        RECT 77.290 132.790 77.610 132.850 ;
        RECT 80.050 132.790 80.370 133.050 ;
        RECT 80.510 132.790 80.830 133.050 ;
        RECT 89.710 132.790 90.030 133.050 ;
        RECT 91.090 132.990 91.410 133.050 ;
        RECT 91.565 132.990 91.855 133.035 ;
        RECT 91.090 132.850 91.855 132.990 ;
        RECT 91.090 132.790 91.410 132.850 ;
        RECT 91.565 132.805 91.855 132.850 ;
        RECT 14.660 132.170 127.820 132.650 ;
        RECT 30.830 131.770 31.150 132.030 ;
        RECT 38.190 131.970 38.510 132.030 ;
        RECT 38.665 131.970 38.955 132.015 ;
        RECT 38.190 131.830 38.955 131.970 ;
        RECT 38.190 131.770 38.510 131.830 ;
        RECT 38.665 131.785 38.955 131.830 ;
        RECT 43.250 131.770 43.570 132.030 ;
        RECT 46.485 131.970 46.775 132.015 ;
        RECT 46.930 131.970 47.250 132.030 ;
        RECT 46.485 131.830 47.250 131.970 ;
        RECT 46.485 131.785 46.775 131.830 ;
        RECT 46.930 131.770 47.250 131.830 ;
        RECT 66.495 131.970 66.785 132.015 ;
        RECT 69.470 131.970 69.790 132.030 ;
        RECT 66.495 131.830 69.790 131.970 ;
        RECT 66.495 131.785 66.785 131.830 ;
        RECT 69.470 131.770 69.790 131.830 ;
        RECT 69.930 131.970 70.250 132.030 ;
        RECT 69.930 131.830 79.360 131.970 ;
        RECT 69.930 131.770 70.250 131.830 ;
        RECT 70.360 131.630 70.650 131.675 ;
        RECT 73.140 131.630 73.430 131.675 ;
        RECT 75.000 131.630 75.290 131.675 ;
        RECT 70.360 131.490 75.290 131.630 ;
        RECT 79.220 131.630 79.360 131.830 ;
        RECT 79.590 131.770 79.910 132.030 ;
        RECT 85.355 131.970 85.645 132.015 ;
        RECT 86.030 131.970 86.350 132.030 ;
        RECT 85.355 131.830 86.350 131.970 ;
        RECT 85.355 131.785 85.645 131.830 ;
        RECT 86.030 131.770 86.350 131.830 ;
        RECT 88.880 131.830 95.920 131.970 ;
        RECT 88.880 131.630 89.020 131.830 ;
        RECT 79.220 131.490 89.020 131.630 ;
        RECT 89.220 131.630 89.510 131.675 ;
        RECT 92.000 131.630 92.290 131.675 ;
        RECT 93.860 131.630 94.150 131.675 ;
        RECT 89.220 131.490 94.150 131.630 ;
        RECT 70.360 131.445 70.650 131.490 ;
        RECT 73.140 131.445 73.430 131.490 ;
        RECT 75.000 131.445 75.290 131.490 ;
        RECT 89.220 131.445 89.510 131.490 ;
        RECT 92.000 131.445 92.290 131.490 ;
        RECT 93.860 131.445 94.150 131.490 ;
        RECT 35.905 131.290 36.195 131.335 ;
        RECT 37.270 131.290 37.590 131.350 ;
        RECT 35.905 131.150 37.590 131.290 ;
        RECT 35.905 131.105 36.195 131.150 ;
        RECT 37.270 131.090 37.590 131.150 ;
        RECT 57.510 131.090 57.830 131.350 ;
        RECT 75.450 131.090 75.770 131.350 ;
        RECT 80.525 131.290 80.815 131.335 ;
        RECT 81.430 131.290 81.750 131.350 ;
        RECT 80.525 131.150 81.750 131.290 ;
        RECT 80.525 131.105 80.815 131.150 ;
        RECT 81.430 131.090 81.750 131.150 ;
        RECT 91.090 131.290 91.410 131.350 ;
        RECT 92.485 131.290 92.775 131.335 ;
        RECT 91.090 131.150 92.775 131.290 ;
        RECT 91.090 131.090 91.410 131.150 ;
        RECT 92.485 131.105 92.775 131.150 ;
        RECT 94.325 131.290 94.615 131.335 ;
        RECT 95.230 131.290 95.550 131.350 ;
        RECT 94.325 131.150 95.550 131.290 ;
        RECT 95.780 131.290 95.920 131.830 ;
        RECT 96.150 131.770 96.470 132.030 ;
        RECT 97.530 131.770 97.850 132.030 ;
        RECT 105.350 131.770 105.670 132.030 ;
        RECT 104.890 131.630 105.210 131.690 ;
        RECT 107.665 131.630 107.955 131.675 ;
        RECT 104.890 131.490 107.955 131.630 ;
        RECT 104.890 131.430 105.210 131.490 ;
        RECT 107.665 131.445 107.955 131.490 ;
        RECT 95.780 131.150 104.660 131.290 ;
        RECT 94.325 131.105 94.615 131.150 ;
        RECT 95.230 131.090 95.550 131.150 ;
        RECT 31.290 130.950 31.610 131.010 ;
        RECT 31.765 130.950 32.055 130.995 ;
        RECT 31.290 130.810 32.055 130.950 ;
        RECT 31.290 130.750 31.610 130.810 ;
        RECT 31.765 130.765 32.055 130.810 ;
        RECT 36.810 130.750 37.130 131.010 ;
        RECT 37.730 130.950 38.050 131.010 ;
        RECT 39.110 130.950 39.430 131.010 ;
        RECT 42.805 130.950 43.095 130.995 ;
        RECT 37.730 130.810 43.095 130.950 ;
        RECT 37.730 130.750 38.050 130.810 ;
        RECT 39.110 130.750 39.430 130.810 ;
        RECT 42.805 130.765 43.095 130.810 ;
        RECT 45.550 130.750 45.870 131.010 ;
        RECT 55.670 130.750 55.990 131.010 ;
        RECT 58.890 130.750 59.210 131.010 ;
        RECT 70.360 130.950 70.650 130.995 ;
        RECT 73.625 130.950 73.915 130.995 ;
        RECT 70.360 130.810 72.895 130.950 ;
        RECT 70.360 130.765 70.650 130.810 ;
        RECT 29.910 130.610 30.230 130.670 ;
        RECT 68.550 130.655 68.870 130.670 ;
        RECT 72.680 130.655 72.895 130.810 ;
        RECT 73.625 130.810 76.600 130.950 ;
        RECT 73.625 130.765 73.915 130.810 ;
        RECT 36.365 130.610 36.655 130.655 ;
        RECT 29.910 130.470 36.655 130.610 ;
        RECT 29.910 130.410 30.230 130.470 ;
        RECT 36.365 130.425 36.655 130.470 ;
        RECT 68.500 130.610 68.870 130.655 ;
        RECT 71.760 130.610 72.050 130.655 ;
        RECT 68.500 130.470 72.050 130.610 ;
        RECT 68.500 130.425 68.870 130.470 ;
        RECT 71.760 130.425 72.050 130.470 ;
        RECT 72.680 130.610 72.970 130.655 ;
        RECT 74.540 130.610 74.830 130.655 ;
        RECT 72.680 130.470 74.830 130.610 ;
        RECT 72.680 130.425 72.970 130.470 ;
        RECT 74.540 130.425 74.830 130.470 ;
        RECT 68.550 130.410 68.870 130.425 ;
        RECT 56.130 130.070 56.450 130.330 ;
        RECT 56.590 130.270 56.910 130.330 ;
        RECT 58.445 130.270 58.735 130.315 ;
        RECT 56.590 130.130 58.735 130.270 ;
        RECT 56.590 130.070 56.910 130.130 ;
        RECT 58.445 130.085 58.735 130.130 ;
        RECT 60.745 130.270 61.035 130.315 ;
        RECT 64.410 130.270 64.730 130.330 ;
        RECT 76.460 130.315 76.600 130.810 ;
        RECT 77.290 130.750 77.610 131.010 ;
        RECT 79.605 130.950 79.895 130.995 ;
        RECT 80.050 130.950 80.370 131.010 ;
        RECT 79.605 130.810 80.370 130.950 ;
        RECT 79.605 130.765 79.895 130.810 ;
        RECT 80.050 130.750 80.370 130.810 ;
        RECT 80.970 130.750 81.290 131.010 ;
        RECT 98.540 130.995 98.680 131.150 ;
        RECT 89.220 130.950 89.510 130.995 ;
        RECT 89.220 130.810 91.755 130.950 ;
        RECT 89.220 130.765 89.510 130.810 ;
        RECT 87.360 130.610 87.650 130.655 ;
        RECT 89.710 130.610 90.030 130.670 ;
        RECT 91.540 130.655 91.755 130.810 ;
        RECT 95.705 130.765 95.995 130.995 ;
        RECT 98.465 130.765 98.755 130.995 ;
        RECT 90.620 130.610 90.910 130.655 ;
        RECT 87.360 130.470 90.910 130.610 ;
        RECT 87.360 130.425 87.650 130.470 ;
        RECT 89.710 130.410 90.030 130.470 ;
        RECT 90.620 130.425 90.910 130.470 ;
        RECT 91.540 130.610 91.830 130.655 ;
        RECT 93.400 130.610 93.690 130.655 ;
        RECT 91.540 130.470 93.690 130.610 ;
        RECT 91.540 130.425 91.830 130.470 ;
        RECT 93.400 130.425 93.690 130.470 ;
        RECT 60.745 130.130 64.730 130.270 ;
        RECT 60.745 130.085 61.035 130.130 ;
        RECT 64.410 130.070 64.730 130.130 ;
        RECT 76.385 130.085 76.675 130.315 ;
        RECT 81.905 130.270 82.195 130.315 ;
        RECT 82.350 130.270 82.670 130.330 ;
        RECT 81.905 130.130 82.670 130.270 ;
        RECT 81.905 130.085 82.195 130.130 ;
        RECT 82.350 130.070 82.670 130.130 ;
        RECT 90.170 130.270 90.490 130.330 ;
        RECT 95.780 130.270 95.920 130.765 ;
        RECT 99.370 130.750 99.690 131.010 ;
        RECT 104.520 130.995 104.660 131.150 ;
        RECT 103.985 130.765 104.275 130.995 ;
        RECT 104.445 130.950 104.735 130.995 ;
        RECT 106.270 130.950 106.590 131.010 ;
        RECT 108.585 130.950 108.875 130.995 ;
        RECT 104.445 130.810 108.875 130.950 ;
        RECT 104.445 130.765 104.735 130.810 ;
        RECT 104.060 130.610 104.200 130.765 ;
        RECT 106.270 130.750 106.590 130.810 ;
        RECT 108.585 130.765 108.875 130.810 ;
        RECT 109.030 130.750 109.350 131.010 ;
        RECT 104.890 130.610 105.210 130.670 ;
        RECT 104.060 130.470 105.210 130.610 ;
        RECT 104.890 130.410 105.210 130.470 ;
        RECT 103.970 130.270 104.290 130.330 ;
        RECT 90.170 130.130 104.290 130.270 ;
        RECT 90.170 130.070 90.490 130.130 ;
        RECT 103.970 130.070 104.290 130.130 ;
        RECT 14.660 129.450 127.820 129.930 ;
        RECT 53.615 129.250 53.905 129.295 ;
        RECT 56.590 129.250 56.910 129.310 ;
        RECT 52.080 129.110 56.910 129.250 ;
        RECT 18.360 128.910 18.650 128.955 ;
        RECT 18.870 128.910 19.190 128.970 ;
        RECT 21.620 128.910 21.910 128.955 ;
        RECT 18.360 128.770 21.910 128.910 ;
        RECT 18.360 128.725 18.650 128.770 ;
        RECT 18.870 128.710 19.190 128.770 ;
        RECT 21.620 128.725 21.910 128.770 ;
        RECT 22.540 128.910 22.830 128.955 ;
        RECT 24.400 128.910 24.690 128.955 ;
        RECT 22.540 128.770 24.690 128.910 ;
        RECT 22.540 128.725 22.830 128.770 ;
        RECT 24.400 128.725 24.690 128.770 ;
        RECT 37.270 128.910 37.590 128.970 ;
        RECT 44.185 128.910 44.475 128.955 ;
        RECT 37.270 128.770 44.475 128.910 ;
        RECT 20.220 128.570 20.510 128.615 ;
        RECT 22.540 128.570 22.755 128.725 ;
        RECT 37.270 128.710 37.590 128.770 ;
        RECT 44.185 128.725 44.475 128.770 ;
        RECT 46.945 128.910 47.235 128.955 ;
        RECT 49.705 128.910 49.995 128.955 ;
        RECT 46.945 128.770 49.995 128.910 ;
        RECT 46.945 128.725 47.235 128.770 ;
        RECT 49.705 128.725 49.995 128.770 ;
        RECT 20.220 128.430 22.755 128.570 ;
        RECT 23.010 128.570 23.330 128.630 ;
        RECT 23.485 128.570 23.775 128.615 ;
        RECT 23.010 128.430 23.775 128.570 ;
        RECT 20.220 128.385 20.510 128.430 ;
        RECT 23.010 128.370 23.330 128.430 ;
        RECT 23.485 128.385 23.775 128.430 ;
        RECT 25.310 128.370 25.630 128.630 ;
        RECT 46.025 128.385 46.315 128.615 ;
        RECT 48.325 128.570 48.615 128.615 ;
        RECT 49.230 128.570 49.550 128.630 ;
        RECT 48.325 128.430 49.550 128.570 ;
        RECT 48.325 128.385 48.615 128.430 ;
        RECT 20.220 127.890 20.510 127.935 ;
        RECT 23.000 127.890 23.290 127.935 ;
        RECT 24.860 127.890 25.150 127.935 ;
        RECT 20.220 127.750 25.150 127.890 ;
        RECT 46.100 127.890 46.240 128.385 ;
        RECT 49.230 128.370 49.550 128.430 ;
        RECT 51.085 128.385 51.375 128.615 ;
        RECT 47.865 128.230 48.155 128.275 ;
        RECT 49.690 128.230 50.010 128.290 ;
        RECT 47.865 128.090 50.010 128.230 ;
        RECT 51.160 128.230 51.300 128.385 ;
        RECT 51.530 128.370 51.850 128.630 ;
        RECT 52.080 128.615 52.220 129.110 ;
        RECT 53.615 129.065 53.905 129.110 ;
        RECT 56.590 129.050 56.910 129.110 ;
        RECT 68.550 129.050 68.870 129.310 ;
        RECT 72.690 129.250 73.010 129.310 ;
        RECT 69.100 129.110 73.010 129.250 ;
        RECT 55.620 128.910 55.910 128.955 ;
        RECT 56.130 128.910 56.450 128.970 ;
        RECT 58.880 128.910 59.170 128.955 ;
        RECT 55.620 128.770 59.170 128.910 ;
        RECT 55.620 128.725 55.910 128.770 ;
        RECT 56.130 128.710 56.450 128.770 ;
        RECT 58.880 128.725 59.170 128.770 ;
        RECT 59.800 128.910 60.090 128.955 ;
        RECT 61.660 128.910 61.950 128.955 ;
        RECT 59.800 128.770 61.950 128.910 ;
        RECT 59.800 128.725 60.090 128.770 ;
        RECT 61.660 128.725 61.950 128.770 ;
        RECT 52.005 128.385 52.295 128.615 ;
        RECT 52.925 128.570 53.215 128.615 ;
        RECT 54.750 128.570 55.070 128.630 ;
        RECT 52.925 128.430 55.070 128.570 ;
        RECT 52.925 128.385 53.215 128.430 ;
        RECT 54.750 128.370 55.070 128.430 ;
        RECT 57.480 128.570 57.770 128.615 ;
        RECT 59.800 128.570 60.015 128.725 ;
        RECT 57.480 128.430 60.015 128.570 ;
        RECT 60.270 128.570 60.590 128.630 ;
        RECT 62.585 128.570 62.875 128.615 ;
        RECT 63.950 128.570 64.270 128.630 ;
        RECT 60.270 128.430 64.270 128.570 ;
        RECT 57.480 128.385 57.770 128.430 ;
        RECT 60.270 128.370 60.590 128.430 ;
        RECT 62.585 128.385 62.875 128.430 ;
        RECT 63.950 128.370 64.270 128.430 ;
        RECT 64.410 128.370 64.730 128.630 ;
        RECT 67.170 128.570 67.490 128.630 ;
        RECT 68.105 128.570 68.395 128.615 ;
        RECT 69.100 128.570 69.240 129.110 ;
        RECT 72.690 129.050 73.010 129.110 ;
        RECT 79.590 129.050 79.910 129.310 ;
        RECT 80.510 129.250 80.830 129.310 ;
        RECT 81.905 129.250 82.195 129.295 ;
        RECT 80.510 129.110 82.195 129.250 ;
        RECT 80.510 129.050 80.830 129.110 ;
        RECT 81.905 129.065 82.195 129.110 ;
        RECT 104.430 129.250 104.750 129.310 ;
        RECT 105.365 129.250 105.655 129.295 ;
        RECT 104.430 129.110 105.655 129.250 ;
        RECT 104.430 129.050 104.750 129.110 ;
        RECT 105.365 129.065 105.655 129.110 ;
        RECT 105.810 129.250 106.130 129.310 ;
        RECT 107.665 129.250 107.955 129.295 ;
        RECT 109.965 129.250 110.255 129.295 ;
        RECT 105.810 129.110 107.955 129.250 ;
        RECT 105.810 129.050 106.130 129.110 ;
        RECT 107.665 129.065 107.955 129.110 ;
        RECT 108.200 129.110 110.255 129.250 ;
        RECT 70.850 128.910 71.170 128.970 ;
        RECT 70.020 128.770 71.170 128.910 ;
        RECT 70.020 128.615 70.160 128.770 ;
        RECT 70.850 128.710 71.170 128.770 ;
        RECT 102.590 128.910 102.910 128.970 ;
        RECT 108.200 128.910 108.340 129.110 ;
        RECT 109.965 129.065 110.255 129.110 ;
        RECT 116.405 128.910 116.695 128.955 ;
        RECT 117.310 128.910 117.630 128.970 ;
        RECT 102.590 128.770 108.340 128.910 ;
        RECT 109.580 128.770 117.630 128.910 ;
        RECT 102.590 128.710 102.910 128.770 ;
        RECT 67.170 128.430 69.240 128.570 ;
        RECT 67.170 128.370 67.490 128.430 ;
        RECT 68.105 128.385 68.395 128.430 ;
        RECT 69.945 128.385 70.235 128.615 ;
        RECT 70.390 128.370 70.710 128.630 ;
        RECT 72.245 128.570 72.535 128.615 ;
        RECT 71.400 128.430 72.535 128.570 ;
        RECT 53.370 128.230 53.690 128.290 ;
        RECT 51.160 128.090 53.690 128.230 ;
        RECT 47.865 128.045 48.155 128.090 ;
        RECT 49.690 128.030 50.010 128.090 ;
        RECT 52.080 127.950 52.220 128.090 ;
        RECT 53.370 128.030 53.690 128.090 ;
        RECT 60.745 128.230 61.035 128.275 ;
        RECT 60.745 128.090 63.720 128.230 ;
        RECT 60.745 128.045 61.035 128.090 ;
        RECT 46.100 127.750 50.840 127.890 ;
        RECT 20.220 127.705 20.510 127.750 ;
        RECT 23.000 127.705 23.290 127.750 ;
        RECT 24.860 127.705 25.150 127.750 ;
        RECT 16.355 127.550 16.645 127.595 ;
        RECT 21.630 127.550 21.950 127.610 ;
        RECT 16.355 127.410 21.950 127.550 ;
        RECT 16.355 127.365 16.645 127.410 ;
        RECT 21.630 127.350 21.950 127.410 ;
        RECT 46.470 127.550 46.790 127.610 ;
        RECT 46.945 127.550 47.235 127.595 ;
        RECT 46.470 127.410 47.235 127.550 ;
        RECT 46.470 127.350 46.790 127.410 ;
        RECT 46.945 127.365 47.235 127.410 ;
        RECT 49.245 127.550 49.535 127.595 ;
        RECT 50.150 127.550 50.470 127.610 ;
        RECT 49.245 127.410 50.470 127.550 ;
        RECT 50.700 127.550 50.840 127.750 ;
        RECT 51.990 127.690 52.310 127.950 ;
        RECT 63.580 127.935 63.720 128.090 ;
        RECT 57.480 127.890 57.770 127.935 ;
        RECT 60.260 127.890 60.550 127.935 ;
        RECT 62.120 127.890 62.410 127.935 ;
        RECT 57.480 127.750 62.410 127.890 ;
        RECT 57.480 127.705 57.770 127.750 ;
        RECT 60.260 127.705 60.550 127.750 ;
        RECT 62.120 127.705 62.410 127.750 ;
        RECT 63.505 127.705 63.795 127.935 ;
        RECT 71.400 127.595 71.540 128.430 ;
        RECT 72.245 128.385 72.535 128.430 ;
        RECT 73.610 128.570 73.930 128.630 ;
        RECT 77.750 128.570 78.070 128.630 ;
        RECT 80.525 128.570 80.815 128.615 ;
        RECT 82.825 128.570 83.115 128.615 ;
        RECT 73.610 128.430 83.115 128.570 ;
        RECT 73.610 128.370 73.930 128.430 ;
        RECT 77.750 128.370 78.070 128.430 ;
        RECT 80.525 128.385 80.815 128.430 ;
        RECT 82.825 128.385 83.115 128.430 ;
        RECT 106.270 128.570 106.590 128.630 ;
        RECT 109.580 128.615 109.720 128.770 ;
        RECT 116.405 128.725 116.695 128.770 ;
        RECT 117.310 128.710 117.630 128.770 ;
        RECT 108.585 128.570 108.875 128.615 ;
        RECT 106.270 128.430 108.875 128.570 ;
        RECT 106.270 128.370 106.590 128.430 ;
        RECT 108.585 128.385 108.875 128.430 ;
        RECT 109.505 128.385 109.795 128.615 ;
        RECT 110.885 128.385 111.175 128.615 ;
        RECT 81.445 128.230 81.735 128.275 ;
        RECT 83.270 128.230 83.590 128.290 ;
        RECT 81.445 128.090 83.590 128.230 ;
        RECT 81.445 128.045 81.735 128.090 ;
        RECT 83.270 128.030 83.590 128.090 ;
        RECT 83.730 128.030 84.050 128.290 ;
        RECT 107.205 128.045 107.495 128.275 ;
        RECT 108.660 128.230 108.800 128.385 ;
        RECT 110.960 128.230 111.100 128.385 ;
        RECT 116.850 128.370 117.170 128.630 ;
        RECT 108.660 128.090 111.100 128.230 ;
        RECT 111.805 128.230 112.095 128.275 ;
        RECT 112.710 128.230 113.030 128.290 ;
        RECT 111.805 128.090 113.030 128.230 ;
        RECT 111.805 128.045 112.095 128.090 ;
        RECT 106.270 127.890 106.590 127.950 ;
        RECT 107.280 127.890 107.420 128.045 ;
        RECT 112.710 128.030 113.030 128.090 ;
        RECT 115.470 128.030 115.790 128.290 ;
        RECT 106.270 127.750 107.420 127.890 ;
        RECT 106.270 127.690 106.590 127.750 ;
        RECT 71.325 127.550 71.615 127.595 ;
        RECT 50.700 127.410 71.615 127.550 ;
        RECT 49.245 127.365 49.535 127.410 ;
        RECT 50.150 127.350 50.470 127.410 ;
        RECT 71.325 127.365 71.615 127.410 ;
        RECT 73.625 127.550 73.915 127.595 ;
        RECT 76.370 127.550 76.690 127.610 ;
        RECT 73.625 127.410 76.690 127.550 ;
        RECT 73.625 127.365 73.915 127.410 ;
        RECT 76.370 127.350 76.690 127.410 ;
        RECT 118.230 127.550 118.550 127.610 ;
        RECT 118.705 127.550 118.995 127.595 ;
        RECT 118.230 127.410 118.995 127.550 ;
        RECT 118.230 127.350 118.550 127.410 ;
        RECT 118.705 127.365 118.995 127.410 ;
        RECT 14.660 126.730 127.820 127.210 ;
        RECT 39.570 126.330 39.890 126.590 ;
        RECT 43.250 126.330 43.570 126.590 ;
        RECT 43.725 126.345 44.015 126.575 ;
        RECT 42.330 126.190 42.650 126.250 ;
        RECT 43.800 126.190 43.940 126.345 ;
        RECT 51.990 126.190 52.310 126.250 ;
        RECT 42.330 126.050 43.940 126.190 ;
        RECT 47.940 126.050 52.310 126.190 ;
        RECT 42.330 125.990 42.650 126.050 ;
        RECT 25.310 125.850 25.630 125.910 ;
        RECT 25.310 125.710 30.140 125.850 ;
        RECT 25.310 125.650 25.630 125.710 ;
        RECT 30.000 125.570 30.140 125.710 ;
        RECT 44.260 125.710 45.780 125.850 ;
        RECT 29.450 125.310 29.770 125.570 ;
        RECT 29.910 125.510 30.230 125.570 ;
        RECT 32.670 125.510 32.990 125.570 ;
        RECT 29.910 125.370 32.990 125.510 ;
        RECT 29.910 125.310 30.230 125.370 ;
        RECT 32.670 125.310 32.990 125.370 ;
        RECT 38.650 125.510 38.970 125.570 ;
        RECT 39.125 125.510 39.415 125.555 ;
        RECT 38.650 125.370 39.415 125.510 ;
        RECT 38.650 125.310 38.970 125.370 ;
        RECT 39.125 125.325 39.415 125.370 ;
        RECT 39.585 125.510 39.875 125.555 ;
        RECT 40.030 125.510 40.350 125.570 ;
        RECT 39.585 125.370 40.350 125.510 ;
        RECT 39.585 125.325 39.875 125.370 ;
        RECT 40.030 125.310 40.350 125.370 ;
        RECT 41.870 125.310 42.190 125.570 ;
        RECT 42.345 125.510 42.635 125.555 ;
        RECT 42.790 125.510 43.110 125.570 ;
        RECT 42.345 125.370 43.110 125.510 ;
        RECT 42.345 125.325 42.635 125.370 ;
        RECT 42.790 125.310 43.110 125.370 ;
        RECT 43.725 125.510 44.015 125.555 ;
        RECT 44.260 125.510 44.400 125.710 ;
        RECT 43.725 125.370 44.400 125.510 ;
        RECT 43.725 125.325 44.015 125.370 ;
        RECT 44.630 125.310 44.950 125.570 ;
        RECT 45.090 125.310 45.410 125.570 ;
        RECT 45.640 125.510 45.780 125.710 ;
        RECT 47.940 125.555 48.080 126.050 ;
        RECT 51.990 125.990 52.310 126.050 ;
        RECT 62.540 126.190 62.830 126.235 ;
        RECT 65.320 126.190 65.610 126.235 ;
        RECT 67.180 126.190 67.470 126.235 ;
        RECT 85.110 126.190 85.430 126.250 ;
        RECT 115.470 126.190 115.790 126.250 ;
        RECT 62.540 126.050 67.470 126.190 ;
        RECT 62.540 126.005 62.830 126.050 ;
        RECT 65.320 126.005 65.610 126.050 ;
        RECT 67.180 126.005 67.470 126.050 ;
        RECT 81.980 126.050 98.220 126.190 ;
        RECT 51.530 125.850 51.850 125.910 ;
        RECT 55.225 125.850 55.515 125.895 ;
        RECT 57.510 125.850 57.830 125.910 ;
        RECT 48.400 125.710 52.680 125.850 ;
        RECT 48.400 125.555 48.540 125.710 ;
        RECT 51.530 125.650 51.850 125.710 ;
        RECT 52.540 125.570 52.680 125.710 ;
        RECT 55.225 125.710 57.830 125.850 ;
        RECT 55.225 125.665 55.515 125.710 ;
        RECT 57.510 125.650 57.830 125.710 ;
        RECT 63.950 125.850 64.270 125.910 ;
        RECT 63.950 125.710 65.560 125.850 ;
        RECT 63.950 125.650 64.270 125.710 ;
        RECT 45.640 125.370 47.160 125.510 ;
        RECT 40.490 124.970 40.810 125.230 ;
        RECT 43.265 125.170 43.555 125.215 ;
        RECT 46.485 125.170 46.775 125.215 ;
        RECT 43.265 125.030 46.775 125.170 ;
        RECT 47.020 125.170 47.160 125.370 ;
        RECT 47.865 125.325 48.155 125.555 ;
        RECT 48.325 125.325 48.615 125.555 ;
        RECT 48.785 125.510 49.075 125.555 ;
        RECT 49.230 125.510 49.550 125.570 ;
        RECT 48.785 125.370 49.550 125.510 ;
        RECT 48.785 125.325 49.075 125.370 ;
        RECT 49.230 125.310 49.550 125.370 ;
        RECT 49.705 125.510 49.995 125.555 ;
        RECT 49.705 125.370 51.760 125.510 ;
        RECT 49.705 125.325 49.995 125.370 ;
        RECT 50.625 125.170 50.915 125.215 ;
        RECT 47.020 125.030 50.915 125.170 ;
        RECT 43.265 124.985 43.555 125.030 ;
        RECT 46.485 124.985 46.775 125.030 ;
        RECT 50.625 124.985 50.915 125.030 ;
        RECT 30.370 124.630 30.690 124.890 ;
        RECT 38.190 124.630 38.510 124.890 ;
        RECT 40.950 124.630 41.270 124.890 ;
        RECT 46.010 124.630 46.330 124.890 ;
        RECT 51.620 124.830 51.760 125.370 ;
        RECT 51.990 125.310 52.310 125.570 ;
        RECT 52.450 125.310 52.770 125.570 ;
        RECT 52.925 125.325 53.215 125.555 ;
        RECT 53.845 125.510 54.135 125.555 ;
        RECT 54.750 125.510 55.070 125.570 ;
        RECT 53.845 125.370 55.070 125.510 ;
        RECT 53.845 125.325 54.135 125.370 ;
        RECT 53.000 125.170 53.140 125.325 ;
        RECT 54.750 125.310 55.070 125.370 ;
        RECT 56.145 125.510 56.435 125.555 ;
        RECT 56.590 125.510 56.910 125.570 ;
        RECT 56.145 125.370 56.910 125.510 ;
        RECT 56.145 125.325 56.435 125.370 ;
        RECT 56.590 125.310 56.910 125.370 ;
        RECT 62.540 125.510 62.830 125.555 ;
        RECT 65.420 125.510 65.560 125.710 ;
        RECT 65.790 125.650 66.110 125.910 ;
        RECT 76.370 125.850 76.690 125.910 ;
        RECT 81.980 125.895 82.120 126.050 ;
        RECT 85.110 125.990 85.430 126.050 ;
        RECT 81.905 125.850 82.195 125.895 ;
        RECT 76.370 125.710 82.195 125.850 ;
        RECT 76.370 125.650 76.690 125.710 ;
        RECT 81.905 125.665 82.195 125.710 ;
        RECT 83.820 125.710 86.260 125.850 ;
        RECT 67.645 125.510 67.935 125.555 ;
        RECT 62.540 125.370 65.075 125.510 ;
        RECT 65.420 125.370 67.935 125.510 ;
        RECT 62.540 125.325 62.830 125.370 ;
        RECT 55.685 125.170 55.975 125.215 ;
        RECT 57.510 125.170 57.830 125.230 ;
        RECT 58.675 125.170 58.965 125.215 ;
        RECT 53.000 125.030 58.965 125.170 ;
        RECT 55.685 124.985 55.975 125.030 ;
        RECT 57.510 124.970 57.830 125.030 ;
        RECT 58.675 124.985 58.965 125.030 ;
        RECT 60.680 125.170 60.970 125.215 ;
        RECT 61.650 125.170 61.970 125.230 ;
        RECT 64.860 125.215 65.075 125.370 ;
        RECT 67.645 125.325 67.935 125.370 ;
        RECT 75.910 125.510 76.230 125.570 ;
        RECT 77.305 125.510 77.595 125.555 ;
        RECT 75.910 125.370 77.595 125.510 ;
        RECT 75.910 125.310 76.230 125.370 ;
        RECT 77.305 125.325 77.595 125.370 ;
        RECT 77.750 125.510 78.070 125.570 ;
        RECT 78.225 125.510 78.515 125.555 ;
        RECT 77.750 125.370 78.515 125.510 ;
        RECT 77.750 125.310 78.070 125.370 ;
        RECT 78.225 125.325 78.515 125.370 ;
        RECT 63.940 125.170 64.230 125.215 ;
        RECT 60.680 125.030 64.230 125.170 ;
        RECT 60.680 124.985 60.970 125.030 ;
        RECT 61.650 124.970 61.970 125.030 ;
        RECT 63.940 124.985 64.230 125.030 ;
        RECT 64.860 125.170 65.150 125.215 ;
        RECT 66.720 125.170 67.010 125.215 ;
        RECT 64.860 125.030 67.010 125.170 ;
        RECT 78.300 125.170 78.440 125.325 ;
        RECT 79.130 125.310 79.450 125.570 ;
        RECT 83.820 125.510 83.960 125.710 ;
        RECT 79.680 125.370 83.960 125.510 ;
        RECT 84.190 125.510 84.510 125.570 ;
        RECT 85.585 125.510 85.875 125.555 ;
        RECT 84.190 125.370 85.875 125.510 ;
        RECT 86.120 125.510 86.260 125.710 ;
        RECT 87.410 125.650 87.730 125.910 ;
        RECT 98.080 125.895 98.220 126.050 ;
        RECT 105.900 126.050 115.790 126.190 ;
        RECT 105.900 125.895 106.040 126.050 ;
        RECT 115.470 125.990 115.790 126.050 ;
        RECT 118.200 126.190 118.490 126.235 ;
        RECT 120.980 126.190 121.270 126.235 ;
        RECT 122.840 126.190 123.130 126.235 ;
        RECT 118.200 126.050 123.130 126.190 ;
        RECT 118.200 126.005 118.490 126.050 ;
        RECT 120.980 126.005 121.270 126.050 ;
        RECT 122.840 126.005 123.130 126.050 ;
        RECT 98.005 125.850 98.295 125.895 ;
        RECT 105.825 125.850 106.115 125.895 ;
        RECT 98.005 125.710 106.115 125.850 ;
        RECT 98.005 125.665 98.295 125.710 ;
        RECT 105.825 125.665 106.115 125.710 ;
        RECT 106.745 125.850 107.035 125.895 ;
        RECT 109.030 125.850 109.350 125.910 ;
        RECT 114.335 125.850 114.625 125.895 ;
        RECT 116.850 125.850 117.170 125.910 ;
        RECT 106.745 125.710 117.170 125.850 ;
        RECT 106.745 125.665 107.035 125.710 ;
        RECT 109.030 125.650 109.350 125.710 ;
        RECT 114.335 125.665 114.625 125.710 ;
        RECT 116.850 125.650 117.170 125.710 ;
        RECT 86.505 125.510 86.795 125.555 ;
        RECT 86.120 125.370 86.795 125.510 ;
        RECT 79.680 125.170 79.820 125.370 ;
        RECT 84.190 125.310 84.510 125.370 ;
        RECT 85.585 125.325 85.875 125.370 ;
        RECT 86.505 125.325 86.795 125.370 ;
        RECT 103.970 125.510 104.290 125.570 ;
        RECT 112.725 125.510 113.015 125.555 ;
        RECT 113.630 125.510 113.950 125.570 ;
        RECT 103.970 125.370 113.950 125.510 ;
        RECT 103.970 125.310 104.290 125.370 ;
        RECT 112.725 125.325 113.015 125.370 ;
        RECT 113.630 125.310 113.950 125.370 ;
        RECT 118.200 125.510 118.490 125.555 ;
        RECT 118.200 125.370 120.735 125.510 ;
        RECT 118.200 125.325 118.490 125.370 ;
        RECT 78.300 125.030 79.820 125.170 ;
        RECT 82.825 125.170 83.115 125.215 ;
        RECT 83.730 125.170 84.050 125.230 ;
        RECT 88.790 125.170 89.110 125.230 ;
        RECT 120.520 125.215 120.735 125.370 ;
        RECT 121.450 125.310 121.770 125.570 ;
        RECT 123.305 125.510 123.595 125.555 ;
        RECT 125.590 125.510 125.910 125.570 ;
        RECT 123.305 125.370 125.910 125.510 ;
        RECT 123.305 125.325 123.595 125.370 ;
        RECT 125.590 125.310 125.910 125.370 ;
        RECT 82.825 125.030 89.110 125.170 ;
        RECT 64.860 124.985 65.150 125.030 ;
        RECT 66.720 124.985 67.010 125.030 ;
        RECT 82.825 124.985 83.115 125.030 ;
        RECT 83.730 124.970 84.050 125.030 ;
        RECT 88.790 124.970 89.110 125.030 ;
        RECT 98.925 125.170 99.215 125.215 ;
        RECT 113.185 125.170 113.475 125.215 ;
        RECT 116.340 125.170 116.630 125.215 ;
        RECT 119.600 125.170 119.890 125.215 ;
        RECT 98.925 125.030 105.120 125.170 ;
        RECT 98.925 124.985 99.215 125.030 ;
        RECT 104.980 124.890 105.120 125.030 ;
        RECT 113.185 125.030 119.890 125.170 ;
        RECT 113.185 124.985 113.475 125.030 ;
        RECT 116.340 124.985 116.630 125.030 ;
        RECT 119.600 124.985 119.890 125.030 ;
        RECT 120.520 125.170 120.810 125.215 ;
        RECT 122.380 125.170 122.670 125.215 ;
        RECT 120.520 125.030 122.670 125.170 ;
        RECT 120.520 124.985 120.810 125.030 ;
        RECT 122.380 124.985 122.670 125.030 ;
        RECT 54.750 124.830 55.070 124.890 ;
        RECT 51.620 124.690 55.070 124.830 ;
        RECT 54.750 124.630 55.070 124.690 ;
        RECT 57.985 124.830 58.275 124.875 ;
        RECT 62.110 124.830 62.430 124.890 ;
        RECT 57.985 124.690 62.430 124.830 ;
        RECT 57.985 124.645 58.275 124.690 ;
        RECT 62.110 124.630 62.430 124.690 ;
        RECT 83.270 124.630 83.590 124.890 ;
        RECT 85.125 124.830 85.415 124.875 ;
        RECT 86.950 124.830 87.270 124.890 ;
        RECT 85.125 124.690 87.270 124.830 ;
        RECT 85.125 124.645 85.415 124.690 ;
        RECT 86.950 124.630 87.270 124.690 ;
        RECT 93.850 124.830 94.170 124.890 ;
        RECT 99.370 124.830 99.690 124.890 ;
        RECT 93.850 124.690 99.690 124.830 ;
        RECT 93.850 124.630 94.170 124.690 ;
        RECT 99.370 124.630 99.690 124.690 ;
        RECT 101.210 124.630 101.530 124.890 ;
        RECT 104.430 124.630 104.750 124.890 ;
        RECT 104.890 124.830 105.210 124.890 ;
        RECT 107.205 124.830 107.495 124.875 ;
        RECT 104.890 124.690 107.495 124.830 ;
        RECT 104.890 124.630 105.210 124.690 ;
        RECT 107.205 124.645 107.495 124.690 ;
        RECT 109.030 124.630 109.350 124.890 ;
        RECT 14.660 124.010 127.820 124.490 ;
        RECT 23.010 123.610 23.330 123.870 ;
        RECT 39.570 123.610 39.890 123.870 ;
        RECT 40.030 123.810 40.350 123.870 ;
        RECT 41.885 123.810 42.175 123.855 ;
        RECT 42.330 123.810 42.650 123.870 ;
        RECT 40.030 123.670 41.180 123.810 ;
        RECT 40.030 123.610 40.350 123.670 ;
        RECT 19.330 123.470 19.650 123.530 ;
        RECT 25.720 123.470 26.010 123.515 ;
        RECT 28.980 123.470 29.270 123.515 ;
        RECT 19.330 123.330 29.270 123.470 ;
        RECT 19.330 123.270 19.650 123.330 ;
        RECT 25.720 123.285 26.010 123.330 ;
        RECT 28.980 123.285 29.270 123.330 ;
        RECT 29.900 123.470 30.190 123.515 ;
        RECT 31.760 123.470 32.050 123.515 ;
        RECT 41.040 123.470 41.180 123.670 ;
        RECT 41.885 123.670 42.650 123.810 ;
        RECT 41.885 123.625 42.175 123.670 ;
        RECT 42.330 123.610 42.650 123.670 ;
        RECT 43.250 123.810 43.570 123.870 ;
        RECT 44.185 123.810 44.475 123.855 ;
        RECT 43.250 123.670 44.475 123.810 ;
        RECT 43.250 123.610 43.570 123.670 ;
        RECT 44.185 123.625 44.475 123.670 ;
        RECT 46.470 123.610 46.790 123.870 ;
        RECT 61.650 123.610 61.970 123.870 ;
        RECT 64.885 123.810 65.175 123.855 ;
        RECT 65.790 123.810 66.110 123.870 ;
        RECT 64.885 123.670 66.110 123.810 ;
        RECT 64.885 123.625 65.175 123.670 ;
        RECT 65.790 123.610 66.110 123.670 ;
        RECT 102.375 123.810 102.665 123.855 ;
        RECT 104.890 123.810 105.210 123.870 ;
        RECT 102.375 123.670 105.210 123.810 ;
        RECT 102.375 123.625 102.665 123.670 ;
        RECT 104.890 123.610 105.210 123.670 ;
        RECT 116.175 123.810 116.465 123.855 ;
        RECT 117.310 123.810 117.630 123.870 ;
        RECT 116.175 123.670 117.630 123.810 ;
        RECT 116.175 123.625 116.465 123.670 ;
        RECT 117.310 123.610 117.630 123.670 ;
        RECT 55.670 123.470 55.990 123.530 ;
        RECT 90.170 123.470 90.490 123.530 ;
        RECT 97.990 123.515 98.310 123.530 ;
        RECT 104.430 123.515 104.750 123.530 ;
        RECT 94.720 123.470 95.010 123.515 ;
        RECT 97.980 123.470 98.310 123.515 ;
        RECT 29.900 123.330 32.050 123.470 ;
        RECT 29.900 123.285 30.190 123.330 ;
        RECT 31.760 123.285 32.050 123.330 ;
        RECT 35.060 123.330 40.720 123.470 ;
        RECT 22.105 123.130 22.395 123.175 ;
        RECT 24.850 123.130 25.170 123.190 ;
        RECT 22.105 122.990 25.170 123.130 ;
        RECT 22.105 122.945 22.395 122.990 ;
        RECT 24.850 122.930 25.170 122.990 ;
        RECT 27.580 123.130 27.870 123.175 ;
        RECT 29.900 123.130 30.115 123.285 ;
        RECT 35.060 123.190 35.200 123.330 ;
        RECT 27.580 122.990 30.115 123.130 ;
        RECT 30.370 123.130 30.690 123.190 ;
        RECT 30.845 123.130 31.135 123.175 ;
        RECT 30.370 122.990 31.135 123.130 ;
        RECT 27.580 122.945 27.870 122.990 ;
        RECT 30.370 122.930 30.690 122.990 ;
        RECT 30.845 122.945 31.135 122.990 ;
        RECT 32.670 122.930 32.990 123.190 ;
        RECT 34.970 122.930 35.290 123.190 ;
        RECT 35.445 123.130 35.735 123.175 ;
        RECT 37.270 123.130 37.590 123.190 ;
        RECT 38.665 123.130 38.955 123.175 ;
        RECT 39.570 123.130 39.890 123.190 ;
        RECT 40.580 123.175 40.720 123.330 ;
        RECT 41.040 123.330 43.480 123.470 ;
        RECT 41.040 123.175 41.180 123.330 ;
        RECT 35.445 122.990 38.420 123.130 ;
        RECT 35.445 122.945 35.735 122.990 ;
        RECT 37.270 122.930 37.590 122.990 ;
        RECT 28.070 122.790 28.390 122.850 ;
        RECT 36.365 122.790 36.655 122.835 ;
        RECT 36.810 122.790 37.130 122.850 ;
        RECT 28.070 122.650 37.130 122.790 ;
        RECT 28.070 122.590 28.390 122.650 ;
        RECT 36.365 122.605 36.655 122.650 ;
        RECT 36.810 122.590 37.130 122.650 ;
        RECT 37.745 122.605 38.035 122.835 ;
        RECT 38.280 122.790 38.420 122.990 ;
        RECT 38.665 122.990 39.890 123.130 ;
        RECT 38.665 122.945 38.955 122.990 ;
        RECT 39.570 122.930 39.890 122.990 ;
        RECT 40.505 122.945 40.795 123.175 ;
        RECT 40.965 122.945 41.255 123.175 ;
        RECT 41.870 123.130 42.190 123.190 ;
        RECT 43.340 123.175 43.480 123.330 ;
        RECT 55.670 123.330 61.420 123.470 ;
        RECT 55.670 123.270 55.990 123.330 ;
        RECT 42.345 123.130 42.635 123.175 ;
        RECT 41.870 122.990 42.635 123.130 ;
        RECT 41.870 122.930 42.190 122.990 ;
        RECT 42.345 122.945 42.635 122.990 ;
        RECT 43.265 123.130 43.555 123.175 ;
        RECT 45.550 123.130 45.870 123.190 ;
        RECT 43.265 122.990 45.870 123.130 ;
        RECT 43.265 122.945 43.555 122.990 ;
        RECT 45.550 122.930 45.870 122.990 ;
        RECT 56.130 122.930 56.450 123.190 ;
        RECT 61.280 123.175 61.420 123.330 ;
        RECT 74.160 123.330 91.320 123.470 ;
        RECT 74.160 123.190 74.300 123.330 ;
        RECT 90.170 123.270 90.490 123.330 ;
        RECT 61.205 122.945 61.495 123.175 ;
        RECT 62.110 123.130 62.430 123.190 ;
        RECT 63.965 123.130 64.255 123.175 ;
        RECT 62.110 122.990 64.255 123.130 ;
        RECT 62.110 122.930 62.430 122.990 ;
        RECT 63.965 122.945 64.255 122.990 ;
        RECT 74.070 122.930 74.390 123.190 ;
        RECT 75.910 123.130 76.230 123.190 ;
        RECT 77.305 123.130 77.595 123.175 ;
        RECT 75.910 122.990 77.595 123.130 ;
        RECT 75.910 122.930 76.230 122.990 ;
        RECT 77.305 122.945 77.595 122.990 ;
        RECT 88.330 122.930 88.650 123.190 ;
        RECT 91.180 123.175 91.320 123.330 ;
        RECT 94.720 123.330 98.310 123.470 ;
        RECT 94.720 123.285 95.010 123.330 ;
        RECT 97.980 123.285 98.310 123.330 ;
        RECT 97.990 123.270 98.310 123.285 ;
        RECT 98.900 123.470 99.190 123.515 ;
        RECT 100.760 123.470 101.050 123.515 ;
        RECT 98.900 123.330 101.050 123.470 ;
        RECT 98.900 123.285 99.190 123.330 ;
        RECT 100.760 123.285 101.050 123.330 ;
        RECT 104.380 123.470 104.750 123.515 ;
        RECT 107.640 123.470 107.930 123.515 ;
        RECT 104.380 123.330 107.930 123.470 ;
        RECT 104.380 123.285 104.750 123.330 ;
        RECT 107.640 123.285 107.930 123.330 ;
        RECT 108.560 123.470 108.850 123.515 ;
        RECT 110.420 123.470 110.710 123.515 ;
        RECT 108.560 123.330 110.710 123.470 ;
        RECT 108.560 123.285 108.850 123.330 ;
        RECT 110.420 123.285 110.710 123.330 ;
        RECT 113.645 123.470 113.935 123.515 ;
        RECT 118.180 123.470 118.470 123.515 ;
        RECT 121.440 123.470 121.730 123.515 ;
        RECT 113.645 123.330 121.730 123.470 ;
        RECT 113.645 123.285 113.935 123.330 ;
        RECT 118.180 123.285 118.470 123.330 ;
        RECT 121.440 123.285 121.730 123.330 ;
        RECT 122.360 123.470 122.650 123.515 ;
        RECT 124.220 123.470 124.510 123.515 ;
        RECT 122.360 123.330 124.510 123.470 ;
        RECT 122.360 123.285 122.650 123.330 ;
        RECT 124.220 123.285 124.510 123.330 ;
        RECT 91.105 122.945 91.395 123.175 ;
        RECT 96.580 123.130 96.870 123.175 ;
        RECT 98.900 123.130 99.115 123.285 ;
        RECT 104.430 123.270 104.750 123.285 ;
        RECT 96.580 122.990 99.115 123.130 ;
        RECT 96.580 122.945 96.870 122.990 ;
        RECT 99.830 122.930 100.150 123.190 ;
        RECT 106.240 123.130 106.530 123.175 ;
        RECT 108.560 123.130 108.775 123.285 ;
        RECT 106.240 122.990 108.775 123.130 ;
        RECT 113.185 123.130 113.475 123.175 ;
        RECT 120.040 123.130 120.330 123.175 ;
        RECT 122.360 123.130 122.575 123.285 ;
        RECT 113.185 122.990 113.860 123.130 ;
        RECT 106.240 122.945 106.530 122.990 ;
        RECT 113.185 122.945 113.475 122.990 ;
        RECT 113.720 122.850 113.860 122.990 ;
        RECT 120.040 122.990 122.575 123.130 ;
        RECT 123.305 123.130 123.595 123.175 ;
        RECT 124.670 123.130 124.990 123.190 ;
        RECT 123.305 122.990 124.990 123.130 ;
        RECT 120.040 122.945 120.330 122.990 ;
        RECT 123.305 122.945 123.595 122.990 ;
        RECT 124.670 122.930 124.990 122.990 ;
        RECT 125.145 123.130 125.435 123.175 ;
        RECT 125.590 123.130 125.910 123.190 ;
        RECT 125.145 122.990 125.910 123.130 ;
        RECT 125.145 122.945 125.435 122.990 ;
        RECT 44.645 122.790 44.935 122.835 ;
        RECT 38.280 122.650 44.935 122.790 ;
        RECT 44.645 122.605 44.935 122.650 ;
        RECT 27.580 122.450 27.870 122.495 ;
        RECT 30.360 122.450 30.650 122.495 ;
        RECT 32.220 122.450 32.510 122.495 ;
        RECT 37.820 122.450 37.960 122.605 ;
        RECT 76.370 122.590 76.690 122.850 ;
        RECT 76.845 122.790 77.135 122.835 ;
        RECT 78.210 122.790 78.530 122.850 ;
        RECT 83.270 122.790 83.590 122.850 ;
        RECT 76.845 122.650 83.590 122.790 ;
        RECT 76.845 122.605 77.135 122.650 ;
        RECT 78.210 122.590 78.530 122.650 ;
        RECT 83.270 122.590 83.590 122.650 ;
        RECT 95.230 122.790 95.550 122.850 ;
        RECT 101.685 122.790 101.975 122.835 ;
        RECT 95.230 122.650 101.975 122.790 ;
        RECT 95.230 122.590 95.550 122.650 ;
        RECT 101.685 122.605 101.975 122.650 ;
        RECT 109.505 122.790 109.795 122.835 ;
        RECT 109.950 122.790 110.270 122.850 ;
        RECT 109.505 122.650 110.270 122.790 ;
        RECT 109.505 122.605 109.795 122.650 ;
        RECT 109.950 122.590 110.270 122.650 ;
        RECT 111.345 122.790 111.635 122.835 ;
        RECT 111.790 122.790 112.110 122.850 ;
        RECT 111.345 122.650 112.110 122.790 ;
        RECT 111.345 122.605 111.635 122.650 ;
        RECT 111.790 122.590 112.110 122.650 ;
        RECT 113.630 122.590 113.950 122.850 ;
        RECT 119.150 122.790 119.470 122.850 ;
        RECT 125.220 122.790 125.360 122.945 ;
        RECT 125.590 122.930 125.910 122.990 ;
        RECT 119.150 122.650 125.360 122.790 ;
        RECT 119.150 122.590 119.470 122.650 ;
        RECT 27.580 122.310 32.510 122.450 ;
        RECT 27.580 122.265 27.870 122.310 ;
        RECT 30.360 122.265 30.650 122.310 ;
        RECT 32.220 122.265 32.510 122.310 ;
        RECT 32.760 122.310 37.960 122.450 ;
        RECT 49.690 122.450 50.010 122.510 ;
        RECT 63.950 122.450 64.270 122.510 ;
        RECT 49.690 122.310 64.270 122.450 ;
        RECT 23.715 122.110 24.005 122.155 ;
        RECT 25.310 122.110 25.630 122.170 ;
        RECT 23.715 121.970 25.630 122.110 ;
        RECT 23.715 121.925 24.005 121.970 ;
        RECT 25.310 121.910 25.630 121.970 ;
        RECT 26.690 122.110 27.010 122.170 ;
        RECT 32.760 122.110 32.900 122.310 ;
        RECT 49.690 122.250 50.010 122.310 ;
        RECT 63.950 122.250 64.270 122.310 ;
        RECT 96.580 122.450 96.870 122.495 ;
        RECT 99.360 122.450 99.650 122.495 ;
        RECT 101.220 122.450 101.510 122.495 ;
        RECT 96.580 122.310 101.510 122.450 ;
        RECT 96.580 122.265 96.870 122.310 ;
        RECT 99.360 122.265 99.650 122.310 ;
        RECT 101.220 122.265 101.510 122.310 ;
        RECT 106.240 122.450 106.530 122.495 ;
        RECT 109.020 122.450 109.310 122.495 ;
        RECT 110.880 122.450 111.170 122.495 ;
        RECT 106.240 122.310 111.170 122.450 ;
        RECT 106.240 122.265 106.530 122.310 ;
        RECT 109.020 122.265 109.310 122.310 ;
        RECT 110.880 122.265 111.170 122.310 ;
        RECT 120.040 122.450 120.330 122.495 ;
        RECT 122.820 122.450 123.110 122.495 ;
        RECT 124.680 122.450 124.970 122.495 ;
        RECT 120.040 122.310 124.970 122.450 ;
        RECT 120.040 122.265 120.330 122.310 ;
        RECT 122.820 122.265 123.110 122.310 ;
        RECT 124.680 122.265 124.970 122.310 ;
        RECT 26.690 121.970 32.900 122.110 ;
        RECT 33.145 122.110 33.435 122.155 ;
        RECT 34.050 122.110 34.370 122.170 ;
        RECT 33.145 121.970 34.370 122.110 ;
        RECT 26.690 121.910 27.010 121.970 ;
        RECT 33.145 121.925 33.435 121.970 ;
        RECT 34.050 121.910 34.370 121.970 ;
        RECT 73.150 122.110 73.470 122.170 ;
        RECT 73.625 122.110 73.915 122.155 ;
        RECT 73.150 121.970 73.915 122.110 ;
        RECT 73.150 121.910 73.470 121.970 ;
        RECT 73.625 121.925 73.915 121.970 ;
        RECT 79.130 121.910 79.450 122.170 ;
        RECT 81.890 121.910 82.210 122.170 ;
        RECT 91.090 122.110 91.410 122.170 ;
        RECT 91.565 122.110 91.855 122.155 ;
        RECT 91.090 121.970 91.855 122.110 ;
        RECT 91.090 121.910 91.410 121.970 ;
        RECT 91.565 121.925 91.855 121.970 ;
        RECT 92.715 122.110 93.005 122.155 ;
        RECT 93.850 122.110 94.170 122.170 ;
        RECT 92.715 121.970 94.170 122.110 ;
        RECT 92.715 121.925 93.005 121.970 ;
        RECT 93.850 121.910 94.170 121.970 ;
        RECT 14.660 121.290 127.820 121.770 ;
        RECT 19.330 120.890 19.650 121.150 ;
        RECT 24.850 120.890 25.170 121.150 ;
        RECT 25.310 121.090 25.630 121.150 ;
        RECT 31.290 121.090 31.610 121.150 ;
        RECT 40.490 121.090 40.810 121.150 ;
        RECT 50.625 121.090 50.915 121.135 ;
        RECT 25.310 120.950 38.420 121.090 ;
        RECT 25.310 120.890 25.630 120.950 ;
        RECT 16.585 120.750 16.875 120.795 ;
        RECT 18.870 120.750 19.190 120.810 ;
        RECT 16.585 120.610 19.190 120.750 ;
        RECT 16.585 120.565 16.875 120.610 ;
        RECT 18.870 120.550 19.190 120.610 ;
        RECT 21.185 120.225 21.475 120.455 ;
        RECT 21.630 120.410 21.950 120.470 ;
        RECT 27.165 120.410 27.455 120.455 ;
        RECT 27.700 120.410 27.840 120.950 ;
        RECT 31.290 120.890 31.610 120.950 ;
        RECT 33.100 120.750 33.390 120.795 ;
        RECT 35.880 120.750 36.170 120.795 ;
        RECT 37.740 120.750 38.030 120.795 ;
        RECT 33.100 120.610 38.030 120.750 ;
        RECT 38.280 120.750 38.420 120.950 ;
        RECT 40.490 120.950 50.915 121.090 ;
        RECT 40.490 120.890 40.810 120.950 ;
        RECT 50.625 120.905 50.915 120.950 ;
        RECT 57.970 120.890 58.290 121.150 ;
        RECT 75.235 121.090 75.525 121.135 ;
        RECT 75.910 121.090 76.230 121.150 ;
        RECT 75.235 120.950 76.230 121.090 ;
        RECT 75.235 120.905 75.525 120.950 ;
        RECT 75.910 120.890 76.230 120.950 ;
        RECT 76.615 121.090 76.905 121.135 ;
        RECT 78.210 121.090 78.530 121.150 ;
        RECT 76.615 120.950 78.530 121.090 ;
        RECT 76.615 120.905 76.905 120.950 ;
        RECT 78.210 120.890 78.530 120.950 ;
        RECT 90.170 121.090 90.490 121.150 ;
        RECT 90.170 120.950 97.760 121.090 ;
        RECT 90.170 120.890 90.490 120.950 ;
        RECT 41.870 120.750 42.190 120.810 ;
        RECT 38.280 120.610 42.190 120.750 ;
        RECT 33.100 120.565 33.390 120.610 ;
        RECT 35.880 120.565 36.170 120.610 ;
        RECT 37.740 120.565 38.030 120.610 ;
        RECT 41.870 120.550 42.190 120.610 ;
        RECT 49.230 120.750 49.550 120.810 ;
        RECT 58.060 120.750 58.200 120.890 ;
        RECT 58.430 120.750 58.750 120.810 ;
        RECT 63.490 120.750 63.810 120.810 ;
        RECT 49.230 120.610 55.440 120.750 ;
        RECT 49.230 120.550 49.550 120.610 ;
        RECT 21.630 120.270 23.010 120.410 ;
        RECT 17.045 120.070 17.335 120.115 ;
        RECT 17.505 120.070 17.795 120.115 ;
        RECT 18.885 120.070 19.175 120.115 ;
        RECT 17.045 119.930 20.940 120.070 ;
        RECT 17.045 119.885 17.335 119.930 ;
        RECT 17.505 119.885 17.795 119.930 ;
        RECT 18.885 119.885 19.175 119.930 ;
        RECT 17.965 119.390 18.255 119.435 ;
        RECT 20.250 119.390 20.570 119.450 ;
        RECT 17.965 119.250 20.570 119.390 ;
        RECT 20.800 119.390 20.940 119.930 ;
        RECT 21.260 119.730 21.400 120.225 ;
        RECT 21.630 120.210 21.950 120.270 ;
        RECT 22.870 120.070 23.010 120.270 ;
        RECT 27.165 120.270 27.840 120.410 ;
        RECT 27.165 120.225 27.455 120.270 ;
        RECT 28.070 120.210 28.390 120.470 ;
        RECT 29.910 120.410 30.230 120.470 ;
        RECT 29.910 120.270 36.120 120.410 ;
        RECT 29.910 120.210 30.230 120.270 ;
        RECT 26.690 120.070 27.010 120.130 ;
        RECT 22.870 119.930 27.010 120.070 ;
        RECT 26.690 119.870 27.010 119.930 ;
        RECT 28.160 119.730 28.300 120.210 ;
        RECT 33.100 120.070 33.390 120.115 ;
        RECT 35.980 120.070 36.120 120.270 ;
        RECT 36.350 120.210 36.670 120.470 ;
        RECT 36.810 120.410 37.130 120.470 ;
        RECT 42.345 120.410 42.635 120.455 ;
        RECT 54.750 120.410 55.070 120.470 ;
        RECT 36.810 120.270 42.635 120.410 ;
        RECT 36.810 120.210 37.130 120.270 ;
        RECT 42.345 120.225 42.635 120.270 ;
        RECT 53.920 120.270 55.070 120.410 ;
        RECT 55.300 120.410 55.440 120.610 ;
        RECT 56.680 120.610 63.810 120.750 ;
        RECT 56.680 120.455 56.820 120.610 ;
        RECT 58.430 120.550 58.750 120.610 ;
        RECT 63.490 120.550 63.810 120.610 ;
        RECT 66.730 120.750 67.020 120.795 ;
        RECT 68.590 120.750 68.880 120.795 ;
        RECT 71.370 120.750 71.660 120.795 ;
        RECT 66.730 120.610 71.660 120.750 ;
        RECT 66.730 120.565 67.020 120.610 ;
        RECT 68.590 120.565 68.880 120.610 ;
        RECT 71.370 120.565 71.660 120.610 ;
        RECT 80.480 120.750 80.770 120.795 ;
        RECT 83.260 120.750 83.550 120.795 ;
        RECT 85.120 120.750 85.410 120.795 ;
        RECT 80.480 120.610 85.410 120.750 ;
        RECT 80.480 120.565 80.770 120.610 ;
        RECT 83.260 120.565 83.550 120.610 ;
        RECT 85.120 120.565 85.410 120.610 ;
        RECT 91.980 120.750 92.270 120.795 ;
        RECT 94.760 120.750 95.050 120.795 ;
        RECT 96.620 120.750 96.910 120.795 ;
        RECT 91.980 120.610 96.910 120.750 ;
        RECT 91.980 120.565 92.270 120.610 ;
        RECT 94.760 120.565 95.050 120.610 ;
        RECT 96.620 120.565 96.910 120.610 ;
        RECT 55.300 120.270 56.360 120.410 ;
        RECT 38.205 120.070 38.495 120.115 ;
        RECT 33.100 119.930 35.635 120.070 ;
        RECT 35.980 119.930 38.495 120.070 ;
        RECT 33.100 119.885 33.390 119.930 ;
        RECT 21.260 119.590 28.300 119.730 ;
        RECT 28.530 119.730 28.850 119.790 ;
        RECT 35.420 119.775 35.635 119.930 ;
        RECT 38.205 119.885 38.495 119.930 ;
        RECT 41.410 120.070 41.730 120.130 ;
        RECT 42.805 120.070 43.095 120.115 ;
        RECT 41.410 119.930 43.095 120.070 ;
        RECT 41.410 119.870 41.730 119.930 ;
        RECT 42.805 119.885 43.095 119.930 ;
        RECT 49.690 119.870 50.010 120.130 ;
        RECT 51.990 119.870 52.310 120.130 ;
        RECT 52.450 119.870 52.770 120.130 ;
        RECT 53.920 120.115 54.060 120.270 ;
        RECT 54.750 120.210 55.070 120.270 ;
        RECT 52.925 119.885 53.215 120.115 ;
        RECT 53.845 119.885 54.135 120.115 ;
        RECT 54.305 120.070 54.595 120.115 ;
        RECT 55.670 120.070 55.990 120.130 ;
        RECT 54.305 119.930 55.990 120.070 ;
        RECT 56.220 120.070 56.360 120.270 ;
        RECT 56.605 120.225 56.895 120.455 ;
        RECT 57.065 120.410 57.355 120.455 ;
        RECT 57.970 120.410 58.290 120.470 ;
        RECT 57.065 120.270 58.290 120.410 ;
        RECT 57.065 120.225 57.355 120.270 ;
        RECT 57.140 120.070 57.280 120.225 ;
        RECT 57.970 120.210 58.290 120.270 ;
        RECT 63.950 120.410 64.270 120.470 ;
        RECT 66.265 120.410 66.555 120.455 ;
        RECT 63.950 120.270 66.555 120.410 ;
        RECT 63.950 120.210 64.270 120.270 ;
        RECT 66.265 120.225 66.555 120.270 ;
        RECT 81.890 120.410 82.210 120.470 ;
        RECT 85.585 120.410 85.875 120.455 ;
        RECT 94.310 120.410 94.630 120.470 ;
        RECT 81.890 120.270 94.630 120.410 ;
        RECT 81.890 120.210 82.210 120.270 ;
        RECT 85.585 120.225 85.875 120.270 ;
        RECT 94.310 120.210 94.630 120.270 ;
        RECT 95.245 120.225 95.535 120.455 ;
        RECT 95.690 120.410 96.010 120.470 ;
        RECT 97.070 120.410 97.390 120.470 ;
        RECT 95.690 120.270 97.390 120.410 ;
        RECT 56.220 119.930 57.280 120.070 ;
        RECT 54.305 119.885 54.595 119.930 ;
        RECT 31.240 119.730 31.530 119.775 ;
        RECT 34.500 119.730 34.790 119.775 ;
        RECT 28.530 119.590 34.790 119.730 ;
        RECT 28.530 119.530 28.850 119.590 ;
        RECT 31.240 119.545 31.530 119.590 ;
        RECT 34.500 119.545 34.790 119.590 ;
        RECT 35.420 119.730 35.710 119.775 ;
        RECT 37.280 119.730 37.570 119.775 ;
        RECT 35.420 119.590 37.570 119.730 ;
        RECT 35.420 119.545 35.710 119.590 ;
        RECT 37.280 119.545 37.570 119.590 ;
        RECT 37.730 119.730 38.050 119.790 ;
        RECT 43.265 119.730 43.555 119.775 ;
        RECT 37.730 119.590 43.555 119.730 ;
        RECT 53.000 119.730 53.140 119.885 ;
        RECT 55.670 119.870 55.990 119.930 ;
        RECT 57.510 119.870 57.830 120.130 ;
        RECT 68.090 119.870 68.410 120.130 ;
        RECT 71.370 120.070 71.660 120.115 ;
        RECT 69.125 119.930 71.660 120.070 ;
        RECT 57.050 119.730 57.370 119.790 ;
        RECT 69.125 119.775 69.340 119.930 ;
        RECT 71.370 119.885 71.660 119.930 ;
        RECT 80.480 120.070 80.770 120.115 ;
        RECT 83.745 120.070 84.035 120.115 ;
        RECT 80.480 119.930 83.015 120.070 ;
        RECT 80.480 119.885 80.770 119.930 ;
        RECT 73.150 119.775 73.470 119.790 ;
        RECT 53.000 119.590 57.370 119.730 ;
        RECT 37.730 119.530 38.050 119.590 ;
        RECT 43.265 119.545 43.555 119.590 ;
        RECT 57.050 119.530 57.370 119.590 ;
        RECT 67.190 119.730 67.480 119.775 ;
        RECT 69.050 119.730 69.340 119.775 ;
        RECT 67.190 119.590 69.340 119.730 ;
        RECT 67.190 119.545 67.480 119.590 ;
        RECT 69.050 119.545 69.340 119.590 ;
        RECT 69.970 119.730 70.260 119.775 ;
        RECT 73.150 119.730 73.520 119.775 ;
        RECT 69.970 119.590 73.520 119.730 ;
        RECT 69.970 119.545 70.260 119.590 ;
        RECT 73.150 119.545 73.520 119.590 ;
        RECT 76.370 119.730 76.690 119.790 ;
        RECT 82.800 119.775 83.015 119.930 ;
        RECT 83.745 119.930 86.260 120.070 ;
        RECT 83.745 119.885 84.035 119.930 ;
        RECT 78.620 119.730 78.910 119.775 ;
        RECT 81.880 119.730 82.170 119.775 ;
        RECT 76.370 119.590 82.170 119.730 ;
        RECT 73.150 119.530 73.470 119.545 ;
        RECT 76.370 119.530 76.690 119.590 ;
        RECT 78.620 119.545 78.910 119.590 ;
        RECT 81.880 119.545 82.170 119.590 ;
        RECT 82.800 119.730 83.090 119.775 ;
        RECT 84.660 119.730 84.950 119.775 ;
        RECT 82.800 119.590 84.950 119.730 ;
        RECT 82.800 119.545 83.090 119.590 ;
        RECT 84.660 119.545 84.950 119.590 ;
        RECT 21.630 119.390 21.950 119.450 ;
        RECT 20.800 119.250 21.950 119.390 ;
        RECT 17.965 119.205 18.255 119.250 ;
        RECT 20.250 119.190 20.570 119.250 ;
        RECT 21.630 119.190 21.950 119.250 ;
        RECT 22.090 119.190 22.410 119.450 ;
        RECT 23.010 119.390 23.330 119.450 ;
        RECT 23.945 119.390 24.235 119.435 ;
        RECT 23.010 119.250 24.235 119.390 ;
        RECT 23.010 119.190 23.330 119.250 ;
        RECT 23.945 119.205 24.235 119.250 ;
        RECT 29.235 119.390 29.525 119.435 ;
        RECT 30.370 119.390 30.690 119.450 ;
        RECT 34.970 119.390 35.290 119.450 ;
        RECT 29.235 119.250 35.290 119.390 ;
        RECT 29.235 119.205 29.525 119.250 ;
        RECT 30.370 119.190 30.690 119.250 ;
        RECT 34.970 119.190 35.290 119.250 ;
        RECT 44.630 119.390 44.950 119.450 ;
        RECT 45.105 119.390 45.395 119.435 ;
        RECT 44.630 119.250 45.395 119.390 ;
        RECT 44.630 119.190 44.950 119.250 ;
        RECT 45.105 119.205 45.395 119.250 ;
        RECT 54.750 119.190 55.070 119.450 ;
        RECT 59.365 119.390 59.655 119.435 ;
        RECT 62.110 119.390 62.430 119.450 ;
        RECT 86.120 119.435 86.260 119.930 ;
        RECT 86.950 119.870 87.270 120.130 ;
        RECT 91.980 120.070 92.270 120.115 ;
        RECT 95.320 120.070 95.460 120.225 ;
        RECT 95.690 120.210 96.010 120.270 ;
        RECT 97.070 120.210 97.390 120.270 ;
        RECT 97.620 120.115 97.760 120.950 ;
        RECT 97.990 120.890 98.310 121.150 ;
        RECT 99.830 121.090 100.150 121.150 ;
        RECT 100.305 121.090 100.595 121.135 ;
        RECT 99.830 120.950 100.595 121.090 ;
        RECT 99.830 120.890 100.150 120.950 ;
        RECT 100.305 120.905 100.595 120.950 ;
        RECT 120.545 121.090 120.835 121.135 ;
        RECT 121.450 121.090 121.770 121.150 ;
        RECT 120.545 120.950 121.770 121.090 ;
        RECT 120.545 120.905 120.835 120.950 ;
        RECT 121.450 120.890 121.770 120.950 ;
        RECT 121.925 121.090 122.215 121.135 ;
        RECT 124.670 121.090 124.990 121.150 ;
        RECT 121.925 120.950 124.990 121.090 ;
        RECT 121.925 120.905 122.215 120.950 ;
        RECT 124.670 120.890 124.990 120.950 ;
        RECT 119.165 120.750 119.455 120.795 ;
        RECT 117.860 120.610 119.455 120.750 ;
        RECT 115.470 120.410 115.790 120.470 ;
        RECT 115.945 120.410 116.235 120.455 ;
        RECT 115.470 120.270 116.235 120.410 ;
        RECT 115.470 120.210 115.790 120.270 ;
        RECT 115.945 120.225 116.235 120.270 ;
        RECT 91.980 119.930 94.515 120.070 ;
        RECT 95.320 119.930 97.300 120.070 ;
        RECT 91.980 119.885 92.270 119.930 ;
        RECT 90.120 119.730 90.410 119.775 ;
        RECT 91.090 119.730 91.410 119.790 ;
        RECT 94.300 119.775 94.515 119.930 ;
        RECT 93.380 119.730 93.670 119.775 ;
        RECT 90.120 119.590 93.670 119.730 ;
        RECT 90.120 119.545 90.410 119.590 ;
        RECT 91.090 119.530 91.410 119.590 ;
        RECT 93.380 119.545 93.670 119.590 ;
        RECT 94.300 119.730 94.590 119.775 ;
        RECT 96.160 119.730 96.450 119.775 ;
        RECT 94.300 119.590 96.450 119.730 ;
        RECT 97.160 119.730 97.300 119.930 ;
        RECT 97.545 119.885 97.835 120.115 ;
        RECT 98.450 120.070 98.770 120.130 ;
        RECT 99.845 120.070 100.135 120.115 ;
        RECT 98.450 119.930 100.135 120.070 ;
        RECT 98.450 119.870 98.770 119.930 ;
        RECT 99.845 119.885 100.135 119.930 ;
        RECT 101.210 119.870 101.530 120.130 ;
        RECT 102.130 119.870 102.450 120.130 ;
        RECT 112.710 120.070 113.030 120.130 ;
        RECT 116.865 120.070 117.155 120.115 ;
        RECT 112.710 119.930 117.155 120.070 ;
        RECT 112.710 119.870 113.030 119.930 ;
        RECT 116.865 119.885 117.155 119.930 ;
        RECT 117.310 119.870 117.630 120.130 ;
        RECT 110.885 119.730 111.175 119.775 ;
        RECT 111.790 119.730 112.110 119.790 ;
        RECT 113.185 119.730 113.475 119.775 ;
        RECT 97.160 119.590 99.140 119.730 ;
        RECT 94.300 119.545 94.590 119.590 ;
        RECT 96.160 119.545 96.450 119.590 ;
        RECT 59.365 119.250 62.430 119.390 ;
        RECT 59.365 119.205 59.655 119.250 ;
        RECT 62.110 119.190 62.430 119.250 ;
        RECT 86.045 119.205 86.335 119.435 ;
        RECT 88.115 119.390 88.405 119.435 ;
        RECT 88.790 119.390 89.110 119.450 ;
        RECT 99.000 119.435 99.140 119.590 ;
        RECT 110.885 119.590 113.475 119.730 ;
        RECT 117.860 119.730 118.000 120.610 ;
        RECT 119.165 120.565 119.455 120.610 ;
        RECT 118.230 120.070 118.550 120.130 ;
        RECT 119.625 120.070 119.915 120.115 ;
        RECT 118.230 119.930 119.915 120.070 ;
        RECT 118.230 119.870 118.550 119.930 ;
        RECT 119.625 119.885 119.915 119.930 ;
        RECT 121.005 119.885 121.295 120.115 ;
        RECT 121.080 119.730 121.220 119.885 ;
        RECT 117.860 119.590 121.220 119.730 ;
        RECT 110.885 119.545 111.175 119.590 ;
        RECT 111.790 119.530 112.110 119.590 ;
        RECT 113.185 119.545 113.475 119.590 ;
        RECT 88.115 119.250 89.110 119.390 ;
        RECT 88.115 119.205 88.405 119.250 ;
        RECT 88.790 119.190 89.110 119.250 ;
        RECT 98.925 119.205 99.215 119.435 ;
        RECT 113.260 119.390 113.400 119.545 ;
        RECT 119.150 119.390 119.470 119.450 ;
        RECT 113.260 119.250 119.470 119.390 ;
        RECT 119.150 119.190 119.470 119.250 ;
        RECT 14.660 118.570 127.820 119.050 ;
        RECT 18.195 118.370 18.485 118.415 ;
        RECT 22.090 118.370 22.410 118.430 ;
        RECT 18.195 118.230 22.410 118.370 ;
        RECT 18.195 118.185 18.485 118.230 ;
        RECT 22.090 118.170 22.410 118.230 ;
        RECT 29.910 118.170 30.230 118.430 ;
        RECT 37.270 118.370 37.590 118.430 ;
        RECT 37.975 118.370 38.265 118.415 ;
        RECT 37.270 118.230 38.265 118.370 ;
        RECT 37.270 118.170 37.590 118.230 ;
        RECT 37.975 118.185 38.265 118.230 ;
        RECT 49.230 118.370 49.550 118.430 ;
        RECT 51.775 118.370 52.065 118.415 ;
        RECT 49.230 118.230 52.065 118.370 ;
        RECT 49.230 118.170 49.550 118.230 ;
        RECT 51.775 118.185 52.065 118.230 ;
        RECT 61.205 118.185 61.495 118.415 ;
        RECT 66.250 118.370 66.570 118.430 ;
        RECT 67.185 118.370 67.475 118.415 ;
        RECT 66.250 118.230 67.475 118.370 ;
        RECT 20.250 118.075 20.570 118.090 ;
        RECT 20.200 118.030 20.570 118.075 ;
        RECT 23.460 118.030 23.750 118.075 ;
        RECT 20.200 117.890 23.750 118.030 ;
        RECT 20.200 117.845 20.570 117.890 ;
        RECT 23.460 117.845 23.750 117.890 ;
        RECT 24.380 118.030 24.670 118.075 ;
        RECT 26.240 118.030 26.530 118.075 ;
        RECT 24.380 117.890 26.530 118.030 ;
        RECT 24.380 117.845 24.670 117.890 ;
        RECT 26.240 117.845 26.530 117.890 ;
        RECT 20.250 117.830 20.570 117.845 ;
        RECT 22.060 117.690 22.350 117.735 ;
        RECT 24.380 117.690 24.595 117.845 ;
        RECT 22.060 117.550 24.595 117.690 ;
        RECT 27.165 117.690 27.455 117.735 ;
        RECT 30.000 117.690 30.140 118.170 ;
        RECT 36.350 117.830 36.670 118.090 ;
        RECT 40.030 118.075 40.350 118.090 ;
        RECT 39.980 118.030 40.350 118.075 ;
        RECT 43.240 118.030 43.530 118.075 ;
        RECT 39.980 117.890 43.530 118.030 ;
        RECT 39.980 117.845 40.350 117.890 ;
        RECT 43.240 117.845 43.530 117.890 ;
        RECT 44.160 118.030 44.450 118.075 ;
        RECT 46.020 118.030 46.310 118.075 ;
        RECT 44.160 117.890 46.310 118.030 ;
        RECT 44.160 117.845 44.450 117.890 ;
        RECT 46.020 117.845 46.310 117.890 ;
        RECT 53.780 118.030 54.070 118.075 ;
        RECT 54.750 118.030 55.070 118.090 ;
        RECT 57.040 118.030 57.330 118.075 ;
        RECT 53.780 117.890 57.330 118.030 ;
        RECT 53.780 117.845 54.070 117.890 ;
        RECT 40.030 117.830 40.350 117.845 ;
        RECT 27.165 117.550 30.140 117.690 ;
        RECT 41.840 117.690 42.130 117.735 ;
        RECT 44.160 117.690 44.375 117.845 ;
        RECT 54.750 117.830 55.070 117.890 ;
        RECT 57.040 117.845 57.330 117.890 ;
        RECT 57.960 118.030 58.250 118.075 ;
        RECT 59.820 118.030 60.110 118.075 ;
        RECT 57.960 117.890 60.110 118.030 ;
        RECT 57.960 117.845 58.250 117.890 ;
        RECT 59.820 117.845 60.110 117.890 ;
        RECT 41.840 117.550 44.375 117.690 ;
        RECT 46.945 117.690 47.235 117.735 ;
        RECT 49.230 117.690 49.550 117.750 ;
        RECT 46.945 117.550 49.550 117.690 ;
        RECT 22.060 117.505 22.350 117.550 ;
        RECT 27.165 117.505 27.455 117.550 ;
        RECT 41.840 117.505 42.130 117.550 ;
        RECT 46.945 117.505 47.235 117.550 ;
        RECT 49.230 117.490 49.550 117.550 ;
        RECT 49.705 117.505 49.995 117.735 ;
        RECT 55.640 117.690 55.930 117.735 ;
        RECT 57.960 117.690 58.175 117.845 ;
        RECT 55.640 117.550 58.175 117.690 ;
        RECT 58.905 117.690 59.195 117.735 ;
        RECT 61.280 117.690 61.420 118.185 ;
        RECT 66.250 118.170 66.570 118.230 ;
        RECT 67.185 118.185 67.475 118.230 ;
        RECT 69.485 118.185 69.775 118.415 ;
        RECT 76.370 118.370 76.690 118.430 ;
        RECT 76.845 118.370 77.135 118.415 ;
        RECT 76.370 118.230 77.135 118.370 ;
        RECT 58.905 117.550 61.420 117.690 ;
        RECT 55.640 117.505 55.930 117.550 ;
        RECT 58.905 117.505 59.195 117.550 ;
        RECT 25.310 117.150 25.630 117.410 ;
        RECT 45.090 117.150 45.410 117.410 ;
        RECT 48.325 117.165 48.615 117.395 ;
        RECT 22.060 117.010 22.350 117.055 ;
        RECT 24.840 117.010 25.130 117.055 ;
        RECT 26.700 117.010 26.990 117.055 ;
        RECT 22.060 116.870 26.990 117.010 ;
        RECT 22.060 116.825 22.350 116.870 ;
        RECT 24.840 116.825 25.130 116.870 ;
        RECT 26.700 116.825 26.990 116.870 ;
        RECT 41.840 117.010 42.130 117.055 ;
        RECT 44.620 117.010 44.910 117.055 ;
        RECT 46.480 117.010 46.770 117.055 ;
        RECT 41.840 116.870 46.770 117.010 ;
        RECT 41.840 116.825 42.130 116.870 ;
        RECT 44.620 116.825 44.910 116.870 ;
        RECT 46.480 116.825 46.770 116.870 ;
        RECT 36.810 116.670 37.130 116.730 ;
        RECT 39.110 116.670 39.430 116.730 ;
        RECT 48.400 116.670 48.540 117.165 ;
        RECT 49.780 117.070 49.920 117.505 ;
        RECT 62.110 117.490 62.430 117.750 ;
        RECT 63.490 117.690 63.810 117.750 ;
        RECT 63.490 117.550 66.480 117.690 ;
        RECT 63.490 117.490 63.810 117.550 ;
        RECT 60.745 117.350 61.035 117.395 ;
        RECT 63.950 117.350 64.270 117.410 ;
        RECT 66.340 117.395 66.480 117.550 ;
        RECT 67.645 117.505 67.935 117.735 ;
        RECT 69.560 117.690 69.700 118.185 ;
        RECT 76.370 118.170 76.690 118.230 ;
        RECT 76.845 118.185 77.135 118.230 ;
        RECT 88.790 118.370 89.110 118.430 ;
        RECT 93.405 118.370 93.695 118.415 ;
        RECT 88.790 118.230 93.695 118.370 ;
        RECT 88.790 118.170 89.110 118.230 ;
        RECT 93.405 118.185 93.695 118.230 ;
        RECT 95.245 118.370 95.535 118.415 ;
        RECT 98.450 118.370 98.770 118.430 ;
        RECT 95.245 118.230 98.770 118.370 ;
        RECT 95.245 118.185 95.535 118.230 ;
        RECT 98.450 118.170 98.770 118.230 ;
        RECT 106.285 118.185 106.575 118.415 ;
        RECT 79.130 118.030 79.450 118.090 ;
        RECT 78.760 117.890 79.450 118.030 ;
        RECT 70.405 117.690 70.695 117.735 ;
        RECT 69.560 117.550 70.695 117.690 ;
        RECT 70.405 117.505 70.695 117.550 ;
        RECT 74.070 117.690 74.390 117.750 ;
        RECT 78.760 117.735 78.900 117.890 ;
        RECT 79.130 117.830 79.450 117.890 ;
        RECT 80.070 118.030 80.360 118.075 ;
        RECT 81.930 118.030 82.220 118.075 ;
        RECT 80.070 117.890 82.220 118.030 ;
        RECT 80.070 117.845 80.360 117.890 ;
        RECT 81.930 117.845 82.220 117.890 ;
        RECT 82.850 118.030 83.140 118.075 ;
        RECT 86.110 118.030 86.400 118.075 ;
        RECT 89.725 118.030 90.015 118.075 ;
        RECT 82.850 117.890 90.015 118.030 ;
        RECT 82.850 117.845 83.140 117.890 ;
        RECT 86.110 117.845 86.400 117.890 ;
        RECT 89.725 117.845 90.015 117.890 ;
        RECT 92.945 118.030 93.235 118.075 ;
        RECT 93.850 118.030 94.170 118.090 ;
        RECT 106.360 118.030 106.500 118.185 ;
        RECT 109.950 118.170 110.270 118.430 ;
        RECT 112.265 118.370 112.555 118.415 ;
        RECT 112.710 118.370 113.030 118.430 ;
        RECT 112.265 118.230 113.030 118.370 ;
        RECT 112.265 118.185 112.555 118.230 ;
        RECT 112.710 118.170 113.030 118.230 ;
        RECT 111.805 118.030 112.095 118.075 ;
        RECT 92.945 117.890 94.170 118.030 ;
        RECT 92.945 117.845 93.235 117.890 ;
        RECT 76.385 117.690 76.675 117.735 ;
        RECT 74.070 117.550 76.675 117.690 ;
        RECT 60.745 117.210 64.270 117.350 ;
        RECT 60.745 117.165 61.035 117.210 ;
        RECT 63.950 117.150 64.270 117.210 ;
        RECT 66.265 117.165 66.555 117.395 ;
        RECT 49.690 116.810 50.010 117.070 ;
        RECT 55.640 117.010 55.930 117.055 ;
        RECT 58.420 117.010 58.710 117.055 ;
        RECT 60.280 117.010 60.570 117.055 ;
        RECT 55.640 116.870 60.570 117.010 ;
        RECT 55.640 116.825 55.930 116.870 ;
        RECT 58.420 116.825 58.710 116.870 ;
        RECT 60.280 116.825 60.570 116.870 ;
        RECT 36.810 116.530 48.540 116.670 ;
        RECT 57.050 116.670 57.370 116.730 ;
        RECT 67.720 116.670 67.860 117.505 ;
        RECT 74.070 117.490 74.390 117.550 ;
        RECT 76.385 117.505 76.675 117.550 ;
        RECT 78.685 117.505 78.975 117.735 ;
        RECT 80.970 117.490 81.290 117.750 ;
        RECT 82.005 117.690 82.220 117.845 ;
        RECT 93.850 117.830 94.170 117.890 ;
        RECT 94.400 117.890 106.500 118.030 ;
        RECT 106.820 117.890 112.095 118.030 ;
        RECT 84.250 117.690 84.540 117.735 ;
        RECT 82.005 117.550 84.540 117.690 ;
        RECT 84.250 117.505 84.540 117.550 ;
        RECT 90.170 117.490 90.490 117.750 ;
        RECT 94.400 117.690 94.540 117.890 ;
        RECT 92.100 117.550 94.540 117.690 ;
        RECT 103.525 117.690 103.815 117.735 ;
        RECT 103.970 117.690 104.290 117.750 ;
        RECT 103.525 117.550 104.290 117.690 ;
        RECT 74.530 117.350 74.850 117.410 ;
        RECT 79.145 117.350 79.435 117.395 ;
        RECT 81.890 117.350 82.210 117.410 ;
        RECT 74.530 117.210 82.210 117.350 ;
        RECT 74.530 117.150 74.850 117.210 ;
        RECT 79.145 117.165 79.435 117.210 ;
        RECT 81.890 117.150 82.210 117.210 ;
        RECT 86.950 117.350 87.270 117.410 ;
        RECT 88.115 117.350 88.405 117.395 ;
        RECT 92.100 117.350 92.240 117.550 ;
        RECT 103.525 117.505 103.815 117.550 ;
        RECT 103.970 117.490 104.290 117.550 ;
        RECT 106.270 117.690 106.590 117.750 ;
        RECT 106.820 117.735 106.960 117.890 ;
        RECT 111.805 117.845 112.095 117.890 ;
        RECT 106.745 117.690 107.035 117.735 ;
        RECT 106.270 117.550 107.035 117.690 ;
        RECT 106.270 117.490 106.590 117.550 ;
        RECT 106.745 117.505 107.035 117.550 ;
        RECT 109.030 117.490 109.350 117.750 ;
        RECT 113.630 117.690 113.950 117.750 ;
        RECT 117.325 117.690 117.615 117.735 ;
        RECT 113.630 117.550 117.615 117.690 ;
        RECT 113.630 117.490 113.950 117.550 ;
        RECT 117.325 117.505 117.615 117.550 ;
        RECT 118.705 117.505 118.995 117.735 ;
        RECT 86.950 117.210 92.240 117.350 ;
        RECT 92.485 117.350 92.775 117.395 ;
        RECT 105.825 117.350 106.115 117.395 ;
        RECT 110.885 117.350 111.175 117.395 ;
        RECT 118.780 117.350 118.920 117.505 ;
        RECT 92.485 117.210 111.175 117.350 ;
        RECT 86.950 117.150 87.270 117.210 ;
        RECT 88.115 117.165 88.405 117.210 ;
        RECT 92.485 117.165 92.775 117.210 ;
        RECT 105.825 117.165 106.115 117.210 ;
        RECT 110.885 117.165 111.175 117.210 ;
        RECT 114.180 117.210 118.920 117.350 ;
        RECT 68.090 117.010 68.410 117.070 ;
        RECT 77.765 117.010 78.055 117.055 ;
        RECT 68.090 116.870 78.055 117.010 ;
        RECT 68.090 116.810 68.410 116.870 ;
        RECT 77.765 116.825 78.055 116.870 ;
        RECT 79.610 117.010 79.900 117.055 ;
        RECT 81.470 117.010 81.760 117.055 ;
        RECT 84.250 117.010 84.540 117.055 ;
        RECT 79.610 116.870 84.540 117.010 ;
        RECT 79.610 116.825 79.900 116.870 ;
        RECT 81.470 116.825 81.760 116.870 ;
        RECT 84.250 116.825 84.540 116.870 ;
        RECT 85.110 117.010 85.430 117.070 ;
        RECT 92.560 117.010 92.700 117.165 ;
        RECT 114.180 117.055 114.320 117.210 ;
        RECT 85.110 116.870 92.700 117.010 ;
        RECT 85.110 116.810 85.430 116.870 ;
        RECT 114.105 116.825 114.395 117.055 ;
        RECT 57.050 116.530 67.860 116.670 ;
        RECT 36.810 116.470 37.130 116.530 ;
        RECT 39.110 116.470 39.430 116.530 ;
        RECT 57.050 116.470 57.370 116.530 ;
        RECT 71.310 116.470 71.630 116.730 ;
        RECT 103.970 116.470 104.290 116.730 ;
        RECT 108.585 116.670 108.875 116.715 ;
        RECT 109.030 116.670 109.350 116.730 ;
        RECT 108.585 116.530 109.350 116.670 ;
        RECT 108.585 116.485 108.875 116.530 ;
        RECT 109.030 116.470 109.350 116.530 ;
        RECT 116.865 116.670 117.155 116.715 ;
        RECT 117.310 116.670 117.630 116.730 ;
        RECT 116.865 116.530 117.630 116.670 ;
        RECT 116.865 116.485 117.155 116.530 ;
        RECT 117.310 116.470 117.630 116.530 ;
        RECT 119.625 116.670 119.915 116.715 ;
        RECT 120.070 116.670 120.390 116.730 ;
        RECT 119.625 116.530 120.390 116.670 ;
        RECT 119.625 116.485 119.915 116.530 ;
        RECT 120.070 116.470 120.390 116.530 ;
        RECT 14.660 115.850 127.820 116.330 ;
        RECT 23.945 115.650 24.235 115.695 ;
        RECT 25.310 115.650 25.630 115.710 ;
        RECT 23.945 115.510 25.630 115.650 ;
        RECT 23.945 115.465 24.235 115.510 ;
        RECT 25.310 115.450 25.630 115.510 ;
        RECT 28.530 115.450 28.850 115.710 ;
        RECT 29.450 115.450 29.770 115.710 ;
        RECT 35.445 115.650 35.735 115.695 ;
        RECT 35.890 115.650 36.210 115.710 ;
        RECT 35.445 115.510 36.210 115.650 ;
        RECT 35.445 115.465 35.735 115.510 ;
        RECT 35.890 115.450 36.210 115.510 ;
        RECT 36.365 115.650 36.655 115.695 ;
        RECT 40.030 115.650 40.350 115.710 ;
        RECT 36.365 115.510 40.350 115.650 ;
        RECT 36.365 115.465 36.655 115.510 ;
        RECT 40.030 115.450 40.350 115.510 ;
        RECT 45.090 115.650 45.410 115.710 ;
        RECT 45.565 115.650 45.855 115.695 ;
        RECT 45.090 115.510 45.855 115.650 ;
        RECT 45.090 115.450 45.410 115.510 ;
        RECT 45.565 115.465 45.855 115.510 ;
        RECT 65.575 115.650 65.865 115.695 ;
        RECT 66.250 115.650 66.570 115.710 ;
        RECT 65.575 115.510 66.570 115.650 ;
        RECT 65.575 115.465 65.865 115.510 ;
        RECT 66.250 115.450 66.570 115.510 ;
        RECT 80.970 115.650 81.290 115.710 ;
        RECT 89.265 115.650 89.555 115.695 ;
        RECT 80.970 115.510 89.555 115.650 ;
        RECT 80.970 115.450 81.290 115.510 ;
        RECT 89.265 115.465 89.555 115.510 ;
        RECT 102.835 115.650 103.125 115.695 ;
        RECT 106.270 115.650 106.590 115.710 ;
        RECT 102.835 115.510 106.590 115.650 ;
        RECT 102.835 115.465 103.125 115.510 ;
        RECT 106.270 115.450 106.590 115.510 ;
        RECT 112.710 115.695 113.030 115.710 ;
        RECT 112.710 115.465 113.245 115.695 ;
        RECT 112.710 115.450 113.030 115.465 ;
        RECT 58.430 115.310 58.750 115.370 ;
        RECT 56.680 115.170 58.750 115.310 ;
        RECT 21.630 114.970 21.950 115.030 ;
        RECT 30.370 114.970 30.690 115.030 ;
        RECT 31.765 114.970 32.055 115.015 ;
        RECT 21.630 114.830 28.300 114.970 ;
        RECT 21.630 114.770 21.950 114.830 ;
        RECT 23.010 114.430 23.330 114.690 ;
        RECT 28.160 114.675 28.300 114.830 ;
        RECT 30.370 114.830 32.055 114.970 ;
        RECT 30.370 114.770 30.690 114.830 ;
        RECT 31.765 114.785 32.055 114.830 ;
        RECT 32.685 114.970 32.975 115.015 ;
        RECT 36.350 114.970 36.670 115.030 ;
        RECT 56.680 115.015 56.820 115.170 ;
        RECT 58.430 115.110 58.750 115.170 ;
        RECT 69.440 115.310 69.730 115.355 ;
        RECT 72.220 115.310 72.510 115.355 ;
        RECT 74.080 115.310 74.370 115.355 ;
        RECT 69.440 115.170 74.370 115.310 ;
        RECT 69.440 115.125 69.730 115.170 ;
        RECT 72.220 115.125 72.510 115.170 ;
        RECT 74.080 115.125 74.370 115.170 ;
        RECT 106.700 115.310 106.990 115.355 ;
        RECT 109.480 115.310 109.770 115.355 ;
        RECT 111.340 115.310 111.630 115.355 ;
        RECT 106.700 115.170 111.630 115.310 ;
        RECT 106.700 115.125 106.990 115.170 ;
        RECT 109.480 115.125 109.770 115.170 ;
        RECT 111.340 115.125 111.630 115.170 ;
        RECT 116.820 115.310 117.110 115.355 ;
        RECT 119.600 115.310 119.890 115.355 ;
        RECT 121.460 115.310 121.750 115.355 ;
        RECT 116.820 115.170 121.750 115.310 ;
        RECT 116.820 115.125 117.110 115.170 ;
        RECT 119.600 115.125 119.890 115.170 ;
        RECT 121.460 115.125 121.750 115.170 ;
        RECT 32.685 114.830 36.670 114.970 ;
        RECT 32.685 114.785 32.975 114.830 ;
        RECT 36.350 114.770 36.670 114.830 ;
        RECT 56.605 114.785 56.895 115.015 ;
        RECT 57.050 114.770 57.370 115.030 ;
        RECT 71.310 114.970 71.630 115.030 ;
        RECT 72.705 114.970 72.995 115.015 ;
        RECT 71.310 114.830 72.995 114.970 ;
        RECT 71.310 114.770 71.630 114.830 ;
        RECT 72.705 114.785 72.995 114.830 ;
        RECT 74.530 114.770 74.850 115.030 ;
        RECT 85.110 114.970 85.430 115.030 ;
        RECT 85.585 114.970 85.875 115.015 ;
        RECT 85.110 114.830 85.875 114.970 ;
        RECT 85.110 114.770 85.430 114.830 ;
        RECT 85.585 114.785 85.875 114.830 ;
        RECT 111.790 114.770 112.110 115.030 ;
        RECT 119.150 114.970 119.470 115.030 ;
        RECT 119.150 114.830 119.840 114.970 ;
        RECT 119.150 114.770 119.470 114.830 ;
        RECT 28.085 114.445 28.375 114.675 ;
        RECT 28.160 114.290 28.300 114.445 ;
        RECT 31.290 114.430 31.610 114.690 ;
        RECT 34.050 114.630 34.370 114.690 ;
        RECT 34.525 114.630 34.815 114.675 ;
        RECT 34.050 114.490 34.815 114.630 ;
        RECT 34.050 114.430 34.370 114.490 ;
        RECT 34.525 114.445 34.815 114.490 ;
        RECT 35.905 114.630 36.195 114.675 ;
        RECT 36.810 114.630 37.130 114.690 ;
        RECT 35.905 114.490 37.130 114.630 ;
        RECT 35.905 114.445 36.195 114.490 ;
        RECT 35.980 114.290 36.120 114.445 ;
        RECT 36.810 114.430 37.130 114.490 ;
        RECT 44.630 114.430 44.950 114.690 ;
        RECT 57.525 114.630 57.815 114.675 ;
        RECT 57.970 114.630 58.290 114.690 ;
        RECT 57.525 114.490 58.290 114.630 ;
        RECT 57.525 114.445 57.815 114.490 ;
        RECT 57.970 114.430 58.290 114.490 ;
        RECT 69.440 114.630 69.730 114.675 ;
        RECT 75.910 114.630 76.230 114.690 ;
        RECT 86.505 114.630 86.795 114.675 ;
        RECT 69.440 114.490 71.975 114.630 ;
        RECT 69.440 114.445 69.730 114.490 ;
        RECT 28.160 114.150 36.120 114.290 ;
        RECT 67.580 114.290 67.870 114.335 ;
        RECT 69.930 114.290 70.250 114.350 ;
        RECT 71.760 114.335 71.975 114.490 ;
        RECT 75.910 114.490 86.795 114.630 ;
        RECT 75.910 114.430 76.230 114.490 ;
        RECT 86.505 114.445 86.795 114.490 ;
        RECT 86.950 114.430 87.270 114.690 ;
        RECT 90.185 114.630 90.475 114.675 ;
        RECT 88.880 114.490 90.475 114.630 ;
        RECT 70.840 114.290 71.130 114.335 ;
        RECT 67.580 114.150 71.130 114.290 ;
        RECT 67.580 114.105 67.870 114.150 ;
        RECT 69.930 114.090 70.250 114.150 ;
        RECT 70.840 114.105 71.130 114.150 ;
        RECT 71.760 114.290 72.050 114.335 ;
        RECT 73.620 114.290 73.910 114.335 ;
        RECT 71.760 114.150 73.910 114.290 ;
        RECT 71.760 114.105 72.050 114.150 ;
        RECT 73.620 114.105 73.910 114.150 ;
        RECT 59.350 113.750 59.670 114.010 ;
        RECT 88.880 113.995 89.020 114.490 ;
        RECT 90.185 114.445 90.475 114.490 ;
        RECT 106.700 114.630 106.990 114.675 ;
        RECT 109.490 114.630 109.810 114.690 ;
        RECT 109.965 114.630 110.255 114.675 ;
        RECT 106.700 114.490 109.235 114.630 ;
        RECT 106.700 114.445 106.990 114.490 ;
        RECT 103.970 114.290 104.290 114.350 ;
        RECT 109.020 114.335 109.235 114.490 ;
        RECT 109.490 114.490 110.255 114.630 ;
        RECT 109.490 114.430 109.810 114.490 ;
        RECT 109.965 114.445 110.255 114.490 ;
        RECT 116.820 114.630 117.110 114.675 ;
        RECT 119.700 114.630 119.840 114.830 ;
        RECT 120.070 114.770 120.390 115.030 ;
        RECT 121.925 114.630 122.215 114.675 ;
        RECT 126.050 114.630 126.370 114.690 ;
        RECT 116.820 114.490 119.355 114.630 ;
        RECT 119.700 114.490 126.370 114.630 ;
        RECT 116.820 114.445 117.110 114.490 ;
        RECT 104.840 114.290 105.130 114.335 ;
        RECT 108.100 114.290 108.390 114.335 ;
        RECT 103.970 114.150 108.390 114.290 ;
        RECT 103.970 114.090 104.290 114.150 ;
        RECT 104.840 114.105 105.130 114.150 ;
        RECT 108.100 114.105 108.390 114.150 ;
        RECT 109.020 114.290 109.310 114.335 ;
        RECT 110.880 114.290 111.170 114.335 ;
        RECT 109.020 114.150 111.170 114.290 ;
        RECT 109.020 114.105 109.310 114.150 ;
        RECT 110.880 114.105 111.170 114.150 ;
        RECT 114.960 114.290 115.250 114.335 ;
        RECT 117.310 114.290 117.630 114.350 ;
        RECT 119.140 114.335 119.355 114.490 ;
        RECT 121.925 114.445 122.215 114.490 ;
        RECT 126.050 114.430 126.370 114.490 ;
        RECT 118.220 114.290 118.510 114.335 ;
        RECT 114.960 114.150 118.510 114.290 ;
        RECT 114.960 114.105 115.250 114.150 ;
        RECT 117.310 114.090 117.630 114.150 ;
        RECT 118.220 114.105 118.510 114.150 ;
        RECT 119.140 114.290 119.430 114.335 ;
        RECT 121.000 114.290 121.290 114.335 ;
        RECT 119.140 114.150 121.290 114.290 ;
        RECT 119.140 114.105 119.430 114.150 ;
        RECT 121.000 114.105 121.290 114.150 ;
        RECT 88.805 113.765 89.095 113.995 ;
        RECT 14.660 113.130 127.820 113.610 ;
        RECT 53.155 112.930 53.445 112.975 ;
        RECT 57.050 112.930 57.370 112.990 ;
        RECT 53.155 112.790 57.370 112.930 ;
        RECT 53.155 112.745 53.445 112.790 ;
        RECT 57.050 112.730 57.370 112.790 ;
        RECT 69.485 112.930 69.775 112.975 ;
        RECT 69.930 112.930 70.250 112.990 ;
        RECT 69.485 112.790 70.250 112.930 ;
        RECT 69.485 112.745 69.775 112.790 ;
        RECT 69.930 112.730 70.250 112.790 ;
        RECT 109.490 112.730 109.810 112.990 ;
        RECT 118.690 112.930 119.010 112.990 ;
        RECT 122.385 112.930 122.675 112.975 ;
        RECT 118.690 112.790 122.675 112.930 ;
        RECT 118.690 112.730 119.010 112.790 ;
        RECT 122.385 112.745 122.675 112.790 ;
        RECT 22.205 112.590 22.495 112.635 ;
        RECT 25.445 112.590 26.095 112.635 ;
        RECT 22.205 112.450 26.095 112.590 ;
        RECT 22.205 112.405 22.795 112.450 ;
        RECT 25.445 112.405 26.095 112.450 ;
        RECT 55.160 112.590 55.450 112.635 ;
        RECT 56.590 112.590 56.910 112.650 ;
        RECT 58.420 112.590 58.710 112.635 ;
        RECT 55.160 112.450 58.710 112.590 ;
        RECT 55.160 112.405 55.450 112.450 ;
        RECT 22.505 112.310 22.795 112.405 ;
        RECT 56.590 112.390 56.910 112.450 ;
        RECT 58.420 112.405 58.710 112.450 ;
        RECT 59.340 112.590 59.630 112.635 ;
        RECT 61.200 112.590 61.490 112.635 ;
        RECT 59.340 112.450 61.490 112.590 ;
        RECT 59.340 112.405 59.630 112.450 ;
        RECT 61.200 112.405 61.490 112.450 ;
        RECT 119.610 112.590 119.930 112.650 ;
        RECT 119.610 112.450 123.520 112.590 ;
        RECT 22.505 112.090 22.870 112.310 ;
        RECT 22.550 112.050 22.870 112.090 ;
        RECT 23.585 112.250 23.875 112.295 ;
        RECT 27.165 112.250 27.455 112.295 ;
        RECT 29.000 112.250 29.290 112.295 ;
        RECT 23.585 112.110 29.290 112.250 ;
        RECT 23.585 112.065 23.875 112.110 ;
        RECT 27.165 112.065 27.455 112.110 ;
        RECT 29.000 112.065 29.290 112.110 ;
        RECT 29.465 112.250 29.755 112.295 ;
        RECT 29.910 112.250 30.230 112.310 ;
        RECT 29.465 112.110 30.230 112.250 ;
        RECT 29.465 112.065 29.755 112.110 ;
        RECT 29.910 112.050 30.230 112.110 ;
        RECT 38.190 112.250 38.510 112.310 ;
        RECT 41.885 112.250 42.175 112.295 ;
        RECT 38.190 112.110 42.175 112.250 ;
        RECT 38.190 112.050 38.510 112.110 ;
        RECT 41.885 112.065 42.175 112.110 ;
        RECT 57.020 112.250 57.310 112.295 ;
        RECT 59.340 112.250 59.555 112.405 ;
        RECT 119.610 112.390 119.930 112.450 ;
        RECT 57.020 112.110 59.555 112.250 ;
        RECT 62.125 112.250 62.415 112.295 ;
        RECT 63.950 112.250 64.270 112.310 ;
        RECT 62.125 112.110 64.270 112.250 ;
        RECT 57.020 112.065 57.310 112.110 ;
        RECT 62.125 112.065 62.415 112.110 ;
        RECT 63.950 112.050 64.270 112.110 ;
        RECT 67.170 112.250 67.490 112.310 ;
        RECT 69.930 112.250 70.250 112.310 ;
        RECT 67.170 112.110 70.250 112.250 ;
        RECT 67.170 112.050 67.490 112.110 ;
        RECT 69.930 112.050 70.250 112.110 ;
        RECT 98.910 112.050 99.230 112.310 ;
        RECT 108.585 112.250 108.875 112.295 ;
        RECT 109.030 112.250 109.350 112.310 ;
        RECT 108.585 112.110 109.350 112.250 ;
        RECT 108.585 112.065 108.875 112.110 ;
        RECT 109.030 112.050 109.350 112.110 ;
        RECT 120.530 112.250 120.850 112.310 ;
        RECT 123.380 112.295 123.520 112.450 ;
        RECT 121.005 112.250 121.295 112.295 ;
        RECT 120.530 112.110 121.295 112.250 ;
        RECT 120.530 112.050 120.850 112.110 ;
        RECT 121.005 112.065 121.295 112.110 ;
        RECT 123.305 112.065 123.595 112.295 ;
        RECT 20.710 111.710 21.030 111.970 ;
        RECT 60.270 111.710 60.590 111.970 ;
        RECT 23.585 111.570 23.875 111.615 ;
        RECT 26.705 111.570 26.995 111.615 ;
        RECT 28.595 111.570 28.885 111.615 ;
        RECT 23.585 111.430 28.885 111.570 ;
        RECT 23.585 111.385 23.875 111.430 ;
        RECT 26.705 111.385 26.995 111.430 ;
        RECT 28.595 111.385 28.885 111.430 ;
        RECT 46.010 111.570 46.330 111.630 ;
        RECT 49.230 111.570 49.550 111.630 ;
        RECT 46.010 111.430 49.550 111.570 ;
        RECT 46.010 111.370 46.330 111.430 ;
        RECT 49.230 111.370 49.550 111.430 ;
        RECT 57.020 111.570 57.310 111.615 ;
        RECT 59.800 111.570 60.090 111.615 ;
        RECT 61.660 111.570 61.950 111.615 ;
        RECT 57.020 111.430 61.950 111.570 ;
        RECT 57.020 111.385 57.310 111.430 ;
        RECT 59.800 111.385 60.090 111.430 ;
        RECT 61.660 111.385 61.950 111.430 ;
        RECT 28.180 111.230 28.470 111.275 ;
        RECT 28.990 111.230 29.310 111.290 ;
        RECT 28.180 111.090 29.310 111.230 ;
        RECT 28.180 111.045 28.470 111.090 ;
        RECT 28.990 111.030 29.310 111.090 ;
        RECT 42.790 111.030 43.110 111.290 ;
        RECT 99.830 111.030 100.150 111.290 ;
        RECT 121.925 111.230 122.215 111.275 ;
        RECT 124.670 111.230 124.990 111.290 ;
        RECT 121.925 111.090 124.990 111.230 ;
        RECT 121.925 111.045 122.215 111.090 ;
        RECT 124.670 111.030 124.990 111.090 ;
        RECT 14.660 110.410 127.820 110.890 ;
        RECT 22.550 110.210 22.870 110.270 ;
        RECT 23.485 110.210 23.775 110.255 ;
        RECT 22.550 110.070 23.775 110.210 ;
        RECT 22.550 110.010 22.870 110.070 ;
        RECT 23.485 110.025 23.775 110.070 ;
        RECT 40.950 110.210 41.270 110.270 ;
        RECT 40.950 110.070 45.320 110.210 ;
        RECT 40.950 110.010 41.270 110.070 ;
        RECT 28.990 109.870 29.310 109.930 ;
        RECT 32.685 109.870 32.975 109.915 ;
        RECT 28.990 109.730 32.975 109.870 ;
        RECT 28.990 109.670 29.310 109.730 ;
        RECT 32.685 109.685 32.975 109.730 ;
        RECT 38.305 109.870 38.595 109.915 ;
        RECT 41.425 109.870 41.715 109.915 ;
        RECT 43.315 109.870 43.605 109.915 ;
        RECT 38.305 109.730 43.605 109.870 ;
        RECT 38.305 109.685 38.595 109.730 ;
        RECT 41.425 109.685 41.715 109.730 ;
        RECT 43.315 109.685 43.605 109.730 ;
        RECT 34.970 109.530 35.290 109.590 ;
        RECT 33.680 109.390 35.290 109.530 ;
        RECT 18.870 109.190 19.190 109.250 ;
        RECT 23.025 109.190 23.315 109.235 ;
        RECT 26.245 109.190 26.535 109.235 ;
        RECT 18.870 109.050 26.535 109.190 ;
        RECT 18.870 108.990 19.190 109.050 ;
        RECT 23.025 109.005 23.315 109.050 ;
        RECT 26.245 109.005 26.535 109.050 ;
        RECT 26.705 109.190 26.995 109.235 ;
        RECT 27.610 109.190 27.930 109.250 ;
        RECT 26.705 109.050 27.930 109.190 ;
        RECT 26.705 109.005 26.995 109.050 ;
        RECT 26.320 108.850 26.460 109.005 ;
        RECT 27.610 108.990 27.930 109.050 ;
        RECT 29.925 109.005 30.215 109.235 ;
        RECT 30.830 109.190 31.150 109.250 ;
        RECT 33.680 109.235 33.820 109.390 ;
        RECT 34.970 109.330 35.290 109.390 ;
        RECT 35.445 109.530 35.735 109.575 ;
        RECT 37.730 109.530 38.050 109.590 ;
        RECT 35.445 109.390 38.050 109.530 ;
        RECT 35.445 109.345 35.735 109.390 ;
        RECT 37.730 109.330 38.050 109.390 ;
        RECT 42.790 109.330 43.110 109.590 ;
        RECT 32.225 109.190 32.515 109.235 ;
        RECT 30.830 109.050 32.515 109.190 ;
        RECT 30.000 108.850 30.140 109.005 ;
        RECT 30.830 108.990 31.150 109.050 ;
        RECT 32.225 109.005 32.515 109.050 ;
        RECT 33.605 109.005 33.895 109.235 ;
        RECT 34.065 109.190 34.355 109.235 ;
        RECT 34.510 109.190 34.830 109.250 ;
        RECT 45.180 109.235 45.320 110.070 ;
        RECT 56.590 110.010 56.910 110.270 ;
        RECT 60.270 110.010 60.590 110.270 ;
        RECT 70.850 110.210 71.170 110.270 ;
        RECT 75.005 110.210 75.295 110.255 ;
        RECT 70.850 110.070 75.295 110.210 ;
        RECT 70.850 110.010 71.170 110.070 ;
        RECT 75.005 110.025 75.295 110.070 ;
        RECT 95.345 109.870 95.635 109.915 ;
        RECT 98.465 109.870 98.755 109.915 ;
        RECT 100.355 109.870 100.645 109.915 ;
        RECT 95.345 109.730 100.645 109.870 ;
        RECT 95.345 109.685 95.635 109.730 ;
        RECT 98.465 109.685 98.755 109.730 ;
        RECT 100.355 109.685 100.645 109.730 ;
        RECT 120.185 109.870 120.475 109.915 ;
        RECT 123.305 109.870 123.595 109.915 ;
        RECT 125.195 109.870 125.485 109.915 ;
        RECT 120.185 109.730 125.485 109.870 ;
        RECT 120.185 109.685 120.475 109.730 ;
        RECT 123.305 109.685 123.595 109.730 ;
        RECT 125.195 109.685 125.485 109.730 ;
        RECT 69.930 109.530 70.250 109.590 ;
        RECT 84.650 109.530 84.970 109.590 ;
        RECT 92.485 109.530 92.775 109.575 ;
        RECT 97.990 109.530 98.310 109.590 ;
        RECT 56.220 109.390 70.250 109.530 ;
        RECT 34.065 109.050 34.830 109.190 ;
        RECT 34.065 109.005 34.355 109.050 ;
        RECT 34.510 108.990 34.830 109.050 ;
        RECT 35.890 108.850 36.210 108.910 ;
        RECT 37.225 108.895 37.515 109.210 ;
        RECT 38.305 109.190 38.595 109.235 ;
        RECT 41.885 109.190 42.175 109.235 ;
        RECT 43.720 109.190 44.010 109.235 ;
        RECT 38.305 109.050 44.010 109.190 ;
        RECT 38.305 109.005 38.595 109.050 ;
        RECT 41.885 109.005 42.175 109.050 ;
        RECT 43.720 109.005 44.010 109.050 ;
        RECT 44.185 109.005 44.475 109.235 ;
        RECT 45.105 109.005 45.395 109.235 ;
        RECT 49.690 109.190 50.010 109.250 ;
        RECT 56.220 109.235 56.360 109.390 ;
        RECT 69.930 109.330 70.250 109.390 ;
        RECT 79.220 109.390 82.580 109.530 ;
        RECT 56.145 109.190 56.435 109.235 ;
        RECT 49.690 109.050 56.435 109.190 ;
        RECT 26.320 108.710 36.210 108.850 ;
        RECT 35.890 108.650 36.210 108.710 ;
        RECT 36.925 108.850 37.515 108.895 ;
        RECT 39.110 108.850 39.430 108.910 ;
        RECT 40.165 108.850 40.815 108.895 ;
        RECT 36.925 108.710 40.815 108.850 ;
        RECT 36.925 108.665 37.215 108.710 ;
        RECT 39.110 108.650 39.430 108.710 ;
        RECT 40.165 108.665 40.815 108.710 ;
        RECT 25.770 108.310 26.090 108.570 ;
        RECT 27.625 108.510 27.915 108.555 ;
        RECT 28.530 108.510 28.850 108.570 ;
        RECT 27.625 108.370 28.850 108.510 ;
        RECT 27.625 108.325 27.915 108.370 ;
        RECT 28.530 108.310 28.850 108.370 ;
        RECT 30.370 108.310 30.690 108.570 ;
        RECT 31.290 108.310 31.610 108.570 ;
        RECT 34.970 108.310 35.290 108.570 ;
        RECT 35.430 108.510 35.750 108.570 ;
        RECT 44.260 108.510 44.400 109.005 ;
        RECT 49.690 108.990 50.010 109.050 ;
        RECT 56.145 109.005 56.435 109.050 ;
        RECT 59.350 108.990 59.670 109.250 ;
        RECT 67.630 108.990 67.950 109.250 ;
        RECT 48.325 108.850 48.615 108.895 ;
        RECT 70.020 108.850 70.160 109.330 ;
        RECT 75.465 109.190 75.755 109.235 ;
        RECT 76.370 109.190 76.690 109.250 ;
        RECT 79.220 109.235 79.360 109.390 ;
        RECT 75.465 109.050 76.690 109.190 ;
        RECT 75.465 109.005 75.755 109.050 ;
        RECT 76.370 108.990 76.690 109.050 ;
        RECT 79.145 109.005 79.435 109.235 ;
        RECT 79.590 108.990 79.910 109.250 ;
        RECT 82.440 109.235 82.580 109.390 ;
        RECT 84.650 109.390 91.320 109.530 ;
        RECT 84.650 109.330 84.970 109.390 ;
        RECT 80.985 109.005 81.275 109.235 ;
        RECT 82.365 109.190 82.655 109.235 ;
        RECT 86.965 109.190 87.255 109.235 ;
        RECT 89.710 109.190 90.030 109.250 ;
        RECT 91.180 109.235 91.320 109.390 ;
        RECT 92.485 109.390 98.310 109.530 ;
        RECT 92.485 109.345 92.775 109.390 ;
        RECT 97.990 109.330 98.310 109.390 ;
        RECT 99.830 109.330 100.150 109.590 ;
        RECT 101.225 109.530 101.515 109.575 ;
        RECT 109.490 109.530 109.810 109.590 ;
        RECT 101.225 109.390 109.810 109.530 ;
        RECT 101.225 109.345 101.515 109.390 ;
        RECT 109.490 109.330 109.810 109.390 ;
        RECT 117.325 109.530 117.615 109.575 ;
        RECT 121.450 109.530 121.770 109.590 ;
        RECT 117.325 109.390 121.770 109.530 ;
        RECT 117.325 109.345 117.615 109.390 ;
        RECT 121.450 109.330 121.770 109.390 ;
        RECT 124.670 109.330 124.990 109.590 ;
        RECT 126.050 109.330 126.370 109.590 ;
        RECT 82.365 109.050 90.030 109.190 ;
        RECT 82.365 109.005 82.655 109.050 ;
        RECT 86.965 109.005 87.255 109.050 ;
        RECT 81.060 108.850 81.200 109.005 ;
        RECT 89.710 108.990 90.030 109.050 ;
        RECT 91.105 109.005 91.395 109.235 ;
        RECT 94.265 108.895 94.555 109.210 ;
        RECT 95.345 109.190 95.635 109.235 ;
        RECT 98.925 109.190 99.215 109.235 ;
        RECT 100.760 109.190 101.050 109.235 ;
        RECT 95.345 109.050 101.050 109.190 ;
        RECT 95.345 109.005 95.635 109.050 ;
        RECT 98.925 109.005 99.215 109.050 ;
        RECT 100.760 109.005 101.050 109.050 ;
        RECT 103.525 109.005 103.815 109.235 ;
        RECT 103.970 109.190 104.290 109.250 ;
        RECT 104.445 109.190 104.735 109.235 ;
        RECT 103.970 109.050 104.735 109.190 ;
        RECT 97.530 108.895 97.850 108.910 ;
        RECT 48.325 108.710 49.920 108.850 ;
        RECT 70.020 108.710 81.200 108.850 ;
        RECT 93.965 108.850 94.555 108.895 ;
        RECT 97.205 108.850 97.855 108.895 ;
        RECT 93.965 108.710 97.855 108.850 ;
        RECT 48.325 108.665 48.615 108.710 ;
        RECT 49.780 108.570 49.920 108.710 ;
        RECT 93.965 108.665 94.255 108.710 ;
        RECT 97.205 108.665 97.855 108.710 ;
        RECT 99.370 108.850 99.690 108.910 ;
        RECT 103.600 108.850 103.740 109.005 ;
        RECT 103.970 108.990 104.290 109.050 ;
        RECT 104.445 109.005 104.735 109.050 ;
        RECT 108.125 109.005 108.415 109.235 ;
        RECT 115.945 109.190 116.235 109.235 ;
        RECT 111.880 109.050 116.235 109.190 ;
        RECT 108.200 108.850 108.340 109.005 ;
        RECT 111.880 108.910 112.020 109.050 ;
        RECT 115.945 109.005 116.235 109.050 ;
        RECT 111.790 108.850 112.110 108.910 ;
        RECT 99.370 108.710 112.110 108.850 ;
        RECT 97.530 108.650 97.850 108.665 ;
        RECT 99.370 108.650 99.690 108.710 ;
        RECT 111.790 108.650 112.110 108.710 ;
        RECT 112.250 108.850 112.570 108.910 ;
        RECT 119.105 108.895 119.395 109.210 ;
        RECT 120.185 109.190 120.475 109.235 ;
        RECT 123.765 109.190 124.055 109.235 ;
        RECT 125.600 109.190 125.890 109.235 ;
        RECT 120.185 109.050 125.890 109.190 ;
        RECT 120.185 109.005 120.475 109.050 ;
        RECT 123.765 109.005 124.055 109.050 ;
        RECT 125.600 109.005 125.890 109.050 ;
        RECT 118.805 108.850 119.395 108.895 ;
        RECT 122.045 108.850 122.695 108.895 ;
        RECT 112.250 108.710 122.695 108.850 ;
        RECT 112.250 108.650 112.570 108.710 ;
        RECT 118.805 108.665 119.095 108.710 ;
        RECT 122.045 108.665 122.695 108.710 ;
        RECT 35.430 108.370 44.400 108.510 ;
        RECT 46.025 108.510 46.315 108.555 ;
        RECT 46.470 108.510 46.790 108.570 ;
        RECT 46.025 108.370 46.790 108.510 ;
        RECT 35.430 108.310 35.750 108.370 ;
        RECT 46.025 108.325 46.315 108.370 ;
        RECT 46.470 108.310 46.790 108.370 ;
        RECT 49.690 108.310 50.010 108.570 ;
        RECT 68.565 108.510 68.855 108.555 ;
        RECT 70.850 108.510 71.170 108.570 ;
        RECT 68.565 108.370 71.170 108.510 ;
        RECT 68.565 108.325 68.855 108.370 ;
        RECT 70.850 108.310 71.170 108.370 ;
        RECT 78.685 108.510 78.975 108.555 ;
        RECT 79.130 108.510 79.450 108.570 ;
        RECT 78.685 108.370 79.450 108.510 ;
        RECT 78.685 108.325 78.975 108.370 ;
        RECT 79.130 108.310 79.450 108.370 ;
        RECT 80.510 108.310 80.830 108.570 ;
        RECT 87.410 108.310 87.730 108.570 ;
        RECT 90.170 108.310 90.490 108.570 ;
        RECT 92.025 108.510 92.315 108.555 ;
        RECT 96.610 108.510 96.930 108.570 ;
        RECT 92.025 108.370 96.930 108.510 ;
        RECT 92.025 108.325 92.315 108.370 ;
        RECT 96.610 108.310 96.930 108.370 ;
        RECT 103.065 108.510 103.355 108.555 ;
        RECT 103.510 108.510 103.830 108.570 ;
        RECT 103.065 108.370 103.830 108.510 ;
        RECT 103.065 108.325 103.355 108.370 ;
        RECT 103.510 108.310 103.830 108.370 ;
        RECT 105.365 108.510 105.655 108.555 ;
        RECT 105.810 108.510 106.130 108.570 ;
        RECT 105.365 108.370 106.130 108.510 ;
        RECT 105.365 108.325 105.655 108.370 ;
        RECT 105.810 108.310 106.130 108.370 ;
        RECT 106.270 108.510 106.590 108.570 ;
        RECT 107.665 108.510 107.955 108.555 ;
        RECT 106.270 108.370 107.955 108.510 ;
        RECT 106.270 108.310 106.590 108.370 ;
        RECT 107.665 108.325 107.955 108.370 ;
        RECT 116.405 108.510 116.695 108.555 ;
        RECT 120.990 108.510 121.310 108.570 ;
        RECT 116.405 108.370 121.310 108.510 ;
        RECT 116.405 108.325 116.695 108.370 ;
        RECT 120.990 108.310 121.310 108.370 ;
        RECT 14.660 107.690 127.820 108.170 ;
        RECT 31.290 107.490 31.610 107.550 ;
        RECT 26.320 107.350 31.610 107.490 ;
        RECT 20.365 107.150 20.655 107.195 ;
        RECT 23.605 107.150 24.255 107.195 ;
        RECT 25.770 107.150 26.090 107.210 ;
        RECT 26.320 107.195 26.460 107.350 ;
        RECT 31.290 107.290 31.610 107.350 ;
        RECT 42.330 107.490 42.650 107.550 ;
        RECT 48.785 107.490 49.075 107.535 ;
        RECT 42.330 107.350 49.075 107.490 ;
        RECT 42.330 107.290 42.650 107.350 ;
        RECT 48.785 107.305 49.075 107.350 ;
        RECT 52.465 107.490 52.755 107.535 ;
        RECT 52.910 107.490 53.230 107.550 ;
        RECT 52.465 107.350 53.230 107.490 ;
        RECT 52.465 107.305 52.755 107.350 ;
        RECT 52.910 107.290 53.230 107.350 ;
        RECT 79.130 107.290 79.450 107.550 ;
        RECT 97.530 107.490 97.850 107.550 ;
        RECT 98.925 107.490 99.215 107.535 ;
        RECT 97.530 107.350 99.215 107.490 ;
        RECT 97.530 107.290 97.850 107.350 ;
        RECT 98.925 107.305 99.215 107.350 ;
        RECT 112.250 107.290 112.570 107.550 ;
        RECT 20.365 107.010 26.090 107.150 ;
        RECT 20.365 106.965 20.955 107.010 ;
        RECT 23.605 106.965 24.255 107.010 ;
        RECT 18.425 106.810 18.715 106.855 ;
        RECT 18.870 106.810 19.190 106.870 ;
        RECT 18.425 106.670 19.190 106.810 ;
        RECT 18.425 106.625 18.715 106.670 ;
        RECT 18.870 106.610 19.190 106.670 ;
        RECT 20.665 106.650 20.955 106.965 ;
        RECT 25.770 106.950 26.090 107.010 ;
        RECT 26.245 106.965 26.535 107.195 ;
        RECT 29.565 107.150 29.855 107.195 ;
        RECT 30.370 107.150 30.690 107.210 ;
        RECT 32.805 107.150 33.455 107.195 ;
        RECT 29.565 107.010 33.455 107.150 ;
        RECT 29.565 106.965 30.155 107.010 ;
        RECT 21.745 106.810 22.035 106.855 ;
        RECT 25.325 106.810 25.615 106.855 ;
        RECT 27.160 106.810 27.450 106.855 ;
        RECT 21.745 106.670 27.450 106.810 ;
        RECT 21.745 106.625 22.035 106.670 ;
        RECT 25.325 106.625 25.615 106.670 ;
        RECT 27.160 106.625 27.450 106.670 ;
        RECT 29.865 106.650 30.155 106.965 ;
        RECT 30.370 106.950 30.690 107.010 ;
        RECT 32.805 106.965 33.455 107.010 ;
        RECT 34.970 107.150 35.290 107.210 ;
        RECT 35.445 107.150 35.735 107.195 ;
        RECT 34.970 107.010 35.735 107.150 ;
        RECT 34.970 106.950 35.290 107.010 ;
        RECT 35.445 106.965 35.735 107.010 ;
        RECT 35.890 107.150 36.210 107.210 ;
        RECT 38.665 107.150 38.955 107.195 ;
        RECT 41.065 107.150 41.355 107.195 ;
        RECT 44.305 107.150 44.955 107.195 ;
        RECT 35.890 107.010 38.420 107.150 ;
        RECT 35.890 106.950 36.210 107.010 ;
        RECT 38.280 106.855 38.420 107.010 ;
        RECT 38.665 107.010 44.955 107.150 ;
        RECT 38.665 106.965 38.955 107.010 ;
        RECT 41.065 106.965 41.655 107.010 ;
        RECT 44.305 106.965 44.955 107.010 ;
        RECT 46.470 107.150 46.790 107.210 ;
        RECT 46.945 107.150 47.235 107.195 ;
        RECT 46.470 107.010 47.235 107.150 ;
        RECT 30.945 106.810 31.235 106.855 ;
        RECT 34.525 106.810 34.815 106.855 ;
        RECT 36.360 106.810 36.650 106.855 ;
        RECT 30.945 106.670 36.650 106.810 ;
        RECT 30.945 106.625 31.235 106.670 ;
        RECT 34.525 106.625 34.815 106.670 ;
        RECT 36.360 106.625 36.650 106.670 ;
        RECT 38.205 106.810 38.495 106.855 ;
        RECT 38.205 106.670 38.880 106.810 ;
        RECT 38.205 106.625 38.495 106.670 ;
        RECT 38.740 106.530 38.880 106.670 ;
        RECT 41.365 106.650 41.655 106.965 ;
        RECT 46.470 106.950 46.790 107.010 ;
        RECT 46.945 106.965 47.235 107.010 ;
        RECT 50.150 107.150 50.470 107.210 ;
        RECT 64.985 107.150 65.275 107.195 ;
        RECT 68.225 107.150 68.875 107.195 ;
        RECT 50.150 107.010 54.980 107.150 ;
        RECT 50.150 106.950 50.470 107.010 ;
        RECT 42.445 106.810 42.735 106.855 ;
        RECT 46.025 106.810 46.315 106.855 ;
        RECT 47.860 106.810 48.150 106.855 ;
        RECT 42.445 106.670 48.150 106.810 ;
        RECT 42.445 106.625 42.735 106.670 ;
        RECT 46.025 106.625 46.315 106.670 ;
        RECT 47.860 106.625 48.150 106.670 ;
        RECT 49.230 106.810 49.550 106.870 ;
        RECT 49.705 106.810 49.995 106.855 ;
        RECT 49.230 106.670 49.995 106.810 ;
        RECT 49.230 106.610 49.550 106.670 ;
        RECT 49.705 106.625 49.995 106.670 ;
        RECT 51.070 106.810 51.390 106.870 ;
        RECT 54.840 106.855 54.980 107.010 ;
        RECT 64.985 107.010 68.875 107.150 ;
        RECT 64.985 106.965 65.575 107.010 ;
        RECT 68.225 106.965 68.875 107.010 ;
        RECT 65.285 106.870 65.575 106.965 ;
        RECT 70.850 106.950 71.170 107.210 ;
        RECT 75.105 107.150 75.395 107.195 ;
        RECT 78.345 107.150 78.995 107.195 ;
        RECT 79.220 107.150 79.360 107.290 ;
        RECT 75.105 107.010 79.360 107.150 ;
        RECT 80.510 107.150 80.830 107.210 ;
        RECT 80.985 107.150 81.275 107.195 ;
        RECT 80.510 107.010 81.275 107.150 ;
        RECT 75.105 106.965 75.695 107.010 ;
        RECT 78.345 106.965 78.995 107.010 ;
        RECT 51.545 106.810 51.835 106.855 ;
        RECT 51.070 106.670 51.835 106.810 ;
        RECT 51.070 106.610 51.390 106.670 ;
        RECT 51.545 106.625 51.835 106.670 ;
        RECT 54.765 106.625 55.055 106.855 ;
        RECT 55.670 106.810 55.990 106.870 ;
        RECT 61.665 106.810 61.955 106.855 ;
        RECT 55.670 106.670 61.955 106.810 ;
        RECT 55.670 106.610 55.990 106.670 ;
        RECT 61.665 106.625 61.955 106.670 ;
        RECT 65.285 106.650 65.650 106.870 ;
        RECT 65.330 106.610 65.650 106.650 ;
        RECT 66.365 106.810 66.655 106.855 ;
        RECT 69.945 106.810 70.235 106.855 ;
        RECT 71.780 106.810 72.070 106.855 ;
        RECT 66.365 106.670 72.070 106.810 ;
        RECT 66.365 106.625 66.655 106.670 ;
        RECT 69.945 106.625 70.235 106.670 ;
        RECT 71.780 106.625 72.070 106.670 ;
        RECT 75.405 106.650 75.695 106.965 ;
        RECT 80.510 106.950 80.830 107.010 ;
        RECT 80.985 106.965 81.275 107.010 ;
        RECT 82.350 107.150 82.670 107.210 ;
        RECT 90.170 107.150 90.490 107.210 ;
        RECT 90.745 107.150 91.035 107.195 ;
        RECT 93.985 107.150 94.635 107.195 ;
        RECT 82.350 107.010 86.720 107.150 ;
        RECT 82.350 106.950 82.670 107.010 ;
        RECT 76.485 106.810 76.775 106.855 ;
        RECT 80.065 106.810 80.355 106.855 ;
        RECT 81.900 106.810 82.190 106.855 ;
        RECT 76.485 106.670 82.190 106.810 ;
        RECT 76.485 106.625 76.775 106.670 ;
        RECT 80.065 106.625 80.355 106.670 ;
        RECT 81.900 106.625 82.190 106.670 ;
        RECT 82.810 106.610 83.130 106.870 ;
        RECT 86.580 106.855 86.720 107.010 ;
        RECT 90.170 107.010 94.635 107.150 ;
        RECT 90.170 106.950 90.490 107.010 ;
        RECT 90.745 106.965 91.335 107.010 ;
        RECT 93.985 106.965 94.635 107.010 ;
        RECT 85.125 106.625 85.415 106.855 ;
        RECT 86.505 106.625 86.795 106.855 ;
        RECT 91.045 106.650 91.335 106.965 ;
        RECT 96.610 106.950 96.930 107.210 ;
        RECT 97.070 107.150 97.390 107.210 ;
        RECT 101.325 107.150 101.615 107.195 ;
        RECT 103.510 107.150 103.830 107.210 ;
        RECT 104.565 107.150 105.215 107.195 ;
        RECT 97.070 107.010 98.220 107.150 ;
        RECT 97.070 106.950 97.390 107.010 ;
        RECT 98.080 106.855 98.220 107.010 ;
        RECT 101.325 107.010 105.215 107.150 ;
        RECT 101.325 106.965 101.915 107.010 ;
        RECT 92.125 106.810 92.415 106.855 ;
        RECT 95.705 106.810 95.995 106.855 ;
        RECT 97.540 106.810 97.830 106.855 ;
        RECT 92.125 106.670 97.830 106.810 ;
        RECT 92.125 106.625 92.415 106.670 ;
        RECT 95.705 106.625 95.995 106.670 ;
        RECT 97.540 106.625 97.830 106.670 ;
        RECT 98.005 106.625 98.295 106.855 ;
        RECT 99.370 106.810 99.690 106.870 ;
        RECT 98.770 106.670 99.690 106.810 ;
        RECT 27.625 106.470 27.915 106.515 ;
        RECT 30.370 106.470 30.690 106.530 ;
        RECT 35.430 106.470 35.750 106.530 ;
        RECT 36.825 106.470 37.115 106.515 ;
        RECT 27.625 106.330 37.115 106.470 ;
        RECT 27.625 106.285 27.915 106.330 ;
        RECT 30.370 106.270 30.690 106.330 ;
        RECT 35.430 106.270 35.750 106.330 ;
        RECT 36.825 106.285 37.115 106.330 ;
        RECT 38.650 106.270 38.970 106.530 ;
        RECT 48.325 106.470 48.615 106.515 ;
        RECT 50.150 106.470 50.470 106.530 ;
        RECT 48.325 106.330 50.470 106.470 ;
        RECT 48.325 106.285 48.615 106.330 ;
        RECT 50.150 106.270 50.470 106.330 ;
        RECT 72.245 106.470 72.535 106.515 ;
        RECT 75.910 106.470 76.230 106.530 ;
        RECT 82.365 106.470 82.655 106.515 ;
        RECT 72.245 106.330 82.655 106.470 ;
        RECT 85.200 106.470 85.340 106.625 ;
        RECT 89.710 106.470 90.030 106.530 ;
        RECT 98.770 106.470 98.910 106.670 ;
        RECT 99.370 106.610 99.690 106.670 ;
        RECT 101.625 106.650 101.915 106.965 ;
        RECT 103.510 106.950 103.830 107.010 ;
        RECT 104.565 106.965 105.215 107.010 ;
        RECT 105.810 107.150 106.130 107.210 ;
        RECT 107.205 107.150 107.495 107.195 ;
        RECT 105.810 107.010 107.495 107.150 ;
        RECT 105.810 106.950 106.130 107.010 ;
        RECT 107.205 106.965 107.495 107.010 ;
        RECT 111.880 107.010 115.240 107.150 ;
        RECT 111.880 106.870 112.020 107.010 ;
        RECT 102.705 106.810 102.995 106.855 ;
        RECT 106.285 106.810 106.575 106.855 ;
        RECT 108.120 106.810 108.410 106.855 ;
        RECT 102.705 106.670 108.410 106.810 ;
        RECT 102.705 106.625 102.995 106.670 ;
        RECT 106.285 106.625 106.575 106.670 ;
        RECT 108.120 106.625 108.410 106.670 ;
        RECT 109.045 106.810 109.335 106.855 ;
        RECT 110.410 106.810 110.730 106.870 ;
        RECT 109.045 106.670 110.730 106.810 ;
        RECT 109.045 106.625 109.335 106.670 ;
        RECT 110.410 106.610 110.730 106.670 ;
        RECT 111.790 106.610 112.110 106.870 ;
        RECT 112.710 106.810 113.030 106.870 ;
        RECT 115.100 106.855 115.240 107.010 ;
        RECT 118.690 106.950 119.010 107.210 ;
        RECT 120.990 107.195 121.310 107.210 ;
        RECT 120.985 107.150 121.635 107.195 ;
        RECT 124.585 107.150 124.875 107.195 ;
        RECT 120.985 107.010 124.875 107.150 ;
        RECT 120.985 106.965 121.635 107.010 ;
        RECT 124.285 106.965 124.875 107.010 ;
        RECT 120.990 106.950 121.310 106.965 ;
        RECT 113.185 106.810 113.475 106.855 ;
        RECT 112.710 106.670 113.475 106.810 ;
        RECT 112.710 106.610 113.030 106.670 ;
        RECT 113.185 106.625 113.475 106.670 ;
        RECT 115.025 106.625 115.315 106.855 ;
        RECT 117.790 106.810 118.080 106.855 ;
        RECT 119.625 106.810 119.915 106.855 ;
        RECT 123.205 106.810 123.495 106.855 ;
        RECT 117.790 106.670 123.495 106.810 ;
        RECT 117.790 106.625 118.080 106.670 ;
        RECT 119.625 106.625 119.915 106.670 ;
        RECT 123.205 106.625 123.495 106.670 ;
        RECT 124.285 106.650 124.575 106.965 ;
        RECT 135.660 106.690 136.800 133.400 ;
        RECT 133.100 106.600 136.850 106.690 ;
        RECT 85.200 106.330 98.910 106.470 ;
        RECT 108.585 106.470 108.875 106.515 ;
        RECT 109.490 106.470 109.810 106.530 ;
        RECT 112.250 106.470 112.570 106.530 ;
        RECT 117.325 106.470 117.615 106.515 ;
        RECT 124.670 106.470 124.990 106.530 ;
        RECT 126.050 106.470 126.370 106.530 ;
        RECT 108.585 106.330 126.370 106.470 ;
        RECT 72.245 106.285 72.535 106.330 ;
        RECT 75.910 106.270 76.230 106.330 ;
        RECT 82.365 106.285 82.655 106.330 ;
        RECT 89.710 106.270 90.030 106.330 ;
        RECT 108.585 106.285 108.875 106.330 ;
        RECT 109.490 106.270 109.810 106.330 ;
        RECT 112.250 106.270 112.570 106.330 ;
        RECT 117.325 106.285 117.615 106.330 ;
        RECT 124.670 106.270 124.990 106.330 ;
        RECT 126.050 106.270 126.370 106.330 ;
        RECT 21.745 106.130 22.035 106.175 ;
        RECT 24.865 106.130 25.155 106.175 ;
        RECT 26.755 106.130 27.045 106.175 ;
        RECT 21.745 105.990 27.045 106.130 ;
        RECT 21.745 105.945 22.035 105.990 ;
        RECT 24.865 105.945 25.155 105.990 ;
        RECT 26.755 105.945 27.045 105.990 ;
        RECT 30.945 106.130 31.235 106.175 ;
        RECT 34.065 106.130 34.355 106.175 ;
        RECT 35.955 106.130 36.245 106.175 ;
        RECT 30.945 105.990 36.245 106.130 ;
        RECT 30.945 105.945 31.235 105.990 ;
        RECT 34.065 105.945 34.355 105.990 ;
        RECT 35.955 105.945 36.245 105.990 ;
        RECT 42.445 106.130 42.735 106.175 ;
        RECT 45.565 106.130 45.855 106.175 ;
        RECT 47.455 106.130 47.745 106.175 ;
        RECT 42.445 105.990 47.745 106.130 ;
        RECT 42.445 105.945 42.735 105.990 ;
        RECT 45.565 105.945 45.855 105.990 ;
        RECT 47.455 105.945 47.745 105.990 ;
        RECT 66.365 106.130 66.655 106.175 ;
        RECT 69.485 106.130 69.775 106.175 ;
        RECT 71.375 106.130 71.665 106.175 ;
        RECT 66.365 105.990 71.665 106.130 ;
        RECT 66.365 105.945 66.655 105.990 ;
        RECT 69.485 105.945 69.775 105.990 ;
        RECT 71.375 105.945 71.665 105.990 ;
        RECT 76.485 106.130 76.775 106.175 ;
        RECT 79.605 106.130 79.895 106.175 ;
        RECT 81.495 106.130 81.785 106.175 ;
        RECT 76.485 105.990 81.785 106.130 ;
        RECT 76.485 105.945 76.775 105.990 ;
        RECT 79.605 105.945 79.895 105.990 ;
        RECT 81.495 105.945 81.785 105.990 ;
        RECT 92.125 106.130 92.415 106.175 ;
        RECT 95.245 106.130 95.535 106.175 ;
        RECT 97.135 106.130 97.425 106.175 ;
        RECT 92.125 105.990 97.425 106.130 ;
        RECT 92.125 105.945 92.415 105.990 ;
        RECT 95.245 105.945 95.535 105.990 ;
        RECT 97.135 105.945 97.425 105.990 ;
        RECT 102.705 106.130 102.995 106.175 ;
        RECT 105.825 106.130 106.115 106.175 ;
        RECT 107.715 106.130 108.005 106.175 ;
        RECT 102.705 105.990 108.005 106.130 ;
        RECT 102.705 105.945 102.995 105.990 ;
        RECT 105.825 105.945 106.115 105.990 ;
        RECT 107.715 105.945 108.005 105.990 ;
        RECT 118.195 106.130 118.485 106.175 ;
        RECT 120.085 106.130 120.375 106.175 ;
        RECT 123.205 106.130 123.495 106.175 ;
        RECT 118.195 105.990 123.495 106.130 ;
        RECT 118.195 105.945 118.485 105.990 ;
        RECT 120.085 105.945 120.375 105.990 ;
        RECT 123.205 105.945 123.495 105.990 ;
        RECT 17.950 105.590 18.270 105.850 ;
        RECT 18.885 105.790 19.175 105.835 ;
        RECT 26.230 105.790 26.550 105.850 ;
        RECT 18.885 105.650 26.550 105.790 ;
        RECT 18.885 105.605 19.175 105.650 ;
        RECT 26.230 105.590 26.550 105.650 ;
        RECT 28.085 105.790 28.375 105.835 ;
        RECT 30.370 105.790 30.690 105.850 ;
        RECT 28.085 105.650 30.690 105.790 ;
        RECT 28.085 105.605 28.375 105.650 ;
        RECT 30.370 105.590 30.690 105.650 ;
        RECT 39.585 105.790 39.875 105.835 ;
        RECT 44.170 105.790 44.490 105.850 ;
        RECT 39.585 105.650 44.490 105.790 ;
        RECT 39.585 105.605 39.875 105.650 ;
        RECT 44.170 105.590 44.490 105.650 ;
        RECT 52.450 105.790 52.770 105.850 ;
        RECT 53.845 105.790 54.135 105.835 ;
        RECT 52.450 105.650 54.135 105.790 ;
        RECT 52.450 105.590 52.770 105.650 ;
        RECT 53.845 105.605 54.135 105.650 ;
        RECT 56.145 105.790 56.435 105.835 ;
        RECT 57.510 105.790 57.830 105.850 ;
        RECT 56.145 105.650 57.830 105.790 ;
        RECT 56.145 105.605 56.435 105.650 ;
        RECT 57.510 105.590 57.830 105.650 ;
        RECT 61.190 105.790 61.510 105.850 ;
        RECT 62.125 105.790 62.415 105.835 ;
        RECT 61.190 105.650 62.415 105.790 ;
        RECT 61.190 105.590 61.510 105.650 ;
        RECT 62.125 105.605 62.415 105.650 ;
        RECT 63.505 105.790 63.795 105.835 ;
        RECT 68.090 105.790 68.410 105.850 ;
        RECT 63.505 105.650 68.410 105.790 ;
        RECT 63.505 105.605 63.795 105.650 ;
        RECT 68.090 105.590 68.410 105.650 ;
        RECT 73.625 105.790 73.915 105.835 ;
        RECT 74.070 105.790 74.390 105.850 ;
        RECT 73.625 105.650 74.390 105.790 ;
        RECT 73.625 105.605 73.915 105.650 ;
        RECT 74.070 105.590 74.390 105.650 ;
        RECT 83.730 105.590 84.050 105.850 ;
        RECT 84.190 105.790 84.510 105.850 ;
        RECT 84.665 105.790 84.955 105.835 ;
        RECT 84.190 105.650 84.955 105.790 ;
        RECT 84.190 105.590 84.510 105.650 ;
        RECT 84.665 105.605 84.955 105.650 ;
        RECT 87.425 105.790 87.715 105.835 ;
        RECT 87.870 105.790 88.190 105.850 ;
        RECT 87.425 105.650 88.190 105.790 ;
        RECT 87.425 105.605 87.715 105.650 ;
        RECT 87.870 105.590 88.190 105.650 ;
        RECT 89.265 105.790 89.555 105.835 ;
        RECT 93.850 105.790 94.170 105.850 ;
        RECT 89.265 105.650 94.170 105.790 ;
        RECT 89.265 105.605 89.555 105.650 ;
        RECT 93.850 105.590 94.170 105.650 ;
        RECT 99.845 105.790 100.135 105.835 ;
        RECT 103.970 105.790 104.290 105.850 ;
        RECT 99.845 105.650 104.290 105.790 ;
        RECT 99.845 105.605 100.135 105.650 ;
        RECT 103.970 105.590 104.290 105.650 ;
        RECT 109.965 105.790 110.255 105.835 ;
        RECT 111.790 105.790 112.110 105.850 ;
        RECT 109.965 105.650 112.110 105.790 ;
        RECT 109.965 105.605 110.255 105.650 ;
        RECT 111.790 105.590 112.110 105.650 ;
        RECT 114.090 105.590 114.410 105.850 ;
        RECT 115.470 105.590 115.790 105.850 ;
        RECT 126.065 105.790 126.355 105.835 ;
        RECT 127.890 105.790 128.210 105.850 ;
        RECT 126.065 105.650 128.210 105.790 ;
        RECT 126.065 105.605 126.355 105.650 ;
        RECT 127.890 105.590 128.210 105.650 ;
        RECT 129.700 105.630 136.850 106.600 ;
        RECT 133.100 105.500 136.850 105.630 ;
        RECT 14.660 104.970 127.820 105.450 ;
        RECT 38.665 104.770 38.955 104.815 ;
        RECT 39.110 104.770 39.430 104.830 ;
        RECT 38.665 104.630 39.430 104.770 ;
        RECT 38.665 104.585 38.955 104.630 ;
        RECT 39.110 104.570 39.430 104.630 ;
        RECT 50.150 104.770 50.470 104.830 ;
        RECT 63.950 104.770 64.270 104.830 ;
        RECT 50.150 104.630 57.740 104.770 ;
        RECT 50.150 104.570 50.470 104.630 ;
        RECT 27.725 104.430 28.015 104.475 ;
        RECT 30.845 104.430 31.135 104.475 ;
        RECT 32.735 104.430 33.025 104.475 ;
        RECT 27.725 104.290 33.025 104.430 ;
        RECT 27.725 104.245 28.015 104.290 ;
        RECT 30.845 104.245 31.135 104.290 ;
        RECT 32.735 104.245 33.025 104.290 ;
        RECT 41.835 104.430 42.125 104.475 ;
        RECT 43.725 104.430 44.015 104.475 ;
        RECT 46.845 104.430 47.135 104.475 ;
        RECT 41.835 104.290 47.135 104.430 ;
        RECT 41.835 104.245 42.125 104.290 ;
        RECT 43.725 104.245 44.015 104.290 ;
        RECT 46.845 104.245 47.135 104.290 ;
        RECT 28.530 104.090 28.850 104.150 ;
        RECT 32.225 104.090 32.515 104.135 ;
        RECT 28.530 103.950 32.515 104.090 ;
        RECT 28.530 103.890 28.850 103.950 ;
        RECT 32.225 103.905 32.515 103.950 ;
        RECT 33.605 104.090 33.895 104.135 ;
        RECT 35.430 104.090 35.750 104.150 ;
        RECT 40.965 104.090 41.255 104.135 ;
        RECT 33.605 103.950 41.255 104.090 ;
        RECT 33.605 103.905 33.895 103.950 ;
        RECT 35.430 103.890 35.750 103.950 ;
        RECT 40.965 103.905 41.255 103.950 ;
        RECT 42.330 103.890 42.650 104.150 ;
        RECT 51.160 104.135 51.300 104.630 ;
        RECT 51.955 104.430 52.245 104.475 ;
        RECT 53.845 104.430 54.135 104.475 ;
        RECT 56.965 104.430 57.255 104.475 ;
        RECT 51.955 104.290 57.255 104.430 ;
        RECT 57.600 104.430 57.740 104.630 ;
        RECT 60.820 104.630 69.240 104.770 ;
        RECT 60.820 104.430 60.960 104.630 ;
        RECT 63.950 104.570 64.270 104.630 ;
        RECT 57.600 104.290 60.960 104.430 ;
        RECT 63.145 104.430 63.435 104.475 ;
        RECT 66.265 104.430 66.555 104.475 ;
        RECT 68.155 104.430 68.445 104.475 ;
        RECT 63.145 104.290 68.445 104.430 ;
        RECT 51.955 104.245 52.245 104.290 ;
        RECT 53.845 104.245 54.135 104.290 ;
        RECT 56.965 104.245 57.255 104.290 ;
        RECT 63.145 104.245 63.435 104.290 ;
        RECT 66.265 104.245 66.555 104.290 ;
        RECT 68.155 104.245 68.445 104.290 ;
        RECT 51.085 103.905 51.375 104.135 ;
        RECT 52.450 103.890 52.770 104.150 ;
        RECT 52.910 104.090 53.230 104.150 ;
        RECT 69.100 104.135 69.240 104.630 ;
        RECT 85.200 104.630 94.540 104.770 ;
        RECT 79.245 104.430 79.535 104.475 ;
        RECT 82.365 104.430 82.655 104.475 ;
        RECT 84.255 104.430 84.545 104.475 ;
        RECT 79.245 104.290 84.545 104.430 ;
        RECT 79.245 104.245 79.535 104.290 ;
        RECT 82.365 104.245 82.655 104.290 ;
        RECT 84.255 104.245 84.545 104.290 ;
        RECT 67.645 104.090 67.935 104.135 ;
        RECT 52.910 103.950 67.935 104.090 ;
        RECT 52.910 103.890 53.230 103.950 ;
        RECT 67.645 103.905 67.935 103.950 ;
        RECT 69.025 103.905 69.315 104.135 ;
        RECT 83.730 103.890 84.050 104.150 ;
        RECT 85.200 104.135 85.340 104.630 ;
        RECT 88.445 104.430 88.735 104.475 ;
        RECT 91.565 104.430 91.855 104.475 ;
        RECT 93.455 104.430 93.745 104.475 ;
        RECT 88.445 104.290 93.745 104.430 ;
        RECT 88.445 104.245 88.735 104.290 ;
        RECT 91.565 104.245 91.855 104.290 ;
        RECT 93.455 104.245 93.745 104.290 ;
        RECT 85.125 103.905 85.415 104.135 ;
        RECT 87.870 104.090 88.190 104.150 ;
        RECT 94.400 104.135 94.540 104.630 ;
        RECT 112.710 104.570 113.030 104.830 ;
        RECT 107.305 104.430 107.595 104.475 ;
        RECT 110.425 104.430 110.715 104.475 ;
        RECT 112.315 104.430 112.605 104.475 ;
        RECT 107.305 104.290 112.605 104.430 ;
        RECT 107.305 104.245 107.595 104.290 ;
        RECT 110.425 104.245 110.715 104.290 ;
        RECT 112.315 104.245 112.605 104.290 ;
        RECT 92.945 104.090 93.235 104.135 ;
        RECT 87.870 103.950 93.235 104.090 ;
        RECT 87.870 103.890 88.190 103.950 ;
        RECT 92.945 103.905 93.235 103.950 ;
        RECT 94.325 104.090 94.615 104.135 ;
        RECT 97.070 104.090 97.390 104.150 ;
        RECT 94.325 103.950 97.390 104.090 ;
        RECT 94.325 103.905 94.615 103.950 ;
        RECT 97.070 103.890 97.390 103.950 ;
        RECT 111.790 103.890 112.110 104.150 ;
        RECT 112.800 104.090 112.940 104.570 ;
        RECT 116.505 104.430 116.795 104.475 ;
        RECT 119.625 104.430 119.915 104.475 ;
        RECT 121.515 104.430 121.805 104.475 ;
        RECT 116.505 104.290 121.805 104.430 ;
        RECT 116.505 104.245 116.795 104.290 ;
        RECT 119.625 104.245 119.915 104.290 ;
        RECT 121.515 104.245 121.805 104.290 ;
        RECT 113.185 104.090 113.475 104.135 ;
        RECT 112.800 103.950 113.475 104.090 ;
        RECT 113.185 103.905 113.475 103.950 ;
        RECT 114.090 104.090 114.410 104.150 ;
        RECT 121.005 104.090 121.295 104.135 ;
        RECT 114.090 103.950 121.295 104.090 ;
        RECT 114.090 103.890 114.410 103.950 ;
        RECT 121.005 103.905 121.295 103.950 ;
        RECT 122.385 104.090 122.675 104.135 ;
        RECT 124.670 104.090 124.990 104.150 ;
        RECT 122.385 103.950 124.990 104.090 ;
        RECT 122.385 103.905 122.675 103.950 ;
        RECT 124.670 103.890 124.990 103.950 ;
        RECT 17.950 103.410 18.270 103.470 ;
        RECT 26.645 103.455 26.935 103.770 ;
        RECT 27.725 103.750 28.015 103.795 ;
        RECT 31.305 103.750 31.595 103.795 ;
        RECT 33.140 103.750 33.430 103.795 ;
        RECT 27.725 103.610 33.430 103.750 ;
        RECT 27.725 103.565 28.015 103.610 ;
        RECT 31.305 103.565 31.595 103.610 ;
        RECT 33.140 103.565 33.430 103.610 ;
        RECT 38.650 103.750 38.970 103.810 ;
        RECT 39.125 103.750 39.415 103.795 ;
        RECT 38.650 103.610 39.415 103.750 ;
        RECT 38.650 103.550 38.970 103.610 ;
        RECT 39.125 103.565 39.415 103.610 ;
        RECT 41.430 103.750 41.720 103.795 ;
        RECT 43.265 103.750 43.555 103.795 ;
        RECT 46.845 103.750 47.135 103.795 ;
        RECT 41.430 103.610 47.135 103.750 ;
        RECT 41.430 103.565 41.720 103.610 ;
        RECT 43.265 103.565 43.555 103.610 ;
        RECT 46.845 103.565 47.135 103.610 ;
        RECT 26.345 103.410 26.935 103.455 ;
        RECT 29.585 103.410 30.235 103.455 ;
        RECT 17.950 103.270 30.235 103.410 ;
        RECT 17.950 103.210 18.270 103.270 ;
        RECT 26.345 103.225 26.635 103.270 ;
        RECT 29.585 103.225 30.235 103.270 ;
        RECT 14.270 103.070 14.590 103.130 ;
        RECT 24.865 103.070 25.155 103.115 ;
        RECT 14.270 102.930 25.155 103.070 ;
        RECT 39.200 103.070 39.340 103.565 ;
        RECT 44.625 103.410 45.275 103.455 ;
        RECT 46.010 103.410 46.330 103.470 ;
        RECT 47.925 103.455 48.215 103.770 ;
        RECT 51.550 103.750 51.840 103.795 ;
        RECT 53.385 103.750 53.675 103.795 ;
        RECT 56.965 103.750 57.255 103.795 ;
        RECT 51.550 103.610 57.255 103.750 ;
        RECT 51.550 103.565 51.840 103.610 ;
        RECT 53.385 103.565 53.675 103.610 ;
        RECT 56.965 103.565 57.255 103.610 ;
        RECT 47.925 103.410 48.515 103.455 ;
        RECT 44.625 103.270 48.515 103.410 ;
        RECT 44.625 103.225 45.275 103.270 ;
        RECT 46.010 103.210 46.330 103.270 ;
        RECT 48.225 103.225 48.515 103.270 ;
        RECT 54.745 103.410 55.395 103.455 ;
        RECT 57.510 103.410 57.830 103.470 ;
        RECT 58.045 103.455 58.335 103.770 ;
        RECT 58.045 103.410 58.635 103.455 ;
        RECT 54.745 103.270 58.635 103.410 ;
        RECT 54.745 103.225 55.395 103.270 ;
        RECT 57.510 103.210 57.830 103.270 ;
        RECT 58.345 103.225 58.635 103.270 ;
        RECT 61.190 103.410 61.510 103.470 ;
        RECT 62.065 103.455 62.355 103.770 ;
        RECT 63.145 103.750 63.435 103.795 ;
        RECT 66.725 103.750 67.015 103.795 ;
        RECT 68.560 103.750 68.850 103.795 ;
        RECT 63.145 103.610 68.850 103.750 ;
        RECT 63.145 103.565 63.435 103.610 ;
        RECT 66.725 103.565 67.015 103.610 ;
        RECT 68.560 103.565 68.850 103.610 ;
        RECT 78.165 103.455 78.455 103.770 ;
        RECT 79.245 103.750 79.535 103.795 ;
        RECT 82.825 103.750 83.115 103.795 ;
        RECT 84.660 103.750 84.950 103.795 ;
        RECT 87.410 103.770 87.730 103.810 ;
        RECT 79.245 103.610 84.950 103.750 ;
        RECT 79.245 103.565 79.535 103.610 ;
        RECT 82.825 103.565 83.115 103.610 ;
        RECT 84.660 103.565 84.950 103.610 ;
        RECT 87.365 103.550 87.730 103.770 ;
        RECT 88.445 103.750 88.735 103.795 ;
        RECT 92.025 103.750 92.315 103.795 ;
        RECT 93.860 103.750 94.150 103.795 ;
        RECT 106.270 103.770 106.590 103.810 ;
        RECT 88.445 103.610 94.150 103.750 ;
        RECT 88.445 103.565 88.735 103.610 ;
        RECT 92.025 103.565 92.315 103.610 ;
        RECT 93.860 103.565 94.150 103.610 ;
        RECT 106.225 103.550 106.590 103.770 ;
        RECT 107.305 103.750 107.595 103.795 ;
        RECT 110.885 103.750 111.175 103.795 ;
        RECT 112.720 103.750 113.010 103.795 ;
        RECT 115.470 103.770 115.790 103.810 ;
        RECT 107.305 103.610 113.010 103.750 ;
        RECT 107.305 103.565 107.595 103.610 ;
        RECT 110.885 103.565 111.175 103.610 ;
        RECT 112.720 103.565 113.010 103.610 ;
        RECT 115.425 103.550 115.790 103.770 ;
        RECT 116.505 103.750 116.795 103.795 ;
        RECT 120.085 103.750 120.375 103.795 ;
        RECT 121.920 103.750 122.210 103.795 ;
        RECT 116.505 103.610 122.210 103.750 ;
        RECT 116.505 103.565 116.795 103.610 ;
        RECT 120.085 103.565 120.375 103.610 ;
        RECT 121.920 103.565 122.210 103.610 ;
        RECT 126.065 103.750 126.355 103.795 ;
        RECT 126.510 103.750 126.830 103.810 ;
        RECT 126.065 103.610 126.830 103.750 ;
        RECT 126.065 103.565 126.355 103.610 ;
        RECT 126.510 103.550 126.830 103.610 ;
        RECT 61.765 103.410 62.355 103.455 ;
        RECT 65.005 103.410 65.655 103.455 ;
        RECT 61.190 103.270 65.655 103.410 ;
        RECT 61.190 103.210 61.510 103.270 ;
        RECT 61.765 103.225 62.055 103.270 ;
        RECT 65.005 103.225 65.655 103.270 ;
        RECT 77.865 103.410 78.455 103.455 ;
        RECT 81.105 103.410 81.755 103.455 ;
        RECT 84.190 103.410 84.510 103.470 ;
        RECT 87.365 103.455 87.655 103.550 ;
        RECT 106.225 103.455 106.515 103.550 ;
        RECT 115.425 103.455 115.715 103.550 ;
        RECT 77.865 103.270 84.510 103.410 ;
        RECT 77.865 103.225 78.155 103.270 ;
        RECT 81.105 103.225 81.755 103.270 ;
        RECT 84.190 103.210 84.510 103.270 ;
        RECT 87.065 103.410 87.655 103.455 ;
        RECT 90.305 103.410 90.955 103.455 ;
        RECT 87.065 103.270 90.955 103.410 ;
        RECT 87.065 103.225 87.355 103.270 ;
        RECT 90.305 103.225 90.955 103.270 ;
        RECT 105.925 103.410 106.515 103.455 ;
        RECT 109.165 103.410 109.815 103.455 ;
        RECT 105.925 103.270 109.815 103.410 ;
        RECT 105.925 103.225 106.215 103.270 ;
        RECT 109.165 103.225 109.815 103.270 ;
        RECT 115.125 103.410 115.715 103.455 ;
        RECT 118.365 103.410 119.015 103.455 ;
        RECT 115.125 103.270 119.015 103.410 ;
        RECT 115.125 103.225 115.415 103.270 ;
        RECT 118.365 103.225 119.015 103.270 ;
        RECT 49.230 103.070 49.550 103.130 ;
        RECT 39.200 102.930 49.550 103.070 ;
        RECT 14.270 102.870 14.590 102.930 ;
        RECT 24.865 102.885 25.155 102.930 ;
        RECT 49.230 102.870 49.550 102.930 ;
        RECT 49.690 102.870 50.010 103.130 ;
        RECT 56.130 103.070 56.450 103.130 ;
        RECT 59.825 103.070 60.115 103.115 ;
        RECT 56.130 102.930 60.115 103.070 ;
        RECT 56.130 102.870 56.450 102.930 ;
        RECT 59.825 102.885 60.115 102.930 ;
        RECT 60.285 103.070 60.575 103.115 ;
        RECT 60.730 103.070 61.050 103.130 ;
        RECT 60.285 102.930 61.050 103.070 ;
        RECT 60.285 102.885 60.575 102.930 ;
        RECT 60.730 102.870 61.050 102.930 ;
        RECT 76.385 103.070 76.675 103.115 ;
        RECT 80.050 103.070 80.370 103.130 ;
        RECT 76.385 102.930 80.370 103.070 ;
        RECT 76.385 102.885 76.675 102.930 ;
        RECT 80.050 102.870 80.370 102.930 ;
        RECT 85.570 102.870 85.890 103.130 ;
        RECT 104.445 103.070 104.735 103.115 ;
        RECT 109.950 103.070 110.270 103.130 ;
        RECT 104.445 102.930 110.270 103.070 ;
        RECT 104.445 102.885 104.735 102.930 ;
        RECT 109.950 102.870 110.270 102.930 ;
        RECT 113.645 103.070 113.935 103.115 ;
        RECT 115.930 103.070 116.250 103.130 ;
        RECT 113.645 102.930 116.250 103.070 ;
        RECT 113.645 102.885 113.935 102.930 ;
        RECT 115.930 102.870 116.250 102.930 ;
        RECT 125.130 102.870 125.450 103.130 ;
        RECT 14.660 102.250 127.820 102.730 ;
        RECT 46.010 102.050 46.330 102.110 ;
        RECT 47.405 102.050 47.695 102.095 ;
        RECT 46.010 101.910 47.695 102.050 ;
        RECT 46.010 101.850 46.330 101.910 ;
        RECT 47.405 101.865 47.695 101.910 ;
        RECT 64.885 102.050 65.175 102.095 ;
        RECT 65.330 102.050 65.650 102.110 ;
        RECT 64.885 101.910 65.650 102.050 ;
        RECT 64.885 101.865 65.175 101.910 ;
        RECT 65.330 101.850 65.650 101.910 ;
        RECT 76.370 102.050 76.690 102.110 ;
        RECT 125.130 102.050 125.450 102.110 ;
        RECT 76.370 101.910 125.450 102.050 ;
        RECT 76.370 101.850 76.690 101.910 ;
        RECT 125.130 101.850 125.450 101.910 ;
        RECT 47.865 101.370 48.155 101.415 ;
        RECT 49.230 101.370 49.550 101.430 ;
        RECT 55.670 101.370 55.990 101.430 ;
        RECT 64.425 101.370 64.715 101.415 ;
        RECT 47.865 101.230 64.715 101.370 ;
        RECT 47.865 101.185 48.155 101.230 ;
        RECT 49.230 101.170 49.550 101.230 ;
        RECT 55.670 101.170 55.990 101.230 ;
        RECT 64.425 101.185 64.715 101.230 ;
        RECT 14.660 99.530 127.820 100.010 ;
        RECT 133.330 76.630 136.060 77.830 ;
        RECT 137.920 77.810 143.450 77.960 ;
        RECT 21.115 74.380 23.065 74.390 ;
        RECT 19.415 73.240 23.065 74.380 ;
        RECT 19.415 73.230 21.125 73.240 ;
        RECT 28.135 73.230 30.305 74.410 ;
        RECT 32.315 74.390 34.265 74.400 ;
        RECT 30.615 73.250 34.265 74.390 ;
        RECT 30.615 73.240 32.325 73.250 ;
        RECT 39.425 73.200 41.595 74.380 ;
        RECT 43.535 74.360 45.485 74.370 ;
        RECT 41.835 73.220 45.485 74.360 ;
        RECT 54.785 74.340 56.735 74.350 ;
        RECT 41.835 73.210 43.545 73.220 ;
        RECT 3.910 73.080 6.100 73.190 ;
        RECT 50.005 73.140 52.175 74.320 ;
        RECT 53.085 73.200 56.735 74.340 ;
        RECT 53.085 73.190 54.795 73.200 ;
        RECT 61.425 73.170 63.595 74.350 ;
        RECT 66.005 74.330 67.955 74.340 ;
        RECT 64.305 73.190 67.955 74.330 ;
        RECT 64.305 73.180 66.015 73.190 ;
        RECT 72.535 73.180 74.705 74.360 ;
        RECT 77.245 74.320 79.195 74.330 ;
        RECT 75.545 73.180 79.195 74.320 ;
        RECT 75.545 73.170 77.255 73.180 ;
        RECT 83.805 73.170 85.975 74.350 ;
        RECT 88.495 74.330 90.445 74.340 ;
        RECT 86.795 73.190 90.445 74.330 ;
        RECT 99.775 74.320 101.725 74.330 ;
        RECT 86.795 73.180 88.505 73.190 ;
        RECT 94.995 73.110 97.165 74.290 ;
        RECT 98.075 73.180 101.725 74.320 ;
        RECT 98.075 73.170 99.785 73.180 ;
        RECT 106.405 73.160 108.575 74.340 ;
        RECT 111.045 74.320 112.995 74.330 ;
        RECT 109.345 73.180 112.995 74.320 ;
        RECT 109.345 73.170 111.055 73.180 ;
        RECT 117.605 73.160 119.775 74.340 ;
        RECT 122.295 74.320 124.245 74.330 ;
        RECT 120.595 73.180 124.245 74.320 ;
        RECT 129.455 73.240 131.625 74.420 ;
        RECT 120.595 73.170 122.305 73.180 ;
        RECT 3.910 72.820 12.240 73.080 ;
        RECT 29.635 72.840 43.235 72.850 ;
        RECT 18.435 72.820 43.235 72.840 ;
        RECT 3.910 72.800 54.455 72.820 ;
        RECT 3.910 72.790 65.705 72.800 ;
        RECT 133.960 72.790 135.640 76.630 ;
        RECT 137.190 76.610 143.450 77.810 ;
        RECT 137.920 75.460 143.450 76.610 ;
        RECT 3.910 72.780 76.925 72.790 ;
        RECT 85.815 72.780 99.415 72.790 ;
        RECT 132.085 72.780 140.600 72.790 ;
        RECT 3.910 71.700 140.600 72.780 ;
        RECT 3.910 71.690 32.035 71.700 ;
        RECT 3.910 71.670 19.135 71.690 ;
        RECT 40.855 71.670 140.600 71.700 ;
        RECT 3.910 71.500 12.240 71.670 ;
        RECT 52.105 71.650 140.600 71.670 ;
        RECT 63.325 71.640 140.600 71.650 ;
        RECT 74.565 71.630 88.165 71.640 ;
        RECT 97.095 71.630 133.215 71.640 ;
        RECT 3.910 71.370 6.100 71.500 ;
        RECT 10.800 71.180 11.950 71.500 ;
        RECT 10.800 69.480 11.915 71.180 ;
        RECT 29.635 71.170 43.285 71.180 ;
        RECT 15.510 71.155 17.040 71.160 ;
        RECT 18.435 71.155 43.285 71.170 ;
        RECT 12.285 71.150 43.285 71.155 ;
        RECT 12.285 71.130 54.505 71.150 ;
        RECT 141.810 71.140 143.230 75.460 ;
        RECT 12.285 71.120 65.755 71.130 ;
        RECT 12.285 71.110 76.975 71.120 ;
        RECT 85.815 71.110 99.465 71.120 ;
        RECT 140.220 71.110 143.240 71.140 ;
        RECT 12.285 70.030 143.240 71.110 ;
        RECT 12.285 70.020 32.085 70.030 ;
        RECT 12.285 70.005 19.375 70.020 ;
        RECT 10.800 13.800 11.950 69.480 ;
        RECT 12.320 15.450 13.470 70.005 ;
        RECT 15.510 68.660 17.040 70.005 ;
        RECT 40.855 70.000 143.240 70.030 ;
        RECT 52.105 69.980 143.240 70.000 ;
        RECT 63.325 69.970 143.240 69.980 ;
        RECT 74.565 69.960 88.215 69.970 ;
        RECT 97.095 69.960 143.240 69.970 ;
        RECT 140.220 69.910 143.240 69.960 ;
        RECT 29.645 69.670 43.315 69.680 ;
        RECT 18.445 69.650 43.315 69.670 ;
        RECT 18.445 69.630 54.535 69.650 ;
        RECT 18.445 69.620 65.785 69.630 ;
        RECT 139.590 69.620 150.610 69.640 ;
        RECT 18.445 69.610 77.005 69.620 ;
        RECT 85.825 69.610 99.495 69.620 ;
        RECT 132.155 69.610 150.610 69.620 ;
        RECT 18.445 69.570 150.610 69.610 ;
        RECT 18.445 68.530 150.740 69.570 ;
        RECT 18.445 68.520 32.115 68.530 ;
        RECT 40.865 68.500 150.740 68.530 ;
        RECT 52.115 68.490 143.320 68.500 ;
        RECT 52.115 68.480 140.670 68.490 ;
        RECT 63.335 68.470 140.670 68.480 ;
        RECT 74.575 68.460 88.245 68.470 ;
        RECT 97.105 68.460 133.295 68.470 ;
        RECT 141.080 68.450 142.300 68.490 ;
        RECT 149.360 68.470 150.740 68.500 ;
        RECT 29.655 68.100 43.325 68.110 ;
        RECT 13.950 68.080 43.325 68.100 ;
        RECT 13.950 68.060 54.545 68.080 ;
        RECT 13.950 68.050 65.795 68.060 ;
        RECT 13.950 68.040 77.015 68.050 ;
        RECT 85.835 68.040 99.505 68.050 ;
        RECT 139.530 68.040 143.320 68.060 ;
        RECT 13.950 66.960 152.870 68.040 ;
        RECT 13.950 66.950 32.125 66.960 ;
        RECT 13.950 18.530 15.100 66.950 ;
        RECT 40.875 66.930 152.870 66.960 ;
        RECT 52.125 66.910 152.870 66.930 ;
        RECT 63.345 66.900 152.870 66.910 ;
        RECT 74.585 66.890 88.255 66.900 ;
        RECT 97.115 66.890 143.320 66.900 ;
        RECT 141.030 66.770 142.490 66.890 ;
        RECT 21.405 65.510 26.555 65.790 ;
        RECT 27.815 65.490 28.965 65.800 ;
        RECT 32.605 65.520 37.755 65.800 ;
        RECT 39.015 65.500 40.165 65.810 ;
        RECT 43.825 65.490 48.975 65.770 ;
        RECT 50.235 65.470 51.385 65.780 ;
        RECT 149.460 65.760 150.600 65.780 ;
        RECT 55.075 65.470 60.225 65.750 ;
        RECT 61.485 65.450 62.635 65.760 ;
        RECT 66.295 65.460 71.445 65.740 ;
        RECT 72.705 65.440 73.855 65.750 ;
        RECT 77.535 65.450 82.685 65.730 ;
        RECT 83.945 65.430 85.095 65.740 ;
        RECT 88.785 65.460 93.935 65.740 ;
        RECT 95.195 65.440 96.345 65.750 ;
        RECT 100.065 65.450 105.215 65.730 ;
        RECT 106.475 65.430 107.625 65.740 ;
        RECT 111.335 65.450 116.485 65.730 ;
        RECT 117.745 65.430 118.895 65.740 ;
        RECT 122.585 65.450 127.735 65.730 ;
        RECT 128.995 65.430 130.145 65.740 ;
        RECT 133.315 65.430 138.455 65.690 ;
        RECT 21.205 65.140 21.435 65.320 ;
        RECT 26.495 65.190 26.725 65.320 ;
        RECT 21.125 55.220 21.485 65.140 ;
        RECT 26.435 55.240 26.805 65.190 ;
        RECT 27.635 65.150 27.865 65.320 ;
        RECT 27.565 55.200 27.935 65.150 ;
        RECT 28.925 65.140 29.155 65.320 ;
        RECT 32.405 65.150 32.635 65.330 ;
        RECT 37.695 65.200 37.925 65.330 ;
        RECT 28.835 55.250 29.255 65.140 ;
        RECT 32.325 55.230 32.685 65.150 ;
        RECT 37.635 55.250 38.005 65.200 ;
        RECT 38.835 65.160 39.065 65.330 ;
        RECT 38.765 55.210 39.135 65.160 ;
        RECT 40.125 65.150 40.355 65.330 ;
        RECT 40.035 55.260 40.455 65.150 ;
        RECT 43.625 65.120 43.855 65.300 ;
        RECT 48.915 65.170 49.145 65.300 ;
        RECT 43.545 55.200 43.905 65.120 ;
        RECT 48.855 55.220 49.225 65.170 ;
        RECT 50.055 65.130 50.285 65.300 ;
        RECT 49.985 55.180 50.355 65.130 ;
        RECT 51.345 65.120 51.575 65.300 ;
        RECT 51.255 55.230 51.675 65.120 ;
        RECT 54.875 65.100 55.105 65.280 ;
        RECT 60.165 65.150 60.395 65.280 ;
        RECT 54.795 55.180 55.155 65.100 ;
        RECT 60.105 55.200 60.475 65.150 ;
        RECT 61.305 65.110 61.535 65.280 ;
        RECT 61.235 55.160 61.605 65.110 ;
        RECT 62.595 65.100 62.825 65.280 ;
        RECT 62.505 55.210 62.925 65.100 ;
        RECT 66.095 65.090 66.325 65.270 ;
        RECT 71.385 65.140 71.615 65.270 ;
        RECT 66.015 55.170 66.375 65.090 ;
        RECT 71.325 55.190 71.695 65.140 ;
        RECT 72.525 65.100 72.755 65.270 ;
        RECT 72.455 55.150 72.825 65.100 ;
        RECT 73.815 65.090 74.045 65.270 ;
        RECT 73.725 55.200 74.145 65.090 ;
        RECT 77.335 65.080 77.565 65.260 ;
        RECT 82.625 65.130 82.855 65.260 ;
        RECT 77.255 55.160 77.615 65.080 ;
        RECT 82.565 55.180 82.935 65.130 ;
        RECT 83.765 65.090 83.995 65.260 ;
        RECT 83.695 55.140 84.065 65.090 ;
        RECT 85.055 65.080 85.285 65.260 ;
        RECT 88.585 65.090 88.815 65.270 ;
        RECT 93.875 65.140 94.105 65.270 ;
        RECT 84.965 55.190 85.385 65.080 ;
        RECT 88.505 55.170 88.865 65.090 ;
        RECT 93.815 55.190 94.185 65.140 ;
        RECT 95.015 65.100 95.245 65.270 ;
        RECT 94.945 55.150 95.315 65.100 ;
        RECT 96.305 65.090 96.535 65.270 ;
        RECT 96.215 55.200 96.635 65.090 ;
        RECT 99.865 65.080 100.095 65.260 ;
        RECT 105.155 65.130 105.385 65.260 ;
        RECT 99.785 55.160 100.145 65.080 ;
        RECT 105.095 55.180 105.465 65.130 ;
        RECT 106.295 65.090 106.525 65.260 ;
        RECT 106.225 55.140 106.595 65.090 ;
        RECT 107.585 65.080 107.815 65.260 ;
        RECT 111.135 65.080 111.365 65.260 ;
        RECT 116.425 65.130 116.655 65.260 ;
        RECT 107.495 55.190 107.915 65.080 ;
        RECT 111.055 55.160 111.415 65.080 ;
        RECT 116.365 55.180 116.735 65.130 ;
        RECT 117.565 65.090 117.795 65.260 ;
        RECT 117.495 55.140 117.865 65.090 ;
        RECT 118.855 65.080 119.085 65.260 ;
        RECT 122.385 65.080 122.615 65.260 ;
        RECT 127.675 65.130 127.905 65.260 ;
        RECT 118.765 55.190 119.185 65.080 ;
        RECT 122.305 55.160 122.665 65.080 ;
        RECT 127.615 55.180 127.985 65.130 ;
        RECT 128.815 65.090 129.045 65.260 ;
        RECT 128.745 55.140 129.115 65.090 ;
        RECT 130.105 65.080 130.335 65.260 ;
        RECT 133.135 65.130 133.365 65.230 ;
        RECT 130.015 55.190 130.435 65.080 ;
        RECT 133.005 55.240 133.405 65.130 ;
        RECT 138.425 65.100 138.655 65.230 ;
        RECT 133.135 55.230 133.365 55.240 ;
        RECT 138.345 55.130 138.725 65.100 ;
        RECT 149.340 64.660 150.720 65.760 ;
        RECT 20.815 54.230 25.555 54.530 ;
        RECT 32.015 54.240 36.755 54.540 ;
        RECT 43.235 54.210 47.975 54.510 ;
        RECT 54.485 54.190 59.225 54.490 ;
        RECT 65.705 54.180 70.445 54.480 ;
        RECT 76.945 54.170 81.685 54.470 ;
        RECT 88.195 54.180 92.935 54.480 ;
        RECT 99.475 54.170 104.215 54.470 ;
        RECT 110.745 54.170 115.485 54.470 ;
        RECT 121.995 54.170 126.735 54.470 ;
        RECT 21.655 52.320 22.115 52.550 ;
        RECT 25.625 52.280 26.255 52.560 ;
        RECT 25.735 52.240 26.195 52.280 ;
        RECT 27.665 52.240 28.125 52.470 ;
        RECT 32.855 52.330 33.315 52.560 ;
        RECT 36.825 52.290 37.455 52.570 ;
        RECT 36.935 52.250 37.395 52.290 ;
        RECT 38.865 52.250 39.325 52.480 ;
        RECT 44.075 52.300 44.535 52.530 ;
        RECT 48.045 52.260 48.675 52.540 ;
        RECT 48.155 52.220 48.615 52.260 ;
        RECT 50.085 52.220 50.545 52.450 ;
        RECT 55.325 52.280 55.785 52.510 ;
        RECT 59.295 52.240 59.925 52.520 ;
        RECT 59.405 52.200 59.865 52.240 ;
        RECT 61.335 52.200 61.795 52.430 ;
        RECT 66.545 52.270 67.005 52.500 ;
        RECT 70.515 52.230 71.145 52.510 ;
        RECT 70.625 52.190 71.085 52.230 ;
        RECT 72.555 52.190 73.015 52.420 ;
        RECT 77.785 52.260 78.245 52.490 ;
        RECT 81.755 52.220 82.385 52.500 ;
        RECT 81.865 52.180 82.325 52.220 ;
        RECT 83.795 52.180 84.255 52.410 ;
        RECT 89.035 52.270 89.495 52.500 ;
        RECT 93.005 52.230 93.635 52.510 ;
        RECT 93.115 52.190 93.575 52.230 ;
        RECT 95.045 52.190 95.505 52.420 ;
        RECT 100.315 52.260 100.775 52.490 ;
        RECT 104.285 52.220 104.915 52.500 ;
        RECT 104.395 52.180 104.855 52.220 ;
        RECT 106.325 52.180 106.785 52.410 ;
        RECT 111.585 52.260 112.045 52.490 ;
        RECT 115.555 52.220 116.185 52.500 ;
        RECT 115.665 52.180 116.125 52.220 ;
        RECT 117.595 52.180 118.055 52.410 ;
        RECT 122.835 52.260 123.295 52.490 ;
        RECT 126.805 52.220 127.435 52.500 ;
        RECT 126.915 52.180 127.375 52.220 ;
        RECT 128.845 52.180 129.305 52.410 ;
        RECT 21.375 52.010 21.605 52.115 ;
        RECT 21.245 50.290 21.615 52.010 ;
        RECT 22.165 51.890 22.395 52.115 ;
        RECT 25.455 51.980 25.685 52.035 ;
        RECT 21.375 50.115 21.605 50.290 ;
        RECT 22.155 50.210 22.525 51.890 ;
        RECT 22.165 50.115 22.395 50.210 ;
        RECT 21.525 49.670 22.245 49.930 ;
        RECT 19.295 46.650 20.065 47.720 ;
        RECT 21.385 47.490 22.105 47.750 ;
        RECT 21.225 47.200 21.455 47.340 ;
        RECT 21.085 46.430 21.475 47.200 ;
        RECT 22.015 47.190 22.245 47.340 ;
        RECT 22.005 46.450 22.375 47.190 ;
        RECT 25.305 47.010 25.735 51.980 ;
        RECT 26.245 51.970 26.475 52.035 ;
        RECT 27.385 51.970 27.615 52.035 ;
        RECT 26.185 46.970 26.585 51.970 ;
        RECT 27.265 46.970 27.665 51.970 ;
        RECT 28.175 51.940 28.405 52.035 ;
        RECT 32.575 52.020 32.805 52.125 ;
        RECT 28.115 46.970 28.545 51.940 ;
        RECT 32.445 50.300 32.815 52.020 ;
        RECT 33.365 51.900 33.595 52.125 ;
        RECT 36.655 51.990 36.885 52.045 ;
        RECT 32.575 50.125 32.805 50.300 ;
        RECT 33.355 50.220 33.725 51.900 ;
        RECT 33.365 50.125 33.595 50.220 ;
        RECT 32.725 49.680 33.445 49.940 ;
        RECT 25.735 46.600 26.195 46.830 ;
        RECT 27.665 46.710 28.125 46.830 ;
        RECT 27.515 46.600 28.125 46.710 ;
        RECT 30.495 46.660 31.265 47.730 ;
        RECT 32.585 47.500 33.305 47.760 ;
        RECT 32.425 47.210 32.655 47.350 ;
        RECT 21.225 46.340 21.455 46.430 ;
        RECT 22.015 46.340 22.245 46.450 ;
        RECT 27.515 46.430 28.095 46.600 ;
        RECT 32.285 46.440 32.675 47.210 ;
        RECT 33.215 47.200 33.445 47.350 ;
        RECT 33.205 46.460 33.575 47.200 ;
        RECT 36.505 47.020 36.935 51.990 ;
        RECT 37.445 51.980 37.675 52.045 ;
        RECT 38.585 51.980 38.815 52.045 ;
        RECT 37.385 46.980 37.785 51.980 ;
        RECT 38.465 46.980 38.865 51.980 ;
        RECT 39.375 51.950 39.605 52.045 ;
        RECT 43.795 51.990 44.025 52.095 ;
        RECT 39.315 46.980 39.745 51.950 ;
        RECT 43.665 50.270 44.035 51.990 ;
        RECT 44.585 51.870 44.815 52.095 ;
        RECT 47.875 51.960 48.105 52.015 ;
        RECT 43.795 50.095 44.025 50.270 ;
        RECT 44.575 50.190 44.945 51.870 ;
        RECT 44.585 50.095 44.815 50.190 ;
        RECT 43.945 49.650 44.665 49.910 ;
        RECT 36.935 46.610 37.395 46.840 ;
        RECT 38.865 46.720 39.325 46.840 ;
        RECT 38.715 46.610 39.325 46.720 ;
        RECT 41.715 46.630 42.485 47.700 ;
        RECT 43.805 47.470 44.525 47.730 ;
        RECT 43.645 47.180 43.875 47.320 ;
        RECT 32.425 46.350 32.655 46.440 ;
        RECT 33.215 46.350 33.445 46.460 ;
        RECT 38.715 46.440 39.295 46.610 ;
        RECT 43.505 46.410 43.895 47.180 ;
        RECT 44.435 47.170 44.665 47.320 ;
        RECT 44.425 46.430 44.795 47.170 ;
        RECT 47.725 46.990 48.155 51.960 ;
        RECT 48.665 51.950 48.895 52.015 ;
        RECT 49.805 51.950 50.035 52.015 ;
        RECT 48.605 46.950 49.005 51.950 ;
        RECT 49.685 46.950 50.085 51.950 ;
        RECT 50.595 51.920 50.825 52.015 ;
        RECT 55.045 51.970 55.275 52.075 ;
        RECT 50.535 46.950 50.965 51.920 ;
        RECT 54.915 50.250 55.285 51.970 ;
        RECT 55.835 51.850 56.065 52.075 ;
        RECT 59.125 51.940 59.355 51.995 ;
        RECT 55.045 50.075 55.275 50.250 ;
        RECT 55.825 50.170 56.195 51.850 ;
        RECT 55.835 50.075 56.065 50.170 ;
        RECT 55.195 49.630 55.915 49.890 ;
        RECT 48.155 46.580 48.615 46.810 ;
        RECT 50.085 46.690 50.545 46.810 ;
        RECT 49.935 46.580 50.545 46.690 ;
        RECT 52.965 46.610 53.735 47.680 ;
        RECT 55.055 47.450 55.775 47.710 ;
        RECT 54.895 47.160 55.125 47.300 ;
        RECT 43.645 46.320 43.875 46.410 ;
        RECT 44.435 46.320 44.665 46.430 ;
        RECT 49.935 46.410 50.515 46.580 ;
        RECT 54.755 46.390 55.145 47.160 ;
        RECT 55.685 47.150 55.915 47.300 ;
        RECT 55.675 46.410 56.045 47.150 ;
        RECT 58.975 46.970 59.405 51.940 ;
        RECT 59.915 51.930 60.145 51.995 ;
        RECT 61.055 51.930 61.285 51.995 ;
        RECT 59.855 46.930 60.255 51.930 ;
        RECT 60.935 46.930 61.335 51.930 ;
        RECT 61.845 51.900 62.075 51.995 ;
        RECT 66.265 51.960 66.495 52.065 ;
        RECT 61.785 46.930 62.215 51.900 ;
        RECT 66.135 50.240 66.505 51.960 ;
        RECT 67.055 51.840 67.285 52.065 ;
        RECT 70.345 51.930 70.575 51.985 ;
        RECT 66.265 50.065 66.495 50.240 ;
        RECT 67.045 50.160 67.415 51.840 ;
        RECT 67.055 50.065 67.285 50.160 ;
        RECT 66.415 49.620 67.135 49.880 ;
        RECT 59.405 46.560 59.865 46.790 ;
        RECT 61.335 46.670 61.795 46.790 ;
        RECT 61.185 46.560 61.795 46.670 ;
        RECT 64.185 46.600 64.955 47.670 ;
        RECT 66.275 47.440 66.995 47.700 ;
        RECT 66.115 47.150 66.345 47.290 ;
        RECT 54.895 46.300 55.125 46.390 ;
        RECT 55.685 46.300 55.915 46.410 ;
        RECT 61.185 46.390 61.765 46.560 ;
        RECT 65.975 46.380 66.365 47.150 ;
        RECT 66.905 47.140 67.135 47.290 ;
        RECT 66.895 46.400 67.265 47.140 ;
        RECT 70.195 46.960 70.625 51.930 ;
        RECT 71.135 51.920 71.365 51.985 ;
        RECT 72.275 51.920 72.505 51.985 ;
        RECT 71.075 46.920 71.475 51.920 ;
        RECT 72.155 46.920 72.555 51.920 ;
        RECT 73.065 51.890 73.295 51.985 ;
        RECT 77.505 51.950 77.735 52.055 ;
        RECT 73.005 46.920 73.435 51.890 ;
        RECT 77.375 50.230 77.745 51.950 ;
        RECT 78.295 51.830 78.525 52.055 ;
        RECT 81.585 51.920 81.815 51.975 ;
        RECT 77.505 50.055 77.735 50.230 ;
        RECT 78.285 50.150 78.655 51.830 ;
        RECT 78.295 50.055 78.525 50.150 ;
        RECT 77.655 49.610 78.375 49.870 ;
        RECT 70.625 46.550 71.085 46.780 ;
        RECT 72.555 46.660 73.015 46.780 ;
        RECT 72.405 46.550 73.015 46.660 ;
        RECT 75.425 46.590 76.195 47.660 ;
        RECT 77.515 47.430 78.235 47.690 ;
        RECT 77.355 47.140 77.585 47.280 ;
        RECT 66.115 46.290 66.345 46.380 ;
        RECT 66.905 46.290 67.135 46.400 ;
        RECT 72.405 46.380 72.985 46.550 ;
        RECT 77.215 46.370 77.605 47.140 ;
        RECT 78.145 47.130 78.375 47.280 ;
        RECT 78.135 46.390 78.505 47.130 ;
        RECT 81.435 46.950 81.865 51.920 ;
        RECT 82.375 51.910 82.605 51.975 ;
        RECT 83.515 51.910 83.745 51.975 ;
        RECT 82.315 46.910 82.715 51.910 ;
        RECT 83.395 46.910 83.795 51.910 ;
        RECT 84.305 51.880 84.535 51.975 ;
        RECT 88.755 51.960 88.985 52.065 ;
        RECT 84.245 46.910 84.675 51.880 ;
        RECT 88.625 50.240 88.995 51.960 ;
        RECT 89.545 51.840 89.775 52.065 ;
        RECT 92.835 51.930 93.065 51.985 ;
        RECT 88.755 50.065 88.985 50.240 ;
        RECT 89.535 50.160 89.905 51.840 ;
        RECT 89.545 50.065 89.775 50.160 ;
        RECT 88.905 49.620 89.625 49.880 ;
        RECT 81.865 46.540 82.325 46.770 ;
        RECT 83.795 46.650 84.255 46.770 ;
        RECT 83.645 46.540 84.255 46.650 ;
        RECT 86.675 46.600 87.445 47.670 ;
        RECT 88.765 47.440 89.485 47.700 ;
        RECT 88.605 47.150 88.835 47.290 ;
        RECT 77.355 46.280 77.585 46.370 ;
        RECT 78.145 46.280 78.375 46.390 ;
        RECT 83.645 46.370 84.225 46.540 ;
        RECT 88.465 46.380 88.855 47.150 ;
        RECT 89.395 47.140 89.625 47.290 ;
        RECT 89.385 46.400 89.755 47.140 ;
        RECT 92.685 46.960 93.115 51.930 ;
        RECT 93.625 51.920 93.855 51.985 ;
        RECT 94.765 51.920 94.995 51.985 ;
        RECT 93.565 46.920 93.965 51.920 ;
        RECT 94.645 46.920 95.045 51.920 ;
        RECT 95.555 51.890 95.785 51.985 ;
        RECT 100.035 51.950 100.265 52.055 ;
        RECT 95.495 46.920 95.925 51.890 ;
        RECT 99.905 50.230 100.275 51.950 ;
        RECT 100.825 51.830 101.055 52.055 ;
        RECT 104.115 51.920 104.345 51.975 ;
        RECT 100.035 50.055 100.265 50.230 ;
        RECT 100.815 50.150 101.185 51.830 ;
        RECT 100.825 50.055 101.055 50.150 ;
        RECT 100.185 49.610 100.905 49.870 ;
        RECT 93.115 46.550 93.575 46.780 ;
        RECT 95.045 46.660 95.505 46.780 ;
        RECT 94.895 46.550 95.505 46.660 ;
        RECT 97.955 46.590 98.725 47.660 ;
        RECT 100.045 47.430 100.765 47.690 ;
        RECT 99.885 47.140 100.115 47.280 ;
        RECT 88.605 46.290 88.835 46.380 ;
        RECT 89.395 46.290 89.625 46.400 ;
        RECT 94.895 46.380 95.475 46.550 ;
        RECT 99.745 46.370 100.135 47.140 ;
        RECT 100.675 47.130 100.905 47.280 ;
        RECT 100.665 46.390 101.035 47.130 ;
        RECT 103.965 46.950 104.395 51.920 ;
        RECT 104.905 51.910 105.135 51.975 ;
        RECT 106.045 51.910 106.275 51.975 ;
        RECT 104.845 46.910 105.245 51.910 ;
        RECT 105.925 46.910 106.325 51.910 ;
        RECT 106.835 51.880 107.065 51.975 ;
        RECT 111.305 51.950 111.535 52.055 ;
        RECT 106.775 46.910 107.205 51.880 ;
        RECT 111.175 50.230 111.545 51.950 ;
        RECT 112.095 51.830 112.325 52.055 ;
        RECT 115.385 51.920 115.615 51.975 ;
        RECT 111.305 50.055 111.535 50.230 ;
        RECT 112.085 50.150 112.455 51.830 ;
        RECT 112.095 50.055 112.325 50.150 ;
        RECT 111.455 49.610 112.175 49.870 ;
        RECT 104.395 46.540 104.855 46.770 ;
        RECT 106.325 46.650 106.785 46.770 ;
        RECT 106.175 46.540 106.785 46.650 ;
        RECT 109.225 46.590 109.995 47.660 ;
        RECT 111.315 47.430 112.035 47.690 ;
        RECT 111.155 47.140 111.385 47.280 ;
        RECT 99.885 46.280 100.115 46.370 ;
        RECT 100.675 46.280 100.905 46.390 ;
        RECT 106.175 46.370 106.755 46.540 ;
        RECT 111.015 46.370 111.405 47.140 ;
        RECT 111.945 47.130 112.175 47.280 ;
        RECT 111.935 46.390 112.305 47.130 ;
        RECT 115.235 46.950 115.665 51.920 ;
        RECT 116.175 51.910 116.405 51.975 ;
        RECT 117.315 51.910 117.545 51.975 ;
        RECT 116.115 46.910 116.515 51.910 ;
        RECT 117.195 46.910 117.595 51.910 ;
        RECT 118.105 51.880 118.335 51.975 ;
        RECT 122.555 51.950 122.785 52.055 ;
        RECT 118.045 46.910 118.475 51.880 ;
        RECT 122.425 50.230 122.795 51.950 ;
        RECT 123.345 51.830 123.575 52.055 ;
        RECT 126.635 51.920 126.865 51.975 ;
        RECT 122.555 50.055 122.785 50.230 ;
        RECT 123.335 50.150 123.705 51.830 ;
        RECT 123.345 50.055 123.575 50.150 ;
        RECT 122.705 49.610 123.425 49.870 ;
        RECT 115.665 46.540 116.125 46.770 ;
        RECT 117.595 46.650 118.055 46.770 ;
        RECT 117.445 46.540 118.055 46.650 ;
        RECT 120.475 46.590 121.245 47.660 ;
        RECT 122.565 47.430 123.285 47.690 ;
        RECT 122.405 47.140 122.635 47.280 ;
        RECT 111.155 46.280 111.385 46.370 ;
        RECT 111.945 46.280 112.175 46.390 ;
        RECT 117.445 46.370 118.025 46.540 ;
        RECT 122.265 46.370 122.655 47.140 ;
        RECT 123.195 47.130 123.425 47.280 ;
        RECT 123.185 46.390 123.555 47.130 ;
        RECT 126.485 46.950 126.915 51.920 ;
        RECT 127.425 51.910 127.655 51.975 ;
        RECT 128.565 51.910 128.795 51.975 ;
        RECT 127.365 46.910 127.765 51.910 ;
        RECT 128.445 46.910 128.845 51.910 ;
        RECT 129.355 51.880 129.585 51.975 ;
        RECT 129.295 46.910 129.725 51.880 ;
        RECT 126.915 46.540 127.375 46.770 ;
        RECT 128.845 46.650 129.305 46.770 ;
        RECT 128.695 46.540 129.305 46.650 ;
        RECT 122.405 46.280 122.635 46.370 ;
        RECT 123.195 46.280 123.425 46.390 ;
        RECT 128.695 46.370 129.275 46.540 ;
        RECT 21.505 45.950 21.965 46.180 ;
        RECT 32.705 45.960 33.165 46.190 ;
        RECT 43.925 45.930 44.385 46.160 ;
        RECT 55.175 45.910 55.635 46.140 ;
        RECT 66.395 45.900 66.855 46.130 ;
        RECT 77.635 45.890 78.095 46.120 ;
        RECT 88.885 45.900 89.345 46.130 ;
        RECT 100.165 45.890 100.625 46.120 ;
        RECT 111.435 45.890 111.895 46.120 ;
        RECT 122.685 45.890 123.145 46.120 ;
        RECT 29.055 45.020 41.225 45.030 ;
        RECT 17.855 45.005 41.225 45.020 ;
        RECT 15.900 45.000 41.225 45.005 ;
        RECT 15.900 44.980 52.445 45.000 ;
        RECT 15.900 44.970 63.695 44.980 ;
        RECT 15.900 44.960 74.915 44.970 ;
        RECT 85.235 44.960 97.405 44.970 ;
        RECT 15.900 43.880 131.205 44.960 ;
        RECT 15.900 43.870 30.025 43.880 ;
        RECT 15.900 43.855 18.690 43.870 ;
        RECT 15.900 41.620 17.050 43.855 ;
        RECT 40.275 43.850 131.205 43.880 ;
        RECT 51.525 43.830 131.205 43.850 ;
        RECT 62.745 43.820 131.205 43.830 ;
        RECT 73.985 43.810 86.155 43.820 ;
        RECT 96.515 43.810 131.205 43.820 ;
        RECT 29.015 43.330 41.185 43.340 ;
        RECT 17.815 43.310 41.185 43.330 ;
        RECT 142.830 43.320 144.150 43.340 ;
        RECT 17.815 43.290 52.405 43.310 ;
        RECT 140.750 43.300 144.150 43.320 ;
        RECT 17.815 43.280 63.655 43.290 ;
        RECT 119.895 43.280 144.150 43.300 ;
        RECT 17.815 43.270 74.875 43.280 ;
        RECT 85.195 43.270 97.365 43.280 ;
        RECT 108.685 43.270 144.150 43.280 ;
        RECT 17.815 42.180 144.150 43.270 ;
        RECT 18.755 42.150 144.150 42.180 ;
        RECT 18.755 42.120 131.165 42.150 ;
        RECT 18.755 42.090 109.655 42.120 ;
        RECT 18.755 42.080 98.445 42.090 ;
        RECT 41.325 42.070 98.445 42.080 ;
        RECT 142.830 42.070 144.150 42.150 ;
        RECT 41.325 42.060 87.205 42.070 ;
        RECT 75.035 42.050 87.205 42.060 ;
        RECT 15.900 41.540 19.685 41.620 ;
        RECT 142.070 41.610 146.210 41.640 ;
        RECT 119.855 41.590 146.210 41.610 ;
        RECT 108.645 41.550 146.210 41.590 ;
        RECT 15.900 41.520 42.165 41.540 ;
        RECT 97.445 41.530 146.210 41.550 ;
        RECT 15.900 41.510 75.875 41.520 ;
        RECT 86.235 41.510 146.210 41.530 ;
        RECT 15.900 40.500 146.210 41.510 ;
        RECT 15.900 40.480 142.320 40.500 ;
        RECT 15.900 40.470 140.920 40.480 ;
        RECT 18.715 40.460 140.920 40.470 ;
        RECT 142.070 40.460 142.250 40.480 ;
        RECT 18.715 40.440 120.815 40.460 ;
        RECT 18.715 40.400 109.615 40.440 ;
        RECT 18.715 40.390 98.405 40.400 ;
        RECT 41.285 40.380 98.405 40.390 ;
        RECT 41.285 40.370 87.165 40.380 ;
        RECT 74.995 40.360 87.165 40.370 ;
        RECT 26.775 39.230 27.235 39.460 ;
        RECT 38.055 39.230 38.515 39.460 ;
        RECT 49.345 39.210 49.805 39.440 ;
        RECT 60.565 39.210 61.025 39.440 ;
        RECT 71.765 39.210 72.225 39.440 ;
        RECT 83.055 39.200 83.515 39.430 ;
        RECT 94.295 39.220 94.755 39.450 ;
        RECT 105.505 39.240 105.965 39.470 ;
        RECT 116.705 39.280 117.165 39.510 ;
        RECT 127.915 39.300 128.375 39.530 ;
        RECT 20.645 38.810 21.225 38.980 ;
        RECT 26.495 38.960 26.725 39.070 ;
        RECT 27.285 38.980 27.515 39.070 ;
        RECT 20.615 38.700 21.225 38.810 ;
        RECT 20.615 38.580 21.075 38.700 ;
        RECT 22.545 38.580 23.005 38.810 ;
        RECT 20.195 33.470 20.625 38.440 ;
        RECT 20.335 33.375 20.565 33.470 ;
        RECT 21.075 33.440 21.475 38.440 ;
        RECT 22.155 33.440 22.555 38.440 ;
        RECT 21.125 33.375 21.355 33.440 ;
        RECT 22.265 33.375 22.495 33.440 ;
        RECT 23.005 33.430 23.435 38.400 ;
        RECT 26.365 38.220 26.735 38.960 ;
        RECT 26.495 38.070 26.725 38.220 ;
        RECT 27.265 38.210 27.655 38.980 ;
        RECT 31.925 38.810 32.505 38.980 ;
        RECT 37.775 38.960 38.005 39.070 ;
        RECT 38.565 38.980 38.795 39.070 ;
        RECT 27.285 38.070 27.515 38.210 ;
        RECT 26.635 37.660 27.355 37.920 ;
        RECT 28.675 37.690 29.445 38.760 ;
        RECT 31.895 38.700 32.505 38.810 ;
        RECT 31.895 38.580 32.355 38.700 ;
        RECT 33.825 38.580 34.285 38.810 ;
        RECT 26.495 35.480 27.215 35.740 ;
        RECT 26.345 35.200 26.575 35.295 ;
        RECT 26.215 33.520 26.585 35.200 ;
        RECT 27.135 35.120 27.365 35.295 ;
        RECT 23.055 33.375 23.285 33.430 ;
        RECT 26.345 33.295 26.575 33.520 ;
        RECT 27.125 33.400 27.495 35.120 ;
        RECT 31.475 33.470 31.905 38.440 ;
        RECT 27.135 33.295 27.365 33.400 ;
        RECT 31.615 33.375 31.845 33.470 ;
        RECT 32.355 33.440 32.755 38.440 ;
        RECT 33.435 33.440 33.835 38.440 ;
        RECT 32.405 33.375 32.635 33.440 ;
        RECT 33.545 33.375 33.775 33.440 ;
        RECT 34.285 33.430 34.715 38.400 ;
        RECT 37.645 38.220 38.015 38.960 ;
        RECT 37.775 38.070 38.005 38.220 ;
        RECT 38.545 38.210 38.935 38.980 ;
        RECT 43.215 38.790 43.795 38.960 ;
        RECT 49.065 38.940 49.295 39.050 ;
        RECT 49.855 38.960 50.085 39.050 ;
        RECT 38.565 38.070 38.795 38.210 ;
        RECT 37.915 37.660 38.635 37.920 ;
        RECT 39.955 37.690 40.725 38.760 ;
        RECT 43.185 38.680 43.795 38.790 ;
        RECT 43.185 38.560 43.645 38.680 ;
        RECT 45.115 38.560 45.575 38.790 ;
        RECT 37.775 35.480 38.495 35.740 ;
        RECT 37.625 35.200 37.855 35.295 ;
        RECT 37.495 33.520 37.865 35.200 ;
        RECT 38.415 35.120 38.645 35.295 ;
        RECT 34.335 33.375 34.565 33.430 ;
        RECT 37.625 33.295 37.855 33.520 ;
        RECT 38.405 33.400 38.775 35.120 ;
        RECT 42.765 33.450 43.195 38.420 ;
        RECT 38.415 33.295 38.645 33.400 ;
        RECT 42.905 33.355 43.135 33.450 ;
        RECT 43.645 33.420 44.045 38.420 ;
        RECT 44.725 33.420 45.125 38.420 ;
        RECT 43.695 33.355 43.925 33.420 ;
        RECT 44.835 33.355 45.065 33.420 ;
        RECT 45.575 33.410 46.005 38.380 ;
        RECT 48.935 38.200 49.305 38.940 ;
        RECT 49.065 38.050 49.295 38.200 ;
        RECT 49.835 38.190 50.225 38.960 ;
        RECT 54.435 38.790 55.015 38.960 ;
        RECT 60.285 38.940 60.515 39.050 ;
        RECT 61.075 38.960 61.305 39.050 ;
        RECT 49.855 38.050 50.085 38.190 ;
        RECT 49.205 37.640 49.925 37.900 ;
        RECT 51.245 37.670 52.015 38.740 ;
        RECT 54.405 38.680 55.015 38.790 ;
        RECT 54.405 38.560 54.865 38.680 ;
        RECT 56.335 38.560 56.795 38.790 ;
        RECT 49.065 35.460 49.785 35.720 ;
        RECT 48.915 35.180 49.145 35.275 ;
        RECT 48.785 33.500 49.155 35.180 ;
        RECT 49.705 35.100 49.935 35.275 ;
        RECT 45.625 33.355 45.855 33.410 ;
        RECT 48.915 33.275 49.145 33.500 ;
        RECT 49.695 33.380 50.065 35.100 ;
        RECT 53.985 33.450 54.415 38.420 ;
        RECT 49.705 33.275 49.935 33.380 ;
        RECT 54.125 33.355 54.355 33.450 ;
        RECT 54.865 33.420 55.265 38.420 ;
        RECT 55.945 33.420 56.345 38.420 ;
        RECT 54.915 33.355 55.145 33.420 ;
        RECT 56.055 33.355 56.285 33.420 ;
        RECT 56.795 33.410 57.225 38.380 ;
        RECT 60.155 38.200 60.525 38.940 ;
        RECT 60.285 38.050 60.515 38.200 ;
        RECT 61.055 38.190 61.445 38.960 ;
        RECT 65.635 38.790 66.215 38.960 ;
        RECT 71.485 38.940 71.715 39.050 ;
        RECT 72.275 38.960 72.505 39.050 ;
        RECT 61.075 38.050 61.305 38.190 ;
        RECT 60.425 37.640 61.145 37.900 ;
        RECT 62.465 37.670 63.235 38.740 ;
        RECT 65.605 38.680 66.215 38.790 ;
        RECT 65.605 38.560 66.065 38.680 ;
        RECT 67.535 38.560 67.995 38.790 ;
        RECT 60.285 35.460 61.005 35.720 ;
        RECT 60.135 35.180 60.365 35.275 ;
        RECT 60.005 33.500 60.375 35.180 ;
        RECT 60.925 35.100 61.155 35.275 ;
        RECT 56.845 33.355 57.075 33.410 ;
        RECT 60.135 33.275 60.365 33.500 ;
        RECT 60.915 33.380 61.285 35.100 ;
        RECT 65.185 33.450 65.615 38.420 ;
        RECT 60.925 33.275 61.155 33.380 ;
        RECT 65.325 33.355 65.555 33.450 ;
        RECT 66.065 33.420 66.465 38.420 ;
        RECT 67.145 33.420 67.545 38.420 ;
        RECT 66.115 33.355 66.345 33.420 ;
        RECT 67.255 33.355 67.485 33.420 ;
        RECT 67.995 33.410 68.425 38.380 ;
        RECT 71.355 38.200 71.725 38.940 ;
        RECT 71.485 38.050 71.715 38.200 ;
        RECT 72.255 38.190 72.645 38.960 ;
        RECT 76.925 38.780 77.505 38.950 ;
        RECT 82.775 38.930 83.005 39.040 ;
        RECT 83.565 38.950 83.795 39.040 ;
        RECT 72.275 38.050 72.505 38.190 ;
        RECT 71.625 37.640 72.345 37.900 ;
        RECT 73.665 37.670 74.435 38.740 ;
        RECT 76.895 38.670 77.505 38.780 ;
        RECT 76.895 38.550 77.355 38.670 ;
        RECT 78.825 38.550 79.285 38.780 ;
        RECT 71.485 35.460 72.205 35.720 ;
        RECT 71.335 35.180 71.565 35.275 ;
        RECT 71.205 33.500 71.575 35.180 ;
        RECT 72.125 35.100 72.355 35.275 ;
        RECT 68.045 33.355 68.275 33.410 ;
        RECT 71.335 33.275 71.565 33.500 ;
        RECT 72.115 33.380 72.485 35.100 ;
        RECT 76.475 33.440 76.905 38.410 ;
        RECT 72.125 33.275 72.355 33.380 ;
        RECT 76.615 33.345 76.845 33.440 ;
        RECT 77.355 33.410 77.755 38.410 ;
        RECT 78.435 33.410 78.835 38.410 ;
        RECT 77.405 33.345 77.635 33.410 ;
        RECT 78.545 33.345 78.775 33.410 ;
        RECT 79.285 33.400 79.715 38.370 ;
        RECT 82.645 38.190 83.015 38.930 ;
        RECT 82.775 38.040 83.005 38.190 ;
        RECT 83.545 38.180 83.935 38.950 ;
        RECT 88.165 38.800 88.745 38.970 ;
        RECT 94.015 38.950 94.245 39.060 ;
        RECT 94.805 38.970 95.035 39.060 ;
        RECT 83.565 38.040 83.795 38.180 ;
        RECT 82.915 37.630 83.635 37.890 ;
        RECT 84.955 37.660 85.725 38.730 ;
        RECT 88.135 38.690 88.745 38.800 ;
        RECT 88.135 38.570 88.595 38.690 ;
        RECT 90.065 38.570 90.525 38.800 ;
        RECT 82.775 35.450 83.495 35.710 ;
        RECT 82.625 35.170 82.855 35.265 ;
        RECT 82.495 33.490 82.865 35.170 ;
        RECT 83.415 35.090 83.645 35.265 ;
        RECT 79.335 33.345 79.565 33.400 ;
        RECT 82.625 33.265 82.855 33.490 ;
        RECT 83.405 33.370 83.775 35.090 ;
        RECT 87.715 33.460 88.145 38.430 ;
        RECT 83.415 33.265 83.645 33.370 ;
        RECT 87.855 33.365 88.085 33.460 ;
        RECT 88.595 33.430 88.995 38.430 ;
        RECT 89.675 33.430 90.075 38.430 ;
        RECT 88.645 33.365 88.875 33.430 ;
        RECT 89.785 33.365 90.015 33.430 ;
        RECT 90.525 33.420 90.955 38.390 ;
        RECT 93.885 38.210 94.255 38.950 ;
        RECT 94.015 38.060 94.245 38.210 ;
        RECT 94.785 38.200 95.175 38.970 ;
        RECT 99.375 38.820 99.955 38.990 ;
        RECT 105.225 38.970 105.455 39.080 ;
        RECT 106.015 38.990 106.245 39.080 ;
        RECT 94.805 38.060 95.035 38.200 ;
        RECT 94.155 37.650 94.875 37.910 ;
        RECT 96.195 37.680 96.965 38.750 ;
        RECT 99.345 38.710 99.955 38.820 ;
        RECT 99.345 38.590 99.805 38.710 ;
        RECT 101.275 38.590 101.735 38.820 ;
        RECT 94.015 35.470 94.735 35.730 ;
        RECT 93.865 35.190 94.095 35.285 ;
        RECT 93.735 33.510 94.105 35.190 ;
        RECT 94.655 35.110 94.885 35.285 ;
        RECT 90.575 33.365 90.805 33.420 ;
        RECT 93.865 33.285 94.095 33.510 ;
        RECT 94.645 33.390 95.015 35.110 ;
        RECT 98.925 33.480 99.355 38.450 ;
        RECT 94.655 33.285 94.885 33.390 ;
        RECT 99.065 33.385 99.295 33.480 ;
        RECT 99.805 33.450 100.205 38.450 ;
        RECT 100.885 33.450 101.285 38.450 ;
        RECT 99.855 33.385 100.085 33.450 ;
        RECT 100.995 33.385 101.225 33.450 ;
        RECT 101.735 33.440 102.165 38.410 ;
        RECT 105.095 38.230 105.465 38.970 ;
        RECT 105.225 38.080 105.455 38.230 ;
        RECT 105.995 38.220 106.385 38.990 ;
        RECT 110.575 38.860 111.155 39.030 ;
        RECT 116.425 39.010 116.655 39.120 ;
        RECT 117.215 39.030 117.445 39.120 ;
        RECT 106.015 38.080 106.245 38.220 ;
        RECT 105.365 37.670 106.085 37.930 ;
        RECT 107.405 37.700 108.175 38.770 ;
        RECT 110.545 38.750 111.155 38.860 ;
        RECT 110.545 38.630 111.005 38.750 ;
        RECT 112.475 38.630 112.935 38.860 ;
        RECT 105.225 35.490 105.945 35.750 ;
        RECT 105.075 35.210 105.305 35.305 ;
        RECT 104.945 33.530 105.315 35.210 ;
        RECT 105.865 35.130 106.095 35.305 ;
        RECT 101.785 33.385 102.015 33.440 ;
        RECT 105.075 33.305 105.305 33.530 ;
        RECT 105.855 33.410 106.225 35.130 ;
        RECT 110.125 33.520 110.555 38.490 ;
        RECT 110.265 33.425 110.495 33.520 ;
        RECT 111.005 33.490 111.405 38.490 ;
        RECT 112.085 33.490 112.485 38.490 ;
        RECT 111.055 33.425 111.285 33.490 ;
        RECT 112.195 33.425 112.425 33.490 ;
        RECT 112.935 33.480 113.365 38.450 ;
        RECT 116.295 38.270 116.665 39.010 ;
        RECT 116.425 38.120 116.655 38.270 ;
        RECT 117.195 38.260 117.585 39.030 ;
        RECT 121.785 38.880 122.365 39.050 ;
        RECT 127.635 39.030 127.865 39.140 ;
        RECT 128.425 39.050 128.655 39.140 ;
        RECT 117.215 38.120 117.445 38.260 ;
        RECT 116.565 37.710 117.285 37.970 ;
        RECT 118.605 37.740 119.375 38.810 ;
        RECT 121.755 38.770 122.365 38.880 ;
        RECT 121.755 38.650 122.215 38.770 ;
        RECT 123.685 38.650 124.145 38.880 ;
        RECT 116.425 35.530 117.145 35.790 ;
        RECT 116.275 35.250 116.505 35.345 ;
        RECT 116.145 33.570 116.515 35.250 ;
        RECT 117.065 35.170 117.295 35.345 ;
        RECT 112.985 33.425 113.215 33.480 ;
        RECT 105.865 33.305 106.095 33.410 ;
        RECT 116.275 33.345 116.505 33.570 ;
        RECT 117.055 33.450 117.425 35.170 ;
        RECT 121.335 33.540 121.765 38.510 ;
        RECT 117.065 33.345 117.295 33.450 ;
        RECT 121.475 33.445 121.705 33.540 ;
        RECT 122.215 33.510 122.615 38.510 ;
        RECT 123.295 33.510 123.695 38.510 ;
        RECT 122.265 33.445 122.495 33.510 ;
        RECT 123.405 33.445 123.635 33.510 ;
        RECT 124.145 33.500 124.575 38.470 ;
        RECT 127.505 38.290 127.875 39.030 ;
        RECT 127.635 38.140 127.865 38.290 ;
        RECT 128.405 38.280 128.795 39.050 ;
        RECT 128.425 38.140 128.655 38.280 ;
        RECT 127.775 37.730 128.495 37.990 ;
        RECT 129.815 37.760 130.585 38.830 ;
        RECT 142.850 37.630 144.170 38.900 ;
        RECT 127.635 35.550 128.355 35.810 ;
        RECT 127.485 35.270 127.715 35.365 ;
        RECT 127.355 33.590 127.725 35.270 ;
        RECT 128.275 35.190 128.505 35.365 ;
        RECT 124.195 33.445 124.425 33.500 ;
        RECT 127.485 33.365 127.715 33.590 ;
        RECT 128.265 33.470 128.635 35.190 ;
        RECT 128.275 33.365 128.505 33.470 ;
        RECT 20.615 32.940 21.075 33.170 ;
        RECT 22.545 33.130 23.005 33.170 ;
        RECT 22.485 32.850 23.115 33.130 ;
        RECT 26.625 32.860 27.085 33.090 ;
        RECT 31.895 32.940 32.355 33.170 ;
        RECT 33.825 33.130 34.285 33.170 ;
        RECT 33.765 32.850 34.395 33.130 ;
        RECT 37.905 32.860 38.365 33.090 ;
        RECT 43.185 32.920 43.645 33.150 ;
        RECT 45.115 33.110 45.575 33.150 ;
        RECT 45.055 32.830 45.685 33.110 ;
        RECT 49.195 32.840 49.655 33.070 ;
        RECT 54.405 32.920 54.865 33.150 ;
        RECT 56.335 33.110 56.795 33.150 ;
        RECT 56.275 32.830 56.905 33.110 ;
        RECT 60.415 32.840 60.875 33.070 ;
        RECT 65.605 32.920 66.065 33.150 ;
        RECT 67.535 33.110 67.995 33.150 ;
        RECT 67.475 32.830 68.105 33.110 ;
        RECT 71.615 32.840 72.075 33.070 ;
        RECT 76.895 32.910 77.355 33.140 ;
        RECT 78.825 33.100 79.285 33.140 ;
        RECT 78.765 32.820 79.395 33.100 ;
        RECT 82.905 32.830 83.365 33.060 ;
        RECT 88.135 32.930 88.595 33.160 ;
        RECT 90.065 33.120 90.525 33.160 ;
        RECT 90.005 32.840 90.635 33.120 ;
        RECT 94.145 32.850 94.605 33.080 ;
        RECT 99.345 32.950 99.805 33.180 ;
        RECT 101.275 33.140 101.735 33.180 ;
        RECT 101.215 32.860 101.845 33.140 ;
        RECT 105.355 32.870 105.815 33.100 ;
        RECT 110.545 32.990 111.005 33.220 ;
        RECT 112.475 33.180 112.935 33.220 ;
        RECT 112.415 32.900 113.045 33.180 ;
        RECT 116.555 32.910 117.015 33.140 ;
        RECT 121.755 33.010 122.215 33.240 ;
        RECT 123.685 33.200 124.145 33.240 ;
        RECT 123.625 32.920 124.255 33.200 ;
        RECT 127.765 32.930 128.225 33.160 ;
        RECT 23.185 30.880 27.925 31.180 ;
        RECT 34.465 30.880 39.205 31.180 ;
        RECT 45.755 30.860 50.495 31.160 ;
        RECT 56.975 30.860 61.715 31.160 ;
        RECT 68.175 30.860 72.915 31.160 ;
        RECT 79.465 30.850 84.205 31.150 ;
        RECT 90.705 30.870 95.445 31.170 ;
        RECT 101.915 30.890 106.655 31.190 ;
        RECT 113.115 30.930 117.855 31.230 ;
        RECT 124.325 30.950 129.065 31.250 ;
        RECT 19.485 20.270 19.905 30.160 ;
        RECT 19.585 20.090 19.815 20.270 ;
        RECT 20.805 20.260 21.175 30.210 ;
        RECT 20.875 20.090 21.105 20.260 ;
        RECT 21.935 20.220 22.305 30.170 ;
        RECT 27.255 20.270 27.615 30.190 ;
        RECT 30.765 20.270 31.185 30.160 ;
        RECT 22.015 20.090 22.245 20.220 ;
        RECT 27.305 20.090 27.535 20.270 ;
        RECT 30.865 20.090 31.095 20.270 ;
        RECT 32.085 20.260 32.455 30.210 ;
        RECT 32.155 20.090 32.385 20.260 ;
        RECT 33.215 20.220 33.585 30.170 ;
        RECT 38.535 20.270 38.895 30.190 ;
        RECT 33.295 20.090 33.525 20.220 ;
        RECT 38.585 20.090 38.815 20.270 ;
        RECT 42.055 20.250 42.475 30.140 ;
        RECT 42.155 20.070 42.385 20.250 ;
        RECT 43.375 20.240 43.745 30.190 ;
        RECT 43.445 20.070 43.675 20.240 ;
        RECT 44.505 20.200 44.875 30.150 ;
        RECT 49.825 20.250 50.185 30.170 ;
        RECT 53.275 20.250 53.695 30.140 ;
        RECT 44.585 20.070 44.815 20.200 ;
        RECT 49.875 20.070 50.105 20.250 ;
        RECT 53.375 20.070 53.605 20.250 ;
        RECT 54.595 20.240 54.965 30.190 ;
        RECT 54.665 20.070 54.895 20.240 ;
        RECT 55.725 20.200 56.095 30.150 ;
        RECT 61.045 20.250 61.405 30.170 ;
        RECT 64.475 20.250 64.895 30.140 ;
        RECT 55.805 20.070 56.035 20.200 ;
        RECT 61.095 20.070 61.325 20.250 ;
        RECT 64.575 20.070 64.805 20.250 ;
        RECT 65.795 20.240 66.165 30.190 ;
        RECT 65.865 20.070 66.095 20.240 ;
        RECT 66.925 20.200 67.295 30.150 ;
        RECT 72.245 20.250 72.605 30.170 ;
        RECT 67.005 20.070 67.235 20.200 ;
        RECT 72.295 20.070 72.525 20.250 ;
        RECT 75.765 20.240 76.185 30.130 ;
        RECT 75.865 20.060 76.095 20.240 ;
        RECT 77.085 20.230 77.455 30.180 ;
        RECT 77.155 20.060 77.385 20.230 ;
        RECT 78.215 20.190 78.585 30.140 ;
        RECT 83.535 20.240 83.895 30.160 ;
        RECT 87.005 20.260 87.425 30.150 ;
        RECT 78.295 20.060 78.525 20.190 ;
        RECT 83.585 20.060 83.815 20.240 ;
        RECT 87.105 20.080 87.335 20.260 ;
        RECT 88.325 20.250 88.695 30.200 ;
        RECT 88.395 20.080 88.625 20.250 ;
        RECT 89.455 20.210 89.825 30.160 ;
        RECT 94.775 20.260 95.135 30.180 ;
        RECT 98.215 20.280 98.635 30.170 ;
        RECT 89.535 20.080 89.765 20.210 ;
        RECT 94.825 20.080 95.055 20.260 ;
        RECT 98.315 20.100 98.545 20.280 ;
        RECT 99.535 20.270 99.905 30.220 ;
        RECT 99.605 20.100 99.835 20.270 ;
        RECT 100.665 20.230 101.035 30.180 ;
        RECT 105.985 20.280 106.345 30.200 ;
        RECT 109.415 20.320 109.835 30.210 ;
        RECT 100.745 20.100 100.975 20.230 ;
        RECT 106.035 20.100 106.265 20.280 ;
        RECT 109.515 20.140 109.745 20.320 ;
        RECT 110.735 20.310 111.105 30.260 ;
        RECT 110.805 20.140 111.035 20.310 ;
        RECT 111.865 20.270 112.235 30.220 ;
        RECT 117.185 20.320 117.545 30.240 ;
        RECT 120.625 20.340 121.045 30.230 ;
        RECT 111.945 20.140 112.175 20.270 ;
        RECT 117.235 20.140 117.465 20.320 ;
        RECT 120.725 20.160 120.955 20.340 ;
        RECT 121.945 20.330 122.315 30.280 ;
        RECT 122.015 20.160 122.245 20.330 ;
        RECT 123.075 20.290 123.445 30.240 ;
        RECT 128.395 20.340 128.755 30.260 ;
        RECT 123.155 20.160 123.385 20.290 ;
        RECT 128.445 20.160 128.675 20.340 ;
        RECT 132.345 20.170 132.755 30.180 ;
        RECT 137.735 30.120 137.965 30.130 ;
        RECT 132.445 20.130 132.675 20.170 ;
        RECT 137.665 20.080 138.055 30.120 ;
        RECT 19.775 19.610 20.925 19.920 ;
        RECT 22.185 19.620 27.335 19.900 ;
        RECT 31.055 19.610 32.205 19.920 ;
        RECT 33.465 19.620 38.615 19.900 ;
        RECT 42.345 19.590 43.495 19.900 ;
        RECT 44.755 19.600 49.905 19.880 ;
        RECT 53.565 19.590 54.715 19.900 ;
        RECT 55.975 19.600 61.125 19.880 ;
        RECT 64.765 19.590 65.915 19.900 ;
        RECT 67.175 19.600 72.325 19.880 ;
        RECT 76.055 19.580 77.205 19.890 ;
        RECT 78.465 19.590 83.615 19.870 ;
        RECT 87.295 19.600 88.445 19.910 ;
        RECT 89.705 19.610 94.855 19.890 ;
        RECT 98.505 19.620 99.655 19.930 ;
        RECT 100.915 19.630 106.065 19.910 ;
        RECT 109.705 19.660 110.855 19.970 ;
        RECT 112.115 19.670 117.265 19.950 ;
        RECT 120.915 19.680 122.065 19.990 ;
        RECT 123.325 19.690 128.475 19.970 ;
        RECT 132.635 19.640 138.025 19.930 ;
        RECT 142.940 19.110 144.080 37.630 ;
        RECT 13.940 18.460 17.635 18.530 ;
        RECT 117.755 18.510 131.425 18.530 ;
        RECT 106.545 18.470 131.425 18.510 ;
        RECT 13.940 18.440 41.565 18.460 ;
        RECT 95.345 18.450 131.425 18.470 ;
        RECT 13.940 18.430 75.275 18.440 ;
        RECT 84.135 18.430 131.425 18.450 ;
        RECT 13.940 17.380 131.425 18.430 ;
        RECT 142.890 17.990 144.140 19.110 ;
        RECT 145.070 18.880 146.210 40.500 ;
        RECT 145.030 17.960 146.250 18.880 ;
        RECT 13.950 17.370 15.100 17.380 ;
        RECT 16.615 17.360 120.215 17.380 ;
        RECT 16.615 17.320 109.015 17.360 ;
        RECT 16.615 17.310 97.805 17.320 ;
        RECT 39.185 17.300 97.805 17.310 ;
        RECT 39.185 17.290 86.565 17.300 ;
        RECT 72.895 17.280 86.565 17.290 ;
        RECT 117.765 16.950 140.620 16.960 ;
        RECT 142.040 16.950 148.010 16.980 ;
        RECT 117.765 16.940 148.010 16.950 ;
        RECT 106.555 16.900 148.010 16.940 ;
        RECT 16.625 16.870 41.575 16.890 ;
        RECT 95.355 16.880 148.010 16.900 ;
        RECT 16.625 16.860 75.285 16.870 ;
        RECT 84.145 16.860 148.010 16.880 ;
        RECT 16.625 15.840 148.010 16.860 ;
        RECT 16.625 15.820 142.660 15.840 ;
        RECT 16.625 15.810 140.620 15.820 ;
        RECT 142.040 15.810 142.660 15.820 ;
        RECT 16.625 15.790 120.225 15.810 ;
        RECT 16.625 15.750 109.025 15.790 ;
        RECT 16.625 15.740 97.815 15.750 ;
        RECT 39.195 15.730 97.815 15.740 ;
        RECT 39.195 15.720 86.575 15.730 ;
        RECT 72.905 15.710 86.575 15.720 ;
        RECT 131.215 15.460 132.585 15.470 ;
        RECT 12.290 15.390 17.625 15.450 ;
        RECT 117.795 15.440 132.785 15.460 ;
        RECT 106.585 15.400 132.785 15.440 ;
        RECT 12.290 15.370 41.585 15.390 ;
        RECT 95.385 15.380 132.785 15.400 ;
        RECT 12.290 15.360 75.295 15.370 ;
        RECT 84.175 15.360 132.785 15.380 ;
        RECT 12.290 14.320 132.785 15.360 ;
        RECT 142.905 15.040 144.045 15.050 ;
        RECT 12.290 14.310 131.445 14.320 ;
        RECT 12.290 14.300 120.235 14.310 ;
        RECT 12.320 14.280 13.470 14.300 ;
        RECT 16.655 14.290 120.235 14.300 ;
        RECT 16.655 14.250 109.035 14.290 ;
        RECT 16.655 14.240 97.825 14.250 ;
        RECT 39.225 14.230 97.825 14.240 ;
        RECT 39.225 14.220 86.585 14.230 ;
        RECT 72.935 14.210 86.585 14.220 ;
        RECT 142.850 13.920 144.100 15.040 ;
        RECT 145.020 14.870 146.160 14.980 ;
        RECT 144.980 13.950 146.200 14.870 ;
        RECT 16.965 13.800 17.435 13.810 ;
        RECT 10.800 13.780 17.435 13.800 ;
        RECT 10.800 13.720 17.555 13.780 ;
        RECT 117.845 13.770 131.445 13.790 ;
        RECT 106.635 13.730 131.445 13.770 ;
        RECT 10.800 13.700 41.585 13.720 ;
        RECT 95.435 13.710 131.445 13.730 ;
        RECT 10.800 13.690 75.295 13.700 ;
        RECT 84.225 13.690 131.445 13.710 ;
        RECT 10.800 12.650 131.445 13.690 ;
        RECT 16.705 12.640 131.445 12.650 ;
        RECT 16.705 12.620 120.235 12.640 ;
        RECT 16.705 12.580 109.035 12.620 ;
        RECT 16.705 12.570 97.825 12.580 ;
        RECT 39.275 12.560 97.825 12.570 ;
        RECT 39.275 12.550 86.585 12.560 ;
        RECT 72.985 12.540 86.585 12.550 ;
        RECT 128.755 12.240 130.465 12.250 ;
        RECT 117.545 12.220 119.255 12.230 ;
        RECT 106.345 12.180 108.055 12.190 ;
        RECT 27.615 12.170 29.325 12.180 ;
        RECT 38.895 12.170 40.605 12.180 ;
        RECT 25.675 11.030 29.325 12.170 ;
        RECT 36.955 11.030 40.605 12.170 ;
        RECT 95.135 12.160 96.845 12.170 ;
        RECT 50.185 12.150 51.895 12.160 ;
        RECT 61.405 12.150 63.115 12.160 ;
        RECT 72.605 12.150 74.315 12.160 ;
        RECT 25.675 11.020 27.625 11.030 ;
        RECT 36.955 11.020 38.905 11.030 ;
        RECT 48.245 11.010 51.895 12.150 ;
        RECT 59.465 11.010 63.115 12.150 ;
        RECT 70.665 11.010 74.315 12.150 ;
        RECT 83.895 12.140 85.605 12.150 ;
        RECT 48.245 11.000 50.195 11.010 ;
        RECT 59.465 11.000 61.415 11.010 ;
        RECT 70.665 11.000 72.615 11.010 ;
        RECT 81.955 11.000 85.605 12.140 ;
        RECT 93.195 11.020 96.845 12.160 ;
        RECT 104.405 11.040 108.055 12.180 ;
        RECT 115.605 11.080 119.255 12.220 ;
        RECT 126.815 11.100 130.465 12.240 ;
        RECT 126.815 11.090 128.765 11.100 ;
        RECT 115.605 11.070 117.555 11.080 ;
        RECT 104.405 11.030 106.355 11.040 ;
        RECT 93.195 11.010 95.145 11.020 ;
        RECT 81.955 10.990 83.905 11.000 ;
        RECT 142.905 8.580 144.045 13.920 ;
        RECT 74.420 7.440 144.045 8.580 ;
        RECT 74.420 1.410 75.560 7.440 ;
        RECT 145.020 6.630 146.160 13.950 ;
        RECT 93.650 5.490 146.160 6.630 ;
        RECT 93.650 1.480 94.790 5.490 ;
        RECT 146.870 4.560 148.010 15.840 ;
        RECT 113.130 3.420 148.010 4.560 ;
        RECT 113.130 1.610 114.270 3.420 ;
        RECT 149.460 2.770 150.600 64.660 ;
        RECT 131.940 1.880 150.600 2.770 ;
        RECT 131.800 1.630 150.600 1.880 ;
        RECT 74.290 0.160 75.680 1.410 ;
        RECT 93.500 0.230 94.890 1.480 ;
        RECT 112.900 0.360 114.290 1.610 ;
        RECT 131.800 1.380 133.490 1.630 ;
        RECT 151.730 1.420 152.870 66.900 ;
        RECT 131.800 0.430 133.540 1.380 ;
        RECT 113.130 0.330 114.270 0.360 ;
        RECT 151.600 0.300 152.970 1.420 ;
        RECT 93.650 0.150 94.790 0.230 ;
      LAYER met2 ;
        RECT 135.390 223.830 136.740 225.230 ;
        RECT 138.180 223.760 139.530 225.160 ;
        RECT 143.230 223.790 144.580 225.190 ;
        RECT 16.880 211.105 18.760 211.475 ;
        RECT 46.880 211.105 48.760 211.475 ;
        RECT 76.880 211.105 78.760 211.475 ;
        RECT 106.880 211.105 108.760 211.475 ;
        RECT 31.880 208.385 33.760 208.755 ;
        RECT 61.880 208.385 63.760 208.755 ;
        RECT 91.880 208.385 93.760 208.755 ;
        RECT 121.880 208.385 123.760 208.755 ;
        RECT 16.880 205.665 18.760 206.035 ;
        RECT 46.880 205.665 48.760 206.035 ;
        RECT 76.880 205.665 78.760 206.035 ;
        RECT 106.880 205.665 108.760 206.035 ;
        RECT 31.880 202.945 33.760 203.315 ;
        RECT 61.880 202.945 63.760 203.315 ;
        RECT 91.880 202.945 93.760 203.315 ;
        RECT 121.880 202.945 123.760 203.315 ;
        RECT 64.440 201.780 64.700 202.100 ;
        RECT 62.600 201.100 62.860 201.420 ;
        RECT 16.880 200.225 18.760 200.595 ;
        RECT 46.880 200.225 48.760 200.595 ;
        RECT 62.660 200.060 62.800 201.100 ;
        RECT 62.600 199.740 62.860 200.060 ;
        RECT 63.980 198.040 64.240 198.360 ;
        RECT 31.880 197.505 33.760 197.875 ;
        RECT 61.880 197.505 63.760 197.875 ;
        RECT 43.280 196.000 43.540 196.320 ;
        RECT 16.880 194.785 18.760 195.155 ;
        RECT 43.340 194.620 43.480 196.000 ;
        RECT 64.040 195.980 64.180 198.040 ;
        RECT 64.500 197.340 64.640 201.780 ;
        RECT 68.580 201.440 68.840 201.760 ;
        RECT 67.200 198.040 67.460 198.360 ;
        RECT 64.440 197.020 64.700 197.340 ;
        RECT 63.980 195.660 64.240 195.980 ;
        RECT 44.200 195.320 44.460 195.640 ;
        RECT 43.280 194.300 43.540 194.620 ;
        RECT 44.260 194.280 44.400 195.320 ;
        RECT 46.880 194.785 48.760 195.155 ;
        RECT 44.200 193.960 44.460 194.280 ;
        RECT 56.160 193.960 56.420 194.280 ;
        RECT 45.580 193.620 45.840 193.940 ;
        RECT 24.880 193.280 25.140 193.600 ;
        RECT 39.140 193.280 39.400 193.600 ;
        RECT 16.880 189.345 18.760 189.715 ;
        RECT 24.940 188.160 25.080 193.280 ;
        RECT 31.880 192.065 33.760 192.435 ;
        RECT 39.200 191.900 39.340 193.280 ;
        RECT 42.820 192.600 43.080 192.920 ;
        RECT 39.140 191.580 39.400 191.900 ;
        RECT 36.380 191.240 36.640 191.560 ;
        RECT 26.260 190.560 26.520 190.880 ;
        RECT 26.320 188.500 26.460 190.560 ;
        RECT 31.320 189.880 31.580 190.200 ;
        RECT 33.620 189.880 33.880 190.200 ;
        RECT 35.460 189.880 35.720 190.200 ;
        RECT 35.920 189.880 36.180 190.200 ;
        RECT 31.380 188.840 31.520 189.880 ;
        RECT 33.680 189.180 33.820 189.880 ;
        RECT 33.620 188.860 33.880 189.180 ;
        RECT 31.320 188.520 31.580 188.840 ;
        RECT 26.260 188.180 26.520 188.500 ;
        RECT 30.400 188.180 30.660 188.500 ;
        RECT 24.880 187.840 25.140 188.160 ;
        RECT 24.940 185.780 25.080 187.840 ;
        RECT 26.320 187.740 26.460 188.180 ;
        RECT 30.460 187.740 30.600 188.180 ;
        RECT 25.860 187.600 26.460 187.740 ;
        RECT 30.000 187.600 30.600 187.740 ;
        RECT 24.880 185.690 25.140 185.780 ;
        RECT 24.480 185.550 25.140 185.690 ;
        RECT 16.880 183.905 18.760 184.275 ;
        RECT 16.880 178.465 18.760 178.835 ;
        RECT 23.960 177.640 24.220 177.960 ;
        RECT 24.020 175.580 24.160 177.640 ;
        RECT 24.480 177.280 24.620 185.550 ;
        RECT 24.880 185.460 25.140 185.550 ;
        RECT 25.860 180.000 26.000 187.600 ;
        RECT 30.000 185.100 30.140 187.600 ;
        RECT 31.880 186.625 33.760 186.995 ;
        RECT 26.260 184.780 26.520 185.100 ;
        RECT 29.940 184.780 30.200 185.100 ;
        RECT 26.320 183.740 26.460 184.780 ;
        RECT 35.520 184.760 35.660 189.880 ;
        RECT 35.980 187.480 36.120 189.880 ;
        RECT 35.920 187.160 36.180 187.480 ;
        RECT 34.080 184.440 34.340 184.760 ;
        RECT 35.460 184.440 35.720 184.760 ;
        RECT 26.260 183.420 26.520 183.740 ;
        RECT 34.140 183.060 34.280 184.440 ;
        RECT 30.860 182.740 31.120 183.060 ;
        RECT 34.080 182.740 34.340 183.060 ;
        RECT 25.800 179.680 26.060 180.000 ;
        RECT 24.420 176.960 24.680 177.280 ;
        RECT 23.960 175.260 24.220 175.580 ;
        RECT 24.480 174.900 24.620 176.960 ;
        RECT 24.420 174.580 24.680 174.900 ;
        RECT 23.960 174.240 24.220 174.560 ;
        RECT 16.880 173.025 18.760 173.395 ;
        RECT 16.880 167.585 18.760 167.955 ;
        RECT 19.360 166.760 19.620 167.080 ;
        RECT 19.420 164.700 19.560 166.760 ;
        RECT 19.820 166.080 20.080 166.400 ;
        RECT 19.360 164.380 19.620 164.700 ;
        RECT 18.900 163.360 19.160 163.680 ;
        RECT 16.880 162.145 18.760 162.515 ;
        RECT 18.960 161.300 19.100 163.360 ;
        RECT 18.900 160.980 19.160 161.300 ;
        RECT 19.880 159.260 20.020 166.080 ;
        RECT 24.020 165.720 24.160 174.240 ;
        RECT 24.480 172.180 24.620 174.580 ;
        RECT 25.860 174.560 26.000 179.680 ;
        RECT 30.920 178.300 31.060 182.740 ;
        RECT 31.880 181.185 33.760 181.555 ;
        RECT 30.860 177.980 31.120 178.300 ;
        RECT 26.260 177.640 26.520 177.960 ;
        RECT 30.400 177.640 30.660 177.960 ;
        RECT 26.320 175.240 26.460 177.640 ;
        RECT 26.260 174.920 26.520 175.240 ;
        RECT 25.800 174.240 26.060 174.560 ;
        RECT 26.720 174.240 26.980 174.560 ;
        RECT 26.780 172.860 26.920 174.240 ;
        RECT 26.720 172.540 26.980 172.860 ;
        RECT 24.420 171.860 24.680 172.180 ;
        RECT 24.480 169.460 24.620 171.860 ;
        RECT 24.420 169.140 24.680 169.460 ;
        RECT 24.480 166.400 24.620 169.140 ;
        RECT 30.460 169.120 30.600 177.640 ;
        RECT 30.860 176.620 31.120 176.940 ;
        RECT 30.400 168.800 30.660 169.120 ;
        RECT 24.420 166.080 24.680 166.400 ;
        RECT 22.580 165.400 22.840 165.720 ;
        RECT 23.960 165.400 24.220 165.720 ;
        RECT 22.120 163.700 22.380 164.020 ;
        RECT 21.660 163.020 21.920 163.340 ;
        RECT 21.720 161.980 21.860 163.020 ;
        RECT 21.660 161.660 21.920 161.980 ;
        RECT 20.740 160.980 21.000 161.300 ;
        RECT 19.820 158.940 20.080 159.260 ;
        RECT 20.800 158.240 20.940 160.980 ;
        RECT 22.180 158.580 22.320 163.700 ;
        RECT 22.640 163.000 22.780 165.400 ;
        RECT 24.480 163.000 24.620 166.080 ;
        RECT 28.560 165.400 28.820 165.720 ;
        RECT 25.340 164.040 25.600 164.360 ;
        RECT 22.580 162.680 22.840 163.000 ;
        RECT 24.420 162.680 24.680 163.000 ;
        RECT 22.120 158.260 22.380 158.580 ;
        RECT 20.740 157.920 21.000 158.240 ;
        RECT 16.880 156.705 18.760 157.075 ;
        RECT 19.360 155.880 19.620 156.200 ;
        RECT 16.880 151.265 18.760 151.635 ;
        RECT 19.420 151.100 19.560 155.880 ;
        RECT 19.360 150.780 19.620 151.100 ;
        RECT 20.800 150.420 20.940 157.920 ;
        RECT 21.660 157.240 21.920 157.560 ;
        RECT 21.720 154.840 21.860 157.240 ;
        RECT 21.660 154.520 21.920 154.840 ;
        RECT 21.720 152.120 21.860 154.520 ;
        RECT 22.180 153.480 22.320 158.260 ;
        RECT 22.640 157.560 22.780 162.680 ;
        RECT 24.480 160.960 24.620 162.680 ;
        RECT 25.400 161.300 25.540 164.040 ;
        RECT 28.620 163.680 28.760 165.400 ;
        RECT 28.560 163.360 28.820 163.680 ;
        RECT 25.340 160.980 25.600 161.300 ;
        RECT 24.420 160.640 24.680 160.960 ;
        RECT 26.260 160.640 26.520 160.960 ;
        RECT 22.580 157.240 22.840 157.560 ;
        RECT 26.320 155.520 26.460 160.640 ;
        RECT 24.420 155.200 24.680 155.520 ;
        RECT 26.260 155.200 26.520 155.520 ;
        RECT 29.020 155.200 29.280 155.520 ;
        RECT 22.120 153.160 22.380 153.480 ;
        RECT 22.120 152.140 22.380 152.460 ;
        RECT 21.660 151.800 21.920 152.120 ;
        RECT 20.740 150.100 21.000 150.420 ;
        RECT 21.720 149.400 21.860 151.800 ;
        RECT 22.180 150.080 22.320 152.140 ;
        RECT 23.960 151.800 24.220 152.120 ;
        RECT 22.120 149.760 22.380 150.080 ;
        RECT 21.660 149.080 21.920 149.400 ;
        RECT 24.020 147.360 24.160 151.800 ;
        RECT 24.480 148.380 24.620 155.200 ;
        RECT 28.560 151.800 28.820 152.120 ;
        RECT 28.620 150.760 28.760 151.800 ;
        RECT 28.560 150.440 28.820 150.760 ;
        RECT 29.080 150.420 29.220 155.200 ;
        RECT 30.400 151.800 30.660 152.120 ;
        RECT 30.460 150.420 30.600 151.800 ;
        RECT 29.020 150.100 29.280 150.420 ;
        RECT 30.400 150.100 30.660 150.420 ;
        RECT 24.420 148.060 24.680 148.380 ;
        RECT 23.960 147.040 24.220 147.360 ;
        RECT 27.640 146.360 27.900 146.680 ;
        RECT 16.880 145.825 18.760 146.195 ;
        RECT 18.900 145.000 19.160 145.320 ;
        RECT 16.880 140.385 18.760 140.755 ;
        RECT 18.960 137.500 19.100 145.000 ;
        RECT 21.200 144.320 21.460 144.640 ;
        RECT 25.340 144.320 25.600 144.640 ;
        RECT 20.740 141.600 21.000 141.920 ;
        RECT 19.360 139.560 19.620 139.880 ;
        RECT 19.420 137.500 19.560 139.560 ;
        RECT 18.900 137.180 19.160 137.500 ;
        RECT 19.360 137.180 19.620 137.500 ;
        RECT 16.880 134.945 18.760 135.315 ;
        RECT 20.800 133.760 20.940 141.600 ;
        RECT 21.260 134.780 21.400 144.320 ;
        RECT 21.660 143.640 21.920 143.960 ;
        RECT 21.720 140.220 21.860 143.640 ;
        RECT 21.660 139.900 21.920 140.220 ;
        RECT 21.720 136.820 21.860 139.900 ;
        RECT 25.400 139.540 25.540 144.320 ;
        RECT 25.340 139.220 25.600 139.540 ;
        RECT 24.880 138.880 25.140 139.200 ;
        RECT 22.120 138.200 22.380 138.520 ;
        RECT 21.660 136.500 21.920 136.820 ;
        RECT 21.720 134.780 21.860 136.500 ;
        RECT 22.180 136.480 22.320 138.200 ;
        RECT 24.940 137.500 25.080 138.880 ;
        RECT 24.880 137.180 25.140 137.500 ;
        RECT 23.040 136.500 23.300 136.820 ;
        RECT 22.120 136.160 22.380 136.480 ;
        RECT 21.200 134.460 21.460 134.780 ;
        RECT 21.660 134.460 21.920 134.780 ;
        RECT 23.100 133.760 23.240 136.500 ;
        RECT 25.400 133.760 25.540 139.220 ;
        RECT 26.260 137.180 26.520 137.500 ;
        RECT 26.320 136.820 26.460 137.180 ;
        RECT 26.260 136.500 26.520 136.820 ;
        RECT 25.800 136.160 26.060 136.480 ;
        RECT 25.860 135.800 26.000 136.160 ;
        RECT 25.800 135.480 26.060 135.800 ;
        RECT 27.180 135.480 27.440 135.800 ;
        RECT 27.240 134.440 27.380 135.480 ;
        RECT 27.180 134.120 27.440 134.440 ;
        RECT 20.740 133.440 21.000 133.760 ;
        RECT 22.120 133.440 22.380 133.760 ;
        RECT 23.040 133.440 23.300 133.760 ;
        RECT 25.340 133.440 25.600 133.760 ;
        RECT 16.880 129.505 18.760 129.875 ;
        RECT 18.900 128.680 19.160 129.000 ;
        RECT 16.880 124.065 18.760 124.435 ;
        RECT 18.960 120.840 19.100 128.680 ;
        RECT 21.660 127.320 21.920 127.640 ;
        RECT 19.360 123.240 19.620 123.560 ;
        RECT 19.420 121.180 19.560 123.240 ;
        RECT 19.360 120.860 19.620 121.180 ;
        RECT 18.900 120.520 19.160 120.840 ;
        RECT 21.720 120.500 21.860 127.320 ;
        RECT 21.660 120.180 21.920 120.500 ;
        RECT 22.180 119.480 22.320 133.440 ;
        RECT 25.400 128.660 25.540 133.440 ;
        RECT 23.040 128.340 23.300 128.660 ;
        RECT 25.340 128.340 25.600 128.660 ;
        RECT 23.100 123.900 23.240 128.340 ;
        RECT 25.400 125.940 25.540 128.340 ;
        RECT 25.340 125.620 25.600 125.940 ;
        RECT 23.040 123.580 23.300 123.900 ;
        RECT 24.880 122.900 25.140 123.220 ;
        RECT 24.940 121.180 25.080 122.900 ;
        RECT 25.340 121.880 25.600 122.200 ;
        RECT 26.720 121.880 26.980 122.200 ;
        RECT 25.400 121.180 25.540 121.880 ;
        RECT 24.880 120.860 25.140 121.180 ;
        RECT 25.340 120.860 25.600 121.180 ;
        RECT 26.780 120.160 26.920 121.880 ;
        RECT 26.720 119.840 26.980 120.160 ;
        RECT 20.280 119.160 20.540 119.480 ;
        RECT 21.660 119.160 21.920 119.480 ;
        RECT 22.120 119.160 22.380 119.480 ;
        RECT 23.040 119.160 23.300 119.480 ;
        RECT 16.880 118.625 18.760 118.995 ;
        RECT 20.340 118.120 20.480 119.160 ;
        RECT 20.280 117.800 20.540 118.120 ;
        RECT 21.720 115.060 21.860 119.160 ;
        RECT 22.180 118.460 22.320 119.160 ;
        RECT 22.120 118.140 22.380 118.460 ;
        RECT 21.660 114.740 21.920 115.060 ;
        RECT 23.100 114.720 23.240 119.160 ;
        RECT 25.340 117.120 25.600 117.440 ;
        RECT 25.400 115.740 25.540 117.120 ;
        RECT 25.340 115.420 25.600 115.740 ;
        RECT 23.040 114.400 23.300 114.720 ;
        RECT 16.880 113.185 18.760 113.555 ;
        RECT 22.580 112.020 22.840 112.340 ;
        RECT 20.740 111.680 21.000 112.000 ;
        RECT 18.900 108.960 19.160 109.280 ;
        RECT 16.880 107.745 18.760 108.115 ;
        RECT 18.960 106.900 19.100 108.960 ;
        RECT 18.900 106.580 19.160 106.900 ;
        RECT 17.980 105.560 18.240 105.880 ;
        RECT 18.040 103.500 18.180 105.560 ;
        RECT 17.980 103.180 18.240 103.500 ;
        RECT 14.300 102.840 14.560 103.160 ;
        RECT 14.360 89.420 14.500 102.840 ;
        RECT 16.880 102.305 18.760 102.675 ;
        RECT 20.800 89.850 20.940 111.680 ;
        RECT 22.640 110.300 22.780 112.020 ;
        RECT 22.580 109.980 22.840 110.300 ;
        RECT 27.700 109.280 27.840 146.360 ;
        RECT 30.920 144.640 31.060 176.620 ;
        RECT 31.320 176.280 31.580 176.600 ;
        RECT 31.380 174.900 31.520 176.280 ;
        RECT 31.880 175.745 33.760 176.115 ;
        RECT 31.320 174.580 31.580 174.900 ;
        RECT 34.140 171.500 34.280 182.740 ;
        RECT 36.440 182.720 36.580 191.240 ;
        RECT 42.880 191.220 43.020 192.600 ;
        RECT 42.820 190.900 43.080 191.220 ;
        RECT 42.880 190.540 43.020 190.900 ;
        RECT 45.640 190.880 45.780 193.620 ;
        RECT 50.180 192.600 50.440 192.920 ;
        RECT 45.580 190.560 45.840 190.880 ;
        RECT 49.260 190.560 49.520 190.880 ;
        RECT 38.220 190.220 38.480 190.540 ;
        RECT 42.820 190.220 43.080 190.540 ;
        RECT 35.460 182.400 35.720 182.720 ;
        RECT 36.380 182.400 36.640 182.720 ;
        RECT 34.540 177.300 34.800 177.620 ;
        RECT 34.600 172.860 34.740 177.300 ;
        RECT 35.520 174.900 35.660 182.400 ;
        RECT 35.920 177.640 36.180 177.960 ;
        RECT 35.460 174.580 35.720 174.900 ;
        RECT 35.000 173.560 35.260 173.880 ;
        RECT 34.540 172.540 34.800 172.860 ;
        RECT 35.060 172.180 35.200 173.560 ;
        RECT 35.000 171.860 35.260 172.180 ;
        RECT 34.080 171.180 34.340 171.500 ;
        RECT 31.880 170.305 33.760 170.675 ;
        RECT 35.060 169.120 35.200 171.860 ;
        RECT 35.520 171.840 35.660 174.580 ;
        RECT 35.980 171.840 36.120 177.640 ;
        RECT 36.380 176.960 36.640 177.280 ;
        RECT 36.440 175.580 36.580 176.960 ;
        RECT 36.380 175.260 36.640 175.580 ;
        RECT 36.370 174.045 36.650 174.415 ;
        RECT 35.460 171.520 35.720 171.840 ;
        RECT 35.920 171.520 36.180 171.840 ;
        RECT 35.000 168.800 35.260 169.120 ;
        RECT 35.460 169.030 35.720 169.120 ;
        RECT 35.980 169.030 36.120 171.520 ;
        RECT 35.460 168.890 36.120 169.030 ;
        RECT 35.460 168.800 35.720 168.890 ;
        RECT 36.440 168.780 36.580 174.045 ;
        RECT 38.280 172.520 38.420 190.220 ;
        RECT 40.060 187.160 40.320 187.480 ;
        RECT 40.120 183.400 40.260 187.160 ;
        RECT 40.060 183.080 40.320 183.400 ;
        RECT 41.440 182.060 41.700 182.380 ;
        RECT 39.140 172.540 39.400 172.860 ;
        RECT 38.220 172.200 38.480 172.520 ;
        RECT 39.200 172.180 39.340 172.540 ;
        RECT 39.140 171.860 39.400 172.180 ;
        RECT 40.980 171.860 41.240 172.180 ;
        RECT 37.300 170.840 37.560 171.160 ;
        RECT 36.380 168.460 36.640 168.780 ;
        RECT 36.840 168.180 37.100 168.440 ;
        RECT 36.440 168.120 37.100 168.180 ;
        RECT 36.440 168.040 37.040 168.120 ;
        RECT 31.880 164.865 33.760 165.235 ;
        RECT 35.460 164.380 35.720 164.700 ;
        RECT 35.520 164.020 35.660 164.380 ;
        RECT 35.000 163.700 35.260 164.020 ;
        RECT 35.460 163.700 35.720 164.020 ;
        RECT 31.320 161.320 31.580 161.640 ;
        RECT 31.380 159.260 31.520 161.320 ;
        RECT 31.880 159.425 33.760 159.795 ;
        RECT 31.320 158.940 31.580 159.260 ;
        RECT 31.780 157.920 32.040 158.240 ;
        RECT 31.320 157.240 31.580 157.560 ;
        RECT 31.380 152.710 31.520 157.240 ;
        RECT 31.840 155.520 31.980 157.920 ;
        RECT 35.060 157.900 35.200 163.700 ;
        RECT 35.000 157.580 35.260 157.900 ;
        RECT 31.780 155.200 32.040 155.520 ;
        RECT 31.880 153.985 33.760 154.355 ;
        RECT 35.520 153.140 35.660 163.700 ;
        RECT 35.920 159.960 36.180 160.280 ;
        RECT 35.980 157.560 36.120 159.960 ;
        RECT 35.920 157.240 36.180 157.560 ;
        RECT 35.460 152.820 35.720 153.140 ;
        RECT 32.240 152.710 32.500 152.800 ;
        RECT 31.380 152.570 32.500 152.710 ;
        RECT 32.240 152.480 32.500 152.570 ;
        RECT 32.700 152.480 32.960 152.800 ;
        RECT 32.760 151.100 32.900 152.480 ;
        RECT 33.620 152.140 33.880 152.460 ;
        RECT 32.700 150.780 32.960 151.100 ;
        RECT 33.680 150.420 33.820 152.140 ;
        RECT 34.080 151.800 34.340 152.120 ;
        RECT 35.000 151.800 35.260 152.120 ;
        RECT 33.620 150.100 33.880 150.420 ;
        RECT 31.880 148.545 33.760 148.915 ;
        RECT 34.140 144.980 34.280 151.800 ;
        RECT 35.060 147.360 35.200 151.800 ;
        RECT 35.520 149.740 35.660 152.820 ;
        RECT 35.460 149.420 35.720 149.740 ;
        RECT 35.920 149.080 36.180 149.400 ;
        RECT 35.460 148.060 35.720 148.380 ;
        RECT 35.000 147.040 35.260 147.360 ;
        RECT 35.000 146.360 35.260 146.680 ;
        RECT 34.080 144.660 34.340 144.980 ;
        RECT 30.860 144.320 31.120 144.640 ;
        RECT 30.400 143.640 30.660 143.960 ;
        RECT 34.080 143.640 34.340 143.960 ;
        RECT 29.940 138.540 30.200 138.860 ;
        RECT 30.000 135.800 30.140 138.540 ;
        RECT 29.940 135.480 30.200 135.800 ;
        RECT 30.000 134.780 30.140 135.480 ;
        RECT 29.940 134.460 30.200 134.780 ;
        RECT 30.000 130.700 30.140 134.460 ;
        RECT 30.460 131.460 30.600 143.640 ;
        RECT 31.880 143.105 33.760 143.475 ;
        RECT 33.160 141.600 33.420 141.920 ;
        RECT 33.220 139.540 33.360 141.600 ;
        RECT 34.140 140.220 34.280 143.640 ;
        RECT 34.540 140.920 34.800 141.240 ;
        RECT 34.080 139.900 34.340 140.220 ;
        RECT 33.160 139.220 33.420 139.540 ;
        RECT 31.880 137.665 33.760 138.035 ;
        RECT 31.780 136.160 32.040 136.480 ;
        RECT 31.320 135.480 31.580 135.800 ;
        RECT 30.860 133.780 31.120 134.100 ;
        RECT 30.920 132.060 31.060 133.780 ;
        RECT 30.860 131.740 31.120 132.060 ;
        RECT 30.460 131.320 31.060 131.460 ;
        RECT 29.940 130.380 30.200 130.700 ;
        RECT 29.480 125.280 29.740 125.600 ;
        RECT 29.940 125.280 30.200 125.600 ;
        RECT 28.100 122.560 28.360 122.880 ;
        RECT 28.160 120.500 28.300 122.560 ;
        RECT 28.100 120.180 28.360 120.500 ;
        RECT 28.560 119.500 28.820 119.820 ;
        RECT 28.620 115.740 28.760 119.500 ;
        RECT 29.540 115.740 29.680 125.280 ;
        RECT 30.000 120.500 30.140 125.280 ;
        RECT 30.400 124.600 30.660 124.920 ;
        RECT 30.460 123.220 30.600 124.600 ;
        RECT 30.400 122.900 30.660 123.220 ;
        RECT 29.940 120.180 30.200 120.500 ;
        RECT 30.000 118.460 30.140 120.180 ;
        RECT 30.400 119.160 30.660 119.480 ;
        RECT 29.940 118.140 30.200 118.460 ;
        RECT 28.560 115.420 28.820 115.740 ;
        RECT 29.480 115.420 29.740 115.740 ;
        RECT 30.000 112.340 30.140 118.140 ;
        RECT 30.460 115.060 30.600 119.160 ;
        RECT 30.400 114.740 30.660 115.060 ;
        RECT 29.940 112.020 30.200 112.340 ;
        RECT 29.020 111.000 29.280 111.320 ;
        RECT 29.080 109.960 29.220 111.000 ;
        RECT 29.020 109.640 29.280 109.960 ;
        RECT 27.640 108.960 27.900 109.280 ;
        RECT 25.800 108.280 26.060 108.600 ;
        RECT 28.560 108.280 28.820 108.600 ;
        RECT 25.860 107.240 26.000 108.280 ;
        RECT 25.800 106.920 26.060 107.240 ;
        RECT 26.260 105.560 26.520 105.880 ;
        RECT 13.920 85.550 15.140 89.420 ;
        RECT 19.910 85.980 21.130 89.850 ;
        RECT 26.320 89.170 26.460 105.560 ;
        RECT 28.620 104.180 28.760 108.280 ;
        RECT 30.000 106.300 30.140 112.020 ;
        RECT 30.920 109.280 31.060 131.320 ;
        RECT 31.380 131.040 31.520 135.480 ;
        RECT 31.840 134.100 31.980 136.160 ;
        RECT 31.780 133.780 32.040 134.100 ;
        RECT 31.880 132.225 33.760 132.595 ;
        RECT 31.320 130.720 31.580 131.040 ;
        RECT 31.880 126.785 33.760 127.155 ;
        RECT 32.700 125.280 32.960 125.600 ;
        RECT 32.760 123.220 32.900 125.280 ;
        RECT 32.700 122.900 32.960 123.220 ;
        RECT 34.080 121.880 34.340 122.200 ;
        RECT 31.880 121.345 33.760 121.715 ;
        RECT 31.320 120.860 31.580 121.180 ;
        RECT 31.380 114.720 31.520 120.860 ;
        RECT 31.880 115.905 33.760 116.275 ;
        RECT 34.140 114.720 34.280 121.880 ;
        RECT 31.320 114.400 31.580 114.720 ;
        RECT 34.080 114.400 34.340 114.720 ;
        RECT 31.880 110.465 33.760 110.835 ;
        RECT 34.600 109.280 34.740 140.920 ;
        RECT 35.060 140.130 35.200 146.360 ;
        RECT 35.520 140.980 35.660 148.060 ;
        RECT 35.980 141.920 36.120 149.080 ;
        RECT 36.440 142.260 36.580 168.040 ;
        RECT 36.840 157.240 37.100 157.560 ;
        RECT 36.900 156.540 37.040 157.240 ;
        RECT 36.840 156.220 37.100 156.540 ;
        RECT 36.840 152.480 37.100 152.800 ;
        RECT 36.900 151.100 37.040 152.480 ;
        RECT 36.840 150.780 37.100 151.100 ;
        RECT 36.900 150.080 37.040 150.780 ;
        RECT 36.840 149.760 37.100 150.080 ;
        RECT 37.360 147.700 37.500 170.840 ;
        RECT 39.200 169.120 39.340 171.860 ;
        RECT 41.040 169.460 41.180 171.860 ;
        RECT 40.980 169.140 41.240 169.460 ;
        RECT 39.140 168.800 39.400 169.120 ;
        RECT 37.760 163.020 38.020 163.340 ;
        RECT 37.820 162.060 37.960 163.020 ;
        RECT 39.140 162.680 39.400 163.000 ;
        RECT 37.820 161.980 38.420 162.060 ;
        RECT 37.820 161.920 38.480 161.980 ;
        RECT 38.220 161.660 38.480 161.920 ;
        RECT 39.200 161.300 39.340 162.680 ;
        RECT 38.680 160.980 38.940 161.300 ;
        RECT 39.140 160.980 39.400 161.300 ;
        RECT 38.740 159.260 38.880 160.980 ;
        RECT 38.680 158.940 38.940 159.260 ;
        RECT 40.980 157.920 41.240 158.240 ;
        RECT 40.060 157.240 40.320 157.560 ;
        RECT 37.760 156.220 38.020 156.540 ;
        RECT 37.820 152.800 37.960 156.220 ;
        RECT 39.600 154.860 39.860 155.180 ;
        RECT 39.660 153.480 39.800 154.860 ;
        RECT 38.210 152.965 38.490 153.335 ;
        RECT 39.600 153.160 39.860 153.480 ;
        RECT 38.280 152.800 38.420 152.965 ;
        RECT 37.760 152.480 38.020 152.800 ;
        RECT 38.220 152.480 38.480 152.800 ;
        RECT 37.760 152.030 38.020 152.120 ;
        RECT 38.280 152.030 38.420 152.480 ;
        RECT 37.760 151.890 38.420 152.030 ;
        RECT 37.760 151.800 38.020 151.890 ;
        RECT 39.660 150.420 39.800 153.160 ;
        RECT 39.600 150.100 39.860 150.420 ;
        RECT 38.680 149.080 38.940 149.400 ;
        RECT 37.300 147.380 37.560 147.700 ;
        RECT 36.840 144.660 37.100 144.980 ;
        RECT 36.900 142.600 37.040 144.660 ;
        RECT 36.840 142.280 37.100 142.600 ;
        RECT 36.380 141.940 36.640 142.260 ;
        RECT 35.920 141.600 36.180 141.920 ;
        RECT 35.520 140.840 36.580 140.980 ;
        RECT 36.440 140.220 36.580 140.840 ;
        RECT 35.060 139.990 35.660 140.130 ;
        RECT 35.000 139.220 35.260 139.540 ;
        RECT 35.060 138.520 35.200 139.220 ;
        RECT 35.000 138.200 35.260 138.520 ;
        RECT 35.060 136.820 35.200 138.200 ;
        RECT 35.000 136.500 35.260 136.820 ;
        RECT 35.000 122.900 35.260 123.220 ;
        RECT 35.060 119.480 35.200 122.900 ;
        RECT 35.000 119.160 35.260 119.480 ;
        RECT 35.520 111.840 35.660 139.990 ;
        RECT 36.380 139.900 36.640 140.220 ;
        RECT 36.380 139.220 36.640 139.540 ;
        RECT 35.920 135.820 36.180 136.140 ;
        RECT 35.980 134.780 36.120 135.820 ;
        RECT 35.920 134.460 36.180 134.780 ;
        RECT 36.440 133.420 36.580 139.220 ;
        RECT 37.300 136.500 37.560 136.820 ;
        RECT 36.840 135.480 37.100 135.800 ;
        RECT 36.380 133.100 36.640 133.420 ;
        RECT 36.900 131.040 37.040 135.480 ;
        RECT 37.360 131.380 37.500 136.500 ;
        RECT 37.760 133.780 38.020 134.100 ;
        RECT 38.220 133.780 38.480 134.100 ;
        RECT 37.300 131.060 37.560 131.380 ;
        RECT 36.840 130.720 37.100 131.040 ;
        RECT 37.360 129.000 37.500 131.060 ;
        RECT 37.820 131.040 37.960 133.780 ;
        RECT 38.280 132.060 38.420 133.780 ;
        RECT 38.220 131.740 38.480 132.060 ;
        RECT 37.760 130.720 38.020 131.040 ;
        RECT 37.300 128.680 37.560 129.000 ;
        RECT 37.360 123.980 37.500 128.680 ;
        RECT 38.740 125.600 38.880 149.080 ;
        RECT 39.140 148.060 39.400 148.380 ;
        RECT 39.200 139.200 39.340 148.060 ;
        RECT 40.120 147.700 40.260 157.240 ;
        RECT 41.040 153.140 41.180 157.920 ;
        RECT 40.980 152.820 41.240 153.140 ;
        RECT 40.520 150.780 40.780 151.100 ;
        RECT 40.060 147.380 40.320 147.700 ;
        RECT 40.580 147.100 40.720 150.780 ;
        RECT 41.500 149.820 41.640 182.060 ;
        RECT 42.880 177.620 43.020 190.220 ;
        RECT 44.660 189.880 44.920 190.200 ;
        RECT 44.720 188.840 44.860 189.880 ;
        RECT 44.660 188.520 44.920 188.840 ;
        RECT 45.640 185.100 45.780 190.560 ;
        RECT 46.500 189.880 46.760 190.200 ;
        RECT 46.560 189.180 46.700 189.880 ;
        RECT 46.880 189.345 48.760 189.715 ;
        RECT 46.500 188.860 46.760 189.180 ;
        RECT 48.800 187.160 49.060 187.480 ;
        RECT 48.860 185.860 49.000 187.160 ;
        RECT 49.320 186.460 49.460 190.560 ;
        RECT 50.240 190.200 50.380 192.600 ;
        RECT 56.220 191.900 56.360 193.960 ;
        RECT 58.000 193.280 58.260 193.600 ;
        RECT 56.160 191.580 56.420 191.900 ;
        RECT 50.640 190.900 50.900 191.220 ;
        RECT 50.180 189.880 50.440 190.200 ;
        RECT 49.260 186.140 49.520 186.460 ;
        RECT 48.860 185.720 49.460 185.860 ;
        RECT 49.320 185.440 49.460 185.720 ;
        RECT 46.040 185.120 46.300 185.440 ;
        RECT 49.260 185.120 49.520 185.440 ;
        RECT 45.580 184.780 45.840 185.100 ;
        RECT 45.120 182.740 45.380 183.060 ;
        RECT 43.740 182.400 44.000 182.720 ;
        RECT 43.800 179.320 43.940 182.400 ;
        RECT 43.740 179.000 44.000 179.320 ;
        RECT 43.280 177.980 43.540 178.300 ;
        RECT 42.820 177.300 43.080 177.620 ;
        RECT 42.820 173.900 43.080 174.220 ;
        RECT 42.880 171.580 43.020 173.900 ;
        RECT 43.340 172.860 43.480 177.980 ;
        RECT 43.800 174.560 43.940 179.000 ;
        RECT 45.180 177.620 45.320 182.740 ;
        RECT 44.200 177.300 44.460 177.620 ;
        RECT 45.120 177.300 45.380 177.620 ;
        RECT 45.580 177.300 45.840 177.620 ;
        RECT 44.260 174.980 44.400 177.300 ;
        RECT 44.660 176.960 44.920 177.280 ;
        RECT 44.720 175.580 44.860 176.960 ;
        RECT 45.120 176.280 45.380 176.600 ;
        RECT 44.660 175.260 44.920 175.580 ;
        RECT 44.260 174.840 44.860 174.980 ;
        RECT 43.740 174.300 44.000 174.560 ;
        RECT 43.740 174.240 44.400 174.300 ;
        RECT 43.800 174.160 44.400 174.240 ;
        RECT 43.280 172.540 43.540 172.860 ;
        RECT 43.340 172.180 43.480 172.540 ;
        RECT 44.260 172.180 44.400 174.160 ;
        RECT 44.720 173.880 44.860 174.840 ;
        RECT 44.660 173.560 44.920 173.880 ;
        RECT 44.720 172.860 44.860 173.560 ;
        RECT 44.660 172.540 44.920 172.860 ;
        RECT 43.280 171.860 43.540 172.180 ;
        RECT 44.200 171.860 44.460 172.180 ;
        RECT 42.880 171.440 44.860 171.580 ;
        RECT 41.900 170.840 42.160 171.160 ;
        RECT 41.960 151.100 42.100 170.840 ;
        RECT 43.280 169.140 43.540 169.460 ;
        RECT 43.340 164.700 43.480 169.140 ;
        RECT 44.200 165.400 44.460 165.720 ;
        RECT 43.280 164.380 43.540 164.700 ;
        RECT 43.340 158.240 43.480 164.380 ;
        RECT 44.260 163.680 44.400 165.400 ;
        RECT 43.740 163.360 44.000 163.680 ;
        RECT 44.200 163.360 44.460 163.680 ;
        RECT 43.800 161.980 43.940 163.360 ;
        RECT 44.200 162.680 44.460 163.000 ;
        RECT 43.740 161.660 44.000 161.980 ;
        RECT 43.280 157.920 43.540 158.240 ;
        RECT 43.800 157.560 43.940 161.660 ;
        RECT 44.260 161.640 44.400 162.680 ;
        RECT 44.200 161.320 44.460 161.640 ;
        RECT 44.200 158.260 44.460 158.580 ;
        RECT 43.740 157.240 44.000 157.560 ;
        RECT 42.360 155.880 42.620 156.200 ;
        RECT 41.900 150.780 42.160 151.100 ;
        RECT 42.420 150.420 42.560 155.880 ;
        RECT 43.280 152.820 43.540 153.140 ;
        RECT 42.820 152.480 43.080 152.800 ;
        RECT 42.880 150.760 43.020 152.480 ;
        RECT 42.820 150.440 43.080 150.760 ;
        RECT 43.340 150.420 43.480 152.820 ;
        RECT 43.800 152.800 43.940 157.240 ;
        RECT 44.260 153.820 44.400 158.260 ;
        RECT 44.200 153.500 44.460 153.820 ;
        RECT 44.260 152.800 44.400 153.500 ;
        RECT 43.740 152.480 44.000 152.800 ;
        RECT 44.200 152.480 44.460 152.800 ;
        RECT 43.740 151.800 44.000 152.120 ;
        RECT 42.360 150.100 42.620 150.420 ;
        RECT 43.280 150.100 43.540 150.420 ;
        RECT 41.500 149.680 43.020 149.820 ;
        RECT 43.800 149.740 43.940 151.800 ;
        RECT 44.190 151.605 44.470 151.975 ;
        RECT 41.900 149.080 42.160 149.400 ;
        RECT 40.120 146.960 40.720 147.100 ;
        RECT 39.140 138.880 39.400 139.200 ;
        RECT 39.140 136.160 39.400 136.480 ;
        RECT 39.200 134.780 39.340 136.160 ;
        RECT 39.140 134.460 39.400 134.780 ;
        RECT 39.140 130.720 39.400 131.040 ;
        RECT 38.680 125.280 38.940 125.600 ;
        RECT 38.220 124.600 38.480 124.920 ;
        RECT 36.900 123.840 37.500 123.980 ;
        RECT 36.900 122.880 37.040 123.840 ;
        RECT 37.300 122.900 37.560 123.220 ;
        RECT 36.840 122.560 37.100 122.880 ;
        RECT 36.900 120.500 37.040 122.560 ;
        RECT 36.380 120.410 36.640 120.500 ;
        RECT 35.980 120.270 36.640 120.410 ;
        RECT 35.980 115.740 36.120 120.270 ;
        RECT 36.380 120.180 36.640 120.270 ;
        RECT 36.840 120.180 37.100 120.500 ;
        RECT 36.370 119.645 36.650 120.015 ;
        RECT 36.440 118.120 36.580 119.645 ;
        RECT 36.380 117.800 36.640 118.120 ;
        RECT 36.900 117.180 37.040 120.180 ;
        RECT 37.360 119.730 37.500 122.900 ;
        RECT 37.760 119.730 38.020 119.820 ;
        RECT 37.360 119.590 38.020 119.730 ;
        RECT 37.360 118.460 37.500 119.590 ;
        RECT 37.760 119.500 38.020 119.590 ;
        RECT 37.300 118.140 37.560 118.460 ;
        RECT 36.440 117.040 37.040 117.180 ;
        RECT 35.920 115.420 36.180 115.740 ;
        RECT 36.440 115.060 36.580 117.040 ;
        RECT 36.840 116.440 37.100 116.760 ;
        RECT 36.380 114.740 36.640 115.060 ;
        RECT 36.900 114.720 37.040 116.440 ;
        RECT 36.840 114.400 37.100 114.720 ;
        RECT 38.280 112.340 38.420 124.600 ;
        RECT 39.200 116.760 39.340 130.720 ;
        RECT 39.600 126.300 39.860 126.620 ;
        RECT 39.660 123.900 39.800 126.300 ;
        RECT 40.120 125.600 40.260 146.960 ;
        RECT 41.440 136.160 41.700 136.480 ;
        RECT 41.500 133.760 41.640 136.160 ;
        RECT 41.440 133.440 41.700 133.760 ;
        RECT 41.440 132.760 41.700 133.080 ;
        RECT 40.060 125.280 40.320 125.600 ;
        RECT 40.520 124.940 40.780 125.260 ;
        RECT 39.600 123.580 39.860 123.900 ;
        RECT 40.060 123.580 40.320 123.900 ;
        RECT 39.600 123.130 39.860 123.220 ;
        RECT 40.120 123.130 40.260 123.580 ;
        RECT 39.600 122.990 40.260 123.130 ;
        RECT 39.600 122.900 39.860 122.990 ;
        RECT 40.580 121.180 40.720 124.940 ;
        RECT 40.980 124.600 41.240 124.920 ;
        RECT 40.520 120.860 40.780 121.180 ;
        RECT 40.060 117.800 40.320 118.120 ;
        RECT 39.140 116.440 39.400 116.760 ;
        RECT 40.120 115.740 40.260 117.800 ;
        RECT 40.060 115.420 40.320 115.740 ;
        RECT 38.220 112.020 38.480 112.340 ;
        RECT 35.060 111.700 35.660 111.840 ;
        RECT 35.060 109.620 35.200 111.700 ;
        RECT 41.040 110.300 41.180 124.600 ;
        RECT 41.500 120.160 41.640 132.760 ;
        RECT 41.960 125.600 42.100 149.080 ;
        RECT 42.360 138.880 42.620 139.200 ;
        RECT 42.420 136.480 42.560 138.880 ;
        RECT 42.360 136.160 42.620 136.480 ;
        RECT 42.420 133.080 42.560 136.160 ;
        RECT 42.360 132.760 42.620 133.080 ;
        RECT 42.360 125.960 42.620 126.280 ;
        RECT 41.900 125.280 42.160 125.600 ;
        RECT 42.420 123.900 42.560 125.960 ;
        RECT 42.880 125.600 43.020 149.680 ;
        RECT 43.740 149.420 44.000 149.740 ;
        RECT 44.260 147.360 44.400 151.605 ;
        RECT 44.200 147.040 44.460 147.360 ;
        RECT 43.280 134.120 43.540 134.440 ;
        RECT 43.340 132.060 43.480 134.120 ;
        RECT 43.280 131.740 43.540 132.060 ;
        RECT 43.280 126.300 43.540 126.620 ;
        RECT 42.820 125.280 43.080 125.600 ;
        RECT 43.340 123.900 43.480 126.300 ;
        RECT 44.720 125.600 44.860 171.440 ;
        RECT 45.180 144.640 45.320 176.280 ;
        RECT 45.640 174.415 45.780 177.300 ;
        RECT 46.100 175.240 46.240 185.120 ;
        RECT 46.500 184.440 46.760 184.760 ;
        RECT 46.560 183.400 46.700 184.440 ;
        RECT 46.880 183.905 48.760 184.275 ;
        RECT 49.320 183.740 49.460 185.120 ;
        RECT 46.960 183.420 47.220 183.740 ;
        RECT 49.260 183.420 49.520 183.740 ;
        RECT 46.500 183.080 46.760 183.400 ;
        RECT 47.020 182.630 47.160 183.420 ;
        RECT 46.560 182.490 47.160 182.630 ;
        RECT 46.560 176.600 46.700 182.490 ;
        RECT 49.720 182.400 49.980 182.720 ;
        RECT 47.880 181.720 48.140 182.040 ;
        RECT 47.940 180.000 48.080 181.720 ;
        RECT 47.880 179.680 48.140 180.000 ;
        RECT 49.260 179.340 49.520 179.660 ;
        RECT 46.880 178.465 48.760 178.835 ;
        RECT 48.340 176.960 48.600 177.280 ;
        RECT 46.500 176.280 46.760 176.600 ;
        RECT 46.040 174.920 46.300 175.240 ;
        RECT 46.560 174.560 46.700 176.280 ;
        RECT 47.880 175.260 48.140 175.580 ;
        RECT 47.940 174.560 48.080 175.260 ;
        RECT 45.570 174.045 45.850 174.415 ;
        RECT 46.500 174.240 46.760 174.560 ;
        RECT 47.880 174.240 48.140 174.560 ;
        RECT 45.580 173.560 45.840 173.880 ;
        RECT 46.040 173.560 46.300 173.880 ;
        RECT 45.640 154.840 45.780 173.560 ;
        RECT 46.100 172.520 46.240 173.560 ;
        RECT 46.040 172.200 46.300 172.520 ;
        RECT 46.560 172.180 46.700 174.240 ;
        RECT 48.400 173.880 48.540 176.960 ;
        RECT 49.320 174.900 49.460 179.340 ;
        RECT 49.780 175.580 49.920 182.400 ;
        RECT 50.240 179.660 50.380 189.880 ;
        RECT 50.700 185.780 50.840 190.900 ;
        RECT 51.560 188.520 51.820 188.840 ;
        RECT 51.620 186.460 51.760 188.520 ;
        RECT 58.060 188.500 58.200 193.280 ;
        RECT 64.500 192.920 64.640 197.020 ;
        RECT 67.260 196.660 67.400 198.040 ;
        RECT 68.640 196.660 68.780 201.440 ;
        RECT 69.040 201.100 69.300 201.420 ;
        RECT 69.100 197.000 69.240 201.100 ;
        RECT 76.880 200.225 78.760 200.595 ;
        RECT 106.880 200.225 108.760 200.595 ;
        RECT 70.880 199.400 71.140 199.720 ;
        RECT 71.340 199.400 71.600 199.720 ;
        RECT 77.320 199.400 77.580 199.720 ;
        RECT 70.420 198.040 70.680 198.360 ;
        RECT 69.040 196.680 69.300 197.000 ;
        RECT 70.480 196.660 70.620 198.040 ;
        RECT 67.200 196.340 67.460 196.660 ;
        RECT 68.580 196.340 68.840 196.660 ;
        RECT 70.420 196.340 70.680 196.660 ;
        RECT 67.660 195.320 67.920 195.640 ;
        RECT 67.720 193.940 67.860 195.320 ;
        RECT 67.660 193.620 67.920 193.940 ;
        RECT 67.720 193.340 67.860 193.620 ;
        RECT 66.800 193.200 67.860 193.340 ;
        RECT 68.120 193.510 68.380 193.600 ;
        RECT 68.640 193.510 68.780 196.340 ;
        RECT 69.960 193.620 70.220 193.940 ;
        RECT 68.120 193.370 68.780 193.510 ;
        RECT 68.120 193.280 68.380 193.370 ;
        RECT 69.040 193.280 69.300 193.600 ;
        RECT 64.440 192.600 64.700 192.920 ;
        RECT 61.880 192.065 63.760 192.435 ;
        RECT 58.000 188.180 58.260 188.500 ;
        RECT 55.700 187.160 55.960 187.480 ;
        RECT 55.760 186.460 55.900 187.160 ;
        RECT 51.560 186.140 51.820 186.460 ;
        RECT 55.700 186.140 55.960 186.460 ;
        RECT 50.640 185.460 50.900 185.780 ;
        RECT 50.700 182.720 50.840 185.460 ;
        RECT 53.400 185.120 53.660 185.440 ;
        RECT 53.460 183.740 53.600 185.120 ;
        RECT 57.540 184.440 57.800 184.760 ;
        RECT 53.400 183.420 53.660 183.740 ;
        RECT 57.600 183.400 57.740 184.440 ;
        RECT 57.540 183.080 57.800 183.400 ;
        RECT 53.860 182.740 54.120 183.060 ;
        RECT 50.640 182.400 50.900 182.720 ;
        RECT 53.920 182.040 54.060 182.740 ;
        RECT 58.060 182.720 58.200 188.180 ;
        RECT 61.880 186.625 63.760 186.995 ;
        RECT 63.980 185.120 64.240 185.440 ;
        RECT 61.220 183.080 61.480 183.400 ;
        RECT 58.000 182.400 58.260 182.720 ;
        RECT 54.780 182.060 55.040 182.380 ;
        RECT 53.860 181.720 54.120 182.040 ;
        RECT 50.180 179.340 50.440 179.660 ;
        RECT 53.920 179.320 54.060 181.720 ;
        RECT 54.840 180.340 54.980 182.060 ;
        RECT 54.320 180.020 54.580 180.340 ;
        RECT 54.780 180.020 55.040 180.340 ;
        RECT 57.080 180.020 57.340 180.340 ;
        RECT 53.860 179.000 54.120 179.320 ;
        RECT 49.720 175.260 49.980 175.580 ;
        RECT 49.260 174.580 49.520 174.900 ;
        RECT 48.340 173.560 48.600 173.880 ;
        RECT 46.880 173.025 48.760 173.395 ;
        RECT 49.780 172.860 49.920 175.260 ;
        RECT 50.630 174.725 50.910 175.095 ;
        RECT 50.180 174.240 50.440 174.560 ;
        RECT 47.420 172.540 47.680 172.860 ;
        RECT 49.720 172.540 49.980 172.860 ;
        RECT 47.480 172.180 47.620 172.540 ;
        RECT 50.240 172.520 50.380 174.240 ;
        RECT 50.180 172.200 50.440 172.520 ;
        RECT 46.500 171.860 46.760 172.180 ;
        RECT 47.420 171.860 47.680 172.180 ;
        RECT 46.040 170.840 46.300 171.160 ;
        RECT 45.580 154.520 45.840 154.840 ;
        RECT 46.100 153.730 46.240 170.840 ;
        RECT 46.560 167.420 46.700 171.860 ;
        RECT 50.240 171.160 50.380 172.200 ;
        RECT 50.700 171.160 50.840 174.725 ;
        RECT 53.920 174.560 54.060 179.000 ;
        RECT 54.380 177.960 54.520 180.020 ;
        RECT 54.320 177.640 54.580 177.960 ;
        RECT 53.400 174.240 53.660 174.560 ;
        RECT 53.860 174.240 54.120 174.560 ;
        RECT 51.100 173.560 51.360 173.880 ;
        RECT 50.180 170.840 50.440 171.160 ;
        RECT 50.640 170.840 50.900 171.160 ;
        RECT 51.160 170.220 51.300 173.560 ;
        RECT 52.940 171.860 53.200 172.180 ;
        RECT 50.700 170.080 51.300 170.220 ;
        RECT 46.880 167.585 48.760 167.955 ;
        RECT 46.500 167.100 46.760 167.420 ;
        RECT 49.260 165.400 49.520 165.720 ;
        RECT 49.320 163.340 49.460 165.400 ;
        RECT 49.260 163.020 49.520 163.340 ;
        RECT 46.500 162.680 46.760 163.000 ;
        RECT 45.640 153.590 46.240 153.730 ;
        RECT 45.640 152.655 45.780 153.590 ;
        RECT 46.040 152.820 46.300 153.140 ;
        RECT 45.570 152.285 45.850 152.655 ;
        RECT 45.580 151.800 45.840 152.120 ;
        RECT 45.120 144.320 45.380 144.640 ;
        RECT 45.640 143.870 45.780 151.800 ;
        RECT 46.100 144.980 46.240 152.820 ;
        RECT 46.560 152.710 46.700 162.680 ;
        RECT 46.880 162.145 48.760 162.515 ;
        RECT 49.320 161.890 49.460 163.020 ;
        RECT 48.860 161.750 49.460 161.890 ;
        RECT 48.860 157.470 49.000 161.750 ;
        RECT 49.720 160.980 49.980 161.300 ;
        RECT 49.780 159.260 49.920 160.980 ;
        RECT 49.720 158.940 49.980 159.260 ;
        RECT 50.700 158.150 50.840 170.080 ;
        RECT 52.480 168.800 52.740 169.120 ;
        RECT 52.540 163.680 52.680 168.800 ;
        RECT 53.000 165.720 53.140 171.860 ;
        RECT 53.460 171.160 53.600 174.240 ;
        RECT 54.380 172.180 54.520 177.640 ;
        RECT 54.780 176.280 55.040 176.600 ;
        RECT 54.840 174.560 54.980 176.280 ;
        RECT 57.140 175.580 57.280 180.020 ;
        RECT 58.060 177.960 58.200 182.400 ;
        RECT 61.280 181.020 61.420 183.080 ;
        RECT 61.880 181.185 63.760 181.555 ;
        RECT 61.220 180.700 61.480 181.020 ;
        RECT 58.000 177.640 58.260 177.960 ;
        RECT 61.880 175.745 63.760 176.115 ;
        RECT 57.080 175.260 57.340 175.580 ;
        RECT 54.780 174.240 55.040 174.560 ;
        RECT 54.320 171.860 54.580 172.180 ;
        RECT 53.400 170.840 53.660 171.160 ;
        RECT 53.860 168.460 54.120 168.780 ;
        RECT 52.940 165.400 53.200 165.720 ;
        RECT 53.920 164.700 54.060 168.460 ;
        RECT 53.860 164.380 54.120 164.700 ;
        RECT 52.480 163.360 52.740 163.680 ;
        RECT 52.540 161.300 52.680 163.360 ;
        RECT 53.860 162.680 54.120 163.000 ;
        RECT 53.920 161.980 54.060 162.680 ;
        RECT 53.860 161.660 54.120 161.980 ;
        RECT 54.380 161.640 54.520 171.860 ;
        RECT 61.880 170.305 63.760 170.675 ;
        RECT 61.220 168.800 61.480 169.120 ;
        RECT 55.700 168.120 55.960 168.440 ;
        RECT 59.380 168.120 59.640 168.440 ;
        RECT 55.760 167.080 55.900 168.120 ;
        RECT 59.440 167.080 59.580 168.120 ;
        RECT 55.700 166.760 55.960 167.080 ;
        RECT 59.380 166.760 59.640 167.080 ;
        RECT 60.760 166.080 61.020 166.400 ;
        RECT 54.780 163.700 55.040 164.020 ;
        RECT 59.380 163.700 59.640 164.020 ;
        RECT 54.320 161.320 54.580 161.640 ;
        RECT 52.480 160.980 52.740 161.300 ;
        RECT 52.940 160.980 53.200 161.300 ;
        RECT 52.480 159.960 52.740 160.280 ;
        RECT 51.100 158.260 51.360 158.580 ;
        RECT 49.780 158.010 50.840 158.150 ;
        RECT 49.260 157.470 49.520 157.560 ;
        RECT 48.860 157.330 49.520 157.470 ;
        RECT 49.260 157.240 49.520 157.330 ;
        RECT 46.880 156.705 48.760 157.075 ;
        RECT 47.420 154.520 47.680 154.840 ;
        RECT 46.960 152.710 47.220 152.800 ;
        RECT 46.560 152.570 47.220 152.710 ;
        RECT 46.960 152.480 47.220 152.570 ;
        RECT 47.480 152.030 47.620 154.520 ;
        RECT 47.880 153.500 48.140 153.820 ;
        RECT 47.940 152.800 48.080 153.500 ;
        RECT 48.340 153.160 48.600 153.480 ;
        RECT 48.400 152.800 48.540 153.160 ;
        RECT 47.880 152.480 48.140 152.800 ;
        RECT 48.340 152.480 48.600 152.800 ;
        RECT 46.560 151.890 47.620 152.030 ;
        RECT 46.040 144.660 46.300 144.980 ;
        RECT 45.180 143.730 45.780 143.870 ;
        RECT 45.180 125.600 45.320 143.730 ;
        RECT 46.040 143.640 46.300 143.960 ;
        RECT 46.100 137.500 46.240 143.640 ;
        RECT 46.560 140.130 46.700 151.890 ;
        RECT 46.880 151.265 48.760 151.635 ;
        RECT 49.320 150.760 49.460 157.240 ;
        RECT 49.260 150.440 49.520 150.760 ;
        RECT 49.260 149.080 49.520 149.400 ;
        RECT 46.880 145.825 48.760 146.195 ;
        RECT 46.960 143.640 47.220 143.960 ;
        RECT 47.020 142.940 47.160 143.640 ;
        RECT 46.960 142.620 47.220 142.940 ;
        RECT 46.880 140.385 48.760 140.755 ;
        RECT 46.560 139.990 47.160 140.130 ;
        RECT 46.500 139.220 46.760 139.540 ;
        RECT 46.040 137.180 46.300 137.500 ;
        RECT 46.040 136.390 46.300 136.480 ;
        RECT 46.560 136.390 46.700 139.220 ;
        RECT 47.020 139.200 47.160 139.990 ;
        RECT 46.960 138.880 47.220 139.200 ;
        RECT 46.040 136.250 46.700 136.390 ;
        RECT 46.040 136.160 46.300 136.250 ;
        RECT 45.580 135.480 45.840 135.800 ;
        RECT 45.640 131.040 45.780 135.480 ;
        RECT 45.580 130.720 45.840 131.040 ;
        RECT 46.100 130.270 46.240 136.160 ;
        RECT 46.880 134.945 48.760 135.315 ;
        RECT 46.960 133.440 47.220 133.760 ;
        RECT 47.020 132.060 47.160 133.440 ;
        RECT 46.960 131.740 47.220 132.060 ;
        RECT 45.640 130.130 46.240 130.270 ;
        RECT 44.660 125.280 44.920 125.600 ;
        RECT 45.120 125.280 45.380 125.600 ;
        RECT 45.640 125.455 45.780 130.130 ;
        RECT 46.880 129.505 48.760 129.875 ;
        RECT 49.320 128.660 49.460 149.080 ;
        RECT 49.260 128.340 49.520 128.660 ;
        RECT 49.780 128.320 49.920 158.010 ;
        RECT 50.180 157.240 50.440 157.560 ;
        RECT 50.240 155.180 50.380 157.240 ;
        RECT 50.180 154.860 50.440 155.180 ;
        RECT 50.640 153.500 50.900 153.820 ;
        RECT 50.180 151.800 50.440 152.120 ;
        RECT 50.240 139.620 50.380 151.800 ;
        RECT 50.700 150.420 50.840 153.500 ;
        RECT 51.160 152.800 51.300 158.260 ;
        RECT 52.540 157.900 52.680 159.960 ;
        RECT 53.000 159.260 53.140 160.980 ;
        RECT 54.840 160.700 54.980 163.700 ;
        RECT 59.440 161.980 59.580 163.700 ;
        RECT 60.820 163.340 60.960 166.080 ;
        RECT 60.760 163.020 61.020 163.340 ;
        RECT 59.380 161.660 59.640 161.980 ;
        RECT 60.820 161.640 60.960 163.020 ;
        RECT 60.760 161.320 61.020 161.640 ;
        RECT 57.540 160.870 57.800 160.960 ;
        RECT 54.380 160.560 54.980 160.700 ;
        RECT 57.140 160.730 57.800 160.870 ;
        RECT 54.380 160.280 54.520 160.560 ;
        RECT 54.320 160.140 54.580 160.280 ;
        RECT 53.920 160.000 54.580 160.140 ;
        RECT 52.940 158.940 53.200 159.260 ;
        RECT 52.480 157.580 52.740 157.900 ;
        RECT 53.000 155.860 53.140 158.940 ;
        RECT 53.920 158.920 54.060 160.000 ;
        RECT 54.320 159.960 54.580 160.000 ;
        RECT 53.860 158.600 54.120 158.920 ;
        RECT 52.940 155.540 53.200 155.860 ;
        RECT 51.560 155.200 51.820 155.520 ;
        RECT 51.620 154.840 51.760 155.200 ;
        RECT 51.560 154.520 51.820 154.840 ;
        RECT 52.480 153.500 52.740 153.820 ;
        RECT 52.540 152.800 52.680 153.500 ;
        RECT 53.000 152.800 53.140 155.540 ;
        RECT 53.920 155.520 54.060 158.600 ;
        RECT 53.860 155.200 54.120 155.520 ;
        RECT 57.140 154.840 57.280 160.730 ;
        RECT 57.540 160.640 57.800 160.730 ;
        RECT 60.820 158.240 60.960 161.320 ;
        RECT 61.280 161.210 61.420 168.800 ;
        RECT 61.880 164.865 63.760 165.235 ;
        RECT 64.040 164.360 64.180 185.120 ;
        RECT 66.800 183.400 66.940 193.200 ;
        RECT 67.200 192.600 67.460 192.920 ;
        RECT 67.720 192.830 67.860 193.200 ;
        RECT 68.120 192.830 68.380 192.920 ;
        RECT 67.720 192.690 68.380 192.830 ;
        RECT 68.120 192.600 68.380 192.690 ;
        RECT 66.740 183.080 67.000 183.400 ;
        RECT 66.800 180.680 66.940 183.080 ;
        RECT 64.440 180.360 64.700 180.680 ;
        RECT 66.740 180.360 67.000 180.680 ;
        RECT 64.500 174.900 64.640 180.360 ;
        RECT 66.740 177.980 67.000 178.300 ;
        RECT 64.900 177.300 65.160 177.620 ;
        RECT 66.280 177.300 66.540 177.620 ;
        RECT 64.960 175.580 65.100 177.300 ;
        RECT 65.820 176.960 66.080 177.280 ;
        RECT 64.900 175.260 65.160 175.580 ;
        RECT 64.440 174.580 64.700 174.900 ;
        RECT 64.960 172.180 65.100 175.260 ;
        RECT 65.880 174.900 66.020 176.960 ;
        RECT 65.820 174.580 66.080 174.900 ;
        RECT 66.340 174.220 66.480 177.300 ;
        RECT 66.280 173.900 66.540 174.220 ;
        RECT 66.340 172.520 66.480 173.900 ;
        RECT 66.280 172.200 66.540 172.520 ;
        RECT 64.900 171.860 65.160 172.180 ;
        RECT 64.900 165.400 65.160 165.720 ;
        RECT 63.980 164.040 64.240 164.360 ;
        RECT 63.980 163.360 64.240 163.680 ;
        RECT 61.680 161.210 61.940 161.300 ;
        RECT 61.280 161.070 61.940 161.210 ;
        RECT 61.680 160.980 61.940 161.070 ;
        RECT 61.880 159.425 63.760 159.795 ;
        RECT 61.220 158.600 61.480 158.920 ;
        RECT 60.760 157.920 61.020 158.240 ;
        RECT 59.380 157.580 59.640 157.900 ;
        RECT 59.440 156.540 59.580 157.580 ;
        RECT 59.380 156.220 59.640 156.540 ;
        RECT 53.400 154.520 53.660 154.840 ;
        RECT 57.080 154.520 57.340 154.840 ;
        RECT 51.100 152.480 51.360 152.800 ;
        RECT 52.480 152.480 52.740 152.800 ;
        RECT 52.940 152.480 53.200 152.800 ;
        RECT 50.640 150.100 50.900 150.420 ;
        RECT 51.160 149.740 51.300 152.480 ;
        RECT 51.100 149.420 51.360 149.740 ;
        RECT 53.460 147.360 53.600 154.520 ;
        RECT 53.860 152.480 54.120 152.800 ;
        RECT 53.920 151.100 54.060 152.480 ;
        RECT 53.860 150.780 54.120 151.100 ;
        RECT 59.380 149.080 59.640 149.400 ;
        RECT 60.300 149.080 60.560 149.400 ;
        RECT 58.460 147.380 58.720 147.700 ;
        RECT 53.400 147.100 53.660 147.360 ;
        RECT 53.400 147.040 54.060 147.100 ;
        RECT 53.460 146.960 54.060 147.040 ;
        RECT 53.400 146.360 53.660 146.680 ;
        RECT 53.460 145.320 53.600 146.360 ;
        RECT 53.400 145.000 53.660 145.320 ;
        RECT 50.630 144.125 50.910 144.495 ;
        RECT 53.390 144.125 53.670 144.495 ;
        RECT 50.640 143.980 50.900 144.125 ;
        RECT 51.100 139.900 51.360 140.220 ;
        RECT 50.240 139.540 50.840 139.620 ;
        RECT 50.240 139.480 50.900 139.540 ;
        RECT 50.640 139.220 50.900 139.480 ;
        RECT 49.720 128.000 49.980 128.320 ;
        RECT 46.500 127.320 46.760 127.640 ;
        RECT 50.180 127.320 50.440 127.640 ;
        RECT 45.570 125.085 45.850 125.455 ;
        RECT 42.360 123.580 42.620 123.900 ;
        RECT 43.280 123.580 43.540 123.900 ;
        RECT 45.640 123.220 45.780 125.085 ;
        RECT 46.040 124.600 46.300 124.920 ;
        RECT 41.900 122.900 42.160 123.220 ;
        RECT 45.580 122.900 45.840 123.220 ;
        RECT 41.960 120.840 42.100 122.900 ;
        RECT 41.900 120.520 42.160 120.840 ;
        RECT 41.440 119.840 41.700 120.160 ;
        RECT 44.660 119.160 44.920 119.480 ;
        RECT 44.720 114.720 44.860 119.160 ;
        RECT 45.120 117.120 45.380 117.440 ;
        RECT 45.180 115.740 45.320 117.120 ;
        RECT 45.120 115.420 45.380 115.740 ;
        RECT 44.660 114.400 44.920 114.720 ;
        RECT 46.100 111.660 46.240 124.600 ;
        RECT 46.560 123.900 46.700 127.320 ;
        RECT 49.260 125.280 49.520 125.600 ;
        RECT 46.880 124.065 48.760 124.435 ;
        RECT 46.500 123.580 46.760 123.900 ;
        RECT 49.320 120.840 49.460 125.280 ;
        RECT 49.720 122.220 49.980 122.540 ;
        RECT 49.260 120.520 49.520 120.840 ;
        RECT 46.880 118.625 48.760 118.995 ;
        RECT 49.320 118.460 49.460 120.520 ;
        RECT 49.780 120.160 49.920 122.220 ;
        RECT 49.720 119.840 49.980 120.160 ;
        RECT 49.260 118.140 49.520 118.460 ;
        RECT 49.780 117.860 49.920 119.840 ;
        RECT 49.320 117.780 49.920 117.860 ;
        RECT 49.260 117.720 49.920 117.780 ;
        RECT 49.260 117.460 49.520 117.720 ;
        RECT 49.720 116.780 49.980 117.100 ;
        RECT 46.880 113.185 48.760 113.555 ;
        RECT 46.040 111.340 46.300 111.660 ;
        RECT 49.260 111.340 49.520 111.660 ;
        RECT 42.820 111.000 43.080 111.320 ;
        RECT 40.980 109.980 41.240 110.300 ;
        RECT 42.880 109.620 43.020 111.000 ;
        RECT 35.000 109.300 35.260 109.620 ;
        RECT 37.760 109.300 38.020 109.620 ;
        RECT 42.820 109.300 43.080 109.620 ;
        RECT 30.860 108.960 31.120 109.280 ;
        RECT 34.540 108.960 34.800 109.280 ;
        RECT 37.820 109.020 37.960 109.300 ;
        RECT 35.920 108.620 36.180 108.940 ;
        RECT 37.820 108.880 38.420 109.020 ;
        RECT 30.400 108.280 30.660 108.600 ;
        RECT 31.320 108.280 31.580 108.600 ;
        RECT 35.000 108.280 35.260 108.600 ;
        RECT 35.460 108.280 35.720 108.600 ;
        RECT 30.460 107.240 30.600 108.280 ;
        RECT 31.380 107.580 31.520 108.280 ;
        RECT 31.320 107.260 31.580 107.580 ;
        RECT 35.060 107.240 35.200 108.280 ;
        RECT 30.400 106.920 30.660 107.240 ;
        RECT 35.000 106.920 35.260 107.240 ;
        RECT 35.520 106.560 35.660 108.280 ;
        RECT 35.980 107.240 36.120 108.620 ;
        RECT 35.920 106.920 36.180 107.240 ;
        RECT 30.400 106.300 30.660 106.560 ;
        RECT 30.000 106.240 30.660 106.300 ;
        RECT 35.460 106.240 35.720 106.560 ;
        RECT 30.000 106.160 30.600 106.240 ;
        RECT 30.400 105.560 30.660 105.880 ;
        RECT 28.560 103.860 28.820 104.180 ;
        RECT 26.250 88.990 26.530 89.170 ;
        RECT 25.730 85.120 26.950 88.990 ;
        RECT 30.460 88.620 30.600 105.560 ;
        RECT 31.880 105.025 33.760 105.395 ;
        RECT 35.520 104.180 35.660 106.240 ;
        RECT 35.460 103.860 35.720 104.180 ;
        RECT 31.880 99.585 33.760 99.955 ;
        RECT 31.780 88.620 33.000 89.380 ;
        RECT 38.280 89.290 38.420 108.880 ;
        RECT 39.140 108.620 39.400 108.940 ;
        RECT 38.680 106.240 38.940 106.560 ;
        RECT 38.740 103.840 38.880 106.240 ;
        RECT 39.200 104.860 39.340 108.620 ;
        RECT 46.500 108.280 46.760 108.600 ;
        RECT 42.360 107.260 42.620 107.580 ;
        RECT 39.140 104.540 39.400 104.860 ;
        RECT 42.420 104.180 42.560 107.260 ;
        RECT 46.560 107.240 46.700 108.280 ;
        RECT 46.880 107.745 48.760 108.115 ;
        RECT 46.500 106.920 46.760 107.240 ;
        RECT 49.320 106.900 49.460 111.340 ;
        RECT 49.780 109.280 49.920 116.780 ;
        RECT 49.720 108.960 49.980 109.280 ;
        RECT 49.720 108.280 49.980 108.600 ;
        RECT 49.260 106.580 49.520 106.900 ;
        RECT 49.780 106.300 49.920 108.280 ;
        RECT 50.240 107.240 50.380 127.320 ;
        RECT 50.180 106.920 50.440 107.240 ;
        RECT 51.160 106.900 51.300 139.900 ;
        RECT 53.460 139.540 53.600 144.125 ;
        RECT 51.560 139.220 51.820 139.540 ;
        RECT 53.400 139.220 53.660 139.540 ;
        RECT 51.620 128.660 51.760 139.220 ;
        RECT 51.560 128.340 51.820 128.660 ;
        RECT 51.620 125.940 51.760 128.340 ;
        RECT 53.460 128.320 53.600 139.220 ;
        RECT 53.920 134.100 54.060 146.960 ;
        RECT 54.780 145.340 55.040 145.660 ;
        RECT 54.840 139.880 54.980 145.340 ;
        RECT 55.240 144.320 55.500 144.640 ;
        RECT 54.780 139.560 55.040 139.880 ;
        RECT 55.300 139.540 55.440 144.320 ;
        RECT 58.000 143.640 58.260 143.960 ;
        RECT 57.540 141.940 57.800 142.260 ;
        RECT 57.600 141.580 57.740 141.940 ;
        RECT 57.540 141.260 57.800 141.580 ;
        RECT 57.600 139.880 57.740 141.260 ;
        RECT 58.060 141.240 58.200 143.640 ;
        RECT 58.520 141.920 58.660 147.380 ;
        RECT 59.440 147.020 59.580 149.080 ;
        RECT 60.360 147.700 60.500 149.080 ;
        RECT 60.820 147.700 60.960 157.920 ;
        RECT 61.280 156.200 61.420 158.600 ;
        RECT 61.220 155.880 61.480 156.200 ;
        RECT 61.880 153.985 63.760 154.355 ;
        RECT 64.040 152.800 64.180 163.360 ;
        RECT 64.440 152.820 64.700 153.140 ;
        RECT 63.980 152.655 64.240 152.800 ;
        RECT 63.970 152.285 64.250 152.655 ;
        RECT 64.500 152.460 64.640 152.820 ;
        RECT 64.440 152.140 64.700 152.460 ;
        RECT 63.980 151.800 64.240 152.120 ;
        RECT 61.680 150.100 61.940 150.420 ;
        RECT 61.740 149.400 61.880 150.100 ;
        RECT 61.680 149.080 61.940 149.400 ;
        RECT 61.880 148.545 63.760 148.915 ;
        RECT 60.300 147.380 60.560 147.700 ;
        RECT 60.760 147.380 61.020 147.700 ;
        RECT 59.380 146.700 59.640 147.020 ;
        RECT 60.360 146.680 60.500 147.380 ;
        RECT 64.040 147.020 64.180 151.800 ;
        RECT 64.500 149.740 64.640 152.140 ;
        RECT 64.960 150.420 65.100 165.400 ;
        RECT 66.800 164.100 66.940 177.980 ;
        RECT 67.260 169.120 67.400 192.600 ;
        RECT 69.100 191.220 69.240 193.280 ;
        RECT 70.020 191.900 70.160 193.620 ;
        RECT 70.480 191.900 70.620 196.340 ;
        RECT 70.940 194.620 71.080 199.400 ;
        RECT 71.400 195.640 71.540 199.400 ;
        RECT 75.940 199.060 76.200 199.380 ;
        RECT 71.800 198.040 72.060 198.360 ;
        RECT 71.340 195.320 71.600 195.640 ;
        RECT 71.400 194.620 71.540 195.320 ;
        RECT 70.880 194.300 71.140 194.620 ;
        RECT 71.340 194.300 71.600 194.620 ;
        RECT 70.880 192.600 71.140 192.920 ;
        RECT 70.940 191.900 71.080 192.600 ;
        RECT 69.960 191.580 70.220 191.900 ;
        RECT 70.420 191.580 70.680 191.900 ;
        RECT 70.880 191.580 71.140 191.900 ;
        RECT 69.040 190.900 69.300 191.220 ;
        RECT 67.660 184.440 67.920 184.760 ;
        RECT 67.720 182.630 67.860 184.440 ;
        RECT 69.100 183.740 69.240 190.900 ;
        RECT 70.420 190.790 70.680 190.880 ;
        RECT 71.860 190.790 72.000 198.040 ;
        RECT 76.000 196.320 76.140 199.060 ;
        RECT 77.380 197.340 77.520 199.400 ;
        RECT 111.820 199.060 112.080 199.380 ;
        RECT 82.380 198.720 82.640 199.040 ;
        RECT 93.880 198.720 94.140 199.040 ;
        RECT 82.440 197.340 82.580 198.720 ;
        RECT 91.880 197.505 93.760 197.875 ;
        RECT 77.320 197.020 77.580 197.340 ;
        RECT 82.380 197.020 82.640 197.340 ;
        RECT 76.400 196.340 76.660 196.660 ;
        RECT 91.580 196.340 91.840 196.660 ;
        RECT 75.940 196.000 76.200 196.320 ;
        RECT 73.640 195.660 73.900 195.980 ;
        RECT 73.700 194.620 73.840 195.660 ;
        RECT 75.020 195.320 75.280 195.640 ;
        RECT 73.640 194.300 73.900 194.620 ;
        RECT 72.260 193.280 72.520 193.600 ;
        RECT 72.320 191.220 72.460 193.280 ;
        RECT 73.700 192.920 73.840 194.300 ;
        RECT 75.080 194.280 75.220 195.320 ;
        RECT 75.020 193.960 75.280 194.280 ;
        RECT 73.640 192.600 73.900 192.920 ;
        RECT 74.560 192.600 74.820 192.920 ;
        RECT 75.480 192.600 75.740 192.920 ;
        RECT 76.000 192.830 76.140 196.000 ;
        RECT 76.460 194.280 76.600 196.340 ;
        RECT 86.520 195.660 86.780 195.980 ;
        RECT 86.060 195.320 86.320 195.640 ;
        RECT 76.880 194.785 78.760 195.155 ;
        RECT 76.400 193.960 76.660 194.280 ;
        RECT 76.860 193.620 77.120 193.940 ;
        RECT 77.780 193.620 78.040 193.940 ;
        RECT 76.400 192.830 76.660 192.920 ;
        RECT 76.000 192.690 76.660 192.830 ;
        RECT 76.400 192.600 76.660 192.690 ;
        RECT 72.260 190.900 72.520 191.220 ;
        RECT 70.420 190.650 72.000 190.790 ;
        RECT 70.420 190.560 70.680 190.650 ;
        RECT 69.040 183.420 69.300 183.740 ;
        RECT 68.120 182.630 68.380 182.720 ;
        RECT 67.720 182.490 68.380 182.630 ;
        RECT 68.120 182.400 68.380 182.490 ;
        RECT 68.580 182.400 68.840 182.720 ;
        RECT 68.180 180.340 68.320 182.400 ;
        RECT 68.640 182.040 68.780 182.400 ;
        RECT 68.580 181.720 68.840 182.040 ;
        RECT 68.120 180.020 68.380 180.340 ;
        RECT 69.100 177.280 69.240 183.420 ;
        RECT 70.420 182.740 70.680 183.060 ;
        RECT 69.500 181.720 69.760 182.040 ;
        RECT 69.560 180.000 69.700 181.720 ;
        RECT 69.500 179.680 69.760 180.000 ;
        RECT 69.500 179.000 69.760 179.320 ;
        RECT 69.960 179.000 70.220 179.320 ;
        RECT 69.040 176.960 69.300 177.280 ;
        RECT 68.580 175.260 68.840 175.580 ;
        RECT 67.200 168.800 67.460 169.120 ;
        RECT 68.120 168.460 68.380 168.780 ;
        RECT 66.340 164.020 66.940 164.100 ;
        RECT 66.280 163.960 66.940 164.020 ;
        RECT 66.280 163.700 66.540 163.960 ;
        RECT 66.740 163.360 67.000 163.680 ;
        RECT 66.800 161.300 66.940 163.360 ;
        RECT 66.740 160.980 67.000 161.300 ;
        RECT 66.740 157.240 67.000 157.560 ;
        RECT 66.800 156.200 66.940 157.240 ;
        RECT 66.740 155.880 67.000 156.200 ;
        RECT 66.800 153.820 66.940 155.880 ;
        RECT 67.660 154.520 67.920 154.840 ;
        RECT 66.740 153.500 67.000 153.820 ;
        RECT 66.740 152.480 67.000 152.800 ;
        RECT 65.360 151.800 65.620 152.120 ;
        RECT 64.900 150.100 65.160 150.420 ;
        RECT 64.440 149.420 64.700 149.740 ;
        RECT 63.980 146.700 64.240 147.020 ;
        RECT 60.300 146.360 60.560 146.680 ;
        RECT 61.220 144.660 61.480 144.980 ;
        RECT 59.840 144.320 60.100 144.640 ;
        RECT 58.920 142.620 59.180 142.940 ;
        RECT 58.460 141.600 58.720 141.920 ;
        RECT 58.980 141.580 59.120 142.620 ;
        RECT 58.920 141.260 59.180 141.580 ;
        RECT 58.000 140.920 58.260 141.240 ;
        RECT 58.060 140.220 58.200 140.920 ;
        RECT 58.000 139.900 58.260 140.220 ;
        RECT 57.540 139.560 57.800 139.880 ;
        RECT 55.240 139.220 55.500 139.540 ;
        RECT 55.300 138.520 55.440 139.220 ;
        RECT 55.240 138.430 55.500 138.520 ;
        RECT 54.840 138.290 55.500 138.430 ;
        RECT 53.860 133.780 54.120 134.100 ;
        RECT 54.840 128.660 54.980 138.290 ;
        RECT 55.240 138.200 55.500 138.290 ;
        RECT 55.700 133.780 55.960 134.100 ;
        RECT 55.760 131.040 55.900 133.780 ;
        RECT 57.600 131.380 57.740 139.560 ;
        RECT 58.920 138.880 59.180 139.200 ;
        RECT 58.000 135.820 58.260 136.140 ;
        RECT 58.060 134.780 58.200 135.820 ;
        RECT 58.980 135.800 59.120 138.880 ;
        RECT 59.900 136.820 60.040 144.320 ;
        RECT 60.760 143.640 61.020 143.960 ;
        RECT 60.820 142.260 60.960 143.640 ;
        RECT 61.280 142.940 61.420 144.660 ;
        RECT 64.500 143.960 64.640 149.420 ;
        RECT 64.900 149.255 65.160 149.400 ;
        RECT 64.890 148.885 65.170 149.255 ;
        RECT 65.420 148.380 65.560 151.800 ;
        RECT 66.800 150.760 66.940 152.480 ;
        RECT 66.740 150.440 67.000 150.760 ;
        RECT 65.820 150.100 66.080 150.420 ;
        RECT 65.360 148.060 65.620 148.380 ;
        RECT 65.880 145.570 66.020 150.100 ;
        RECT 66.800 149.400 66.940 150.440 ;
        RECT 66.740 149.080 67.000 149.400 ;
        RECT 65.420 145.430 66.020 145.570 ;
        RECT 65.420 144.300 65.560 145.430 ;
        RECT 65.820 144.660 66.080 144.980 ;
        RECT 66.280 144.660 66.540 144.980 ;
        RECT 65.360 143.980 65.620 144.300 ;
        RECT 64.440 143.640 64.700 143.960 ;
        RECT 61.880 143.105 63.760 143.475 ;
        RECT 61.220 142.620 61.480 142.940 ;
        RECT 60.760 141.940 61.020 142.260 ;
        RECT 64.500 141.920 64.640 143.640 ;
        RECT 65.420 141.920 65.560 143.980 ;
        RECT 65.880 143.960 66.020 144.660 ;
        RECT 65.820 143.640 66.080 143.960 ;
        RECT 64.440 141.600 64.700 141.920 ;
        RECT 64.900 141.600 65.160 141.920 ;
        RECT 65.360 141.600 65.620 141.920 ;
        RECT 64.960 140.220 65.100 141.600 ;
        RECT 64.900 139.900 65.160 140.220 ;
        RECT 61.220 138.200 61.480 138.520 ;
        RECT 59.840 136.730 60.100 136.820 ;
        RECT 59.840 136.590 60.500 136.730 ;
        RECT 59.840 136.500 60.100 136.590 ;
        RECT 58.920 135.480 59.180 135.800 ;
        RECT 58.000 134.460 58.260 134.780 ;
        RECT 57.540 131.060 57.800 131.380 ;
        RECT 55.700 130.720 55.960 131.040 ;
        RECT 54.780 128.340 55.040 128.660 ;
        RECT 53.400 128.000 53.660 128.320 ;
        RECT 52.020 127.660 52.280 127.980 ;
        RECT 52.080 126.280 52.220 127.660 ;
        RECT 52.020 125.960 52.280 126.280 ;
        RECT 51.560 125.620 51.820 125.940 ;
        RECT 52.080 125.600 52.220 125.960 ;
        RECT 54.840 125.600 54.980 128.340 ;
        RECT 52.020 125.280 52.280 125.600 ;
        RECT 52.480 125.280 52.740 125.600 ;
        RECT 54.780 125.280 55.040 125.600 ;
        RECT 52.080 120.160 52.220 125.280 ;
        RECT 52.540 120.160 52.680 125.280 ;
        RECT 54.840 124.920 54.980 125.280 ;
        RECT 54.780 124.600 55.040 124.920 ;
        RECT 54.840 120.500 54.980 124.600 ;
        RECT 55.760 123.560 55.900 130.720 ;
        RECT 56.160 130.040 56.420 130.360 ;
        RECT 56.620 130.040 56.880 130.360 ;
        RECT 56.220 129.000 56.360 130.040 ;
        RECT 56.680 129.340 56.820 130.040 ;
        RECT 56.620 129.020 56.880 129.340 ;
        RECT 56.160 128.680 56.420 129.000 ;
        RECT 56.680 125.600 56.820 129.020 ;
        RECT 57.600 126.020 57.740 131.060 ;
        RECT 58.980 131.040 59.120 135.480 ;
        RECT 60.360 133.760 60.500 136.590 ;
        RECT 61.280 136.480 61.420 138.200 ;
        RECT 61.880 137.665 63.760 138.035 ;
        RECT 61.220 136.160 61.480 136.480 ;
        RECT 66.340 134.100 66.480 144.660 ;
        RECT 66.800 144.640 66.940 149.080 ;
        RECT 66.740 144.320 67.000 144.640 ;
        RECT 66.800 142.260 66.940 144.320 ;
        RECT 67.720 142.600 67.860 154.520 ;
        RECT 67.660 142.280 67.920 142.600 ;
        RECT 66.740 141.940 67.000 142.260 ;
        RECT 67.660 141.260 67.920 141.580 ;
        RECT 66.280 133.780 66.540 134.100 ;
        RECT 60.300 133.440 60.560 133.760 ;
        RECT 58.920 130.720 59.180 131.040 ;
        RECT 60.360 128.660 60.500 133.440 ;
        RECT 61.880 132.225 63.760 132.595 ;
        RECT 64.440 130.040 64.700 130.360 ;
        RECT 64.500 128.660 64.640 130.040 ;
        RECT 60.300 128.340 60.560 128.660 ;
        RECT 63.980 128.340 64.240 128.660 ;
        RECT 64.440 128.340 64.700 128.660 ;
        RECT 61.880 126.785 63.760 127.155 ;
        RECT 57.600 125.940 58.200 126.020 ;
        RECT 64.040 125.940 64.180 128.340 ;
        RECT 57.540 125.880 58.200 125.940 ;
        RECT 57.540 125.620 57.800 125.880 ;
        RECT 56.620 125.280 56.880 125.600 ;
        RECT 57.540 124.940 57.800 125.260 ;
        RECT 55.700 123.240 55.960 123.560 ;
        RECT 54.780 120.180 55.040 120.500 ;
        RECT 55.760 120.160 55.900 123.240 ;
        RECT 56.160 122.900 56.420 123.220 ;
        RECT 56.220 122.735 56.360 122.900 ;
        RECT 56.150 122.365 56.430 122.735 ;
        RECT 52.020 119.840 52.280 120.160 ;
        RECT 52.480 119.840 52.740 120.160 ;
        RECT 55.700 119.840 55.960 120.160 ;
        RECT 56.220 120.015 56.360 122.365 ;
        RECT 57.600 120.160 57.740 124.940 ;
        RECT 58.060 121.180 58.200 125.880 ;
        RECT 63.980 125.620 64.240 125.940 ;
        RECT 65.820 125.620 66.080 125.940 ;
        RECT 61.680 124.940 61.940 125.260 ;
        RECT 61.740 123.900 61.880 124.940 ;
        RECT 62.140 124.600 62.400 124.920 ;
        RECT 61.680 123.580 61.940 123.900 ;
        RECT 62.200 123.220 62.340 124.600 ;
        RECT 62.140 122.900 62.400 123.220 ;
        RECT 64.040 122.540 64.180 125.620 ;
        RECT 65.880 123.900 66.020 125.620 ;
        RECT 65.820 123.580 66.080 123.900 ;
        RECT 63.980 122.220 64.240 122.540 ;
        RECT 61.880 121.345 63.760 121.715 ;
        RECT 58.000 120.860 58.260 121.180 ;
        RECT 58.460 120.520 58.720 120.840 ;
        RECT 63.520 120.520 63.780 120.840 ;
        RECT 58.000 120.180 58.260 120.500 ;
        RECT 56.150 119.645 56.430 120.015 ;
        RECT 57.540 119.840 57.800 120.160 ;
        RECT 57.080 119.500 57.340 119.820 ;
        RECT 54.780 119.160 55.040 119.480 ;
        RECT 54.840 118.120 54.980 119.160 ;
        RECT 54.780 117.800 55.040 118.120 ;
        RECT 57.140 116.760 57.280 119.500 ;
        RECT 57.080 116.440 57.340 116.760 ;
        RECT 57.140 115.060 57.280 116.440 ;
        RECT 57.080 114.740 57.340 115.060 ;
        RECT 57.140 113.020 57.280 114.740 ;
        RECT 58.060 114.720 58.200 120.180 ;
        RECT 58.520 115.400 58.660 120.520 ;
        RECT 62.140 119.160 62.400 119.480 ;
        RECT 62.200 117.780 62.340 119.160 ;
        RECT 63.580 117.780 63.720 120.520 ;
        RECT 64.040 120.500 64.180 122.220 ;
        RECT 63.980 120.180 64.240 120.500 ;
        RECT 62.140 117.460 62.400 117.780 ;
        RECT 63.520 117.460 63.780 117.780 ;
        RECT 64.040 117.440 64.180 120.180 ;
        RECT 66.340 118.460 66.480 133.780 ;
        RECT 67.200 128.340 67.460 128.660 ;
        RECT 66.280 118.140 66.540 118.460 ;
        RECT 63.980 117.120 64.240 117.440 ;
        RECT 61.880 115.905 63.760 116.275 ;
        RECT 58.460 115.080 58.720 115.400 ;
        RECT 58.000 114.400 58.260 114.720 ;
        RECT 59.380 113.720 59.640 114.040 ;
        RECT 57.080 112.700 57.340 113.020 ;
        RECT 56.620 112.360 56.880 112.680 ;
        RECT 56.680 110.300 56.820 112.360 ;
        RECT 56.620 109.980 56.880 110.300 ;
        RECT 59.440 109.280 59.580 113.720 ;
        RECT 64.040 112.340 64.180 117.120 ;
        RECT 66.340 115.740 66.480 118.140 ;
        RECT 66.280 115.420 66.540 115.740 ;
        RECT 67.260 112.340 67.400 128.340 ;
        RECT 63.980 112.020 64.240 112.340 ;
        RECT 67.200 112.020 67.460 112.340 ;
        RECT 60.300 111.680 60.560 112.000 ;
        RECT 60.360 110.300 60.500 111.680 ;
        RECT 61.880 110.465 63.760 110.835 ;
        RECT 60.300 109.980 60.560 110.300 ;
        RECT 59.380 108.960 59.640 109.280 ;
        RECT 52.940 107.260 53.200 107.580 ;
        RECT 51.100 106.580 51.360 106.900 ;
        RECT 49.320 106.160 49.920 106.300 ;
        RECT 50.180 106.240 50.440 106.560 ;
        RECT 44.200 105.560 44.460 105.880 ;
        RECT 42.360 103.860 42.620 104.180 ;
        RECT 38.680 103.520 38.940 103.840 ;
        RECT 44.260 89.530 44.400 105.560 ;
        RECT 46.040 103.180 46.300 103.500 ;
        RECT 46.100 102.140 46.240 103.180 ;
        RECT 49.320 103.160 49.460 106.160 ;
        RECT 50.240 104.860 50.380 106.240 ;
        RECT 52.480 105.560 52.740 105.880 ;
        RECT 50.180 104.540 50.440 104.860 ;
        RECT 52.540 104.180 52.680 105.560 ;
        RECT 53.000 104.180 53.140 107.260 ;
        RECT 55.700 106.580 55.960 106.900 ;
        RECT 52.480 103.860 52.740 104.180 ;
        RECT 52.940 103.860 53.200 104.180 ;
        RECT 49.260 102.840 49.520 103.160 ;
        RECT 49.720 102.840 49.980 103.160 ;
        RECT 46.880 102.305 48.760 102.675 ;
        RECT 46.040 101.820 46.300 102.140 ;
        RECT 49.320 101.460 49.460 102.840 ;
        RECT 49.260 101.140 49.520 101.460 ;
        RECT 37.750 88.780 38.970 89.290 ;
        RECT 30.460 88.480 33.000 88.620 ;
        RECT 31.780 85.510 33.000 88.480 ;
        RECT 37.680 88.620 38.970 88.780 ;
        RECT 43.810 88.630 45.030 89.530 ;
        RECT 49.780 89.040 49.920 102.840 ;
        RECT 55.760 101.460 55.900 106.580 ;
        RECT 57.540 105.560 57.800 105.880 ;
        RECT 61.220 105.560 61.480 105.880 ;
        RECT 57.600 103.500 57.740 105.560 ;
        RECT 61.280 103.500 61.420 105.560 ;
        RECT 61.880 105.025 63.760 105.395 ;
        RECT 64.040 104.860 64.180 112.020 ;
        RECT 67.720 109.280 67.860 141.260 ;
        RECT 68.180 134.440 68.320 168.460 ;
        RECT 68.640 163.340 68.780 175.260 ;
        RECT 69.100 174.900 69.240 176.960 ;
        RECT 69.040 174.580 69.300 174.900 ;
        RECT 69.040 173.900 69.300 174.220 ;
        RECT 69.100 164.700 69.240 173.900 ;
        RECT 69.560 164.700 69.700 179.000 ;
        RECT 70.020 178.300 70.160 179.000 ;
        RECT 69.960 177.980 70.220 178.300 ;
        RECT 69.960 177.300 70.220 177.620 ;
        RECT 70.020 173.880 70.160 177.300 ;
        RECT 69.960 173.560 70.220 173.880 ;
        RECT 70.020 172.520 70.160 173.560 ;
        RECT 69.960 172.200 70.220 172.520 ;
        RECT 69.960 171.520 70.220 171.840 ;
        RECT 70.020 166.060 70.160 171.520 ;
        RECT 69.960 165.740 70.220 166.060 ;
        RECT 69.040 164.380 69.300 164.700 ;
        RECT 69.500 164.380 69.760 164.700 ;
        RECT 68.580 163.020 68.840 163.340 ;
        RECT 68.640 158.580 68.780 163.020 ;
        RECT 69.100 161.980 69.240 164.380 ;
        RECT 69.040 161.660 69.300 161.980 ;
        RECT 68.580 158.260 68.840 158.580 ;
        RECT 69.560 158.240 69.700 164.380 ;
        RECT 69.960 163.535 70.220 163.680 ;
        RECT 69.950 163.165 70.230 163.535 ;
        RECT 69.500 157.920 69.760 158.240 ;
        RECT 70.480 155.860 70.620 182.740 ;
        RECT 70.880 180.360 71.140 180.680 ;
        RECT 70.940 175.580 71.080 180.360 ;
        RECT 71.400 180.340 71.540 190.650 ;
        RECT 72.320 190.200 72.460 190.900 ;
        RECT 72.260 189.880 72.520 190.200 ;
        RECT 72.260 187.840 72.520 188.160 ;
        RECT 72.320 183.400 72.460 187.840 ;
        RECT 72.260 183.080 72.520 183.400 ;
        RECT 73.700 182.720 73.840 192.600 ;
        RECT 74.620 188.500 74.760 192.600 ;
        RECT 75.540 191.900 75.680 192.600 ;
        RECT 75.480 191.580 75.740 191.900 ;
        RECT 75.020 190.900 75.280 191.220 ;
        RECT 74.560 188.180 74.820 188.500 ;
        RECT 74.100 187.160 74.360 187.480 ;
        RECT 74.160 185.780 74.300 187.160 ;
        RECT 74.100 185.460 74.360 185.780 ;
        RECT 73.640 182.400 73.900 182.720 ;
        RECT 71.340 180.020 71.600 180.340 ;
        RECT 72.260 179.340 72.520 179.660 ;
        RECT 70.880 175.260 71.140 175.580 ;
        RECT 71.340 175.260 71.600 175.580 ;
        RECT 70.940 174.900 71.080 175.260 ;
        RECT 70.880 174.580 71.140 174.900 ;
        RECT 71.400 172.520 71.540 175.260 ;
        RECT 72.320 174.900 72.460 179.340 ;
        RECT 72.720 176.960 72.980 177.280 ;
        RECT 72.780 174.900 72.920 176.960 ;
        RECT 73.700 175.240 73.840 182.400 ;
        RECT 75.080 180.000 75.220 190.900 ;
        RECT 76.460 188.160 76.600 192.600 ;
        RECT 76.920 191.220 77.060 193.620 ;
        RECT 76.860 190.900 77.120 191.220 ;
        RECT 77.840 190.880 77.980 193.620 ;
        RECT 86.120 193.600 86.260 195.320 ;
        RECT 85.140 193.280 85.400 193.600 ;
        RECT 86.060 193.280 86.320 193.600 ;
        RECT 85.200 191.900 85.340 193.280 ;
        RECT 85.140 191.580 85.400 191.900 ;
        RECT 77.780 190.560 78.040 190.880 ;
        RECT 76.880 189.345 78.760 189.715 ;
        RECT 76.400 187.840 76.660 188.160 ;
        RECT 76.460 185.440 76.600 187.840 ;
        RECT 85.200 185.780 85.340 191.580 ;
        RECT 86.120 191.220 86.260 193.280 ;
        RECT 86.060 190.900 86.320 191.220 ;
        RECT 85.140 185.460 85.400 185.780 ;
        RECT 75.480 185.120 75.740 185.440 ;
        RECT 76.400 185.120 76.660 185.440 ;
        RECT 75.540 182.720 75.680 185.120 ;
        RECT 75.480 182.400 75.740 182.720 ;
        RECT 76.460 181.100 76.600 185.120 ;
        RECT 84.680 184.780 84.940 185.100 ;
        RECT 76.880 183.905 78.760 184.275 ;
        RECT 77.320 183.080 77.580 183.400 ;
        RECT 76.460 180.960 77.060 181.100 ;
        RECT 77.380 181.020 77.520 183.080 ;
        RECT 84.740 183.060 84.880 184.780 ;
        RECT 84.680 182.740 84.940 183.060 ;
        RECT 76.400 180.020 76.660 180.340 ;
        RECT 75.020 179.680 75.280 180.000 ;
        RECT 76.460 178.300 76.600 180.020 ;
        RECT 76.920 179.660 77.060 180.960 ;
        RECT 77.320 180.700 77.580 181.020 ;
        RECT 84.740 180.680 84.880 182.740 ;
        RECT 85.200 182.720 85.340 185.460 ;
        RECT 85.140 182.400 85.400 182.720 ;
        RECT 85.200 181.020 85.340 182.400 ;
        RECT 85.140 180.700 85.400 181.020 ;
        RECT 81.460 180.360 81.720 180.680 ;
        RECT 84.680 180.360 84.940 180.680 ;
        RECT 76.860 179.340 77.120 179.660 ;
        RECT 76.880 178.465 78.760 178.835 ;
        RECT 76.400 177.980 76.660 178.300 ;
        RECT 77.320 177.980 77.580 178.300 ;
        RECT 77.380 177.620 77.520 177.980 ;
        RECT 81.520 177.960 81.660 180.360 ;
        RECT 85.200 180.340 85.340 180.700 ;
        RECT 85.140 180.020 85.400 180.340 ;
        RECT 84.680 179.680 84.940 180.000 ;
        RECT 81.460 177.640 81.720 177.960 ;
        RECT 84.740 177.620 84.880 179.680 ;
        RECT 76.400 177.300 76.660 177.620 ;
        RECT 77.320 177.300 77.580 177.620 ;
        RECT 78.700 177.300 78.960 177.620 ;
        RECT 79.160 177.300 79.420 177.620 ;
        RECT 84.680 177.300 84.940 177.620 ;
        RECT 73.640 174.920 73.900 175.240 ;
        RECT 72.260 174.580 72.520 174.900 ;
        RECT 72.720 174.580 72.980 174.900 ;
        RECT 71.340 172.200 71.600 172.520 ;
        RECT 70.880 171.860 71.140 172.180 ;
        RECT 70.420 155.540 70.680 155.860 ;
        RECT 68.580 154.860 68.840 155.180 ;
        RECT 68.640 153.335 68.780 154.860 ;
        RECT 69.500 154.520 69.760 154.840 ;
        RECT 68.570 152.965 68.850 153.335 ;
        RECT 68.640 152.800 68.780 152.965 ;
        RECT 68.580 152.480 68.840 152.800 ;
        RECT 69.040 151.800 69.300 152.120 ;
        RECT 68.580 149.420 68.840 149.740 ;
        RECT 68.640 145.660 68.780 149.420 ;
        RECT 69.100 147.020 69.240 151.800 ;
        RECT 69.560 149.740 69.700 154.520 ;
        RECT 70.480 152.800 70.620 155.540 ;
        RECT 70.940 153.820 71.080 171.860 ;
        RECT 71.400 169.460 71.540 172.200 ;
        RECT 72.320 171.500 72.460 174.580 ;
        RECT 72.780 172.180 72.920 174.580 ;
        RECT 73.700 172.860 73.840 174.920 ;
        RECT 76.460 174.560 76.600 177.300 ;
        RECT 78.760 176.940 78.900 177.300 ;
        RECT 78.700 176.620 78.960 176.940 ;
        RECT 78.760 174.560 78.900 176.620 ;
        RECT 79.220 175.095 79.360 177.300 ;
        RECT 81.000 176.960 81.260 177.280 ;
        RECT 80.080 176.280 80.340 176.600 ;
        RECT 80.540 176.455 80.800 176.600 ;
        RECT 80.140 175.580 80.280 176.280 ;
        RECT 80.530 176.085 80.810 176.455 ;
        RECT 80.080 175.260 80.340 175.580 ;
        RECT 79.150 174.725 79.430 175.095 ;
        RECT 81.060 174.900 81.200 176.960 ;
        RECT 82.840 176.280 83.100 176.600 ;
        RECT 79.220 174.560 79.360 174.725 ;
        RECT 81.000 174.580 81.260 174.900 ;
        RECT 76.400 174.240 76.660 174.560 ;
        RECT 78.700 174.240 78.960 174.560 ;
        RECT 79.160 174.240 79.420 174.560 ;
        RECT 73.640 172.540 73.900 172.860 ;
        RECT 72.720 171.860 72.980 172.180 ;
        RECT 71.800 171.180 72.060 171.500 ;
        RECT 72.260 171.180 72.520 171.500 ;
        RECT 71.860 170.140 72.000 171.180 ;
        RECT 71.800 169.820 72.060 170.140 ;
        RECT 71.340 169.140 71.600 169.460 ;
        RECT 71.860 166.740 72.000 169.820 ;
        RECT 72.780 169.120 72.920 171.860 ;
        RECT 73.700 169.460 73.840 172.540 ;
        RECT 76.460 171.500 76.600 174.240 ;
        RECT 76.880 173.025 78.760 173.395 ;
        RECT 79.220 172.180 79.360 174.240 ;
        RECT 79.620 173.900 79.880 174.220 ;
        RECT 80.540 173.900 80.800 174.220 ;
        RECT 79.680 172.520 79.820 173.900 ;
        RECT 79.620 172.200 79.880 172.520 ;
        RECT 79.160 171.860 79.420 172.180 ;
        RECT 76.400 171.180 76.660 171.500 ;
        RECT 73.640 169.140 73.900 169.460 ;
        RECT 72.720 168.800 72.980 169.120 ;
        RECT 76.460 167.420 76.600 171.180 ;
        RECT 79.680 171.160 79.820 172.200 ;
        RECT 79.620 170.840 79.880 171.160 ;
        RECT 80.080 170.840 80.340 171.160 ;
        RECT 76.880 167.585 78.760 167.955 ;
        RECT 76.400 167.100 76.660 167.420 ;
        RECT 71.800 166.420 72.060 166.740 ;
        RECT 71.340 165.740 71.600 166.060 ;
        RECT 71.400 164.020 71.540 165.740 ;
        RECT 71.340 163.700 71.600 164.020 ;
        RECT 71.860 163.930 72.000 166.420 ;
        RECT 74.100 164.040 74.360 164.360 ;
        RECT 72.260 163.930 72.520 164.020 ;
        RECT 71.860 163.790 72.520 163.930 ;
        RECT 71.860 161.300 72.000 163.790 ;
        RECT 72.260 163.700 72.520 163.790 ;
        RECT 73.180 163.590 73.440 163.680 ;
        RECT 73.180 163.450 73.840 163.590 ;
        RECT 73.180 163.360 73.440 163.450 ;
        RECT 72.260 162.680 72.520 163.000 ;
        RECT 72.320 161.640 72.460 162.680 ;
        RECT 72.260 161.320 72.520 161.640 ;
        RECT 71.800 160.980 72.060 161.300 ;
        RECT 71.860 155.860 72.000 160.980 ;
        RECT 71.800 155.540 72.060 155.860 ;
        RECT 72.260 155.200 72.520 155.520 ;
        RECT 72.320 154.840 72.460 155.200 ;
        RECT 72.260 154.520 72.520 154.840 ;
        RECT 70.880 153.500 71.140 153.820 ;
        RECT 70.420 152.480 70.680 152.800 ;
        RECT 69.960 152.140 70.220 152.460 ;
        RECT 69.500 149.420 69.760 149.740 ;
        RECT 69.040 146.700 69.300 147.020 ;
        RECT 68.580 145.340 68.840 145.660 ;
        RECT 68.640 144.495 68.780 145.340 ;
        RECT 69.100 144.640 69.240 146.700 ;
        RECT 70.020 144.640 70.160 152.140 ;
        RECT 70.480 150.760 70.620 152.480 ;
        RECT 72.320 151.100 72.460 154.520 ;
        RECT 73.180 153.500 73.440 153.820 ;
        RECT 72.710 152.285 72.990 152.655 ;
        RECT 72.260 150.780 72.520 151.100 ;
        RECT 70.420 150.440 70.680 150.760 ;
        RECT 72.260 150.100 72.520 150.420 ;
        RECT 71.800 149.080 72.060 149.400 ;
        RECT 70.880 147.380 71.140 147.700 ;
        RECT 70.420 145.000 70.680 145.320 ;
        RECT 68.570 144.125 68.850 144.495 ;
        RECT 69.040 144.320 69.300 144.640 ;
        RECT 69.960 144.320 70.220 144.640 ;
        RECT 68.580 142.280 68.840 142.600 ;
        RECT 68.640 139.880 68.780 142.280 ;
        RECT 69.100 141.240 69.240 144.320 ;
        RECT 70.020 142.940 70.160 144.320 ;
        RECT 69.960 142.620 70.220 142.940 ;
        RECT 69.040 140.920 69.300 141.240 ;
        RECT 68.580 139.560 68.840 139.880 ;
        RECT 68.120 134.120 68.380 134.440 ;
        RECT 69.100 133.760 69.240 140.920 ;
        RECT 70.480 140.220 70.620 145.000 ;
        RECT 69.500 139.900 69.760 140.220 ;
        RECT 70.420 139.900 70.680 140.220 ;
        RECT 69.560 134.780 69.700 139.900 ;
        RECT 69.500 134.460 69.760 134.780 ;
        RECT 69.040 133.440 69.300 133.760 ;
        RECT 69.560 132.060 69.700 134.460 ;
        RECT 70.420 134.120 70.680 134.440 ;
        RECT 69.960 132.760 70.220 133.080 ;
        RECT 70.020 132.060 70.160 132.760 ;
        RECT 69.500 131.740 69.760 132.060 ;
        RECT 69.960 131.740 70.220 132.060 ;
        RECT 68.580 130.380 68.840 130.700 ;
        RECT 68.640 129.340 68.780 130.380 ;
        RECT 68.580 129.020 68.840 129.340 ;
        RECT 70.480 128.660 70.620 134.120 ;
        RECT 70.940 129.000 71.080 147.380 ;
        RECT 71.860 145.660 72.000 149.080 ;
        RECT 72.320 146.535 72.460 150.100 ;
        RECT 72.250 146.165 72.530 146.535 ;
        RECT 71.800 145.340 72.060 145.660 ;
        RECT 71.860 144.300 72.000 145.340 ;
        RECT 71.800 143.980 72.060 144.300 ;
        RECT 71.800 141.260 72.060 141.580 ;
        RECT 71.860 140.220 72.000 141.260 ;
        RECT 71.800 139.900 72.060 140.220 ;
        RECT 72.780 139.540 72.920 152.285 ;
        RECT 73.240 150.420 73.380 153.500 ;
        RECT 73.700 153.140 73.840 163.450 ;
        RECT 73.640 152.820 73.900 153.140 ;
        RECT 73.180 150.100 73.440 150.420 ;
        RECT 73.700 147.700 73.840 152.820 ;
        RECT 73.640 147.380 73.900 147.700 ;
        RECT 72.720 139.220 72.980 139.540 ;
        RECT 72.780 129.340 72.920 139.220 ;
        RECT 73.640 133.100 73.900 133.420 ;
        RECT 72.720 129.020 72.980 129.340 ;
        RECT 70.880 128.680 71.140 129.000 ;
        RECT 70.420 128.340 70.680 128.660 ;
        RECT 68.120 119.840 68.380 120.160 ;
        RECT 68.180 117.100 68.320 119.840 ;
        RECT 68.120 116.780 68.380 117.100 ;
        RECT 69.960 114.060 70.220 114.380 ;
        RECT 70.020 113.020 70.160 114.060 ;
        RECT 69.960 112.700 70.220 113.020 ;
        RECT 69.960 112.020 70.220 112.340 ;
        RECT 70.020 109.620 70.160 112.020 ;
        RECT 70.940 110.300 71.080 128.680 ;
        RECT 73.700 128.660 73.840 133.100 ;
        RECT 73.640 128.340 73.900 128.660 ;
        RECT 74.160 123.220 74.300 164.040 ;
        RECT 79.620 163.360 79.880 163.680 ;
        RECT 76.880 162.145 78.760 162.515 ;
        RECT 79.680 160.960 79.820 163.360 ;
        RECT 79.620 160.640 79.880 160.960 ;
        RECT 79.160 158.940 79.420 159.260 ;
        RECT 76.880 156.705 78.760 157.075 ;
        RECT 79.220 155.860 79.360 158.940 ;
        RECT 79.620 155.880 79.880 156.200 ;
        RECT 74.560 155.540 74.820 155.860 ;
        RECT 79.160 155.540 79.420 155.860 ;
        RECT 74.620 153.140 74.760 155.540 ;
        RECT 79.220 153.480 79.360 155.540 ;
        RECT 79.680 153.820 79.820 155.880 ;
        RECT 79.620 153.500 79.880 153.820 ;
        RECT 79.160 153.160 79.420 153.480 ;
        RECT 74.560 152.820 74.820 153.140 ;
        RECT 79.220 152.800 79.360 153.160 ;
        RECT 79.680 152.800 79.820 153.500 ;
        RECT 79.160 152.480 79.420 152.800 ;
        RECT 79.620 152.480 79.880 152.800 ;
        RECT 75.020 151.800 75.280 152.120 ;
        RECT 76.400 151.800 76.660 152.120 ;
        RECT 79.160 151.800 79.420 152.120 ;
        RECT 75.080 150.760 75.220 151.800 ;
        RECT 75.020 150.440 75.280 150.760 ;
        RECT 74.560 143.640 74.820 143.960 ;
        RECT 74.620 142.260 74.760 143.640 ;
        RECT 74.560 141.940 74.820 142.260 ;
        RECT 76.460 141.920 76.600 151.800 ;
        RECT 76.880 151.265 78.760 151.635 ;
        RECT 76.880 145.825 78.760 146.195 ;
        RECT 79.220 144.980 79.360 151.800 ;
        RECT 79.680 150.760 79.820 152.480 ;
        RECT 79.620 150.440 79.880 150.760 ;
        RECT 79.620 149.080 79.880 149.400 ;
        RECT 79.160 144.660 79.420 144.980 ;
        RECT 78.240 143.815 78.500 143.960 ;
        RECT 78.230 143.445 78.510 143.815 ;
        RECT 79.160 142.620 79.420 142.940 ;
        RECT 75.480 141.600 75.740 141.920 ;
        RECT 76.400 141.600 76.660 141.920 ;
        RECT 75.540 139.540 75.680 141.600 ;
        RECT 76.880 140.385 78.760 140.755 ;
        RECT 75.480 139.220 75.740 139.540 ;
        RECT 75.540 131.380 75.680 139.220 ;
        RECT 76.880 134.945 78.760 135.315 ;
        RECT 77.320 132.760 77.580 133.080 ;
        RECT 75.480 131.060 75.740 131.380 ;
        RECT 77.380 131.040 77.520 132.760 ;
        RECT 77.320 130.720 77.580 131.040 ;
        RECT 76.880 129.505 78.760 129.875 ;
        RECT 77.780 128.340 78.040 128.660 ;
        RECT 76.400 127.320 76.660 127.640 ;
        RECT 76.460 125.940 76.600 127.320 ;
        RECT 76.400 125.620 76.660 125.940 ;
        RECT 75.940 125.280 76.200 125.600 ;
        RECT 76.000 123.220 76.140 125.280 ;
        RECT 74.100 122.900 74.360 123.220 ;
        RECT 75.940 122.900 76.200 123.220 ;
        RECT 73.180 121.880 73.440 122.200 ;
        RECT 73.240 119.820 73.380 121.880 ;
        RECT 73.180 119.500 73.440 119.820 ;
        RECT 74.160 117.780 74.300 122.900 ;
        RECT 76.000 121.180 76.140 122.900 ;
        RECT 76.460 122.880 76.600 125.620 ;
        RECT 77.840 125.600 77.980 128.340 ;
        RECT 79.220 125.600 79.360 142.620 ;
        RECT 79.680 134.100 79.820 149.080 ;
        RECT 79.620 133.780 79.880 134.100 ;
        RECT 80.140 133.760 80.280 170.840 ;
        RECT 80.600 144.640 80.740 173.900 ;
        RECT 81.460 168.120 81.720 168.440 ;
        RECT 81.000 166.420 81.260 166.740 ;
        RECT 81.060 165.720 81.200 166.420 ;
        RECT 81.000 165.400 81.260 165.720 ;
        RECT 81.520 163.000 81.660 168.120 ;
        RECT 81.460 162.680 81.720 163.000 ;
        RECT 81.520 161.980 81.660 162.680 ;
        RECT 81.460 161.890 81.720 161.980 ;
        RECT 81.460 161.750 82.120 161.890 ;
        RECT 81.460 161.660 81.720 161.750 ;
        RECT 81.460 160.980 81.720 161.300 ;
        RECT 81.520 157.900 81.660 160.980 ;
        RECT 81.460 157.580 81.720 157.900 ;
        RECT 81.520 156.200 81.660 157.580 ;
        RECT 81.460 155.880 81.720 156.200 ;
        RECT 81.000 154.520 81.260 154.840 ;
        RECT 80.540 144.320 80.800 144.640 ;
        RECT 80.540 142.620 80.800 142.940 ;
        RECT 80.600 139.880 80.740 142.620 ;
        RECT 80.540 139.560 80.800 139.880 ;
        RECT 80.080 133.440 80.340 133.760 ;
        RECT 80.080 132.760 80.340 133.080 ;
        RECT 80.540 132.760 80.800 133.080 ;
        RECT 79.620 131.740 79.880 132.060 ;
        RECT 79.680 129.340 79.820 131.740 ;
        RECT 80.140 131.040 80.280 132.760 ;
        RECT 80.080 130.720 80.340 131.040 ;
        RECT 80.600 129.340 80.740 132.760 ;
        RECT 81.060 131.040 81.200 154.520 ;
        RECT 81.460 153.160 81.720 153.480 ;
        RECT 81.520 149.740 81.660 153.160 ;
        RECT 81.980 153.140 82.120 161.750 ;
        RECT 82.380 155.540 82.640 155.860 ;
        RECT 81.920 152.820 82.180 153.140 ;
        RECT 82.440 150.420 82.580 155.540 ;
        RECT 82.900 154.580 83.040 176.280 ;
        RECT 86.120 175.240 86.260 190.900 ;
        RECT 86.580 189.180 86.720 195.660 ;
        RECT 91.640 194.620 91.780 196.340 ;
        RECT 93.940 196.320 94.080 198.720 ;
        RECT 109.980 198.040 110.240 198.360 ;
        RECT 93.880 196.000 94.140 196.320 ;
        RECT 100.320 196.000 100.580 196.320 ;
        RECT 91.580 194.300 91.840 194.620 ;
        RECT 86.980 193.960 87.240 194.280 ;
        RECT 87.040 190.200 87.180 193.960 ;
        RECT 91.880 192.065 93.760 192.435 ;
        RECT 93.940 190.880 94.080 196.000 ;
        RECT 100.380 191.900 100.520 196.000 ;
        RECT 110.040 195.980 110.180 198.040 ;
        RECT 111.360 196.340 111.620 196.660 ;
        RECT 109.980 195.660 110.240 195.980 ;
        RECT 102.620 195.320 102.880 195.640 ;
        RECT 106.300 195.320 106.560 195.640 ;
        RECT 102.680 194.280 102.820 195.320 ;
        RECT 102.620 193.960 102.880 194.280 ;
        RECT 106.360 193.940 106.500 195.320 ;
        RECT 106.880 194.785 108.760 195.155 ;
        RECT 106.760 193.960 107.020 194.280 ;
        RECT 106.300 193.620 106.560 193.940 ;
        RECT 105.840 193.280 106.100 193.600 ;
        RECT 106.820 193.340 106.960 193.960 ;
        RECT 105.380 192.940 105.640 193.260 ;
        RECT 100.320 191.580 100.580 191.900 ;
        RECT 105.440 191.220 105.580 192.940 ;
        RECT 103.080 190.900 103.340 191.220 ;
        RECT 105.380 190.900 105.640 191.220 ;
        RECT 91.580 190.560 91.840 190.880 ;
        RECT 93.880 190.560 94.140 190.880 ;
        RECT 87.900 190.220 88.160 190.540 ;
        RECT 86.980 189.880 87.240 190.200 ;
        RECT 86.520 188.860 86.780 189.180 ;
        RECT 87.040 184.760 87.180 189.880 ;
        RECT 87.960 189.180 88.100 190.220 ;
        RECT 91.640 189.180 91.780 190.560 ;
        RECT 87.900 188.860 88.160 189.180 ;
        RECT 91.580 188.860 91.840 189.180 ;
        RECT 89.740 188.180 90.000 188.500 ;
        RECT 90.660 188.180 90.920 188.500 ;
        RECT 89.800 186.460 89.940 188.180 ;
        RECT 89.740 186.140 90.000 186.460 ;
        RECT 86.980 184.440 87.240 184.760 ;
        RECT 86.520 182.740 86.780 183.060 ;
        RECT 86.060 174.920 86.320 175.240 ;
        RECT 86.580 172.520 86.720 182.740 ;
        RECT 87.040 177.280 87.180 184.440 ;
        RECT 90.720 179.660 90.860 188.180 ;
        RECT 91.880 186.625 93.760 186.995 ;
        RECT 93.940 182.380 94.080 190.560 ;
        RECT 98.480 187.160 98.740 187.480 ;
        RECT 98.540 185.440 98.680 187.160 ;
        RECT 103.140 185.780 103.280 190.900 ;
        RECT 105.900 188.160 106.040 193.280 ;
        RECT 106.360 193.200 106.960 193.340 ;
        RECT 109.980 193.280 110.240 193.600 ;
        RECT 106.360 190.200 106.500 193.200 ;
        RECT 110.040 190.200 110.180 193.280 ;
        RECT 111.420 191.220 111.560 196.340 ;
        RECT 111.880 192.920 112.020 199.060 ;
        RECT 115.500 198.040 115.760 198.360 ;
        RECT 115.560 195.980 115.700 198.040 ;
        RECT 121.880 197.505 123.760 197.875 ;
        RECT 116.420 196.340 116.680 196.660 ;
        RECT 112.280 195.660 112.540 195.980 ;
        RECT 115.500 195.660 115.760 195.980 ;
        RECT 112.340 194.620 112.480 195.660 ;
        RECT 116.480 194.620 116.620 196.340 ;
        RECT 124.240 195.320 124.500 195.640 ;
        RECT 112.280 194.300 112.540 194.620 ;
        RECT 116.420 194.300 116.680 194.620 ;
        RECT 115.500 193.620 115.760 193.940 ;
        RECT 111.820 192.600 112.080 192.920 ;
        RECT 111.360 190.900 111.620 191.220 ;
        RECT 106.300 189.880 106.560 190.200 ;
        RECT 109.980 189.880 110.240 190.200 ;
        RECT 105.840 187.840 106.100 188.160 ;
        RECT 103.080 185.460 103.340 185.780 ;
        RECT 98.480 185.120 98.740 185.440 ;
        RECT 95.260 182.740 95.520 183.060 ;
        RECT 93.880 182.060 94.140 182.380 ;
        RECT 91.120 181.720 91.380 182.040 ;
        RECT 91.180 180.420 91.320 181.720 ;
        RECT 91.880 181.185 93.760 181.555 ;
        RECT 91.180 180.340 91.780 180.420 ;
        RECT 91.180 180.280 91.840 180.340 ;
        RECT 91.580 180.020 91.840 180.280 ;
        RECT 93.940 180.000 94.080 182.060 ;
        RECT 95.320 181.020 95.460 182.740 ;
        RECT 97.560 182.400 97.820 182.720 ;
        RECT 95.260 180.700 95.520 181.020 ;
        RECT 97.620 180.340 97.760 182.400 ;
        RECT 97.560 180.020 97.820 180.340 ;
        RECT 98.540 180.000 98.680 185.120 ;
        RECT 101.240 184.440 101.500 184.760 ;
        RECT 100.780 182.400 101.040 182.720 ;
        RECT 100.840 181.020 100.980 182.400 ;
        RECT 100.780 180.700 101.040 181.020 ;
        RECT 93.880 179.680 94.140 180.000 ;
        RECT 98.480 179.680 98.740 180.000 ;
        RECT 88.360 179.340 88.620 179.660 ;
        RECT 90.660 179.340 90.920 179.660 ;
        RECT 88.420 178.300 88.560 179.340 ;
        RECT 88.360 177.980 88.620 178.300 ;
        RECT 90.720 177.620 90.860 179.340 ;
        RECT 90.660 177.300 90.920 177.620 ;
        RECT 86.980 176.960 87.240 177.280 ;
        RECT 91.880 175.745 93.760 176.115 ;
        RECT 93.940 175.240 94.080 179.680 ;
        RECT 92.040 174.920 92.300 175.240 ;
        RECT 93.880 174.920 94.140 175.240 ;
        RECT 86.520 172.200 86.780 172.520 ;
        RECT 92.100 172.180 92.240 174.920 ;
        RECT 98.540 174.900 98.680 179.680 ;
        RECT 99.860 177.640 100.120 177.960 ;
        RECT 99.400 176.960 99.660 177.280 ;
        RECT 98.480 174.580 98.740 174.900 ;
        RECT 99.460 174.560 99.600 176.960 ;
        RECT 99.920 175.580 100.060 177.640 ;
        RECT 101.300 177.620 101.440 184.440 ;
        RECT 103.140 182.720 103.280 185.460 ;
        RECT 105.900 183.060 106.040 187.840 ;
        RECT 105.840 182.740 106.100 183.060 ;
        RECT 103.080 182.400 103.340 182.720 ;
        RECT 105.380 179.680 105.640 180.000 ;
        RECT 105.440 177.620 105.580 179.680 ;
        RECT 100.780 177.300 101.040 177.620 ;
        RECT 101.240 177.300 101.500 177.620 ;
        RECT 105.380 177.300 105.640 177.620 ;
        RECT 100.840 176.940 100.980 177.300 ;
        RECT 105.900 177.020 106.040 182.740 ;
        RECT 106.360 177.620 106.500 189.880 ;
        RECT 106.880 189.345 108.760 189.715 ;
        RECT 106.760 187.160 107.020 187.480 ;
        RECT 106.820 186.460 106.960 187.160 ;
        RECT 106.760 186.140 107.020 186.460 ;
        RECT 106.880 183.905 108.760 184.275 ;
        RECT 109.060 179.000 109.320 179.320 ;
        RECT 109.520 179.000 109.780 179.320 ;
        RECT 106.880 178.465 108.760 178.835 ;
        RECT 106.300 177.300 106.560 177.620 ;
        RECT 108.600 177.300 108.860 177.620 ;
        RECT 100.780 176.620 101.040 176.940 ;
        RECT 105.900 176.880 106.500 177.020 ;
        RECT 106.760 176.960 107.020 177.280 ;
        RECT 99.860 175.260 100.120 175.580 ;
        RECT 99.920 174.560 100.060 175.260 ;
        RECT 100.840 174.560 100.980 176.620 ;
        RECT 101.700 176.280 101.960 176.600 ;
        RECT 104.000 176.280 104.260 176.600 ;
        RECT 104.920 176.280 105.180 176.600 ;
        RECT 92.950 174.045 93.230 174.415 ;
        RECT 99.400 174.240 99.660 174.560 ;
        RECT 99.860 174.240 100.120 174.560 ;
        RECT 100.780 174.240 101.040 174.560 ;
        RECT 92.960 173.900 93.220 174.045 ;
        RECT 97.560 173.900 97.820 174.220 ;
        RECT 92.040 171.860 92.300 172.180 ;
        RECT 96.180 171.860 96.440 172.180 ;
        RECT 91.880 170.305 93.760 170.675 ;
        RECT 90.200 169.480 90.460 169.800 ;
        RECT 83.300 169.140 83.560 169.460 ;
        RECT 83.360 164.020 83.500 169.140 ;
        RECT 88.820 168.800 89.080 169.120 ;
        RECT 83.760 168.460 84.020 168.780 ;
        RECT 83.820 167.420 83.960 168.460 ;
        RECT 84.680 168.120 84.940 168.440 ;
        RECT 83.760 167.100 84.020 167.420 ;
        RECT 83.300 163.700 83.560 164.020 ;
        RECT 83.360 160.960 83.500 163.700 ;
        RECT 83.300 160.640 83.560 160.960 ;
        RECT 83.360 155.520 83.500 160.640 ;
        RECT 83.300 155.200 83.560 155.520 ;
        RECT 82.900 154.440 83.500 154.580 ;
        RECT 82.380 150.100 82.640 150.420 ;
        RECT 81.460 149.420 81.720 149.740 ;
        RECT 81.460 145.340 81.720 145.660 ;
        RECT 82.840 145.340 83.100 145.660 ;
        RECT 81.520 141.580 81.660 145.340 ;
        RECT 81.920 144.660 82.180 144.980 ;
        RECT 81.980 141.920 82.120 144.660 ;
        RECT 82.900 141.920 83.040 145.340 ;
        RECT 83.360 142.260 83.500 154.440 ;
        RECT 83.820 152.800 83.960 167.100 ;
        RECT 84.740 167.080 84.880 168.120 ;
        RECT 84.680 166.760 84.940 167.080 ;
        RECT 84.740 166.060 85.340 166.140 ;
        RECT 86.060 166.080 86.320 166.400 ;
        RECT 84.740 166.000 85.400 166.060 ;
        RECT 84.740 164.020 84.880 166.000 ;
        RECT 85.140 165.740 85.400 166.000 ;
        RECT 86.120 164.020 86.260 166.080 ;
        RECT 84.680 163.700 84.940 164.020 ;
        RECT 86.060 163.700 86.320 164.020 ;
        RECT 84.220 160.300 84.480 160.620 ;
        RECT 84.280 155.520 84.420 160.300 ;
        RECT 84.680 159.960 84.940 160.280 ;
        RECT 84.740 157.900 84.880 159.960 ;
        RECT 86.120 158.580 86.260 163.700 ;
        RECT 88.880 163.680 89.020 168.800 ;
        RECT 90.260 166.740 90.400 169.480 ;
        RECT 94.340 168.120 94.600 168.440 ;
        RECT 90.200 166.420 90.460 166.740 ;
        RECT 94.400 166.400 94.540 168.120 ;
        RECT 96.240 167.420 96.380 171.860 ;
        RECT 97.100 170.840 97.360 171.160 ;
        RECT 97.160 169.460 97.300 170.840 ;
        RECT 97.100 169.140 97.360 169.460 ;
        RECT 96.180 167.100 96.440 167.420 ;
        RECT 94.340 166.080 94.600 166.400 ;
        RECT 91.880 164.865 93.760 165.235 ;
        RECT 87.440 163.360 87.700 163.680 ;
        RECT 88.820 163.360 89.080 163.680 ;
        RECT 87.500 161.980 87.640 163.360 ;
        RECT 87.440 161.660 87.700 161.980 ;
        RECT 88.880 161.640 89.020 163.360 ;
        RECT 93.880 162.680 94.140 163.000 ;
        RECT 88.820 161.320 89.080 161.640 ;
        RECT 86.980 160.980 87.240 161.300 ;
        RECT 86.060 158.260 86.320 158.580 ;
        RECT 84.680 157.580 84.940 157.900 ;
        RECT 87.040 156.540 87.180 160.980 ;
        RECT 93.940 160.620 94.080 162.680 ;
        RECT 93.880 160.300 94.140 160.620 ;
        RECT 94.400 160.280 94.540 166.080 ;
        RECT 95.720 165.740 95.980 166.060 ;
        RECT 95.780 164.020 95.920 165.740 ;
        RECT 95.720 163.700 95.980 164.020 ;
        RECT 95.720 163.020 95.980 163.340 ;
        RECT 95.260 161.320 95.520 161.640 ;
        RECT 88.360 159.960 88.620 160.280 ;
        RECT 94.340 159.960 94.600 160.280 ;
        RECT 88.420 158.580 88.560 159.960 ;
        RECT 91.880 159.425 93.760 159.795 ;
        RECT 95.320 159.260 95.460 161.320 ;
        RECT 94.340 158.940 94.600 159.260 ;
        RECT 95.260 158.940 95.520 159.260 ;
        RECT 88.360 158.260 88.620 158.580 ;
        RECT 94.400 156.540 94.540 158.940 ;
        RECT 95.260 158.150 95.520 158.240 ;
        RECT 95.780 158.150 95.920 163.020 ;
        RECT 97.620 160.140 97.760 173.900 ;
        RECT 99.860 171.520 100.120 171.840 ;
        RECT 99.920 168.860 100.060 171.520 ;
        RECT 100.320 168.860 100.580 169.120 ;
        RECT 99.920 168.800 100.580 168.860 ;
        RECT 99.920 168.720 100.520 168.800 ;
        RECT 99.920 164.360 100.060 168.720 ;
        RECT 100.780 166.420 101.040 166.740 ;
        RECT 99.860 164.040 100.120 164.360 ;
        RECT 99.920 160.960 100.060 164.040 ;
        RECT 100.840 164.020 100.980 166.420 ;
        RECT 100.780 163.700 101.040 164.020 ;
        RECT 99.860 160.640 100.120 160.960 ;
        RECT 95.260 158.010 95.920 158.150 ;
        RECT 97.160 160.000 97.760 160.140 ;
        RECT 95.260 157.920 95.520 158.010 ;
        RECT 86.980 156.220 87.240 156.540 ;
        RECT 94.340 156.220 94.600 156.540 ;
        RECT 84.220 155.200 84.480 155.520 ;
        RECT 84.680 154.860 84.940 155.180 ;
        RECT 84.740 152.800 84.880 154.860 ;
        RECT 91.880 153.985 93.760 154.355 ;
        RECT 90.660 152.820 90.920 153.140 ;
        RECT 83.760 152.480 84.020 152.800 ;
        RECT 84.680 152.480 84.940 152.800 ;
        RECT 84.740 152.120 84.880 152.480 ;
        RECT 84.680 151.800 84.940 152.120 ;
        RECT 84.740 150.420 84.880 151.800 ;
        RECT 85.140 150.780 85.400 151.100 ;
        RECT 84.680 150.100 84.940 150.420 ;
        RECT 83.760 144.660 84.020 144.980 ;
        RECT 83.820 142.940 83.960 144.660 ;
        RECT 85.200 144.640 85.340 150.780 ;
        RECT 90.720 150.420 90.860 152.820 ;
        RECT 95.320 152.800 95.460 157.920 ;
        RECT 95.260 152.480 95.520 152.800 ;
        RECT 96.640 152.480 96.900 152.800 ;
        RECT 96.180 151.800 96.440 152.120 ;
        RECT 95.720 150.780 95.980 151.100 ;
        RECT 90.660 150.100 90.920 150.420 ;
        RECT 91.120 150.100 91.380 150.420 ;
        RECT 90.660 149.080 90.920 149.400 ;
        RECT 90.720 147.020 90.860 149.080 ;
        RECT 90.660 146.700 90.920 147.020 ;
        RECT 86.060 146.360 86.320 146.680 ;
        RECT 86.120 145.320 86.260 146.360 ;
        RECT 91.180 145.660 91.320 150.100 ;
        RECT 93.880 149.080 94.140 149.400 ;
        RECT 91.880 148.545 93.760 148.915 ;
        RECT 93.940 147.700 94.080 149.080 ;
        RECT 93.880 147.380 94.140 147.700 ;
        RECT 95.260 147.040 95.520 147.360 ;
        RECT 91.120 145.340 91.380 145.660 ;
        RECT 86.060 145.000 86.320 145.320 ;
        RECT 85.140 144.320 85.400 144.640 ;
        RECT 84.220 143.640 84.480 143.960 ;
        RECT 83.760 142.620 84.020 142.940 ;
        RECT 83.300 141.940 83.560 142.260 ;
        RECT 83.820 141.920 83.960 142.620 ;
        RECT 81.920 141.600 82.180 141.920 ;
        RECT 82.840 141.600 83.100 141.920 ;
        RECT 83.760 141.600 84.020 141.920 ;
        RECT 81.460 141.260 81.720 141.580 ;
        RECT 81.520 136.140 81.660 141.260 ;
        RECT 81.980 136.480 82.120 141.600 ;
        RECT 82.380 140.920 82.640 141.240 ;
        RECT 82.440 139.620 82.580 140.920 ;
        RECT 82.900 140.220 83.040 141.600 ;
        RECT 82.840 139.900 83.100 140.220 ;
        RECT 82.440 139.480 83.040 139.620 ;
        RECT 81.920 136.220 82.180 136.480 ;
        RECT 81.920 136.160 82.580 136.220 ;
        RECT 81.460 135.820 81.720 136.140 ;
        RECT 81.980 136.080 82.580 136.160 ;
        RECT 81.520 134.780 81.660 135.820 ;
        RECT 81.920 135.480 82.180 135.800 ;
        RECT 81.460 134.460 81.720 134.780 ;
        RECT 81.980 134.440 82.120 135.480 ;
        RECT 81.920 134.120 82.180 134.440 ;
        RECT 82.440 134.100 82.580 136.080 ;
        RECT 82.380 133.780 82.640 134.100 ;
        RECT 81.450 131.885 81.730 132.255 ;
        RECT 81.520 131.380 81.660 131.885 ;
        RECT 81.460 131.060 81.720 131.380 ;
        RECT 81.000 130.720 81.260 131.040 ;
        RECT 82.380 130.040 82.640 130.360 ;
        RECT 79.620 129.020 79.880 129.340 ;
        RECT 80.540 129.020 80.800 129.340 ;
        RECT 77.780 125.455 78.040 125.600 ;
        RECT 77.770 125.085 78.050 125.455 ;
        RECT 79.160 125.280 79.420 125.600 ;
        RECT 76.880 124.065 78.760 124.435 ;
        RECT 76.400 122.560 76.660 122.880 ;
        RECT 78.240 122.560 78.500 122.880 ;
        RECT 78.300 121.180 78.440 122.560 ;
        RECT 79.160 121.880 79.420 122.200 ;
        RECT 81.920 121.880 82.180 122.200 ;
        RECT 75.940 120.860 76.200 121.180 ;
        RECT 78.240 120.860 78.500 121.180 ;
        RECT 74.100 117.460 74.360 117.780 ;
        RECT 74.560 117.120 74.820 117.440 ;
        RECT 71.340 116.440 71.600 116.760 ;
        RECT 71.400 115.060 71.540 116.440 ;
        RECT 74.620 115.060 74.760 117.120 ;
        RECT 71.340 114.740 71.600 115.060 ;
        RECT 74.560 114.740 74.820 115.060 ;
        RECT 74.620 111.840 74.760 114.740 ;
        RECT 76.000 114.720 76.140 120.860 ;
        RECT 76.400 119.500 76.660 119.820 ;
        RECT 76.460 118.460 76.600 119.500 ;
        RECT 76.880 118.625 78.760 118.995 ;
        RECT 76.400 118.140 76.660 118.460 ;
        RECT 79.220 118.120 79.360 121.880 ;
        RECT 81.980 120.500 82.120 121.880 ;
        RECT 81.920 120.180 82.180 120.500 ;
        RECT 79.160 117.800 79.420 118.120 ;
        RECT 81.000 117.460 81.260 117.780 ;
        RECT 81.060 115.740 81.200 117.460 ;
        RECT 81.980 117.440 82.120 120.180 ;
        RECT 81.920 117.120 82.180 117.440 ;
        RECT 81.000 115.420 81.260 115.740 ;
        RECT 75.940 114.400 76.200 114.720 ;
        RECT 76.880 113.185 78.760 113.555 ;
        RECT 74.620 111.700 75.680 111.840 ;
        RECT 70.880 109.980 71.140 110.300 ;
        RECT 69.960 109.300 70.220 109.620 ;
        RECT 67.660 108.960 67.920 109.280 ;
        RECT 70.880 108.280 71.140 108.600 ;
        RECT 70.940 107.240 71.080 108.280 ;
        RECT 70.880 106.920 71.140 107.240 ;
        RECT 65.360 106.580 65.620 106.900 ;
        RECT 63.980 104.540 64.240 104.860 ;
        RECT 57.540 103.180 57.800 103.500 ;
        RECT 61.220 103.180 61.480 103.500 ;
        RECT 56.160 102.840 56.420 103.160 ;
        RECT 60.760 102.840 61.020 103.160 ;
        RECT 55.700 101.140 55.960 101.460 ;
        RECT 56.220 89.190 56.360 102.840 ;
        RECT 50.170 89.040 50.450 89.170 ;
        RECT 49.740 88.640 50.960 89.040 ;
        RECT 37.680 86.810 39.070 88.620 ;
        RECT 37.750 85.420 38.970 86.810 ;
        RECT 43.810 86.720 45.140 88.630 ;
        RECT 49.740 86.920 51.010 88.640 ;
        RECT 43.810 85.660 45.030 86.720 ;
        RECT 49.740 85.170 50.960 86.920 ;
        RECT 55.530 85.320 56.750 89.190 ;
        RECT 60.820 88.620 60.960 102.840 ;
        RECT 65.420 102.140 65.560 106.580 ;
        RECT 75.540 106.470 75.680 111.700 ;
        RECT 79.610 111.485 79.890 111.855 ;
        RECT 79.680 109.280 79.820 111.485 ;
        RECT 76.400 108.960 76.660 109.280 ;
        RECT 79.620 108.960 79.880 109.280 ;
        RECT 75.940 106.470 76.200 106.560 ;
        RECT 75.540 106.330 76.200 106.470 ;
        RECT 75.940 106.240 76.200 106.330 ;
        RECT 68.120 105.560 68.380 105.880 ;
        RECT 74.100 105.560 74.360 105.880 ;
        RECT 65.360 101.820 65.620 102.140 ;
        RECT 61.880 99.585 63.760 99.955 ;
        RECT 68.180 89.840 68.320 105.560 ;
        RECT 67.730 89.640 68.670 89.840 ;
        RECT 61.740 89.170 62.340 89.300 ;
        RECT 61.740 89.160 62.410 89.170 ;
        RECT 61.740 88.870 61.880 89.160 ;
        RECT 62.130 88.870 62.410 89.160 ;
        RECT 61.720 88.640 62.940 88.870 ;
        RECT 61.720 88.620 63.130 88.640 ;
        RECT 60.820 88.480 63.130 88.620 ;
        RECT 61.720 86.600 63.130 88.480 ;
        RECT 61.720 85.000 62.940 86.600 ;
        RECT 67.580 85.770 68.800 89.640 ;
        RECT 74.160 89.170 74.300 105.560 ;
        RECT 76.460 102.140 76.600 108.960 ;
        RECT 79.160 108.280 79.420 108.600 ;
        RECT 80.540 108.280 80.800 108.600 ;
        RECT 76.880 107.745 78.760 108.115 ;
        RECT 79.220 107.580 79.360 108.280 ;
        RECT 79.160 107.260 79.420 107.580 ;
        RECT 80.600 107.240 80.740 108.280 ;
        RECT 82.440 107.240 82.580 130.040 ;
        RECT 80.540 106.920 80.800 107.240 ;
        RECT 82.380 106.920 82.640 107.240 ;
        RECT 82.900 106.900 83.040 139.480 ;
        RECT 83.820 137.160 83.960 141.600 ;
        RECT 83.760 136.840 84.020 137.160 ;
        RECT 83.820 134.100 83.960 136.840 ;
        RECT 83.760 133.780 84.020 134.100 ;
        RECT 83.300 128.000 83.560 128.320 ;
        RECT 83.760 128.000 84.020 128.320 ;
        RECT 83.360 124.920 83.500 128.000 ;
        RECT 83.820 125.260 83.960 128.000 ;
        RECT 84.280 125.600 84.420 143.640 ;
        RECT 85.200 142.260 85.340 144.320 ;
        RECT 91.880 143.105 93.760 143.475 ;
        RECT 85.140 141.940 85.400 142.260 ;
        RECT 84.680 141.260 84.940 141.580 ;
        RECT 84.740 139.880 84.880 141.260 ;
        RECT 84.680 139.560 84.940 139.880 ;
        RECT 85.200 137.160 85.340 141.940 ;
        RECT 89.740 141.600 90.000 141.920 ;
        RECT 86.060 140.920 86.320 141.240 ;
        RECT 85.140 136.840 85.400 137.160 ;
        RECT 84.680 136.160 84.940 136.480 ;
        RECT 84.740 134.440 84.880 136.160 ;
        RECT 84.680 134.120 84.940 134.440 ;
        RECT 85.200 133.760 85.340 136.840 ;
        RECT 86.120 134.780 86.260 140.920 ;
        RECT 86.060 134.460 86.320 134.780 ;
        RECT 84.680 133.440 84.940 133.760 ;
        RECT 85.140 133.440 85.400 133.760 ;
        RECT 84.220 125.280 84.480 125.600 ;
        RECT 83.760 124.940 84.020 125.260 ;
        RECT 83.300 124.600 83.560 124.920 ;
        RECT 83.360 122.880 83.500 124.600 ;
        RECT 83.300 122.560 83.560 122.880 ;
        RECT 84.740 109.620 84.880 133.440 ;
        RECT 86.120 132.060 86.260 134.460 ;
        RECT 89.800 134.180 89.940 141.600 ;
        RECT 90.200 140.920 90.460 141.240 ;
        RECT 90.260 139.540 90.400 140.920 ;
        RECT 90.200 139.220 90.460 139.540 ;
        RECT 95.320 139.200 95.460 147.040 ;
        RECT 95.780 146.680 95.920 150.780 ;
        RECT 96.240 150.760 96.380 151.800 ;
        RECT 96.180 150.440 96.440 150.760 ;
        RECT 95.720 146.360 95.980 146.680 ;
        RECT 95.780 145.660 95.920 146.360 ;
        RECT 96.700 145.660 96.840 152.480 ;
        RECT 95.720 145.340 95.980 145.660 ;
        RECT 96.640 145.340 96.900 145.660 ;
        RECT 97.160 139.200 97.300 160.000 ;
        RECT 99.400 157.240 99.660 157.560 ;
        RECT 99.460 155.860 99.600 157.240 ;
        RECT 99.400 155.540 99.660 155.860 ;
        RECT 98.020 154.520 98.280 154.840 ;
        RECT 98.080 139.540 98.220 154.520 ;
        RECT 98.480 151.800 98.740 152.120 ;
        RECT 98.540 150.760 98.680 151.800 ;
        RECT 98.480 150.440 98.740 150.760 ;
        RECT 99.920 150.080 100.060 160.640 ;
        RECT 100.840 155.860 100.980 163.700 ;
        RECT 101.240 162.680 101.500 163.000 ;
        RECT 101.300 161.300 101.440 162.680 ;
        RECT 101.240 160.980 101.500 161.300 ;
        RECT 101.760 160.140 101.900 176.280 ;
        RECT 102.620 168.800 102.880 169.120 ;
        RECT 102.680 167.420 102.820 168.800 ;
        RECT 102.620 167.100 102.880 167.420 ;
        RECT 101.300 160.000 101.900 160.140 ;
        RECT 100.780 155.540 101.040 155.860 ;
        RECT 99.860 149.760 100.120 150.080 ;
        RECT 100.780 149.080 101.040 149.400 ;
        RECT 100.320 143.980 100.580 144.300 ;
        RECT 98.940 139.900 99.200 140.220 ;
        RECT 98.020 139.220 98.280 139.540 ;
        RECT 95.260 138.880 95.520 139.200 ;
        RECT 97.100 138.880 97.360 139.200 ;
        RECT 91.880 137.665 93.760 138.035 ;
        RECT 89.800 134.100 90.400 134.180 ;
        RECT 89.800 134.040 90.460 134.100 ;
        RECT 90.200 133.780 90.460 134.040 ;
        RECT 89.740 132.760 90.000 133.080 ;
        RECT 86.060 131.740 86.320 132.060 ;
        RECT 89.800 130.700 89.940 132.760 ;
        RECT 89.740 130.380 90.000 130.700 ;
        RECT 90.260 130.360 90.400 133.780 ;
        RECT 91.120 132.760 91.380 133.080 ;
        RECT 91.180 131.380 91.320 132.760 ;
        RECT 91.880 132.225 93.760 132.595 ;
        RECT 95.320 131.380 95.460 138.880 ;
        RECT 97.560 138.200 97.820 138.520 ;
        RECT 96.180 134.120 96.440 134.440 ;
        RECT 96.240 132.060 96.380 134.120 ;
        RECT 97.620 132.060 97.760 138.200 ;
        RECT 98.020 135.480 98.280 135.800 ;
        RECT 98.080 133.760 98.220 135.480 ;
        RECT 98.020 133.440 98.280 133.760 ;
        RECT 96.180 131.740 96.440 132.060 ;
        RECT 97.560 131.740 97.820 132.060 ;
        RECT 91.120 131.060 91.380 131.380 ;
        RECT 95.260 131.060 95.520 131.380 ;
        RECT 90.200 130.040 90.460 130.360 ;
        RECT 91.880 126.785 93.760 127.155 ;
        RECT 85.140 125.960 85.400 126.280 ;
        RECT 85.200 117.100 85.340 125.960 ;
        RECT 87.440 125.620 87.700 125.940 ;
        RECT 86.980 124.600 87.240 124.920 ;
        RECT 87.040 120.160 87.180 124.600 ;
        RECT 86.980 119.840 87.240 120.160 ;
        RECT 87.500 119.220 87.640 125.620 ;
        RECT 88.820 124.940 89.080 125.260 ;
        RECT 88.360 122.900 88.620 123.220 ;
        RECT 88.420 122.735 88.560 122.900 ;
        RECT 88.350 122.365 88.630 122.735 ;
        RECT 88.880 119.480 89.020 124.940 ;
        RECT 93.880 124.600 94.140 124.920 ;
        RECT 90.200 123.240 90.460 123.560 ;
        RECT 90.260 121.180 90.400 123.240 ;
        RECT 93.940 122.200 94.080 124.600 ;
        RECT 95.320 122.880 95.460 131.060 ;
        RECT 98.020 123.240 98.280 123.560 ;
        RECT 95.260 122.560 95.520 122.880 ;
        RECT 91.120 121.880 91.380 122.200 ;
        RECT 93.880 121.880 94.140 122.200 ;
        RECT 90.200 120.860 90.460 121.180 ;
        RECT 87.040 119.080 87.640 119.220 ;
        RECT 88.820 119.160 89.080 119.480 ;
        RECT 87.040 117.440 87.180 119.080 ;
        RECT 88.880 118.460 89.020 119.160 ;
        RECT 88.820 118.140 89.080 118.460 ;
        RECT 90.260 117.780 90.400 120.860 ;
        RECT 91.180 119.820 91.320 121.880 ;
        RECT 91.880 121.345 93.760 121.715 ;
        RECT 91.120 119.500 91.380 119.820 ;
        RECT 93.940 118.120 94.080 121.880 ;
        RECT 95.320 120.580 95.460 122.560 ;
        RECT 98.080 121.180 98.220 123.240 ;
        RECT 98.020 120.860 98.280 121.180 ;
        RECT 94.400 120.500 95.920 120.580 ;
        RECT 94.340 120.440 95.980 120.500 ;
        RECT 94.340 120.180 94.600 120.440 ;
        RECT 95.720 120.180 95.980 120.440 ;
        RECT 97.100 120.180 97.360 120.500 ;
        RECT 93.880 117.800 94.140 118.120 ;
        RECT 90.200 117.460 90.460 117.780 ;
        RECT 86.980 117.120 87.240 117.440 ;
        RECT 85.140 116.780 85.400 117.100 ;
        RECT 85.200 115.060 85.340 116.780 ;
        RECT 85.140 114.740 85.400 115.060 ;
        RECT 87.040 114.720 87.180 117.120 ;
        RECT 91.880 115.905 93.760 116.275 ;
        RECT 86.980 114.400 87.240 114.720 ;
        RECT 91.880 110.465 93.760 110.835 ;
        RECT 84.680 109.300 84.940 109.620 ;
        RECT 89.740 108.960 90.000 109.280 ;
        RECT 87.440 108.280 87.700 108.600 ;
        RECT 82.840 106.580 83.100 106.900 ;
        RECT 83.760 105.560 84.020 105.880 ;
        RECT 84.220 105.560 84.480 105.880 ;
        RECT 83.820 104.180 83.960 105.560 ;
        RECT 83.760 103.860 84.020 104.180 ;
        RECT 84.280 103.500 84.420 105.560 ;
        RECT 87.500 103.840 87.640 108.280 ;
        RECT 89.800 106.560 89.940 108.960 ;
        RECT 90.200 108.280 90.460 108.600 ;
        RECT 96.640 108.280 96.900 108.600 ;
        RECT 90.260 107.240 90.400 108.280 ;
        RECT 96.700 107.240 96.840 108.280 ;
        RECT 97.160 107.240 97.300 120.180 ;
        RECT 98.480 119.840 98.740 120.160 ;
        RECT 98.540 118.460 98.680 119.840 ;
        RECT 98.480 118.140 98.740 118.460 ;
        RECT 99.000 112.340 99.140 139.900 ;
        RECT 100.380 139.880 100.520 143.980 ;
        RECT 100.320 139.560 100.580 139.880 ;
        RECT 100.840 139.540 100.980 149.080 ;
        RECT 100.780 139.220 101.040 139.540 ;
        RECT 101.300 138.860 101.440 160.000 ;
        RECT 102.160 158.600 102.420 158.920 ;
        RECT 102.220 153.480 102.360 158.600 ;
        RECT 103.080 157.580 103.340 157.900 ;
        RECT 103.140 156.200 103.280 157.580 ;
        RECT 103.540 157.240 103.800 157.560 ;
        RECT 102.610 155.685 102.890 156.055 ;
        RECT 103.080 155.880 103.340 156.200 ;
        RECT 102.620 155.540 102.880 155.685 ;
        RECT 103.080 154.520 103.340 154.840 ;
        RECT 102.160 153.160 102.420 153.480 ;
        RECT 102.220 143.960 102.360 153.160 ;
        RECT 102.620 149.080 102.880 149.400 ;
        RECT 102.160 143.640 102.420 143.960 ;
        RECT 102.160 142.280 102.420 142.600 ;
        RECT 102.220 139.540 102.360 142.280 ;
        RECT 101.700 139.220 101.960 139.540 ;
        RECT 102.160 139.220 102.420 139.540 ;
        RECT 101.760 138.860 101.900 139.220 ;
        RECT 101.240 138.540 101.500 138.860 ;
        RECT 101.700 138.540 101.960 138.860 ;
        RECT 101.760 136.480 101.900 138.540 ;
        RECT 101.700 136.160 101.960 136.480 ;
        RECT 99.400 130.720 99.660 131.040 ;
        RECT 99.460 124.920 99.600 130.720 ;
        RECT 102.680 129.000 102.820 149.080 ;
        RECT 103.140 139.540 103.280 154.520 ;
        RECT 103.600 147.360 103.740 157.240 ;
        RECT 104.060 147.700 104.200 176.280 ;
        RECT 104.460 168.120 104.720 168.440 ;
        RECT 104.520 166.740 104.660 168.120 ;
        RECT 104.460 166.420 104.720 166.740 ;
        RECT 104.520 160.620 104.660 166.420 ;
        RECT 104.460 160.300 104.720 160.620 ;
        RECT 104.460 158.260 104.720 158.580 ;
        RECT 104.520 156.540 104.660 158.260 ;
        RECT 104.460 156.220 104.720 156.540 ;
        RECT 104.460 153.500 104.720 153.820 ;
        RECT 104.520 150.420 104.660 153.500 ;
        RECT 104.980 150.420 105.120 176.280 ;
        RECT 106.360 174.560 106.500 176.880 ;
        RECT 106.820 174.560 106.960 176.960 ;
        RECT 108.660 174.560 108.800 177.300 ;
        RECT 106.300 174.240 106.560 174.560 ;
        RECT 106.760 174.240 107.020 174.560 ;
        RECT 108.600 174.240 108.860 174.560 ;
        RECT 105.380 173.900 105.640 174.220 ;
        RECT 104.460 150.100 104.720 150.420 ;
        RECT 104.920 150.100 105.180 150.420 ;
        RECT 104.460 148.060 104.720 148.380 ;
        RECT 104.000 147.380 104.260 147.700 ;
        RECT 103.540 147.040 103.800 147.360 ;
        RECT 104.000 143.640 104.260 143.960 ;
        RECT 103.540 139.900 103.800 140.220 ;
        RECT 103.080 139.220 103.340 139.540 ;
        RECT 103.080 135.480 103.340 135.800 ;
        RECT 103.140 134.100 103.280 135.480 ;
        RECT 103.080 133.780 103.340 134.100 ;
        RECT 102.620 128.680 102.880 129.000 ;
        RECT 99.400 124.600 99.660 124.920 ;
        RECT 101.240 124.600 101.500 124.920 ;
        RECT 99.860 122.900 100.120 123.220 ;
        RECT 99.920 121.180 100.060 122.900 ;
        RECT 99.860 120.860 100.120 121.180 ;
        RECT 101.300 120.160 101.440 124.600 ;
        RECT 102.150 122.365 102.430 122.735 ;
        RECT 102.220 120.160 102.360 122.365 ;
        RECT 101.240 119.840 101.500 120.160 ;
        RECT 102.160 119.840 102.420 120.160 ;
        RECT 98.940 112.020 99.200 112.340 ;
        RECT 103.600 111.840 103.740 139.900 ;
        RECT 104.060 134.100 104.200 143.640 ;
        RECT 104.000 133.780 104.260 134.100 ;
        RECT 104.060 130.360 104.200 133.780 ;
        RECT 104.000 130.040 104.260 130.360 ;
        RECT 104.060 125.600 104.200 130.040 ;
        RECT 104.520 129.340 104.660 148.060 ;
        RECT 104.920 142.620 105.180 142.940 ;
        RECT 104.980 131.720 105.120 142.620 ;
        RECT 105.440 142.260 105.580 173.900 ;
        RECT 105.830 173.365 106.110 173.735 ;
        RECT 105.900 172.520 106.040 173.365 ;
        RECT 106.360 172.860 106.500 174.240 ;
        RECT 106.880 173.025 108.760 173.395 ;
        RECT 106.300 172.540 106.560 172.860 ;
        RECT 105.840 172.200 106.100 172.520 ;
        RECT 106.360 170.140 106.500 172.540 ;
        RECT 106.300 169.820 106.560 170.140 ;
        RECT 109.120 169.540 109.260 179.000 ;
        RECT 109.580 174.560 109.720 179.000 ;
        RECT 110.040 177.620 110.180 189.880 ;
        RECT 111.420 180.000 111.560 190.900 ;
        RECT 111.880 185.780 112.020 192.600 ;
        RECT 115.560 191.900 115.700 193.620 ;
        RECT 121.880 192.065 123.760 192.435 ;
        RECT 115.500 191.580 115.760 191.900 ;
        RECT 119.180 188.520 119.440 188.840 ;
        RECT 112.280 187.840 112.540 188.160 ;
        RECT 111.820 185.460 112.080 185.780 ;
        RECT 111.820 184.440 112.080 184.760 ;
        RECT 111.880 183.740 112.020 184.440 ;
        RECT 111.820 183.420 112.080 183.740 ;
        RECT 112.340 183.060 112.480 187.840 ;
        RECT 119.240 186.460 119.380 188.520 ;
        RECT 124.300 188.500 124.440 195.320 ;
        RECT 124.240 188.180 124.500 188.500 ;
        RECT 121.020 187.160 121.280 187.480 ;
        RECT 121.080 186.460 121.220 187.160 ;
        RECT 121.880 186.625 123.760 186.995 ;
        RECT 119.180 186.140 119.440 186.460 ;
        RECT 121.020 186.140 121.280 186.460 ;
        RECT 124.300 185.780 124.440 188.180 ;
        RECT 113.200 185.460 113.460 185.780 ;
        RECT 124.240 185.460 124.500 185.780 ;
        RECT 113.260 184.760 113.400 185.460 ;
        RECT 120.560 185.350 120.820 185.440 ;
        RECT 119.240 185.210 120.820 185.350 ;
        RECT 118.260 184.780 118.520 185.100 ;
        RECT 113.200 184.440 113.460 184.760 ;
        RECT 118.320 183.740 118.460 184.780 ;
        RECT 118.260 183.420 118.520 183.740 ;
        RECT 112.280 182.740 112.540 183.060 ;
        RECT 111.820 182.400 112.080 182.720 ;
        RECT 111.880 180.340 112.020 182.400 ;
        RECT 111.820 180.020 112.080 180.340 ;
        RECT 110.440 179.680 110.700 180.000 ;
        RECT 111.360 179.680 111.620 180.000 ;
        RECT 109.980 177.300 110.240 177.620 ;
        RECT 110.500 177.280 110.640 179.680 ;
        RECT 110.900 179.340 111.160 179.660 ;
        RECT 110.960 178.300 111.100 179.340 ;
        RECT 112.340 179.320 112.480 182.740 ;
        RECT 119.240 181.020 119.380 185.210 ;
        RECT 120.560 185.120 120.820 185.210 ;
        RECT 121.880 181.185 123.760 181.555 ;
        RECT 119.180 180.700 119.440 181.020 ;
        RECT 118.720 179.680 118.980 180.000 ;
        RECT 112.280 179.000 112.540 179.320 ;
        RECT 110.900 177.980 111.160 178.300 ;
        RECT 110.440 176.960 110.700 177.280 ;
        RECT 118.780 177.190 118.920 179.680 ;
        RECT 119.180 179.000 119.440 179.320 ;
        RECT 119.240 177.960 119.380 179.000 ;
        RECT 119.180 177.640 119.440 177.960 ;
        RECT 124.300 177.280 124.440 185.460 ;
        RECT 118.780 177.050 119.380 177.190 ;
        RECT 109.980 176.280 110.240 176.600 ;
        RECT 109.520 174.240 109.780 174.560 ;
        RECT 110.040 172.180 110.180 176.280 ;
        RECT 110.500 174.560 110.640 176.960 ;
        RECT 114.120 174.580 114.380 174.900 ;
        RECT 110.440 174.240 110.700 174.560 ;
        RECT 114.180 172.860 114.320 174.580 ;
        RECT 119.240 174.560 119.380 177.050 ;
        RECT 121.020 176.960 121.280 177.280 ;
        RECT 124.240 176.960 124.500 177.280 ;
        RECT 125.620 176.960 125.880 177.280 ;
        RECT 121.080 175.580 121.220 176.960 ;
        RECT 121.880 175.745 123.760 176.115 ;
        RECT 121.020 175.260 121.280 175.580 ;
        RECT 119.180 174.240 119.440 174.560 ;
        RECT 118.260 173.560 118.520 173.880 ;
        RECT 114.120 172.540 114.380 172.860 ;
        RECT 118.320 172.520 118.460 173.560 ;
        RECT 118.260 172.200 118.520 172.520 ;
        RECT 109.980 171.860 110.240 172.180 ;
        RECT 115.500 171.860 115.760 172.180 ;
        RECT 105.900 169.400 109.260 169.540 ;
        RECT 105.900 151.010 106.040 169.400 ;
        RECT 106.880 167.585 108.760 167.955 ;
        RECT 110.040 166.740 110.180 171.860 ;
        RECT 110.440 171.520 110.700 171.840 ;
        RECT 109.980 166.420 110.240 166.740 ;
        RECT 107.680 166.080 107.940 166.400 ;
        RECT 106.300 165.400 106.560 165.720 ;
        RECT 106.360 161.300 106.500 165.400 ;
        RECT 107.740 164.700 107.880 166.080 ;
        RECT 107.680 164.380 107.940 164.700 ;
        RECT 109.520 163.360 109.780 163.680 ;
        RECT 106.880 162.145 108.760 162.515 ;
        RECT 109.580 161.980 109.720 163.360 ;
        RECT 109.520 161.660 109.780 161.980 ;
        RECT 106.300 160.980 106.560 161.300 ;
        RECT 106.300 160.300 106.560 160.620 ;
        RECT 106.360 155.860 106.500 160.300 ;
        RECT 106.760 159.960 107.020 160.280 ;
        RECT 106.820 158.240 106.960 159.960 ;
        RECT 106.760 157.920 107.020 158.240 ;
        RECT 109.520 157.920 109.780 158.240 ;
        RECT 106.880 156.705 108.760 157.075 ;
        RECT 109.060 156.220 109.320 156.540 ;
        RECT 106.300 155.540 106.560 155.860 ;
        RECT 106.750 155.685 107.030 156.055 ;
        RECT 109.120 155.860 109.260 156.220 ;
        RECT 109.580 156.055 109.720 157.920 ;
        RECT 106.760 155.540 107.020 155.685 ;
        RECT 108.600 155.540 108.860 155.860 ;
        RECT 109.060 155.540 109.320 155.860 ;
        RECT 109.510 155.685 109.790 156.055 ;
        RECT 110.040 155.860 110.180 166.420 ;
        RECT 110.500 165.720 110.640 171.520 ;
        RECT 115.560 171.160 115.700 171.860 ;
        RECT 115.500 170.840 115.760 171.160 ;
        RECT 111.360 169.140 111.620 169.460 ;
        RECT 110.440 165.400 110.700 165.720 ;
        RECT 110.500 164.700 110.640 165.400 ;
        RECT 110.440 164.380 110.700 164.700 ;
        RECT 111.420 164.020 111.560 169.140 ;
        RECT 111.820 168.460 112.080 168.780 ;
        RECT 111.880 167.420 112.020 168.460 ;
        RECT 111.820 167.100 112.080 167.420 ;
        RECT 115.560 166.740 115.700 170.840 ;
        RECT 118.720 168.800 118.980 169.120 ;
        RECT 118.780 167.420 118.920 168.800 ;
        RECT 118.720 167.100 118.980 167.420 ;
        RECT 119.240 166.740 119.380 174.240 ;
        RECT 125.680 171.840 125.820 176.960 ;
        RECT 135.630 173.380 136.780 174.600 ;
        RECT 121.480 171.520 121.740 171.840 ;
        RECT 125.620 171.520 125.880 171.840 ;
        RECT 121.540 170.140 121.680 171.520 ;
        RECT 121.880 170.305 123.760 170.675 ;
        RECT 121.480 169.820 121.740 170.140 ;
        RECT 125.680 169.460 125.820 171.520 ;
        RECT 130.210 171.325 130.490 171.695 ;
        RECT 125.620 169.140 125.880 169.460 ;
        RECT 119.640 168.460 119.900 168.780 ;
        RECT 115.500 166.420 115.760 166.740 ;
        RECT 116.880 166.420 117.140 166.740 ;
        RECT 119.180 166.420 119.440 166.740 ;
        RECT 111.360 163.700 111.620 164.020 ;
        RECT 113.200 163.020 113.460 163.340 ;
        RECT 110.900 162.680 111.160 163.000 ;
        RECT 110.960 158.580 111.100 162.680 ;
        RECT 110.900 158.260 111.160 158.580 ;
        RECT 111.820 157.580 112.080 157.900 ;
        RECT 111.880 156.200 112.020 157.580 ;
        RECT 111.820 155.880 112.080 156.200 ;
        RECT 113.260 155.860 113.400 163.020 ;
        RECT 108.660 152.800 108.800 155.540 ;
        RECT 109.120 153.480 109.260 155.540 ;
        RECT 109.580 155.260 109.720 155.685 ;
        RECT 109.980 155.540 110.240 155.860 ;
        RECT 113.200 155.540 113.460 155.860 ;
        RECT 109.580 155.180 110.180 155.260 ;
        RECT 109.580 155.120 110.240 155.180 ;
        RECT 109.980 154.860 110.240 155.120 ;
        RECT 109.520 154.520 109.780 154.840 ;
        RECT 109.060 153.160 109.320 153.480 ;
        RECT 108.600 152.480 108.860 152.800 ;
        RECT 109.060 151.800 109.320 152.120 ;
        RECT 106.880 151.265 108.760 151.635 ;
        RECT 105.900 150.870 107.420 151.010 ;
        RECT 107.280 150.420 107.420 150.870 ;
        RECT 109.120 150.420 109.260 151.800 ;
        RECT 106.760 150.100 107.020 150.420 ;
        RECT 107.220 150.100 107.480 150.420 ;
        RECT 109.060 150.100 109.320 150.420 ;
        RECT 105.840 149.420 106.100 149.740 ;
        RECT 105.900 147.700 106.040 149.420 ;
        RECT 106.300 149.080 106.560 149.400 ;
        RECT 105.840 147.380 106.100 147.700 ;
        RECT 105.840 146.700 106.100 147.020 ;
        RECT 105.900 144.300 106.040 146.700 ;
        RECT 105.840 143.980 106.100 144.300 ;
        RECT 105.380 141.940 105.640 142.260 ;
        RECT 106.360 141.660 106.500 149.080 ;
        RECT 106.820 148.380 106.960 150.100 ;
        RECT 106.760 148.060 107.020 148.380 ;
        RECT 106.760 147.100 107.020 147.360 ;
        RECT 106.760 147.040 108.340 147.100 ;
        RECT 109.060 147.040 109.320 147.360 ;
        RECT 106.820 147.020 108.340 147.040 ;
        RECT 106.820 146.960 108.400 147.020 ;
        RECT 108.140 146.700 108.400 146.960 ;
        RECT 106.880 145.825 108.760 146.195 ;
        RECT 109.120 145.320 109.260 147.040 ;
        RECT 109.060 145.000 109.320 145.320 ;
        RECT 108.140 143.980 108.400 144.300 ;
        RECT 107.220 143.640 107.480 143.960 ;
        RECT 107.280 141.920 107.420 143.640 ;
        RECT 108.200 141.920 108.340 143.980 ;
        RECT 109.120 141.920 109.260 145.000 ;
        RECT 109.580 142.600 109.720 154.520 ;
        RECT 110.040 152.710 110.180 154.860 ;
        RECT 110.900 154.520 111.160 154.840 ;
        RECT 110.960 153.820 111.100 154.520 ;
        RECT 110.900 153.500 111.160 153.820 ;
        RECT 115.560 153.140 115.700 166.420 ;
        RECT 115.950 163.165 116.230 163.535 ;
        RECT 116.940 163.340 117.080 166.420 ;
        RECT 117.340 163.360 117.600 163.680 ;
        RECT 116.020 161.300 116.160 163.165 ;
        RECT 116.880 163.020 117.140 163.340 ;
        RECT 115.960 160.980 116.220 161.300 ;
        RECT 116.020 158.240 116.160 160.980 ;
        RECT 117.400 160.960 117.540 163.360 ;
        RECT 119.700 161.300 119.840 168.460 ;
        RECT 121.020 166.420 121.280 166.740 ;
        RECT 120.100 165.400 120.360 165.720 ;
        RECT 120.160 163.340 120.300 165.400 ;
        RECT 121.080 164.700 121.220 166.420 ;
        RECT 121.480 165.400 121.740 165.720 ;
        RECT 121.020 164.380 121.280 164.700 ;
        RECT 121.540 164.020 121.680 165.400 ;
        RECT 121.880 164.865 123.760 165.235 ;
        RECT 121.480 163.700 121.740 164.020 ;
        RECT 125.680 163.680 125.820 169.140 ;
        RECT 130.280 169.120 130.420 171.325 ;
        RECT 133.750 170.070 134.880 172.730 ;
        RECT 130.220 168.800 130.480 169.120 ;
        RECT 135.630 166.640 136.740 173.380 ;
        RECT 135.630 165.420 136.780 166.640 ;
        RECT 125.620 163.360 125.880 163.680 ;
        RECT 120.100 163.020 120.360 163.340 ;
        RECT 119.640 160.980 119.900 161.300 ;
        RECT 117.340 160.640 117.600 160.960 ;
        RECT 115.960 157.920 116.220 158.240 ;
        RECT 117.400 155.860 117.540 160.640 ;
        RECT 121.880 159.425 123.760 159.795 ;
        RECT 124.240 155.880 124.500 156.200 ;
        RECT 117.340 155.540 117.600 155.860 ;
        RECT 116.420 154.520 116.680 154.840 ;
        RECT 115.500 152.820 115.760 153.140 ;
        RECT 110.440 152.710 110.700 152.800 ;
        RECT 110.040 152.570 110.700 152.710 ;
        RECT 110.440 152.480 110.700 152.570 ;
        RECT 116.480 152.120 116.620 154.520 ;
        RECT 117.400 153.480 117.540 155.540 ;
        RECT 121.880 153.985 123.760 154.355 ;
        RECT 124.300 153.820 124.440 155.880 ;
        RECT 125.680 155.520 125.820 163.360 ;
        RECT 125.620 155.200 125.880 155.520 ;
        RECT 124.240 153.500 124.500 153.820 ;
        RECT 117.340 153.160 117.600 153.480 ;
        RECT 117.340 152.480 117.600 152.800 ;
        RECT 121.020 152.480 121.280 152.800 ;
        RECT 121.480 152.480 121.740 152.800 ;
        RECT 116.420 151.800 116.680 152.120 ;
        RECT 116.880 151.800 117.140 152.120 ;
        RECT 110.500 150.420 111.100 150.500 ;
        RECT 109.980 150.100 110.240 150.420 ;
        RECT 110.500 150.360 111.160 150.420 ;
        RECT 110.040 147.020 110.180 150.100 ;
        RECT 110.500 147.100 110.640 150.360 ;
        RECT 110.900 150.100 111.160 150.360 ;
        RECT 112.280 150.100 112.540 150.420 ;
        RECT 110.900 149.420 111.160 149.740 ;
        RECT 110.960 148.040 111.100 149.420 ;
        RECT 110.900 147.720 111.160 148.040 ;
        RECT 112.340 147.360 112.480 150.100 ;
        RECT 116.480 150.080 116.620 151.800 ;
        RECT 116.420 149.760 116.680 150.080 ;
        RECT 112.740 149.080 113.000 149.400 ;
        RECT 110.900 147.100 111.160 147.360 ;
        RECT 110.500 147.040 111.160 147.100 ;
        RECT 112.280 147.040 112.540 147.360 ;
        RECT 109.980 146.700 110.240 147.020 ;
        RECT 110.500 146.960 111.100 147.040 ;
        RECT 110.040 144.980 110.180 146.700 ;
        RECT 110.960 145.060 111.100 146.960 ;
        RECT 112.340 145.320 112.480 147.040 ;
        RECT 110.500 144.980 111.100 145.060 ;
        RECT 112.280 145.000 112.540 145.320 ;
        RECT 109.980 144.660 110.240 144.980 ;
        RECT 110.440 144.920 111.100 144.980 ;
        RECT 110.440 144.660 110.700 144.920 ;
        RECT 109.520 142.280 109.780 142.600 ;
        RECT 110.040 142.260 110.180 144.660 ;
        RECT 109.980 141.940 110.240 142.260 ;
        RECT 112.280 141.940 112.540 142.260 ;
        RECT 105.900 141.520 106.500 141.660 ;
        RECT 107.220 141.600 107.480 141.920 ;
        RECT 108.140 141.600 108.400 141.920 ;
        RECT 109.060 141.600 109.320 141.920 ;
        RECT 105.380 138.200 105.640 138.520 ;
        RECT 105.440 132.060 105.580 138.200 ;
        RECT 105.380 131.740 105.640 132.060 ;
        RECT 104.920 131.400 105.180 131.720 ;
        RECT 104.920 130.380 105.180 130.700 ;
        RECT 104.460 129.020 104.720 129.340 ;
        RECT 104.000 125.280 104.260 125.600 ;
        RECT 104.060 117.780 104.200 125.280 ;
        RECT 104.980 124.920 105.120 130.380 ;
        RECT 105.900 129.340 106.040 141.520 ;
        RECT 106.300 140.920 106.560 141.240 ;
        RECT 106.360 139.880 106.500 140.920 ;
        RECT 106.880 140.385 108.760 140.755 ;
        RECT 109.120 140.220 109.260 141.600 ;
        RECT 110.440 140.920 110.700 141.240 ;
        RECT 109.060 139.900 109.320 140.220 ;
        RECT 106.300 139.560 106.560 139.880 ;
        RECT 108.140 138.880 108.400 139.200 ;
        RECT 108.200 137.160 108.340 138.880 ;
        RECT 108.140 136.840 108.400 137.160 ;
        RECT 109.520 135.820 109.780 136.140 ;
        RECT 106.880 134.945 108.760 135.315 ;
        RECT 109.580 134.780 109.720 135.820 ;
        RECT 109.520 134.460 109.780 134.780 ;
        RECT 106.300 130.720 106.560 131.040 ;
        RECT 109.060 130.720 109.320 131.040 ;
        RECT 105.840 129.020 106.100 129.340 ;
        RECT 106.360 128.660 106.500 130.720 ;
        RECT 106.880 129.505 108.760 129.875 ;
        RECT 106.300 128.340 106.560 128.660 ;
        RECT 106.300 127.660 106.560 127.980 ;
        RECT 104.460 124.600 104.720 124.920 ;
        RECT 104.920 124.600 105.180 124.920 ;
        RECT 104.520 123.560 104.660 124.600 ;
        RECT 104.980 123.900 105.120 124.600 ;
        RECT 104.920 123.580 105.180 123.900 ;
        RECT 104.460 123.240 104.720 123.560 ;
        RECT 106.360 117.780 106.500 127.660 ;
        RECT 109.120 125.940 109.260 130.720 ;
        RECT 109.060 125.620 109.320 125.940 ;
        RECT 109.060 124.600 109.320 124.920 ;
        RECT 106.880 124.065 108.760 124.435 ;
        RECT 106.880 118.625 108.760 118.995 ;
        RECT 109.120 117.780 109.260 124.600 ;
        RECT 109.980 122.560 110.240 122.880 ;
        RECT 110.040 118.460 110.180 122.560 ;
        RECT 109.980 118.140 110.240 118.460 ;
        RECT 104.000 117.460 104.260 117.780 ;
        RECT 106.300 117.460 106.560 117.780 ;
        RECT 109.060 117.460 109.320 117.780 ;
        RECT 104.000 116.440 104.260 116.760 ;
        RECT 104.060 114.380 104.200 116.440 ;
        RECT 106.360 115.740 106.500 117.460 ;
        RECT 109.060 116.440 109.320 116.760 ;
        RECT 106.300 115.420 106.560 115.740 ;
        RECT 104.000 114.060 104.260 114.380 ;
        RECT 106.880 113.185 108.760 113.555 ;
        RECT 109.120 112.340 109.260 116.440 ;
        RECT 109.520 114.400 109.780 114.720 ;
        RECT 109.580 113.020 109.720 114.400 ;
        RECT 109.520 112.700 109.780 113.020 ;
        RECT 109.060 112.020 109.320 112.340 ;
        RECT 103.600 111.700 104.200 111.840 ;
        RECT 99.860 111.000 100.120 111.320 ;
        RECT 99.920 109.620 100.060 111.000 ;
        RECT 98.020 109.300 98.280 109.620 ;
        RECT 99.860 109.300 100.120 109.620 ;
        RECT 97.560 108.620 97.820 108.940 ;
        RECT 97.620 107.580 97.760 108.620 ;
        RECT 97.560 107.260 97.820 107.580 ;
        RECT 90.200 106.920 90.460 107.240 ;
        RECT 96.640 106.920 96.900 107.240 ;
        RECT 97.100 106.920 97.360 107.240 ;
        RECT 89.740 106.240 90.000 106.560 ;
        RECT 87.900 105.560 88.160 105.880 ;
        RECT 93.880 105.560 94.140 105.880 ;
        RECT 87.960 104.180 88.100 105.560 ;
        RECT 91.880 105.025 93.760 105.395 ;
        RECT 87.900 103.860 88.160 104.180 ;
        RECT 87.440 103.520 87.700 103.840 ;
        RECT 84.220 103.180 84.480 103.500 ;
        RECT 80.080 102.840 80.340 103.160 ;
        RECT 85.600 102.840 85.860 103.160 ;
        RECT 76.880 102.305 78.760 102.675 ;
        RECT 76.400 101.820 76.660 102.140 ;
        RECT 80.140 89.170 80.280 102.840 ;
        RECT 74.090 88.160 74.370 89.170 ;
        RECT 80.070 88.180 80.350 89.170 ;
        RECT 85.660 88.620 85.800 102.840 ;
        RECT 91.880 99.585 93.760 99.955 ;
        RECT 86.050 88.620 86.330 89.170 ;
        RECT 85.660 88.480 86.330 88.620 ;
        RECT 73.850 84.290 75.070 88.160 ;
        RECT 79.730 84.310 80.950 88.180 ;
        RECT 86.050 87.970 86.330 88.480 ;
        RECT 92.030 88.620 92.310 89.170 ;
        RECT 93.940 88.620 94.080 105.560 ;
        RECT 97.160 104.180 97.300 106.920 ;
        RECT 97.100 103.860 97.360 104.180 ;
        RECT 98.080 89.170 98.220 109.300 ;
        RECT 104.060 109.280 104.200 111.700 ;
        RECT 109.520 109.300 109.780 109.620 ;
        RECT 104.000 108.960 104.260 109.280 ;
        RECT 99.400 108.620 99.660 108.940 ;
        RECT 99.460 106.900 99.600 108.620 ;
        RECT 103.540 108.280 103.800 108.600 ;
        RECT 105.840 108.280 106.100 108.600 ;
        RECT 106.300 108.280 106.560 108.600 ;
        RECT 103.600 107.240 103.740 108.280 ;
        RECT 105.900 107.240 106.040 108.280 ;
        RECT 103.540 106.920 103.800 107.240 ;
        RECT 105.840 106.920 106.100 107.240 ;
        RECT 99.400 106.580 99.660 106.900 ;
        RECT 104.000 105.560 104.260 105.880 ;
        RECT 104.060 89.170 104.200 105.560 ;
        RECT 106.360 103.840 106.500 108.280 ;
        RECT 106.880 107.745 108.760 108.115 ;
        RECT 109.580 106.560 109.720 109.300 ;
        RECT 110.500 106.900 110.640 140.920 ;
        RECT 112.340 139.540 112.480 141.940 ;
        RECT 112.280 139.220 112.540 139.540 ;
        RECT 112.800 138.940 112.940 149.080 ;
        RECT 116.480 147.360 116.620 149.760 ;
        RECT 116.940 147.700 117.080 151.800 ;
        RECT 117.400 147.700 117.540 152.480 ;
        RECT 120.100 151.800 120.360 152.120 ;
        RECT 120.160 150.760 120.300 151.800 ;
        RECT 120.560 150.780 120.820 151.100 ;
        RECT 120.100 150.440 120.360 150.760 ;
        RECT 119.640 149.420 119.900 149.740 ;
        RECT 118.260 149.080 118.520 149.400 ;
        RECT 116.880 147.380 117.140 147.700 ;
        RECT 117.340 147.380 117.600 147.700 ;
        RECT 116.420 147.040 116.680 147.360 ;
        RECT 114.120 144.320 114.380 144.640 ;
        RECT 114.180 141.920 114.320 144.320 ;
        RECT 117.400 142.940 117.540 147.380 ;
        RECT 118.320 146.680 118.460 149.080 ;
        RECT 118.260 146.360 118.520 146.680 ;
        RECT 117.340 142.620 117.600 142.940 ;
        RECT 115.960 142.280 116.220 142.600 ;
        RECT 114.120 141.600 114.380 141.920 ;
        RECT 113.200 140.920 113.460 141.240 ;
        RECT 113.260 139.540 113.400 140.920 ;
        RECT 114.180 140.220 114.320 141.600 ;
        RECT 114.580 141.260 114.840 141.580 ;
        RECT 114.120 139.900 114.380 140.220 ;
        RECT 114.640 139.880 114.780 141.260 ;
        RECT 114.580 139.560 114.840 139.880 ;
        RECT 113.200 139.220 113.460 139.540 ;
        RECT 112.800 138.800 113.400 138.940 ;
        RECT 111.360 138.200 111.620 138.520 ;
        RECT 111.420 134.100 111.560 138.200 ;
        RECT 112.280 136.500 112.540 136.820 ;
        RECT 111.820 136.160 112.080 136.480 ;
        RECT 111.360 133.780 111.620 134.100 ;
        RECT 111.880 133.760 112.020 136.160 ;
        RECT 112.340 134.780 112.480 136.500 ;
        RECT 112.280 134.460 112.540 134.780 ;
        RECT 111.820 133.440 112.080 133.760 ;
        RECT 112.740 128.000 113.000 128.320 ;
        RECT 111.820 122.560 112.080 122.880 ;
        RECT 111.880 119.820 112.020 122.560 ;
        RECT 112.800 120.160 112.940 128.000 ;
        RECT 112.740 119.840 113.000 120.160 ;
        RECT 111.820 119.500 112.080 119.820 ;
        RECT 111.880 115.060 112.020 119.500 ;
        RECT 112.800 118.460 112.940 119.840 ;
        RECT 112.740 118.140 113.000 118.460 ;
        RECT 112.800 115.740 112.940 118.140 ;
        RECT 112.740 115.420 113.000 115.740 ;
        RECT 111.820 114.740 112.080 115.060 ;
        RECT 113.260 111.840 113.400 138.800 ;
        RECT 114.640 137.500 114.780 139.560 ;
        RECT 115.500 139.220 115.760 139.540 ;
        RECT 114.580 137.180 114.840 137.500 ;
        RECT 115.560 136.140 115.700 139.220 ;
        RECT 115.500 135.820 115.760 136.140 ;
        RECT 116.020 134.100 116.160 142.280 ;
        RECT 118.320 141.920 118.460 146.360 ;
        RECT 118.260 141.600 118.520 141.920 ;
        RECT 115.960 133.780 116.220 134.100 ;
        RECT 117.340 128.680 117.600 129.000 ;
        RECT 116.880 128.340 117.140 128.660 ;
        RECT 115.500 128.000 115.760 128.320 ;
        RECT 115.560 126.280 115.700 128.000 ;
        RECT 115.500 125.960 115.760 126.280 ;
        RECT 113.660 125.280 113.920 125.600 ;
        RECT 113.720 122.880 113.860 125.280 ;
        RECT 113.660 122.560 113.920 122.880 ;
        RECT 113.720 117.780 113.860 122.560 ;
        RECT 115.560 120.500 115.700 125.960 ;
        RECT 116.940 125.940 117.080 128.340 ;
        RECT 116.880 125.620 117.140 125.940 ;
        RECT 117.400 123.900 117.540 128.680 ;
        RECT 118.260 127.320 118.520 127.640 ;
        RECT 117.340 123.580 117.600 123.900 ;
        RECT 115.500 120.180 115.760 120.500 ;
        RECT 117.400 120.160 117.540 123.580 ;
        RECT 118.320 120.160 118.460 127.320 ;
        RECT 119.180 122.560 119.440 122.880 ;
        RECT 117.340 119.840 117.600 120.160 ;
        RECT 118.260 119.840 118.520 120.160 ;
        RECT 119.240 119.480 119.380 122.560 ;
        RECT 119.180 119.160 119.440 119.480 ;
        RECT 113.660 117.460 113.920 117.780 ;
        RECT 117.340 116.440 117.600 116.760 ;
        RECT 117.400 114.380 117.540 116.440 ;
        RECT 119.240 115.060 119.380 119.160 ;
        RECT 119.180 114.740 119.440 115.060 ;
        RECT 117.340 114.060 117.600 114.380 ;
        RECT 118.720 112.700 118.980 113.020 ;
        RECT 112.800 111.700 113.400 111.840 ;
        RECT 111.820 108.620 112.080 108.940 ;
        RECT 112.280 108.620 112.540 108.940 ;
        RECT 111.880 106.900 112.020 108.620 ;
        RECT 112.340 107.580 112.480 108.620 ;
        RECT 112.280 107.260 112.540 107.580 ;
        RECT 112.800 106.900 112.940 111.700 ;
        RECT 118.780 107.240 118.920 112.700 ;
        RECT 119.700 112.680 119.840 149.420 ;
        RECT 120.100 141.600 120.360 141.920 ;
        RECT 120.160 140.220 120.300 141.600 ;
        RECT 120.100 139.900 120.360 140.220 ;
        RECT 120.100 116.440 120.360 116.760 ;
        RECT 120.160 115.060 120.300 116.440 ;
        RECT 120.100 114.740 120.360 115.060 ;
        RECT 119.640 112.360 119.900 112.680 ;
        RECT 120.620 112.340 120.760 150.780 ;
        RECT 121.080 141.920 121.220 152.480 ;
        RECT 121.540 148.380 121.680 152.480 ;
        RECT 123.780 151.800 124.040 152.120 ;
        RECT 123.840 150.420 123.980 151.800 ;
        RECT 125.680 150.420 125.820 155.200 ;
        RECT 123.780 150.100 124.040 150.420 ;
        RECT 125.620 150.100 125.880 150.420 ;
        RECT 121.880 148.545 123.760 148.915 ;
        RECT 121.480 148.060 121.740 148.380 ;
        RECT 121.880 143.105 123.760 143.475 ;
        RECT 121.020 141.600 121.280 141.920 ;
        RECT 121.020 140.920 121.280 141.240 ;
        RECT 135.630 141.200 136.780 141.270 ;
        RECT 121.080 139.880 121.220 140.920 ;
        RECT 135.630 140.180 136.800 141.200 ;
        RECT 121.020 139.560 121.280 139.880 ;
        RECT 125.620 138.880 125.880 139.200 ;
        RECT 121.880 137.665 123.760 138.035 ;
        RECT 125.680 136.820 125.820 138.880 ;
        RECT 129.140 138.175 134.100 139.455 ;
        RECT 123.320 136.500 123.580 136.820 ;
        RECT 125.620 136.500 125.880 136.820 ;
        RECT 123.380 134.780 123.520 136.500 ;
        RECT 123.320 134.460 123.580 134.780 ;
        RECT 121.880 132.225 123.760 132.595 ;
        RECT 121.880 126.785 123.760 127.155 ;
        RECT 125.680 125.600 125.820 136.500 ;
        RECT 135.640 133.320 136.800 140.180 ;
        RECT 121.480 125.280 121.740 125.600 ;
        RECT 125.620 125.280 125.880 125.600 ;
        RECT 121.540 121.180 121.680 125.280 ;
        RECT 125.680 123.220 125.820 125.280 ;
        RECT 124.700 122.900 124.960 123.220 ;
        RECT 125.620 122.900 125.880 123.220 ;
        RECT 121.880 121.345 123.760 121.715 ;
        RECT 124.760 121.180 124.900 122.900 ;
        RECT 121.480 120.860 121.740 121.180 ;
        RECT 124.700 120.860 124.960 121.180 ;
        RECT 121.880 115.905 123.760 116.275 ;
        RECT 126.080 114.400 126.340 114.720 ;
        RECT 120.560 112.020 120.820 112.340 ;
        RECT 124.700 111.000 124.960 111.320 ;
        RECT 121.880 110.465 123.760 110.835 ;
        RECT 124.760 109.620 124.900 111.000 ;
        RECT 126.140 109.620 126.280 114.400 ;
        RECT 121.480 109.300 121.740 109.620 ;
        RECT 124.700 109.300 124.960 109.620 ;
        RECT 126.080 109.300 126.340 109.620 ;
        RECT 121.020 108.280 121.280 108.600 ;
        RECT 121.080 107.240 121.220 108.280 ;
        RECT 118.720 106.920 118.980 107.240 ;
        RECT 121.020 106.920 121.280 107.240 ;
        RECT 110.440 106.580 110.700 106.900 ;
        RECT 111.820 106.580 112.080 106.900 ;
        RECT 112.740 106.580 113.000 106.900 ;
        RECT 109.520 106.240 109.780 106.560 ;
        RECT 112.280 106.240 112.540 106.560 ;
        RECT 111.820 105.560 112.080 105.880 ;
        RECT 111.880 104.180 112.020 105.560 ;
        RECT 112.340 104.940 112.480 106.240 ;
        RECT 114.120 105.560 114.380 105.880 ;
        RECT 115.500 105.560 115.760 105.880 ;
        RECT 112.340 104.860 112.940 104.940 ;
        RECT 112.340 104.800 113.000 104.860 ;
        RECT 112.740 104.540 113.000 104.800 ;
        RECT 114.180 104.180 114.320 105.560 ;
        RECT 111.820 103.860 112.080 104.180 ;
        RECT 114.120 103.860 114.380 104.180 ;
        RECT 115.560 103.840 115.700 105.560 ;
        RECT 106.300 103.520 106.560 103.840 ;
        RECT 115.500 103.520 115.760 103.840 ;
        RECT 109.980 102.840 110.240 103.160 ;
        RECT 115.960 102.840 116.220 103.160 ;
        RECT 106.880 102.305 108.760 102.675 ;
        RECT 110.040 89.290 110.180 102.840 ;
        RECT 116.020 89.570 116.160 102.840 ;
        RECT 121.540 98.820 121.680 109.300 ;
        RECT 126.140 106.560 126.280 109.300 ;
        RECT 124.700 106.240 124.960 106.560 ;
        RECT 126.080 106.240 126.340 106.560 ;
        RECT 121.880 105.025 123.760 105.395 ;
        RECT 124.760 104.180 124.900 106.240 ;
        RECT 126.530 106.045 126.810 106.415 ;
        RECT 124.700 103.860 124.960 104.180 ;
        RECT 126.600 103.840 126.740 106.045 ;
        RECT 127.920 105.560 128.180 105.880 ;
        RECT 129.750 105.580 133.160 106.650 ;
        RECT 126.540 103.520 126.800 103.840 ;
        RECT 125.160 102.840 125.420 103.160 ;
        RECT 125.220 102.140 125.360 102.840 ;
        RECT 125.160 101.820 125.420 102.140 ;
        RECT 121.880 99.585 123.760 99.955 ;
        RECT 121.540 98.680 122.140 98.820 ;
        RECT 122.000 89.570 122.140 98.680 ;
        RECT 92.030 88.480 94.080 88.620 ;
        RECT 98.010 88.500 98.290 89.170 ;
        RECT 103.990 88.610 104.270 89.170 ;
        RECT 92.030 88.320 92.310 88.480 ;
        RECT 74.090 80.440 74.370 84.290 ;
        RECT 20.140 80.160 74.370 80.440 ;
        RECT 20.140 75.650 20.420 80.160 ;
        RECT 80.070 79.800 80.350 84.310 ;
        RECT 85.470 84.100 86.690 87.970 ;
        RECT 91.460 84.500 92.680 88.320 ;
        RECT 97.600 84.630 98.820 88.500 ;
        RECT 103.650 84.740 104.870 88.610 ;
        RECT 109.620 85.420 110.840 89.290 ;
        RECT 115.740 85.700 116.960 89.570 ;
        RECT 121.520 85.700 122.740 89.570 ;
        RECT 127.980 89.380 128.120 105.560 ;
        RECT 31.380 79.520 80.350 79.800 ;
        RECT 31.380 75.850 31.660 79.520 ;
        RECT 86.050 79.170 86.330 84.100 ;
        RECT 42.510 78.890 86.330 79.170 ;
        RECT 3.960 71.320 6.050 73.240 ;
        RECT 19.330 73.120 21.890 75.650 ;
        RECT 28.185 73.180 30.255 74.460 ;
        RECT 30.670 73.320 33.230 75.850 ;
        RECT 42.510 75.750 42.790 78.890 ;
        RECT 92.030 78.570 92.310 84.500 ;
        RECT 53.830 78.290 92.310 78.570 ;
        RECT 53.830 75.820 54.110 78.290 ;
        RECT 98.010 77.990 98.290 84.630 ;
        RECT 64.900 77.710 98.290 77.990 ;
        RECT 19.005 71.800 19.865 72.640 ;
        RECT 15.560 68.610 16.990 71.210 ;
        RECT 19.305 68.570 19.845 71.800 ;
        RECT 20.145 70.600 20.555 73.120 ;
        RECT 30.205 71.810 31.065 72.650 ;
        RECT 19.325 47.770 19.825 68.570 ;
        RECT 20.165 49.090 20.555 70.600 ;
        RECT 20.955 70.010 21.845 70.740 ;
        RECT 21.055 65.190 21.315 70.010 ;
        RECT 22.695 68.620 25.405 69.470 ;
        RECT 22.895 65.840 24.825 68.620 ;
        RECT 30.505 68.580 31.045 71.810 ;
        RECT 31.345 70.610 31.755 73.320 ;
        RECT 39.475 73.150 41.545 74.430 ;
        RECT 41.910 73.220 44.470 75.750 ;
        RECT 41.425 71.780 42.285 72.620 ;
        RECT 27.795 67.130 28.915 67.810 ;
        RECT 28.075 65.850 28.745 67.130 ;
        RECT 21.455 65.460 26.505 65.840 ;
        RECT 27.865 65.440 28.915 65.850 ;
        RECT 21.055 63.640 21.435 65.190 ;
        RECT 21.175 55.800 21.435 63.640 ;
        RECT 26.485 63.200 26.755 65.240 ;
        RECT 27.615 63.200 27.885 65.200 ;
        RECT 26.485 56.510 27.885 63.200 ;
        RECT 21.085 55.290 21.445 55.800 ;
        RECT 21.065 54.860 21.445 55.290 ;
        RECT 26.485 55.190 26.755 56.510 ;
        RECT 27.615 55.150 27.885 56.510 ;
        RECT 28.885 55.260 29.205 65.190 ;
        RECT 28.885 55.200 29.215 55.260 ;
        RECT 21.065 54.580 21.315 54.860 ;
        RECT 20.865 54.180 25.505 54.580 ;
        RECT 26.405 54.290 27.535 54.300 ;
        RECT 28.895 54.290 29.215 55.200 ;
        RECT 21.065 52.060 21.315 54.180 ;
        RECT 25.765 53.490 26.125 54.110 ;
        RECT 25.845 52.610 26.105 53.490 ;
        RECT 26.385 53.240 29.215 54.290 ;
        RECT 25.675 52.230 26.205 52.610 ;
        RECT 21.065 51.970 21.565 52.060 ;
        RECT 21.055 51.240 21.565 51.970 ;
        RECT 21.295 50.240 21.565 51.240 ;
        RECT 22.205 50.990 22.475 51.940 ;
        RECT 22.205 50.840 22.675 50.990 ;
        RECT 22.205 50.160 22.765 50.840 ;
        RECT 22.285 50.150 22.765 50.160 ;
        RECT 21.575 49.620 22.195 49.980 ;
        RECT 21.615 49.090 22.045 49.620 ;
        RECT 20.165 48.670 22.045 49.090 ;
        RECT 22.535 48.960 22.765 50.150 ;
        RECT 21.615 47.800 22.045 48.670 ;
        RECT 22.455 48.360 22.835 48.960 ;
        RECT 19.325 47.060 20.015 47.770 ;
        RECT 21.435 47.440 22.055 47.800 ;
        RECT 21.135 47.060 21.425 47.250 ;
        RECT 19.325 46.620 21.425 47.060 ;
        RECT 19.325 46.600 20.015 46.620 ;
        RECT 21.135 46.380 21.425 46.620 ;
        RECT 22.055 46.990 22.325 47.240 ;
        RECT 22.535 46.990 22.765 48.360 ;
        RECT 25.355 47.010 25.685 52.030 ;
        RECT 26.405 52.020 27.535 53.240 ;
        RECT 28.895 53.220 29.215 53.240 ;
        RECT 22.055 46.880 22.765 46.990 ;
        RECT 25.345 46.960 25.685 47.010 ;
        RECT 26.235 47.780 27.615 52.020 ;
        RECT 22.055 46.570 22.715 46.880 ;
        RECT 22.055 46.400 22.325 46.570 ;
        RECT 25.345 45.000 25.625 46.960 ;
        RECT 26.235 46.920 26.535 47.780 ;
        RECT 27.315 46.920 27.615 47.780 ;
        RECT 28.165 46.920 28.495 51.990 ;
        RECT 27.565 46.380 28.045 46.760 ;
        RECT 27.665 45.760 27.915 46.380 ;
        RECT 27.565 45.160 27.945 45.760 ;
        RECT 24.825 44.230 25.925 45.000 ;
        RECT 28.215 44.930 28.495 46.920 ;
        RECT 30.525 47.780 31.025 68.580 ;
        RECT 31.365 49.100 31.755 70.610 ;
        RECT 32.155 70.020 33.045 70.750 ;
        RECT 32.255 65.200 32.515 70.020 ;
        RECT 33.895 68.630 36.605 69.480 ;
        RECT 34.095 65.850 36.025 68.630 ;
        RECT 41.725 68.550 42.265 71.780 ;
        RECT 42.565 70.580 42.975 73.220 ;
        RECT 50.055 73.090 52.125 74.370 ;
        RECT 53.150 73.290 55.710 75.820 ;
        RECT 64.900 75.810 65.180 77.710 ;
        RECT 103.990 77.230 104.270 84.740 ;
        RECT 76.140 76.950 104.270 77.230 ;
        RECT 52.675 71.760 53.535 72.600 ;
        RECT 38.995 67.140 40.115 67.820 ;
        RECT 39.275 65.860 39.945 67.140 ;
        RECT 32.655 65.470 37.705 65.850 ;
        RECT 39.065 65.450 40.115 65.860 ;
        RECT 32.255 63.650 32.635 65.200 ;
        RECT 32.375 55.810 32.635 63.650 ;
        RECT 37.685 63.210 37.955 65.250 ;
        RECT 38.815 63.210 39.085 65.210 ;
        RECT 37.685 56.520 39.085 63.210 ;
        RECT 32.285 55.300 32.645 55.810 ;
        RECT 32.265 54.870 32.645 55.300 ;
        RECT 37.685 55.200 37.955 56.520 ;
        RECT 38.815 55.160 39.085 56.520 ;
        RECT 40.085 55.270 40.405 65.200 ;
        RECT 40.085 55.210 40.415 55.270 ;
        RECT 32.265 54.590 32.515 54.870 ;
        RECT 32.065 54.190 36.705 54.590 ;
        RECT 37.605 54.300 38.735 54.310 ;
        RECT 40.095 54.300 40.415 55.210 ;
        RECT 32.265 52.070 32.515 54.190 ;
        RECT 36.965 53.500 37.325 54.120 ;
        RECT 37.045 52.620 37.305 53.500 ;
        RECT 37.585 53.250 40.415 54.300 ;
        RECT 36.875 52.240 37.405 52.620 ;
        RECT 32.265 51.980 32.765 52.070 ;
        RECT 32.255 51.250 32.765 51.980 ;
        RECT 32.495 50.250 32.765 51.250 ;
        RECT 33.405 51.000 33.675 51.950 ;
        RECT 33.405 50.850 33.875 51.000 ;
        RECT 33.405 50.170 33.965 50.850 ;
        RECT 33.485 50.160 33.965 50.170 ;
        RECT 32.775 49.630 33.395 49.990 ;
        RECT 32.815 49.100 33.245 49.630 ;
        RECT 31.365 48.680 33.245 49.100 ;
        RECT 33.735 48.970 33.965 50.160 ;
        RECT 32.815 47.810 33.245 48.680 ;
        RECT 33.655 48.370 34.035 48.970 ;
        RECT 30.525 47.070 31.215 47.780 ;
        RECT 32.635 47.450 33.255 47.810 ;
        RECT 32.335 47.070 32.625 47.260 ;
        RECT 30.525 46.630 32.625 47.070 ;
        RECT 30.525 46.610 31.215 46.630 ;
        RECT 32.335 46.390 32.625 46.630 ;
        RECT 33.255 47.000 33.525 47.250 ;
        RECT 33.735 47.000 33.965 48.370 ;
        RECT 36.555 47.020 36.885 52.040 ;
        RECT 37.605 52.030 38.735 53.250 ;
        RECT 40.095 53.230 40.415 53.250 ;
        RECT 33.255 46.890 33.965 47.000 ;
        RECT 36.545 46.970 36.885 47.020 ;
        RECT 37.435 47.790 38.815 52.030 ;
        RECT 33.255 46.580 33.915 46.890 ;
        RECT 33.255 46.410 33.525 46.580 ;
        RECT 36.545 45.010 36.825 46.970 ;
        RECT 37.435 46.930 37.735 47.790 ;
        RECT 38.515 46.930 38.815 47.790 ;
        RECT 39.365 46.930 39.695 52.000 ;
        RECT 38.765 46.390 39.245 46.770 ;
        RECT 38.865 45.770 39.115 46.390 ;
        RECT 38.765 45.170 39.145 45.770 ;
        RECT 28.215 43.200 28.515 44.930 ;
        RECT 36.025 44.240 37.125 45.010 ;
        RECT 39.415 44.940 39.695 46.930 ;
        RECT 41.745 47.750 42.245 68.550 ;
        RECT 42.585 49.070 42.975 70.580 ;
        RECT 43.375 69.990 44.265 70.720 ;
        RECT 43.475 65.170 43.735 69.990 ;
        RECT 45.115 68.600 47.825 69.450 ;
        RECT 45.315 65.820 47.245 68.600 ;
        RECT 52.975 68.530 53.515 71.760 ;
        RECT 53.815 70.560 54.225 73.290 ;
        RECT 61.475 73.120 63.545 74.400 ;
        RECT 64.400 73.280 66.960 75.810 ;
        RECT 76.140 75.740 76.420 76.950 ;
        RECT 109.970 76.610 110.250 85.420 ;
        RECT 87.580 76.330 110.250 76.610 ;
        RECT 87.580 75.760 87.860 76.330 ;
        RECT 115.950 76.030 116.230 85.700 ;
        RECT 98.850 75.840 116.230 76.030 ;
        RECT 63.895 71.750 64.755 72.590 ;
        RECT 50.215 67.110 51.335 67.790 ;
        RECT 50.495 65.830 51.165 67.110 ;
        RECT 43.875 65.440 48.925 65.820 ;
        RECT 50.285 65.420 51.335 65.830 ;
        RECT 43.475 63.620 43.855 65.170 ;
        RECT 43.595 55.780 43.855 63.620 ;
        RECT 48.905 63.180 49.175 65.220 ;
        RECT 50.035 63.180 50.305 65.180 ;
        RECT 48.905 56.490 50.305 63.180 ;
        RECT 43.505 55.270 43.865 55.780 ;
        RECT 43.485 54.840 43.865 55.270 ;
        RECT 48.905 55.170 49.175 56.490 ;
        RECT 50.035 55.130 50.305 56.490 ;
        RECT 51.305 55.240 51.625 65.170 ;
        RECT 51.305 55.180 51.635 55.240 ;
        RECT 43.485 54.560 43.735 54.840 ;
        RECT 43.285 54.160 47.925 54.560 ;
        RECT 48.825 54.270 49.955 54.280 ;
        RECT 51.315 54.270 51.635 55.180 ;
        RECT 43.485 52.040 43.735 54.160 ;
        RECT 48.185 53.470 48.545 54.090 ;
        RECT 48.265 52.590 48.525 53.470 ;
        RECT 48.805 53.220 51.635 54.270 ;
        RECT 48.095 52.210 48.625 52.590 ;
        RECT 43.485 51.950 43.985 52.040 ;
        RECT 43.475 51.220 43.985 51.950 ;
        RECT 43.715 50.220 43.985 51.220 ;
        RECT 44.625 50.970 44.895 51.920 ;
        RECT 44.625 50.820 45.095 50.970 ;
        RECT 44.625 50.140 45.185 50.820 ;
        RECT 44.705 50.130 45.185 50.140 ;
        RECT 43.995 49.600 44.615 49.960 ;
        RECT 44.035 49.070 44.465 49.600 ;
        RECT 42.585 48.650 44.465 49.070 ;
        RECT 44.955 48.940 45.185 50.130 ;
        RECT 44.035 47.780 44.465 48.650 ;
        RECT 44.875 48.340 45.255 48.940 ;
        RECT 41.745 47.040 42.435 47.750 ;
        RECT 43.855 47.420 44.475 47.780 ;
        RECT 43.555 47.040 43.845 47.230 ;
        RECT 41.745 46.600 43.845 47.040 ;
        RECT 41.745 46.580 42.435 46.600 ;
        RECT 43.555 46.360 43.845 46.600 ;
        RECT 44.475 46.970 44.745 47.220 ;
        RECT 44.955 46.970 45.185 48.340 ;
        RECT 47.775 46.990 48.105 52.010 ;
        RECT 48.825 52.000 49.955 53.220 ;
        RECT 51.315 53.200 51.635 53.220 ;
        RECT 44.475 46.860 45.185 46.970 ;
        RECT 47.765 46.940 48.105 46.990 ;
        RECT 48.655 47.760 50.035 52.000 ;
        RECT 44.475 46.550 45.135 46.860 ;
        RECT 44.475 46.380 44.745 46.550 ;
        RECT 47.765 44.980 48.045 46.940 ;
        RECT 48.655 46.900 48.955 47.760 ;
        RECT 49.735 46.900 50.035 47.760 ;
        RECT 50.585 46.900 50.915 51.970 ;
        RECT 49.985 46.360 50.465 46.740 ;
        RECT 50.085 45.740 50.335 46.360 ;
        RECT 49.985 45.140 50.365 45.740 ;
        RECT 39.415 43.210 39.715 44.940 ;
        RECT 47.245 44.210 48.345 44.980 ;
        RECT 50.635 44.910 50.915 46.900 ;
        RECT 52.995 47.730 53.495 68.530 ;
        RECT 53.835 49.050 54.225 70.560 ;
        RECT 54.625 69.970 55.515 70.700 ;
        RECT 54.725 65.150 54.985 69.970 ;
        RECT 56.365 68.580 59.075 69.430 ;
        RECT 56.565 65.800 58.495 68.580 ;
        RECT 64.195 68.520 64.735 71.750 ;
        RECT 65.035 70.550 65.445 73.280 ;
        RECT 72.585 73.130 74.655 74.410 ;
        RECT 75.550 73.210 78.110 75.740 ;
        RECT 75.135 71.740 75.995 72.580 ;
        RECT 61.465 67.090 62.585 67.770 ;
        RECT 61.745 65.810 62.415 67.090 ;
        RECT 55.125 65.420 60.175 65.800 ;
        RECT 61.535 65.400 62.585 65.810 ;
        RECT 54.725 63.600 55.105 65.150 ;
        RECT 54.845 55.760 55.105 63.600 ;
        RECT 60.155 63.160 60.425 65.200 ;
        RECT 61.285 63.160 61.555 65.160 ;
        RECT 60.155 56.470 61.555 63.160 ;
        RECT 54.755 55.250 55.115 55.760 ;
        RECT 54.735 54.820 55.115 55.250 ;
        RECT 60.155 55.150 60.425 56.470 ;
        RECT 61.285 55.110 61.555 56.470 ;
        RECT 62.555 55.220 62.875 65.150 ;
        RECT 62.555 55.160 62.885 55.220 ;
        RECT 54.735 54.540 54.985 54.820 ;
        RECT 54.535 54.140 59.175 54.540 ;
        RECT 60.075 54.250 61.205 54.260 ;
        RECT 62.565 54.250 62.885 55.160 ;
        RECT 54.735 52.020 54.985 54.140 ;
        RECT 59.435 53.450 59.795 54.070 ;
        RECT 59.515 52.570 59.775 53.450 ;
        RECT 60.055 53.200 62.885 54.250 ;
        RECT 59.345 52.190 59.875 52.570 ;
        RECT 54.735 51.930 55.235 52.020 ;
        RECT 54.725 51.200 55.235 51.930 ;
        RECT 54.965 50.200 55.235 51.200 ;
        RECT 55.875 50.950 56.145 51.900 ;
        RECT 55.875 50.800 56.345 50.950 ;
        RECT 55.875 50.120 56.435 50.800 ;
        RECT 55.955 50.110 56.435 50.120 ;
        RECT 55.245 49.580 55.865 49.940 ;
        RECT 55.285 49.050 55.715 49.580 ;
        RECT 53.835 48.630 55.715 49.050 ;
        RECT 56.205 48.920 56.435 50.110 ;
        RECT 55.285 47.760 55.715 48.630 ;
        RECT 56.125 48.320 56.505 48.920 ;
        RECT 52.995 47.020 53.685 47.730 ;
        RECT 55.105 47.400 55.725 47.760 ;
        RECT 54.805 47.020 55.095 47.210 ;
        RECT 52.995 46.580 55.095 47.020 ;
        RECT 52.995 46.560 53.685 46.580 ;
        RECT 54.805 46.340 55.095 46.580 ;
        RECT 55.725 46.950 55.995 47.200 ;
        RECT 56.205 46.950 56.435 48.320 ;
        RECT 59.025 46.970 59.355 51.990 ;
        RECT 60.075 51.980 61.205 53.200 ;
        RECT 62.565 53.180 62.885 53.200 ;
        RECT 55.725 46.840 56.435 46.950 ;
        RECT 59.015 46.920 59.355 46.970 ;
        RECT 59.905 47.740 61.285 51.980 ;
        RECT 55.725 46.530 56.385 46.840 ;
        RECT 55.725 46.360 55.995 46.530 ;
        RECT 59.015 44.960 59.295 46.920 ;
        RECT 59.905 46.880 60.205 47.740 ;
        RECT 60.985 46.880 61.285 47.740 ;
        RECT 61.835 46.880 62.165 51.950 ;
        RECT 61.235 46.340 61.715 46.720 ;
        RECT 61.335 45.720 61.585 46.340 ;
        RECT 61.235 45.120 61.615 45.720 ;
        RECT 19.865 42.210 21.245 42.780 ;
        RECT 27.495 42.630 28.875 43.200 ;
        RECT 31.145 42.210 32.525 42.780 ;
        RECT 38.695 42.640 40.075 43.210 ;
        RECT 50.635 43.180 50.935 44.910 ;
        RECT 58.495 44.190 59.595 44.960 ;
        RECT 61.885 44.890 62.165 46.880 ;
        RECT 64.215 47.720 64.715 68.520 ;
        RECT 65.055 49.040 65.445 70.550 ;
        RECT 65.845 69.960 66.735 70.690 ;
        RECT 65.945 65.140 66.205 69.960 ;
        RECT 67.585 68.570 70.295 69.420 ;
        RECT 67.785 65.790 69.715 68.570 ;
        RECT 75.435 68.510 75.975 71.740 ;
        RECT 76.275 70.540 76.685 73.210 ;
        RECT 83.855 73.120 85.925 74.400 ;
        RECT 86.850 73.230 89.410 75.760 ;
        RECT 98.150 75.750 116.230 75.840 ;
        RECT 86.385 71.750 87.245 72.590 ;
        RECT 72.685 67.080 73.805 67.760 ;
        RECT 72.965 65.800 73.635 67.080 ;
        RECT 66.345 65.410 71.395 65.790 ;
        RECT 72.755 65.390 73.805 65.800 ;
        RECT 65.945 63.590 66.325 65.140 ;
        RECT 66.065 55.750 66.325 63.590 ;
        RECT 71.375 63.150 71.645 65.190 ;
        RECT 72.505 63.150 72.775 65.150 ;
        RECT 71.375 56.460 72.775 63.150 ;
        RECT 65.975 55.240 66.335 55.750 ;
        RECT 65.955 54.810 66.335 55.240 ;
        RECT 71.375 55.140 71.645 56.460 ;
        RECT 72.505 55.100 72.775 56.460 ;
        RECT 73.775 55.210 74.095 65.140 ;
        RECT 73.775 55.150 74.105 55.210 ;
        RECT 65.955 54.530 66.205 54.810 ;
        RECT 65.755 54.130 70.395 54.530 ;
        RECT 71.295 54.240 72.425 54.250 ;
        RECT 73.785 54.240 74.105 55.150 ;
        RECT 65.955 52.010 66.205 54.130 ;
        RECT 70.655 53.440 71.015 54.060 ;
        RECT 70.735 52.560 70.995 53.440 ;
        RECT 71.275 53.190 74.105 54.240 ;
        RECT 70.565 52.180 71.095 52.560 ;
        RECT 65.955 51.920 66.455 52.010 ;
        RECT 65.945 51.190 66.455 51.920 ;
        RECT 66.185 50.190 66.455 51.190 ;
        RECT 67.095 50.940 67.365 51.890 ;
        RECT 67.095 50.790 67.565 50.940 ;
        RECT 67.095 50.110 67.655 50.790 ;
        RECT 67.175 50.100 67.655 50.110 ;
        RECT 66.465 49.570 67.085 49.930 ;
        RECT 66.505 49.040 66.935 49.570 ;
        RECT 65.055 48.620 66.935 49.040 ;
        RECT 67.425 48.910 67.655 50.100 ;
        RECT 66.505 47.750 66.935 48.620 ;
        RECT 67.345 48.310 67.725 48.910 ;
        RECT 64.215 47.010 64.905 47.720 ;
        RECT 66.325 47.390 66.945 47.750 ;
        RECT 66.025 47.010 66.315 47.200 ;
        RECT 64.215 46.570 66.315 47.010 ;
        RECT 64.215 46.550 64.905 46.570 ;
        RECT 66.025 46.330 66.315 46.570 ;
        RECT 66.945 46.940 67.215 47.190 ;
        RECT 67.425 46.940 67.655 48.310 ;
        RECT 70.245 46.960 70.575 51.980 ;
        RECT 71.295 51.970 72.425 53.190 ;
        RECT 73.785 53.170 74.105 53.190 ;
        RECT 66.945 46.830 67.655 46.940 ;
        RECT 70.235 46.910 70.575 46.960 ;
        RECT 71.125 47.730 72.505 51.970 ;
        RECT 66.945 46.520 67.605 46.830 ;
        RECT 66.945 46.350 67.215 46.520 ;
        RECT 70.235 44.950 70.515 46.910 ;
        RECT 71.125 46.870 71.425 47.730 ;
        RECT 72.205 46.870 72.505 47.730 ;
        RECT 73.055 46.870 73.385 51.940 ;
        RECT 72.455 46.330 72.935 46.710 ;
        RECT 72.555 45.710 72.805 46.330 ;
        RECT 72.455 45.110 72.835 45.710 ;
        RECT 20.225 40.480 20.525 42.210 ;
        RECT 20.245 38.490 20.525 40.480 ;
        RECT 22.815 40.410 23.915 41.180 ;
        RECT 31.505 40.480 31.805 42.210 ;
        RECT 42.435 42.190 43.815 42.760 ;
        RECT 49.915 42.610 51.295 43.180 ;
        RECT 61.885 43.160 62.185 44.890 ;
        RECT 69.715 44.180 70.815 44.950 ;
        RECT 73.105 44.880 73.385 46.870 ;
        RECT 75.455 47.710 75.955 68.510 ;
        RECT 76.295 49.030 76.685 70.540 ;
        RECT 77.085 69.950 77.975 70.680 ;
        RECT 77.185 65.130 77.445 69.950 ;
        RECT 78.825 68.560 81.535 69.410 ;
        RECT 79.025 65.780 80.955 68.560 ;
        RECT 86.685 68.520 87.225 71.750 ;
        RECT 87.525 70.550 87.935 73.230 ;
        RECT 95.045 73.060 97.115 74.340 ;
        RECT 98.150 73.310 100.710 75.750 ;
        RECT 109.390 75.480 111.950 75.560 ;
        RECT 121.930 75.480 122.210 85.700 ;
        RECT 127.550 85.510 128.770 89.380 ;
        RECT 127.910 76.040 128.190 85.510 ;
        RECT 133.380 76.580 136.010 77.880 ;
        RECT 137.240 76.560 139.870 77.860 ;
        RECT 109.390 75.200 122.210 75.480 ;
        RECT 97.665 71.740 98.525 72.580 ;
        RECT 83.925 67.070 85.045 67.750 ;
        RECT 84.205 65.790 84.875 67.070 ;
        RECT 77.585 65.400 82.635 65.780 ;
        RECT 83.995 65.380 85.045 65.790 ;
        RECT 77.185 63.580 77.565 65.130 ;
        RECT 77.305 55.740 77.565 63.580 ;
        RECT 82.615 63.140 82.885 65.180 ;
        RECT 83.745 63.140 84.015 65.140 ;
        RECT 82.615 56.450 84.015 63.140 ;
        RECT 77.215 55.230 77.575 55.740 ;
        RECT 77.195 54.800 77.575 55.230 ;
        RECT 82.615 55.130 82.885 56.450 ;
        RECT 83.745 55.090 84.015 56.450 ;
        RECT 85.015 55.200 85.335 65.130 ;
        RECT 85.015 55.140 85.345 55.200 ;
        RECT 77.195 54.520 77.445 54.800 ;
        RECT 76.995 54.120 81.635 54.520 ;
        RECT 82.535 54.230 83.665 54.240 ;
        RECT 85.025 54.230 85.345 55.140 ;
        RECT 77.195 52.000 77.445 54.120 ;
        RECT 81.895 53.430 82.255 54.050 ;
        RECT 81.975 52.550 82.235 53.430 ;
        RECT 82.515 53.180 85.345 54.230 ;
        RECT 81.805 52.170 82.335 52.550 ;
        RECT 77.195 51.910 77.695 52.000 ;
        RECT 77.185 51.180 77.695 51.910 ;
        RECT 77.425 50.180 77.695 51.180 ;
        RECT 78.335 50.930 78.605 51.880 ;
        RECT 78.335 50.780 78.805 50.930 ;
        RECT 78.335 50.100 78.895 50.780 ;
        RECT 78.415 50.090 78.895 50.100 ;
        RECT 77.705 49.560 78.325 49.920 ;
        RECT 77.745 49.030 78.175 49.560 ;
        RECT 76.295 48.610 78.175 49.030 ;
        RECT 78.665 48.900 78.895 50.090 ;
        RECT 77.745 47.740 78.175 48.610 ;
        RECT 78.585 48.300 78.965 48.900 ;
        RECT 75.455 47.000 76.145 47.710 ;
        RECT 77.565 47.380 78.185 47.740 ;
        RECT 77.265 47.000 77.555 47.190 ;
        RECT 75.455 46.560 77.555 47.000 ;
        RECT 75.455 46.540 76.145 46.560 ;
        RECT 77.265 46.320 77.555 46.560 ;
        RECT 78.185 46.930 78.455 47.180 ;
        RECT 78.665 46.930 78.895 48.300 ;
        RECT 81.485 46.950 81.815 51.970 ;
        RECT 82.535 51.960 83.665 53.180 ;
        RECT 85.025 53.160 85.345 53.180 ;
        RECT 78.185 46.820 78.895 46.930 ;
        RECT 81.475 46.900 81.815 46.950 ;
        RECT 82.365 47.720 83.745 51.960 ;
        RECT 78.185 46.510 78.845 46.820 ;
        RECT 78.185 46.340 78.455 46.510 ;
        RECT 81.475 44.940 81.755 46.900 ;
        RECT 82.365 46.860 82.665 47.720 ;
        RECT 83.445 46.860 83.745 47.720 ;
        RECT 84.295 46.860 84.625 51.930 ;
        RECT 83.695 46.320 84.175 46.700 ;
        RECT 83.795 45.700 84.045 46.320 ;
        RECT 83.695 45.100 84.075 45.700 ;
        RECT 53.655 42.190 55.035 42.760 ;
        RECT 61.165 42.590 62.545 43.160 ;
        RECT 73.105 43.150 73.405 44.880 ;
        RECT 80.955 44.170 82.055 44.940 ;
        RECT 84.345 44.870 84.625 46.860 ;
        RECT 86.705 47.720 87.205 68.520 ;
        RECT 87.545 49.040 87.935 70.550 ;
        RECT 88.335 69.960 89.225 70.690 ;
        RECT 88.435 65.140 88.695 69.960 ;
        RECT 90.075 68.570 92.785 69.420 ;
        RECT 90.275 65.790 92.205 68.570 ;
        RECT 97.965 68.510 98.505 71.740 ;
        RECT 98.805 70.540 99.215 73.310 ;
        RECT 106.455 73.110 108.525 74.390 ;
        RECT 109.390 73.030 111.950 75.200 ;
        RECT 125.760 74.810 128.190 76.040 ;
        RECT 121.290 74.790 128.190 74.810 ;
        RECT 120.600 74.530 128.190 74.790 ;
        RECT 117.655 73.110 119.725 74.390 ;
        RECT 120.600 73.180 128.160 74.530 ;
        RECT 129.505 73.190 131.575 74.470 ;
        RECT 120.600 73.110 126.160 73.180 ;
        RECT 108.935 71.740 109.795 72.580 ;
        RECT 95.175 67.080 96.295 67.760 ;
        RECT 95.455 65.800 96.125 67.080 ;
        RECT 88.835 65.410 93.885 65.790 ;
        RECT 95.245 65.390 96.295 65.800 ;
        RECT 88.435 63.590 88.815 65.140 ;
        RECT 88.555 55.750 88.815 63.590 ;
        RECT 93.865 63.150 94.135 65.190 ;
        RECT 94.995 63.150 95.265 65.150 ;
        RECT 93.865 56.460 95.265 63.150 ;
        RECT 88.465 55.240 88.825 55.750 ;
        RECT 88.445 54.810 88.825 55.240 ;
        RECT 93.865 55.140 94.135 56.460 ;
        RECT 94.995 55.100 95.265 56.460 ;
        RECT 96.265 55.210 96.585 65.140 ;
        RECT 96.265 55.150 96.595 55.210 ;
        RECT 88.445 54.530 88.695 54.810 ;
        RECT 88.245 54.130 92.885 54.530 ;
        RECT 93.785 54.240 94.915 54.250 ;
        RECT 96.275 54.240 96.595 55.150 ;
        RECT 88.445 52.010 88.695 54.130 ;
        RECT 93.145 53.440 93.505 54.060 ;
        RECT 93.225 52.560 93.485 53.440 ;
        RECT 93.765 53.190 96.595 54.240 ;
        RECT 93.055 52.180 93.585 52.560 ;
        RECT 88.445 51.920 88.945 52.010 ;
        RECT 88.435 51.190 88.945 51.920 ;
        RECT 88.675 50.190 88.945 51.190 ;
        RECT 89.585 50.940 89.855 51.890 ;
        RECT 89.585 50.790 90.055 50.940 ;
        RECT 89.585 50.110 90.145 50.790 ;
        RECT 89.665 50.100 90.145 50.110 ;
        RECT 88.955 49.570 89.575 49.930 ;
        RECT 88.995 49.040 89.425 49.570 ;
        RECT 87.545 48.620 89.425 49.040 ;
        RECT 89.915 48.910 90.145 50.100 ;
        RECT 88.995 47.750 89.425 48.620 ;
        RECT 89.835 48.310 90.215 48.910 ;
        RECT 86.705 47.010 87.395 47.720 ;
        RECT 88.815 47.390 89.435 47.750 ;
        RECT 88.515 47.010 88.805 47.200 ;
        RECT 86.705 46.570 88.805 47.010 ;
        RECT 86.705 46.550 87.395 46.570 ;
        RECT 88.515 46.330 88.805 46.570 ;
        RECT 89.435 46.940 89.705 47.190 ;
        RECT 89.915 46.940 90.145 48.310 ;
        RECT 92.735 46.960 93.065 51.980 ;
        RECT 93.785 51.970 94.915 53.190 ;
        RECT 96.275 53.170 96.595 53.190 ;
        RECT 89.435 46.830 90.145 46.940 ;
        RECT 92.725 46.910 93.065 46.960 ;
        RECT 93.615 47.730 94.995 51.970 ;
        RECT 89.435 46.520 90.095 46.830 ;
        RECT 89.435 46.350 89.705 46.520 ;
        RECT 92.725 44.950 93.005 46.910 ;
        RECT 93.615 46.870 93.915 47.730 ;
        RECT 94.695 46.870 94.995 47.730 ;
        RECT 95.545 46.870 95.875 51.940 ;
        RECT 94.945 46.330 95.425 46.710 ;
        RECT 95.045 45.710 95.295 46.330 ;
        RECT 94.945 45.110 95.325 45.710 ;
        RECT 64.855 42.190 66.235 42.760 ;
        RECT 72.385 42.580 73.765 43.150 ;
        RECT 84.345 43.140 84.645 44.870 ;
        RECT 92.205 44.180 93.305 44.950 ;
        RECT 95.595 44.880 95.875 46.870 ;
        RECT 97.985 47.710 98.485 68.510 ;
        RECT 98.825 49.030 99.215 70.540 ;
        RECT 99.615 69.950 100.505 70.680 ;
        RECT 99.715 65.130 99.975 69.950 ;
        RECT 101.355 68.560 104.065 69.410 ;
        RECT 101.555 65.780 103.485 68.560 ;
        RECT 109.235 68.510 109.775 71.740 ;
        RECT 110.075 70.540 110.485 73.030 ;
        RECT 120.185 71.740 121.045 72.580 ;
        RECT 106.455 67.070 107.575 67.750 ;
        RECT 106.735 65.790 107.405 67.070 ;
        RECT 100.115 65.400 105.165 65.780 ;
        RECT 106.525 65.380 107.575 65.790 ;
        RECT 99.715 63.580 100.095 65.130 ;
        RECT 99.835 55.740 100.095 63.580 ;
        RECT 105.145 63.140 105.415 65.180 ;
        RECT 106.275 63.140 106.545 65.140 ;
        RECT 105.145 56.450 106.545 63.140 ;
        RECT 99.745 55.230 100.105 55.740 ;
        RECT 99.725 54.800 100.105 55.230 ;
        RECT 105.145 55.130 105.415 56.450 ;
        RECT 106.275 55.090 106.545 56.450 ;
        RECT 107.545 55.200 107.865 65.130 ;
        RECT 107.545 55.140 107.875 55.200 ;
        RECT 99.725 54.520 99.975 54.800 ;
        RECT 99.525 54.120 104.165 54.520 ;
        RECT 105.065 54.230 106.195 54.240 ;
        RECT 107.555 54.230 107.875 55.140 ;
        RECT 99.725 52.000 99.975 54.120 ;
        RECT 104.425 53.430 104.785 54.050 ;
        RECT 104.505 52.550 104.765 53.430 ;
        RECT 105.045 53.180 107.875 54.230 ;
        RECT 104.335 52.170 104.865 52.550 ;
        RECT 99.725 51.910 100.225 52.000 ;
        RECT 99.715 51.180 100.225 51.910 ;
        RECT 99.955 50.180 100.225 51.180 ;
        RECT 100.865 50.930 101.135 51.880 ;
        RECT 100.865 50.780 101.335 50.930 ;
        RECT 100.865 50.100 101.425 50.780 ;
        RECT 100.945 50.090 101.425 50.100 ;
        RECT 100.235 49.560 100.855 49.920 ;
        RECT 100.275 49.030 100.705 49.560 ;
        RECT 98.825 48.610 100.705 49.030 ;
        RECT 101.195 48.900 101.425 50.090 ;
        RECT 100.275 47.740 100.705 48.610 ;
        RECT 101.115 48.300 101.495 48.900 ;
        RECT 97.985 47.000 98.675 47.710 ;
        RECT 100.095 47.380 100.715 47.740 ;
        RECT 99.795 47.000 100.085 47.190 ;
        RECT 97.985 46.560 100.085 47.000 ;
        RECT 97.985 46.540 98.675 46.560 ;
        RECT 99.795 46.320 100.085 46.560 ;
        RECT 100.715 46.930 100.985 47.180 ;
        RECT 101.195 46.930 101.425 48.300 ;
        RECT 104.015 46.950 104.345 51.970 ;
        RECT 105.065 51.960 106.195 53.180 ;
        RECT 107.555 53.160 107.875 53.180 ;
        RECT 100.715 46.820 101.425 46.930 ;
        RECT 104.005 46.900 104.345 46.950 ;
        RECT 104.895 47.720 106.275 51.960 ;
        RECT 100.715 46.510 101.375 46.820 ;
        RECT 100.715 46.340 100.985 46.510 ;
        RECT 104.005 44.940 104.285 46.900 ;
        RECT 104.895 46.860 105.195 47.720 ;
        RECT 105.975 46.860 106.275 47.720 ;
        RECT 106.825 46.860 107.155 51.930 ;
        RECT 106.225 46.320 106.705 46.700 ;
        RECT 106.325 45.700 106.575 46.320 ;
        RECT 106.225 45.100 106.605 45.700 ;
        RECT 95.595 43.150 95.895 44.880 ;
        RECT 103.485 44.170 104.585 44.940 ;
        RECT 106.875 44.870 107.155 46.860 ;
        RECT 109.255 47.710 109.755 68.510 ;
        RECT 110.095 49.030 110.485 70.540 ;
        RECT 110.885 69.950 111.775 70.680 ;
        RECT 110.985 65.130 111.245 69.950 ;
        RECT 112.625 68.560 115.335 69.410 ;
        RECT 112.825 65.780 114.755 68.560 ;
        RECT 120.485 68.510 121.025 71.740 ;
        RECT 121.325 70.540 121.735 73.110 ;
        RECT 132.925 70.810 133.225 70.900 ;
        RECT 117.725 67.070 118.845 67.750 ;
        RECT 118.005 65.790 118.675 67.070 ;
        RECT 111.385 65.400 116.435 65.780 ;
        RECT 117.795 65.380 118.845 65.790 ;
        RECT 110.985 63.580 111.365 65.130 ;
        RECT 111.105 55.740 111.365 63.580 ;
        RECT 116.415 63.140 116.685 65.180 ;
        RECT 117.545 63.140 117.815 65.140 ;
        RECT 116.415 56.450 117.815 63.140 ;
        RECT 111.015 55.230 111.375 55.740 ;
        RECT 110.995 54.800 111.375 55.230 ;
        RECT 116.415 55.130 116.685 56.450 ;
        RECT 117.545 55.090 117.815 56.450 ;
        RECT 118.815 55.200 119.135 65.130 ;
        RECT 118.815 55.140 119.145 55.200 ;
        RECT 110.995 54.520 111.245 54.800 ;
        RECT 110.795 54.120 115.435 54.520 ;
        RECT 116.335 54.230 117.465 54.240 ;
        RECT 118.825 54.230 119.145 55.140 ;
        RECT 110.995 52.000 111.245 54.120 ;
        RECT 115.695 53.430 116.055 54.050 ;
        RECT 115.775 52.550 116.035 53.430 ;
        RECT 116.315 53.180 119.145 54.230 ;
        RECT 115.605 52.170 116.135 52.550 ;
        RECT 110.995 51.910 111.495 52.000 ;
        RECT 110.985 51.180 111.495 51.910 ;
        RECT 111.225 50.180 111.495 51.180 ;
        RECT 112.135 50.930 112.405 51.880 ;
        RECT 112.135 50.780 112.605 50.930 ;
        RECT 112.135 50.100 112.695 50.780 ;
        RECT 112.215 50.090 112.695 50.100 ;
        RECT 111.505 49.560 112.125 49.920 ;
        RECT 111.545 49.030 111.975 49.560 ;
        RECT 110.095 48.610 111.975 49.030 ;
        RECT 112.465 48.900 112.695 50.090 ;
        RECT 111.545 47.740 111.975 48.610 ;
        RECT 112.385 48.300 112.765 48.900 ;
        RECT 109.255 47.000 109.945 47.710 ;
        RECT 111.365 47.380 111.985 47.740 ;
        RECT 111.065 47.000 111.355 47.190 ;
        RECT 109.255 46.560 111.355 47.000 ;
        RECT 109.255 46.540 109.945 46.560 ;
        RECT 111.065 46.320 111.355 46.560 ;
        RECT 111.985 46.930 112.255 47.180 ;
        RECT 112.465 46.930 112.695 48.300 ;
        RECT 115.285 46.950 115.615 51.970 ;
        RECT 116.335 51.960 117.465 53.180 ;
        RECT 118.825 53.160 119.145 53.180 ;
        RECT 111.985 46.820 112.695 46.930 ;
        RECT 115.275 46.900 115.615 46.950 ;
        RECT 116.165 47.720 117.545 51.960 ;
        RECT 111.985 46.510 112.645 46.820 ;
        RECT 111.985 46.340 112.255 46.510 ;
        RECT 115.275 44.940 115.555 46.900 ;
        RECT 116.165 46.860 116.465 47.720 ;
        RECT 117.245 46.860 117.545 47.720 ;
        RECT 118.095 46.860 118.425 51.930 ;
        RECT 117.495 46.320 117.975 46.700 ;
        RECT 117.595 45.700 117.845 46.320 ;
        RECT 117.495 45.100 117.875 45.700 ;
        RECT 20.795 39.650 21.175 40.250 ;
        RECT 20.825 39.030 21.075 39.650 ;
        RECT 20.695 38.650 21.175 39.030 ;
        RECT 20.245 33.420 20.575 38.490 ;
        RECT 21.125 37.630 21.425 38.490 ;
        RECT 22.205 37.630 22.505 38.490 ;
        RECT 23.115 38.450 23.395 40.410 ;
        RECT 26.415 38.840 26.685 39.010 ;
        RECT 26.025 38.530 26.685 38.840 ;
        RECT 21.125 33.390 22.505 37.630 ;
        RECT 23.055 38.400 23.395 38.450 ;
        RECT 25.975 38.420 26.685 38.530 ;
        RECT 19.525 32.170 19.845 32.190 ;
        RECT 21.205 32.170 22.335 33.390 ;
        RECT 23.055 33.380 23.385 38.400 ;
        RECT 25.975 37.050 26.205 38.420 ;
        RECT 26.415 38.170 26.685 38.420 ;
        RECT 27.315 38.790 27.605 39.030 ;
        RECT 28.725 38.790 29.415 38.810 ;
        RECT 27.315 38.350 29.415 38.790 ;
        RECT 27.315 38.160 27.605 38.350 ;
        RECT 26.685 37.610 27.305 37.970 ;
        RECT 28.725 37.640 29.415 38.350 ;
        RECT 25.905 36.450 26.285 37.050 ;
        RECT 26.695 36.740 27.125 37.610 ;
        RECT 25.975 35.260 26.205 36.450 ;
        RECT 26.695 36.320 28.575 36.740 ;
        RECT 26.695 35.790 27.125 36.320 ;
        RECT 26.545 35.430 27.165 35.790 ;
        RECT 25.975 35.250 26.455 35.260 ;
        RECT 25.975 34.570 26.535 35.250 ;
        RECT 26.065 34.420 26.535 34.570 ;
        RECT 26.265 33.470 26.535 34.420 ;
        RECT 27.175 34.170 27.445 35.170 ;
        RECT 27.175 33.440 27.685 34.170 ;
        RECT 27.175 33.350 27.675 33.440 ;
        RECT 22.535 32.800 23.065 33.180 ;
        RECT 19.525 31.120 22.355 32.170 ;
        RECT 22.635 31.920 22.895 32.800 ;
        RECT 22.615 31.300 22.975 31.920 ;
        RECT 27.425 31.230 27.675 33.350 ;
        RECT 19.525 30.210 19.845 31.120 ;
        RECT 21.205 31.110 22.335 31.120 ;
        RECT 23.235 30.830 27.875 31.230 ;
        RECT 27.425 30.550 27.675 30.830 ;
        RECT 19.525 30.150 19.855 30.210 ;
        RECT 19.535 20.220 19.855 30.150 ;
        RECT 20.855 28.900 21.125 30.260 ;
        RECT 21.985 28.900 22.255 30.220 ;
        RECT 27.295 30.120 27.675 30.550 ;
        RECT 27.295 29.610 27.655 30.120 ;
        RECT 20.855 22.210 22.255 28.900 ;
        RECT 20.855 20.210 21.125 22.210 ;
        RECT 21.985 20.170 22.255 22.210 ;
        RECT 27.305 21.770 27.565 29.610 ;
        RECT 27.305 20.220 27.685 21.770 ;
        RECT 19.825 19.560 20.875 19.970 ;
        RECT 22.235 19.570 27.285 19.950 ;
        RECT 19.995 18.280 20.665 19.560 ;
        RECT 19.825 17.600 20.945 18.280 ;
        RECT 23.915 16.790 25.845 19.570 ;
        RECT 23.335 15.940 26.045 16.790 ;
        RECT 27.425 15.400 27.685 20.220 ;
        RECT 26.895 14.670 27.785 15.400 ;
        RECT 28.185 14.810 28.575 36.320 ;
        RECT 28.915 16.840 29.415 37.640 ;
        RECT 31.525 38.490 31.805 40.480 ;
        RECT 34.095 40.410 35.195 41.180 ;
        RECT 42.795 40.460 43.095 42.190 ;
        RECT 32.075 39.650 32.455 40.250 ;
        RECT 32.105 39.030 32.355 39.650 ;
        RECT 31.975 38.650 32.455 39.030 ;
        RECT 31.525 33.420 31.855 38.490 ;
        RECT 32.405 37.630 32.705 38.490 ;
        RECT 33.485 37.630 33.785 38.490 ;
        RECT 34.395 38.450 34.675 40.410 ;
        RECT 37.695 38.840 37.965 39.010 ;
        RECT 37.305 38.530 37.965 38.840 ;
        RECT 32.405 33.390 33.785 37.630 ;
        RECT 34.335 38.400 34.675 38.450 ;
        RECT 37.255 38.420 37.965 38.530 ;
        RECT 30.805 32.170 31.125 32.190 ;
        RECT 32.485 32.170 33.615 33.390 ;
        RECT 34.335 33.380 34.665 38.400 ;
        RECT 37.255 37.050 37.485 38.420 ;
        RECT 37.695 38.170 37.965 38.420 ;
        RECT 38.595 38.790 38.885 39.030 ;
        RECT 40.005 38.790 40.695 38.810 ;
        RECT 38.595 38.350 40.695 38.790 ;
        RECT 38.595 38.160 38.885 38.350 ;
        RECT 37.965 37.610 38.585 37.970 ;
        RECT 40.005 37.640 40.695 38.350 ;
        RECT 37.185 36.450 37.565 37.050 ;
        RECT 37.975 36.740 38.405 37.610 ;
        RECT 37.255 35.260 37.485 36.450 ;
        RECT 37.975 36.320 39.855 36.740 ;
        RECT 37.975 35.790 38.405 36.320 ;
        RECT 37.825 35.430 38.445 35.790 ;
        RECT 37.255 35.250 37.735 35.260 ;
        RECT 37.255 34.570 37.815 35.250 ;
        RECT 37.345 34.420 37.815 34.570 ;
        RECT 37.545 33.470 37.815 34.420 ;
        RECT 38.455 34.170 38.725 35.170 ;
        RECT 38.455 33.440 38.965 34.170 ;
        RECT 38.455 33.350 38.955 33.440 ;
        RECT 33.815 32.800 34.345 33.180 ;
        RECT 30.805 31.120 33.635 32.170 ;
        RECT 33.915 31.920 34.175 32.800 ;
        RECT 33.895 31.300 34.255 31.920 ;
        RECT 38.705 31.230 38.955 33.350 ;
        RECT 30.805 30.210 31.125 31.120 ;
        RECT 32.485 31.110 33.615 31.120 ;
        RECT 34.515 30.830 39.155 31.230 ;
        RECT 38.705 30.550 38.955 30.830 ;
        RECT 30.805 30.150 31.135 30.210 ;
        RECT 30.815 20.220 31.135 30.150 ;
        RECT 32.135 28.900 32.405 30.260 ;
        RECT 33.265 28.900 33.535 30.220 ;
        RECT 38.575 30.120 38.955 30.550 ;
        RECT 38.575 29.610 38.935 30.120 ;
        RECT 32.135 22.210 33.535 28.900 ;
        RECT 32.135 20.210 32.405 22.210 ;
        RECT 33.265 20.170 33.535 22.210 ;
        RECT 38.585 21.770 38.845 29.610 ;
        RECT 38.585 20.220 38.965 21.770 ;
        RECT 31.105 19.560 32.155 19.970 ;
        RECT 33.515 19.570 38.565 19.950 ;
        RECT 31.275 18.280 31.945 19.560 ;
        RECT 31.105 17.600 32.225 18.280 ;
        RECT 28.185 12.290 28.595 14.810 ;
        RECT 28.895 13.610 29.435 16.840 ;
        RECT 35.195 16.790 37.125 19.570 ;
        RECT 34.615 15.940 37.325 16.790 ;
        RECT 38.705 15.400 38.965 20.220 ;
        RECT 38.175 14.670 39.065 15.400 ;
        RECT 39.465 14.810 39.855 36.320 ;
        RECT 40.195 16.840 40.695 37.640 ;
        RECT 42.815 38.470 43.095 40.460 ;
        RECT 45.385 40.390 46.485 41.160 ;
        RECT 54.015 40.460 54.315 42.190 ;
        RECT 43.365 39.630 43.745 40.230 ;
        RECT 43.395 39.010 43.645 39.630 ;
        RECT 43.265 38.630 43.745 39.010 ;
        RECT 42.815 33.400 43.145 38.470 ;
        RECT 43.695 37.610 43.995 38.470 ;
        RECT 44.775 37.610 45.075 38.470 ;
        RECT 45.685 38.430 45.965 40.390 ;
        RECT 48.985 38.820 49.255 38.990 ;
        RECT 48.595 38.510 49.255 38.820 ;
        RECT 43.695 33.370 45.075 37.610 ;
        RECT 45.625 38.380 45.965 38.430 ;
        RECT 48.545 38.400 49.255 38.510 ;
        RECT 42.095 32.150 42.415 32.170 ;
        RECT 43.775 32.150 44.905 33.370 ;
        RECT 45.625 33.360 45.955 38.380 ;
        RECT 48.545 37.030 48.775 38.400 ;
        RECT 48.985 38.150 49.255 38.400 ;
        RECT 49.885 38.770 50.175 39.010 ;
        RECT 51.295 38.770 51.985 38.790 ;
        RECT 49.885 38.330 51.985 38.770 ;
        RECT 49.885 38.140 50.175 38.330 ;
        RECT 49.255 37.590 49.875 37.950 ;
        RECT 51.295 37.620 51.985 38.330 ;
        RECT 48.475 36.430 48.855 37.030 ;
        RECT 49.265 36.720 49.695 37.590 ;
        RECT 48.545 35.240 48.775 36.430 ;
        RECT 49.265 36.300 51.145 36.720 ;
        RECT 49.265 35.770 49.695 36.300 ;
        RECT 49.115 35.410 49.735 35.770 ;
        RECT 48.545 35.230 49.025 35.240 ;
        RECT 48.545 34.550 49.105 35.230 ;
        RECT 48.635 34.400 49.105 34.550 ;
        RECT 48.835 33.450 49.105 34.400 ;
        RECT 49.745 34.150 50.015 35.150 ;
        RECT 49.745 33.420 50.255 34.150 ;
        RECT 49.745 33.330 50.245 33.420 ;
        RECT 45.105 32.780 45.635 33.160 ;
        RECT 42.095 31.100 44.925 32.150 ;
        RECT 45.205 31.900 45.465 32.780 ;
        RECT 45.185 31.280 45.545 31.900 ;
        RECT 49.995 31.210 50.245 33.330 ;
        RECT 42.095 30.190 42.415 31.100 ;
        RECT 43.775 31.090 44.905 31.100 ;
        RECT 45.805 30.810 50.445 31.210 ;
        RECT 49.995 30.530 50.245 30.810 ;
        RECT 42.095 30.130 42.425 30.190 ;
        RECT 42.105 20.200 42.425 30.130 ;
        RECT 43.425 28.880 43.695 30.240 ;
        RECT 44.555 28.880 44.825 30.200 ;
        RECT 49.865 30.100 50.245 30.530 ;
        RECT 49.865 29.590 50.225 30.100 ;
        RECT 43.425 22.190 44.825 28.880 ;
        RECT 43.425 20.190 43.695 22.190 ;
        RECT 44.555 20.150 44.825 22.190 ;
        RECT 49.875 21.750 50.135 29.590 ;
        RECT 49.875 20.200 50.255 21.750 ;
        RECT 42.395 19.540 43.445 19.950 ;
        RECT 44.805 19.550 49.855 19.930 ;
        RECT 42.565 18.260 43.235 19.540 ;
        RECT 42.395 17.580 43.515 18.260 ;
        RECT 28.875 12.770 29.735 13.610 ;
        RECT 28.185 11.950 30.415 12.290 ;
        RECT 39.465 11.990 39.875 14.810 ;
        RECT 40.175 13.610 40.715 16.840 ;
        RECT 46.485 16.770 48.415 19.550 ;
        RECT 45.905 15.920 48.615 16.770 ;
        RECT 49.995 15.380 50.255 20.200 ;
        RECT 49.465 14.650 50.355 15.380 ;
        RECT 50.755 14.790 51.145 36.300 ;
        RECT 51.485 16.820 51.985 37.620 ;
        RECT 54.035 38.470 54.315 40.460 ;
        RECT 56.605 40.390 57.705 41.160 ;
        RECT 65.215 40.460 65.515 42.190 ;
        RECT 76.145 42.180 77.525 42.750 ;
        RECT 83.625 42.570 85.005 43.140 ;
        RECT 87.385 42.200 88.765 42.770 ;
        RECT 94.875 42.580 96.255 43.150 ;
        RECT 106.875 43.140 107.175 44.870 ;
        RECT 114.755 44.170 115.855 44.940 ;
        RECT 118.145 44.870 118.425 46.860 ;
        RECT 120.505 47.710 121.005 68.510 ;
        RECT 121.345 49.030 121.735 70.540 ;
        RECT 122.135 69.950 123.025 70.680 ;
        RECT 132.615 70.040 134.265 70.810 ;
        RECT 122.235 65.130 122.495 69.950 ;
        RECT 123.875 68.560 126.585 69.410 ;
        RECT 124.075 65.780 126.005 68.560 ;
        RECT 128.975 67.070 130.095 67.750 ;
        RECT 129.255 65.790 129.925 67.070 ;
        RECT 122.635 65.400 127.685 65.780 ;
        RECT 129.045 65.380 130.095 65.790 ;
        RECT 132.925 65.180 133.225 70.040 ;
        RECT 137.675 68.690 139.075 69.460 ;
        RECT 138.385 65.740 138.645 68.690 ;
        RECT 149.410 68.420 150.690 69.620 ;
        RECT 149.480 65.810 150.640 68.420 ;
        RECT 133.365 65.380 138.645 65.740 ;
        RECT 122.235 63.580 122.615 65.130 ;
        RECT 122.355 55.740 122.615 63.580 ;
        RECT 127.665 63.140 127.935 65.180 ;
        RECT 128.795 63.140 129.065 65.140 ;
        RECT 127.665 56.450 129.065 63.140 ;
        RECT 122.265 55.230 122.625 55.740 ;
        RECT 122.245 54.800 122.625 55.230 ;
        RECT 127.665 55.130 127.935 56.450 ;
        RECT 128.795 55.090 129.065 56.450 ;
        RECT 130.065 55.200 130.385 65.130 ;
        RECT 132.925 61.010 133.355 65.180 ;
        RECT 138.385 65.150 138.645 65.380 ;
        RECT 138.385 64.770 138.675 65.150 ;
        RECT 130.065 55.140 130.395 55.200 ;
        RECT 133.055 55.190 133.355 61.010 ;
        RECT 122.245 54.520 122.495 54.800 ;
        RECT 122.045 54.120 126.685 54.520 ;
        RECT 127.585 54.230 128.715 54.240 ;
        RECT 130.075 54.230 130.395 55.140 ;
        RECT 138.395 55.080 138.675 64.770 ;
        RECT 149.390 64.610 150.670 65.810 ;
        RECT 122.245 52.000 122.495 54.120 ;
        RECT 126.945 53.430 127.305 54.050 ;
        RECT 127.025 52.550 127.285 53.430 ;
        RECT 127.565 53.180 130.395 54.230 ;
        RECT 126.855 52.170 127.385 52.550 ;
        RECT 122.245 51.910 122.745 52.000 ;
        RECT 122.235 51.180 122.745 51.910 ;
        RECT 122.475 50.180 122.745 51.180 ;
        RECT 123.385 50.930 123.655 51.880 ;
        RECT 123.385 50.780 123.855 50.930 ;
        RECT 123.385 50.100 123.945 50.780 ;
        RECT 123.465 50.090 123.945 50.100 ;
        RECT 122.755 49.560 123.375 49.920 ;
        RECT 122.795 49.030 123.225 49.560 ;
        RECT 121.345 48.610 123.225 49.030 ;
        RECT 123.715 48.900 123.945 50.090 ;
        RECT 122.795 47.740 123.225 48.610 ;
        RECT 123.635 48.300 124.015 48.900 ;
        RECT 120.505 47.000 121.195 47.710 ;
        RECT 122.615 47.380 123.235 47.740 ;
        RECT 122.315 47.000 122.605 47.190 ;
        RECT 120.505 46.560 122.605 47.000 ;
        RECT 120.505 46.540 121.195 46.560 ;
        RECT 122.315 46.320 122.605 46.560 ;
        RECT 123.235 46.930 123.505 47.180 ;
        RECT 123.715 46.930 123.945 48.300 ;
        RECT 126.535 46.950 126.865 51.970 ;
        RECT 127.585 51.960 128.715 53.180 ;
        RECT 130.075 53.160 130.395 53.180 ;
        RECT 123.235 46.820 123.945 46.930 ;
        RECT 126.525 46.900 126.865 46.950 ;
        RECT 127.415 47.720 128.795 51.960 ;
        RECT 123.235 46.510 123.895 46.820 ;
        RECT 123.235 46.340 123.505 46.510 ;
        RECT 126.525 44.940 126.805 46.900 ;
        RECT 127.415 46.860 127.715 47.720 ;
        RECT 128.495 46.860 128.795 47.720 ;
        RECT 129.345 46.860 129.675 51.930 ;
        RECT 128.745 46.320 129.225 46.700 ;
        RECT 128.845 45.700 129.095 46.320 ;
        RECT 128.745 45.100 129.125 45.700 ;
        RECT 118.145 43.140 118.445 44.870 ;
        RECT 126.005 44.170 127.105 44.940 ;
        RECT 129.395 44.870 129.675 46.860 ;
        RECT 129.395 43.140 129.695 44.870 ;
        RECT 98.595 42.220 99.975 42.790 ;
        RECT 106.155 42.570 107.535 43.140 ;
        RECT 109.795 42.260 111.175 42.830 ;
        RECT 117.425 42.570 118.805 43.140 ;
        RECT 121.005 42.280 122.385 42.850 ;
        RECT 128.675 42.570 130.055 43.140 ;
        RECT 54.585 39.630 54.965 40.230 ;
        RECT 54.615 39.010 54.865 39.630 ;
        RECT 54.485 38.630 54.965 39.010 ;
        RECT 54.035 33.400 54.365 38.470 ;
        RECT 54.915 37.610 55.215 38.470 ;
        RECT 55.995 37.610 56.295 38.470 ;
        RECT 56.905 38.430 57.185 40.390 ;
        RECT 60.205 38.820 60.475 38.990 ;
        RECT 59.815 38.510 60.475 38.820 ;
        RECT 54.915 33.370 56.295 37.610 ;
        RECT 56.845 38.380 57.185 38.430 ;
        RECT 59.765 38.400 60.475 38.510 ;
        RECT 53.315 32.150 53.635 32.170 ;
        RECT 54.995 32.150 56.125 33.370 ;
        RECT 56.845 33.360 57.175 38.380 ;
        RECT 59.765 37.030 59.995 38.400 ;
        RECT 60.205 38.150 60.475 38.400 ;
        RECT 61.105 38.770 61.395 39.010 ;
        RECT 62.515 38.770 63.205 38.790 ;
        RECT 61.105 38.330 63.205 38.770 ;
        RECT 61.105 38.140 61.395 38.330 ;
        RECT 60.475 37.590 61.095 37.950 ;
        RECT 62.515 37.620 63.205 38.330 ;
        RECT 59.695 36.430 60.075 37.030 ;
        RECT 60.485 36.720 60.915 37.590 ;
        RECT 59.765 35.240 59.995 36.430 ;
        RECT 60.485 36.300 62.365 36.720 ;
        RECT 60.485 35.770 60.915 36.300 ;
        RECT 60.335 35.410 60.955 35.770 ;
        RECT 59.765 35.230 60.245 35.240 ;
        RECT 59.765 34.550 60.325 35.230 ;
        RECT 59.855 34.400 60.325 34.550 ;
        RECT 60.055 33.450 60.325 34.400 ;
        RECT 60.965 34.150 61.235 35.150 ;
        RECT 60.965 33.420 61.475 34.150 ;
        RECT 60.965 33.330 61.465 33.420 ;
        RECT 56.325 32.780 56.855 33.160 ;
        RECT 53.315 31.100 56.145 32.150 ;
        RECT 56.425 31.900 56.685 32.780 ;
        RECT 56.405 31.280 56.765 31.900 ;
        RECT 61.215 31.210 61.465 33.330 ;
        RECT 53.315 30.190 53.635 31.100 ;
        RECT 54.995 31.090 56.125 31.100 ;
        RECT 57.025 30.810 61.665 31.210 ;
        RECT 61.215 30.530 61.465 30.810 ;
        RECT 53.315 30.130 53.645 30.190 ;
        RECT 53.325 20.200 53.645 30.130 ;
        RECT 54.645 28.880 54.915 30.240 ;
        RECT 55.775 28.880 56.045 30.200 ;
        RECT 61.085 30.100 61.465 30.530 ;
        RECT 61.085 29.590 61.445 30.100 ;
        RECT 54.645 22.190 56.045 28.880 ;
        RECT 54.645 20.190 54.915 22.190 ;
        RECT 55.775 20.150 56.045 22.190 ;
        RECT 61.095 21.750 61.355 29.590 ;
        RECT 61.095 20.200 61.475 21.750 ;
        RECT 53.615 19.540 54.665 19.950 ;
        RECT 56.025 19.550 61.075 19.930 ;
        RECT 53.785 18.260 54.455 19.540 ;
        RECT 53.615 17.580 54.735 18.260 ;
        RECT 40.155 12.770 41.015 13.610 ;
        RECT 50.755 12.170 51.165 14.790 ;
        RECT 51.465 13.590 52.005 16.820 ;
        RECT 57.705 16.770 59.635 19.550 ;
        RECT 57.125 15.920 59.835 16.770 ;
        RECT 61.215 15.380 61.475 20.200 ;
        RECT 60.685 14.650 61.575 15.380 ;
        RECT 61.975 14.790 62.365 36.300 ;
        RECT 62.705 16.820 63.205 37.620 ;
        RECT 65.235 38.470 65.515 40.460 ;
        RECT 67.805 40.390 68.905 41.160 ;
        RECT 76.505 40.450 76.805 42.180 ;
        RECT 65.785 39.630 66.165 40.230 ;
        RECT 65.815 39.010 66.065 39.630 ;
        RECT 65.685 38.630 66.165 39.010 ;
        RECT 65.235 33.400 65.565 38.470 ;
        RECT 66.115 37.610 66.415 38.470 ;
        RECT 67.195 37.610 67.495 38.470 ;
        RECT 68.105 38.430 68.385 40.390 ;
        RECT 71.405 38.820 71.675 38.990 ;
        RECT 71.015 38.510 71.675 38.820 ;
        RECT 66.115 33.370 67.495 37.610 ;
        RECT 68.045 38.380 68.385 38.430 ;
        RECT 70.965 38.400 71.675 38.510 ;
        RECT 64.515 32.150 64.835 32.170 ;
        RECT 66.195 32.150 67.325 33.370 ;
        RECT 68.045 33.360 68.375 38.380 ;
        RECT 70.965 37.030 71.195 38.400 ;
        RECT 71.405 38.150 71.675 38.400 ;
        RECT 72.305 38.770 72.595 39.010 ;
        RECT 73.715 38.770 74.405 38.790 ;
        RECT 72.305 38.330 74.405 38.770 ;
        RECT 72.305 38.140 72.595 38.330 ;
        RECT 71.675 37.590 72.295 37.950 ;
        RECT 73.715 37.620 74.405 38.330 ;
        RECT 70.895 36.430 71.275 37.030 ;
        RECT 71.685 36.720 72.115 37.590 ;
        RECT 70.965 35.240 71.195 36.430 ;
        RECT 71.685 36.300 73.565 36.720 ;
        RECT 71.685 35.770 72.115 36.300 ;
        RECT 71.535 35.410 72.155 35.770 ;
        RECT 70.965 35.230 71.445 35.240 ;
        RECT 70.965 34.550 71.525 35.230 ;
        RECT 71.055 34.400 71.525 34.550 ;
        RECT 71.255 33.450 71.525 34.400 ;
        RECT 72.165 34.150 72.435 35.150 ;
        RECT 72.165 33.420 72.675 34.150 ;
        RECT 72.165 33.330 72.665 33.420 ;
        RECT 67.525 32.780 68.055 33.160 ;
        RECT 64.515 31.100 67.345 32.150 ;
        RECT 67.625 31.900 67.885 32.780 ;
        RECT 67.605 31.280 67.965 31.900 ;
        RECT 72.415 31.210 72.665 33.330 ;
        RECT 64.515 30.190 64.835 31.100 ;
        RECT 66.195 31.090 67.325 31.100 ;
        RECT 68.225 30.810 72.865 31.210 ;
        RECT 72.415 30.530 72.665 30.810 ;
        RECT 64.515 30.130 64.845 30.190 ;
        RECT 64.525 20.200 64.845 30.130 ;
        RECT 65.845 28.880 66.115 30.240 ;
        RECT 66.975 28.880 67.245 30.200 ;
        RECT 72.285 30.100 72.665 30.530 ;
        RECT 72.285 29.590 72.645 30.100 ;
        RECT 65.845 22.190 67.245 28.880 ;
        RECT 65.845 20.190 66.115 22.190 ;
        RECT 66.975 20.150 67.245 22.190 ;
        RECT 72.295 21.750 72.555 29.590 ;
        RECT 72.295 20.200 72.675 21.750 ;
        RECT 64.815 19.540 65.865 19.950 ;
        RECT 67.225 19.550 72.275 19.930 ;
        RECT 64.985 18.260 65.655 19.540 ;
        RECT 64.815 17.580 65.935 18.260 ;
        RECT 51.445 12.750 52.305 13.590 ;
        RECT 27.865 11.130 30.415 11.950 ;
        RECT 28.395 11.090 30.415 11.130 ;
        RECT 39.115 10.980 41.565 11.990 ;
        RECT 50.335 10.970 52.355 12.170 ;
        RECT 61.975 12.160 62.385 14.790 ;
        RECT 62.685 13.590 63.225 16.820 ;
        RECT 68.905 16.770 70.835 19.550 ;
        RECT 68.325 15.920 71.035 16.770 ;
        RECT 72.415 15.380 72.675 20.200 ;
        RECT 71.885 14.650 72.775 15.380 ;
        RECT 73.175 14.790 73.565 36.300 ;
        RECT 73.905 16.820 74.405 37.620 ;
        RECT 76.525 38.460 76.805 40.450 ;
        RECT 79.095 40.380 80.195 41.150 ;
        RECT 87.745 40.470 88.045 42.200 ;
        RECT 77.075 39.620 77.455 40.220 ;
        RECT 77.105 39.000 77.355 39.620 ;
        RECT 76.975 38.620 77.455 39.000 ;
        RECT 76.525 33.390 76.855 38.460 ;
        RECT 77.405 37.600 77.705 38.460 ;
        RECT 78.485 37.600 78.785 38.460 ;
        RECT 79.395 38.420 79.675 40.380 ;
        RECT 82.695 38.810 82.965 38.980 ;
        RECT 82.305 38.500 82.965 38.810 ;
        RECT 77.405 33.360 78.785 37.600 ;
        RECT 79.335 38.370 79.675 38.420 ;
        RECT 82.255 38.390 82.965 38.500 ;
        RECT 75.805 32.140 76.125 32.160 ;
        RECT 77.485 32.140 78.615 33.360 ;
        RECT 79.335 33.350 79.665 38.370 ;
        RECT 82.255 37.020 82.485 38.390 ;
        RECT 82.695 38.140 82.965 38.390 ;
        RECT 83.595 38.760 83.885 39.000 ;
        RECT 85.005 38.760 85.695 38.780 ;
        RECT 83.595 38.320 85.695 38.760 ;
        RECT 83.595 38.130 83.885 38.320 ;
        RECT 82.965 37.580 83.585 37.940 ;
        RECT 85.005 37.610 85.695 38.320 ;
        RECT 82.185 36.420 82.565 37.020 ;
        RECT 82.975 36.710 83.405 37.580 ;
        RECT 82.255 35.230 82.485 36.420 ;
        RECT 82.975 36.290 84.855 36.710 ;
        RECT 82.975 35.760 83.405 36.290 ;
        RECT 82.825 35.400 83.445 35.760 ;
        RECT 82.255 35.220 82.735 35.230 ;
        RECT 82.255 34.540 82.815 35.220 ;
        RECT 82.345 34.390 82.815 34.540 ;
        RECT 82.545 33.440 82.815 34.390 ;
        RECT 83.455 34.140 83.725 35.140 ;
        RECT 83.455 33.410 83.965 34.140 ;
        RECT 83.455 33.320 83.955 33.410 ;
        RECT 78.815 32.770 79.345 33.150 ;
        RECT 75.805 31.090 78.635 32.140 ;
        RECT 78.915 31.890 79.175 32.770 ;
        RECT 78.895 31.270 79.255 31.890 ;
        RECT 83.705 31.200 83.955 33.320 ;
        RECT 75.805 30.180 76.125 31.090 ;
        RECT 77.485 31.080 78.615 31.090 ;
        RECT 79.515 30.800 84.155 31.200 ;
        RECT 83.705 30.520 83.955 30.800 ;
        RECT 75.805 30.120 76.135 30.180 ;
        RECT 75.815 20.190 76.135 30.120 ;
        RECT 77.135 28.870 77.405 30.230 ;
        RECT 78.265 28.870 78.535 30.190 ;
        RECT 83.575 30.090 83.955 30.520 ;
        RECT 83.575 29.580 83.935 30.090 ;
        RECT 77.135 22.180 78.535 28.870 ;
        RECT 77.135 20.180 77.405 22.180 ;
        RECT 78.265 20.140 78.535 22.180 ;
        RECT 83.585 21.740 83.845 29.580 ;
        RECT 83.585 20.190 83.965 21.740 ;
        RECT 76.105 19.530 77.155 19.940 ;
        RECT 78.515 19.540 83.565 19.920 ;
        RECT 76.275 18.250 76.945 19.530 ;
        RECT 76.105 17.570 77.225 18.250 ;
        RECT 62.665 12.750 63.525 13.590 ;
        RECT 73.175 12.190 73.585 14.790 ;
        RECT 73.885 13.590 74.425 16.820 ;
        RECT 80.195 16.760 82.125 19.540 ;
        RECT 79.615 15.910 82.325 16.760 ;
        RECT 83.705 15.370 83.965 20.190 ;
        RECT 83.175 14.640 84.065 15.370 ;
        RECT 84.465 14.780 84.855 36.290 ;
        RECT 85.195 16.810 85.695 37.610 ;
        RECT 87.765 38.480 88.045 40.470 ;
        RECT 90.335 40.400 91.435 41.170 ;
        RECT 98.955 40.490 99.255 42.220 ;
        RECT 88.315 39.640 88.695 40.240 ;
        RECT 88.345 39.020 88.595 39.640 ;
        RECT 88.215 38.640 88.695 39.020 ;
        RECT 87.765 33.410 88.095 38.480 ;
        RECT 88.645 37.620 88.945 38.480 ;
        RECT 89.725 37.620 90.025 38.480 ;
        RECT 90.635 38.440 90.915 40.400 ;
        RECT 93.935 38.830 94.205 39.000 ;
        RECT 93.545 38.520 94.205 38.830 ;
        RECT 88.645 33.380 90.025 37.620 ;
        RECT 90.575 38.390 90.915 38.440 ;
        RECT 93.495 38.410 94.205 38.520 ;
        RECT 87.045 32.160 87.365 32.180 ;
        RECT 88.725 32.160 89.855 33.380 ;
        RECT 90.575 33.370 90.905 38.390 ;
        RECT 93.495 37.040 93.725 38.410 ;
        RECT 93.935 38.160 94.205 38.410 ;
        RECT 94.835 38.780 95.125 39.020 ;
        RECT 96.245 38.780 96.935 38.800 ;
        RECT 94.835 38.340 96.935 38.780 ;
        RECT 94.835 38.150 95.125 38.340 ;
        RECT 94.205 37.600 94.825 37.960 ;
        RECT 96.245 37.630 96.935 38.340 ;
        RECT 93.425 36.440 93.805 37.040 ;
        RECT 94.215 36.730 94.645 37.600 ;
        RECT 93.495 35.250 93.725 36.440 ;
        RECT 94.215 36.310 96.095 36.730 ;
        RECT 94.215 35.780 94.645 36.310 ;
        RECT 94.065 35.420 94.685 35.780 ;
        RECT 93.495 35.240 93.975 35.250 ;
        RECT 93.495 34.560 94.055 35.240 ;
        RECT 93.585 34.410 94.055 34.560 ;
        RECT 93.785 33.460 94.055 34.410 ;
        RECT 94.695 34.160 94.965 35.160 ;
        RECT 94.695 33.430 95.205 34.160 ;
        RECT 94.695 33.340 95.195 33.430 ;
        RECT 90.055 32.790 90.585 33.170 ;
        RECT 87.045 31.110 89.875 32.160 ;
        RECT 90.155 31.910 90.415 32.790 ;
        RECT 90.135 31.290 90.495 31.910 ;
        RECT 94.945 31.220 95.195 33.340 ;
        RECT 87.045 30.200 87.365 31.110 ;
        RECT 88.725 31.100 89.855 31.110 ;
        RECT 90.755 30.820 95.395 31.220 ;
        RECT 94.945 30.540 95.195 30.820 ;
        RECT 87.045 30.140 87.375 30.200 ;
        RECT 87.055 20.210 87.375 30.140 ;
        RECT 88.375 28.890 88.645 30.250 ;
        RECT 89.505 28.890 89.775 30.210 ;
        RECT 94.815 30.110 95.195 30.540 ;
        RECT 94.815 29.600 95.175 30.110 ;
        RECT 88.375 22.200 89.775 28.890 ;
        RECT 88.375 20.200 88.645 22.200 ;
        RECT 89.505 20.160 89.775 22.200 ;
        RECT 94.825 21.760 95.085 29.600 ;
        RECT 94.825 20.210 95.205 21.760 ;
        RECT 87.345 19.550 88.395 19.960 ;
        RECT 89.755 19.560 94.805 19.940 ;
        RECT 87.515 18.270 88.185 19.550 ;
        RECT 87.345 17.590 88.465 18.270 ;
        RECT 73.865 12.750 74.725 13.590 ;
        RECT 61.415 10.960 63.435 12.160 ;
        RECT 72.725 10.990 74.745 12.190 ;
        RECT 84.465 12.180 84.875 14.780 ;
        RECT 85.175 13.580 85.715 16.810 ;
        RECT 91.435 16.780 93.365 19.560 ;
        RECT 90.855 15.930 93.565 16.780 ;
        RECT 94.945 15.390 95.205 20.210 ;
        RECT 94.415 14.660 95.305 15.390 ;
        RECT 95.705 14.800 96.095 36.310 ;
        RECT 96.435 16.830 96.935 37.630 ;
        RECT 98.975 38.500 99.255 40.490 ;
        RECT 101.545 40.420 102.645 41.190 ;
        RECT 110.155 40.530 110.455 42.260 ;
        RECT 99.525 39.660 99.905 40.260 ;
        RECT 99.555 39.040 99.805 39.660 ;
        RECT 99.425 38.660 99.905 39.040 ;
        RECT 98.975 33.430 99.305 38.500 ;
        RECT 99.855 37.640 100.155 38.500 ;
        RECT 100.935 37.640 101.235 38.500 ;
        RECT 101.845 38.460 102.125 40.420 ;
        RECT 105.145 38.850 105.415 39.020 ;
        RECT 104.755 38.540 105.415 38.850 ;
        RECT 99.855 33.400 101.235 37.640 ;
        RECT 101.785 38.410 102.125 38.460 ;
        RECT 104.705 38.430 105.415 38.540 ;
        RECT 98.255 32.180 98.575 32.200 ;
        RECT 99.935 32.180 101.065 33.400 ;
        RECT 101.785 33.390 102.115 38.410 ;
        RECT 104.705 37.060 104.935 38.430 ;
        RECT 105.145 38.180 105.415 38.430 ;
        RECT 106.045 38.800 106.335 39.040 ;
        RECT 107.455 38.800 108.145 38.820 ;
        RECT 106.045 38.360 108.145 38.800 ;
        RECT 106.045 38.170 106.335 38.360 ;
        RECT 105.415 37.620 106.035 37.980 ;
        RECT 107.455 37.650 108.145 38.360 ;
        RECT 104.635 36.460 105.015 37.060 ;
        RECT 105.425 36.750 105.855 37.620 ;
        RECT 104.705 35.270 104.935 36.460 ;
        RECT 105.425 36.330 107.305 36.750 ;
        RECT 105.425 35.800 105.855 36.330 ;
        RECT 105.275 35.440 105.895 35.800 ;
        RECT 104.705 35.260 105.185 35.270 ;
        RECT 104.705 34.580 105.265 35.260 ;
        RECT 104.795 34.430 105.265 34.580 ;
        RECT 104.995 33.480 105.265 34.430 ;
        RECT 105.905 34.180 106.175 35.180 ;
        RECT 105.905 33.450 106.415 34.180 ;
        RECT 105.905 33.360 106.405 33.450 ;
        RECT 101.265 32.810 101.795 33.190 ;
        RECT 98.255 31.130 101.085 32.180 ;
        RECT 101.365 31.930 101.625 32.810 ;
        RECT 101.345 31.310 101.705 31.930 ;
        RECT 106.155 31.240 106.405 33.360 ;
        RECT 98.255 30.220 98.575 31.130 ;
        RECT 99.935 31.120 101.065 31.130 ;
        RECT 101.965 30.840 106.605 31.240 ;
        RECT 106.155 30.560 106.405 30.840 ;
        RECT 98.255 30.160 98.585 30.220 ;
        RECT 98.265 20.230 98.585 30.160 ;
        RECT 99.585 28.910 99.855 30.270 ;
        RECT 100.715 28.910 100.985 30.230 ;
        RECT 106.025 30.130 106.405 30.560 ;
        RECT 106.025 29.620 106.385 30.130 ;
        RECT 99.585 22.220 100.985 28.910 ;
        RECT 99.585 20.220 99.855 22.220 ;
        RECT 100.715 20.180 100.985 22.220 ;
        RECT 106.035 21.780 106.295 29.620 ;
        RECT 106.035 20.230 106.415 21.780 ;
        RECT 98.555 19.570 99.605 19.980 ;
        RECT 100.965 19.580 106.015 19.960 ;
        RECT 98.725 18.290 99.395 19.570 ;
        RECT 98.555 17.610 99.675 18.290 ;
        RECT 85.155 12.740 86.015 13.580 ;
        RECT 95.705 12.180 96.115 14.800 ;
        RECT 96.415 13.600 96.955 16.830 ;
        RECT 102.645 16.800 104.575 19.580 ;
        RECT 102.065 15.950 104.775 16.800 ;
        RECT 106.155 15.410 106.415 20.230 ;
        RECT 105.625 14.680 106.515 15.410 ;
        RECT 106.915 14.820 107.305 36.330 ;
        RECT 107.645 16.850 108.145 37.650 ;
        RECT 110.175 38.540 110.455 40.530 ;
        RECT 112.745 40.460 113.845 41.230 ;
        RECT 121.365 40.550 121.665 42.280 ;
        RECT 142.880 42.020 144.100 43.390 ;
        RECT 110.725 39.700 111.105 40.300 ;
        RECT 110.755 39.080 111.005 39.700 ;
        RECT 110.625 38.700 111.105 39.080 ;
        RECT 110.175 33.470 110.505 38.540 ;
        RECT 111.055 37.680 111.355 38.540 ;
        RECT 112.135 37.680 112.435 38.540 ;
        RECT 113.045 38.500 113.325 40.460 ;
        RECT 116.345 38.890 116.615 39.060 ;
        RECT 115.955 38.580 116.615 38.890 ;
        RECT 111.055 33.440 112.435 37.680 ;
        RECT 112.985 38.450 113.325 38.500 ;
        RECT 115.905 38.470 116.615 38.580 ;
        RECT 109.455 32.220 109.775 32.240 ;
        RECT 111.135 32.220 112.265 33.440 ;
        RECT 112.985 33.430 113.315 38.450 ;
        RECT 115.905 37.100 116.135 38.470 ;
        RECT 116.345 38.220 116.615 38.470 ;
        RECT 117.245 38.840 117.535 39.080 ;
        RECT 118.655 38.840 119.345 38.860 ;
        RECT 117.245 38.400 119.345 38.840 ;
        RECT 117.245 38.210 117.535 38.400 ;
        RECT 116.615 37.660 117.235 38.020 ;
        RECT 118.655 37.690 119.345 38.400 ;
        RECT 115.835 36.500 116.215 37.100 ;
        RECT 116.625 36.790 117.055 37.660 ;
        RECT 115.905 35.310 116.135 36.500 ;
        RECT 116.625 36.370 118.505 36.790 ;
        RECT 116.625 35.840 117.055 36.370 ;
        RECT 116.475 35.480 117.095 35.840 ;
        RECT 115.905 35.300 116.385 35.310 ;
        RECT 115.905 34.620 116.465 35.300 ;
        RECT 115.995 34.470 116.465 34.620 ;
        RECT 116.195 33.520 116.465 34.470 ;
        RECT 117.105 34.220 117.375 35.220 ;
        RECT 117.105 33.490 117.615 34.220 ;
        RECT 117.105 33.400 117.605 33.490 ;
        RECT 112.465 32.850 112.995 33.230 ;
        RECT 109.455 31.170 112.285 32.220 ;
        RECT 112.565 31.970 112.825 32.850 ;
        RECT 112.545 31.350 112.905 31.970 ;
        RECT 117.355 31.280 117.605 33.400 ;
        RECT 109.455 30.260 109.775 31.170 ;
        RECT 111.135 31.160 112.265 31.170 ;
        RECT 113.165 30.880 117.805 31.280 ;
        RECT 117.355 30.600 117.605 30.880 ;
        RECT 109.455 30.200 109.785 30.260 ;
        RECT 109.465 20.270 109.785 30.200 ;
        RECT 110.785 28.950 111.055 30.310 ;
        RECT 111.915 28.950 112.185 30.270 ;
        RECT 117.225 30.170 117.605 30.600 ;
        RECT 117.225 29.660 117.585 30.170 ;
        RECT 110.785 22.260 112.185 28.950 ;
        RECT 110.785 20.260 111.055 22.260 ;
        RECT 111.915 20.220 112.185 22.260 ;
        RECT 117.235 21.820 117.495 29.660 ;
        RECT 117.235 20.270 117.615 21.820 ;
        RECT 109.755 19.610 110.805 20.020 ;
        RECT 112.165 19.620 117.215 20.000 ;
        RECT 109.925 18.330 110.595 19.610 ;
        RECT 109.755 17.650 110.875 18.330 ;
        RECT 96.395 12.760 97.255 13.600 ;
        RECT 106.915 12.230 107.325 14.820 ;
        RECT 107.625 13.620 108.165 16.850 ;
        RECT 113.845 16.840 115.775 19.620 ;
        RECT 113.265 15.990 115.975 16.840 ;
        RECT 117.355 15.450 117.615 20.270 ;
        RECT 116.825 14.720 117.715 15.450 ;
        RECT 118.115 14.860 118.505 36.370 ;
        RECT 118.845 16.890 119.345 37.690 ;
        RECT 121.385 38.560 121.665 40.550 ;
        RECT 123.955 40.480 125.055 41.250 ;
        RECT 121.935 39.720 122.315 40.320 ;
        RECT 121.965 39.100 122.215 39.720 ;
        RECT 121.835 38.720 122.315 39.100 ;
        RECT 121.385 33.490 121.715 38.560 ;
        RECT 122.265 37.700 122.565 38.560 ;
        RECT 123.345 37.700 123.645 38.560 ;
        RECT 124.255 38.520 124.535 40.480 ;
        RECT 127.555 38.910 127.825 39.080 ;
        RECT 127.165 38.600 127.825 38.910 ;
        RECT 122.265 33.460 123.645 37.700 ;
        RECT 124.195 38.470 124.535 38.520 ;
        RECT 127.115 38.490 127.825 38.600 ;
        RECT 120.665 32.240 120.985 32.260 ;
        RECT 122.345 32.240 123.475 33.460 ;
        RECT 124.195 33.450 124.525 38.470 ;
        RECT 127.115 37.120 127.345 38.490 ;
        RECT 127.555 38.240 127.825 38.490 ;
        RECT 128.455 38.860 128.745 39.100 ;
        RECT 142.940 38.950 144.100 42.020 ;
        RECT 129.865 38.860 130.555 38.880 ;
        RECT 128.455 38.420 130.555 38.860 ;
        RECT 128.455 38.230 128.745 38.420 ;
        RECT 127.825 37.680 128.445 38.040 ;
        RECT 129.865 37.710 130.555 38.420 ;
        RECT 127.045 36.520 127.425 37.120 ;
        RECT 127.835 36.810 128.265 37.680 ;
        RECT 127.115 35.330 127.345 36.520 ;
        RECT 127.835 36.390 129.715 36.810 ;
        RECT 127.835 35.860 128.265 36.390 ;
        RECT 127.685 35.500 128.305 35.860 ;
        RECT 127.115 35.320 127.595 35.330 ;
        RECT 127.115 34.640 127.675 35.320 ;
        RECT 127.205 34.490 127.675 34.640 ;
        RECT 127.405 33.540 127.675 34.490 ;
        RECT 128.315 34.240 128.585 35.240 ;
        RECT 128.315 33.510 128.825 34.240 ;
        RECT 128.315 33.420 128.815 33.510 ;
        RECT 123.675 32.870 124.205 33.250 ;
        RECT 120.665 31.190 123.495 32.240 ;
        RECT 123.775 31.990 124.035 32.870 ;
        RECT 123.755 31.370 124.115 31.990 ;
        RECT 128.565 31.300 128.815 33.420 ;
        RECT 120.665 30.280 120.985 31.190 ;
        RECT 122.345 31.180 123.475 31.190 ;
        RECT 124.375 30.900 129.015 31.300 ;
        RECT 128.565 30.620 128.815 30.900 ;
        RECT 120.665 30.220 120.995 30.280 ;
        RECT 120.675 20.290 120.995 30.220 ;
        RECT 121.995 28.970 122.265 30.330 ;
        RECT 123.125 28.970 123.395 30.290 ;
        RECT 128.435 30.190 128.815 30.620 ;
        RECT 128.435 29.680 128.795 30.190 ;
        RECT 121.995 22.280 123.395 28.970 ;
        RECT 121.995 20.280 122.265 22.280 ;
        RECT 123.125 20.240 123.395 22.280 ;
        RECT 128.445 21.840 128.705 29.680 ;
        RECT 128.445 20.290 128.825 21.840 ;
        RECT 120.965 19.630 122.015 20.040 ;
        RECT 123.375 19.640 128.425 20.020 ;
        RECT 121.135 18.350 121.805 19.630 ;
        RECT 120.965 17.670 122.085 18.350 ;
        RECT 107.605 12.780 108.465 13.620 ;
        RECT 118.115 12.230 118.525 14.860 ;
        RECT 118.825 13.660 119.365 16.890 ;
        RECT 125.055 16.860 126.985 19.640 ;
        RECT 124.475 16.010 127.185 16.860 ;
        RECT 128.565 15.470 128.825 20.290 ;
        RECT 128.035 14.740 128.925 15.470 ;
        RECT 129.325 14.880 129.715 36.390 ;
        RECT 130.055 16.910 130.555 37.710 ;
        RECT 142.900 37.580 144.120 38.950 ;
        RECT 132.395 24.340 132.705 30.230 ;
        RECT 132.195 20.120 132.705 24.340 ;
        RECT 118.805 12.820 119.665 13.660 ;
        RECT 129.325 12.260 129.735 14.880 ;
        RECT 130.035 13.680 130.575 16.910 ;
        RECT 132.195 15.510 132.505 20.120 ;
        RECT 137.715 19.980 138.005 30.170 ;
        RECT 132.685 19.590 138.005 19.980 ;
        RECT 137.715 16.940 138.005 19.590 ;
        RECT 142.940 17.940 144.090 19.160 ;
        RECT 145.080 18.760 146.200 18.930 ;
        RECT 137.395 15.890 138.295 16.940 ;
        RECT 137.715 15.720 138.005 15.890 ;
        RECT 131.975 14.270 132.735 15.510 ;
        RECT 142.940 15.090 144.050 17.940 ;
        RECT 142.900 13.870 144.050 15.090 ;
        RECT 145.070 14.920 146.200 18.760 ;
        RECT 145.030 13.970 146.200 14.920 ;
        RECT 145.030 13.900 146.150 13.970 ;
        RECT 130.015 12.840 130.875 13.680 ;
        RECT 83.845 10.980 85.865 12.180 ;
        RECT 95.145 10.980 97.165 12.180 ;
        RECT 106.335 11.030 108.355 12.230 ;
        RECT 117.565 11.030 119.585 12.230 ;
        RECT 128.865 11.060 130.885 12.260 ;
        RECT 74.340 0.110 75.630 1.460 ;
        RECT 93.550 0.180 94.840 1.530 ;
        RECT 112.950 0.310 114.240 1.660 ;
        RECT 131.850 0.380 133.490 1.930 ;
        RECT 151.650 0.250 152.920 1.470 ;
      LAYER met3 ;
        RECT 135.340 223.855 136.790 225.205 ;
        RECT 138.130 223.785 139.580 225.135 ;
        RECT 143.180 223.815 144.630 225.165 ;
        RECT 16.830 211.125 18.810 211.455 ;
        RECT 46.830 211.125 48.810 211.455 ;
        RECT 76.830 211.125 78.810 211.455 ;
        RECT 106.830 211.125 108.810 211.455 ;
        RECT 31.830 208.405 33.810 208.735 ;
        RECT 61.830 208.405 63.810 208.735 ;
        RECT 91.830 208.405 93.810 208.735 ;
        RECT 121.830 208.405 123.810 208.735 ;
        RECT 16.830 205.685 18.810 206.015 ;
        RECT 46.830 205.685 48.810 206.015 ;
        RECT 76.830 205.685 78.810 206.015 ;
        RECT 106.830 205.685 108.810 206.015 ;
        RECT 31.830 202.965 33.810 203.295 ;
        RECT 61.830 202.965 63.810 203.295 ;
        RECT 91.830 202.965 93.810 203.295 ;
        RECT 121.830 202.965 123.810 203.295 ;
        RECT 16.830 200.245 18.810 200.575 ;
        RECT 46.830 200.245 48.810 200.575 ;
        RECT 76.830 200.245 78.810 200.575 ;
        RECT 106.830 200.245 108.810 200.575 ;
        RECT 31.830 197.525 33.810 197.855 ;
        RECT 61.830 197.525 63.810 197.855 ;
        RECT 91.830 197.525 93.810 197.855 ;
        RECT 121.830 197.525 123.810 197.855 ;
        RECT 16.830 194.805 18.810 195.135 ;
        RECT 46.830 194.805 48.810 195.135 ;
        RECT 76.830 194.805 78.810 195.135 ;
        RECT 106.830 194.805 108.810 195.135 ;
        RECT 31.830 192.085 33.810 192.415 ;
        RECT 61.830 192.085 63.810 192.415 ;
        RECT 91.830 192.085 93.810 192.415 ;
        RECT 121.830 192.085 123.810 192.415 ;
        RECT 16.830 189.365 18.810 189.695 ;
        RECT 46.830 189.365 48.810 189.695 ;
        RECT 76.830 189.365 78.810 189.695 ;
        RECT 106.830 189.365 108.810 189.695 ;
        RECT 31.830 186.645 33.810 186.975 ;
        RECT 61.830 186.645 63.810 186.975 ;
        RECT 91.830 186.645 93.810 186.975 ;
        RECT 121.830 186.645 123.810 186.975 ;
        RECT 16.830 183.925 18.810 184.255 ;
        RECT 46.830 183.925 48.810 184.255 ;
        RECT 76.830 183.925 78.810 184.255 ;
        RECT 106.830 183.925 108.810 184.255 ;
        RECT 31.830 181.205 33.810 181.535 ;
        RECT 61.830 181.205 63.810 181.535 ;
        RECT 91.830 181.205 93.810 181.535 ;
        RECT 121.830 181.205 123.810 181.535 ;
        RECT 16.830 178.485 18.810 178.815 ;
        RECT 46.830 178.485 48.810 178.815 ;
        RECT 76.830 178.485 78.810 178.815 ;
        RECT 106.830 178.485 108.810 178.815 ;
        RECT 80.505 176.420 80.835 176.435 ;
        RECT 81.170 176.420 81.550 176.430 ;
        RECT 80.505 176.120 81.550 176.420 ;
        RECT 80.505 176.105 80.835 176.120 ;
        RECT 81.170 176.110 81.550 176.120 ;
        RECT 31.830 175.765 33.810 176.095 ;
        RECT 61.830 175.765 63.810 176.095 ;
        RECT 91.830 175.765 93.810 176.095 ;
        RECT 121.830 175.765 123.810 176.095 ;
        RECT 50.605 175.060 50.935 175.075 ;
        RECT 79.125 175.060 79.455 175.075 ;
        RECT 50.605 174.760 79.455 175.060 ;
        RECT 50.605 174.745 50.935 174.760 ;
        RECT 79.125 174.745 79.455 174.760 ;
        RECT 36.345 174.380 36.675 174.395 ;
        RECT 45.545 174.380 45.875 174.395 ;
        RECT 64.610 174.380 64.990 174.390 ;
        RECT 92.925 174.380 93.255 174.395 ;
        RECT 36.345 174.080 98.990 174.380 ;
        RECT 36.345 174.065 36.675 174.080 ;
        RECT 45.545 174.065 45.875 174.080 ;
        RECT 64.610 174.070 64.990 174.080 ;
        RECT 92.925 174.065 93.255 174.080 ;
        RECT 98.690 173.700 98.990 174.080 ;
        RECT 105.805 173.700 106.135 173.715 ;
        RECT 98.690 173.400 106.135 173.700 ;
        RECT 105.805 173.385 106.135 173.400 ;
        RECT 16.830 173.045 18.810 173.375 ;
        RECT 46.830 173.045 48.810 173.375 ;
        RECT 76.830 173.045 78.810 173.375 ;
        RECT 106.830 173.045 108.810 173.375 ;
        RECT 133.700 172.500 134.930 172.705 ;
        RECT 31.830 170.325 33.810 170.655 ;
        RECT 61.830 170.325 63.810 170.655 ;
        RECT 91.830 170.325 93.810 170.655 ;
        RECT 121.830 170.325 123.810 170.655 ;
        RECT 129.030 170.130 134.930 172.500 ;
        RECT 133.700 170.095 134.930 170.130 ;
        RECT 16.830 167.605 18.810 167.935 ;
        RECT 46.830 167.605 48.810 167.935 ;
        RECT 76.830 167.605 78.810 167.935 ;
        RECT 106.830 167.605 108.810 167.935 ;
        RECT 31.830 164.885 33.810 165.215 ;
        RECT 61.830 164.885 63.810 165.215 ;
        RECT 91.830 164.885 93.810 165.215 ;
        RECT 121.830 164.885 123.810 165.215 ;
        RECT 69.925 163.500 70.255 163.515 ;
        RECT 115.925 163.500 116.255 163.515 ;
        RECT 69.925 163.200 116.255 163.500 ;
        RECT 69.925 163.185 70.255 163.200 ;
        RECT 115.925 163.185 116.255 163.200 ;
        RECT 16.830 162.165 18.810 162.495 ;
        RECT 46.830 162.165 48.810 162.495 ;
        RECT 76.830 162.165 78.810 162.495 ;
        RECT 106.830 162.165 108.810 162.495 ;
        RECT 31.830 159.445 33.810 159.775 ;
        RECT 61.830 159.445 63.810 159.775 ;
        RECT 91.830 159.445 93.810 159.775 ;
        RECT 121.830 159.445 123.810 159.775 ;
        RECT 16.830 156.725 18.810 157.055 ;
        RECT 46.830 156.725 48.810 157.055 ;
        RECT 76.830 156.725 78.810 157.055 ;
        RECT 106.830 156.725 108.810 157.055 ;
        RECT 102.585 156.020 102.915 156.035 ;
        RECT 106.725 156.020 107.055 156.035 ;
        RECT 109.485 156.020 109.815 156.035 ;
        RECT 102.585 155.720 109.815 156.020 ;
        RECT 102.585 155.705 102.915 155.720 ;
        RECT 106.725 155.705 107.055 155.720 ;
        RECT 109.485 155.705 109.815 155.720 ;
        RECT 31.830 154.005 33.810 154.335 ;
        RECT 61.830 154.005 63.810 154.335 ;
        RECT 91.830 154.005 93.810 154.335 ;
        RECT 121.830 154.005 123.810 154.335 ;
        RECT 38.185 153.300 38.515 153.315 ;
        RECT 68.545 153.300 68.875 153.315 ;
        RECT 38.185 153.000 68.875 153.300 ;
        RECT 38.185 152.985 38.515 153.000 ;
        RECT 68.545 152.985 68.875 153.000 ;
        RECT 45.545 152.620 45.875 152.635 ;
        RECT 45.330 152.305 45.875 152.620 ;
        RECT 63.945 152.620 64.275 152.635 ;
        RECT 72.685 152.620 73.015 152.635 ;
        RECT 63.945 152.320 73.015 152.620 ;
        RECT 63.945 152.305 64.275 152.320 ;
        RECT 72.685 152.305 73.015 152.320 ;
        RECT 44.165 151.940 44.495 151.955 ;
        RECT 45.330 151.940 45.630 152.305 ;
        RECT 44.165 151.640 45.630 151.940 ;
        RECT 44.165 151.625 44.495 151.640 ;
        RECT 16.830 151.285 18.810 151.615 ;
        RECT 46.830 151.285 48.810 151.615 ;
        RECT 76.830 151.285 78.810 151.615 ;
        RECT 106.830 151.285 108.810 151.615 ;
        RECT 64.865 149.230 65.195 149.235 ;
        RECT 64.610 149.220 65.195 149.230 ;
        RECT 64.610 148.920 65.420 149.220 ;
        RECT 64.610 148.910 65.195 148.920 ;
        RECT 64.865 148.905 65.195 148.910 ;
        RECT 31.830 148.565 33.810 148.895 ;
        RECT 61.830 148.565 63.810 148.895 ;
        RECT 91.830 148.565 93.810 148.895 ;
        RECT 121.830 148.565 123.810 148.895 ;
        RECT 72.225 146.500 72.555 146.515 ;
        RECT 75.650 146.500 76.030 146.510 ;
        RECT 72.225 146.200 76.030 146.500 ;
        RECT 72.225 146.185 72.555 146.200 ;
        RECT 75.650 146.190 76.030 146.200 ;
        RECT 16.830 145.845 18.810 146.175 ;
        RECT 46.830 145.845 48.810 146.175 ;
        RECT 76.830 145.845 78.810 146.175 ;
        RECT 106.830 145.845 108.810 146.175 ;
        RECT 50.605 144.460 50.935 144.475 ;
        RECT 53.365 144.460 53.695 144.475 ;
        RECT 68.545 144.460 68.875 144.475 ;
        RECT 50.605 144.160 68.875 144.460 ;
        RECT 50.605 144.145 50.935 144.160 ;
        RECT 53.365 144.145 53.695 144.160 ;
        RECT 68.545 144.145 68.875 144.160 ;
        RECT 78.205 143.780 78.535 143.795 ;
        RECT 80.250 143.780 80.630 143.790 ;
        RECT 78.205 143.480 80.630 143.780 ;
        RECT 78.205 143.465 78.535 143.480 ;
        RECT 80.250 143.470 80.630 143.480 ;
        RECT 31.830 143.125 33.810 143.455 ;
        RECT 61.830 143.125 63.810 143.455 ;
        RECT 91.830 143.125 93.810 143.455 ;
        RECT 121.830 143.125 123.810 143.455 ;
        RECT 16.830 140.405 18.810 140.735 ;
        RECT 46.830 140.405 48.810 140.735 ;
        RECT 76.830 140.405 78.810 140.735 ;
        RECT 106.830 140.405 108.810 140.735 ;
        RECT 75.650 139.020 76.030 139.030 ;
        RECT 129.090 139.020 134.150 139.430 ;
        RECT 75.650 138.720 134.150 139.020 ;
        RECT 75.650 138.710 76.030 138.720 ;
        RECT 129.090 138.200 134.150 138.720 ;
        RECT 31.830 137.685 33.810 138.015 ;
        RECT 61.830 137.685 63.810 138.015 ;
        RECT 91.830 137.685 93.810 138.015 ;
        RECT 121.830 137.685 123.810 138.015 ;
        RECT 16.830 134.965 18.810 135.295 ;
        RECT 46.830 134.965 48.810 135.295 ;
        RECT 76.830 134.965 78.810 135.295 ;
        RECT 106.830 134.965 108.810 135.295 ;
        RECT 31.830 132.245 33.810 132.575 ;
        RECT 61.830 132.245 63.810 132.575 ;
        RECT 91.830 132.245 93.810 132.575 ;
        RECT 121.830 132.245 123.810 132.575 ;
        RECT 81.425 132.230 81.755 132.235 ;
        RECT 81.170 132.220 81.755 132.230 ;
        RECT 80.970 131.920 81.755 132.220 ;
        RECT 81.170 131.910 81.755 131.920 ;
        RECT 81.425 131.905 81.755 131.910 ;
        RECT 16.830 129.525 18.810 129.855 ;
        RECT 46.830 129.525 48.810 129.855 ;
        RECT 76.830 129.525 78.810 129.855 ;
        RECT 106.830 129.525 108.810 129.855 ;
        RECT 31.830 126.805 33.810 127.135 ;
        RECT 61.830 126.805 63.810 127.135 ;
        RECT 91.830 126.805 93.810 127.135 ;
        RECT 121.830 126.805 123.810 127.135 ;
        RECT 45.545 125.420 45.875 125.435 ;
        RECT 77.745 125.420 78.075 125.435 ;
        RECT 45.545 125.120 78.075 125.420 ;
        RECT 45.545 125.105 45.875 125.120 ;
        RECT 77.745 125.105 78.075 125.120 ;
        RECT 16.830 124.085 18.810 124.415 ;
        RECT 46.830 124.085 48.810 124.415 ;
        RECT 76.830 124.085 78.810 124.415 ;
        RECT 106.830 124.085 108.810 124.415 ;
        RECT 56.125 122.700 56.455 122.715 ;
        RECT 64.610 122.700 64.990 122.710 ;
        RECT 88.325 122.700 88.655 122.715 ;
        RECT 102.125 122.700 102.455 122.715 ;
        RECT 56.125 122.400 102.455 122.700 ;
        RECT 56.125 122.385 56.455 122.400 ;
        RECT 64.610 122.390 64.990 122.400 ;
        RECT 88.325 122.385 88.655 122.400 ;
        RECT 102.125 122.385 102.455 122.400 ;
        RECT 31.830 121.365 33.810 121.695 ;
        RECT 61.830 121.365 63.810 121.695 ;
        RECT 91.830 121.365 93.810 121.695 ;
        RECT 121.830 121.365 123.810 121.695 ;
        RECT 36.345 119.980 36.675 119.995 ;
        RECT 56.125 119.980 56.455 119.995 ;
        RECT 36.345 119.680 56.455 119.980 ;
        RECT 36.345 119.665 36.675 119.680 ;
        RECT 56.125 119.665 56.455 119.680 ;
        RECT 16.830 118.645 18.810 118.975 ;
        RECT 46.830 118.645 48.810 118.975 ;
        RECT 76.830 118.645 78.810 118.975 ;
        RECT 106.830 118.645 108.810 118.975 ;
        RECT 31.830 115.925 33.810 116.255 ;
        RECT 61.830 115.925 63.810 116.255 ;
        RECT 91.830 115.925 93.810 116.255 ;
        RECT 121.830 115.925 123.810 116.255 ;
        RECT 16.830 113.205 18.810 113.535 ;
        RECT 46.830 113.205 48.810 113.535 ;
        RECT 76.830 113.205 78.810 113.535 ;
        RECT 106.830 113.205 108.810 113.535 ;
        RECT 79.585 111.820 79.915 111.835 ;
        RECT 80.250 111.820 80.630 111.830 ;
        RECT 79.585 111.520 80.630 111.820 ;
        RECT 79.585 111.505 79.915 111.520 ;
        RECT 80.250 111.510 80.630 111.520 ;
        RECT 31.830 110.485 33.810 110.815 ;
        RECT 61.830 110.485 63.810 110.815 ;
        RECT 91.830 110.485 93.810 110.815 ;
        RECT 121.830 110.485 123.810 110.815 ;
        RECT 16.830 107.765 18.810 108.095 ;
        RECT 46.830 107.765 48.810 108.095 ;
        RECT 76.830 107.765 78.810 108.095 ;
        RECT 106.830 107.765 108.810 108.095 ;
        RECT 129.700 106.530 133.210 106.625 ;
        RECT 126.505 106.380 126.835 106.395 ;
        RECT 129.700 106.380 133.340 106.530 ;
        RECT 126.505 106.080 133.340 106.380 ;
        RECT 126.505 106.065 126.835 106.080 ;
        RECT 129.700 105.930 133.340 106.080 ;
        RECT 129.700 105.605 133.210 105.930 ;
        RECT 31.830 105.045 33.810 105.375 ;
        RECT 61.830 105.045 63.810 105.375 ;
        RECT 91.830 105.045 93.810 105.375 ;
        RECT 121.830 105.045 123.810 105.375 ;
        RECT 16.830 102.325 18.810 102.655 ;
        RECT 46.830 102.325 48.810 102.655 ;
        RECT 76.830 102.325 78.810 102.655 ;
        RECT 106.830 102.325 108.810 102.655 ;
        RECT 31.830 99.605 33.810 99.935 ;
        RECT 61.830 99.605 63.810 99.935 ;
        RECT 91.830 99.605 93.810 99.935 ;
        RECT 121.830 99.605 123.810 99.935 ;
        RECT 37.630 88.620 38.970 88.755 ;
        RECT 13.950 87.980 14.980 88.515 ;
        RECT 13.950 87.500 14.990 87.980 ;
        RECT 13.950 87.175 14.980 87.500 ;
        RECT 14.070 86.570 14.810 87.175 ;
        RECT 20.050 87.105 20.920 88.515 ;
        RECT 14.070 75.715 14.700 86.570 ;
        RECT 20.170 77.115 20.800 87.105 ;
        RECT 25.910 87.055 26.860 88.515 ;
        RECT 26.070 78.385 26.700 87.055 ;
        RECT 31.730 86.965 32.910 88.585 ;
        RECT 32.005 79.615 32.635 86.965 ;
        RECT 37.630 86.835 39.120 88.620 ;
        RECT 38.060 81.125 38.690 86.835 ;
        RECT 43.790 86.745 45.190 88.605 ;
        RECT 49.710 86.945 51.060 88.615 ;
        RECT 44.175 82.625 44.805 86.745 ;
        RECT 50.070 83.875 50.700 86.945 ;
        RECT 55.530 86.785 56.750 88.545 ;
        RECT 55.825 85.115 56.455 86.785 ;
        RECT 61.670 86.625 63.180 88.615 ;
        RECT 67.680 88.305 68.720 89.815 ;
        RECT 67.885 87.225 68.515 88.305 ;
        RECT 62.110 86.175 62.740 86.625 ;
        RECT 67.885 86.595 130.605 87.225 ;
        RECT 62.110 85.545 118.855 86.175 ;
        RECT 55.825 84.485 107.605 85.115 ;
        RECT 50.070 83.245 96.285 83.875 ;
        RECT 44.175 81.995 85.055 82.625 ;
        RECT 38.060 80.495 73.765 81.125 ;
        RECT 32.005 78.985 62.635 79.615 ;
        RECT 26.070 77.755 51.245 78.385 ;
        RECT 20.170 76.485 40.645 77.115 ;
        RECT 14.070 75.660 29.295 75.715 ;
        RECT 40.015 75.710 40.645 76.485 ;
        RECT 14.070 75.085 30.410 75.660 ;
        RECT 27.850 74.670 30.410 75.085 ;
        RECT 3.910 71.345 6.100 73.215 ;
        RECT 27.850 73.120 30.450 74.670 ;
        RECT 39.060 74.510 41.620 75.710 ;
        RECT 50.615 75.580 51.245 77.755 ;
        RECT 62.005 75.690 62.635 78.985 ;
        RECT 49.930 74.650 52.490 75.580 ;
        RECT 0.970 70.330 3.070 70.430 ;
        RECT 15.510 70.330 17.040 71.185 ;
        RECT 0.960 68.750 17.040 70.330 ;
        RECT 0.970 68.710 3.070 68.750 ;
        RECT 15.510 68.635 17.040 68.750 ;
        RECT 20.145 54.060 20.605 54.135 ;
        RECT 25.715 54.060 26.175 54.085 ;
        RECT 20.145 53.620 26.175 54.060 ;
        RECT 20.145 53.565 20.605 53.620 ;
        RECT 25.715 53.515 26.175 53.620 ;
        RECT 22.405 48.870 22.885 48.935 ;
        RECT 22.405 48.550 24.205 48.870 ;
        RECT 22.405 48.385 22.885 48.550 ;
        RECT 23.635 45.710 24.195 48.550 ;
        RECT 27.515 45.710 27.995 45.735 ;
        RECT 23.635 45.290 27.995 45.710 ;
        RECT 23.635 45.280 24.195 45.290 ;
        RECT 27.515 45.185 27.995 45.290 ;
        RECT 20.745 40.120 21.225 40.225 ;
        RECT 24.545 40.120 25.105 40.130 ;
        RECT 20.745 39.700 25.105 40.120 ;
        RECT 20.745 39.675 21.225 39.700 ;
        RECT 24.545 36.860 25.105 39.700 ;
        RECT 25.855 36.860 26.335 37.025 ;
        RECT 24.535 36.540 26.335 36.860 ;
        RECT 25.855 36.475 26.335 36.540 ;
        RECT 22.565 31.790 23.025 31.895 ;
        RECT 28.135 31.790 28.595 31.845 ;
        RECT 22.565 31.350 28.595 31.790 ;
        RECT 22.565 31.325 23.025 31.350 ;
        RECT 28.135 31.275 28.595 31.350 ;
        RECT 29.765 12.265 30.255 73.120 ;
        RECT 38.960 73.080 41.730 74.510 ;
        RECT 31.345 54.070 31.805 54.145 ;
        RECT 36.915 54.070 37.375 54.095 ;
        RECT 31.345 53.630 37.375 54.070 ;
        RECT 31.345 53.575 31.805 53.630 ;
        RECT 36.915 53.525 37.375 53.630 ;
        RECT 33.605 48.880 34.085 48.945 ;
        RECT 33.605 48.560 35.405 48.880 ;
        RECT 33.605 48.395 34.085 48.560 ;
        RECT 34.835 45.720 35.395 48.560 ;
        RECT 38.715 45.720 39.195 45.745 ;
        RECT 34.835 45.300 39.195 45.720 ;
        RECT 34.835 45.290 35.395 45.300 ;
        RECT 38.715 45.195 39.195 45.300 ;
        RECT 32.025 40.120 32.505 40.225 ;
        RECT 35.825 40.120 36.385 40.130 ;
        RECT 32.025 39.700 36.385 40.120 ;
        RECT 32.025 39.675 32.505 39.700 ;
        RECT 35.825 36.860 36.385 39.700 ;
        RECT 37.135 36.860 37.615 37.025 ;
        RECT 35.815 36.540 37.615 36.860 ;
        RECT 37.135 36.475 37.615 36.540 ;
        RECT 33.845 31.790 34.305 31.895 ;
        RECT 39.415 31.790 39.875 31.845 ;
        RECT 33.845 31.350 39.875 31.790 ;
        RECT 33.845 31.325 34.305 31.350 ;
        RECT 39.415 31.275 39.875 31.350 ;
        RECT 41.055 12.360 41.545 73.080 ;
        RECT 49.930 73.030 52.530 74.650 ;
        RECT 61.330 74.530 63.890 75.690 ;
        RECT 73.135 75.580 73.765 80.495 ;
        RECT 84.425 75.690 85.055 81.995 ;
        RECT 72.340 74.980 74.900 75.580 ;
        RECT 42.565 54.040 43.025 54.115 ;
        RECT 48.135 54.040 48.595 54.065 ;
        RECT 42.565 53.600 48.595 54.040 ;
        RECT 42.565 53.545 43.025 53.600 ;
        RECT 48.135 53.495 48.595 53.600 ;
        RECT 44.825 48.850 45.305 48.915 ;
        RECT 44.825 48.530 46.625 48.850 ;
        RECT 44.825 48.365 45.305 48.530 ;
        RECT 46.055 45.690 46.615 48.530 ;
        RECT 49.935 45.690 50.415 45.715 ;
        RECT 46.055 45.270 50.415 45.690 ;
        RECT 46.055 45.260 46.615 45.270 ;
        RECT 49.935 45.165 50.415 45.270 ;
        RECT 43.315 40.100 43.795 40.205 ;
        RECT 47.115 40.100 47.675 40.110 ;
        RECT 43.315 39.680 47.675 40.100 ;
        RECT 43.315 39.655 43.795 39.680 ;
        RECT 47.115 36.840 47.675 39.680 ;
        RECT 48.425 36.840 48.905 37.005 ;
        RECT 47.105 36.520 48.905 36.840 ;
        RECT 48.425 36.455 48.905 36.520 ;
        RECT 45.135 31.770 45.595 31.875 ;
        RECT 50.705 31.770 51.165 31.825 ;
        RECT 45.135 31.330 51.165 31.770 ;
        RECT 45.135 31.305 45.595 31.330 ;
        RECT 50.705 31.255 51.165 31.330 ;
        RECT 41.055 12.350 41.555 12.360 ;
        RECT 28.345 11.115 30.465 12.265 ;
        RECT 41.065 11.965 41.555 12.350 ;
        RECT 51.635 12.145 52.125 73.030 ;
        RECT 61.260 73.010 64.060 74.530 ;
        RECT 72.340 73.050 75.020 74.980 ;
        RECT 83.730 74.540 86.290 75.690 ;
        RECT 95.655 75.580 96.285 83.245 ;
        RECT 106.975 75.640 107.605 84.485 ;
        RECT 118.225 75.650 118.855 85.545 ;
        RECT 129.975 75.650 130.605 86.595 ;
        RECT 133.330 76.605 136.060 77.855 ;
        RECT 137.190 76.585 139.920 77.835 ;
        RECT 53.815 54.020 54.275 54.095 ;
        RECT 59.385 54.020 59.845 54.045 ;
        RECT 53.815 53.580 59.845 54.020 ;
        RECT 53.815 53.525 54.275 53.580 ;
        RECT 59.385 53.475 59.845 53.580 ;
        RECT 56.075 48.830 56.555 48.895 ;
        RECT 56.075 48.510 57.875 48.830 ;
        RECT 56.075 48.345 56.555 48.510 ;
        RECT 57.305 45.670 57.865 48.510 ;
        RECT 61.185 45.670 61.665 45.695 ;
        RECT 57.305 45.250 61.665 45.670 ;
        RECT 57.305 45.240 57.865 45.250 ;
        RECT 61.185 45.145 61.665 45.250 ;
        RECT 54.535 40.100 55.015 40.205 ;
        RECT 58.335 40.100 58.895 40.110 ;
        RECT 54.535 39.680 58.895 40.100 ;
        RECT 54.535 39.655 55.015 39.680 ;
        RECT 58.335 36.840 58.895 39.680 ;
        RECT 59.645 36.840 60.125 37.005 ;
        RECT 58.325 36.520 60.125 36.840 ;
        RECT 59.645 36.455 60.125 36.520 ;
        RECT 56.355 31.770 56.815 31.875 ;
        RECT 61.925 31.770 62.385 31.825 ;
        RECT 56.355 31.330 62.385 31.770 ;
        RECT 56.355 31.305 56.815 31.330 ;
        RECT 61.925 31.255 62.385 31.330 ;
        RECT 29.765 11.100 30.255 11.115 ;
        RECT 39.065 11.005 41.615 11.965 ;
        RECT 50.285 10.995 52.405 12.145 ;
        RECT 62.915 12.135 63.405 73.010 ;
        RECT 65.035 54.010 65.495 54.085 ;
        RECT 70.605 54.010 71.065 54.035 ;
        RECT 65.035 53.570 71.065 54.010 ;
        RECT 65.035 53.515 65.495 53.570 ;
        RECT 70.605 53.465 71.065 53.570 ;
        RECT 67.295 48.820 67.775 48.885 ;
        RECT 67.295 48.500 69.095 48.820 ;
        RECT 67.295 48.335 67.775 48.500 ;
        RECT 68.525 45.660 69.085 48.500 ;
        RECT 72.405 45.660 72.885 45.685 ;
        RECT 68.525 45.240 72.885 45.660 ;
        RECT 68.525 45.230 69.085 45.240 ;
        RECT 72.405 45.135 72.885 45.240 ;
        RECT 65.735 40.100 66.215 40.205 ;
        RECT 69.535 40.100 70.095 40.110 ;
        RECT 65.735 39.680 70.095 40.100 ;
        RECT 65.735 39.655 66.215 39.680 ;
        RECT 69.535 36.840 70.095 39.680 ;
        RECT 70.845 36.840 71.325 37.005 ;
        RECT 69.525 36.520 71.325 36.840 ;
        RECT 70.845 36.455 71.325 36.520 ;
        RECT 67.555 31.770 68.015 31.875 ;
        RECT 73.125 31.770 73.585 31.825 ;
        RECT 67.555 31.330 73.585 31.770 ;
        RECT 67.555 31.305 68.015 31.330 ;
        RECT 73.125 31.255 73.585 31.330 ;
        RECT 74.055 12.165 74.545 73.050 ;
        RECT 83.690 73.000 86.290 74.540 ;
        RECT 94.960 74.710 97.520 75.580 ;
        RECT 94.960 73.020 97.570 74.710 ;
        RECT 106.340 74.460 108.900 75.640 ;
        RECT 117.470 74.720 120.030 75.650 ;
        RECT 76.275 54.000 76.735 54.075 ;
        RECT 81.845 54.000 82.305 54.025 ;
        RECT 76.275 53.560 82.305 54.000 ;
        RECT 76.275 53.505 76.735 53.560 ;
        RECT 81.845 53.455 82.305 53.560 ;
        RECT 78.535 48.810 79.015 48.875 ;
        RECT 78.535 48.490 80.335 48.810 ;
        RECT 78.535 48.325 79.015 48.490 ;
        RECT 79.765 45.650 80.325 48.490 ;
        RECT 83.645 45.650 84.125 45.675 ;
        RECT 79.765 45.230 84.125 45.650 ;
        RECT 79.765 45.220 80.325 45.230 ;
        RECT 83.645 45.125 84.125 45.230 ;
        RECT 77.025 40.090 77.505 40.195 ;
        RECT 80.825 40.090 81.385 40.100 ;
        RECT 77.025 39.670 81.385 40.090 ;
        RECT 77.025 39.645 77.505 39.670 ;
        RECT 80.825 36.830 81.385 39.670 ;
        RECT 82.135 36.830 82.615 36.995 ;
        RECT 80.815 36.510 82.615 36.830 ;
        RECT 82.135 36.445 82.615 36.510 ;
        RECT 78.845 31.760 79.305 31.865 ;
        RECT 84.415 31.760 84.875 31.815 ;
        RECT 78.845 31.320 84.875 31.760 ;
        RECT 78.845 31.295 79.305 31.320 ;
        RECT 84.415 31.245 84.875 31.320 ;
        RECT 61.365 10.985 63.485 12.135 ;
        RECT 72.675 11.015 74.795 12.165 ;
        RECT 85.375 12.155 85.865 73.000 ;
        RECT 87.525 54.010 87.985 54.085 ;
        RECT 93.095 54.010 93.555 54.035 ;
        RECT 87.525 53.570 93.555 54.010 ;
        RECT 87.525 53.515 87.985 53.570 ;
        RECT 93.095 53.465 93.555 53.570 ;
        RECT 89.785 48.820 90.265 48.885 ;
        RECT 89.785 48.500 91.585 48.820 ;
        RECT 89.785 48.335 90.265 48.500 ;
        RECT 91.015 45.660 91.575 48.500 ;
        RECT 94.895 45.660 95.375 45.685 ;
        RECT 91.015 45.240 95.375 45.660 ;
        RECT 91.015 45.230 91.575 45.240 ;
        RECT 94.895 45.135 95.375 45.240 ;
        RECT 88.265 40.110 88.745 40.215 ;
        RECT 92.065 40.110 92.625 40.120 ;
        RECT 88.265 39.690 92.625 40.110 ;
        RECT 88.265 39.665 88.745 39.690 ;
        RECT 92.065 36.850 92.625 39.690 ;
        RECT 93.375 36.850 93.855 37.015 ;
        RECT 92.055 36.530 93.855 36.850 ;
        RECT 93.375 36.465 93.855 36.530 ;
        RECT 90.085 31.780 90.545 31.885 ;
        RECT 95.655 31.780 96.115 31.835 ;
        RECT 90.085 31.340 96.115 31.780 ;
        RECT 90.085 31.315 90.545 31.340 ;
        RECT 95.655 31.265 96.115 31.340 ;
        RECT 96.605 12.155 97.095 73.020 ;
        RECT 106.150 73.000 109.060 74.460 ;
        RECT 117.470 73.070 120.000 74.720 ;
        RECT 129.290 74.650 131.850 75.650 ;
        RECT 129.300 73.140 131.820 74.650 ;
        RECT 98.805 54.000 99.265 54.075 ;
        RECT 104.375 54.000 104.835 54.025 ;
        RECT 98.805 53.560 104.835 54.000 ;
        RECT 98.805 53.505 99.265 53.560 ;
        RECT 104.375 53.455 104.835 53.560 ;
        RECT 101.065 48.810 101.545 48.875 ;
        RECT 101.065 48.490 102.865 48.810 ;
        RECT 101.065 48.325 101.545 48.490 ;
        RECT 102.295 45.650 102.855 48.490 ;
        RECT 106.175 45.650 106.655 45.675 ;
        RECT 102.295 45.230 106.655 45.650 ;
        RECT 102.295 45.220 102.855 45.230 ;
        RECT 106.175 45.125 106.655 45.230 ;
        RECT 99.475 40.130 99.955 40.235 ;
        RECT 103.275 40.130 103.835 40.140 ;
        RECT 99.475 39.710 103.835 40.130 ;
        RECT 99.475 39.685 99.955 39.710 ;
        RECT 103.275 36.870 103.835 39.710 ;
        RECT 104.585 36.870 105.065 37.035 ;
        RECT 103.265 36.550 105.065 36.870 ;
        RECT 104.585 36.485 105.065 36.550 ;
        RECT 101.295 31.800 101.755 31.905 ;
        RECT 106.865 31.800 107.325 31.855 ;
        RECT 101.295 31.360 107.325 31.800 ;
        RECT 101.295 31.335 101.755 31.360 ;
        RECT 106.865 31.285 107.325 31.360 ;
        RECT 107.865 12.205 108.355 73.000 ;
        RECT 110.075 54.000 110.535 54.075 ;
        RECT 115.645 54.000 116.105 54.025 ;
        RECT 110.075 53.560 116.105 54.000 ;
        RECT 110.075 53.505 110.535 53.560 ;
        RECT 115.645 53.455 116.105 53.560 ;
        RECT 112.335 48.810 112.815 48.875 ;
        RECT 112.335 48.490 114.135 48.810 ;
        RECT 112.335 48.325 112.815 48.490 ;
        RECT 113.565 45.650 114.125 48.490 ;
        RECT 117.445 45.650 117.925 45.675 ;
        RECT 113.565 45.230 117.925 45.650 ;
        RECT 113.565 45.220 114.125 45.230 ;
        RECT 117.445 45.125 117.925 45.230 ;
        RECT 110.675 40.170 111.155 40.275 ;
        RECT 114.475 40.170 115.035 40.180 ;
        RECT 110.675 39.750 115.035 40.170 ;
        RECT 110.675 39.725 111.155 39.750 ;
        RECT 114.475 36.910 115.035 39.750 ;
        RECT 115.785 36.910 116.265 37.075 ;
        RECT 114.465 36.590 116.265 36.910 ;
        RECT 115.785 36.525 116.265 36.590 ;
        RECT 112.495 31.840 112.955 31.945 ;
        RECT 118.065 31.840 118.525 31.895 ;
        RECT 112.495 31.400 118.525 31.840 ;
        RECT 112.495 31.375 112.955 31.400 ;
        RECT 118.065 31.325 118.525 31.400 ;
        RECT 119.085 12.205 119.575 73.070 ;
        RECT 121.325 54.000 121.785 54.075 ;
        RECT 126.895 54.000 127.355 54.025 ;
        RECT 121.325 53.560 127.355 54.000 ;
        RECT 121.325 53.505 121.785 53.560 ;
        RECT 126.895 53.455 127.355 53.560 ;
        RECT 123.585 48.810 124.065 48.875 ;
        RECT 123.585 48.490 125.385 48.810 ;
        RECT 123.585 48.325 124.065 48.490 ;
        RECT 124.815 45.650 125.375 48.490 ;
        RECT 128.695 45.650 129.175 45.675 ;
        RECT 124.815 45.230 129.175 45.650 ;
        RECT 124.815 45.220 125.375 45.230 ;
        RECT 128.695 45.125 129.175 45.230 ;
        RECT 121.885 40.190 122.365 40.295 ;
        RECT 125.685 40.190 126.245 40.200 ;
        RECT 121.885 39.770 126.245 40.190 ;
        RECT 121.885 39.745 122.365 39.770 ;
        RECT 125.685 36.930 126.245 39.770 ;
        RECT 126.995 36.930 127.475 37.095 ;
        RECT 125.675 36.610 127.475 36.930 ;
        RECT 126.995 36.545 127.475 36.610 ;
        RECT 123.705 31.860 124.165 31.965 ;
        RECT 129.275 31.860 129.735 31.915 ;
        RECT 123.705 31.420 129.735 31.860 ;
        RECT 123.705 31.395 124.165 31.420 ;
        RECT 129.275 31.345 129.735 31.420 ;
        RECT 130.335 12.235 130.825 73.140 ;
        RECT 74.055 11.010 74.545 11.015 ;
        RECT 83.795 11.005 85.915 12.155 ;
        RECT 95.095 11.005 97.215 12.155 ;
        RECT 106.285 11.055 108.405 12.205 ;
        RECT 117.515 11.055 119.635 12.205 ;
        RECT 128.815 11.085 130.935 12.235 ;
        RECT 107.865 11.010 108.355 11.055 ;
        RECT 119.085 11.050 119.575 11.055 ;
        RECT 85.375 11.000 85.865 11.005 ;
        RECT 96.605 10.980 97.095 11.005 ;
        RECT 74.290 0.135 75.680 1.435 ;
        RECT 93.500 0.205 94.890 1.505 ;
        RECT 112.900 0.335 114.290 1.635 ;
        RECT 131.800 0.405 133.540 1.905 ;
        RECT 151.600 0.275 152.970 1.445 ;
      LAYER met4 ;
        RECT 30.420 225.130 30.670 225.140 ;
        RECT 30.300 224.760 30.670 225.130 ;
        RECT 30.970 224.760 33.430 225.140 ;
        RECT 33.730 224.760 36.190 225.140 ;
        RECT 36.490 224.760 38.950 225.140 ;
        RECT 39.250 224.760 41.710 225.140 ;
        RECT 42.010 224.760 44.470 225.140 ;
        RECT 44.770 224.760 47.230 225.140 ;
        RECT 47.530 224.760 49.990 225.140 ;
        RECT 50.290 224.760 52.750 225.140 ;
        RECT 53.050 224.760 55.510 225.140 ;
        RECT 55.810 224.760 58.270 225.140 ;
        RECT 58.570 224.760 61.030 225.140 ;
        RECT 61.330 224.760 63.790 225.140 ;
        RECT 64.090 224.760 66.550 225.140 ;
        RECT 66.850 224.760 69.310 225.140 ;
        RECT 69.610 224.760 72.070 225.140 ;
        RECT 72.370 224.760 74.830 225.140 ;
        RECT 75.130 224.760 77.590 225.140 ;
        RECT 77.890 224.760 80.350 225.140 ;
        RECT 80.650 224.760 83.110 225.140 ;
        RECT 83.410 224.760 85.870 225.140 ;
        RECT 86.170 224.760 88.630 225.140 ;
        RECT 88.930 224.760 91.390 225.140 ;
        RECT 91.690 224.760 94.150 225.140 ;
        RECT 94.450 224.760 96.910 225.140 ;
        RECT 97.210 224.760 99.670 225.140 ;
        RECT 99.970 224.760 102.430 225.140 ;
        RECT 102.730 224.760 105.190 225.140 ;
        RECT 105.490 224.760 107.950 225.140 ;
        RECT 108.250 224.760 110.710 225.140 ;
        RECT 111.010 224.760 113.470 225.140 ;
        RECT 113.770 224.760 116.230 225.140 ;
        RECT 116.530 224.760 118.990 225.140 ;
        RECT 119.290 224.760 121.750 225.140 ;
        RECT 122.050 224.760 124.510 225.140 ;
        RECT 124.810 224.760 127.270 225.140 ;
        RECT 127.570 224.760 130.030 225.140 ;
        RECT 130.330 224.760 132.790 225.140 ;
        RECT 133.090 224.760 133.520 225.140 ;
        RECT 30.300 224.240 133.520 224.760 ;
        RECT 135.385 224.760 135.550 225.185 ;
        RECT 135.850 224.760 136.745 225.185 ;
        RECT 30.300 219.100 31.660 224.240 ;
        RECT 135.385 223.875 136.745 224.760 ;
        RECT 138.175 224.760 138.310 225.115 ;
        RECT 138.610 224.760 139.535 225.115 ;
        RECT 138.175 223.805 139.535 224.760 ;
        RECT 143.225 224.760 143.830 225.145 ;
        RECT 144.130 224.760 144.585 225.145 ;
        RECT 143.225 223.835 144.585 224.760 ;
        RECT 6.000 218.040 31.660 219.100 ;
        RECT 30.300 217.960 31.660 218.040 ;
        RECT 16.820 99.530 18.820 211.530 ;
        RECT 31.820 99.530 33.820 211.530 ;
        RECT 46.820 99.530 48.820 211.530 ;
        RECT 61.820 99.530 63.820 211.530 ;
        RECT 64.635 174.065 64.965 174.395 ;
        RECT 64.650 149.235 64.950 174.065 ;
        RECT 64.635 148.905 64.965 149.235 ;
        RECT 64.650 122.715 64.950 148.905 ;
        RECT 75.675 146.185 76.005 146.515 ;
        RECT 75.690 139.035 75.990 146.185 ;
        RECT 75.675 138.705 76.005 139.035 ;
        RECT 64.635 122.385 64.965 122.715 ;
        RECT 76.820 99.530 78.820 211.530 ;
        RECT 81.195 176.105 81.525 176.435 ;
        RECT 80.275 143.465 80.605 143.795 ;
        RECT 80.290 111.835 80.590 143.465 ;
        RECT 81.210 132.235 81.510 176.105 ;
        RECT 81.195 131.905 81.525 132.235 ;
        RECT 80.275 111.505 80.605 111.835 ;
        RECT 91.820 99.530 93.820 211.530 ;
        RECT 106.820 99.530 108.820 211.530 ;
        RECT 121.820 99.720 123.820 211.530 ;
        RECT 118.110 97.700 120.130 99.670 ;
        RECT 121.810 97.750 123.830 99.720 ;
        RECT 118.130 93.980 120.130 97.700 ;
        RECT 121.820 96.830 123.820 97.750 ;
        RECT 121.820 94.830 139.410 96.830 ;
        RECT 118.130 91.980 135.580 93.980 ;
        RECT 133.580 77.835 135.580 91.980 ;
        RECT 133.375 76.625 136.015 77.835 ;
        RECT 137.410 77.815 139.410 94.830 ;
        RECT 137.235 76.605 139.875 77.815 ;
        RECT 3.955 71.365 4.000 73.195 ;
        RECT 6.000 71.365 6.055 73.195 ;
        RECT 3.000 68.705 3.025 70.435 ;
        RECT 15.555 68.655 16.995 71.165 ;
        RECT 74.335 1.000 75.635 1.415 ;
        RECT 74.335 0.155 74.530 1.000 ;
        RECT 75.430 0.155 75.635 1.000 ;
        RECT 93.545 1.000 94.845 1.485 ;
        RECT 93.545 0.225 93.850 1.000 ;
        RECT 94.750 0.225 94.845 1.000 ;
        RECT 112.945 1.000 114.245 1.615 ;
        RECT 112.945 0.355 113.170 1.000 ;
        RECT 114.070 0.355 114.245 1.000 ;
        RECT 131.845 1.000 133.495 1.885 ;
        RECT 131.845 0.425 132.490 1.000 ;
        RECT 133.390 0.425 133.495 1.000 ;
        RECT 151.645 1.000 152.925 1.425 ;
        RECT 151.645 0.295 151.810 1.000 ;
        RECT 152.710 0.295 152.925 1.000 ;
  END
END tt_um_08_sws
END LIBRARY

