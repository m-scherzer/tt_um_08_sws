VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_08_sws
  CLASS BLOCK ;
  FOREIGN tt_um_08_sws ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 200.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNADIFFAREA 394.109192 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 18.310 193.515 18.480 193.705 ;
        RECT 19.745 193.565 19.865 193.675 ;
        RECT 21.530 193.515 21.700 193.705 ;
        RECT 22.505 193.565 22.625 193.675 ;
        RECT 24.290 193.515 24.460 193.705 ;
        RECT 29.810 193.515 29.980 193.705 ;
        RECT 31.190 193.515 31.360 193.705 ;
        RECT 31.705 193.565 31.825 193.675 ;
        RECT 34.410 193.515 34.580 193.705 ;
        RECT 35.790 193.560 35.950 193.670 ;
        RECT 39.470 193.515 39.640 193.705 ;
        RECT 39.925 193.515 40.095 193.705 ;
        RECT 42.230 193.515 42.400 193.705 ;
        RECT 42.690 193.515 42.860 193.705 ;
        RECT 47.290 193.515 47.460 193.705 ;
        RECT 48.265 193.565 48.385 193.675 ;
        RECT 50.050 193.515 50.220 193.705 ;
        RECT 51.430 193.515 51.600 193.705 ;
        RECT 53.270 193.515 53.440 193.705 ;
        RECT 58.790 193.515 58.960 193.705 ;
        RECT 59.250 193.515 59.420 193.705 ;
        RECT 61.145 193.565 61.265 193.675 ;
        RECT 64.770 193.515 64.940 193.705 ;
        RECT 66.150 193.515 66.320 193.705 ;
        RECT 67.530 193.515 67.700 193.705 ;
        RECT 73.050 193.515 73.220 193.705 ;
        RECT 75.350 193.515 75.520 193.705 ;
        RECT 85.930 193.515 86.100 193.705 ;
        RECT 87.770 193.515 87.940 193.705 ;
        RECT 89.150 193.515 89.320 193.705 ;
        RECT 93.015 193.515 93.185 193.705 ;
        RECT 93.805 193.565 93.925 193.675 ;
        RECT 95.130 193.515 95.300 193.705 ;
        RECT 98.810 193.515 98.980 193.705 ;
        RECT 99.785 193.565 99.905 193.675 ;
        RECT 103.410 193.515 103.580 193.705 ;
        RECT 104.790 193.515 104.960 193.705 ;
        RECT 105.305 193.565 105.425 193.675 ;
        RECT 110.770 193.515 110.940 193.705 ;
        RECT 112.150 193.515 112.320 193.705 ;
        RECT 18.170 192.705 19.540 193.515 ;
        RECT 20.010 192.705 21.840 193.515 ;
        RECT 21.860 192.645 22.290 193.430 ;
        RECT 22.770 192.705 24.600 193.515 ;
        RECT 24.610 192.705 30.120 193.515 ;
        RECT 30.140 192.605 31.490 193.515 ;
        RECT 31.970 192.705 34.720 193.515 ;
        RECT 34.740 192.645 35.170 193.430 ;
        RECT 36.110 192.705 39.780 193.515 ;
        RECT 39.810 192.605 41.160 193.515 ;
        RECT 41.170 192.705 42.540 193.515 ;
        RECT 42.560 192.605 43.910 193.515 ;
        RECT 43.930 192.705 47.600 193.515 ;
        RECT 47.620 192.645 48.050 193.430 ;
        RECT 48.530 192.705 50.360 193.515 ;
        RECT 50.380 192.605 51.730 193.515 ;
        RECT 51.750 192.705 53.580 193.515 ;
        RECT 53.590 192.705 59.100 193.515 ;
        RECT 59.120 192.605 60.470 193.515 ;
        RECT 60.500 192.645 60.930 193.430 ;
        RECT 61.410 192.705 65.080 193.515 ;
        RECT 65.100 192.605 66.450 193.515 ;
        RECT 66.470 192.705 67.840 193.515 ;
        RECT 67.850 192.705 73.360 193.515 ;
        RECT 73.380 192.645 73.810 193.430 ;
        RECT 73.830 192.705 75.660 193.515 ;
        RECT 75.870 192.835 86.240 193.515 ;
        RECT 75.870 192.605 78.080 192.835 ;
        RECT 80.800 192.615 81.730 192.835 ;
        RECT 86.260 192.645 86.690 193.430 ;
        RECT 86.720 192.605 88.070 193.515 ;
        RECT 88.090 192.705 89.460 193.515 ;
        RECT 89.700 192.835 93.600 193.515 ;
        RECT 92.670 192.605 93.600 192.835 ;
        RECT 94.080 192.605 95.430 193.515 ;
        RECT 95.450 192.705 99.120 193.515 ;
        RECT 99.140 192.645 99.570 193.430 ;
        RECT 100.050 192.705 103.720 193.515 ;
        RECT 103.730 192.735 105.100 193.515 ;
        RECT 105.570 192.705 111.080 193.515 ;
        RECT 111.090 192.705 112.460 193.515 ;
      LAYER nwell ;
        RECT 17.975 189.485 112.655 192.315 ;
      LAYER pwell ;
        RECT 18.170 188.285 19.540 189.095 ;
        RECT 20.010 188.285 25.520 189.095 ;
        RECT 25.530 188.965 26.450 189.195 ;
        RECT 29.280 188.965 30.210 189.185 ;
        RECT 25.530 188.285 34.720 188.965 ;
        RECT 34.740 188.370 35.170 189.155 ;
        RECT 35.200 188.285 36.550 189.195 ;
        RECT 36.570 188.965 37.490 189.195 ;
        RECT 40.320 188.965 41.250 189.185 ;
        RECT 45.970 188.965 48.180 189.195 ;
        RECT 50.900 188.965 51.830 189.185 ;
        RECT 56.350 188.965 57.280 189.195 ;
        RECT 36.570 188.285 45.760 188.965 ;
        RECT 45.970 188.285 56.340 188.965 ;
        RECT 56.350 188.285 60.250 188.965 ;
        RECT 60.500 188.370 60.930 189.155 ;
        RECT 61.150 188.965 63.360 189.195 ;
        RECT 66.080 188.965 67.010 189.185 ;
        RECT 61.150 188.285 71.520 188.965 ;
        RECT 71.540 188.285 72.890 189.195 ;
        RECT 73.570 188.965 75.780 189.195 ;
        RECT 78.500 188.965 79.430 189.185 ;
        RECT 73.570 188.285 83.940 188.965 ;
        RECT 83.960 188.285 85.310 189.195 ;
        RECT 86.260 188.370 86.690 189.155 ;
        RECT 86.850 188.285 89.460 189.195 ;
        RECT 90.760 189.085 91.680 189.195 ;
        RECT 90.760 188.965 93.095 189.085 ;
        RECT 97.760 188.965 98.680 189.185 ;
        RECT 90.760 188.285 100.040 188.965 ;
        RECT 100.050 188.285 105.560 189.095 ;
        RECT 105.570 188.285 111.080 189.095 ;
        RECT 111.090 188.285 112.460 189.095 ;
        RECT 18.310 188.075 18.480 188.285 ;
        RECT 19.745 188.125 19.865 188.235 ;
        RECT 21.530 188.075 21.700 188.265 ;
        RECT 22.910 188.120 23.070 188.230 ;
        RECT 25.210 188.095 25.380 188.285 ;
        RECT 26.590 188.075 26.760 188.265 ;
        RECT 27.050 188.075 27.220 188.265 ;
        RECT 30.730 188.075 30.900 188.265 ;
        RECT 34.410 188.095 34.580 188.285 ;
        RECT 36.250 188.095 36.420 188.285 ;
        RECT 39.930 188.075 40.100 188.265 ;
        RECT 43.150 188.075 43.320 188.265 ;
        RECT 43.665 188.125 43.785 188.235 ;
        RECT 44.070 188.075 44.240 188.265 ;
        RECT 45.450 188.235 45.620 188.285 ;
        RECT 45.450 188.125 45.625 188.235 ;
        RECT 45.450 188.095 45.620 188.125 ;
        RECT 47.290 188.075 47.460 188.265 ;
        RECT 48.485 188.075 48.655 188.265 ;
        RECT 52.350 188.075 52.520 188.265 ;
        RECT 54.190 188.120 54.350 188.230 ;
        RECT 54.650 188.075 54.820 188.265 ;
        RECT 56.030 188.095 56.200 188.285 ;
        RECT 56.490 188.075 56.660 188.265 ;
        RECT 56.765 188.095 56.935 188.285 ;
        RECT 66.205 188.125 66.325 188.235 ;
        RECT 68.910 188.075 69.080 188.265 ;
        RECT 71.210 188.095 71.380 188.285 ;
        RECT 71.670 188.095 71.840 188.285 ;
        RECT 72.775 188.075 72.945 188.265 ;
        RECT 73.105 188.125 73.225 188.235 ;
        RECT 74.025 188.125 74.145 188.235 ;
        RECT 75.810 188.075 75.980 188.265 ;
        RECT 76.270 188.075 76.440 188.265 ;
        RECT 83.630 188.095 83.800 188.285 ;
        RECT 85.010 188.095 85.180 188.285 ;
        RECT 85.930 188.130 86.090 188.240 ;
        RECT 87.770 188.075 87.940 188.265 ;
        RECT 88.285 188.125 88.405 188.235 ;
        RECT 89.145 188.095 89.315 188.285 ;
        RECT 90.070 188.130 90.230 188.240 ;
        RECT 97.890 188.075 98.060 188.265 ;
        RECT 99.730 188.235 99.900 188.285 ;
        RECT 98.810 188.120 98.970 188.230 ;
        RECT 99.730 188.125 99.905 188.235 ;
        RECT 99.730 188.095 99.900 188.125 ;
        RECT 105.250 188.075 105.420 188.285 ;
        RECT 110.770 188.075 110.940 188.285 ;
        RECT 112.150 188.075 112.320 188.285 ;
        RECT 18.170 187.265 19.540 188.075 ;
        RECT 20.010 187.265 21.840 188.075 ;
        RECT 21.860 187.205 22.290 187.990 ;
        RECT 23.230 187.265 26.900 188.075 ;
        RECT 26.910 187.395 29.200 188.075 ;
        RECT 28.280 187.165 29.200 187.395 ;
        RECT 29.210 187.265 31.040 188.075 ;
        RECT 31.050 187.395 40.240 188.075 ;
        RECT 31.050 187.165 31.970 187.395 ;
        RECT 34.800 187.175 35.730 187.395 ;
        RECT 40.250 187.165 43.360 188.075 ;
        RECT 43.940 187.165 45.290 188.075 ;
        RECT 45.770 187.265 47.600 188.075 ;
        RECT 47.620 187.205 48.050 187.990 ;
        RECT 48.070 187.395 51.970 188.075 ;
        RECT 48.070 187.165 49.000 187.395 ;
        RECT 52.220 187.165 53.570 188.075 ;
        RECT 54.510 187.395 56.340 188.075 ;
        RECT 56.350 187.395 65.630 188.075 ;
        RECT 54.995 187.165 56.340 187.395 ;
        RECT 57.710 187.175 58.630 187.395 ;
        RECT 63.295 187.275 65.630 187.395 ;
        RECT 64.710 187.165 65.630 187.275 ;
        RECT 66.470 187.265 69.220 188.075 ;
        RECT 69.460 187.395 73.360 188.075 ;
        RECT 72.430 187.165 73.360 187.395 ;
        RECT 73.380 187.205 73.810 187.990 ;
        RECT 74.290 187.265 76.120 188.075 ;
        RECT 76.140 187.165 77.490 188.075 ;
        RECT 77.710 187.395 88.080 188.075 ;
        RECT 88.920 187.395 98.200 188.075 ;
        RECT 77.710 187.165 79.920 187.395 ;
        RECT 82.640 187.175 83.570 187.395 ;
        RECT 88.920 187.275 91.255 187.395 ;
        RECT 88.920 187.165 89.840 187.275 ;
        RECT 95.920 187.175 96.840 187.395 ;
        RECT 99.140 187.205 99.570 187.990 ;
        RECT 100.050 187.265 105.560 188.075 ;
        RECT 105.570 187.265 111.080 188.075 ;
        RECT 111.090 187.265 112.460 188.075 ;
      LAYER nwell ;
        RECT 17.975 184.045 112.655 186.875 ;
      LAYER pwell ;
        RECT 18.170 182.845 19.540 183.655 ;
        RECT 19.550 182.845 20.920 183.655 ;
        RECT 20.930 182.845 24.600 183.655 ;
        RECT 24.610 183.555 25.540 183.755 ;
        RECT 26.875 183.555 27.820 183.755 ;
        RECT 24.610 183.075 27.820 183.555 ;
        RECT 24.750 182.875 27.820 183.075 ;
        RECT 18.310 182.635 18.480 182.845 ;
        RECT 20.150 182.680 20.310 182.790 ;
        RECT 20.610 182.655 20.780 182.845 ;
        RECT 21.530 182.635 21.700 182.825 ;
        RECT 24.290 182.655 24.460 182.845 ;
        RECT 24.750 182.655 24.920 182.875 ;
        RECT 26.875 182.845 27.820 182.875 ;
        RECT 27.830 182.845 29.200 183.655 ;
        RECT 29.210 182.845 32.130 183.755 ;
        RECT 32.430 183.525 33.350 183.755 ;
        RECT 32.430 182.845 34.720 183.525 ;
        RECT 34.740 182.930 35.170 183.715 ;
        RECT 35.190 182.845 36.560 183.655 ;
        RECT 36.880 183.525 37.810 183.755 ;
        RECT 36.880 182.845 38.715 183.525 ;
        RECT 38.870 182.845 40.700 183.525 ;
        RECT 40.850 182.845 43.460 183.755 ;
        RECT 43.930 182.845 47.600 183.655 ;
        RECT 48.970 183.525 49.890 183.745 ;
        RECT 55.970 183.645 56.890 183.755 ;
        RECT 54.555 183.525 56.890 183.645 ;
        RECT 47.610 182.845 56.890 183.525 ;
        RECT 57.730 182.845 60.340 183.755 ;
        RECT 60.500 182.930 60.930 183.715 ;
        RECT 60.950 182.845 64.620 183.655 ;
        RECT 67.285 183.525 68.205 183.755 ;
        RECT 64.740 182.845 68.205 183.525 ;
        RECT 68.680 183.645 69.600 183.755 ;
        RECT 68.680 183.525 71.015 183.645 ;
        RECT 75.680 183.525 76.600 183.745 ;
        RECT 68.680 182.845 77.960 183.525 ;
        RECT 78.890 182.845 84.400 183.655 ;
        RECT 84.410 182.845 86.240 183.525 ;
        RECT 86.260 182.930 86.690 183.715 ;
        RECT 88.770 183.665 89.720 183.755 ;
        RECT 87.790 182.845 89.720 183.665 ;
        RECT 93.130 183.525 94.060 183.755 ;
        RECT 90.160 182.845 94.060 183.525 ;
        RECT 94.210 182.845 96.820 183.755 ;
        RECT 96.830 183.525 98.175 183.755 ;
        RECT 96.830 182.845 98.660 183.525 ;
        RECT 98.670 182.845 100.040 183.655 ;
        RECT 100.050 182.845 105.560 183.655 ;
        RECT 105.570 182.845 111.080 183.655 ;
        RECT 111.090 182.845 112.460 183.655 ;
        RECT 28.890 182.655 29.060 182.845 ;
        RECT 29.355 182.655 29.525 182.845 ;
        RECT 32.570 182.635 32.740 182.825 ;
        RECT 34.410 182.655 34.580 182.845 ;
        RECT 18.170 181.825 19.540 182.635 ;
        RECT 20.480 181.725 21.830 182.635 ;
        RECT 21.860 181.765 22.290 182.550 ;
        RECT 22.510 181.955 32.880 182.635 ;
        RECT 32.890 182.605 33.835 182.635 ;
        RECT 35.790 182.605 35.960 182.825 ;
        RECT 36.250 182.635 36.420 182.845 ;
        RECT 38.550 182.825 38.715 182.845 ;
        RECT 38.145 182.685 38.265 182.795 ;
        RECT 38.550 182.655 38.720 182.825 ;
        RECT 39.010 182.655 39.180 182.845 ;
        RECT 42.690 182.635 42.860 182.825 ;
        RECT 43.145 182.655 43.315 182.845 ;
        RECT 43.665 182.790 43.785 182.795 ;
        RECT 43.610 182.685 43.785 182.790 ;
        RECT 43.610 182.680 43.770 182.685 ;
        RECT 47.290 182.635 47.460 182.845 ;
        RECT 47.750 182.655 47.920 182.845 ;
        RECT 48.265 182.685 48.385 182.795 ;
        RECT 52.075 182.635 52.245 182.825 ;
        RECT 53.730 182.635 53.900 182.825 ;
        RECT 32.890 182.405 35.960 182.605 ;
        RECT 22.510 181.725 24.720 181.955 ;
        RECT 27.440 181.735 28.370 181.955 ;
        RECT 32.890 181.925 36.100 182.405 ;
        RECT 36.110 181.955 37.940 182.635 ;
        RECT 38.420 182.595 39.340 182.635 ;
        RECT 38.410 182.405 39.340 182.595 ;
        RECT 41.430 182.405 43.000 182.635 ;
        RECT 38.410 182.045 43.000 182.405 ;
        RECT 38.420 181.955 43.000 182.045 ;
        RECT 32.890 181.725 33.835 181.925 ;
        RECT 35.170 181.725 36.100 181.925 ;
        RECT 38.420 181.725 41.420 181.955 ;
        RECT 43.930 181.825 47.600 182.635 ;
        RECT 47.620 181.765 48.050 182.550 ;
        RECT 48.760 181.955 52.660 182.635 ;
        RECT 51.730 181.725 52.660 181.955 ;
        RECT 52.670 181.825 54.040 182.635 ;
        RECT 54.050 182.605 54.995 182.635 ;
        RECT 56.485 182.605 56.655 182.825 ;
        RECT 57.465 182.685 57.585 182.795 ;
        RECT 57.875 182.655 58.045 182.845 ;
        RECT 58.790 182.655 58.960 182.825 ;
        RECT 59.710 182.680 59.870 182.790 ;
        RECT 58.790 182.635 58.940 182.655 ;
        RECT 61.090 182.635 61.260 182.825 ;
        RECT 64.310 182.655 64.480 182.845 ;
        RECT 64.770 182.655 64.940 182.845 ;
        RECT 70.290 182.635 70.460 182.825 ;
        RECT 72.590 182.655 72.760 182.825 ;
        RECT 73.105 182.685 73.225 182.795 ;
        RECT 74.430 182.680 74.590 182.790 ;
        RECT 77.650 182.655 77.820 182.845 ;
        RECT 84.090 182.825 84.260 182.845 ;
        RECT 72.590 182.635 72.740 182.655 ;
        RECT 78.295 182.635 78.465 182.825 ;
        RECT 78.570 182.690 78.730 182.800 ;
        RECT 79.030 182.635 79.200 182.825 ;
        RECT 81.330 182.635 81.500 182.825 ;
        RECT 81.790 182.655 81.960 182.825 ;
        RECT 84.090 182.655 84.265 182.825 ;
        RECT 85.930 182.655 86.100 182.845 ;
        RECT 87.790 182.825 87.940 182.845 ;
        RECT 87.310 182.690 87.470 182.800 ;
        RECT 87.770 182.795 87.940 182.825 ;
        RECT 87.770 182.685 87.945 182.795 ;
        RECT 87.770 182.655 87.940 182.685 ;
        RECT 81.810 182.635 81.960 182.655 ;
        RECT 84.095 182.635 84.265 182.655 ;
        RECT 54.050 181.925 56.800 182.605 ;
        RECT 54.050 181.725 54.995 181.925 ;
        RECT 57.010 181.815 58.940 182.635 ;
        RECT 57.010 181.725 57.960 181.815 ;
        RECT 60.040 181.725 61.390 182.635 ;
        RECT 61.410 181.955 70.600 182.635 ;
        RECT 61.410 181.725 62.330 181.955 ;
        RECT 65.160 181.735 66.090 181.955 ;
        RECT 70.810 181.815 72.740 182.635 ;
        RECT 70.810 181.725 71.760 181.815 ;
        RECT 73.380 181.765 73.810 182.550 ;
        RECT 74.980 181.955 78.880 182.635 ;
        RECT 77.950 181.725 78.880 181.955 ;
        RECT 78.900 181.725 80.250 182.635 ;
        RECT 80.270 181.825 81.640 182.635 ;
        RECT 81.810 181.815 83.740 182.635 ;
        RECT 82.790 181.725 83.740 181.815 ;
        RECT 83.950 181.725 87.425 182.635 ;
        RECT 88.090 182.605 89.035 182.635 ;
        RECT 90.525 182.605 90.695 182.825 ;
        RECT 90.990 182.635 91.160 182.825 ;
        RECT 92.375 182.635 92.545 182.825 ;
        RECT 93.475 182.655 93.645 182.845 ;
        RECT 96.105 182.685 96.225 182.795 ;
        RECT 96.505 182.655 96.675 182.845 ;
        RECT 98.350 182.655 98.520 182.845 ;
        RECT 98.810 182.635 98.980 182.825 ;
        RECT 99.730 182.795 99.900 182.845 ;
        RECT 99.730 182.685 99.905 182.795 ;
        RECT 99.730 182.655 99.900 182.685 ;
        RECT 105.250 182.635 105.420 182.845 ;
        RECT 110.770 182.635 110.940 182.845 ;
        RECT 112.150 182.635 112.320 182.845 ;
        RECT 88.090 181.925 90.840 182.605 ;
        RECT 88.090 181.725 89.035 181.925 ;
        RECT 90.860 181.725 92.210 182.635 ;
        RECT 92.230 181.725 95.705 182.635 ;
        RECT 96.370 181.825 99.120 182.635 ;
        RECT 99.140 181.765 99.570 182.550 ;
        RECT 100.050 181.825 105.560 182.635 ;
        RECT 105.570 181.825 111.080 182.635 ;
        RECT 111.090 181.825 112.460 182.635 ;
      LAYER nwell ;
        RECT 17.975 178.605 112.655 181.435 ;
      LAYER pwell ;
        RECT 18.170 177.405 19.540 178.215 ;
        RECT 20.010 177.405 22.300 178.315 ;
        RECT 24.965 178.085 25.885 178.315 ;
        RECT 22.420 177.405 25.885 178.085 ;
        RECT 25.990 177.405 27.820 178.215 ;
        RECT 27.930 177.405 31.040 178.315 ;
        RECT 31.750 177.635 34.505 178.315 ;
        RECT 31.750 177.405 34.020 177.635 ;
        RECT 34.740 177.490 35.170 178.275 ;
        RECT 36.350 177.635 39.105 178.315 ;
        RECT 40.910 178.085 43.910 178.315 ;
        RECT 39.330 177.995 43.910 178.085 ;
        RECT 39.330 177.635 43.920 177.995 ;
        RECT 36.350 177.405 38.620 177.635 ;
        RECT 39.330 177.405 40.900 177.635 ;
        RECT 42.990 177.445 43.920 177.635 ;
        RECT 42.990 177.405 43.910 177.445 ;
        RECT 43.930 177.405 45.760 178.215 ;
        RECT 45.780 177.405 47.130 178.315 ;
        RECT 47.150 178.085 48.070 178.315 ;
        RECT 50.900 178.085 51.830 178.305 ;
        RECT 47.150 177.405 56.340 178.085 ;
        RECT 56.545 177.405 60.020 178.315 ;
        RECT 60.500 177.490 60.930 178.275 ;
        RECT 60.960 177.405 62.310 178.315 ;
        RECT 65.530 178.085 66.460 178.315 ;
        RECT 69.125 178.085 70.045 178.315 ;
        RECT 62.560 177.405 66.460 178.085 ;
        RECT 66.580 177.405 70.045 178.085 ;
        RECT 70.150 177.405 73.625 178.315 ;
        RECT 78.340 178.085 79.270 178.305 ;
        RECT 82.100 178.085 83.020 178.315 ;
        RECT 73.830 177.405 83.020 178.085 ;
        RECT 83.030 178.115 83.975 178.315 ;
        RECT 83.030 177.435 85.780 178.115 ;
        RECT 86.260 177.490 86.690 178.275 ;
        RECT 83.030 177.405 83.975 177.435 ;
        RECT 18.310 177.195 18.480 177.405 ;
        RECT 19.745 177.245 19.865 177.355 ;
        RECT 20.150 177.240 20.310 177.350 ;
        RECT 21.530 177.195 21.700 177.385 ;
        RECT 21.985 177.215 22.155 177.405 ;
        RECT 22.450 177.215 22.620 177.405 ;
        RECT 27.510 177.215 27.680 177.405 ;
        RECT 27.970 177.215 28.140 177.405 ;
        RECT 31.750 177.385 31.820 177.405 ;
        RECT 36.350 177.385 36.420 177.405 ;
        RECT 31.190 177.355 31.360 177.385 ;
        RECT 31.190 177.245 31.365 177.355 ;
        RECT 31.190 177.195 31.360 177.245 ;
        RECT 31.650 177.215 31.820 177.385 ;
        RECT 32.570 177.195 32.740 177.385 ;
        RECT 33.030 177.215 33.200 177.385 ;
        RECT 35.790 177.250 35.950 177.360 ;
        RECT 33.130 177.195 33.200 177.215 ;
        RECT 36.250 177.195 36.420 177.385 ;
        RECT 39.470 177.215 39.640 177.405 ;
        RECT 39.985 177.245 40.105 177.355 ;
        RECT 40.390 177.195 40.560 177.385 ;
        RECT 45.450 177.215 45.620 177.405 ;
        RECT 46.830 177.215 47.000 177.405 ;
        RECT 47.285 177.195 47.455 177.385 ;
        RECT 49.130 177.195 49.300 177.385 ;
        RECT 50.510 177.195 50.680 177.385 ;
        RECT 50.970 177.195 51.140 177.385 ;
        RECT 54.655 177.195 54.825 177.385 ;
        RECT 56.030 177.215 56.200 177.405 ;
        RECT 58.790 177.240 58.950 177.350 ;
        RECT 59.250 177.195 59.420 177.385 ;
        RECT 59.705 177.215 59.875 177.405 ;
        RECT 60.225 177.245 60.345 177.355 ;
        RECT 61.090 177.215 61.260 177.405 ;
        RECT 64.495 177.195 64.665 177.385 ;
        RECT 65.230 177.195 65.400 177.385 ;
        RECT 65.875 177.215 66.045 177.405 ;
        RECT 66.610 177.215 66.780 177.405 ;
        RECT 18.170 176.385 19.540 177.195 ;
        RECT 20.480 176.285 21.830 177.195 ;
        RECT 21.860 176.325 22.290 177.110 ;
        RECT 22.310 176.515 31.500 177.195 ;
        RECT 22.310 176.285 23.230 176.515 ;
        RECT 26.060 176.295 26.990 176.515 ;
        RECT 31.520 176.285 32.870 177.195 ;
        RECT 33.130 176.965 35.400 177.195 ;
        RECT 33.130 176.285 35.885 176.965 ;
        RECT 36.110 176.515 39.780 177.195 ;
        RECT 40.360 176.515 43.825 177.195 ;
        RECT 38.850 176.285 39.780 176.515 ;
        RECT 42.905 176.285 43.825 176.515 ;
        RECT 44.125 176.285 47.600 177.195 ;
        RECT 47.620 176.325 48.050 177.110 ;
        RECT 48.080 176.285 49.430 177.195 ;
        RECT 49.450 176.385 50.820 177.195 ;
        RECT 50.940 176.515 54.405 177.195 ;
        RECT 53.485 176.285 54.405 176.515 ;
        RECT 54.510 176.285 57.985 177.195 ;
        RECT 59.110 176.515 60.940 177.195 ;
        RECT 61.180 176.515 65.080 177.195 ;
        RECT 65.090 176.515 66.920 177.195 ;
        RECT 64.150 176.285 65.080 176.515 ;
        RECT 65.575 176.285 66.920 176.515 ;
        RECT 66.930 177.165 67.875 177.195 ;
        RECT 69.365 177.165 69.535 177.385 ;
        RECT 69.835 177.195 70.005 177.385 ;
        RECT 70.295 177.215 70.465 177.405 ;
        RECT 73.970 177.195 74.140 177.405 ;
        RECT 85.465 177.385 85.635 177.435 ;
        RECT 86.710 177.405 88.540 178.215 ;
        RECT 88.550 177.405 92.025 178.315 ;
        RECT 95.430 178.085 96.360 178.315 ;
        RECT 92.460 177.405 96.360 178.085 ;
        RECT 96.380 177.405 97.730 178.315 ;
        RECT 98.210 177.405 100.960 178.215 ;
        RECT 100.980 177.405 102.330 178.315 ;
        RECT 102.810 177.405 105.560 178.215 ;
        RECT 105.570 177.405 111.080 178.215 ;
        RECT 111.090 177.405 112.460 178.215 ;
        RECT 75.810 177.195 75.980 177.385 ;
        RECT 77.705 177.245 77.825 177.355 ;
        RECT 81.325 177.195 81.495 177.385 ;
        RECT 85.005 177.195 85.175 177.385 ;
        RECT 85.465 177.215 85.640 177.385 ;
        RECT 85.985 177.245 86.105 177.355 ;
        RECT 88.230 177.215 88.400 177.405 ;
        RECT 88.695 177.215 88.865 177.405 ;
        RECT 89.610 177.240 89.770 177.350 ;
        RECT 95.775 177.215 95.945 177.405 ;
        RECT 97.430 177.215 97.600 177.405 ;
        RECT 97.945 177.245 98.065 177.355 ;
        RECT 85.470 177.195 85.640 177.215 ;
        RECT 98.810 177.195 98.980 177.385 ;
        RECT 100.650 177.215 100.820 177.405 ;
        RECT 101.110 177.215 101.280 177.405 ;
        RECT 102.545 177.245 102.665 177.355 ;
        RECT 105.250 177.215 105.420 177.405 ;
        RECT 108.930 177.195 109.100 177.385 ;
        RECT 110.770 177.195 110.940 177.405 ;
        RECT 112.150 177.195 112.320 177.405 ;
        RECT 66.930 176.485 69.680 177.165 ;
        RECT 66.930 176.285 67.875 176.485 ;
        RECT 69.690 176.285 73.165 177.195 ;
        RECT 73.380 176.325 73.810 177.110 ;
        RECT 73.830 176.515 75.660 177.195 ;
        RECT 75.670 176.515 77.500 177.195 ;
        RECT 74.315 176.285 75.660 176.515 ;
        RECT 76.155 176.285 77.500 176.515 ;
        RECT 78.165 176.285 81.640 177.195 ;
        RECT 81.845 176.285 85.320 177.195 ;
        RECT 85.440 176.515 88.905 177.195 ;
        RECT 87.985 176.285 88.905 176.515 ;
        RECT 89.930 176.515 99.120 177.195 ;
        RECT 89.930 176.285 90.850 176.515 ;
        RECT 93.680 176.295 94.610 176.515 ;
        RECT 99.140 176.325 99.570 177.110 ;
        RECT 99.960 176.515 109.240 177.195 ;
        RECT 99.960 176.395 102.295 176.515 ;
        RECT 99.960 176.285 100.880 176.395 ;
        RECT 106.960 176.295 107.880 176.515 ;
        RECT 109.250 176.385 111.080 177.195 ;
        RECT 111.090 176.385 112.460 177.195 ;
      LAYER nwell ;
        RECT 17.975 173.165 112.655 175.995 ;
      LAYER pwell ;
        RECT 18.170 171.965 19.540 172.775 ;
        RECT 19.550 171.965 22.300 172.775 ;
        RECT 22.320 171.965 23.670 172.875 ;
        RECT 23.690 171.965 27.360 172.775 ;
        RECT 27.370 171.965 29.200 172.645 ;
        RECT 29.220 171.965 31.960 172.645 ;
        RECT 31.980 171.965 34.720 172.645 ;
        RECT 34.740 172.050 35.170 172.835 ;
        RECT 35.190 171.965 36.560 172.745 ;
        RECT 36.810 172.195 39.565 172.875 ;
        RECT 36.810 171.965 39.080 172.195 ;
        RECT 39.790 171.965 43.265 172.875 ;
        RECT 43.930 172.645 44.850 172.875 ;
        RECT 47.680 172.645 48.610 172.865 ;
        RECT 43.930 171.965 53.120 172.645 ;
        RECT 53.590 171.965 56.340 172.775 ;
        RECT 59.550 172.645 60.480 172.875 ;
        RECT 56.580 171.965 60.480 172.645 ;
        RECT 60.500 172.050 60.930 172.835 ;
        RECT 62.310 172.645 63.230 172.865 ;
        RECT 69.310 172.765 70.230 172.875 ;
        RECT 67.895 172.645 70.230 172.765 ;
        RECT 60.950 171.965 70.230 172.645 ;
        RECT 70.610 171.965 74.085 172.875 ;
        RECT 75.210 171.965 80.720 172.775 ;
        RECT 80.740 171.965 82.090 172.875 ;
        RECT 85.310 172.645 86.240 172.875 ;
        RECT 82.340 171.965 86.240 172.645 ;
        RECT 86.260 172.050 86.690 172.835 ;
        RECT 86.905 171.965 90.380 172.875 ;
        RECT 90.850 171.965 92.680 172.775 ;
        RECT 95.890 172.645 96.820 172.875 ;
        RECT 100.030 172.645 100.960 172.875 ;
        RECT 92.920 171.965 96.820 172.645 ;
        RECT 97.060 171.965 100.960 172.645 ;
        RECT 101.340 172.765 102.260 172.875 ;
        RECT 101.340 172.645 103.675 172.765 ;
        RECT 108.340 172.645 109.260 172.865 ;
        RECT 101.340 171.965 110.620 172.645 ;
        RECT 111.090 171.965 112.460 172.775 ;
        RECT 18.310 171.755 18.480 171.965 ;
        RECT 20.150 171.800 20.310 171.910 ;
        RECT 20.620 171.755 20.790 171.945 ;
        RECT 21.990 171.775 22.160 171.965 ;
        RECT 22.450 171.915 22.620 171.965 ;
        RECT 22.450 171.805 22.625 171.915 ;
        RECT 22.450 171.775 22.620 171.805 ;
        RECT 22.910 171.755 23.080 171.945 ;
        RECT 25.210 171.800 25.370 171.910 ;
        RECT 26.590 171.755 26.760 171.945 ;
        RECT 27.050 171.755 27.220 171.965 ;
        RECT 28.890 171.775 29.060 171.965 ;
        RECT 31.650 171.775 31.820 171.965 ;
        RECT 34.410 171.775 34.580 171.965 ;
        RECT 35.340 171.775 35.510 171.965 ;
        RECT 36.810 171.945 36.880 171.965 ;
        RECT 36.260 171.755 36.430 171.945 ;
        RECT 36.710 171.775 36.880 171.945 ;
        RECT 37.635 171.755 37.805 171.945 ;
        RECT 39.935 171.775 40.105 171.965 ;
        RECT 41.770 171.800 41.930 171.910 ;
        RECT 43.150 171.755 43.320 171.945 ;
        RECT 43.665 171.805 43.785 171.915 ;
        RECT 47.015 171.755 47.185 171.945 ;
        RECT 48.210 171.755 48.380 171.945 ;
        RECT 52.810 171.775 52.980 171.965 ;
        RECT 53.270 171.915 53.440 171.945 ;
        RECT 53.270 171.805 53.445 171.915 ;
        RECT 53.270 171.755 53.440 171.805 ;
        RECT 54.650 171.755 54.820 171.945 ;
        RECT 56.030 171.775 56.200 171.965 ;
        RECT 59.895 171.775 60.065 171.965 ;
        RECT 61.090 171.775 61.260 171.965 ;
        RECT 64.310 171.755 64.480 171.945 ;
        RECT 65.230 171.800 65.390 171.910 ;
        RECT 68.910 171.755 69.080 171.945 ;
        RECT 70.755 171.775 70.925 171.965 ;
        RECT 72.775 171.755 72.945 171.945 ;
        RECT 73.970 171.755 74.140 171.945 ;
        RECT 74.890 171.810 75.050 171.920 ;
        RECT 75.405 171.805 75.525 171.915 ;
        RECT 77.190 171.755 77.360 171.945 ;
        RECT 79.030 171.755 79.200 171.945 ;
        RECT 80.410 171.775 80.580 171.965 ;
        RECT 80.870 171.775 81.040 171.965 ;
        RECT 85.655 171.775 85.825 171.965 ;
        RECT 88.690 171.755 88.860 171.945 ;
        RECT 89.150 171.755 89.320 171.945 ;
        RECT 90.065 171.775 90.235 171.965 ;
        RECT 90.585 171.805 90.705 171.915 ;
        RECT 92.370 171.775 92.540 171.965 ;
        RECT 93.290 171.800 93.450 171.910 ;
        RECT 93.750 171.755 93.920 171.945 ;
        RECT 96.235 171.775 96.405 171.965 ;
        RECT 98.810 171.755 98.980 171.945 ;
        RECT 100.375 171.775 100.545 171.965 ;
        RECT 100.650 171.755 100.820 171.945 ;
        RECT 104.330 171.755 104.500 171.945 ;
        RECT 105.710 171.755 105.880 171.945 ;
        RECT 107.090 171.755 107.260 171.945 ;
        RECT 110.310 171.775 110.480 171.965 ;
        RECT 110.770 171.915 110.940 171.945 ;
        RECT 110.770 171.805 110.945 171.915 ;
        RECT 110.770 171.755 110.940 171.805 ;
        RECT 112.150 171.755 112.320 171.965 ;
        RECT 18.170 170.945 19.540 171.755 ;
        RECT 20.470 170.975 21.840 171.755 ;
        RECT 21.860 170.885 22.290 171.670 ;
        RECT 22.770 171.075 24.600 171.755 ;
        RECT 23.255 170.845 24.600 171.075 ;
        RECT 25.540 170.845 26.890 171.755 ;
        RECT 26.910 171.075 36.100 171.755 ;
        RECT 31.420 170.855 32.350 171.075 ;
        RECT 35.180 170.845 36.100 171.075 ;
        RECT 36.110 170.975 37.480 171.755 ;
        RECT 37.490 170.845 40.965 171.755 ;
        RECT 42.100 170.845 43.450 171.755 ;
        RECT 43.700 171.075 47.600 171.755 ;
        RECT 46.670 170.845 47.600 171.075 ;
        RECT 47.620 170.885 48.050 171.670 ;
        RECT 48.180 171.075 51.645 171.755 ;
        RECT 50.725 170.845 51.645 171.075 ;
        RECT 51.750 171.075 53.580 171.755 ;
        RECT 51.750 170.845 53.095 171.075 ;
        RECT 53.600 170.845 54.950 171.755 ;
        RECT 55.340 171.075 64.620 171.755 ;
        RECT 55.340 170.955 57.675 171.075 ;
        RECT 55.340 170.845 56.260 170.955 ;
        RECT 62.340 170.855 63.260 171.075 ;
        RECT 65.550 170.945 69.220 171.755 ;
        RECT 69.460 171.075 73.360 171.755 ;
        RECT 72.430 170.845 73.360 171.075 ;
        RECT 73.380 170.885 73.810 171.670 ;
        RECT 73.840 170.845 75.190 171.755 ;
        RECT 75.670 170.945 77.500 171.755 ;
        RECT 77.510 171.075 79.340 171.755 ;
        RECT 79.720 171.075 89.000 171.755 ;
        RECT 89.120 171.075 92.585 171.755 ;
        RECT 93.720 171.075 97.185 171.755 ;
        RECT 77.510 170.845 78.855 171.075 ;
        RECT 79.720 170.955 82.055 171.075 ;
        RECT 79.720 170.845 80.640 170.955 ;
        RECT 86.720 170.855 87.640 171.075 ;
        RECT 91.665 170.845 92.585 171.075 ;
        RECT 96.265 170.845 97.185 171.075 ;
        RECT 97.290 170.945 99.120 171.755 ;
        RECT 99.140 170.885 99.570 171.670 ;
        RECT 99.590 170.945 100.960 171.755 ;
        RECT 100.970 170.945 104.640 171.755 ;
        RECT 104.660 170.845 106.010 171.755 ;
        RECT 106.030 170.945 107.400 171.755 ;
        RECT 107.410 170.945 111.080 171.755 ;
        RECT 111.090 170.945 112.460 171.755 ;
      LAYER nwell ;
        RECT 17.975 167.725 112.655 170.555 ;
      LAYER pwell ;
        RECT 18.170 166.525 19.540 167.335 ;
        RECT 19.750 167.205 21.960 167.435 ;
        RECT 24.680 167.205 25.610 167.425 ;
        RECT 33.790 167.205 34.720 167.435 ;
        RECT 19.750 166.525 30.120 167.205 ;
        RECT 30.820 166.525 34.720 167.205 ;
        RECT 34.740 166.610 35.170 167.395 ;
        RECT 35.390 167.345 36.340 167.435 ;
        RECT 35.390 166.525 37.320 167.345 ;
        RECT 40.145 167.205 41.065 167.435 ;
        RECT 44.370 167.205 45.300 167.435 ;
        RECT 37.600 166.525 41.065 167.205 ;
        RECT 41.400 166.525 45.300 167.205 ;
        RECT 45.320 166.525 46.670 167.435 ;
        RECT 55.890 167.205 56.820 167.435 ;
        RECT 46.690 166.525 55.795 167.205 ;
        RECT 55.890 166.525 59.790 167.205 ;
        RECT 60.500 166.610 60.930 167.395 ;
        RECT 60.960 166.525 62.310 167.435 ;
        RECT 62.330 166.525 64.160 167.335 ;
        RECT 64.180 166.525 65.530 167.435 ;
        RECT 68.750 167.205 69.680 167.435 ;
        RECT 71.050 167.205 71.970 167.425 ;
        RECT 78.050 167.325 78.970 167.435 ;
        RECT 80.950 167.345 81.900 167.435 ;
        RECT 76.635 167.205 78.970 167.325 ;
        RECT 65.780 166.525 69.680 167.205 ;
        RECT 69.690 166.525 78.970 167.205 ;
        RECT 79.970 166.525 81.900 167.345 ;
        RECT 85.310 167.205 86.240 167.435 ;
        RECT 82.340 166.525 86.240 167.205 ;
        RECT 86.260 166.610 86.690 167.395 ;
        RECT 86.710 167.235 87.655 167.435 ;
        RECT 86.710 166.555 89.460 167.235 ;
        RECT 86.710 166.525 87.655 166.555 ;
        RECT 18.310 166.315 18.480 166.525 ;
        RECT 29.810 166.505 29.980 166.525 ;
        RECT 19.745 166.365 19.865 166.475 ;
        RECT 20.150 166.315 20.320 166.505 ;
        RECT 22.505 166.365 22.625 166.475 ;
        RECT 22.910 166.315 23.080 166.505 ;
        RECT 24.750 166.315 24.920 166.505 ;
        RECT 29.805 166.335 29.980 166.505 ;
        RECT 30.325 166.365 30.445 166.475 ;
        RECT 18.170 165.505 19.540 166.315 ;
        RECT 20.010 165.635 21.840 166.315 ;
        RECT 21.860 165.445 22.290 166.230 ;
        RECT 22.770 165.635 24.600 166.315 ;
        RECT 24.610 165.635 27.350 166.315 ;
        RECT 27.370 166.285 28.315 166.315 ;
        RECT 29.805 166.285 29.975 166.335 ;
        RECT 33.490 166.315 33.660 166.505 ;
        RECT 33.955 166.315 34.125 166.505 ;
        RECT 34.135 166.335 34.305 166.525 ;
        RECT 37.170 166.505 37.320 166.525 ;
        RECT 37.170 166.335 37.340 166.505 ;
        RECT 37.630 166.335 37.800 166.525 ;
        RECT 44.715 166.335 44.885 166.525 ;
        RECT 46.370 166.335 46.540 166.525 ;
        RECT 46.830 166.315 47.000 166.525 ;
        RECT 47.345 166.365 47.465 166.475 ;
        RECT 48.210 166.315 48.380 166.505 ;
        RECT 56.305 166.335 56.475 166.525 ;
        RECT 58.790 166.315 58.960 166.505 ;
        RECT 60.170 166.475 60.340 166.505 ;
        RECT 60.170 166.365 60.345 166.475 ;
        RECT 60.170 166.315 60.340 166.365 ;
        RECT 60.630 166.315 60.800 166.505 ;
        RECT 62.010 166.335 62.180 166.525 ;
        RECT 63.850 166.335 64.020 166.525 ;
        RECT 65.230 166.335 65.400 166.525 ;
        RECT 69.095 166.335 69.265 166.525 ;
        RECT 69.830 166.335 70.000 166.525 ;
        RECT 79.970 166.505 80.120 166.525 ;
        RECT 73.050 166.315 73.220 166.505 ;
        RECT 74.430 166.360 74.590 166.470 ;
        RECT 74.890 166.315 75.060 166.505 ;
        RECT 78.570 166.315 78.740 166.505 ;
        RECT 79.545 166.365 79.665 166.475 ;
        RECT 79.950 166.335 80.120 166.505 ;
        RECT 85.655 166.335 85.825 166.525 ;
        RECT 88.230 166.315 88.400 166.505 ;
        RECT 89.145 166.335 89.315 166.555 ;
        RECT 89.470 166.525 92.945 167.435 ;
        RECT 96.350 167.205 97.280 167.435 ;
        RECT 93.380 166.525 97.280 167.205 ;
        RECT 97.290 166.525 100.040 167.335 ;
        RECT 103.250 167.205 104.180 167.435 ;
        RECT 100.280 166.525 104.180 167.205 ;
        RECT 104.660 166.525 106.010 167.435 ;
        RECT 106.030 166.525 107.400 167.335 ;
        RECT 107.410 166.525 111.080 167.335 ;
        RECT 111.090 166.525 112.460 167.335 ;
        RECT 89.615 166.505 89.785 166.525 ;
        RECT 89.610 166.335 89.785 166.505 ;
        RECT 96.695 166.335 96.865 166.525 ;
        RECT 89.610 166.315 89.780 166.335 ;
        RECT 98.810 166.315 98.980 166.505 ;
        RECT 99.730 166.335 99.900 166.525 ;
        RECT 100.650 166.315 100.820 166.505 ;
        RECT 103.595 166.335 103.765 166.525 ;
        RECT 104.385 166.365 104.505 166.475 ;
        RECT 105.710 166.335 105.880 166.525 ;
        RECT 107.090 166.335 107.260 166.525 ;
        RECT 110.310 166.315 110.480 166.505 ;
        RECT 110.770 166.475 110.940 166.525 ;
        RECT 110.770 166.365 110.945 166.475 ;
        RECT 110.770 166.335 110.940 166.365 ;
        RECT 112.150 166.315 112.320 166.525 ;
        RECT 23.255 165.405 24.600 165.635 ;
        RECT 27.370 165.605 30.120 166.285 ;
        RECT 30.225 165.635 33.690 166.315 ;
        RECT 27.370 165.405 28.315 165.605 ;
        RECT 30.225 165.405 31.145 165.635 ;
        RECT 33.810 165.405 37.285 166.315 ;
        RECT 37.860 165.635 47.140 166.315 ;
        RECT 37.860 165.515 40.195 165.635 ;
        RECT 37.860 165.405 38.780 165.515 ;
        RECT 44.860 165.415 45.780 165.635 ;
        RECT 47.620 165.445 48.050 166.230 ;
        RECT 48.080 165.405 49.430 166.315 ;
        RECT 49.820 165.635 59.100 166.315 ;
        RECT 49.820 165.515 52.155 165.635 ;
        RECT 49.820 165.405 50.740 165.515 ;
        RECT 56.820 165.415 57.740 165.635 ;
        RECT 59.110 165.505 60.480 166.315 ;
        RECT 60.600 165.635 64.065 166.315 ;
        RECT 63.145 165.405 64.065 165.635 ;
        RECT 64.170 165.635 73.360 166.315 ;
        RECT 64.170 165.405 65.090 165.635 ;
        RECT 67.920 165.415 68.850 165.635 ;
        RECT 73.380 165.445 73.810 166.230 ;
        RECT 74.760 165.405 76.110 166.315 ;
        RECT 76.140 165.635 78.880 166.315 ;
        RECT 79.260 165.635 88.540 166.315 ;
        RECT 79.260 165.515 81.595 165.635 ;
        RECT 79.260 165.405 80.180 165.515 ;
        RECT 86.260 165.415 87.180 165.635 ;
        RECT 88.560 165.405 89.910 166.315 ;
        RECT 89.930 165.635 99.120 166.315 ;
        RECT 89.930 165.405 90.850 165.635 ;
        RECT 93.680 165.415 94.610 165.635 ;
        RECT 99.140 165.445 99.570 166.230 ;
        RECT 99.590 165.505 100.960 166.315 ;
        RECT 101.340 165.635 110.620 166.315 ;
        RECT 101.340 165.515 103.675 165.635 ;
        RECT 101.340 165.405 102.260 165.515 ;
        RECT 108.340 165.415 109.260 165.635 ;
        RECT 111.090 165.505 112.460 166.315 ;
      LAYER nwell ;
        RECT 17.975 162.285 112.655 165.115 ;
      LAYER pwell ;
        RECT 18.170 161.085 19.540 161.895 ;
        RECT 20.010 161.765 21.355 161.995 ;
        RECT 24.505 161.765 25.425 161.995 ;
        RECT 20.010 161.085 21.840 161.765 ;
        RECT 21.960 161.085 25.425 161.765 ;
        RECT 25.530 161.765 26.450 161.995 ;
        RECT 29.280 161.765 30.210 161.985 ;
        RECT 25.530 161.085 34.720 161.765 ;
        RECT 34.740 161.170 35.170 161.955 ;
        RECT 47.505 161.765 48.425 161.995 ;
        RECT 51.185 161.765 52.105 161.995 ;
        RECT 55.410 161.765 56.340 161.995 ;
        RECT 35.275 161.085 44.380 161.765 ;
        RECT 44.960 161.085 48.425 161.765 ;
        RECT 48.640 161.085 52.105 161.765 ;
        RECT 52.440 161.085 56.340 161.765 ;
        RECT 57.010 161.085 59.100 161.895 ;
        RECT 59.120 161.085 60.470 161.995 ;
        RECT 60.500 161.170 60.930 161.955 ;
        RECT 64.610 161.765 65.540 161.995 ;
        RECT 61.640 161.085 65.540 161.765 ;
        RECT 65.550 161.085 66.920 161.895 ;
        RECT 69.585 161.765 70.505 161.995 ;
        RECT 80.270 161.765 81.200 161.995 ;
        RECT 67.040 161.085 70.505 161.765 ;
        RECT 71.155 161.085 80.260 161.765 ;
        RECT 80.270 161.085 84.170 161.765 ;
        RECT 84.410 161.085 85.775 161.765 ;
        RECT 86.260 161.170 86.690 161.955 ;
        RECT 99.110 161.765 100.040 161.995 ;
        RECT 86.710 161.085 95.815 161.765 ;
        RECT 96.140 161.085 100.040 161.765 ;
        RECT 100.420 161.885 101.340 161.995 ;
        RECT 100.420 161.765 102.755 161.885 ;
        RECT 107.420 161.765 108.340 161.985 ;
        RECT 100.420 161.085 109.700 161.765 ;
        RECT 109.710 161.085 111.080 161.895 ;
        RECT 111.090 161.085 112.460 161.895 ;
        RECT 18.310 160.875 18.480 161.085 ;
        RECT 19.745 160.925 19.865 161.035 ;
        RECT 20.150 160.920 20.310 161.030 ;
        RECT 21.530 160.875 21.700 161.085 ;
        RECT 21.990 160.895 22.160 161.085 ;
        RECT 32.570 160.875 32.740 161.065 ;
        RECT 33.305 160.875 33.475 161.065 ;
        RECT 34.410 160.895 34.580 161.085 ;
        RECT 18.170 160.065 19.540 160.875 ;
        RECT 20.480 159.965 21.830 160.875 ;
        RECT 21.860 160.005 22.290 160.790 ;
        RECT 22.510 160.195 32.880 160.875 ;
        RECT 32.890 160.195 36.790 160.875 ;
        RECT 37.030 160.845 37.975 160.875 ;
        RECT 39.465 160.845 39.635 161.065 ;
        RECT 39.935 160.875 40.105 161.065 ;
        RECT 44.070 160.895 44.240 161.085 ;
        RECT 44.585 160.925 44.705 161.035 ;
        RECT 44.990 160.895 45.160 161.085 ;
        RECT 47.015 160.875 47.185 161.065 ;
        RECT 48.265 160.925 48.385 161.035 ;
        RECT 48.670 160.895 48.840 161.085 ;
        RECT 55.755 160.895 55.925 161.085 ;
        RECT 57.410 160.875 57.580 161.065 ;
        RECT 58.330 160.920 58.490 161.030 ;
        RECT 58.790 160.895 58.960 161.085 ;
        RECT 59.250 160.895 59.420 161.085 ;
        RECT 61.145 160.925 61.265 161.035 ;
        RECT 64.955 160.895 65.125 161.085 ;
        RECT 66.610 160.895 66.780 161.085 ;
        RECT 67.070 160.895 67.240 161.085 ;
        RECT 67.530 160.875 67.700 161.065 ;
        RECT 67.990 160.875 68.160 161.065 ;
        RECT 70.805 160.925 70.925 161.035 ;
        RECT 72.775 160.875 72.945 161.065 ;
        RECT 79.950 160.895 80.120 161.085 ;
        RECT 80.685 160.895 80.855 161.085 ;
        RECT 86.850 161.065 87.020 161.085 ;
        RECT 83.170 160.875 83.340 161.065 ;
        RECT 85.930 160.895 86.100 161.065 ;
        RECT 86.845 160.895 87.020 161.065 ;
        RECT 87.365 160.925 87.485 161.035 ;
        RECT 86.845 160.875 87.015 160.895 ;
        RECT 87.775 160.875 87.945 161.065 ;
        RECT 91.450 160.875 91.620 161.065 ;
        RECT 98.535 160.875 98.705 161.065 ;
        RECT 99.455 160.895 99.625 161.085 ;
        RECT 102.945 160.875 103.115 161.065 ;
        RECT 103.410 160.875 103.580 161.065 ;
        RECT 105.710 160.875 105.880 161.065 ;
        RECT 107.090 160.875 107.260 161.065 ;
        RECT 109.390 160.895 109.560 161.085 ;
        RECT 110.770 160.875 110.940 161.085 ;
        RECT 112.150 160.875 112.320 161.085 ;
        RECT 22.510 159.965 24.720 160.195 ;
        RECT 27.440 159.975 28.370 160.195 ;
        RECT 32.890 159.965 33.820 160.195 ;
        RECT 37.030 160.165 39.780 160.845 ;
        RECT 37.030 159.965 37.975 160.165 ;
        RECT 39.790 159.965 43.265 160.875 ;
        RECT 43.700 160.195 47.600 160.875 ;
        RECT 46.670 159.965 47.600 160.195 ;
        RECT 47.620 160.005 48.050 160.790 ;
        RECT 48.530 160.195 57.720 160.875 ;
        RECT 58.650 160.195 67.840 160.875 ;
        RECT 48.530 159.965 49.450 160.195 ;
        RECT 52.280 159.975 53.210 160.195 ;
        RECT 58.650 159.965 59.570 160.195 ;
        RECT 62.400 159.975 63.330 160.195 ;
        RECT 67.860 159.965 69.210 160.875 ;
        RECT 69.460 160.195 73.360 160.875 ;
        RECT 72.430 159.965 73.360 160.195 ;
        RECT 73.380 160.005 73.810 160.790 ;
        RECT 74.200 160.195 83.480 160.875 ;
        RECT 74.200 160.075 76.535 160.195 ;
        RECT 74.200 159.965 75.120 160.075 ;
        RECT 81.200 159.975 82.120 160.195 ;
        RECT 83.685 159.965 87.160 160.875 ;
        RECT 87.630 159.965 91.105 160.875 ;
        RECT 91.420 160.195 94.885 160.875 ;
        RECT 95.220 160.195 99.120 160.875 ;
        RECT 93.965 159.965 94.885 160.195 ;
        RECT 98.190 159.965 99.120 160.195 ;
        RECT 99.140 160.005 99.570 160.790 ;
        RECT 99.785 159.965 103.260 160.875 ;
        RECT 103.280 159.965 104.630 160.875 ;
        RECT 104.660 159.965 106.010 160.875 ;
        RECT 106.030 160.065 107.400 160.875 ;
        RECT 107.410 160.065 111.080 160.875 ;
        RECT 111.090 160.065 112.460 160.875 ;
      LAYER nwell ;
        RECT 17.975 156.845 112.655 159.675 ;
      LAYER pwell ;
        RECT 18.170 155.645 19.540 156.455 ;
        RECT 19.550 155.645 22.300 156.455 ;
        RECT 22.310 155.645 23.680 156.425 ;
        RECT 24.150 155.645 29.660 156.455 ;
        RECT 29.680 155.645 31.030 156.555 ;
        RECT 31.245 155.645 34.720 156.555 ;
        RECT 34.740 155.730 35.170 156.515 ;
        RECT 35.190 156.325 36.535 156.555 ;
        RECT 37.230 156.465 38.180 156.555 ;
        RECT 35.190 155.645 37.020 156.325 ;
        RECT 37.230 155.645 39.160 156.465 ;
        RECT 39.330 155.645 42.805 156.555 ;
        RECT 43.010 156.325 43.930 156.555 ;
        RECT 46.760 156.325 47.690 156.545 ;
        RECT 54.865 156.325 55.785 156.555 ;
        RECT 43.010 155.645 52.200 156.325 ;
        RECT 52.320 155.645 55.785 156.325 ;
        RECT 56.810 155.645 60.285 156.555 ;
        RECT 60.500 155.730 60.930 156.515 ;
        RECT 61.410 155.645 64.885 156.555 ;
        RECT 65.090 155.645 66.460 156.455 ;
        RECT 66.840 156.445 67.760 156.555 ;
        RECT 66.840 156.325 69.175 156.445 ;
        RECT 73.840 156.325 74.760 156.545 ;
        RECT 66.840 155.645 76.120 156.325 ;
        RECT 76.600 155.645 77.950 156.555 ;
        RECT 78.430 155.645 81.180 156.455 ;
        RECT 81.200 155.645 82.550 156.555 ;
        RECT 82.765 155.645 86.240 156.555 ;
        RECT 86.260 155.730 86.690 156.515 ;
        RECT 87.850 156.465 88.800 156.555 ;
        RECT 86.870 155.645 88.800 156.465 ;
        RECT 89.010 155.645 92.485 156.555 ;
        RECT 95.890 156.325 96.820 156.555 ;
        RECT 92.920 155.645 96.820 156.325 ;
        RECT 96.830 155.645 98.200 156.455 ;
        RECT 98.580 156.445 99.500 156.555 ;
        RECT 98.580 156.325 100.915 156.445 ;
        RECT 105.580 156.325 106.500 156.545 ;
        RECT 98.580 155.645 107.860 156.325 ;
        RECT 108.330 155.645 111.080 156.455 ;
        RECT 111.090 155.645 112.460 156.455 ;
        RECT 18.310 155.435 18.480 155.645 ;
        RECT 20.150 155.480 20.310 155.590 ;
        RECT 21.530 155.435 21.700 155.625 ;
        RECT 21.990 155.455 22.160 155.645 ;
        RECT 22.460 155.455 22.630 155.645 ;
        RECT 23.885 155.485 24.005 155.595 ;
        RECT 29.350 155.455 29.520 155.645 ;
        RECT 30.730 155.455 30.900 155.645 ;
        RECT 32.570 155.435 32.740 155.625 ;
        RECT 33.490 155.480 33.650 155.590 ;
        RECT 33.950 155.435 34.120 155.625 ;
        RECT 34.405 155.455 34.575 155.645 ;
        RECT 35.340 155.435 35.510 155.625 ;
        RECT 36.710 155.455 36.880 155.645 ;
        RECT 39.010 155.625 39.160 155.645 ;
        RECT 37.630 155.435 37.800 155.625 ;
        RECT 38.090 155.435 38.260 155.625 ;
        RECT 39.010 155.455 39.180 155.625 ;
        RECT 39.475 155.455 39.645 155.645 ;
        RECT 18.170 154.625 19.540 155.435 ;
        RECT 20.480 154.525 21.830 155.435 ;
        RECT 21.860 154.565 22.290 155.350 ;
        RECT 22.510 154.755 32.880 155.435 ;
        RECT 22.510 154.525 24.720 154.755 ;
        RECT 27.440 154.535 28.370 154.755 ;
        RECT 33.820 154.525 35.170 155.435 ;
        RECT 35.190 154.655 36.560 155.435 ;
        RECT 36.570 154.625 37.940 155.435 ;
        RECT 37.950 154.755 39.780 155.435 ;
        RECT 38.435 154.525 39.780 154.755 ;
        RECT 39.790 155.405 40.735 155.435 ;
        RECT 42.225 155.405 42.395 155.625 ;
        RECT 46.095 155.435 46.265 155.625 ;
        RECT 47.290 155.480 47.450 155.590 ;
        RECT 48.215 155.435 48.385 155.625 ;
        RECT 51.890 155.455 52.060 155.645 ;
        RECT 52.350 155.455 52.520 155.645 ;
        RECT 52.810 155.435 52.980 155.625 ;
        RECT 56.490 155.490 56.650 155.600 ;
        RECT 56.955 155.590 57.125 155.645 ;
        RECT 56.950 155.480 57.125 155.590 ;
        RECT 56.955 155.455 57.125 155.480 ;
        RECT 57.415 155.435 57.585 155.625 ;
        RECT 61.145 155.485 61.265 155.595 ;
        RECT 61.555 155.455 61.725 155.645 ;
        RECT 66.150 155.455 66.320 155.645 ;
        RECT 69.830 155.435 70.000 155.625 ;
        RECT 70.345 155.485 70.465 155.595 ;
        RECT 73.050 155.435 73.220 155.625 ;
        RECT 74.430 155.480 74.590 155.590 ;
        RECT 75.810 155.455 75.980 155.645 ;
        RECT 76.325 155.485 76.445 155.595 ;
        RECT 76.730 155.455 76.900 155.645 ;
        RECT 78.165 155.485 78.285 155.595 ;
        RECT 80.870 155.455 81.040 155.645 ;
        RECT 81.330 155.455 81.500 155.645 ;
        RECT 84.090 155.435 84.260 155.625 ;
        RECT 85.010 155.480 85.170 155.590 ;
        RECT 85.925 155.455 86.095 155.645 ;
        RECT 86.870 155.625 87.020 155.645 ;
        RECT 86.850 155.455 87.020 155.625 ;
        RECT 88.875 155.435 89.045 155.625 ;
        RECT 89.155 155.455 89.325 155.645 ;
        RECT 96.235 155.455 96.405 155.645 ;
        RECT 97.890 155.455 98.060 155.645 ;
        RECT 98.810 155.435 98.980 155.625 ;
        RECT 100.190 155.480 100.350 155.590 ;
        RECT 100.650 155.435 100.820 155.625 ;
        RECT 107.550 155.455 107.720 155.645 ;
        RECT 108.065 155.485 108.185 155.595 ;
        RECT 110.770 155.455 110.940 155.645 ;
        RECT 112.150 155.435 112.320 155.645 ;
        RECT 39.790 154.725 42.540 155.405 ;
        RECT 42.780 154.755 46.680 155.435 ;
        RECT 39.790 154.525 40.735 154.725 ;
        RECT 45.750 154.525 46.680 154.755 ;
        RECT 47.620 154.565 48.050 155.350 ;
        RECT 48.070 154.525 51.545 155.435 ;
        RECT 52.780 154.755 56.245 155.435 ;
        RECT 55.325 154.525 56.245 154.755 ;
        RECT 57.270 154.525 60.745 155.435 ;
        RECT 60.950 154.755 70.140 155.435 ;
        RECT 60.950 154.525 61.870 154.755 ;
        RECT 64.700 154.535 65.630 154.755 ;
        RECT 70.610 154.625 73.360 155.435 ;
        RECT 73.380 154.565 73.810 155.350 ;
        RECT 75.120 154.755 84.400 155.435 ;
        RECT 85.560 154.755 89.460 155.435 ;
        RECT 75.120 154.635 77.455 154.755 ;
        RECT 75.120 154.525 76.040 154.635 ;
        RECT 82.120 154.535 83.040 154.755 ;
        RECT 88.530 154.525 89.460 154.755 ;
        RECT 89.840 154.755 99.120 155.435 ;
        RECT 89.840 154.635 92.175 154.755 ;
        RECT 89.840 154.525 90.760 154.635 ;
        RECT 96.840 154.535 97.760 154.755 ;
        RECT 99.140 154.565 99.570 155.350 ;
        RECT 100.510 154.755 110.880 155.435 ;
        RECT 105.020 154.535 105.950 154.755 ;
        RECT 108.670 154.525 110.880 154.755 ;
        RECT 111.090 154.625 112.460 155.435 ;
      LAYER nwell ;
        RECT 17.975 151.405 112.655 154.235 ;
      LAYER pwell ;
        RECT 18.170 150.205 19.540 151.015 ;
        RECT 20.010 150.205 25.520 151.015 ;
        RECT 25.530 150.885 26.450 151.115 ;
        RECT 29.280 150.885 30.210 151.105 ;
        RECT 25.530 150.205 34.720 150.885 ;
        RECT 34.740 150.290 35.170 151.075 ;
        RECT 35.845 150.205 39.320 151.115 ;
        RECT 39.700 151.005 40.620 151.115 ;
        RECT 39.700 150.885 42.035 151.005 ;
        RECT 46.700 150.885 47.620 151.105 ;
        RECT 39.700 150.205 48.980 150.885 ;
        RECT 49.450 150.205 53.120 151.015 ;
        RECT 53.130 150.915 54.075 151.115 ;
        RECT 53.130 150.235 55.880 150.915 ;
        RECT 59.090 150.885 60.020 151.115 ;
        RECT 53.130 150.205 54.075 150.235 ;
        RECT 18.310 149.995 18.480 150.205 ;
        RECT 19.745 150.045 19.865 150.155 ;
        RECT 20.150 150.040 20.310 150.150 ;
        RECT 21.530 149.995 21.700 150.185 ;
        RECT 25.210 150.015 25.380 150.205 ;
        RECT 32.570 149.995 32.740 150.185 ;
        RECT 34.410 150.015 34.580 150.205 ;
        RECT 35.385 150.045 35.505 150.155 ;
        RECT 39.005 150.015 39.175 150.205 ;
        RECT 41.770 149.995 41.940 150.185 ;
        RECT 42.285 150.045 42.405 150.155 ;
        RECT 42.690 149.995 42.860 150.185 ;
        RECT 44.075 149.995 44.245 150.185 ;
        RECT 48.265 150.045 48.385 150.155 ;
        RECT 48.670 150.015 48.840 150.205 ;
        RECT 49.185 150.045 49.305 150.155 ;
        RECT 51.890 149.995 52.060 150.185 ;
        RECT 52.810 150.015 52.980 150.205 ;
        RECT 55.565 150.015 55.735 150.235 ;
        RECT 56.120 150.205 60.020 150.885 ;
        RECT 60.500 150.290 60.930 151.075 ;
        RECT 61.150 151.025 62.100 151.115 ;
        RECT 61.150 150.205 63.080 151.025 ;
        RECT 66.450 150.885 67.380 151.115 ;
        RECT 63.480 150.205 67.380 150.885 ;
        RECT 67.390 150.205 69.220 151.015 ;
        RECT 69.600 151.005 70.520 151.115 ;
        RECT 69.600 150.885 71.935 151.005 ;
        RECT 76.600 150.885 77.520 151.105 ;
        RECT 82.090 150.885 83.020 151.115 ;
        RECT 69.600 150.205 78.880 150.885 ;
        RECT 79.120 150.205 83.020 150.885 ;
        RECT 83.500 150.205 86.240 150.885 ;
        RECT 86.260 150.290 86.690 151.075 ;
        RECT 86.710 150.205 88.080 151.015 ;
        RECT 89.895 150.915 90.840 151.115 ;
        RECT 88.090 150.235 90.840 150.915 ;
        RECT 59.435 150.015 59.605 150.205 ;
        RECT 62.930 150.185 63.080 150.205 ;
        RECT 60.225 150.045 60.345 150.155 ;
        RECT 61.550 149.995 61.720 150.185 ;
        RECT 62.930 150.015 63.100 150.185 ;
        RECT 63.390 149.995 63.560 150.185 ;
        RECT 63.850 149.995 64.020 150.185 ;
        RECT 65.285 150.045 65.405 150.155 ;
        RECT 66.795 150.015 66.965 150.205 ;
        RECT 68.910 149.995 69.080 150.205 ;
        RECT 72.775 149.995 72.945 150.185 ;
        RECT 74.890 149.995 75.060 150.185 ;
        RECT 75.405 150.045 75.525 150.155 ;
        RECT 78.110 149.995 78.280 150.185 ;
        RECT 78.570 150.015 78.740 150.205 ;
        RECT 79.490 149.995 79.660 150.185 ;
        RECT 80.005 150.045 80.125 150.155 ;
        RECT 81.790 149.995 81.960 150.185 ;
        RECT 82.435 150.015 82.605 150.205 ;
        RECT 83.225 150.045 83.345 150.155 ;
        RECT 85.930 150.015 86.100 150.205 ;
        RECT 87.770 150.015 87.940 150.205 ;
        RECT 88.235 150.015 88.405 150.235 ;
        RECT 89.895 150.205 90.840 150.235 ;
        RECT 91.770 150.205 94.510 150.885 ;
        RECT 95.000 150.205 96.350 151.115 ;
        RECT 96.830 150.205 100.500 151.015 ;
        RECT 100.510 150.205 106.020 151.015 ;
        RECT 106.040 150.205 107.390 151.115 ;
        RECT 107.410 150.205 111.080 151.015 ;
        RECT 111.090 150.205 112.460 151.015 ;
        RECT 91.450 149.995 91.620 150.185 ;
        RECT 91.910 150.015 92.080 150.205 ;
        RECT 93.290 149.995 93.460 150.185 ;
        RECT 94.725 150.045 94.845 150.155 ;
        RECT 96.050 150.015 96.220 150.205 ;
        RECT 96.565 150.045 96.685 150.155 ;
        RECT 98.810 149.995 98.980 150.185 ;
        RECT 99.785 150.045 99.905 150.155 ;
        RECT 100.190 150.015 100.360 150.205 ;
        RECT 101.110 149.995 101.280 150.185 ;
        RECT 101.575 149.995 101.745 150.185 ;
        RECT 105.250 149.995 105.420 150.185 ;
        RECT 105.710 150.015 105.880 150.205 ;
        RECT 106.170 150.015 106.340 150.205 ;
        RECT 110.770 149.995 110.940 150.205 ;
        RECT 112.150 149.995 112.320 150.205 ;
        RECT 18.170 149.185 19.540 149.995 ;
        RECT 20.480 149.085 21.830 149.995 ;
        RECT 21.860 149.125 22.290 149.910 ;
        RECT 22.510 149.315 32.880 149.995 ;
        RECT 32.890 149.315 42.080 149.995 ;
        RECT 22.510 149.085 24.720 149.315 ;
        RECT 27.440 149.095 28.370 149.315 ;
        RECT 32.890 149.085 33.810 149.315 ;
        RECT 36.640 149.095 37.570 149.315 ;
        RECT 42.560 149.085 43.910 149.995 ;
        RECT 43.930 149.085 47.405 149.995 ;
        RECT 47.620 149.125 48.050 149.910 ;
        RECT 48.530 149.185 52.200 149.995 ;
        RECT 52.580 149.315 61.860 149.995 ;
        RECT 52.580 149.195 54.915 149.315 ;
        RECT 52.580 149.085 53.500 149.195 ;
        RECT 59.580 149.095 60.500 149.315 ;
        RECT 61.870 149.185 63.700 149.995 ;
        RECT 63.720 149.085 65.070 149.995 ;
        RECT 65.550 149.185 69.220 149.995 ;
        RECT 69.460 149.315 73.360 149.995 ;
        RECT 72.430 149.085 73.360 149.315 ;
        RECT 73.380 149.125 73.810 149.910 ;
        RECT 73.840 149.085 75.190 149.995 ;
        RECT 75.670 149.185 78.420 149.995 ;
        RECT 78.440 149.085 79.790 149.995 ;
        RECT 80.270 149.185 82.100 149.995 ;
        RECT 82.480 149.315 91.760 149.995 ;
        RECT 82.480 149.195 84.815 149.315 ;
        RECT 82.480 149.085 83.400 149.195 ;
        RECT 89.480 149.095 90.400 149.315 ;
        RECT 91.770 149.185 93.600 149.995 ;
        RECT 93.610 149.185 99.120 149.995 ;
        RECT 99.140 149.125 99.570 149.910 ;
        RECT 100.060 149.085 101.410 149.995 ;
        RECT 101.430 149.085 104.040 149.995 ;
        RECT 104.190 149.185 105.560 149.995 ;
        RECT 105.570 149.185 111.080 149.995 ;
        RECT 111.090 149.185 112.460 149.995 ;
      LAYER nwell ;
        RECT 17.975 145.965 112.655 148.795 ;
      LAYER pwell ;
        RECT 18.170 144.765 19.540 145.575 ;
        RECT 20.010 144.765 25.520 145.575 ;
        RECT 28.185 145.445 29.105 145.675 ;
        RECT 25.640 144.765 29.105 145.445 ;
        RECT 29.220 144.765 30.570 145.675 ;
        RECT 33.790 145.445 34.720 145.675 ;
        RECT 30.820 144.765 34.720 145.445 ;
        RECT 34.740 144.850 35.170 145.635 ;
        RECT 38.850 145.445 39.780 145.675 ;
        RECT 43.210 145.585 44.160 145.675 ;
        RECT 35.880 144.765 39.780 145.445 ;
        RECT 40.250 144.765 43.000 145.575 ;
        RECT 43.210 144.765 45.140 145.585 ;
        RECT 46.230 144.765 49.900 145.575 ;
        RECT 53.110 145.445 54.040 145.675 ;
        RECT 50.140 144.765 54.040 145.445 ;
        RECT 54.050 144.765 55.420 145.575 ;
        RECT 55.440 144.765 56.790 145.675 ;
        RECT 56.810 144.765 60.480 145.575 ;
        RECT 60.500 144.850 60.930 145.635 ;
        RECT 61.035 144.765 70.140 145.445 ;
        RECT 70.610 144.765 73.360 145.575 ;
        RECT 73.370 144.765 78.880 145.575 ;
        RECT 78.900 144.765 80.250 145.675 ;
        RECT 80.270 144.765 82.880 145.675 ;
        RECT 83.490 144.765 86.240 145.575 ;
        RECT 86.260 144.850 86.690 145.635 ;
        RECT 86.710 144.765 88.080 145.575 ;
        RECT 88.130 144.765 92.680 145.675 ;
        RECT 92.690 144.765 96.360 145.575 ;
        RECT 96.740 145.565 97.660 145.675 ;
        RECT 96.740 145.445 99.075 145.565 ;
        RECT 103.740 145.445 104.660 145.665 ;
        RECT 96.740 144.765 106.020 145.445 ;
        RECT 106.040 144.765 107.390 145.675 ;
        RECT 107.410 144.765 111.080 145.575 ;
        RECT 111.090 144.765 112.460 145.575 ;
        RECT 18.310 144.555 18.480 144.765 ;
        RECT 19.745 144.605 19.865 144.715 ;
        RECT 21.530 144.555 21.700 144.745 ;
        RECT 25.210 144.575 25.380 144.765 ;
        RECT 25.670 144.555 25.840 144.765 ;
        RECT 30.270 144.575 30.440 144.765 ;
        RECT 31.190 144.555 31.360 144.745 ;
        RECT 34.135 144.575 34.305 144.765 ;
        RECT 34.870 144.555 35.040 144.745 ;
        RECT 35.385 144.605 35.505 144.715 ;
        RECT 39.010 144.555 39.180 144.745 ;
        RECT 39.195 144.575 39.365 144.765 ;
        RECT 39.985 144.605 40.105 144.715 ;
        RECT 42.690 144.575 42.860 144.765 ;
        RECT 44.990 144.745 45.140 144.765 ;
        RECT 44.530 144.555 44.700 144.745 ;
        RECT 44.990 144.555 45.160 144.745 ;
        RECT 45.910 144.610 46.070 144.720 ;
        RECT 46.370 144.555 46.540 144.745 ;
        RECT 48.265 144.605 48.385 144.715 ;
        RECT 49.590 144.575 49.760 144.765 ;
        RECT 53.455 144.575 53.625 144.765 ;
        RECT 55.110 144.575 55.280 144.765 ;
        RECT 55.570 144.575 55.740 144.765 ;
        RECT 57.870 144.555 58.040 144.745 ;
        RECT 59.250 144.555 59.420 144.745 ;
        RECT 60.170 144.575 60.340 144.765 ;
        RECT 68.450 144.555 68.620 144.745 ;
        RECT 68.965 144.605 69.085 144.715 ;
        RECT 69.830 144.575 70.000 144.765 ;
        RECT 70.345 144.605 70.465 144.715 ;
        RECT 72.775 144.555 72.945 144.745 ;
        RECT 73.050 144.575 73.220 144.765 ;
        RECT 73.970 144.555 74.140 144.745 ;
        RECT 78.570 144.575 78.740 144.765 ;
        RECT 79.030 144.575 79.200 144.765 ;
        RECT 80.415 144.575 80.585 144.765 ;
        RECT 83.225 144.605 83.345 144.715 ;
        RECT 84.090 144.600 84.250 144.710 ;
        RECT 84.550 144.555 84.720 144.745 ;
        RECT 85.930 144.575 86.100 144.765 ;
        RECT 87.770 144.575 87.940 144.765 ;
        RECT 89.150 144.555 89.320 144.745 ;
        RECT 92.370 144.575 92.540 144.765 ;
        RECT 94.670 144.555 94.840 144.745 ;
        RECT 96.050 144.575 96.220 144.765 ;
        RECT 98.535 144.555 98.705 144.745 ;
        RECT 99.730 144.555 99.900 144.745 ;
        RECT 105.710 144.575 105.880 144.765 ;
        RECT 107.090 144.575 107.260 144.765 ;
        RECT 109.445 144.605 109.565 144.715 ;
        RECT 110.770 144.555 110.940 144.765 ;
        RECT 112.150 144.555 112.320 144.765 ;
        RECT 18.170 143.745 19.540 144.555 ;
        RECT 20.010 143.745 21.840 144.555 ;
        RECT 21.860 143.685 22.290 144.470 ;
        RECT 22.310 143.745 25.980 144.555 ;
        RECT 25.990 143.745 31.500 144.555 ;
        RECT 31.605 143.875 35.070 144.555 ;
        RECT 31.605 143.645 32.525 143.875 ;
        RECT 35.650 143.745 39.320 144.555 ;
        RECT 39.330 143.745 44.840 144.555 ;
        RECT 44.860 143.645 46.210 144.555 ;
        RECT 46.240 143.645 47.590 144.555 ;
        RECT 47.620 143.685 48.050 144.470 ;
        RECT 48.900 143.875 58.180 144.555 ;
        RECT 48.900 143.755 51.235 143.875 ;
        RECT 48.900 143.645 49.820 143.755 ;
        RECT 55.900 143.655 56.820 143.875 ;
        RECT 58.190 143.745 59.560 144.555 ;
        RECT 59.570 143.875 68.760 144.555 ;
        RECT 69.460 143.875 73.360 144.555 ;
        RECT 59.570 143.645 60.490 143.875 ;
        RECT 63.320 143.655 64.250 143.875 ;
        RECT 72.430 143.645 73.360 143.875 ;
        RECT 73.380 143.685 73.810 144.470 ;
        RECT 73.830 143.875 83.110 144.555 ;
        RECT 75.190 143.655 76.110 143.875 ;
        RECT 80.775 143.755 83.110 143.875 ;
        RECT 82.190 143.645 83.110 143.755 ;
        RECT 84.410 143.645 88.960 144.555 ;
        RECT 89.010 143.645 93.560 144.555 ;
        RECT 93.620 143.645 94.970 144.555 ;
        RECT 95.220 143.875 99.120 144.555 ;
        RECT 98.190 143.645 99.120 143.875 ;
        RECT 99.140 143.685 99.570 144.470 ;
        RECT 99.590 143.875 108.870 144.555 ;
        RECT 100.950 143.655 101.870 143.875 ;
        RECT 106.535 143.755 108.870 143.875 ;
        RECT 109.710 143.775 111.080 144.555 ;
        RECT 107.950 143.645 108.870 143.755 ;
        RECT 111.090 143.745 112.460 144.555 ;
      LAYER nwell ;
        RECT 17.975 140.525 112.655 143.355 ;
      LAYER pwell ;
        RECT 18.170 139.325 19.540 140.135 ;
        RECT 20.470 139.325 24.140 140.135 ;
        RECT 24.150 139.325 29.660 140.135 ;
        RECT 29.680 139.325 31.030 140.235 ;
        RECT 31.050 139.325 34.720 140.135 ;
        RECT 34.740 139.410 35.170 140.195 ;
        RECT 35.660 139.325 37.010 140.235 ;
        RECT 37.490 139.325 40.965 140.235 ;
        RECT 41.170 139.325 44.645 140.235 ;
        RECT 45.220 140.125 46.140 140.235 ;
        RECT 45.220 140.005 47.555 140.125 ;
        RECT 52.220 140.005 53.140 140.225 ;
        RECT 54.510 140.005 55.440 140.235 ;
        RECT 45.220 139.325 54.500 140.005 ;
        RECT 54.510 139.325 58.410 140.005 ;
        RECT 58.660 139.325 60.010 140.235 ;
        RECT 60.500 139.410 60.930 140.195 ;
        RECT 60.960 139.325 62.310 140.235 ;
        RECT 65.530 140.005 66.460 140.235 ;
        RECT 62.560 139.325 66.460 140.005 ;
        RECT 66.470 139.325 67.840 140.135 ;
        RECT 68.220 140.125 69.140 140.235 ;
        RECT 68.220 140.005 70.555 140.125 ;
        RECT 75.220 140.005 76.140 140.225 ;
        RECT 80.625 140.005 81.545 140.235 ;
        RECT 68.220 139.325 77.500 140.005 ;
        RECT 78.080 139.325 81.545 140.005 ;
        RECT 81.660 139.325 83.010 140.235 ;
        RECT 83.030 139.325 86.240 140.235 ;
        RECT 86.260 139.410 86.690 140.195 ;
        RECT 87.850 140.145 88.800 140.235 ;
        RECT 86.870 139.325 88.800 140.145 ;
        RECT 89.010 139.325 92.485 140.235 ;
        RECT 95.890 140.005 96.820 140.235 ;
        RECT 92.920 139.325 96.820 140.005 ;
        RECT 97.200 140.125 98.120 140.235 ;
        RECT 97.200 140.005 99.535 140.125 ;
        RECT 104.200 140.005 105.120 140.225 ;
        RECT 97.200 139.325 106.480 140.005 ;
        RECT 107.410 139.325 111.080 140.135 ;
        RECT 111.090 139.325 112.460 140.135 ;
        RECT 18.310 139.115 18.480 139.325 ;
        RECT 20.150 139.160 20.310 139.280 ;
        RECT 21.530 139.115 21.700 139.305 ;
        RECT 23.370 139.115 23.540 139.305 ;
        RECT 23.830 139.115 24.000 139.325 ;
        RECT 29.350 139.135 29.520 139.325 ;
        RECT 30.730 139.135 30.900 139.325 ;
        RECT 34.410 139.135 34.580 139.325 ;
        RECT 35.385 139.165 35.505 139.275 ;
        RECT 36.710 139.135 36.880 139.325 ;
        RECT 37.225 139.165 37.345 139.275 ;
        RECT 37.635 139.135 37.805 139.325 ;
        RECT 41.315 139.135 41.485 139.325 ;
        RECT 41.770 139.115 41.940 139.305 ;
        RECT 43.610 139.115 43.780 139.305 ;
        RECT 44.075 139.115 44.245 139.305 ;
        RECT 48.670 139.160 48.830 139.270 ;
        RECT 54.190 139.135 54.360 139.325 ;
        RECT 54.925 139.135 55.095 139.325 ;
        RECT 58.330 139.115 58.500 139.305 ;
        RECT 58.790 139.115 58.960 139.305 ;
        RECT 59.710 139.135 59.880 139.325 ;
        RECT 60.225 139.165 60.345 139.275 ;
        RECT 61.090 139.135 61.260 139.325 ;
        RECT 62.475 139.115 62.645 139.305 ;
        RECT 65.875 139.135 66.045 139.325 ;
        RECT 67.530 139.115 67.700 139.325 ;
        RECT 67.995 139.115 68.165 139.305 ;
        RECT 72.590 139.115 72.760 139.305 ;
        RECT 73.105 139.165 73.225 139.275 ;
        RECT 77.190 139.135 77.360 139.325 ;
        RECT 77.375 139.115 77.545 139.305 ;
        RECT 77.705 139.165 77.825 139.275 ;
        RECT 78.110 139.135 78.280 139.325 ;
        RECT 79.030 139.115 79.200 139.305 ;
        RECT 82.710 139.135 82.880 139.325 ;
        RECT 83.170 139.135 83.340 139.325 ;
        RECT 86.870 139.305 87.020 139.325 ;
        RECT 86.850 139.135 87.020 139.305 ;
        RECT 88.690 139.115 88.860 139.305 ;
        RECT 89.155 139.115 89.325 139.325 ;
        RECT 92.885 139.165 93.005 139.275 ;
        RECT 94.670 139.115 94.840 139.305 ;
        RECT 96.235 139.135 96.405 139.325 ;
        RECT 98.535 139.115 98.705 139.305 ;
        RECT 100.190 139.160 100.350 139.270 ;
        RECT 100.650 139.115 100.820 139.305 ;
        RECT 106.170 139.135 106.340 139.325 ;
        RECT 107.090 139.170 107.250 139.280 ;
        RECT 110.770 139.135 110.940 139.325 ;
        RECT 112.150 139.115 112.320 139.325 ;
        RECT 18.170 138.305 19.540 139.115 ;
        RECT 20.480 138.205 21.830 139.115 ;
        RECT 21.860 138.245 22.290 139.030 ;
        RECT 22.310 138.305 23.680 139.115 ;
        RECT 23.690 138.435 32.880 139.115 ;
        RECT 28.200 138.215 29.130 138.435 ;
        RECT 31.960 138.205 32.880 138.435 ;
        RECT 32.890 138.435 42.080 139.115 ;
        RECT 42.090 138.435 43.920 139.115 ;
        RECT 32.890 138.205 33.810 138.435 ;
        RECT 36.640 138.215 37.570 138.435 ;
        RECT 42.090 138.205 43.435 138.435 ;
        RECT 43.930 138.205 47.405 139.115 ;
        RECT 47.620 138.245 48.050 139.030 ;
        RECT 49.360 138.435 58.640 139.115 ;
        RECT 58.760 138.435 62.225 139.115 ;
        RECT 49.360 138.315 51.695 138.435 ;
        RECT 49.360 138.205 50.280 138.315 ;
        RECT 56.360 138.215 57.280 138.435 ;
        RECT 61.305 138.205 62.225 138.435 ;
        RECT 62.330 138.205 65.805 139.115 ;
        RECT 66.010 138.305 67.840 139.115 ;
        RECT 67.850 138.205 71.325 139.115 ;
        RECT 71.540 138.205 72.890 139.115 ;
        RECT 73.380 138.245 73.810 139.030 ;
        RECT 74.060 138.435 77.960 139.115 ;
        RECT 77.030 138.205 77.960 138.435 ;
        RECT 77.970 138.305 79.340 139.115 ;
        RECT 79.720 138.435 89.000 139.115 ;
        RECT 79.720 138.315 82.055 138.435 ;
        RECT 79.720 138.205 80.640 138.315 ;
        RECT 86.720 138.215 87.640 138.435 ;
        RECT 89.010 138.205 92.485 139.115 ;
        RECT 93.150 138.305 94.980 139.115 ;
        RECT 95.220 138.435 99.120 139.115 ;
        RECT 98.190 138.205 99.120 138.435 ;
        RECT 99.140 138.245 99.570 139.030 ;
        RECT 100.510 138.435 110.880 139.115 ;
        RECT 105.020 138.215 105.950 138.435 ;
        RECT 108.670 138.205 110.880 138.435 ;
        RECT 111.090 138.305 112.460 139.115 ;
      LAYER nwell ;
        RECT 17.975 135.085 112.655 137.915 ;
      LAYER pwell ;
        RECT 18.170 133.885 19.540 134.695 ;
        RECT 23.325 134.565 24.245 134.795 ;
        RECT 29.565 134.565 30.485 134.795 ;
        RECT 20.480 133.885 23.220 134.565 ;
        RECT 23.325 133.885 26.790 134.565 ;
        RECT 27.020 133.885 30.485 134.565 ;
        RECT 30.590 134.565 31.520 134.795 ;
        RECT 30.590 133.885 34.490 134.565 ;
        RECT 34.740 133.970 35.170 134.755 ;
        RECT 35.650 134.565 36.995 134.795 ;
        RECT 40.690 134.565 41.620 134.795 ;
        RECT 35.650 133.885 37.480 134.565 ;
        RECT 37.720 133.885 41.620 134.565 ;
        RECT 42.090 133.885 45.565 134.795 ;
        RECT 46.230 133.885 51.740 134.695 ;
        RECT 54.950 134.565 55.880 134.795 ;
        RECT 51.980 133.885 55.880 134.565 ;
        RECT 56.360 133.885 57.710 134.795 ;
        RECT 57.870 133.885 60.480 134.795 ;
        RECT 60.500 133.970 60.930 134.755 ;
        RECT 61.090 133.885 63.700 134.795 ;
        RECT 66.910 134.565 67.840 134.795 ;
        RECT 63.940 133.885 67.840 134.565 ;
        RECT 67.850 133.885 70.590 134.565 ;
        RECT 70.620 133.885 73.360 134.565 ;
        RECT 73.565 133.885 77.040 134.795 ;
        RECT 80.250 134.565 81.180 134.795 ;
        RECT 85.310 134.565 86.240 134.795 ;
        RECT 77.280 133.885 81.180 134.565 ;
        RECT 82.340 133.885 86.240 134.565 ;
        RECT 86.260 133.970 86.690 134.755 ;
        RECT 86.710 133.885 89.450 134.565 ;
        RECT 89.470 133.885 92.945 134.795 ;
        RECT 93.345 133.885 96.820 134.795 ;
        RECT 96.830 133.885 99.580 134.695 ;
        RECT 99.600 133.885 100.950 134.795 ;
        RECT 100.970 133.885 103.710 134.565 ;
        RECT 104.190 133.885 106.020 134.695 ;
        RECT 106.040 133.885 107.390 134.795 ;
        RECT 107.410 133.885 111.080 134.695 ;
        RECT 111.090 133.885 112.460 134.695 ;
        RECT 18.310 133.675 18.480 133.885 ;
        RECT 20.150 133.720 20.310 133.840 ;
        RECT 21.530 133.675 21.700 133.865 ;
        RECT 22.450 133.675 22.620 133.865 ;
        RECT 22.910 133.695 23.080 133.885 ;
        RECT 26.590 133.695 26.760 133.885 ;
        RECT 27.050 133.695 27.220 133.885 ;
        RECT 31.005 133.695 31.175 133.885 ;
        RECT 34.870 133.675 35.040 133.865 ;
        RECT 35.385 133.725 35.505 133.835 ;
        RECT 36.250 133.675 36.420 133.865 ;
        RECT 36.715 133.675 36.885 133.865 ;
        RECT 37.170 133.695 37.340 133.885 ;
        RECT 40.390 133.675 40.560 133.865 ;
        RECT 41.035 133.695 41.205 133.885 ;
        RECT 41.825 133.725 41.945 133.835 ;
        RECT 42.235 133.695 42.405 133.885 ;
        RECT 44.075 133.675 44.245 133.865 ;
        RECT 45.965 133.725 46.085 133.835 ;
        RECT 49.130 133.675 49.300 133.865 ;
        RECT 51.430 133.695 51.600 133.885 ;
        RECT 55.295 133.695 55.465 133.885 ;
        RECT 56.085 133.725 56.205 133.835 ;
        RECT 56.490 133.695 56.660 133.885 ;
        RECT 58.330 133.675 58.500 133.865 ;
        RECT 59.710 133.675 59.880 133.865 ;
        RECT 60.165 133.695 60.335 133.885 ;
        RECT 63.385 133.695 63.555 133.885 ;
        RECT 67.255 133.695 67.425 133.885 ;
        RECT 67.990 133.695 68.160 133.885 ;
        RECT 69.370 133.675 69.540 133.865 ;
        RECT 69.885 133.725 70.005 133.835 ;
        RECT 71.670 133.675 71.840 133.865 ;
        RECT 72.130 133.675 72.300 133.865 ;
        RECT 73.050 133.695 73.220 133.885 ;
        RECT 76.725 133.695 76.895 133.885 ;
        RECT 80.595 133.695 80.765 133.885 ;
        RECT 81.790 133.730 81.950 133.840 ;
        RECT 83.170 133.675 83.340 133.865 ;
        RECT 83.630 133.675 83.800 133.865 ;
        RECT 85.655 133.695 85.825 133.885 ;
        RECT 86.850 133.695 87.020 133.885 ;
        RECT 89.615 133.695 89.785 133.885 ;
        RECT 92.885 133.725 93.005 133.835 ;
        RECT 94.670 133.675 94.840 133.865 ;
        RECT 96.505 133.695 96.675 133.885 ;
        RECT 98.535 133.675 98.705 133.865 ;
        RECT 99.270 133.695 99.440 133.885 ;
        RECT 99.730 133.695 99.900 133.885 ;
        RECT 100.190 133.720 100.350 133.830 ;
        RECT 100.650 133.675 100.820 133.865 ;
        RECT 101.110 133.695 101.280 133.885 ;
        RECT 103.925 133.725 104.045 133.835 ;
        RECT 105.710 133.695 105.880 133.885 ;
        RECT 107.090 133.695 107.260 133.885 ;
        RECT 110.770 133.695 110.940 133.885 ;
        RECT 112.150 133.675 112.320 133.885 ;
        RECT 18.170 132.865 19.540 133.675 ;
        RECT 20.480 132.765 21.830 133.675 ;
        RECT 21.860 132.805 22.290 133.590 ;
        RECT 22.420 132.995 25.885 133.675 ;
        RECT 24.965 132.765 25.885 132.995 ;
        RECT 25.990 132.995 35.180 133.675 ;
        RECT 25.990 132.765 26.910 132.995 ;
        RECT 29.740 132.775 30.670 132.995 ;
        RECT 35.200 132.765 36.550 133.675 ;
        RECT 36.570 132.765 40.045 133.675 ;
        RECT 40.360 132.995 43.825 133.675 ;
        RECT 42.905 132.765 43.825 132.995 ;
        RECT 43.930 132.765 47.405 133.675 ;
        RECT 47.620 132.805 48.050 133.590 ;
        RECT 48.070 132.865 49.440 133.675 ;
        RECT 49.450 132.995 58.640 133.675 ;
        RECT 49.450 132.765 50.370 132.995 ;
        RECT 53.200 132.775 54.130 132.995 ;
        RECT 58.650 132.865 60.020 133.675 ;
        RECT 60.400 132.995 69.680 133.675 ;
        RECT 60.400 132.875 62.735 132.995 ;
        RECT 60.400 132.765 61.320 132.875 ;
        RECT 67.400 132.775 68.320 132.995 ;
        RECT 70.150 132.865 71.980 133.675 ;
        RECT 72.000 132.765 73.350 133.675 ;
        RECT 73.380 132.805 73.810 133.590 ;
        RECT 74.200 132.995 83.480 133.675 ;
        RECT 83.490 132.995 92.595 133.675 ;
        RECT 74.200 132.875 76.535 132.995 ;
        RECT 74.200 132.765 75.120 132.875 ;
        RECT 81.200 132.775 82.120 132.995 ;
        RECT 93.150 132.865 94.980 133.675 ;
        RECT 95.220 132.995 99.120 133.675 ;
        RECT 98.190 132.765 99.120 132.995 ;
        RECT 99.140 132.805 99.570 133.590 ;
        RECT 100.510 132.995 110.880 133.675 ;
        RECT 105.020 132.775 105.950 132.995 ;
        RECT 108.670 132.765 110.880 132.995 ;
        RECT 111.090 132.865 112.460 133.675 ;
      LAYER nwell ;
        RECT 17.975 129.645 112.655 132.475 ;
      LAYER pwell ;
        RECT 18.170 128.445 19.540 129.255 ;
        RECT 19.750 129.125 21.960 129.355 ;
        RECT 24.680 129.125 25.610 129.345 ;
        RECT 33.330 129.125 34.260 129.355 ;
        RECT 19.750 128.445 30.120 129.125 ;
        RECT 30.360 128.445 34.260 129.125 ;
        RECT 34.740 128.530 35.170 129.315 ;
        RECT 35.735 128.445 44.840 129.125 ;
        RECT 45.330 128.445 56.340 129.355 ;
        RECT 56.350 128.445 59.100 129.255 ;
        RECT 59.120 128.445 60.470 129.355 ;
        RECT 60.500 128.530 60.930 129.315 ;
        RECT 64.150 129.125 65.080 129.355 ;
        RECT 61.180 128.445 65.080 129.125 ;
        RECT 65.090 128.445 66.920 129.255 ;
        RECT 66.930 129.125 67.850 129.355 ;
        RECT 70.680 129.125 71.610 129.345 ;
        RECT 76.960 129.245 77.880 129.355 ;
        RECT 76.960 129.125 79.295 129.245 ;
        RECT 83.960 129.125 84.880 129.345 ;
        RECT 66.930 128.445 76.120 129.125 ;
        RECT 76.960 128.445 86.240 129.125 ;
        RECT 86.260 128.530 86.690 129.315 ;
        RECT 87.865 128.445 92.680 129.125 ;
        RECT 92.700 128.445 94.050 129.355 ;
        RECT 94.990 129.125 95.910 129.355 ;
        RECT 98.740 129.125 99.670 129.345 ;
        RECT 94.990 128.445 104.180 129.125 ;
        RECT 104.190 128.445 105.560 129.255 ;
        RECT 105.580 128.445 106.930 129.355 ;
        RECT 107.410 128.445 111.080 129.255 ;
        RECT 111.090 128.445 112.460 129.255 ;
        RECT 18.310 128.235 18.480 128.445 ;
        RECT 20.150 128.280 20.310 128.390 ;
        RECT 21.530 128.235 21.700 128.425 ;
        RECT 29.810 128.255 29.980 128.445 ;
        RECT 32.570 128.235 32.740 128.425 ;
        RECT 33.490 128.280 33.650 128.390 ;
        RECT 33.675 128.255 33.845 128.445 ;
        RECT 33.960 128.235 34.130 128.425 ;
        RECT 34.465 128.285 34.585 128.395 ;
        RECT 35.335 128.235 35.505 128.425 ;
        RECT 39.470 128.280 39.630 128.390 ;
        RECT 39.935 128.235 40.105 128.425 ;
        RECT 44.530 128.255 44.700 128.445 ;
        RECT 45.045 128.285 45.165 128.395 ;
        RECT 47.015 128.235 47.185 128.425 ;
        RECT 48.210 128.235 48.380 128.425 ;
        RECT 50.970 128.280 51.130 128.390 ;
        RECT 51.430 128.235 51.600 128.425 ;
        RECT 56.025 128.255 56.195 128.445 ;
        RECT 56.215 128.235 56.385 128.425 ;
        RECT 58.790 128.255 58.960 128.445 ;
        RECT 59.250 128.255 59.420 128.445 ;
        RECT 64.495 128.255 64.665 128.445 ;
        RECT 66.150 128.235 66.320 128.425 ;
        RECT 66.610 128.255 66.780 128.445 ;
        RECT 67.530 128.235 67.700 128.425 ;
        RECT 68.910 128.235 69.080 128.425 ;
        RECT 72.775 128.235 72.945 128.425 ;
        RECT 75.810 128.255 75.980 128.445 ;
        RECT 76.325 128.285 76.445 128.395 ;
        RECT 82.710 128.235 82.880 128.425 ;
        RECT 83.225 128.285 83.345 128.395 ;
        RECT 85.930 128.255 86.100 128.445 ;
        RECT 87.310 128.290 87.470 128.400 ;
        RECT 92.370 128.255 92.540 128.445 ;
        RECT 92.830 128.235 93.000 128.445 ;
        RECT 93.295 128.235 93.465 128.425 ;
        RECT 94.670 128.290 94.830 128.400 ;
        RECT 97.430 128.280 97.590 128.390 ;
        RECT 98.810 128.235 98.980 128.425 ;
        RECT 99.730 128.235 99.900 128.425 ;
        RECT 103.410 128.235 103.580 128.425 ;
        RECT 103.870 128.255 104.040 128.445 ;
        RECT 105.250 128.255 105.420 128.445 ;
        RECT 105.710 128.255 105.880 128.445 ;
        RECT 107.090 128.395 107.260 128.425 ;
        RECT 107.090 128.285 107.265 128.395 ;
        RECT 107.090 128.235 107.260 128.285 ;
        RECT 110.770 128.235 110.940 128.445 ;
        RECT 112.150 128.235 112.320 128.445 ;
        RECT 18.170 127.425 19.540 128.235 ;
        RECT 20.480 127.325 21.830 128.235 ;
        RECT 21.860 127.365 22.290 128.150 ;
        RECT 22.510 127.555 32.880 128.235 ;
        RECT 22.510 127.325 24.720 127.555 ;
        RECT 27.440 127.335 28.370 127.555 ;
        RECT 33.810 127.455 35.180 128.235 ;
        RECT 35.190 127.325 38.665 128.235 ;
        RECT 39.790 127.325 43.265 128.235 ;
        RECT 43.700 127.555 47.600 128.235 ;
        RECT 46.670 127.325 47.600 127.555 ;
        RECT 47.620 127.365 48.050 128.150 ;
        RECT 48.120 127.325 50.310 128.235 ;
        RECT 51.300 127.325 52.650 128.235 ;
        RECT 52.900 127.555 56.800 128.235 ;
        RECT 55.870 127.325 56.800 127.555 ;
        RECT 57.180 127.555 66.460 128.235 ;
        RECT 57.180 127.435 59.515 127.555 ;
        RECT 57.180 127.325 58.100 127.435 ;
        RECT 64.180 127.335 65.100 127.555 ;
        RECT 66.470 127.425 67.840 128.235 ;
        RECT 67.860 127.325 69.210 128.235 ;
        RECT 69.460 127.555 73.360 128.235 ;
        RECT 72.430 127.325 73.360 127.555 ;
        RECT 73.380 127.365 73.810 128.150 ;
        RECT 73.915 127.555 83.020 128.235 ;
        RECT 83.860 127.555 93.140 128.235 ;
        RECT 83.860 127.435 86.195 127.555 ;
        RECT 83.860 127.325 84.780 127.435 ;
        RECT 90.860 127.335 91.780 127.555 ;
        RECT 93.150 127.325 96.625 128.235 ;
        RECT 97.760 127.325 99.110 128.235 ;
        RECT 99.140 127.365 99.570 128.150 ;
        RECT 99.700 127.555 103.165 128.235 ;
        RECT 103.270 127.555 106.010 128.235 ;
        RECT 102.245 127.325 103.165 127.555 ;
        RECT 106.030 127.425 107.400 128.235 ;
        RECT 107.410 127.425 111.080 128.235 ;
        RECT 111.090 127.425 112.460 128.235 ;
      LAYER nwell ;
        RECT 17.975 124.205 112.655 127.035 ;
      LAYER pwell ;
        RECT 18.170 123.005 19.540 123.815 ;
        RECT 19.550 123.005 21.380 123.815 ;
        RECT 21.400 123.005 22.750 123.915 ;
        RECT 28.185 123.685 29.105 123.915 ;
        RECT 22.780 123.005 25.520 123.685 ;
        RECT 25.640 123.005 29.105 123.685 ;
        RECT 29.210 123.005 30.580 123.815 ;
        RECT 33.790 123.685 34.720 123.915 ;
        RECT 30.820 123.005 34.720 123.685 ;
        RECT 34.740 123.090 35.170 123.875 ;
        RECT 35.190 123.715 36.135 123.915 ;
        RECT 35.190 123.035 37.940 123.715 ;
        RECT 37.950 123.685 38.870 123.915 ;
        RECT 41.700 123.685 42.630 123.905 ;
        RECT 35.190 123.005 36.135 123.035 ;
        RECT 18.310 122.795 18.480 123.005 ;
        RECT 19.745 122.845 19.865 122.955 ;
        RECT 21.070 122.815 21.240 123.005 ;
        RECT 21.530 122.795 21.700 123.005 ;
        RECT 23.370 122.795 23.540 122.985 ;
        RECT 24.750 122.795 24.920 122.985 ;
        RECT 25.210 122.815 25.380 123.005 ;
        RECT 25.670 122.815 25.840 123.005 ;
        RECT 26.130 122.795 26.300 122.985 ;
        RECT 29.805 122.795 29.975 122.985 ;
        RECT 30.270 122.795 30.440 123.005 ;
        RECT 34.135 122.815 34.305 123.005 ;
        RECT 37.625 122.815 37.795 123.035 ;
        RECT 37.950 123.005 47.140 123.685 ;
        RECT 47.150 123.005 56.255 123.685 ;
        RECT 57.005 123.005 60.480 123.915 ;
        RECT 60.500 123.090 60.930 123.875 ;
        RECT 60.950 123.005 64.425 123.915 ;
        RECT 65.090 123.005 67.840 123.815 ;
        RECT 71.050 123.685 71.980 123.915 ;
        RECT 73.350 123.685 74.270 123.905 ;
        RECT 80.350 123.805 81.270 123.915 ;
        RECT 78.935 123.685 81.270 123.805 ;
        RECT 85.310 123.685 86.240 123.915 ;
        RECT 68.080 123.005 71.980 123.685 ;
        RECT 71.990 123.005 81.270 123.685 ;
        RECT 82.340 123.005 86.240 123.685 ;
        RECT 86.260 123.090 86.690 123.875 ;
        RECT 87.825 123.005 91.300 123.915 ;
        RECT 91.310 123.005 93.140 123.815 ;
        RECT 95.805 123.685 96.725 123.915 ;
        RECT 93.260 123.005 96.725 123.685 ;
        RECT 96.830 123.685 97.750 123.915 ;
        RECT 100.580 123.685 101.510 123.905 ;
        RECT 96.830 123.005 106.020 123.685 ;
        RECT 106.030 123.005 107.400 123.815 ;
        RECT 107.410 123.005 111.080 123.815 ;
        RECT 111.090 123.005 112.460 123.815 ;
        RECT 39.525 122.845 39.645 122.955 ;
        RECT 39.930 122.795 40.100 122.985 ;
        RECT 46.830 122.815 47.000 123.005 ;
        RECT 47.015 122.795 47.185 122.985 ;
        RECT 47.290 122.815 47.460 123.005 ;
        RECT 48.265 122.845 48.385 122.955 ;
        RECT 49.590 122.795 49.760 122.985 ;
        RECT 53.455 122.795 53.625 122.985 ;
        RECT 54.650 122.840 54.810 122.950 ;
        RECT 55.110 122.795 55.280 122.985 ;
        RECT 56.545 122.845 56.665 122.955 ;
        RECT 59.250 122.840 59.410 122.950 ;
        RECT 59.715 122.795 59.885 122.985 ;
        RECT 60.165 122.815 60.335 123.005 ;
        RECT 61.095 122.815 61.265 123.005 ;
        RECT 63.390 122.795 63.560 122.985 ;
        RECT 64.825 122.845 64.945 122.955 ;
        RECT 67.345 122.795 67.515 122.985 ;
        RECT 67.530 122.815 67.700 123.005 ;
        RECT 71.265 122.845 71.385 122.955 ;
        RECT 71.395 122.815 71.565 123.005 ;
        RECT 72.130 122.815 72.300 123.005 ;
        RECT 73.050 122.815 73.220 122.985 ;
        RECT 73.970 122.795 74.140 122.985 ;
        RECT 78.570 122.795 78.740 122.985 ;
        RECT 79.030 122.795 79.200 122.985 ;
        RECT 81.845 122.845 81.965 122.955 ;
        RECT 82.710 122.795 82.880 122.985 ;
        RECT 83.175 122.795 83.345 122.985 ;
        RECT 85.655 122.815 85.825 123.005 ;
        RECT 86.855 122.795 87.025 122.985 ;
        RECT 87.310 122.850 87.470 122.960 ;
        RECT 90.985 122.815 91.155 123.005 ;
        RECT 92.830 122.815 93.000 123.005 ;
        RECT 93.290 122.815 93.460 123.005 ;
        RECT 94.665 122.795 94.835 122.985 ;
        RECT 98.535 122.795 98.705 122.985 ;
        RECT 99.730 122.795 99.900 122.985 ;
        RECT 103.410 122.795 103.580 122.985 ;
        RECT 105.250 122.840 105.410 122.950 ;
        RECT 105.710 122.815 105.880 123.005 ;
        RECT 107.090 122.815 107.260 123.005 ;
        RECT 110.770 122.795 110.940 123.005 ;
        RECT 112.150 122.795 112.320 123.005 ;
        RECT 18.170 121.985 19.540 122.795 ;
        RECT 20.010 121.985 21.840 122.795 ;
        RECT 21.860 121.925 22.290 122.710 ;
        RECT 22.310 121.985 23.680 122.795 ;
        RECT 23.700 121.885 25.050 122.795 ;
        RECT 25.070 121.985 26.440 122.795 ;
        RECT 26.645 121.885 30.120 122.795 ;
        RECT 30.130 122.115 39.320 122.795 ;
        RECT 39.900 122.115 43.365 122.795 ;
        RECT 43.700 122.115 47.600 122.795 ;
        RECT 34.640 121.895 35.570 122.115 ;
        RECT 38.400 121.885 39.320 122.115 ;
        RECT 42.445 121.885 43.365 122.115 ;
        RECT 46.670 121.885 47.600 122.115 ;
        RECT 47.620 121.925 48.050 122.710 ;
        RECT 48.540 121.885 49.890 122.795 ;
        RECT 50.140 122.115 54.040 122.795 ;
        RECT 55.080 122.115 58.545 122.795 ;
        RECT 53.110 121.885 54.040 122.115 ;
        RECT 57.625 121.885 58.545 122.115 ;
        RECT 59.570 121.885 63.045 122.795 ;
        RECT 63.360 122.115 66.825 122.795 ;
        RECT 65.905 121.885 66.825 122.115 ;
        RECT 66.930 122.115 70.830 122.795 ;
        RECT 71.530 122.115 72.895 122.795 ;
        RECT 66.930 121.885 67.860 122.115 ;
        RECT 73.380 121.925 73.810 122.710 ;
        RECT 73.840 121.885 75.190 122.795 ;
        RECT 75.305 122.115 78.770 122.795 ;
        RECT 78.890 122.115 81.630 122.795 ;
        RECT 75.305 121.885 76.225 122.115 ;
        RECT 81.650 121.985 83.020 122.795 ;
        RECT 83.030 121.885 86.505 122.795 ;
        RECT 86.710 121.885 90.185 122.795 ;
        RECT 91.505 121.885 94.980 122.795 ;
        RECT 95.220 122.115 99.120 122.795 ;
        RECT 98.190 121.885 99.120 122.115 ;
        RECT 99.140 121.925 99.570 122.710 ;
        RECT 99.700 122.115 103.165 122.795 ;
        RECT 102.245 121.885 103.165 122.115 ;
        RECT 103.280 121.885 104.630 122.795 ;
        RECT 105.570 121.985 111.080 122.795 ;
        RECT 111.090 121.985 112.460 122.795 ;
      LAYER nwell ;
        RECT 17.975 118.765 112.655 121.595 ;
      LAYER pwell ;
        RECT 18.170 117.565 19.540 118.375 ;
        RECT 19.750 118.245 21.960 118.475 ;
        RECT 24.680 118.245 25.610 118.465 ;
        RECT 31.145 118.245 32.065 118.475 ;
        RECT 19.750 117.565 30.120 118.245 ;
        RECT 31.145 117.565 34.610 118.245 ;
        RECT 34.740 117.650 35.170 118.435 ;
        RECT 35.190 117.565 38.665 118.475 ;
        RECT 43.380 118.245 44.310 118.465 ;
        RECT 47.140 118.245 48.060 118.475 ;
        RECT 38.870 117.565 48.060 118.245 ;
        RECT 48.070 118.245 48.990 118.475 ;
        RECT 51.820 118.245 52.750 118.465 ;
        RECT 57.730 118.275 58.675 118.475 ;
        RECT 48.070 117.565 57.260 118.245 ;
        RECT 57.730 117.595 60.480 118.275 ;
        RECT 60.500 117.650 60.930 118.435 ;
        RECT 61.150 118.385 62.100 118.475 ;
        RECT 57.730 117.565 58.675 117.595 ;
        RECT 18.310 117.355 18.480 117.565 ;
        RECT 19.745 117.405 19.865 117.515 ;
        RECT 21.530 117.355 21.700 117.545 ;
        RECT 22.505 117.405 22.625 117.515 ;
        RECT 29.810 117.375 29.980 117.565 ;
        RECT 30.730 117.410 30.890 117.520 ;
        RECT 33.030 117.355 33.200 117.545 ;
        RECT 34.410 117.375 34.580 117.565 ;
        RECT 35.335 117.375 35.505 117.565 ;
        RECT 35.790 117.355 35.960 117.545 ;
        RECT 36.250 117.355 36.420 117.545 ;
        RECT 39.010 117.375 39.180 117.565 ;
        RECT 39.930 117.355 40.100 117.545 ;
        RECT 46.830 117.355 47.000 117.545 ;
        RECT 47.345 117.405 47.465 117.515 ;
        RECT 48.215 117.355 48.385 117.545 ;
        RECT 52.810 117.355 52.980 117.545 ;
        RECT 56.490 117.355 56.660 117.545 ;
        RECT 56.950 117.355 57.120 117.565 ;
        RECT 57.465 117.405 57.585 117.515 ;
        RECT 60.165 117.375 60.335 117.595 ;
        RECT 61.150 117.565 63.080 118.385 ;
        RECT 63.250 118.275 64.195 118.475 ;
        RECT 63.250 117.595 66.000 118.275 ;
        RECT 70.520 118.245 71.450 118.465 ;
        RECT 74.280 118.245 75.200 118.475 ;
        RECT 78.410 118.245 79.340 118.475 ;
        RECT 63.250 117.565 64.195 117.595 ;
        RECT 62.930 117.545 63.080 117.565 ;
        RECT 62.930 117.375 63.100 117.545 ;
        RECT 65.685 117.375 65.855 117.595 ;
        RECT 66.010 117.565 75.200 118.245 ;
        RECT 75.440 117.565 79.340 118.245 ;
        RECT 79.810 117.565 82.550 118.245 ;
        RECT 82.570 117.565 86.045 118.475 ;
        RECT 86.260 117.650 86.690 118.435 ;
        RECT 86.720 117.565 88.070 118.475 ;
        RECT 88.090 117.565 91.565 118.475 ;
        RECT 94.970 118.245 95.900 118.475 ;
        RECT 100.420 118.245 101.350 118.465 ;
        RECT 104.180 118.245 105.100 118.475 ;
        RECT 92.000 117.565 95.900 118.245 ;
        RECT 95.910 117.565 105.100 118.245 ;
        RECT 105.570 117.565 111.080 118.375 ;
        RECT 111.090 117.565 112.460 118.375 ;
        RECT 66.150 117.375 66.320 117.565 ;
        RECT 66.665 117.405 66.785 117.515 ;
        RECT 67.075 117.355 67.245 117.545 ;
        RECT 70.750 117.355 70.920 117.545 ;
        RECT 72.130 117.355 72.300 117.545 ;
        RECT 74.430 117.400 74.590 117.510 ;
        RECT 74.890 117.355 75.060 117.545 ;
        RECT 78.755 117.375 78.925 117.565 ;
        RECT 79.545 117.405 79.665 117.515 ;
        RECT 79.950 117.375 80.120 117.565 ;
        RECT 82.715 117.375 82.885 117.565 ;
        RECT 84.550 117.400 84.710 117.510 ;
        RECT 85.010 117.355 85.180 117.545 ;
        RECT 86.850 117.375 87.020 117.565 ;
        RECT 88.235 117.375 88.405 117.565 ;
        RECT 89.610 117.355 89.780 117.545 ;
        RECT 18.170 116.545 19.540 117.355 ;
        RECT 20.010 116.545 21.840 117.355 ;
        RECT 21.860 116.485 22.290 117.270 ;
        RECT 22.970 116.675 33.340 117.355 ;
        RECT 33.360 116.675 36.100 117.355 ;
        RECT 36.220 116.675 39.685 117.355 ;
        RECT 39.900 116.675 43.365 117.355 ;
        RECT 22.970 116.445 25.180 116.675 ;
        RECT 27.900 116.455 28.830 116.675 ;
        RECT 38.765 116.445 39.685 116.675 ;
        RECT 42.445 116.445 43.365 116.675 ;
        RECT 43.565 116.675 47.030 117.355 ;
        RECT 43.565 116.445 44.485 116.675 ;
        RECT 47.620 116.485 48.050 117.270 ;
        RECT 48.070 116.445 51.545 117.355 ;
        RECT 51.760 116.445 53.110 117.355 ;
        RECT 53.130 116.545 56.800 117.355 ;
        RECT 56.810 116.675 66.090 117.355 ;
        RECT 58.170 116.455 59.090 116.675 ;
        RECT 63.755 116.555 66.090 116.675 ;
        RECT 65.170 116.445 66.090 116.555 ;
        RECT 66.930 116.445 70.405 117.355 ;
        RECT 70.620 116.445 71.970 117.355 ;
        RECT 72.000 116.445 73.350 117.355 ;
        RECT 73.380 116.485 73.810 117.270 ;
        RECT 74.750 116.675 83.940 117.355 ;
        RECT 84.980 116.675 88.445 117.355 ;
        RECT 79.260 116.455 80.190 116.675 ;
        RECT 83.020 116.445 83.940 116.675 ;
        RECT 87.525 116.445 88.445 116.675 ;
        RECT 88.550 116.545 89.920 117.355 ;
        RECT 90.075 117.325 90.245 117.545 ;
        RECT 92.830 117.355 93.000 117.545 ;
        RECT 95.315 117.375 95.485 117.565 ;
        RECT 96.050 117.375 96.220 117.565 ;
        RECT 91.735 117.325 92.680 117.355 ;
        RECT 89.930 116.645 92.680 117.325 ;
        RECT 92.800 116.675 96.265 117.355 ;
        RECT 96.515 117.325 96.685 117.545 ;
        RECT 101.570 117.375 101.740 117.545 ;
        RECT 103.870 117.375 104.040 117.545 ;
        RECT 105.250 117.515 105.420 117.545 ;
        RECT 105.250 117.405 105.425 117.515 ;
        RECT 101.570 117.355 101.720 117.375 ;
        RECT 103.870 117.355 104.020 117.375 ;
        RECT 105.250 117.355 105.420 117.405 ;
        RECT 110.770 117.355 110.940 117.565 ;
        RECT 112.150 117.355 112.320 117.565 ;
        RECT 98.175 117.325 99.120 117.355 ;
        RECT 91.735 116.445 92.680 116.645 ;
        RECT 95.345 116.445 96.265 116.675 ;
        RECT 96.370 116.645 99.120 117.325 ;
        RECT 98.175 116.445 99.120 116.645 ;
        RECT 99.140 116.485 99.570 117.270 ;
        RECT 99.790 116.535 101.720 117.355 ;
        RECT 102.090 116.535 104.020 117.355 ;
        RECT 99.790 116.445 100.740 116.535 ;
        RECT 102.090 116.445 103.040 116.535 ;
        RECT 104.200 116.445 105.550 117.355 ;
        RECT 105.570 116.545 111.080 117.355 ;
        RECT 111.090 116.545 112.460 117.355 ;
      LAYER nwell ;
        RECT 17.975 113.325 112.655 116.155 ;
      LAYER pwell ;
        RECT 18.170 112.125 19.540 112.935 ;
        RECT 20.470 112.125 25.980 112.935 ;
        RECT 26.000 112.125 27.350 113.035 ;
        RECT 28.510 112.945 29.460 113.035 ;
        RECT 30.810 112.945 31.760 113.035 ;
        RECT 27.530 112.125 29.460 112.945 ;
        RECT 29.830 112.125 31.760 112.945 ;
        RECT 31.970 112.835 32.915 113.035 ;
        RECT 31.970 112.155 34.720 112.835 ;
        RECT 34.740 112.210 35.170 112.995 ;
        RECT 31.970 112.125 32.915 112.155 ;
        RECT 18.310 111.915 18.480 112.125 ;
        RECT 19.745 111.965 19.865 112.075 ;
        RECT 20.150 111.970 20.310 112.080 ;
        RECT 21.530 111.915 21.700 112.105 ;
        RECT 24.750 111.915 24.920 112.105 ;
        RECT 25.670 111.935 25.840 112.125 ;
        RECT 26.130 111.935 26.300 112.125 ;
        RECT 27.530 112.105 27.680 112.125 ;
        RECT 29.830 112.105 29.980 112.125 ;
        RECT 27.510 111.935 27.680 112.105 ;
        RECT 29.810 111.935 29.980 112.105 ;
        RECT 30.270 111.915 30.440 112.105 ;
        RECT 30.730 111.915 30.900 112.105 ;
        RECT 18.170 111.105 19.540 111.915 ;
        RECT 20.010 111.105 21.840 111.915 ;
        RECT 21.860 111.045 22.290 111.830 ;
        RECT 22.310 111.105 25.060 111.915 ;
        RECT 25.070 111.105 30.580 111.915 ;
        RECT 30.600 111.005 31.950 111.915 ;
        RECT 31.970 111.885 32.915 111.915 ;
        RECT 34.405 111.885 34.575 112.155 ;
        RECT 35.190 112.125 37.020 112.805 ;
        RECT 37.030 112.125 40.505 113.035 ;
        RECT 43.910 112.805 44.840 113.035 ;
        RECT 40.940 112.125 44.840 112.805 ;
        RECT 45.510 112.945 46.460 113.035 ;
        RECT 45.510 112.125 47.440 112.945 ;
        RECT 47.610 112.125 49.440 112.935 ;
        RECT 49.450 112.125 54.960 112.935 ;
        RECT 54.980 112.125 56.330 113.035 ;
        RECT 59.550 112.805 60.480 113.035 ;
        RECT 56.580 112.125 60.480 112.805 ;
        RECT 60.500 112.210 60.930 112.995 ;
        RECT 67.590 112.945 68.540 113.035 ;
        RECT 71.290 112.945 72.240 113.035 ;
        RECT 61.410 112.125 63.240 112.805 ;
        RECT 63.710 112.125 67.380 112.935 ;
        RECT 67.590 112.125 69.520 112.945 ;
        RECT 35.330 111.935 35.500 112.125 ;
        RECT 37.175 112.105 37.345 112.125 ;
        RECT 37.165 111.935 37.345 112.105 ;
        RECT 44.255 111.935 44.425 112.125 ;
        RECT 47.290 112.105 47.440 112.125 ;
        RECT 45.045 111.965 45.165 112.075 ;
        RECT 34.730 111.885 35.675 111.915 ;
        RECT 37.165 111.885 37.335 111.935 ;
        RECT 46.830 111.915 47.000 112.105 ;
        RECT 47.290 112.075 47.460 112.105 ;
        RECT 47.290 111.965 47.465 112.075 ;
        RECT 47.290 111.935 47.460 111.965 ;
        RECT 49.130 111.915 49.300 112.125 ;
        RECT 49.645 111.965 49.765 112.075 ;
        RECT 53.270 111.915 53.440 112.105 ;
        RECT 54.650 111.935 54.820 112.125 ;
        RECT 55.110 111.935 55.280 112.125 ;
        RECT 59.895 111.935 60.065 112.125 ;
        RECT 61.145 111.965 61.265 112.075 ;
        RECT 61.550 111.935 61.720 112.125 ;
        RECT 62.930 111.915 63.100 112.105 ;
        RECT 63.390 112.075 63.560 112.105 ;
        RECT 63.390 111.965 63.565 112.075 ;
        RECT 64.825 111.965 64.945 112.075 ;
        RECT 63.390 111.915 63.560 111.965 ;
        RECT 67.070 111.935 67.240 112.125 ;
        RECT 69.370 112.105 69.520 112.125 ;
        RECT 70.310 112.125 72.240 112.945 ;
        RECT 75.105 112.805 76.025 113.035 ;
        RECT 72.560 112.125 76.025 112.805 ;
        RECT 76.225 112.805 77.145 113.035 ;
        RECT 81.615 112.835 82.560 113.035 ;
        RECT 76.225 112.125 79.690 112.805 ;
        RECT 79.810 112.155 82.560 112.835 ;
        RECT 70.310 112.105 70.460 112.125 ;
        RECT 67.530 111.915 67.700 112.105 ;
        RECT 68.910 111.915 69.080 112.105 ;
        RECT 69.370 111.935 69.540 112.105 ;
        RECT 69.885 111.965 70.005 112.075 ;
        RECT 70.290 111.935 70.460 112.105 ;
        RECT 72.590 111.935 72.760 112.125 ;
        RECT 72.775 111.915 72.945 112.105 ;
        RECT 77.375 111.915 77.545 112.105 ;
        RECT 78.165 111.965 78.285 112.075 ;
        RECT 78.570 111.935 78.740 112.105 ;
        RECT 79.490 111.935 79.660 112.125 ;
        RECT 79.955 111.935 80.125 112.155 ;
        RECT 81.615 112.125 82.560 112.155 ;
        RECT 83.490 112.835 84.435 113.035 ;
        RECT 83.490 112.155 86.240 112.835 ;
        RECT 86.260 112.210 86.690 112.995 ;
        RECT 83.490 112.125 84.435 112.155 ;
        RECT 83.170 111.970 83.330 112.080 ;
        RECT 85.925 111.935 86.095 112.155 ;
        RECT 86.720 112.125 88.070 113.035 ;
        RECT 91.290 112.805 92.220 113.035 ;
        RECT 88.320 112.125 92.220 112.805 ;
        RECT 92.600 112.925 93.520 113.035 ;
        RECT 92.600 112.805 94.935 112.925 ;
        RECT 99.600 112.805 100.520 113.025 ;
        RECT 92.600 112.125 101.880 112.805 ;
        RECT 101.890 112.125 105.560 112.935 ;
        RECT 105.570 112.125 111.080 112.935 ;
        RECT 111.090 112.125 112.460 112.935 ;
        RECT 87.770 111.935 87.940 112.125 ;
        RECT 78.590 111.915 78.740 111.935 ;
        RECT 90.070 111.915 90.240 112.105 ;
        RECT 90.805 111.915 90.975 112.105 ;
        RECT 91.635 111.935 91.805 112.125 ;
        RECT 98.075 111.915 98.245 112.105 ;
        RECT 98.865 111.965 98.985 112.075 ;
        RECT 99.785 111.965 99.905 112.075 ;
        RECT 101.570 111.935 101.740 112.125 ;
        RECT 105.250 111.915 105.420 112.125 ;
        RECT 110.770 111.915 110.940 112.125 ;
        RECT 112.150 111.915 112.320 112.125 ;
        RECT 31.970 111.205 34.720 111.885 ;
        RECT 34.730 111.205 37.480 111.885 ;
        RECT 37.860 111.235 47.140 111.915 ;
        RECT 31.970 111.005 32.915 111.205 ;
        RECT 34.730 111.005 35.675 111.205 ;
        RECT 37.860 111.115 40.195 111.235 ;
        RECT 37.860 111.005 38.780 111.115 ;
        RECT 44.860 111.015 45.780 111.235 ;
        RECT 47.620 111.045 48.050 111.830 ;
        RECT 48.080 111.005 49.430 111.915 ;
        RECT 49.910 111.105 53.580 111.915 ;
        RECT 53.960 111.235 63.240 111.915 ;
        RECT 53.960 111.115 56.295 111.235 ;
        RECT 53.960 111.005 54.880 111.115 ;
        RECT 60.960 111.015 61.880 111.235 ;
        RECT 63.260 111.005 64.610 111.915 ;
        RECT 65.090 111.105 67.840 111.915 ;
        RECT 67.860 111.005 69.210 111.915 ;
        RECT 69.460 111.235 73.360 111.915 ;
        RECT 72.430 111.005 73.360 111.235 ;
        RECT 73.380 111.045 73.810 111.830 ;
        RECT 74.060 111.235 77.960 111.915 ;
        RECT 77.030 111.005 77.960 111.235 ;
        RECT 78.590 111.095 80.520 111.915 ;
        RECT 79.570 111.005 80.520 111.095 ;
        RECT 81.100 111.235 90.380 111.915 ;
        RECT 90.390 111.235 94.290 111.915 ;
        RECT 94.760 111.235 98.660 111.915 ;
        RECT 81.100 111.115 83.435 111.235 ;
        RECT 81.100 111.005 82.020 111.115 ;
        RECT 88.100 111.015 89.020 111.235 ;
        RECT 90.390 111.005 91.320 111.235 ;
        RECT 97.730 111.005 98.660 111.235 ;
        RECT 99.140 111.045 99.570 111.830 ;
        RECT 100.050 111.105 105.560 111.915 ;
        RECT 105.570 111.105 111.080 111.915 ;
        RECT 111.090 111.105 112.460 111.915 ;
      LAYER nwell ;
        RECT 17.975 107.885 112.655 110.715 ;
      LAYER pwell ;
        RECT 18.170 106.685 19.540 107.495 ;
        RECT 20.010 106.685 25.520 107.495 ;
        RECT 25.530 106.685 31.040 107.495 ;
        RECT 31.060 106.685 32.410 107.595 ;
        RECT 32.630 107.505 33.580 107.595 ;
        RECT 32.630 106.685 34.560 107.505 ;
        RECT 34.740 106.770 35.170 107.555 ;
        RECT 39.310 107.365 40.240 107.595 ;
        RECT 43.450 107.365 44.380 107.595 ;
        RECT 36.340 106.685 40.240 107.365 ;
        RECT 40.480 106.685 44.380 107.365 ;
        RECT 44.760 107.485 45.680 107.595 ;
        RECT 44.760 107.365 47.095 107.485 ;
        RECT 51.760 107.365 52.680 107.585 ;
        RECT 44.760 106.685 54.040 107.365 ;
        RECT 54.510 106.685 56.340 107.495 ;
        RECT 59.550 107.365 60.480 107.595 ;
        RECT 56.580 106.685 60.480 107.365 ;
        RECT 60.500 106.770 60.930 107.555 ;
        RECT 61.435 107.365 62.780 107.595 ;
        RECT 60.950 106.685 62.780 107.365 ;
        RECT 62.790 106.685 65.540 107.495 ;
        RECT 65.920 107.485 66.840 107.595 ;
        RECT 65.920 107.365 68.255 107.485 ;
        RECT 72.920 107.365 73.840 107.585 ;
        RECT 76.570 107.365 77.490 107.585 ;
        RECT 83.570 107.485 84.490 107.595 ;
        RECT 82.155 107.365 84.490 107.485 ;
        RECT 65.920 106.685 75.200 107.365 ;
        RECT 75.210 106.685 84.490 107.365 ;
        RECT 84.880 106.685 86.230 107.595 ;
        RECT 86.260 106.770 86.690 107.555 ;
        RECT 86.710 106.685 89.450 107.365 ;
        RECT 89.480 106.685 90.830 107.595 ;
        RECT 92.210 107.365 93.130 107.585 ;
        RECT 99.210 107.485 100.130 107.595 ;
        RECT 97.795 107.365 100.130 107.485 ;
        RECT 90.850 106.685 100.130 107.365 ;
        RECT 100.520 106.685 101.870 107.595 ;
        RECT 101.890 106.685 105.560 107.495 ;
        RECT 105.570 106.685 111.080 107.495 ;
        RECT 111.090 106.685 112.460 107.495 ;
        RECT 18.310 106.475 18.480 106.685 ;
        RECT 19.745 106.525 19.865 106.635 ;
        RECT 21.530 106.475 21.700 106.665 ;
        RECT 22.910 106.520 23.070 106.630 ;
        RECT 25.210 106.495 25.380 106.685 ;
        RECT 26.590 106.475 26.760 106.665 ;
        RECT 30.730 106.495 30.900 106.685 ;
        RECT 31.190 106.495 31.360 106.685 ;
        RECT 34.410 106.665 34.560 106.685 ;
        RECT 32.110 106.475 32.280 106.665 ;
        RECT 34.410 106.495 34.580 106.665 ;
        RECT 35.790 106.530 35.950 106.640 ;
        RECT 37.630 106.475 37.800 106.665 ;
        RECT 39.655 106.495 39.825 106.685 ;
        RECT 43.795 106.495 43.965 106.685 ;
        RECT 47.290 106.475 47.460 106.665 ;
        RECT 49.130 106.475 49.300 106.665 ;
        RECT 53.730 106.495 53.900 106.685 ;
        RECT 54.245 106.525 54.365 106.635 ;
        RECT 56.030 106.495 56.200 106.685 ;
        RECT 59.710 106.475 59.880 106.665 ;
        RECT 59.895 106.495 60.065 106.685 ;
        RECT 61.090 106.495 61.260 106.685 ;
        RECT 65.230 106.495 65.400 106.685 ;
        RECT 70.290 106.475 70.460 106.665 ;
        RECT 73.050 106.475 73.220 106.665 ;
        RECT 74.025 106.525 74.145 106.635 ;
        RECT 74.430 106.475 74.600 106.665 ;
        RECT 74.890 106.495 75.060 106.685 ;
        RECT 75.350 106.495 75.520 106.685 ;
        RECT 85.930 106.475 86.100 106.685 ;
        RECT 86.850 106.495 87.020 106.685 ;
        RECT 89.610 106.495 89.780 106.685 ;
        RECT 90.990 106.495 91.160 106.685 ;
        RECT 96.510 106.475 96.680 106.665 ;
        RECT 97.025 106.525 97.145 106.635 ;
        RECT 98.810 106.475 98.980 106.665 ;
        RECT 99.785 106.525 99.905 106.635 ;
        RECT 101.570 106.495 101.740 106.685 ;
        RECT 105.250 106.475 105.420 106.685 ;
        RECT 110.770 106.475 110.940 106.685 ;
        RECT 112.150 106.475 112.320 106.685 ;
        RECT 18.170 105.665 19.540 106.475 ;
        RECT 20.010 105.665 21.840 106.475 ;
        RECT 21.860 105.605 22.290 106.390 ;
        RECT 23.230 105.665 26.900 106.475 ;
        RECT 26.910 105.665 32.420 106.475 ;
        RECT 32.430 105.665 37.940 106.475 ;
        RECT 38.320 105.795 47.600 106.475 ;
        RECT 38.320 105.675 40.655 105.795 ;
        RECT 38.320 105.565 39.240 105.675 ;
        RECT 45.320 105.575 46.240 105.795 ;
        RECT 47.620 105.605 48.050 106.390 ;
        RECT 48.070 105.665 49.440 106.475 ;
        RECT 49.650 105.795 60.020 106.475 ;
        RECT 60.230 105.795 70.600 106.475 ;
        RECT 49.650 105.565 51.860 105.795 ;
        RECT 54.580 105.575 55.510 105.795 ;
        RECT 60.230 105.565 62.440 105.795 ;
        RECT 65.160 105.575 66.090 105.795 ;
        RECT 70.610 105.665 73.360 106.475 ;
        RECT 73.380 105.605 73.810 106.390 ;
        RECT 74.300 105.565 75.650 106.475 ;
        RECT 75.870 105.795 86.240 106.475 ;
        RECT 86.450 105.795 96.820 106.475 ;
        RECT 75.870 105.565 78.080 105.795 ;
        RECT 80.800 105.575 81.730 105.795 ;
        RECT 86.450 105.565 88.660 105.795 ;
        RECT 91.380 105.575 92.310 105.795 ;
        RECT 97.290 105.665 99.120 106.475 ;
        RECT 99.140 105.605 99.570 106.390 ;
        RECT 100.050 105.665 105.560 106.475 ;
        RECT 105.570 105.665 111.080 106.475 ;
        RECT 111.090 105.665 112.460 106.475 ;
      LAYER nwell ;
        RECT 17.975 102.445 112.655 105.275 ;
      LAYER pwell ;
        RECT 18.170 101.245 19.540 102.055 ;
        RECT 20.010 101.245 21.840 102.055 ;
        RECT 21.860 101.330 22.290 102.115 ;
        RECT 22.310 101.245 23.680 102.055 ;
        RECT 23.690 101.245 29.200 102.055 ;
        RECT 29.210 101.245 34.720 102.055 ;
        RECT 34.740 101.330 35.170 102.115 ;
        RECT 35.190 101.245 36.560 102.055 ;
        RECT 36.570 101.245 42.080 102.055 ;
        RECT 42.090 101.245 47.600 102.055 ;
        RECT 47.620 101.330 48.050 102.115 ;
        RECT 48.070 101.245 53.580 102.055 ;
        RECT 53.600 101.245 54.950 102.155 ;
        RECT 54.970 101.245 60.480 102.055 ;
        RECT 60.500 101.330 60.930 102.115 ;
        RECT 60.950 101.245 62.320 102.055 ;
        RECT 62.340 101.245 63.690 102.155 ;
        RECT 64.170 101.245 67.840 102.055 ;
        RECT 67.850 101.245 73.360 102.055 ;
        RECT 73.380 101.330 73.810 102.115 ;
        RECT 74.290 101.245 79.800 102.055 ;
        RECT 79.820 101.245 81.170 102.155 ;
        RECT 81.190 101.245 82.560 102.055 ;
        RECT 82.570 101.245 86.240 102.055 ;
        RECT 86.260 101.330 86.690 102.115 ;
        RECT 86.710 101.245 88.080 102.055 ;
        RECT 88.090 101.245 93.600 102.055 ;
        RECT 93.610 101.245 99.120 102.055 ;
        RECT 99.140 101.330 99.570 102.115 ;
        RECT 100.050 101.245 105.560 102.055 ;
        RECT 105.570 101.245 111.080 102.055 ;
        RECT 111.090 101.245 112.460 102.055 ;
        RECT 18.310 101.055 18.480 101.245 ;
        RECT 19.745 101.085 19.865 101.195 ;
        RECT 21.530 101.055 21.700 101.245 ;
        RECT 23.370 101.055 23.540 101.245 ;
        RECT 28.890 101.055 29.060 101.245 ;
        RECT 34.410 101.055 34.580 101.245 ;
        RECT 36.250 101.055 36.420 101.245 ;
        RECT 41.770 101.055 41.940 101.245 ;
        RECT 47.290 101.055 47.460 101.245 ;
        RECT 53.270 101.055 53.440 101.245 ;
        RECT 54.650 101.055 54.820 101.245 ;
        RECT 60.170 101.055 60.340 101.245 ;
        RECT 62.010 101.055 62.180 101.245 ;
        RECT 62.470 101.055 62.640 101.245 ;
        RECT 63.905 101.085 64.025 101.195 ;
        RECT 67.530 101.055 67.700 101.245 ;
        RECT 73.050 101.055 73.220 101.245 ;
        RECT 74.025 101.085 74.145 101.195 ;
        RECT 79.490 101.055 79.660 101.245 ;
        RECT 80.870 101.055 81.040 101.245 ;
        RECT 82.250 101.055 82.420 101.245 ;
        RECT 85.930 101.055 86.100 101.245 ;
        RECT 87.770 101.055 87.940 101.245 ;
        RECT 93.290 101.055 93.460 101.245 ;
        RECT 98.810 101.055 98.980 101.245 ;
        RECT 99.785 101.085 99.905 101.195 ;
        RECT 105.250 101.055 105.420 101.245 ;
        RECT 110.770 101.055 110.940 101.245 ;
        RECT 112.150 101.055 112.320 101.245 ;
      LAYER nwell ;
        RECT 20.485 54.580 29.875 66.420 ;
        RECT 31.685 54.590 41.075 66.430 ;
        RECT 42.905 54.560 52.295 66.400 ;
        RECT 54.155 54.540 63.545 66.380 ;
        RECT 65.375 54.530 74.765 66.370 ;
        RECT 76.615 54.520 86.005 66.360 ;
        RECT 87.865 54.530 97.255 66.370 ;
        RECT 99.145 54.520 108.535 66.360 ;
        RECT 110.415 54.520 119.805 66.360 ;
        RECT 121.665 54.520 131.055 66.360 ;
        RECT 132.415 54.490 139.375 66.330 ;
        RECT 20.655 49.020 23.115 53.210 ;
      LAYER pwell ;
        RECT 20.555 45.340 22.915 48.340 ;
      LAYER nwell ;
        RECT 24.735 45.940 29.125 53.130 ;
        RECT 31.855 49.030 34.315 53.220 ;
      LAYER pwell ;
        RECT 31.755 45.350 34.115 48.350 ;
      LAYER nwell ;
        RECT 35.935 45.950 40.325 53.140 ;
        RECT 43.075 49.000 45.535 53.190 ;
      LAYER pwell ;
        RECT 42.975 45.320 45.335 48.320 ;
      LAYER nwell ;
        RECT 47.155 45.920 51.545 53.110 ;
        RECT 54.325 48.980 56.785 53.170 ;
      LAYER pwell ;
        RECT 54.225 45.300 56.585 48.300 ;
      LAYER nwell ;
        RECT 58.405 45.900 62.795 53.090 ;
        RECT 65.545 48.970 68.005 53.160 ;
      LAYER pwell ;
        RECT 65.445 45.290 67.805 48.290 ;
      LAYER nwell ;
        RECT 69.625 45.890 74.015 53.080 ;
        RECT 76.785 48.960 79.245 53.150 ;
      LAYER pwell ;
        RECT 76.685 45.280 79.045 48.280 ;
      LAYER nwell ;
        RECT 80.865 45.880 85.255 53.070 ;
        RECT 88.035 48.970 90.495 53.160 ;
      LAYER pwell ;
        RECT 87.935 45.290 90.295 48.290 ;
      LAYER nwell ;
        RECT 92.115 45.890 96.505 53.080 ;
        RECT 99.315 48.960 101.775 53.150 ;
      LAYER pwell ;
        RECT 99.215 45.280 101.575 48.280 ;
      LAYER nwell ;
        RECT 103.395 45.880 107.785 53.070 ;
        RECT 110.585 48.960 113.045 53.150 ;
      LAYER pwell ;
        RECT 110.485 45.280 112.845 48.280 ;
      LAYER nwell ;
        RECT 114.665 45.880 119.055 53.070 ;
        RECT 121.835 48.960 124.295 53.150 ;
      LAYER pwell ;
        RECT 121.735 45.280 124.095 48.280 ;
      LAYER nwell ;
        RECT 125.915 45.880 130.305 53.070 ;
        RECT 19.615 32.280 24.005 39.470 ;
      LAYER pwell ;
        RECT 25.825 37.070 28.185 40.070 ;
      LAYER nwell ;
        RECT 25.625 32.200 28.085 36.390 ;
        RECT 30.895 32.280 35.285 39.470 ;
      LAYER pwell ;
        RECT 37.105 37.070 39.465 40.070 ;
      LAYER nwell ;
        RECT 36.905 32.200 39.365 36.390 ;
        RECT 42.185 32.260 46.575 39.450 ;
      LAYER pwell ;
        RECT 48.395 37.050 50.755 40.050 ;
      LAYER nwell ;
        RECT 48.195 32.180 50.655 36.370 ;
        RECT 53.405 32.260 57.795 39.450 ;
      LAYER pwell ;
        RECT 59.615 37.050 61.975 40.050 ;
      LAYER nwell ;
        RECT 59.415 32.180 61.875 36.370 ;
        RECT 64.605 32.260 68.995 39.450 ;
      LAYER pwell ;
        RECT 70.815 37.050 73.175 40.050 ;
      LAYER nwell ;
        RECT 70.615 32.180 73.075 36.370 ;
        RECT 75.895 32.250 80.285 39.440 ;
      LAYER pwell ;
        RECT 82.105 37.040 84.465 40.040 ;
      LAYER nwell ;
        RECT 81.905 32.170 84.365 36.360 ;
        RECT 87.135 32.270 91.525 39.460 ;
      LAYER pwell ;
        RECT 93.345 37.060 95.705 40.060 ;
      LAYER nwell ;
        RECT 93.145 32.190 95.605 36.380 ;
        RECT 98.345 32.290 102.735 39.480 ;
      LAYER pwell ;
        RECT 104.555 37.080 106.915 40.080 ;
      LAYER nwell ;
        RECT 104.355 32.210 106.815 36.400 ;
        RECT 109.545 32.330 113.935 39.520 ;
      LAYER pwell ;
        RECT 115.755 37.120 118.115 40.120 ;
      LAYER nwell ;
        RECT 115.555 32.250 118.015 36.440 ;
        RECT 120.755 32.350 125.145 39.540 ;
      LAYER pwell ;
        RECT 126.965 37.140 129.325 40.140 ;
      LAYER nwell ;
        RECT 126.765 32.270 129.225 36.460 ;
        RECT 18.865 18.990 28.255 30.830 ;
        RECT 30.145 18.990 39.535 30.830 ;
        RECT 41.435 18.970 50.825 30.810 ;
        RECT 52.655 18.970 62.045 30.810 ;
        RECT 63.855 18.970 73.245 30.810 ;
        RECT 75.145 18.960 84.535 30.800 ;
        RECT 86.385 18.980 95.775 30.820 ;
        RECT 97.595 19.000 106.985 30.840 ;
        RECT 108.795 19.040 118.185 30.880 ;
        RECT 120.005 19.060 129.395 30.900 ;
        RECT 131.725 19.030 138.685 30.870 ;
      LAYER li1 ;
        RECT 18.165 193.535 112.465 193.705 ;
        RECT 18.250 192.785 19.460 193.535 ;
        RECT 18.250 192.245 18.770 192.785 ;
        RECT 20.090 192.765 21.760 193.535 ;
        RECT 21.930 192.810 22.220 193.535 ;
        RECT 22.850 192.765 24.520 193.535 ;
        RECT 24.695 192.990 30.040 193.535 ;
        RECT 18.940 192.075 19.460 192.615 ;
        RECT 18.250 190.985 19.460 192.075 ;
        RECT 20.090 192.075 20.840 192.595 ;
        RECT 21.010 192.245 21.760 192.765 ;
        RECT 20.090 190.985 21.760 192.075 ;
        RECT 21.930 190.985 22.220 192.150 ;
        RECT 22.850 192.075 23.600 192.595 ;
        RECT 23.770 192.245 24.520 192.765 ;
        RECT 22.850 190.985 24.520 192.075 ;
        RECT 26.285 191.420 26.635 192.670 ;
        RECT 28.115 192.160 28.455 192.990 ;
        RECT 30.270 192.715 30.480 193.535 ;
        RECT 30.650 192.735 30.980 193.365 ;
        RECT 30.650 192.135 30.900 192.735 ;
        RECT 31.150 192.715 31.380 193.535 ;
        RECT 32.050 192.765 34.640 193.535 ;
        RECT 34.810 192.810 35.100 193.535 ;
        RECT 36.190 192.765 39.700 193.535 ;
        RECT 31.070 192.295 31.400 192.545 ;
        RECT 24.695 190.985 30.040 191.420 ;
        RECT 30.270 190.985 30.480 192.125 ;
        RECT 30.650 191.155 30.980 192.135 ;
        RECT 31.150 190.985 31.380 192.125 ;
        RECT 32.050 192.075 33.260 192.595 ;
        RECT 33.430 192.245 34.640 192.765 ;
        RECT 32.050 190.985 34.640 192.075 ;
        RECT 34.810 190.985 35.100 192.150 ;
        RECT 36.190 192.075 37.880 192.595 ;
        RECT 38.050 192.245 39.700 192.765 ;
        RECT 39.870 192.735 40.180 193.535 ;
        RECT 40.385 192.735 41.080 193.365 ;
        RECT 41.250 192.785 42.460 193.535 ;
        RECT 39.880 192.295 40.215 192.565 ;
        RECT 40.385 192.135 40.555 192.735 ;
        RECT 40.725 192.295 41.060 192.545 ;
        RECT 36.190 190.985 39.700 192.075 ;
        RECT 39.870 190.985 40.150 192.125 ;
        RECT 40.320 191.155 40.650 192.135 ;
        RECT 40.820 190.985 41.080 192.125 ;
        RECT 41.250 192.075 41.770 192.615 ;
        RECT 41.940 192.245 42.460 192.785 ;
        RECT 42.670 192.715 42.900 193.535 ;
        RECT 43.070 192.735 43.400 193.365 ;
        RECT 42.650 192.295 42.980 192.545 ;
        RECT 43.150 192.135 43.400 192.735 ;
        RECT 43.570 192.715 43.780 193.535 ;
        RECT 44.010 192.765 47.520 193.535 ;
        RECT 47.690 192.810 47.980 193.535 ;
        RECT 48.610 192.765 50.280 193.535 ;
        RECT 41.250 190.985 42.460 192.075 ;
        RECT 42.670 190.985 42.900 192.125 ;
        RECT 43.070 191.155 43.400 192.135 ;
        RECT 43.570 190.985 43.780 192.125 ;
        RECT 44.010 192.075 45.700 192.595 ;
        RECT 45.870 192.245 47.520 192.765 ;
        RECT 44.010 190.985 47.520 192.075 ;
        RECT 47.690 190.985 47.980 192.150 ;
        RECT 48.610 192.075 49.360 192.595 ;
        RECT 49.530 192.245 50.280 192.765 ;
        RECT 50.510 192.715 50.720 193.535 ;
        RECT 50.890 192.735 51.220 193.365 ;
        RECT 50.890 192.135 51.140 192.735 ;
        RECT 51.390 192.715 51.620 193.535 ;
        RECT 51.830 192.765 53.500 193.535 ;
        RECT 53.675 192.990 59.020 193.535 ;
        RECT 51.310 192.295 51.640 192.545 ;
        RECT 48.610 190.985 50.280 192.075 ;
        RECT 50.510 190.985 50.720 192.125 ;
        RECT 50.890 191.155 51.220 192.135 ;
        RECT 51.390 190.985 51.620 192.125 ;
        RECT 51.830 192.075 52.580 192.595 ;
        RECT 52.750 192.245 53.500 192.765 ;
        RECT 51.830 190.985 53.500 192.075 ;
        RECT 55.265 191.420 55.615 192.670 ;
        RECT 57.095 192.160 57.435 192.990 ;
        RECT 59.230 192.715 59.460 193.535 ;
        RECT 59.630 192.735 59.960 193.365 ;
        RECT 59.210 192.295 59.540 192.545 ;
        RECT 59.710 192.135 59.960 192.735 ;
        RECT 60.130 192.715 60.340 193.535 ;
        RECT 60.570 192.810 60.860 193.535 ;
        RECT 61.490 192.765 65.000 193.535 ;
        RECT 53.675 190.985 59.020 191.420 ;
        RECT 59.230 190.985 59.460 192.125 ;
        RECT 59.630 191.155 59.960 192.135 ;
        RECT 60.130 190.985 60.340 192.125 ;
        RECT 60.570 190.985 60.860 192.150 ;
        RECT 61.490 192.075 63.180 192.595 ;
        RECT 63.350 192.245 65.000 192.765 ;
        RECT 65.230 192.715 65.440 193.535 ;
        RECT 65.610 192.735 65.940 193.365 ;
        RECT 65.610 192.135 65.860 192.735 ;
        RECT 66.110 192.715 66.340 193.535 ;
        RECT 66.550 192.785 67.760 193.535 ;
        RECT 67.935 192.990 73.280 193.535 ;
        RECT 66.030 192.295 66.360 192.545 ;
        RECT 61.490 190.985 65.000 192.075 ;
        RECT 65.230 190.985 65.440 192.125 ;
        RECT 65.610 191.155 65.940 192.135 ;
        RECT 66.110 190.985 66.340 192.125 ;
        RECT 66.550 192.075 67.070 192.615 ;
        RECT 67.240 192.245 67.760 192.785 ;
        RECT 66.550 190.985 67.760 192.075 ;
        RECT 69.525 191.420 69.875 192.670 ;
        RECT 71.355 192.160 71.695 192.990 ;
        RECT 73.450 192.810 73.740 193.535 ;
        RECT 73.910 192.765 75.580 193.535 ;
        RECT 76.060 193.065 76.230 193.535 ;
        RECT 76.400 192.885 76.730 193.365 ;
        RECT 76.900 193.065 77.070 193.535 ;
        RECT 77.240 192.885 77.570 193.365 ;
        RECT 67.935 190.985 73.280 191.420 ;
        RECT 73.450 190.985 73.740 192.150 ;
        RECT 73.910 192.075 74.660 192.595 ;
        RECT 74.830 192.245 75.580 192.765 ;
        RECT 75.805 192.715 77.570 192.885 ;
        RECT 77.740 192.725 77.910 193.535 ;
        RECT 78.110 193.155 79.180 193.325 ;
        RECT 78.110 192.800 78.430 193.155 ;
        RECT 75.805 192.165 76.215 192.715 ;
        RECT 78.105 192.545 78.430 192.800 ;
        RECT 76.400 192.335 78.430 192.545 ;
        RECT 78.085 192.325 78.430 192.335 ;
        RECT 78.600 192.585 78.840 192.985 ;
        RECT 79.010 192.925 79.180 193.155 ;
        RECT 79.350 193.095 79.540 193.535 ;
        RECT 79.710 193.085 80.660 193.365 ;
        RECT 80.880 193.175 81.230 193.345 ;
        RECT 79.010 192.755 79.540 192.925 ;
        RECT 73.910 190.985 75.580 192.075 ;
        RECT 75.805 191.995 77.530 192.165 ;
        RECT 76.060 190.985 76.230 191.825 ;
        RECT 76.440 191.155 76.690 191.995 ;
        RECT 76.900 190.985 77.070 191.825 ;
        RECT 77.240 191.155 77.530 191.995 ;
        RECT 77.740 190.985 77.910 192.045 ;
        RECT 78.085 191.705 78.255 192.325 ;
        RECT 78.600 192.215 79.140 192.585 ;
        RECT 79.320 192.475 79.540 192.755 ;
        RECT 79.710 192.305 79.880 193.085 ;
        RECT 79.475 192.135 79.880 192.305 ;
        RECT 80.050 192.295 80.400 192.915 ;
        RECT 79.475 192.045 79.645 192.135 ;
        RECT 80.570 192.125 80.780 192.915 ;
        RECT 78.425 191.875 79.645 192.045 ;
        RECT 80.105 191.965 80.780 192.125 ;
        RECT 78.085 191.535 78.885 191.705 ;
        RECT 78.205 190.985 78.535 191.365 ;
        RECT 78.715 191.245 78.885 191.535 ;
        RECT 79.475 191.495 79.645 191.875 ;
        RECT 79.815 191.955 80.780 191.965 ;
        RECT 80.970 192.785 81.230 193.175 ;
        RECT 81.440 193.075 81.770 193.535 ;
        RECT 82.645 193.145 83.500 193.315 ;
        RECT 83.705 193.145 84.200 193.315 ;
        RECT 84.370 193.175 84.700 193.535 ;
        RECT 80.970 192.095 81.140 192.785 ;
        RECT 81.310 192.435 81.480 192.615 ;
        RECT 81.650 192.605 82.440 192.855 ;
        RECT 82.645 192.435 82.815 193.145 ;
        RECT 82.985 192.635 83.340 192.855 ;
        RECT 81.310 192.265 83.000 192.435 ;
        RECT 79.815 191.665 80.275 191.955 ;
        RECT 80.970 191.925 82.470 192.095 ;
        RECT 80.970 191.785 81.140 191.925 ;
        RECT 80.580 191.615 81.140 191.785 ;
        RECT 79.055 190.985 79.305 191.445 ;
        RECT 79.475 191.155 80.345 191.495 ;
        RECT 80.580 191.155 80.750 191.615 ;
        RECT 81.585 191.585 82.660 191.755 ;
        RECT 80.920 190.985 81.290 191.445 ;
        RECT 81.585 191.245 81.755 191.585 ;
        RECT 81.925 190.985 82.255 191.415 ;
        RECT 82.490 191.245 82.660 191.585 ;
        RECT 82.830 191.485 83.000 192.265 ;
        RECT 83.170 192.045 83.340 192.635 ;
        RECT 83.510 192.235 83.860 192.855 ;
        RECT 83.170 191.655 83.635 192.045 ;
        RECT 84.030 191.785 84.200 193.145 ;
        RECT 84.370 191.955 84.830 193.005 ;
        RECT 83.805 191.615 84.200 191.785 ;
        RECT 83.805 191.485 83.975 191.615 ;
        RECT 82.830 191.155 83.510 191.485 ;
        RECT 83.725 191.155 83.975 191.485 ;
        RECT 84.145 190.985 84.395 191.445 ;
        RECT 84.565 191.170 84.890 191.955 ;
        RECT 85.060 191.155 85.230 193.275 ;
        RECT 85.400 193.155 85.730 193.535 ;
        RECT 85.900 192.985 86.155 193.275 ;
        RECT 85.405 192.815 86.155 192.985 ;
        RECT 85.405 191.825 85.635 192.815 ;
        RECT 86.330 192.810 86.620 193.535 ;
        RECT 86.850 192.715 87.060 193.535 ;
        RECT 87.230 192.735 87.560 193.365 ;
        RECT 85.805 191.995 86.155 192.645 ;
        RECT 85.405 191.655 86.155 191.825 ;
        RECT 85.400 190.985 85.730 191.485 ;
        RECT 85.900 191.155 86.155 191.655 ;
        RECT 86.330 190.985 86.620 192.150 ;
        RECT 87.230 192.135 87.480 192.735 ;
        RECT 87.730 192.715 87.960 193.535 ;
        RECT 88.170 192.785 89.380 193.535 ;
        RECT 87.650 192.295 87.980 192.545 ;
        RECT 86.850 190.985 87.060 192.125 ;
        RECT 87.230 191.155 87.560 192.135 ;
        RECT 87.730 190.985 87.960 192.125 ;
        RECT 88.170 192.075 88.690 192.615 ;
        RECT 88.860 192.245 89.380 192.785 ;
        RECT 89.825 192.725 90.070 193.330 ;
        RECT 90.290 193.000 90.800 193.535 ;
        RECT 89.550 192.555 90.780 192.725 ;
        RECT 88.170 190.985 89.380 192.075 ;
        RECT 89.550 191.745 89.890 192.555 ;
        RECT 90.060 191.990 90.810 192.180 ;
        RECT 89.550 191.335 90.065 191.745 ;
        RECT 90.300 190.985 90.470 191.745 ;
        RECT 90.640 191.325 90.810 191.990 ;
        RECT 90.980 192.005 91.170 193.365 ;
        RECT 91.340 192.515 91.615 193.365 ;
        RECT 91.805 193.000 92.335 193.365 ;
        RECT 92.760 193.135 93.090 193.535 ;
        RECT 92.160 192.965 92.335 193.000 ;
        RECT 91.340 192.345 91.620 192.515 ;
        RECT 91.340 192.205 91.615 192.345 ;
        RECT 91.820 192.005 91.990 192.805 ;
        RECT 90.980 191.835 91.990 192.005 ;
        RECT 92.160 192.795 93.090 192.965 ;
        RECT 93.260 192.795 93.515 193.365 ;
        RECT 92.160 191.665 92.330 192.795 ;
        RECT 92.920 192.625 93.090 192.795 ;
        RECT 91.205 191.495 92.330 191.665 ;
        RECT 92.500 192.295 92.695 192.625 ;
        RECT 92.920 192.295 93.175 192.625 ;
        RECT 92.500 191.325 92.670 192.295 ;
        RECT 93.345 192.125 93.515 192.795 ;
        RECT 94.210 192.715 94.420 193.535 ;
        RECT 94.590 192.735 94.920 193.365 ;
        RECT 94.590 192.135 94.840 192.735 ;
        RECT 95.090 192.715 95.320 193.535 ;
        RECT 95.530 192.765 99.040 193.535 ;
        RECT 99.210 192.810 99.500 193.535 ;
        RECT 100.130 192.765 103.640 193.535 ;
        RECT 95.010 192.295 95.340 192.545 ;
        RECT 90.640 191.155 92.670 191.325 ;
        RECT 92.840 190.985 93.010 192.125 ;
        RECT 93.180 191.155 93.515 192.125 ;
        RECT 94.210 190.985 94.420 192.125 ;
        RECT 94.590 191.155 94.920 192.135 ;
        RECT 95.090 190.985 95.320 192.125 ;
        RECT 95.530 192.075 97.220 192.595 ;
        RECT 97.390 192.245 99.040 192.765 ;
        RECT 95.530 190.985 99.040 192.075 ;
        RECT 99.210 190.985 99.500 192.150 ;
        RECT 100.130 192.075 101.820 192.595 ;
        RECT 101.990 192.245 103.640 192.765 ;
        RECT 103.810 192.860 104.070 193.365 ;
        RECT 104.250 193.155 104.580 193.535 ;
        RECT 104.760 192.985 104.930 193.365 ;
        RECT 105.655 192.990 111.000 193.535 ;
        RECT 100.130 190.985 103.640 192.075 ;
        RECT 103.810 192.060 103.980 192.860 ;
        RECT 104.265 192.815 104.930 192.985 ;
        RECT 104.265 192.560 104.435 192.815 ;
        RECT 104.150 192.230 104.435 192.560 ;
        RECT 104.670 192.265 105.000 192.635 ;
        RECT 104.265 192.085 104.435 192.230 ;
        RECT 103.810 191.155 104.080 192.060 ;
        RECT 104.265 191.915 104.930 192.085 ;
        RECT 104.250 190.985 104.580 191.745 ;
        RECT 104.760 191.155 104.930 191.915 ;
        RECT 107.245 191.420 107.595 192.670 ;
        RECT 109.075 192.160 109.415 192.990 ;
        RECT 111.170 192.785 112.380 193.535 ;
        RECT 111.170 192.075 111.690 192.615 ;
        RECT 111.860 192.245 112.380 192.785 ;
        RECT 105.655 190.985 111.000 191.420 ;
        RECT 111.170 190.985 112.380 192.075 ;
        RECT 18.165 190.815 112.465 190.985 ;
        RECT 18.250 189.725 19.460 190.815 ;
        RECT 20.095 190.380 25.440 190.815 ;
        RECT 18.250 189.015 18.770 189.555 ;
        RECT 18.940 189.185 19.460 189.725 ;
        RECT 21.685 189.130 22.035 190.380 ;
        RECT 18.250 188.265 19.460 189.015 ;
        RECT 23.515 188.810 23.855 189.640 ;
        RECT 25.615 189.625 25.870 190.505 ;
        RECT 26.040 189.675 26.345 190.815 ;
        RECT 26.685 190.435 27.015 190.815 ;
        RECT 27.195 190.265 27.365 190.555 ;
        RECT 27.535 190.355 27.785 190.815 ;
        RECT 26.565 190.095 27.365 190.265 ;
        RECT 27.955 190.305 28.825 190.645 ;
        RECT 25.615 188.975 25.825 189.625 ;
        RECT 26.565 189.505 26.735 190.095 ;
        RECT 27.955 189.925 28.125 190.305 ;
        RECT 29.060 190.185 29.230 190.645 ;
        RECT 29.400 190.355 29.770 190.815 ;
        RECT 30.065 190.215 30.235 190.555 ;
        RECT 30.405 190.385 30.735 190.815 ;
        RECT 30.970 190.215 31.140 190.555 ;
        RECT 26.905 189.755 28.125 189.925 ;
        RECT 28.295 189.845 28.755 190.135 ;
        RECT 29.060 190.015 29.620 190.185 ;
        RECT 30.065 190.045 31.140 190.215 ;
        RECT 31.310 190.315 31.990 190.645 ;
        RECT 32.205 190.315 32.455 190.645 ;
        RECT 32.625 190.355 32.875 190.815 ;
        RECT 29.450 189.875 29.620 190.015 ;
        RECT 28.295 189.835 29.260 189.845 ;
        RECT 27.955 189.665 28.125 189.755 ;
        RECT 28.585 189.675 29.260 189.835 ;
        RECT 25.995 189.475 26.735 189.505 ;
        RECT 25.995 189.175 26.910 189.475 ;
        RECT 26.585 189.000 26.910 189.175 ;
        RECT 20.095 188.265 25.440 188.810 ;
        RECT 25.615 188.445 25.870 188.975 ;
        RECT 26.040 188.265 26.345 188.725 ;
        RECT 26.590 188.645 26.910 189.000 ;
        RECT 27.080 189.215 27.620 189.585 ;
        RECT 27.955 189.495 28.360 189.665 ;
        RECT 27.080 188.815 27.320 189.215 ;
        RECT 27.800 189.045 28.020 189.325 ;
        RECT 27.490 188.875 28.020 189.045 ;
        RECT 27.490 188.645 27.660 188.875 ;
        RECT 28.190 188.715 28.360 189.495 ;
        RECT 28.530 188.885 28.880 189.505 ;
        RECT 29.050 188.885 29.260 189.675 ;
        RECT 29.450 189.705 30.950 189.875 ;
        RECT 29.450 189.015 29.620 189.705 ;
        RECT 31.310 189.535 31.480 190.315 ;
        RECT 32.285 190.185 32.455 190.315 ;
        RECT 29.790 189.365 31.480 189.535 ;
        RECT 31.650 189.755 32.115 190.145 ;
        RECT 32.285 190.015 32.680 190.185 ;
        RECT 29.790 189.185 29.960 189.365 ;
        RECT 26.590 188.475 27.660 188.645 ;
        RECT 27.830 188.265 28.020 188.705 ;
        RECT 28.190 188.435 29.140 188.715 ;
        RECT 29.450 188.625 29.710 189.015 ;
        RECT 30.130 188.945 30.920 189.195 ;
        RECT 29.360 188.455 29.710 188.625 ;
        RECT 29.920 188.265 30.250 188.725 ;
        RECT 31.125 188.655 31.295 189.365 ;
        RECT 31.650 189.165 31.820 189.755 ;
        RECT 31.465 188.945 31.820 189.165 ;
        RECT 31.990 188.945 32.340 189.565 ;
        RECT 32.510 188.655 32.680 190.015 ;
        RECT 33.045 189.845 33.370 190.630 ;
        RECT 32.850 188.795 33.310 189.845 ;
        RECT 31.125 188.485 31.980 188.655 ;
        RECT 32.185 188.485 32.680 188.655 ;
        RECT 32.850 188.265 33.180 188.625 ;
        RECT 33.540 188.525 33.710 190.645 ;
        RECT 33.880 190.315 34.210 190.815 ;
        RECT 34.380 190.145 34.635 190.645 ;
        RECT 33.885 189.975 34.635 190.145 ;
        RECT 33.885 188.985 34.115 189.975 ;
        RECT 34.285 189.155 34.635 189.805 ;
        RECT 34.810 189.650 35.100 190.815 ;
        RECT 35.330 189.675 35.540 190.815 ;
        RECT 35.710 189.665 36.040 190.645 ;
        RECT 36.210 189.675 36.440 190.815 ;
        RECT 33.885 188.815 34.635 188.985 ;
        RECT 33.880 188.265 34.210 188.645 ;
        RECT 34.380 188.525 34.635 188.815 ;
        RECT 34.810 188.265 35.100 188.990 ;
        RECT 35.330 188.265 35.540 189.085 ;
        RECT 35.710 189.065 35.960 189.665 ;
        RECT 36.655 189.625 36.910 190.505 ;
        RECT 37.080 189.675 37.385 190.815 ;
        RECT 37.725 190.435 38.055 190.815 ;
        RECT 38.235 190.265 38.405 190.555 ;
        RECT 38.575 190.355 38.825 190.815 ;
        RECT 37.605 190.095 38.405 190.265 ;
        RECT 38.995 190.305 39.865 190.645 ;
        RECT 36.130 189.255 36.460 189.505 ;
        RECT 35.710 188.435 36.040 189.065 ;
        RECT 36.210 188.265 36.440 189.085 ;
        RECT 36.655 188.975 36.865 189.625 ;
        RECT 37.605 189.505 37.775 190.095 ;
        RECT 38.995 189.925 39.165 190.305 ;
        RECT 40.100 190.185 40.270 190.645 ;
        RECT 40.440 190.355 40.810 190.815 ;
        RECT 41.105 190.215 41.275 190.555 ;
        RECT 41.445 190.385 41.775 190.815 ;
        RECT 42.010 190.215 42.180 190.555 ;
        RECT 37.945 189.755 39.165 189.925 ;
        RECT 39.335 189.845 39.795 190.135 ;
        RECT 40.100 190.015 40.660 190.185 ;
        RECT 41.105 190.045 42.180 190.215 ;
        RECT 42.350 190.315 43.030 190.645 ;
        RECT 43.245 190.315 43.495 190.645 ;
        RECT 43.665 190.355 43.915 190.815 ;
        RECT 40.490 189.875 40.660 190.015 ;
        RECT 39.335 189.835 40.300 189.845 ;
        RECT 38.995 189.665 39.165 189.755 ;
        RECT 39.625 189.675 40.300 189.835 ;
        RECT 37.035 189.475 37.775 189.505 ;
        RECT 37.035 189.175 37.950 189.475 ;
        RECT 37.625 189.000 37.950 189.175 ;
        RECT 36.655 188.445 36.910 188.975 ;
        RECT 37.080 188.265 37.385 188.725 ;
        RECT 37.630 188.645 37.950 189.000 ;
        RECT 38.120 189.215 38.660 189.585 ;
        RECT 38.995 189.495 39.400 189.665 ;
        RECT 38.120 188.815 38.360 189.215 ;
        RECT 38.840 189.045 39.060 189.325 ;
        RECT 38.530 188.875 39.060 189.045 ;
        RECT 38.530 188.645 38.700 188.875 ;
        RECT 39.230 188.715 39.400 189.495 ;
        RECT 39.570 188.885 39.920 189.505 ;
        RECT 40.090 188.885 40.300 189.675 ;
        RECT 40.490 189.705 41.990 189.875 ;
        RECT 40.490 189.015 40.660 189.705 ;
        RECT 42.350 189.535 42.520 190.315 ;
        RECT 43.325 190.185 43.495 190.315 ;
        RECT 40.830 189.365 42.520 189.535 ;
        RECT 42.690 189.755 43.155 190.145 ;
        RECT 43.325 190.015 43.720 190.185 ;
        RECT 40.830 189.185 41.000 189.365 ;
        RECT 37.630 188.475 38.700 188.645 ;
        RECT 38.870 188.265 39.060 188.705 ;
        RECT 39.230 188.435 40.180 188.715 ;
        RECT 40.490 188.625 40.750 189.015 ;
        RECT 41.170 188.945 41.960 189.195 ;
        RECT 40.400 188.455 40.750 188.625 ;
        RECT 40.960 188.265 41.290 188.725 ;
        RECT 42.165 188.655 42.335 189.365 ;
        RECT 42.690 189.165 42.860 189.755 ;
        RECT 42.505 188.945 42.860 189.165 ;
        RECT 43.030 188.945 43.380 189.565 ;
        RECT 43.550 188.655 43.720 190.015 ;
        RECT 44.085 189.845 44.410 190.630 ;
        RECT 43.890 188.795 44.350 189.845 ;
        RECT 42.165 188.485 43.020 188.655 ;
        RECT 43.225 188.485 43.720 188.655 ;
        RECT 43.890 188.265 44.220 188.625 ;
        RECT 44.580 188.525 44.750 190.645 ;
        RECT 44.920 190.315 45.250 190.815 ;
        RECT 45.420 190.145 45.675 190.645 ;
        RECT 44.925 189.975 45.675 190.145 ;
        RECT 46.160 189.975 46.330 190.815 ;
        RECT 44.925 188.985 45.155 189.975 ;
        RECT 46.540 189.805 46.790 190.645 ;
        RECT 47.000 189.975 47.170 190.815 ;
        RECT 47.340 189.805 47.630 190.645 ;
        RECT 45.325 189.155 45.675 189.805 ;
        RECT 45.905 189.635 47.630 189.805 ;
        RECT 47.840 189.755 48.010 190.815 ;
        RECT 48.305 190.435 48.635 190.815 ;
        RECT 48.815 190.265 48.985 190.555 ;
        RECT 49.155 190.355 49.405 190.815 ;
        RECT 48.185 190.095 48.985 190.265 ;
        RECT 49.575 190.305 50.445 190.645 ;
        RECT 45.905 189.085 46.315 189.635 ;
        RECT 48.185 189.475 48.355 190.095 ;
        RECT 49.575 189.925 49.745 190.305 ;
        RECT 50.680 190.185 50.850 190.645 ;
        RECT 51.020 190.355 51.390 190.815 ;
        RECT 51.685 190.215 51.855 190.555 ;
        RECT 52.025 190.385 52.355 190.815 ;
        RECT 52.590 190.215 52.760 190.555 ;
        RECT 48.525 189.755 49.745 189.925 ;
        RECT 49.915 189.845 50.375 190.135 ;
        RECT 50.680 190.015 51.240 190.185 ;
        RECT 51.685 190.045 52.760 190.215 ;
        RECT 52.930 190.315 53.610 190.645 ;
        RECT 53.825 190.315 54.075 190.645 ;
        RECT 54.245 190.355 54.495 190.815 ;
        RECT 51.070 189.875 51.240 190.015 ;
        RECT 49.915 189.835 50.880 189.845 ;
        RECT 49.575 189.665 49.745 189.755 ;
        RECT 50.205 189.675 50.880 189.835 ;
        RECT 48.185 189.465 48.530 189.475 ;
        RECT 46.500 189.255 48.530 189.465 ;
        RECT 44.925 188.815 45.675 188.985 ;
        RECT 45.905 188.915 47.670 189.085 ;
        RECT 44.920 188.265 45.250 188.645 ;
        RECT 45.420 188.525 45.675 188.815 ;
        RECT 46.160 188.265 46.330 188.735 ;
        RECT 46.500 188.435 46.830 188.915 ;
        RECT 47.000 188.265 47.170 188.735 ;
        RECT 47.340 188.435 47.670 188.915 ;
        RECT 47.840 188.265 48.010 189.075 ;
        RECT 48.205 189.000 48.530 189.255 ;
        RECT 48.210 188.645 48.530 189.000 ;
        RECT 48.700 189.215 49.240 189.585 ;
        RECT 49.575 189.495 49.980 189.665 ;
        RECT 48.700 188.815 48.940 189.215 ;
        RECT 49.420 189.045 49.640 189.325 ;
        RECT 49.110 188.875 49.640 189.045 ;
        RECT 49.110 188.645 49.280 188.875 ;
        RECT 49.810 188.715 49.980 189.495 ;
        RECT 50.150 188.885 50.500 189.505 ;
        RECT 50.670 188.885 50.880 189.675 ;
        RECT 51.070 189.705 52.570 189.875 ;
        RECT 51.070 189.015 51.240 189.705 ;
        RECT 52.930 189.535 53.100 190.315 ;
        RECT 53.905 190.185 54.075 190.315 ;
        RECT 51.410 189.365 53.100 189.535 ;
        RECT 53.270 189.755 53.735 190.145 ;
        RECT 53.905 190.015 54.300 190.185 ;
        RECT 51.410 189.185 51.580 189.365 ;
        RECT 48.210 188.475 49.280 188.645 ;
        RECT 49.450 188.265 49.640 188.705 ;
        RECT 49.810 188.435 50.760 188.715 ;
        RECT 51.070 188.625 51.330 189.015 ;
        RECT 51.750 188.945 52.540 189.195 ;
        RECT 50.980 188.455 51.330 188.625 ;
        RECT 51.540 188.265 51.870 188.725 ;
        RECT 52.745 188.655 52.915 189.365 ;
        RECT 53.270 189.165 53.440 189.755 ;
        RECT 53.085 188.945 53.440 189.165 ;
        RECT 53.610 188.945 53.960 189.565 ;
        RECT 54.130 188.655 54.300 190.015 ;
        RECT 54.665 189.845 54.990 190.630 ;
        RECT 54.470 188.795 54.930 189.845 ;
        RECT 52.745 188.485 53.600 188.655 ;
        RECT 53.805 188.485 54.300 188.655 ;
        RECT 54.470 188.265 54.800 188.625 ;
        RECT 55.160 188.525 55.330 190.645 ;
        RECT 55.500 190.315 55.830 190.815 ;
        RECT 56.000 190.145 56.255 190.645 ;
        RECT 55.505 189.975 56.255 190.145 ;
        RECT 55.505 188.985 55.735 189.975 ;
        RECT 55.905 189.155 56.255 189.805 ;
        RECT 56.435 189.675 56.770 190.645 ;
        RECT 56.940 189.675 57.110 190.815 ;
        RECT 57.280 190.475 59.310 190.645 ;
        RECT 56.435 189.005 56.605 189.675 ;
        RECT 57.280 189.505 57.450 190.475 ;
        RECT 56.775 189.175 57.030 189.505 ;
        RECT 57.255 189.175 57.450 189.505 ;
        RECT 57.620 190.135 58.745 190.305 ;
        RECT 56.860 189.005 57.030 189.175 ;
        RECT 57.620 189.005 57.790 190.135 ;
        RECT 55.505 188.815 56.255 188.985 ;
        RECT 55.500 188.265 55.830 188.645 ;
        RECT 56.000 188.525 56.255 188.815 ;
        RECT 56.435 188.435 56.690 189.005 ;
        RECT 56.860 188.835 57.790 189.005 ;
        RECT 57.960 189.795 58.970 189.965 ;
        RECT 57.960 188.995 58.130 189.795 ;
        RECT 58.335 189.455 58.610 189.595 ;
        RECT 58.330 189.285 58.610 189.455 ;
        RECT 57.615 188.800 57.790 188.835 ;
        RECT 56.860 188.265 57.190 188.665 ;
        RECT 57.615 188.435 58.145 188.800 ;
        RECT 58.335 188.435 58.610 189.285 ;
        RECT 58.780 188.435 58.970 189.795 ;
        RECT 59.140 189.810 59.310 190.475 ;
        RECT 59.480 190.055 59.650 190.815 ;
        RECT 59.885 190.055 60.400 190.465 ;
        RECT 59.140 189.620 59.890 189.810 ;
        RECT 60.060 189.245 60.400 190.055 ;
        RECT 60.570 189.650 60.860 190.815 ;
        RECT 61.340 189.975 61.510 190.815 ;
        RECT 61.720 189.805 61.970 190.645 ;
        RECT 62.180 189.975 62.350 190.815 ;
        RECT 62.520 189.805 62.810 190.645 ;
        RECT 59.170 189.075 60.400 189.245 ;
        RECT 61.085 189.635 62.810 189.805 ;
        RECT 63.020 189.755 63.190 190.815 ;
        RECT 63.485 190.435 63.815 190.815 ;
        RECT 63.995 190.265 64.165 190.555 ;
        RECT 64.335 190.355 64.585 190.815 ;
        RECT 63.365 190.095 64.165 190.265 ;
        RECT 64.755 190.305 65.625 190.645 ;
        RECT 61.085 189.085 61.495 189.635 ;
        RECT 63.365 189.475 63.535 190.095 ;
        RECT 64.755 189.925 64.925 190.305 ;
        RECT 65.860 190.185 66.030 190.645 ;
        RECT 66.200 190.355 66.570 190.815 ;
        RECT 66.865 190.215 67.035 190.555 ;
        RECT 67.205 190.385 67.535 190.815 ;
        RECT 67.770 190.215 67.940 190.555 ;
        RECT 63.705 189.755 64.925 189.925 ;
        RECT 65.095 189.845 65.555 190.135 ;
        RECT 65.860 190.015 66.420 190.185 ;
        RECT 66.865 190.045 67.940 190.215 ;
        RECT 68.110 190.315 68.790 190.645 ;
        RECT 69.005 190.315 69.255 190.645 ;
        RECT 69.425 190.355 69.675 190.815 ;
        RECT 66.250 189.875 66.420 190.015 ;
        RECT 65.095 189.835 66.060 189.845 ;
        RECT 64.755 189.665 64.925 189.755 ;
        RECT 65.385 189.675 66.060 189.835 ;
        RECT 63.365 189.465 63.710 189.475 ;
        RECT 61.680 189.255 63.710 189.465 ;
        RECT 59.150 188.265 59.660 188.800 ;
        RECT 59.880 188.470 60.125 189.075 ;
        RECT 60.570 188.265 60.860 188.990 ;
        RECT 61.085 188.915 62.850 189.085 ;
        RECT 61.340 188.265 61.510 188.735 ;
        RECT 61.680 188.435 62.010 188.915 ;
        RECT 62.180 188.265 62.350 188.735 ;
        RECT 62.520 188.435 62.850 188.915 ;
        RECT 63.020 188.265 63.190 189.075 ;
        RECT 63.385 189.000 63.710 189.255 ;
        RECT 63.390 188.645 63.710 189.000 ;
        RECT 63.880 189.215 64.420 189.585 ;
        RECT 64.755 189.495 65.160 189.665 ;
        RECT 63.880 188.815 64.120 189.215 ;
        RECT 64.600 189.045 64.820 189.325 ;
        RECT 64.290 188.875 64.820 189.045 ;
        RECT 64.290 188.645 64.460 188.875 ;
        RECT 64.990 188.715 65.160 189.495 ;
        RECT 65.330 188.885 65.680 189.505 ;
        RECT 65.850 188.885 66.060 189.675 ;
        RECT 66.250 189.705 67.750 189.875 ;
        RECT 66.250 189.015 66.420 189.705 ;
        RECT 68.110 189.535 68.280 190.315 ;
        RECT 69.085 190.185 69.255 190.315 ;
        RECT 66.590 189.365 68.280 189.535 ;
        RECT 68.450 189.755 68.915 190.145 ;
        RECT 69.085 190.015 69.480 190.185 ;
        RECT 66.590 189.185 66.760 189.365 ;
        RECT 63.390 188.475 64.460 188.645 ;
        RECT 64.630 188.265 64.820 188.705 ;
        RECT 64.990 188.435 65.940 188.715 ;
        RECT 66.250 188.625 66.510 189.015 ;
        RECT 66.930 188.945 67.720 189.195 ;
        RECT 66.160 188.455 66.510 188.625 ;
        RECT 66.720 188.265 67.050 188.725 ;
        RECT 67.925 188.655 68.095 189.365 ;
        RECT 68.450 189.165 68.620 189.755 ;
        RECT 68.265 188.945 68.620 189.165 ;
        RECT 68.790 188.945 69.140 189.565 ;
        RECT 69.310 188.655 69.480 190.015 ;
        RECT 69.845 189.845 70.170 190.630 ;
        RECT 69.650 188.795 70.110 189.845 ;
        RECT 67.925 188.485 68.780 188.655 ;
        RECT 68.985 188.485 69.480 188.655 ;
        RECT 69.650 188.265 69.980 188.625 ;
        RECT 70.340 188.525 70.510 190.645 ;
        RECT 70.680 190.315 71.010 190.815 ;
        RECT 71.180 190.145 71.435 190.645 ;
        RECT 70.685 189.975 71.435 190.145 ;
        RECT 70.685 188.985 70.915 189.975 ;
        RECT 71.085 189.155 71.435 189.805 ;
        RECT 71.650 189.675 71.880 190.815 ;
        RECT 72.050 189.665 72.380 190.645 ;
        RECT 72.550 189.675 72.760 190.815 ;
        RECT 73.760 189.975 73.930 190.815 ;
        RECT 74.140 189.805 74.390 190.645 ;
        RECT 74.600 189.975 74.770 190.815 ;
        RECT 74.940 189.805 75.230 190.645 ;
        RECT 71.630 189.255 71.960 189.505 ;
        RECT 70.685 188.815 71.435 188.985 ;
        RECT 70.680 188.265 71.010 188.645 ;
        RECT 71.180 188.525 71.435 188.815 ;
        RECT 71.650 188.265 71.880 189.085 ;
        RECT 72.130 189.065 72.380 189.665 ;
        RECT 73.505 189.635 75.230 189.805 ;
        RECT 75.440 189.755 75.610 190.815 ;
        RECT 75.905 190.435 76.235 190.815 ;
        RECT 76.415 190.265 76.585 190.555 ;
        RECT 76.755 190.355 77.005 190.815 ;
        RECT 75.785 190.095 76.585 190.265 ;
        RECT 77.175 190.305 78.045 190.645 ;
        RECT 73.505 189.085 73.915 189.635 ;
        RECT 75.785 189.475 75.955 190.095 ;
        RECT 77.175 189.925 77.345 190.305 ;
        RECT 78.280 190.185 78.450 190.645 ;
        RECT 78.620 190.355 78.990 190.815 ;
        RECT 79.285 190.215 79.455 190.555 ;
        RECT 79.625 190.385 79.955 190.815 ;
        RECT 80.190 190.215 80.360 190.555 ;
        RECT 76.125 189.755 77.345 189.925 ;
        RECT 77.515 189.845 77.975 190.135 ;
        RECT 78.280 190.015 78.840 190.185 ;
        RECT 79.285 190.045 80.360 190.215 ;
        RECT 80.530 190.315 81.210 190.645 ;
        RECT 81.425 190.315 81.675 190.645 ;
        RECT 81.845 190.355 82.095 190.815 ;
        RECT 78.670 189.875 78.840 190.015 ;
        RECT 77.515 189.835 78.480 189.845 ;
        RECT 77.175 189.665 77.345 189.755 ;
        RECT 77.805 189.675 78.480 189.835 ;
        RECT 75.785 189.465 76.130 189.475 ;
        RECT 74.100 189.255 76.130 189.465 ;
        RECT 72.050 188.435 72.380 189.065 ;
        RECT 72.550 188.265 72.760 189.085 ;
        RECT 73.505 188.915 75.270 189.085 ;
        RECT 73.760 188.265 73.930 188.735 ;
        RECT 74.100 188.435 74.430 188.915 ;
        RECT 74.600 188.265 74.770 188.735 ;
        RECT 74.940 188.435 75.270 188.915 ;
        RECT 75.440 188.265 75.610 189.075 ;
        RECT 75.805 189.000 76.130 189.255 ;
        RECT 75.810 188.645 76.130 189.000 ;
        RECT 76.300 189.215 76.840 189.585 ;
        RECT 77.175 189.495 77.580 189.665 ;
        RECT 76.300 188.815 76.540 189.215 ;
        RECT 77.020 189.045 77.240 189.325 ;
        RECT 76.710 188.875 77.240 189.045 ;
        RECT 76.710 188.645 76.880 188.875 ;
        RECT 77.410 188.715 77.580 189.495 ;
        RECT 77.750 188.885 78.100 189.505 ;
        RECT 78.270 188.885 78.480 189.675 ;
        RECT 78.670 189.705 80.170 189.875 ;
        RECT 78.670 189.015 78.840 189.705 ;
        RECT 80.530 189.535 80.700 190.315 ;
        RECT 81.505 190.185 81.675 190.315 ;
        RECT 79.010 189.365 80.700 189.535 ;
        RECT 80.870 189.755 81.335 190.145 ;
        RECT 81.505 190.015 81.900 190.185 ;
        RECT 79.010 189.185 79.180 189.365 ;
        RECT 75.810 188.475 76.880 188.645 ;
        RECT 77.050 188.265 77.240 188.705 ;
        RECT 77.410 188.435 78.360 188.715 ;
        RECT 78.670 188.625 78.930 189.015 ;
        RECT 79.350 188.945 80.140 189.195 ;
        RECT 78.580 188.455 78.930 188.625 ;
        RECT 79.140 188.265 79.470 188.725 ;
        RECT 80.345 188.655 80.515 189.365 ;
        RECT 80.870 189.165 81.040 189.755 ;
        RECT 80.685 188.945 81.040 189.165 ;
        RECT 81.210 188.945 81.560 189.565 ;
        RECT 81.730 188.655 81.900 190.015 ;
        RECT 82.265 189.845 82.590 190.630 ;
        RECT 82.070 188.795 82.530 189.845 ;
        RECT 80.345 188.485 81.200 188.655 ;
        RECT 81.405 188.485 81.900 188.655 ;
        RECT 82.070 188.265 82.400 188.625 ;
        RECT 82.760 188.525 82.930 190.645 ;
        RECT 83.100 190.315 83.430 190.815 ;
        RECT 83.600 190.145 83.855 190.645 ;
        RECT 83.105 189.975 83.855 190.145 ;
        RECT 83.105 188.985 83.335 189.975 ;
        RECT 83.505 189.155 83.855 189.805 ;
        RECT 84.090 189.675 84.300 190.815 ;
        RECT 84.470 189.665 84.800 190.645 ;
        RECT 84.970 189.675 85.200 190.815 ;
        RECT 83.105 188.815 83.855 188.985 ;
        RECT 83.100 188.265 83.430 188.645 ;
        RECT 83.600 188.525 83.855 188.815 ;
        RECT 84.090 188.265 84.300 189.085 ;
        RECT 84.470 189.065 84.720 189.665 ;
        RECT 86.330 189.650 86.620 190.815 ;
        RECT 86.940 189.665 87.270 190.815 ;
        RECT 87.440 189.795 87.610 190.645 ;
        RECT 87.780 190.015 88.110 190.815 ;
        RECT 88.280 189.795 88.450 190.645 ;
        RECT 88.630 190.015 88.870 190.815 ;
        RECT 89.040 189.835 89.370 190.645 ;
        RECT 87.440 189.625 88.450 189.795 ;
        RECT 88.655 189.665 89.370 189.835 ;
        RECT 90.845 189.835 91.100 190.505 ;
        RECT 91.280 190.015 91.565 190.815 ;
        RECT 91.745 190.095 92.075 190.605 ;
        RECT 84.890 189.255 85.220 189.505 ;
        RECT 87.440 189.455 87.935 189.625 ;
        RECT 87.440 189.285 87.940 189.455 ;
        RECT 88.655 189.425 88.825 189.665 ;
        RECT 87.440 189.085 87.935 189.285 ;
        RECT 88.325 189.255 88.825 189.425 ;
        RECT 88.995 189.255 89.375 189.495 ;
        RECT 88.655 189.085 88.825 189.255 ;
        RECT 84.470 188.435 84.800 189.065 ;
        RECT 84.970 188.265 85.200 189.085 ;
        RECT 86.330 188.265 86.620 188.990 ;
        RECT 86.940 188.265 87.270 189.065 ;
        RECT 87.440 188.915 88.450 189.085 ;
        RECT 88.655 188.915 89.290 189.085 ;
        RECT 87.440 188.435 87.610 188.915 ;
        RECT 87.780 188.265 88.110 188.745 ;
        RECT 88.280 188.435 88.450 188.915 ;
        RECT 88.700 188.265 88.940 188.745 ;
        RECT 89.120 188.435 89.290 188.915 ;
        RECT 90.845 188.975 91.025 189.835 ;
        RECT 91.745 189.505 91.995 190.095 ;
        RECT 92.345 189.945 92.515 190.555 ;
        RECT 92.685 190.125 93.015 190.815 ;
        RECT 93.245 190.265 93.485 190.555 ;
        RECT 93.685 190.435 94.105 190.815 ;
        RECT 94.285 190.345 94.915 190.595 ;
        RECT 95.385 190.435 95.715 190.815 ;
        RECT 94.285 190.265 94.455 190.345 ;
        RECT 95.885 190.265 96.055 190.555 ;
        RECT 96.235 190.435 96.615 190.815 ;
        RECT 96.855 190.430 97.685 190.600 ;
        RECT 93.245 190.095 94.455 190.265 ;
        RECT 91.195 189.175 91.995 189.505 ;
        RECT 90.845 188.775 91.100 188.975 ;
        RECT 90.760 188.605 91.100 188.775 ;
        RECT 90.845 188.445 91.100 188.605 ;
        RECT 91.280 188.265 91.565 188.725 ;
        RECT 91.745 188.525 91.995 189.175 ;
        RECT 92.195 189.925 92.515 189.945 ;
        RECT 92.195 189.755 94.115 189.925 ;
        RECT 92.195 188.860 92.385 189.755 ;
        RECT 94.285 189.585 94.455 190.095 ;
        RECT 94.625 189.835 95.145 190.145 ;
        RECT 92.555 189.415 94.455 189.585 ;
        RECT 92.555 189.355 92.885 189.415 ;
        RECT 93.035 189.185 93.365 189.245 ;
        RECT 92.705 188.915 93.365 189.185 ;
        RECT 92.195 188.530 92.515 188.860 ;
        RECT 92.695 188.265 93.355 188.745 ;
        RECT 93.555 188.655 93.725 189.415 ;
        RECT 94.625 189.245 94.805 189.655 ;
        RECT 93.895 189.075 94.225 189.195 ;
        RECT 94.975 189.075 95.145 189.835 ;
        RECT 93.895 188.905 95.145 189.075 ;
        RECT 95.315 190.015 96.685 190.265 ;
        RECT 95.315 189.245 95.505 190.015 ;
        RECT 96.435 189.755 96.685 190.015 ;
        RECT 95.675 189.585 95.925 189.745 ;
        RECT 96.855 189.585 97.025 190.430 ;
        RECT 97.920 190.145 98.090 190.645 ;
        RECT 98.260 190.315 98.590 190.815 ;
        RECT 97.195 189.755 97.695 190.135 ;
        RECT 97.920 189.975 98.615 190.145 ;
        RECT 95.675 189.415 97.025 189.585 ;
        RECT 96.605 189.375 97.025 189.415 ;
        RECT 95.315 188.905 95.735 189.245 ;
        RECT 96.025 188.915 96.435 189.245 ;
        RECT 93.555 188.485 94.405 188.655 ;
        RECT 94.965 188.265 95.285 188.725 ;
        RECT 95.485 188.475 95.735 188.905 ;
        RECT 96.025 188.265 96.435 188.705 ;
        RECT 96.605 188.645 96.775 189.375 ;
        RECT 96.945 188.825 97.295 189.195 ;
        RECT 97.475 188.885 97.695 189.755 ;
        RECT 97.865 189.185 98.275 189.805 ;
        RECT 98.445 189.005 98.615 189.975 ;
        RECT 97.920 188.815 98.615 189.005 ;
        RECT 96.605 188.445 97.620 188.645 ;
        RECT 97.920 188.485 98.090 188.815 ;
        RECT 98.260 188.265 98.590 188.645 ;
        RECT 98.805 188.525 99.030 190.645 ;
        RECT 99.200 190.315 99.530 190.815 ;
        RECT 99.700 190.145 99.870 190.645 ;
        RECT 100.135 190.380 105.480 190.815 ;
        RECT 105.655 190.380 111.000 190.815 ;
        RECT 99.205 189.975 99.870 190.145 ;
        RECT 99.205 188.985 99.435 189.975 ;
        RECT 99.605 189.155 99.955 189.805 ;
        RECT 101.725 189.130 102.075 190.380 ;
        RECT 99.205 188.815 99.870 188.985 ;
        RECT 99.200 188.265 99.530 188.645 ;
        RECT 99.700 188.525 99.870 188.815 ;
        RECT 103.555 188.810 103.895 189.640 ;
        RECT 107.245 189.130 107.595 190.380 ;
        RECT 111.170 189.725 112.380 190.815 ;
        RECT 109.075 188.810 109.415 189.640 ;
        RECT 111.170 189.185 111.690 189.725 ;
        RECT 111.860 189.015 112.380 189.555 ;
        RECT 100.135 188.265 105.480 188.810 ;
        RECT 105.655 188.265 111.000 188.810 ;
        RECT 111.170 188.265 112.380 189.015 ;
        RECT 18.165 188.095 112.465 188.265 ;
        RECT 18.250 187.345 19.460 188.095 ;
        RECT 18.250 186.805 18.770 187.345 ;
        RECT 20.090 187.325 21.760 188.095 ;
        RECT 21.930 187.370 22.220 188.095 ;
        RECT 23.310 187.325 26.820 188.095 ;
        RECT 26.990 187.715 27.880 187.885 ;
        RECT 18.940 186.635 19.460 187.175 ;
        RECT 18.250 185.545 19.460 186.635 ;
        RECT 20.090 186.635 20.840 187.155 ;
        RECT 21.010 186.805 21.760 187.325 ;
        RECT 20.090 185.545 21.760 186.635 ;
        RECT 21.930 185.545 22.220 186.710 ;
        RECT 23.310 186.635 25.000 187.155 ;
        RECT 25.170 186.805 26.820 187.325 ;
        RECT 26.990 187.160 27.540 187.545 ;
        RECT 27.710 186.990 27.880 187.715 ;
        RECT 26.990 186.920 27.880 186.990 ;
        RECT 28.050 187.415 28.270 187.875 ;
        RECT 28.440 187.555 28.690 188.095 ;
        RECT 28.860 187.445 29.120 187.925 ;
        RECT 28.050 187.390 28.300 187.415 ;
        RECT 28.050 186.965 28.380 187.390 ;
        RECT 26.990 186.895 27.885 186.920 ;
        RECT 26.990 186.880 27.895 186.895 ;
        RECT 26.990 186.865 27.900 186.880 ;
        RECT 26.990 186.860 27.910 186.865 ;
        RECT 26.990 186.850 27.915 186.860 ;
        RECT 26.990 186.840 27.920 186.850 ;
        RECT 26.990 186.835 27.930 186.840 ;
        RECT 26.990 186.825 27.940 186.835 ;
        RECT 26.990 186.820 27.950 186.825 ;
        RECT 23.310 185.545 26.820 186.635 ;
        RECT 26.990 186.370 27.250 186.820 ;
        RECT 27.615 186.815 27.950 186.820 ;
        RECT 27.615 186.810 27.965 186.815 ;
        RECT 27.615 186.800 27.980 186.810 ;
        RECT 27.615 186.795 28.005 186.800 ;
        RECT 28.550 186.795 28.780 187.190 ;
        RECT 27.615 186.790 28.780 186.795 ;
        RECT 27.645 186.755 28.780 186.790 ;
        RECT 27.680 186.730 28.780 186.755 ;
        RECT 27.710 186.700 28.780 186.730 ;
        RECT 27.730 186.670 28.780 186.700 ;
        RECT 27.750 186.640 28.780 186.670 ;
        RECT 27.820 186.630 28.780 186.640 ;
        RECT 27.845 186.620 28.780 186.630 ;
        RECT 27.865 186.605 28.780 186.620 ;
        RECT 27.885 186.590 28.780 186.605 ;
        RECT 27.890 186.580 28.675 186.590 ;
        RECT 27.905 186.545 28.675 186.580 ;
        RECT 27.420 186.225 27.750 186.470 ;
        RECT 27.920 186.295 28.675 186.545 ;
        RECT 28.950 186.415 29.120 187.445 ;
        RECT 29.290 187.325 30.960 188.095 ;
        RECT 27.420 186.200 27.605 186.225 ;
        RECT 26.990 186.100 27.605 186.200 ;
        RECT 26.990 185.545 27.595 186.100 ;
        RECT 27.770 185.715 28.250 186.055 ;
        RECT 28.420 185.545 28.675 186.090 ;
        RECT 28.845 185.715 29.120 186.415 ;
        RECT 29.290 186.635 30.040 187.155 ;
        RECT 30.210 186.805 30.960 187.325 ;
        RECT 31.135 187.385 31.390 187.915 ;
        RECT 31.560 187.635 31.865 188.095 ;
        RECT 32.110 187.715 33.180 187.885 ;
        RECT 31.135 186.735 31.345 187.385 ;
        RECT 32.110 187.360 32.430 187.715 ;
        RECT 32.105 187.185 32.430 187.360 ;
        RECT 31.515 186.885 32.430 187.185 ;
        RECT 32.600 187.145 32.840 187.545 ;
        RECT 33.010 187.485 33.180 187.715 ;
        RECT 33.350 187.655 33.540 188.095 ;
        RECT 33.710 187.645 34.660 187.925 ;
        RECT 34.880 187.735 35.230 187.905 ;
        RECT 33.010 187.315 33.540 187.485 ;
        RECT 31.515 186.855 32.255 186.885 ;
        RECT 29.290 185.545 30.960 186.635 ;
        RECT 31.135 185.855 31.390 186.735 ;
        RECT 31.560 185.545 31.865 186.685 ;
        RECT 32.085 186.265 32.255 186.855 ;
        RECT 32.600 186.775 33.140 187.145 ;
        RECT 33.320 187.035 33.540 187.315 ;
        RECT 33.710 186.865 33.880 187.645 ;
        RECT 33.475 186.695 33.880 186.865 ;
        RECT 34.050 186.855 34.400 187.475 ;
        RECT 33.475 186.605 33.645 186.695 ;
        RECT 34.570 186.685 34.780 187.475 ;
        RECT 32.425 186.435 33.645 186.605 ;
        RECT 34.105 186.525 34.780 186.685 ;
        RECT 32.085 186.095 32.885 186.265 ;
        RECT 32.205 185.545 32.535 185.925 ;
        RECT 32.715 185.805 32.885 186.095 ;
        RECT 33.475 186.055 33.645 186.435 ;
        RECT 33.815 186.515 34.780 186.525 ;
        RECT 34.970 187.345 35.230 187.735 ;
        RECT 35.440 187.635 35.770 188.095 ;
        RECT 36.645 187.705 37.500 187.875 ;
        RECT 37.705 187.705 38.200 187.875 ;
        RECT 38.370 187.735 38.700 188.095 ;
        RECT 34.970 186.655 35.140 187.345 ;
        RECT 35.310 186.995 35.480 187.175 ;
        RECT 35.650 187.165 36.440 187.415 ;
        RECT 36.645 186.995 36.815 187.705 ;
        RECT 36.985 187.195 37.340 187.415 ;
        RECT 35.310 186.825 37.000 186.995 ;
        RECT 33.815 186.225 34.275 186.515 ;
        RECT 34.970 186.485 36.470 186.655 ;
        RECT 34.970 186.345 35.140 186.485 ;
        RECT 34.580 186.175 35.140 186.345 ;
        RECT 33.055 185.545 33.305 186.005 ;
        RECT 33.475 185.715 34.345 186.055 ;
        RECT 34.580 185.715 34.750 186.175 ;
        RECT 35.585 186.145 36.660 186.315 ;
        RECT 34.920 185.545 35.290 186.005 ;
        RECT 35.585 185.805 35.755 186.145 ;
        RECT 35.925 185.545 36.255 185.975 ;
        RECT 36.490 185.805 36.660 186.145 ;
        RECT 36.830 186.045 37.000 186.825 ;
        RECT 37.170 186.605 37.340 187.195 ;
        RECT 37.510 186.795 37.860 187.415 ;
        RECT 37.170 186.215 37.635 186.605 ;
        RECT 38.030 186.345 38.200 187.705 ;
        RECT 38.370 186.515 38.830 187.565 ;
        RECT 37.805 186.175 38.200 186.345 ;
        RECT 37.805 186.045 37.975 186.175 ;
        RECT 36.830 185.715 37.510 186.045 ;
        RECT 37.725 185.715 37.975 186.045 ;
        RECT 38.145 185.545 38.395 186.005 ;
        RECT 38.565 185.730 38.890 186.515 ;
        RECT 39.060 185.715 39.230 187.835 ;
        RECT 39.400 187.715 39.730 188.095 ;
        RECT 39.900 187.545 40.155 187.835 ;
        RECT 39.405 187.375 40.155 187.545 ;
        RECT 39.405 186.385 39.635 187.375 ;
        RECT 40.330 187.355 40.650 187.835 ;
        RECT 40.820 187.525 41.050 187.925 ;
        RECT 41.220 187.705 41.570 188.095 ;
        RECT 40.820 187.445 41.330 187.525 ;
        RECT 41.740 187.445 42.070 187.925 ;
        RECT 40.820 187.355 42.070 187.445 ;
        RECT 39.805 186.555 40.155 187.205 ;
        RECT 40.330 186.425 40.500 187.355 ;
        RECT 41.160 187.275 42.070 187.355 ;
        RECT 42.240 187.275 42.410 188.095 ;
        RECT 42.915 187.355 43.380 187.900 ;
        RECT 40.670 186.765 40.840 187.185 ;
        RECT 41.070 186.935 41.670 187.105 ;
        RECT 40.670 186.595 41.330 186.765 ;
        RECT 39.405 186.215 40.155 186.385 ;
        RECT 40.330 186.225 40.990 186.425 ;
        RECT 41.160 186.395 41.330 186.595 ;
        RECT 41.500 186.735 41.670 186.935 ;
        RECT 41.840 186.905 42.535 187.105 ;
        RECT 42.795 186.735 43.040 187.185 ;
        RECT 41.500 186.565 43.040 186.735 ;
        RECT 43.210 186.395 43.380 187.355 ;
        RECT 44.050 187.275 44.280 188.095 ;
        RECT 44.450 187.295 44.780 187.925 ;
        RECT 44.030 186.855 44.360 187.105 ;
        RECT 44.530 186.695 44.780 187.295 ;
        RECT 44.950 187.275 45.160 188.095 ;
        RECT 45.850 187.325 47.520 188.095 ;
        RECT 47.690 187.370 47.980 188.095 ;
        RECT 41.160 186.225 43.380 186.395 ;
        RECT 39.400 185.545 39.730 186.045 ;
        RECT 39.900 185.715 40.155 186.215 ;
        RECT 40.820 186.055 40.990 186.225 ;
        RECT 40.350 185.545 40.650 186.055 ;
        RECT 40.820 185.885 41.200 186.055 ;
        RECT 41.780 185.545 42.410 186.055 ;
        RECT 42.580 185.715 42.910 186.225 ;
        RECT 43.080 185.545 43.380 186.055 ;
        RECT 44.050 185.545 44.280 186.685 ;
        RECT 44.450 185.715 44.780 186.695 ;
        RECT 44.950 185.545 45.160 186.685 ;
        RECT 45.850 186.635 46.600 187.155 ;
        RECT 46.770 186.805 47.520 187.325 ;
        RECT 48.155 187.355 48.410 187.925 ;
        RECT 48.580 187.695 48.910 188.095 ;
        RECT 49.335 187.560 49.865 187.925 ;
        RECT 49.335 187.525 49.510 187.560 ;
        RECT 48.580 187.355 49.510 187.525 ;
        RECT 50.055 187.415 50.330 187.925 ;
        RECT 45.850 185.545 47.520 186.635 ;
        RECT 47.690 185.545 47.980 186.710 ;
        RECT 48.155 186.685 48.325 187.355 ;
        RECT 48.580 187.185 48.750 187.355 ;
        RECT 48.495 186.855 48.750 187.185 ;
        RECT 48.975 186.855 49.170 187.185 ;
        RECT 48.155 185.715 48.490 186.685 ;
        RECT 48.660 185.545 48.830 186.685 ;
        RECT 49.000 185.885 49.170 186.855 ;
        RECT 49.340 186.225 49.510 187.355 ;
        RECT 49.680 186.565 49.850 187.365 ;
        RECT 50.050 187.245 50.330 187.415 ;
        RECT 50.055 186.765 50.330 187.245 ;
        RECT 50.500 186.565 50.690 187.925 ;
        RECT 50.870 187.560 51.380 188.095 ;
        RECT 51.600 187.285 51.845 187.890 ;
        RECT 50.890 187.115 52.120 187.285 ;
        RECT 52.330 187.275 52.560 188.095 ;
        RECT 52.730 187.295 53.060 187.925 ;
        RECT 49.680 186.395 50.690 186.565 ;
        RECT 50.860 186.550 51.610 186.740 ;
        RECT 49.340 186.055 50.465 186.225 ;
        RECT 50.860 185.885 51.030 186.550 ;
        RECT 51.780 186.305 52.120 187.115 ;
        RECT 52.310 186.855 52.640 187.105 ;
        RECT 52.810 186.695 53.060 187.295 ;
        RECT 53.230 187.275 53.440 188.095 ;
        RECT 54.680 187.545 54.850 187.925 ;
        RECT 55.065 187.715 55.395 188.095 ;
        RECT 54.680 187.375 55.395 187.545 ;
        RECT 54.590 186.825 54.945 187.195 ;
        RECT 55.225 187.185 55.395 187.375 ;
        RECT 55.565 187.350 55.820 187.925 ;
        RECT 55.225 186.855 55.480 187.185 ;
        RECT 49.000 185.715 51.030 185.885 ;
        RECT 51.200 185.545 51.370 186.305 ;
        RECT 51.605 185.895 52.120 186.305 ;
        RECT 52.330 185.545 52.560 186.685 ;
        RECT 52.730 185.715 53.060 186.695 ;
        RECT 53.230 185.545 53.440 186.685 ;
        RECT 55.225 186.645 55.395 186.855 ;
        RECT 54.680 186.475 55.395 186.645 ;
        RECT 55.650 186.620 55.820 187.350 ;
        RECT 55.995 187.255 56.255 188.095 ;
        RECT 56.520 187.545 56.690 187.835 ;
        RECT 56.860 187.715 57.190 188.095 ;
        RECT 56.520 187.375 57.185 187.545 ;
        RECT 54.680 185.715 54.850 186.475 ;
        RECT 55.065 185.545 55.395 186.305 ;
        RECT 55.565 185.715 55.820 186.620 ;
        RECT 55.995 185.545 56.255 186.695 ;
        RECT 56.435 186.555 56.785 187.205 ;
        RECT 56.955 186.385 57.185 187.375 ;
        RECT 56.520 186.215 57.185 186.385 ;
        RECT 56.520 185.715 56.690 186.215 ;
        RECT 56.860 185.545 57.190 186.045 ;
        RECT 57.360 185.715 57.585 187.835 ;
        RECT 57.800 187.715 58.130 188.095 ;
        RECT 58.300 187.545 58.470 187.875 ;
        RECT 58.770 187.715 59.785 187.915 ;
        RECT 57.775 187.355 58.470 187.545 ;
        RECT 57.775 186.385 57.945 187.355 ;
        RECT 58.115 186.555 58.525 187.175 ;
        RECT 58.695 186.605 58.915 187.475 ;
        RECT 59.095 187.165 59.445 187.535 ;
        RECT 59.615 186.985 59.785 187.715 ;
        RECT 59.955 187.655 60.365 188.095 ;
        RECT 60.655 187.455 60.905 187.885 ;
        RECT 61.105 187.635 61.425 188.095 ;
        RECT 61.985 187.705 62.835 187.875 ;
        RECT 59.955 187.115 60.365 187.445 ;
        RECT 60.655 187.115 61.075 187.455 ;
        RECT 59.365 186.945 59.785 186.985 ;
        RECT 59.365 186.775 60.715 186.945 ;
        RECT 57.775 186.215 58.470 186.385 ;
        RECT 58.695 186.225 59.195 186.605 ;
        RECT 57.800 185.545 58.130 186.045 ;
        RECT 58.300 185.715 58.470 186.215 ;
        RECT 59.365 185.930 59.535 186.775 ;
        RECT 60.465 186.615 60.715 186.775 ;
        RECT 59.705 186.345 59.955 186.605 ;
        RECT 60.885 186.345 61.075 187.115 ;
        RECT 59.705 186.095 61.075 186.345 ;
        RECT 61.245 187.285 62.495 187.455 ;
        RECT 61.245 186.525 61.415 187.285 ;
        RECT 62.165 187.165 62.495 187.285 ;
        RECT 61.585 186.705 61.765 187.115 ;
        RECT 62.665 186.945 62.835 187.705 ;
        RECT 63.035 187.615 63.695 188.095 ;
        RECT 63.875 187.500 64.195 187.830 ;
        RECT 63.025 187.175 63.685 187.445 ;
        RECT 63.025 187.115 63.355 187.175 ;
        RECT 63.505 186.945 63.835 187.005 ;
        RECT 61.935 186.775 63.835 186.945 ;
        RECT 61.245 186.215 61.765 186.525 ;
        RECT 61.935 186.265 62.105 186.775 ;
        RECT 64.005 186.605 64.195 187.500 ;
        RECT 62.275 186.435 64.195 186.605 ;
        RECT 63.875 186.415 64.195 186.435 ;
        RECT 64.395 187.185 64.645 187.835 ;
        RECT 64.825 187.635 65.110 188.095 ;
        RECT 65.290 187.755 65.545 187.915 ;
        RECT 65.290 187.585 65.630 187.755 ;
        RECT 65.290 187.385 65.545 187.585 ;
        RECT 64.395 186.855 65.195 187.185 ;
        RECT 61.935 186.095 63.145 186.265 ;
        RECT 58.705 185.760 59.535 185.930 ;
        RECT 59.775 185.545 60.155 185.925 ;
        RECT 60.335 185.805 60.505 186.095 ;
        RECT 61.935 186.015 62.105 186.095 ;
        RECT 60.675 185.545 61.005 185.925 ;
        RECT 61.475 185.765 62.105 186.015 ;
        RECT 62.285 185.545 62.705 185.925 ;
        RECT 62.905 185.805 63.145 186.095 ;
        RECT 63.375 185.545 63.705 186.235 ;
        RECT 63.875 185.805 64.045 186.415 ;
        RECT 64.395 186.265 64.645 186.855 ;
        RECT 65.365 186.525 65.545 187.385 ;
        RECT 66.550 187.325 69.140 188.095 ;
        RECT 64.315 185.755 64.645 186.265 ;
        RECT 64.825 185.545 65.110 186.345 ;
        RECT 65.290 185.855 65.545 186.525 ;
        RECT 66.550 186.635 67.760 187.155 ;
        RECT 67.930 186.805 69.140 187.325 ;
        RECT 69.585 187.285 69.830 187.890 ;
        RECT 70.050 187.560 70.560 188.095 ;
        RECT 69.310 187.115 70.540 187.285 ;
        RECT 66.550 185.545 69.140 186.635 ;
        RECT 69.310 186.305 69.650 187.115 ;
        RECT 69.820 186.550 70.570 186.740 ;
        RECT 69.310 185.895 69.825 186.305 ;
        RECT 70.060 185.545 70.230 186.305 ;
        RECT 70.400 185.885 70.570 186.550 ;
        RECT 70.740 186.565 70.930 187.925 ;
        RECT 71.100 187.415 71.375 187.925 ;
        RECT 71.565 187.560 72.095 187.925 ;
        RECT 72.520 187.695 72.850 188.095 ;
        RECT 71.920 187.525 72.095 187.560 ;
        RECT 71.100 187.245 71.380 187.415 ;
        RECT 71.100 186.765 71.375 187.245 ;
        RECT 71.580 186.565 71.750 187.365 ;
        RECT 70.740 186.395 71.750 186.565 ;
        RECT 71.920 187.355 72.850 187.525 ;
        RECT 73.020 187.355 73.275 187.925 ;
        RECT 73.450 187.370 73.740 188.095 ;
        RECT 71.920 186.225 72.090 187.355 ;
        RECT 72.680 187.185 72.850 187.355 ;
        RECT 70.965 186.055 72.090 186.225 ;
        RECT 72.260 186.855 72.455 187.185 ;
        RECT 72.680 186.855 72.935 187.185 ;
        RECT 72.260 185.885 72.430 186.855 ;
        RECT 73.105 186.685 73.275 187.355 ;
        RECT 74.370 187.325 76.040 188.095 ;
        RECT 70.400 185.715 72.430 185.885 ;
        RECT 72.600 185.545 72.770 186.685 ;
        RECT 72.940 185.715 73.275 186.685 ;
        RECT 73.450 185.545 73.740 186.710 ;
        RECT 74.370 186.635 75.120 187.155 ;
        RECT 75.290 186.805 76.040 187.325 ;
        RECT 76.250 187.275 76.480 188.095 ;
        RECT 76.650 187.295 76.980 187.925 ;
        RECT 76.230 186.855 76.560 187.105 ;
        RECT 76.730 186.695 76.980 187.295 ;
        RECT 77.150 187.275 77.360 188.095 ;
        RECT 77.900 187.625 78.070 188.095 ;
        RECT 78.240 187.445 78.570 187.925 ;
        RECT 78.740 187.625 78.910 188.095 ;
        RECT 79.080 187.445 79.410 187.925 ;
        RECT 77.645 187.275 79.410 187.445 ;
        RECT 79.580 187.285 79.750 188.095 ;
        RECT 79.950 187.715 81.020 187.885 ;
        RECT 79.950 187.360 80.270 187.715 ;
        RECT 74.370 185.545 76.040 186.635 ;
        RECT 76.250 185.545 76.480 186.685 ;
        RECT 76.650 185.715 76.980 186.695 ;
        RECT 77.645 186.725 78.055 187.275 ;
        RECT 79.945 187.105 80.270 187.360 ;
        RECT 78.240 186.895 80.270 187.105 ;
        RECT 79.925 186.885 80.270 186.895 ;
        RECT 80.440 187.145 80.680 187.545 ;
        RECT 80.850 187.485 81.020 187.715 ;
        RECT 81.190 187.655 81.380 188.095 ;
        RECT 81.550 187.645 82.500 187.925 ;
        RECT 82.720 187.735 83.070 187.905 ;
        RECT 80.850 187.315 81.380 187.485 ;
        RECT 77.150 185.545 77.360 186.685 ;
        RECT 77.645 186.555 79.370 186.725 ;
        RECT 77.900 185.545 78.070 186.385 ;
        RECT 78.280 185.715 78.530 186.555 ;
        RECT 78.740 185.545 78.910 186.385 ;
        RECT 79.080 185.715 79.370 186.555 ;
        RECT 79.580 185.545 79.750 186.605 ;
        RECT 79.925 186.265 80.095 186.885 ;
        RECT 80.440 186.775 80.980 187.145 ;
        RECT 81.160 187.035 81.380 187.315 ;
        RECT 81.550 186.865 81.720 187.645 ;
        RECT 81.315 186.695 81.720 186.865 ;
        RECT 81.890 186.855 82.240 187.475 ;
        RECT 81.315 186.605 81.485 186.695 ;
        RECT 82.410 186.685 82.620 187.475 ;
        RECT 80.265 186.435 81.485 186.605 ;
        RECT 81.945 186.525 82.620 186.685 ;
        RECT 79.925 186.095 80.725 186.265 ;
        RECT 80.045 185.545 80.375 185.925 ;
        RECT 80.555 185.805 80.725 186.095 ;
        RECT 81.315 186.055 81.485 186.435 ;
        RECT 81.655 186.515 82.620 186.525 ;
        RECT 82.810 187.345 83.070 187.735 ;
        RECT 83.280 187.635 83.610 188.095 ;
        RECT 84.485 187.705 85.340 187.875 ;
        RECT 85.545 187.705 86.040 187.875 ;
        RECT 86.210 187.735 86.540 188.095 ;
        RECT 82.810 186.655 82.980 187.345 ;
        RECT 83.150 186.995 83.320 187.175 ;
        RECT 83.490 187.165 84.280 187.415 ;
        RECT 84.485 186.995 84.655 187.705 ;
        RECT 84.825 187.195 85.180 187.415 ;
        RECT 83.150 186.825 84.840 186.995 ;
        RECT 81.655 186.225 82.115 186.515 ;
        RECT 82.810 186.485 84.310 186.655 ;
        RECT 82.810 186.345 82.980 186.485 ;
        RECT 82.420 186.175 82.980 186.345 ;
        RECT 80.895 185.545 81.145 186.005 ;
        RECT 81.315 185.715 82.185 186.055 ;
        RECT 82.420 185.715 82.590 186.175 ;
        RECT 83.425 186.145 84.500 186.315 ;
        RECT 82.760 185.545 83.130 186.005 ;
        RECT 83.425 185.805 83.595 186.145 ;
        RECT 83.765 185.545 84.095 185.975 ;
        RECT 84.330 185.805 84.500 186.145 ;
        RECT 84.670 186.045 84.840 186.825 ;
        RECT 85.010 186.605 85.180 187.195 ;
        RECT 85.350 186.795 85.700 187.415 ;
        RECT 85.010 186.215 85.475 186.605 ;
        RECT 85.870 186.345 86.040 187.705 ;
        RECT 86.210 186.515 86.670 187.565 ;
        RECT 85.645 186.175 86.040 186.345 ;
        RECT 85.645 186.045 85.815 186.175 ;
        RECT 84.670 185.715 85.350 186.045 ;
        RECT 85.565 185.715 85.815 186.045 ;
        RECT 85.985 185.545 86.235 186.005 ;
        RECT 86.405 185.730 86.730 186.515 ;
        RECT 86.900 185.715 87.070 187.835 ;
        RECT 87.240 187.715 87.570 188.095 ;
        RECT 87.740 187.545 87.995 187.835 ;
        RECT 87.245 187.375 87.995 187.545 ;
        RECT 89.005 187.385 89.260 187.915 ;
        RECT 89.440 187.635 89.725 188.095 ;
        RECT 87.245 186.385 87.475 187.375 ;
        RECT 87.645 186.555 87.995 187.205 ;
        RECT 89.005 186.525 89.185 187.385 ;
        RECT 89.905 187.185 90.155 187.835 ;
        RECT 89.355 186.855 90.155 187.185 ;
        RECT 87.245 186.215 87.995 186.385 ;
        RECT 87.240 185.545 87.570 186.045 ;
        RECT 87.740 185.715 87.995 186.215 ;
        RECT 89.005 186.055 89.260 186.525 ;
        RECT 88.920 185.885 89.260 186.055 ;
        RECT 89.005 185.855 89.260 185.885 ;
        RECT 89.440 185.545 89.725 186.345 ;
        RECT 89.905 186.265 90.155 186.855 ;
        RECT 90.355 187.500 90.675 187.830 ;
        RECT 90.855 187.615 91.515 188.095 ;
        RECT 91.715 187.705 92.565 187.875 ;
        RECT 90.355 186.605 90.545 187.500 ;
        RECT 90.865 187.175 91.525 187.445 ;
        RECT 91.195 187.115 91.525 187.175 ;
        RECT 90.715 186.945 91.045 187.005 ;
        RECT 91.715 186.945 91.885 187.705 ;
        RECT 93.125 187.635 93.445 188.095 ;
        RECT 93.645 187.455 93.895 187.885 ;
        RECT 94.185 187.655 94.595 188.095 ;
        RECT 94.765 187.715 95.780 187.915 ;
        RECT 92.055 187.285 93.305 187.455 ;
        RECT 92.055 187.165 92.385 187.285 ;
        RECT 90.715 186.775 92.615 186.945 ;
        RECT 90.355 186.435 92.275 186.605 ;
        RECT 90.355 186.415 90.675 186.435 ;
        RECT 89.905 185.755 90.235 186.265 ;
        RECT 90.505 185.805 90.675 186.415 ;
        RECT 92.445 186.265 92.615 186.775 ;
        RECT 92.785 186.705 92.965 187.115 ;
        RECT 93.135 186.525 93.305 187.285 ;
        RECT 90.845 185.545 91.175 186.235 ;
        RECT 91.405 186.095 92.615 186.265 ;
        RECT 92.785 186.215 93.305 186.525 ;
        RECT 93.475 187.115 93.895 187.455 ;
        RECT 94.185 187.115 94.595 187.445 ;
        RECT 93.475 186.345 93.665 187.115 ;
        RECT 94.765 186.985 94.935 187.715 ;
        RECT 96.080 187.545 96.250 187.875 ;
        RECT 96.420 187.715 96.750 188.095 ;
        RECT 95.105 187.165 95.455 187.535 ;
        RECT 94.765 186.945 95.185 186.985 ;
        RECT 93.835 186.775 95.185 186.945 ;
        RECT 93.835 186.615 94.085 186.775 ;
        RECT 94.595 186.345 94.845 186.605 ;
        RECT 93.475 186.095 94.845 186.345 ;
        RECT 91.405 185.805 91.645 186.095 ;
        RECT 92.445 186.015 92.615 186.095 ;
        RECT 91.845 185.545 92.265 185.925 ;
        RECT 92.445 185.765 93.075 186.015 ;
        RECT 93.545 185.545 93.875 185.925 ;
        RECT 94.045 185.805 94.215 186.095 ;
        RECT 95.015 185.930 95.185 186.775 ;
        RECT 95.635 186.605 95.855 187.475 ;
        RECT 96.080 187.355 96.775 187.545 ;
        RECT 95.355 186.225 95.855 186.605 ;
        RECT 96.025 186.555 96.435 187.175 ;
        RECT 96.605 186.385 96.775 187.355 ;
        RECT 96.080 186.215 96.775 186.385 ;
        RECT 94.395 185.545 94.775 185.925 ;
        RECT 95.015 185.760 95.845 185.930 ;
        RECT 96.080 185.715 96.250 186.215 ;
        RECT 96.420 185.545 96.750 186.045 ;
        RECT 96.965 185.715 97.190 187.835 ;
        RECT 97.360 187.715 97.690 188.095 ;
        RECT 97.860 187.545 98.030 187.835 ;
        RECT 97.365 187.375 98.030 187.545 ;
        RECT 97.365 186.385 97.595 187.375 ;
        RECT 99.210 187.370 99.500 188.095 ;
        RECT 100.135 187.550 105.480 188.095 ;
        RECT 105.655 187.550 111.000 188.095 ;
        RECT 97.765 186.555 98.115 187.205 ;
        RECT 97.365 186.215 98.030 186.385 ;
        RECT 97.360 185.545 97.690 186.045 ;
        RECT 97.860 185.715 98.030 186.215 ;
        RECT 99.210 185.545 99.500 186.710 ;
        RECT 101.725 185.980 102.075 187.230 ;
        RECT 103.555 186.720 103.895 187.550 ;
        RECT 107.245 185.980 107.595 187.230 ;
        RECT 109.075 186.720 109.415 187.550 ;
        RECT 111.170 187.345 112.380 188.095 ;
        RECT 111.170 186.635 111.690 187.175 ;
        RECT 111.860 186.805 112.380 187.345 ;
        RECT 100.135 185.545 105.480 185.980 ;
        RECT 105.655 185.545 111.000 185.980 ;
        RECT 111.170 185.545 112.380 186.635 ;
        RECT 18.165 185.375 112.465 185.545 ;
        RECT 18.250 184.285 19.460 185.375 ;
        RECT 18.250 183.575 18.770 184.115 ;
        RECT 18.940 183.745 19.460 184.285 ;
        RECT 19.630 184.285 20.840 185.375 ;
        RECT 21.010 184.285 24.520 185.375 ;
        RECT 19.630 183.745 20.150 184.285 ;
        RECT 20.320 183.575 20.840 184.115 ;
        RECT 21.010 183.765 22.700 184.285 ;
        RECT 24.690 184.235 24.950 185.375 ;
        RECT 25.190 184.865 26.805 185.195 ;
        RECT 22.870 183.595 24.520 184.115 ;
        RECT 25.200 184.065 25.370 184.625 ;
        RECT 25.630 184.525 26.805 184.695 ;
        RECT 26.975 184.575 27.255 185.375 ;
        RECT 25.630 184.235 25.960 184.525 ;
        RECT 26.635 184.405 26.805 184.525 ;
        RECT 26.130 184.065 26.375 184.355 ;
        RECT 26.635 184.235 27.295 184.405 ;
        RECT 27.465 184.235 27.740 185.205 ;
        RECT 27.125 184.065 27.295 184.235 ;
        RECT 24.695 183.815 25.030 184.065 ;
        RECT 25.200 183.735 25.915 184.065 ;
        RECT 26.130 183.735 26.955 184.065 ;
        RECT 27.125 183.735 27.400 184.065 ;
        RECT 25.200 183.645 25.450 183.735 ;
        RECT 18.250 182.825 19.460 183.575 ;
        RECT 19.630 182.825 20.840 183.575 ;
        RECT 21.010 182.825 24.520 183.595 ;
        RECT 24.690 182.825 24.950 183.645 ;
        RECT 25.120 183.225 25.450 183.645 ;
        RECT 27.125 183.565 27.295 183.735 ;
        RECT 25.630 183.395 27.295 183.565 ;
        RECT 27.570 183.500 27.740 184.235 ;
        RECT 27.910 184.285 29.120 185.375 ;
        RECT 29.300 184.315 29.630 185.165 ;
        RECT 27.910 183.745 28.430 184.285 ;
        RECT 28.600 183.575 29.120 184.115 ;
        RECT 25.630 182.995 25.890 183.395 ;
        RECT 26.060 182.825 26.390 183.225 ;
        RECT 26.560 183.045 26.730 183.395 ;
        RECT 26.900 182.825 27.275 183.225 ;
        RECT 27.465 183.155 27.740 183.500 ;
        RECT 27.910 182.825 29.120 183.575 ;
        RECT 29.300 183.550 29.490 184.315 ;
        RECT 29.800 184.235 30.050 185.375 ;
        RECT 30.240 184.735 30.490 185.155 ;
        RECT 30.720 184.905 31.050 185.375 ;
        RECT 31.280 184.735 31.530 185.155 ;
        RECT 30.240 184.565 31.530 184.735 ;
        RECT 31.710 184.735 32.040 185.165 ;
        RECT 31.710 184.565 32.165 184.735 ;
        RECT 30.230 184.065 30.445 184.395 ;
        RECT 29.660 183.735 29.970 184.065 ;
        RECT 30.140 183.735 30.445 184.065 ;
        RECT 30.620 183.735 30.905 184.395 ;
        RECT 31.100 183.735 31.365 184.395 ;
        RECT 31.580 183.735 31.825 184.395 ;
        RECT 29.800 183.565 29.970 183.735 ;
        RECT 31.995 183.565 32.165 184.565 ;
        RECT 29.300 183.040 29.630 183.550 ;
        RECT 29.800 183.395 32.165 183.565 ;
        RECT 32.510 184.505 32.785 185.205 ;
        RECT 32.955 184.830 33.210 185.375 ;
        RECT 33.380 184.865 33.860 185.205 ;
        RECT 34.035 184.820 34.640 185.375 ;
        RECT 34.025 184.720 34.640 184.820 ;
        RECT 34.025 184.695 34.210 184.720 ;
        RECT 32.510 183.475 32.680 184.505 ;
        RECT 32.955 184.375 33.710 184.625 ;
        RECT 33.880 184.450 34.210 184.695 ;
        RECT 32.955 184.340 33.725 184.375 ;
        RECT 32.955 184.330 33.740 184.340 ;
        RECT 32.850 184.315 33.745 184.330 ;
        RECT 32.850 184.300 33.765 184.315 ;
        RECT 32.850 184.290 33.785 184.300 ;
        RECT 32.850 184.280 33.810 184.290 ;
        RECT 32.850 184.250 33.880 184.280 ;
        RECT 32.850 184.220 33.900 184.250 ;
        RECT 32.850 184.190 33.920 184.220 ;
        RECT 32.850 184.165 33.950 184.190 ;
        RECT 32.850 184.130 33.985 184.165 ;
        RECT 32.850 184.125 34.015 184.130 ;
        RECT 32.850 183.730 33.080 184.125 ;
        RECT 33.625 184.120 34.015 184.125 ;
        RECT 33.650 184.110 34.015 184.120 ;
        RECT 33.665 184.105 34.015 184.110 ;
        RECT 33.680 184.100 34.015 184.105 ;
        RECT 34.380 184.100 34.640 184.550 ;
        RECT 34.810 184.210 35.100 185.375 ;
        RECT 35.270 184.285 36.480 185.375 ;
        RECT 36.685 184.585 37.220 185.205 ;
        RECT 33.680 184.095 34.640 184.100 ;
        RECT 33.690 184.085 34.640 184.095 ;
        RECT 33.700 184.080 34.640 184.085 ;
        RECT 33.710 184.070 34.640 184.080 ;
        RECT 33.715 184.060 34.640 184.070 ;
        RECT 33.720 184.055 34.640 184.060 ;
        RECT 33.730 184.040 34.640 184.055 ;
        RECT 33.735 184.025 34.640 184.040 ;
        RECT 33.745 184.000 34.640 184.025 ;
        RECT 33.250 183.530 33.580 183.955 ;
        RECT 33.330 183.505 33.580 183.530 ;
        RECT 29.800 182.825 30.130 183.225 ;
        RECT 31.180 183.055 31.510 183.395 ;
        RECT 31.680 182.825 32.010 183.225 ;
        RECT 32.510 182.995 32.770 183.475 ;
        RECT 32.940 182.825 33.190 183.365 ;
        RECT 33.360 183.045 33.580 183.505 ;
        RECT 33.750 183.930 34.640 184.000 ;
        RECT 33.750 183.205 33.920 183.930 ;
        RECT 34.090 183.375 34.640 183.760 ;
        RECT 35.270 183.745 35.790 184.285 ;
        RECT 35.960 183.575 36.480 184.115 ;
        RECT 33.750 183.035 34.640 183.205 ;
        RECT 34.810 182.825 35.100 183.550 ;
        RECT 35.270 182.825 36.480 183.575 ;
        RECT 36.685 183.565 37.000 184.585 ;
        RECT 37.390 184.575 37.720 185.375 ;
        RECT 38.205 184.405 38.595 184.580 ;
        RECT 37.170 184.235 38.595 184.405 ;
        RECT 38.950 184.405 39.220 185.175 ;
        RECT 39.390 184.595 39.720 185.375 ;
        RECT 39.925 184.770 40.110 185.175 ;
        RECT 40.280 184.950 40.615 185.375 ;
        RECT 39.925 184.595 40.590 184.770 ;
        RECT 38.950 184.235 40.080 184.405 ;
        RECT 37.170 183.735 37.340 184.235 ;
        RECT 36.685 182.995 37.300 183.565 ;
        RECT 37.590 183.505 37.855 184.065 ;
        RECT 38.025 183.335 38.195 184.235 ;
        RECT 38.365 183.505 38.720 184.065 ;
        RECT 37.470 182.825 37.685 183.335 ;
        RECT 37.915 183.005 38.195 183.335 ;
        RECT 38.375 182.825 38.615 183.335 ;
        RECT 38.950 183.325 39.120 184.235 ;
        RECT 39.290 183.485 39.650 184.065 ;
        RECT 39.830 183.735 40.080 184.235 ;
        RECT 40.250 183.565 40.590 184.595 ;
        RECT 40.940 184.225 41.270 185.375 ;
        RECT 41.440 184.355 41.610 185.205 ;
        RECT 41.780 184.575 42.110 185.375 ;
        RECT 42.280 184.355 42.450 185.205 ;
        RECT 42.630 184.575 42.870 185.375 ;
        RECT 43.040 184.395 43.370 185.205 ;
        RECT 41.440 184.185 42.450 184.355 ;
        RECT 42.655 184.225 43.370 184.395 ;
        RECT 44.010 184.285 47.520 185.375 ;
        RECT 47.780 184.705 47.950 185.205 ;
        RECT 48.120 184.875 48.450 185.375 ;
        RECT 47.780 184.535 48.445 184.705 ;
        RECT 41.440 183.645 41.935 184.185 ;
        RECT 42.655 183.985 42.825 184.225 ;
        RECT 42.325 183.815 42.825 183.985 ;
        RECT 42.995 183.815 43.375 184.055 ;
        RECT 42.655 183.645 42.825 183.815 ;
        RECT 44.010 183.765 45.700 184.285 ;
        RECT 39.905 183.395 40.590 183.565 ;
        RECT 38.950 182.995 39.210 183.325 ;
        RECT 39.420 182.825 39.695 183.305 ;
        RECT 39.905 182.995 40.110 183.395 ;
        RECT 40.280 182.825 40.615 183.225 ;
        RECT 40.940 182.825 41.270 183.625 ;
        RECT 41.440 183.475 42.450 183.645 ;
        RECT 42.655 183.475 43.290 183.645 ;
        RECT 45.870 183.595 47.520 184.115 ;
        RECT 47.695 183.715 48.045 184.365 ;
        RECT 41.440 182.995 41.610 183.475 ;
        RECT 41.780 182.825 42.110 183.305 ;
        RECT 42.280 182.995 42.450 183.475 ;
        RECT 42.700 182.825 42.940 183.305 ;
        RECT 43.120 182.995 43.290 183.475 ;
        RECT 44.010 182.825 47.520 183.595 ;
        RECT 48.215 183.545 48.445 184.535 ;
        RECT 47.780 183.375 48.445 183.545 ;
        RECT 47.780 183.085 47.950 183.375 ;
        RECT 48.120 182.825 48.450 183.205 ;
        RECT 48.620 183.085 48.845 185.205 ;
        RECT 49.060 184.875 49.390 185.375 ;
        RECT 49.560 184.705 49.730 185.205 ;
        RECT 49.965 184.990 50.795 185.160 ;
        RECT 51.035 184.995 51.415 185.375 ;
        RECT 49.035 184.535 49.730 184.705 ;
        RECT 49.035 183.565 49.205 184.535 ;
        RECT 49.375 183.745 49.785 184.365 ;
        RECT 49.955 184.315 50.455 184.695 ;
        RECT 49.035 183.375 49.730 183.565 ;
        RECT 49.955 183.445 50.175 184.315 ;
        RECT 50.625 184.145 50.795 184.990 ;
        RECT 51.595 184.825 51.765 185.115 ;
        RECT 51.935 184.995 52.265 185.375 ;
        RECT 52.735 184.905 53.365 185.155 ;
        RECT 53.545 184.995 53.965 185.375 ;
        RECT 53.195 184.825 53.365 184.905 ;
        RECT 54.165 184.825 54.405 185.115 ;
        RECT 50.965 184.575 52.335 184.825 ;
        RECT 50.965 184.315 51.215 184.575 ;
        RECT 51.725 184.145 51.975 184.305 ;
        RECT 50.625 183.975 51.975 184.145 ;
        RECT 50.625 183.935 51.045 183.975 ;
        RECT 50.355 183.385 50.705 183.755 ;
        RECT 49.060 182.825 49.390 183.205 ;
        RECT 49.560 183.045 49.730 183.375 ;
        RECT 50.875 183.205 51.045 183.935 ;
        RECT 52.145 183.805 52.335 184.575 ;
        RECT 51.215 183.475 51.625 183.805 ;
        RECT 51.915 183.465 52.335 183.805 ;
        RECT 52.505 184.395 53.025 184.705 ;
        RECT 53.195 184.655 54.405 184.825 ;
        RECT 54.635 184.685 54.965 185.375 ;
        RECT 52.505 183.635 52.675 184.395 ;
        RECT 52.845 183.805 53.025 184.215 ;
        RECT 53.195 184.145 53.365 184.655 ;
        RECT 55.135 184.505 55.305 185.115 ;
        RECT 55.575 184.655 55.905 185.165 ;
        RECT 55.135 184.485 55.455 184.505 ;
        RECT 53.535 184.315 55.455 184.485 ;
        RECT 53.195 183.975 55.095 184.145 ;
        RECT 53.425 183.635 53.755 183.755 ;
        RECT 52.505 183.465 53.755 183.635 ;
        RECT 50.030 183.005 51.045 183.205 ;
        RECT 51.215 182.825 51.625 183.265 ;
        RECT 51.915 183.035 52.165 183.465 ;
        RECT 52.365 182.825 52.685 183.285 ;
        RECT 53.925 183.215 54.095 183.975 ;
        RECT 54.765 183.915 55.095 183.975 ;
        RECT 54.285 183.745 54.615 183.805 ;
        RECT 54.285 183.475 54.945 183.745 ;
        RECT 55.265 183.420 55.455 184.315 ;
        RECT 53.245 183.045 54.095 183.215 ;
        RECT 54.295 182.825 54.955 183.305 ;
        RECT 55.135 183.090 55.455 183.420 ;
        RECT 55.655 184.065 55.905 184.655 ;
        RECT 56.085 184.575 56.370 185.375 ;
        RECT 56.550 185.035 56.805 185.065 ;
        RECT 56.550 184.865 56.890 185.035 ;
        RECT 56.550 184.395 56.805 184.865 ;
        RECT 55.655 183.735 56.455 184.065 ;
        RECT 55.655 183.085 55.905 183.735 ;
        RECT 56.625 183.535 56.805 184.395 ;
        RECT 57.820 184.395 58.150 185.205 ;
        RECT 58.320 184.575 58.560 185.375 ;
        RECT 57.820 184.225 58.535 184.395 ;
        RECT 57.815 183.815 58.195 184.055 ;
        RECT 58.365 183.985 58.535 184.225 ;
        RECT 58.740 184.355 58.910 185.205 ;
        RECT 59.080 184.575 59.410 185.375 ;
        RECT 59.580 184.355 59.750 185.205 ;
        RECT 58.740 184.185 59.750 184.355 ;
        RECT 59.920 184.225 60.250 185.375 ;
        RECT 60.570 184.210 60.860 185.375 ;
        RECT 61.030 184.285 64.540 185.375 ;
        RECT 64.825 184.745 65.110 185.205 ;
        RECT 65.280 184.915 65.550 185.375 ;
        RECT 64.825 184.525 65.780 184.745 ;
        RECT 58.365 183.815 58.865 183.985 ;
        RECT 58.365 183.645 58.535 183.815 ;
        RECT 59.255 183.645 59.750 184.185 ;
        RECT 61.030 183.765 62.720 184.285 ;
        RECT 56.085 182.825 56.370 183.285 ;
        RECT 56.550 183.005 56.805 183.535 ;
        RECT 57.900 183.475 58.535 183.645 ;
        RECT 58.740 183.475 59.750 183.645 ;
        RECT 57.900 182.995 58.070 183.475 ;
        RECT 58.250 182.825 58.490 183.305 ;
        RECT 58.740 182.995 58.910 183.475 ;
        RECT 59.080 182.825 59.410 183.305 ;
        RECT 59.580 182.995 59.750 183.475 ;
        RECT 59.920 182.825 60.250 183.625 ;
        RECT 62.890 183.595 64.540 184.115 ;
        RECT 64.710 183.795 65.400 184.355 ;
        RECT 65.570 183.625 65.780 184.525 ;
        RECT 60.570 182.825 60.860 183.550 ;
        RECT 61.030 182.825 64.540 183.595 ;
        RECT 64.825 183.455 65.780 183.625 ;
        RECT 65.950 184.355 66.350 185.205 ;
        RECT 66.540 184.745 66.820 185.205 ;
        RECT 67.340 184.915 67.665 185.375 ;
        RECT 66.540 184.525 67.665 184.745 ;
        RECT 65.950 183.795 67.045 184.355 ;
        RECT 67.215 184.065 67.665 184.525 ;
        RECT 67.835 184.235 68.220 185.205 ;
        RECT 68.765 185.035 69.020 185.065 ;
        RECT 68.680 184.865 69.020 185.035 ;
        RECT 64.825 182.995 65.110 183.455 ;
        RECT 65.280 182.825 65.550 183.285 ;
        RECT 65.950 182.995 66.350 183.795 ;
        RECT 67.215 183.735 67.770 184.065 ;
        RECT 67.215 183.625 67.665 183.735 ;
        RECT 66.540 183.455 67.665 183.625 ;
        RECT 67.940 183.565 68.220 184.235 ;
        RECT 66.540 182.995 66.820 183.455 ;
        RECT 67.340 182.825 67.665 183.285 ;
        RECT 67.835 182.995 68.220 183.565 ;
        RECT 68.765 184.395 69.020 184.865 ;
        RECT 69.200 184.575 69.485 185.375 ;
        RECT 69.665 184.655 69.995 185.165 ;
        RECT 68.765 183.535 68.945 184.395 ;
        RECT 69.665 184.065 69.915 184.655 ;
        RECT 70.265 184.505 70.435 185.115 ;
        RECT 70.605 184.685 70.935 185.375 ;
        RECT 71.165 184.825 71.405 185.115 ;
        RECT 71.605 184.995 72.025 185.375 ;
        RECT 72.205 184.905 72.835 185.155 ;
        RECT 73.305 184.995 73.635 185.375 ;
        RECT 72.205 184.825 72.375 184.905 ;
        RECT 73.805 184.825 73.975 185.115 ;
        RECT 74.155 184.995 74.535 185.375 ;
        RECT 74.775 184.990 75.605 185.160 ;
        RECT 71.165 184.655 72.375 184.825 ;
        RECT 69.115 183.735 69.915 184.065 ;
        RECT 68.765 183.005 69.020 183.535 ;
        RECT 69.200 182.825 69.485 183.285 ;
        RECT 69.665 183.085 69.915 183.735 ;
        RECT 70.115 184.485 70.435 184.505 ;
        RECT 70.115 184.315 72.035 184.485 ;
        RECT 70.115 183.420 70.305 184.315 ;
        RECT 72.205 184.145 72.375 184.655 ;
        RECT 72.545 184.395 73.065 184.705 ;
        RECT 70.475 183.975 72.375 184.145 ;
        RECT 70.475 183.915 70.805 183.975 ;
        RECT 70.955 183.745 71.285 183.805 ;
        RECT 70.625 183.475 71.285 183.745 ;
        RECT 70.115 183.090 70.435 183.420 ;
        RECT 70.615 182.825 71.275 183.305 ;
        RECT 71.475 183.215 71.645 183.975 ;
        RECT 72.545 183.805 72.725 184.215 ;
        RECT 71.815 183.635 72.145 183.755 ;
        RECT 72.895 183.635 73.065 184.395 ;
        RECT 71.815 183.465 73.065 183.635 ;
        RECT 73.235 184.575 74.605 184.825 ;
        RECT 73.235 183.805 73.425 184.575 ;
        RECT 74.355 184.315 74.605 184.575 ;
        RECT 73.595 184.145 73.845 184.305 ;
        RECT 74.775 184.145 74.945 184.990 ;
        RECT 75.840 184.705 76.010 185.205 ;
        RECT 76.180 184.875 76.510 185.375 ;
        RECT 75.115 184.315 75.615 184.695 ;
        RECT 75.840 184.535 76.535 184.705 ;
        RECT 73.595 183.975 74.945 184.145 ;
        RECT 74.525 183.935 74.945 183.975 ;
        RECT 73.235 183.465 73.655 183.805 ;
        RECT 73.945 183.475 74.355 183.805 ;
        RECT 71.475 183.045 72.325 183.215 ;
        RECT 72.885 182.825 73.205 183.285 ;
        RECT 73.405 183.035 73.655 183.465 ;
        RECT 73.945 182.825 74.355 183.265 ;
        RECT 74.525 183.205 74.695 183.935 ;
        RECT 74.865 183.385 75.215 183.755 ;
        RECT 75.395 183.445 75.615 184.315 ;
        RECT 75.785 183.745 76.195 184.365 ;
        RECT 76.365 183.565 76.535 184.535 ;
        RECT 75.840 183.375 76.535 183.565 ;
        RECT 74.525 183.005 75.540 183.205 ;
        RECT 75.840 183.045 76.010 183.375 ;
        RECT 76.180 182.825 76.510 183.205 ;
        RECT 76.725 183.085 76.950 185.205 ;
        RECT 77.120 184.875 77.450 185.375 ;
        RECT 77.620 184.705 77.790 185.205 ;
        RECT 78.975 184.940 84.320 185.375 ;
        RECT 84.495 184.950 84.830 185.375 ;
        RECT 77.125 184.535 77.790 184.705 ;
        RECT 77.125 183.545 77.355 184.535 ;
        RECT 77.525 183.715 77.875 184.365 ;
        RECT 80.565 183.690 80.915 184.940 ;
        RECT 85.000 184.770 85.185 185.175 ;
        RECT 84.520 184.595 85.185 184.770 ;
        RECT 85.390 184.595 85.720 185.375 ;
        RECT 77.125 183.375 77.790 183.545 ;
        RECT 77.120 182.825 77.450 183.205 ;
        RECT 77.620 183.085 77.790 183.375 ;
        RECT 82.395 183.370 82.735 184.200 ;
        RECT 84.520 183.565 84.860 184.595 ;
        RECT 85.890 184.405 86.160 185.175 ;
        RECT 85.030 184.235 86.160 184.405 ;
        RECT 85.030 183.735 85.280 184.235 ;
        RECT 84.520 183.395 85.205 183.565 ;
        RECT 85.460 183.485 85.820 184.065 ;
        RECT 78.975 182.825 84.320 183.370 ;
        RECT 84.495 182.825 84.830 183.225 ;
        RECT 85.000 182.995 85.205 183.395 ;
        RECT 85.990 183.325 86.160 184.235 ;
        RECT 86.330 184.210 86.620 185.375 ;
        RECT 87.910 184.705 88.190 185.375 ;
        RECT 88.360 184.485 88.660 185.035 ;
        RECT 88.860 184.655 89.190 185.375 ;
        RECT 89.380 184.655 89.840 185.205 ;
        RECT 87.725 184.065 87.990 184.425 ;
        RECT 88.360 184.315 89.300 184.485 ;
        RECT 89.130 184.065 89.300 184.315 ;
        RECT 87.725 183.815 88.400 184.065 ;
        RECT 88.620 183.815 88.960 184.065 ;
        RECT 89.130 183.735 89.420 184.065 ;
        RECT 89.130 183.645 89.300 183.735 ;
        RECT 85.415 182.825 85.690 183.305 ;
        RECT 85.900 182.995 86.160 183.325 ;
        RECT 86.330 182.825 86.620 183.550 ;
        RECT 87.910 183.455 89.300 183.645 ;
        RECT 87.910 183.095 88.240 183.455 ;
        RECT 89.590 183.285 89.840 184.655 ;
        RECT 90.010 184.615 90.525 185.025 ;
        RECT 90.760 184.615 90.930 185.375 ;
        RECT 91.100 185.035 93.130 185.205 ;
        RECT 90.010 183.805 90.350 184.615 ;
        RECT 91.100 184.370 91.270 185.035 ;
        RECT 91.665 184.695 92.790 184.865 ;
        RECT 90.520 184.180 91.270 184.370 ;
        RECT 91.440 184.355 92.450 184.525 ;
        RECT 90.010 183.635 91.240 183.805 ;
        RECT 88.860 182.825 89.110 183.285 ;
        RECT 89.280 182.995 89.840 183.285 ;
        RECT 90.285 183.030 90.530 183.635 ;
        RECT 90.750 182.825 91.260 183.360 ;
        RECT 91.440 182.995 91.630 184.355 ;
        RECT 91.800 184.015 92.075 184.155 ;
        RECT 91.800 183.845 92.080 184.015 ;
        RECT 91.800 182.995 92.075 183.845 ;
        RECT 92.280 183.555 92.450 184.355 ;
        RECT 92.620 183.565 92.790 184.695 ;
        RECT 92.960 184.065 93.130 185.035 ;
        RECT 93.300 184.235 93.470 185.375 ;
        RECT 93.640 184.235 93.975 185.205 ;
        RECT 92.960 183.735 93.155 184.065 ;
        RECT 93.380 183.735 93.635 184.065 ;
        RECT 93.380 183.565 93.550 183.735 ;
        RECT 93.805 183.565 93.975 184.235 ;
        RECT 94.300 184.225 94.630 185.375 ;
        RECT 94.800 184.355 94.970 185.205 ;
        RECT 95.140 184.575 95.470 185.375 ;
        RECT 95.640 184.355 95.810 185.205 ;
        RECT 95.990 184.575 96.230 185.375 ;
        RECT 96.400 184.395 96.730 185.205 ;
        RECT 94.800 184.185 95.810 184.355 ;
        RECT 96.015 184.225 96.730 184.395 ;
        RECT 96.915 184.225 97.175 185.375 ;
        RECT 97.350 184.300 97.605 185.205 ;
        RECT 97.775 184.615 98.105 185.375 ;
        RECT 98.320 184.445 98.490 185.205 ;
        RECT 94.800 183.675 95.295 184.185 ;
        RECT 96.015 183.985 96.185 184.225 ;
        RECT 95.685 183.815 96.185 183.985 ;
        RECT 96.355 183.815 96.735 184.055 ;
        RECT 94.800 183.645 95.300 183.675 ;
        RECT 96.015 183.645 96.185 183.815 ;
        RECT 92.620 183.395 93.550 183.565 ;
        RECT 92.620 183.360 92.795 183.395 ;
        RECT 92.265 182.995 92.795 183.360 ;
        RECT 93.220 182.825 93.550 183.225 ;
        RECT 93.720 182.995 93.975 183.565 ;
        RECT 94.300 182.825 94.630 183.625 ;
        RECT 94.800 183.475 95.810 183.645 ;
        RECT 96.015 183.475 96.650 183.645 ;
        RECT 94.800 182.995 94.970 183.475 ;
        RECT 95.140 182.825 95.470 183.305 ;
        RECT 95.640 182.995 95.810 183.475 ;
        RECT 96.060 182.825 96.300 183.305 ;
        RECT 96.480 182.995 96.650 183.475 ;
        RECT 96.915 182.825 97.175 183.665 ;
        RECT 97.350 183.570 97.520 184.300 ;
        RECT 97.775 184.275 98.490 184.445 ;
        RECT 98.750 184.285 99.960 185.375 ;
        RECT 100.135 184.940 105.480 185.375 ;
        RECT 105.655 184.940 111.000 185.375 ;
        RECT 97.775 184.065 97.945 184.275 ;
        RECT 97.690 183.735 97.945 184.065 ;
        RECT 97.350 182.995 97.605 183.570 ;
        RECT 97.775 183.545 97.945 183.735 ;
        RECT 98.225 183.725 98.580 184.095 ;
        RECT 98.750 183.745 99.270 184.285 ;
        RECT 99.440 183.575 99.960 184.115 ;
        RECT 101.725 183.690 102.075 184.940 ;
        RECT 97.775 183.375 98.490 183.545 ;
        RECT 97.775 182.825 98.105 183.205 ;
        RECT 98.320 182.995 98.490 183.375 ;
        RECT 98.750 182.825 99.960 183.575 ;
        RECT 103.555 183.370 103.895 184.200 ;
        RECT 107.245 183.690 107.595 184.940 ;
        RECT 111.170 184.285 112.380 185.375 ;
        RECT 109.075 183.370 109.415 184.200 ;
        RECT 111.170 183.745 111.690 184.285 ;
        RECT 111.860 183.575 112.380 184.115 ;
        RECT 100.135 182.825 105.480 183.370 ;
        RECT 105.655 182.825 111.000 183.370 ;
        RECT 111.170 182.825 112.380 183.575 ;
        RECT 18.165 182.655 112.465 182.825 ;
        RECT 18.250 181.905 19.460 182.655 ;
        RECT 18.250 181.365 18.770 181.905 ;
        RECT 20.610 181.835 20.820 182.655 ;
        RECT 20.990 181.855 21.320 182.485 ;
        RECT 18.940 181.195 19.460 181.735 ;
        RECT 20.990 181.255 21.240 181.855 ;
        RECT 21.490 181.835 21.720 182.655 ;
        RECT 21.930 181.930 22.220 182.655 ;
        RECT 22.700 182.185 22.870 182.655 ;
        RECT 23.040 182.005 23.370 182.485 ;
        RECT 23.540 182.185 23.710 182.655 ;
        RECT 23.880 182.005 24.210 182.485 ;
        RECT 22.445 181.835 24.210 182.005 ;
        RECT 24.380 181.845 24.550 182.655 ;
        RECT 24.750 182.275 25.820 182.445 ;
        RECT 24.750 181.920 25.070 182.275 ;
        RECT 21.410 181.415 21.740 181.665 ;
        RECT 22.445 181.285 22.855 181.835 ;
        RECT 24.745 181.665 25.070 181.920 ;
        RECT 23.040 181.455 25.070 181.665 ;
        RECT 24.725 181.445 25.070 181.455 ;
        RECT 25.240 181.705 25.480 182.105 ;
        RECT 25.650 182.045 25.820 182.275 ;
        RECT 25.990 182.215 26.180 182.655 ;
        RECT 26.350 182.205 27.300 182.485 ;
        RECT 27.520 182.295 27.870 182.465 ;
        RECT 25.650 181.875 26.180 182.045 ;
        RECT 18.250 180.105 19.460 181.195 ;
        RECT 20.610 180.105 20.820 181.245 ;
        RECT 20.990 180.275 21.320 181.255 ;
        RECT 21.490 180.105 21.720 181.245 ;
        RECT 21.930 180.105 22.220 181.270 ;
        RECT 22.445 181.115 24.170 181.285 ;
        RECT 22.700 180.105 22.870 180.945 ;
        RECT 23.080 180.275 23.330 181.115 ;
        RECT 23.540 180.105 23.710 180.945 ;
        RECT 23.880 180.275 24.170 181.115 ;
        RECT 24.380 180.105 24.550 181.165 ;
        RECT 24.725 180.825 24.895 181.445 ;
        RECT 25.240 181.335 25.780 181.705 ;
        RECT 25.960 181.595 26.180 181.875 ;
        RECT 26.350 181.425 26.520 182.205 ;
        RECT 26.115 181.255 26.520 181.425 ;
        RECT 26.690 181.415 27.040 182.035 ;
        RECT 26.115 181.165 26.285 181.255 ;
        RECT 27.210 181.245 27.420 182.035 ;
        RECT 25.065 180.995 26.285 181.165 ;
        RECT 26.745 181.085 27.420 181.245 ;
        RECT 24.725 180.655 25.525 180.825 ;
        RECT 24.845 180.105 25.175 180.485 ;
        RECT 25.355 180.365 25.525 180.655 ;
        RECT 26.115 180.615 26.285 180.995 ;
        RECT 26.455 181.075 27.420 181.085 ;
        RECT 27.610 181.905 27.870 182.295 ;
        RECT 28.080 182.195 28.410 182.655 ;
        RECT 29.285 182.265 30.140 182.435 ;
        RECT 30.345 182.265 30.840 182.435 ;
        RECT 31.010 182.295 31.340 182.655 ;
        RECT 27.610 181.215 27.780 181.905 ;
        RECT 27.950 181.555 28.120 181.735 ;
        RECT 28.290 181.725 29.080 181.975 ;
        RECT 29.285 181.555 29.455 182.265 ;
        RECT 29.625 181.755 29.980 181.975 ;
        RECT 27.950 181.385 29.640 181.555 ;
        RECT 26.455 180.785 26.915 181.075 ;
        RECT 27.610 181.045 29.110 181.215 ;
        RECT 27.610 180.905 27.780 181.045 ;
        RECT 27.220 180.735 27.780 180.905 ;
        RECT 25.695 180.105 25.945 180.565 ;
        RECT 26.115 180.275 26.985 180.615 ;
        RECT 27.220 180.275 27.390 180.735 ;
        RECT 28.225 180.705 29.300 180.875 ;
        RECT 27.560 180.105 27.930 180.565 ;
        RECT 28.225 180.365 28.395 180.705 ;
        RECT 28.565 180.105 28.895 180.535 ;
        RECT 29.130 180.365 29.300 180.705 ;
        RECT 29.470 180.605 29.640 181.385 ;
        RECT 29.810 181.165 29.980 181.755 ;
        RECT 30.150 181.355 30.500 181.975 ;
        RECT 29.810 180.775 30.275 181.165 ;
        RECT 30.670 180.905 30.840 182.265 ;
        RECT 31.010 181.075 31.470 182.125 ;
        RECT 30.445 180.735 30.840 180.905 ;
        RECT 30.445 180.605 30.615 180.735 ;
        RECT 29.470 180.275 30.150 180.605 ;
        RECT 30.365 180.275 30.615 180.605 ;
        RECT 30.785 180.105 31.035 180.565 ;
        RECT 31.205 180.290 31.530 181.075 ;
        RECT 31.700 180.275 31.870 182.395 ;
        RECT 32.040 182.275 32.370 182.655 ;
        RECT 32.540 182.105 32.795 182.395 ;
        RECT 32.045 181.935 32.795 182.105 ;
        RECT 32.970 181.980 33.245 182.325 ;
        RECT 33.435 182.255 33.810 182.655 ;
        RECT 33.980 182.085 34.150 182.435 ;
        RECT 34.320 182.255 34.650 182.655 ;
        RECT 34.820 182.085 35.080 182.485 ;
        RECT 32.045 180.945 32.275 181.935 ;
        RECT 32.445 181.115 32.795 181.765 ;
        RECT 32.970 181.245 33.140 181.980 ;
        RECT 33.415 181.915 35.080 182.085 ;
        RECT 33.415 181.745 33.585 181.915 ;
        RECT 35.260 181.835 35.590 182.255 ;
        RECT 35.760 181.835 36.020 182.655 ;
        RECT 36.190 182.155 36.450 182.485 ;
        RECT 36.660 182.175 36.935 182.655 ;
        RECT 35.260 181.745 35.510 181.835 ;
        RECT 33.310 181.415 33.585 181.745 ;
        RECT 33.755 181.415 34.580 181.745 ;
        RECT 34.795 181.415 35.510 181.745 ;
        RECT 35.680 181.415 36.015 181.665 ;
        RECT 33.415 181.245 33.585 181.415 ;
        RECT 32.045 180.775 32.795 180.945 ;
        RECT 32.040 180.105 32.370 180.605 ;
        RECT 32.540 180.275 32.795 180.775 ;
        RECT 32.970 180.275 33.245 181.245 ;
        RECT 33.415 181.075 34.075 181.245 ;
        RECT 34.335 181.125 34.580 181.415 ;
        RECT 33.905 180.955 34.075 181.075 ;
        RECT 34.750 180.955 35.080 181.245 ;
        RECT 33.455 180.105 33.735 180.905 ;
        RECT 33.905 180.785 35.080 180.955 ;
        RECT 35.340 180.855 35.510 181.415 ;
        RECT 36.190 181.245 36.360 182.155 ;
        RECT 37.145 182.085 37.350 182.485 ;
        RECT 37.520 182.255 37.855 182.655 ;
        RECT 36.530 181.415 36.890 181.995 ;
        RECT 37.145 181.915 37.830 182.085 ;
        RECT 37.070 181.245 37.320 181.745 ;
        RECT 33.905 180.285 35.520 180.615 ;
        RECT 35.760 180.105 36.020 181.245 ;
        RECT 36.190 181.075 37.320 181.245 ;
        RECT 36.190 180.305 36.460 181.075 ;
        RECT 37.490 180.885 37.830 181.915 ;
        RECT 36.630 180.105 36.960 180.885 ;
        RECT 37.165 180.710 37.830 180.885 ;
        RECT 37.165 180.305 37.350 180.710 ;
        RECT 37.520 180.105 37.855 180.530 ;
        RECT 38.490 180.275 38.750 182.485 ;
        RECT 38.920 182.275 39.250 182.655 ;
        RECT 39.460 181.745 39.655 182.320 ;
        RECT 39.925 181.745 40.110 182.325 ;
        RECT 38.920 180.825 39.090 181.745 ;
        RECT 39.400 181.415 39.655 181.745 ;
        RECT 39.880 181.415 40.110 181.745 ;
        RECT 40.360 182.315 41.840 182.485 ;
        RECT 40.360 181.415 40.530 182.315 ;
        RECT 40.700 181.815 41.250 182.145 ;
        RECT 41.440 181.985 41.840 182.315 ;
        RECT 42.020 182.275 42.350 182.655 ;
        RECT 42.660 182.155 42.920 182.485 ;
        RECT 39.460 181.105 39.655 181.415 ;
        RECT 39.925 181.105 40.110 181.415 ;
        RECT 40.700 180.825 40.870 181.815 ;
        RECT 41.440 181.505 41.610 181.985 ;
        RECT 42.190 181.795 42.400 181.975 ;
        RECT 41.780 181.625 42.400 181.795 ;
        RECT 38.920 180.655 40.870 180.825 ;
        RECT 41.040 181.335 41.610 181.505 ;
        RECT 42.750 181.455 42.920 182.155 ;
        RECT 44.010 181.885 47.520 182.655 ;
        RECT 47.690 181.930 47.980 182.655 ;
        RECT 41.040 180.825 41.210 181.335 ;
        RECT 41.790 181.285 42.920 181.455 ;
        RECT 41.790 181.165 41.960 181.285 ;
        RECT 41.380 180.995 41.960 181.165 ;
        RECT 41.040 180.655 41.780 180.825 ;
        RECT 42.230 180.785 42.580 181.115 ;
        RECT 38.920 180.105 39.250 180.485 ;
        RECT 39.675 180.275 39.845 180.655 ;
        RECT 40.105 180.105 40.435 180.485 ;
        RECT 40.630 180.275 40.800 180.655 ;
        RECT 41.010 180.105 41.340 180.485 ;
        RECT 41.590 180.275 41.780 180.655 ;
        RECT 42.750 180.605 42.920 181.285 ;
        RECT 42.020 180.105 42.350 180.485 ;
        RECT 42.660 180.275 42.920 180.605 ;
        RECT 44.010 181.195 45.700 181.715 ;
        RECT 45.870 181.365 47.520 181.885 ;
        RECT 48.885 181.845 49.130 182.450 ;
        RECT 49.350 182.120 49.860 182.655 ;
        RECT 48.610 181.675 49.840 181.845 ;
        RECT 44.010 180.105 47.520 181.195 ;
        RECT 47.690 180.105 47.980 181.270 ;
        RECT 48.610 180.865 48.950 181.675 ;
        RECT 49.120 181.110 49.870 181.300 ;
        RECT 48.610 180.455 49.125 180.865 ;
        RECT 49.360 180.105 49.530 180.865 ;
        RECT 49.700 180.445 49.870 181.110 ;
        RECT 50.040 181.125 50.230 182.485 ;
        RECT 50.400 181.635 50.675 182.485 ;
        RECT 50.865 182.120 51.395 182.485 ;
        RECT 51.820 182.255 52.150 182.655 ;
        RECT 51.220 182.085 51.395 182.120 ;
        RECT 50.400 181.465 50.680 181.635 ;
        RECT 50.400 181.325 50.675 181.465 ;
        RECT 50.880 181.125 51.050 181.925 ;
        RECT 50.040 180.955 51.050 181.125 ;
        RECT 51.220 181.915 52.150 182.085 ;
        RECT 52.320 181.915 52.575 182.485 ;
        RECT 51.220 180.785 51.390 181.915 ;
        RECT 51.980 181.745 52.150 181.915 ;
        RECT 50.265 180.615 51.390 180.785 ;
        RECT 51.560 181.415 51.755 181.745 ;
        RECT 51.980 181.415 52.235 181.745 ;
        RECT 51.560 180.445 51.730 181.415 ;
        RECT 52.405 181.245 52.575 181.915 ;
        RECT 52.750 181.905 53.960 182.655 ;
        RECT 49.700 180.275 51.730 180.445 ;
        RECT 51.900 180.105 52.070 181.245 ;
        RECT 52.240 180.275 52.575 181.245 ;
        RECT 52.750 181.195 53.270 181.735 ;
        RECT 53.440 181.365 53.960 181.905 ;
        RECT 54.130 181.980 54.400 182.325 ;
        RECT 54.590 182.255 54.970 182.655 ;
        RECT 55.140 182.085 55.310 182.435 ;
        RECT 55.480 182.255 55.810 182.655 ;
        RECT 56.010 182.085 56.180 182.435 ;
        RECT 56.380 182.155 56.710 182.655 ;
        RECT 56.890 182.195 57.450 182.485 ;
        RECT 57.620 182.195 57.870 182.655 ;
        RECT 54.130 181.245 54.300 181.980 ;
        RECT 54.570 181.915 56.180 182.085 ;
        RECT 54.570 181.745 54.740 181.915 ;
        RECT 54.470 181.415 54.740 181.745 ;
        RECT 54.910 181.415 55.315 181.745 ;
        RECT 54.570 181.245 54.740 181.415 ;
        RECT 55.485 181.295 56.195 181.745 ;
        RECT 56.365 181.415 56.715 181.985 ;
        RECT 52.750 180.105 53.960 181.195 ;
        RECT 54.130 180.275 54.400 181.245 ;
        RECT 54.570 181.075 55.295 181.245 ;
        RECT 55.485 181.125 56.200 181.295 ;
        RECT 55.125 180.955 55.295 181.075 ;
        RECT 56.395 180.955 56.715 181.245 ;
        RECT 54.610 180.105 54.890 180.905 ;
        RECT 55.125 180.785 56.715 180.955 ;
        RECT 56.890 180.825 57.140 182.195 ;
        RECT 58.490 182.025 58.820 182.385 ;
        RECT 57.430 181.835 58.820 182.025 ;
        RECT 60.170 181.835 60.380 182.655 ;
        RECT 60.550 181.855 60.880 182.485 ;
        RECT 57.430 181.745 57.600 181.835 ;
        RECT 57.310 181.415 57.600 181.745 ;
        RECT 57.770 181.415 58.110 181.665 ;
        RECT 58.330 181.415 59.005 181.665 ;
        RECT 57.430 181.165 57.600 181.415 ;
        RECT 57.430 180.995 58.370 181.165 ;
        RECT 58.740 181.055 59.005 181.415 ;
        RECT 60.550 181.255 60.800 181.855 ;
        RECT 61.050 181.835 61.280 182.655 ;
        RECT 61.495 181.945 61.750 182.475 ;
        RECT 61.920 182.195 62.225 182.655 ;
        RECT 62.470 182.275 63.540 182.445 ;
        RECT 60.970 181.415 61.300 181.665 ;
        RECT 61.495 181.295 61.705 181.945 ;
        RECT 62.470 181.920 62.790 182.275 ;
        RECT 62.465 181.745 62.790 181.920 ;
        RECT 61.875 181.445 62.790 181.745 ;
        RECT 62.960 181.705 63.200 182.105 ;
        RECT 63.370 182.045 63.540 182.275 ;
        RECT 63.710 182.215 63.900 182.655 ;
        RECT 64.070 182.205 65.020 182.485 ;
        RECT 65.240 182.295 65.590 182.465 ;
        RECT 63.370 181.875 63.900 182.045 ;
        RECT 61.875 181.415 62.615 181.445 ;
        RECT 55.060 180.325 56.715 180.615 ;
        RECT 56.890 180.275 57.350 180.825 ;
        RECT 57.540 180.105 57.870 180.825 ;
        RECT 58.070 180.445 58.370 180.995 ;
        RECT 58.540 180.105 58.820 180.775 ;
        RECT 60.170 180.105 60.380 181.245 ;
        RECT 60.550 180.275 60.880 181.255 ;
        RECT 61.050 180.105 61.280 181.245 ;
        RECT 61.495 180.415 61.750 181.295 ;
        RECT 61.920 180.105 62.225 181.245 ;
        RECT 62.445 180.825 62.615 181.415 ;
        RECT 62.960 181.335 63.500 181.705 ;
        RECT 63.680 181.595 63.900 181.875 ;
        RECT 64.070 181.425 64.240 182.205 ;
        RECT 63.835 181.255 64.240 181.425 ;
        RECT 64.410 181.415 64.760 182.035 ;
        RECT 63.835 181.165 64.005 181.255 ;
        RECT 64.930 181.245 65.140 182.035 ;
        RECT 62.785 180.995 64.005 181.165 ;
        RECT 64.465 181.085 65.140 181.245 ;
        RECT 62.445 180.655 63.245 180.825 ;
        RECT 62.565 180.105 62.895 180.485 ;
        RECT 63.075 180.365 63.245 180.655 ;
        RECT 63.835 180.615 64.005 180.995 ;
        RECT 64.175 181.075 65.140 181.085 ;
        RECT 65.330 181.905 65.590 182.295 ;
        RECT 65.800 182.195 66.130 182.655 ;
        RECT 67.005 182.265 67.860 182.435 ;
        RECT 68.065 182.265 68.560 182.435 ;
        RECT 68.730 182.295 69.060 182.655 ;
        RECT 65.330 181.215 65.500 181.905 ;
        RECT 65.670 181.555 65.840 181.735 ;
        RECT 66.010 181.725 66.800 181.975 ;
        RECT 67.005 181.555 67.175 182.265 ;
        RECT 67.345 181.755 67.700 181.975 ;
        RECT 65.670 181.385 67.360 181.555 ;
        RECT 64.175 180.785 64.635 181.075 ;
        RECT 65.330 181.045 66.830 181.215 ;
        RECT 65.330 180.905 65.500 181.045 ;
        RECT 64.940 180.735 65.500 180.905 ;
        RECT 63.415 180.105 63.665 180.565 ;
        RECT 63.835 180.275 64.705 180.615 ;
        RECT 64.940 180.275 65.110 180.735 ;
        RECT 65.945 180.705 67.020 180.875 ;
        RECT 65.280 180.105 65.650 180.565 ;
        RECT 65.945 180.365 66.115 180.705 ;
        RECT 66.285 180.105 66.615 180.535 ;
        RECT 66.850 180.365 67.020 180.705 ;
        RECT 67.190 180.605 67.360 181.385 ;
        RECT 67.530 181.165 67.700 181.755 ;
        RECT 67.870 181.355 68.220 181.975 ;
        RECT 67.530 180.775 67.995 181.165 ;
        RECT 68.390 180.905 68.560 182.265 ;
        RECT 68.730 181.075 69.190 182.125 ;
        RECT 68.165 180.735 68.560 180.905 ;
        RECT 68.165 180.605 68.335 180.735 ;
        RECT 67.190 180.275 67.870 180.605 ;
        RECT 68.085 180.275 68.335 180.605 ;
        RECT 68.505 180.105 68.755 180.565 ;
        RECT 68.925 180.290 69.250 181.075 ;
        RECT 69.420 180.275 69.590 182.395 ;
        RECT 69.760 182.275 70.090 182.655 ;
        RECT 70.260 182.105 70.515 182.395 ;
        RECT 69.765 181.935 70.515 182.105 ;
        RECT 70.690 182.195 71.250 182.485 ;
        RECT 71.420 182.195 71.670 182.655 ;
        RECT 69.765 180.945 69.995 181.935 ;
        RECT 70.165 181.115 70.515 181.765 ;
        RECT 69.765 180.775 70.515 180.945 ;
        RECT 69.760 180.105 70.090 180.605 ;
        RECT 70.260 180.275 70.515 180.775 ;
        RECT 70.690 180.825 70.940 182.195 ;
        RECT 72.290 182.025 72.620 182.385 ;
        RECT 71.230 181.835 72.620 182.025 ;
        RECT 73.450 181.930 73.740 182.655 ;
        RECT 75.105 181.845 75.350 182.450 ;
        RECT 75.570 182.120 76.080 182.655 ;
        RECT 71.230 181.745 71.400 181.835 ;
        RECT 71.110 181.415 71.400 181.745 ;
        RECT 74.830 181.675 76.060 181.845 ;
        RECT 71.570 181.415 71.910 181.665 ;
        RECT 72.130 181.415 72.805 181.665 ;
        RECT 71.230 181.165 71.400 181.415 ;
        RECT 71.230 180.995 72.170 181.165 ;
        RECT 72.540 181.055 72.805 181.415 ;
        RECT 70.690 180.275 71.150 180.825 ;
        RECT 71.340 180.105 71.670 180.825 ;
        RECT 71.870 180.445 72.170 180.995 ;
        RECT 72.340 180.105 72.620 180.775 ;
        RECT 73.450 180.105 73.740 181.270 ;
        RECT 74.830 180.865 75.170 181.675 ;
        RECT 75.340 181.110 76.090 181.300 ;
        RECT 74.830 180.455 75.345 180.865 ;
        RECT 75.580 180.105 75.750 180.865 ;
        RECT 75.920 180.445 76.090 181.110 ;
        RECT 76.260 181.125 76.450 182.485 ;
        RECT 76.620 181.975 76.895 182.485 ;
        RECT 77.085 182.120 77.615 182.485 ;
        RECT 78.040 182.255 78.370 182.655 ;
        RECT 77.440 182.085 77.615 182.120 ;
        RECT 76.620 181.805 76.900 181.975 ;
        RECT 76.620 181.325 76.895 181.805 ;
        RECT 77.100 181.125 77.270 181.925 ;
        RECT 76.260 180.955 77.270 181.125 ;
        RECT 77.440 181.915 78.370 182.085 ;
        RECT 78.540 181.915 78.795 182.485 ;
        RECT 77.440 180.785 77.610 181.915 ;
        RECT 78.200 181.745 78.370 181.915 ;
        RECT 76.485 180.615 77.610 180.785 ;
        RECT 77.780 181.415 77.975 181.745 ;
        RECT 78.200 181.415 78.455 181.745 ;
        RECT 77.780 180.445 77.950 181.415 ;
        RECT 78.625 181.245 78.795 181.915 ;
        RECT 79.010 181.835 79.240 182.655 ;
        RECT 79.410 181.855 79.740 182.485 ;
        RECT 78.990 181.415 79.320 181.665 ;
        RECT 79.490 181.255 79.740 181.855 ;
        RECT 79.910 181.835 80.120 182.655 ;
        RECT 80.350 181.905 81.560 182.655 ;
        RECT 75.920 180.275 77.950 180.445 ;
        RECT 78.120 180.105 78.290 181.245 ;
        RECT 78.460 180.275 78.795 181.245 ;
        RECT 79.010 180.105 79.240 181.245 ;
        RECT 79.410 180.275 79.740 181.255 ;
        RECT 79.910 180.105 80.120 181.245 ;
        RECT 80.350 181.195 80.870 181.735 ;
        RECT 81.040 181.365 81.560 181.905 ;
        RECT 81.930 182.025 82.260 182.385 ;
        RECT 82.880 182.195 83.130 182.655 ;
        RECT 83.300 182.195 83.860 182.485 ;
        RECT 81.930 181.835 83.320 182.025 ;
        RECT 83.150 181.745 83.320 181.835 ;
        RECT 81.745 181.415 82.420 181.665 ;
        RECT 82.640 181.415 82.980 181.665 ;
        RECT 83.150 181.415 83.440 181.745 ;
        RECT 80.350 180.105 81.560 181.195 ;
        RECT 81.745 181.055 82.010 181.415 ;
        RECT 83.150 181.165 83.320 181.415 ;
        RECT 82.380 180.995 83.320 181.165 ;
        RECT 81.930 180.105 82.210 180.775 ;
        RECT 82.380 180.445 82.680 180.995 ;
        RECT 83.610 180.825 83.860 182.195 ;
        RECT 82.880 180.105 83.210 180.825 ;
        RECT 83.400 180.275 83.860 180.825 ;
        RECT 84.030 181.855 84.370 182.485 ;
        RECT 84.540 181.855 84.790 182.655 ;
        RECT 84.980 182.005 85.310 182.485 ;
        RECT 85.480 182.195 85.705 182.655 ;
        RECT 85.875 182.005 86.205 182.485 ;
        RECT 84.030 181.245 84.205 181.855 ;
        RECT 84.980 181.835 86.205 182.005 ;
        RECT 86.835 181.875 87.335 182.485 ;
        RECT 88.170 181.980 88.440 182.325 ;
        RECT 88.630 182.255 89.010 182.655 ;
        RECT 89.180 182.085 89.350 182.435 ;
        RECT 89.520 182.255 89.850 182.655 ;
        RECT 90.050 182.085 90.220 182.435 ;
        RECT 90.420 182.155 90.750 182.655 ;
        RECT 84.375 181.495 85.070 181.665 ;
        RECT 84.900 181.245 85.070 181.495 ;
        RECT 85.245 181.465 85.665 181.665 ;
        RECT 85.835 181.465 86.165 181.665 ;
        RECT 86.335 181.465 86.665 181.665 ;
        RECT 86.835 181.245 87.005 181.875 ;
        RECT 87.190 181.415 87.540 181.665 ;
        RECT 88.170 181.245 88.340 181.980 ;
        RECT 88.610 181.915 90.220 182.085 ;
        RECT 88.610 181.745 88.780 181.915 ;
        RECT 88.510 181.415 88.780 181.745 ;
        RECT 88.950 181.415 89.355 181.745 ;
        RECT 88.610 181.245 88.780 181.415 ;
        RECT 84.030 180.275 84.370 181.245 ;
        RECT 84.540 180.105 84.710 181.245 ;
        RECT 84.900 181.075 87.335 181.245 ;
        RECT 84.980 180.105 85.230 180.905 ;
        RECT 85.875 180.275 86.205 181.075 ;
        RECT 86.505 180.105 86.835 180.905 ;
        RECT 87.005 180.275 87.335 181.075 ;
        RECT 88.170 180.275 88.440 181.245 ;
        RECT 88.610 181.075 89.335 181.245 ;
        RECT 89.525 181.125 90.235 181.745 ;
        RECT 90.405 181.415 90.755 181.985 ;
        RECT 90.970 181.835 91.200 182.655 ;
        RECT 91.370 181.855 91.700 182.485 ;
        RECT 90.950 181.415 91.280 181.665 ;
        RECT 91.450 181.255 91.700 181.855 ;
        RECT 91.870 181.835 92.080 182.655 ;
        RECT 92.310 181.855 92.650 182.485 ;
        RECT 92.820 181.855 93.070 182.655 ;
        RECT 93.260 182.005 93.590 182.485 ;
        RECT 93.760 182.195 93.985 182.655 ;
        RECT 94.155 182.005 94.485 182.485 ;
        RECT 89.165 180.955 89.335 181.075 ;
        RECT 90.435 180.955 90.755 181.245 ;
        RECT 88.650 180.105 88.930 180.905 ;
        RECT 89.165 180.785 90.755 180.955 ;
        RECT 89.100 180.325 90.755 180.615 ;
        RECT 90.970 180.105 91.200 181.245 ;
        RECT 91.370 180.275 91.700 181.255 ;
        RECT 92.310 181.805 92.540 181.855 ;
        RECT 93.260 181.835 94.485 182.005 ;
        RECT 95.115 181.875 95.615 182.485 ;
        RECT 96.450 181.885 99.040 182.655 ;
        RECT 99.210 181.930 99.500 182.655 ;
        RECT 100.135 182.110 105.480 182.655 ;
        RECT 105.655 182.110 111.000 182.655 ;
        RECT 92.310 181.245 92.485 181.805 ;
        RECT 92.655 181.495 93.350 181.665 ;
        RECT 93.180 181.245 93.350 181.495 ;
        RECT 93.525 181.465 93.945 181.665 ;
        RECT 94.115 181.465 94.445 181.665 ;
        RECT 94.615 181.465 94.945 181.665 ;
        RECT 95.115 181.245 95.285 181.875 ;
        RECT 95.470 181.415 95.820 181.665 ;
        RECT 91.870 180.105 92.080 181.245 ;
        RECT 92.310 180.275 92.650 181.245 ;
        RECT 92.820 180.105 92.990 181.245 ;
        RECT 93.180 181.075 95.615 181.245 ;
        RECT 93.260 180.105 93.510 180.905 ;
        RECT 94.155 180.275 94.485 181.075 ;
        RECT 94.785 180.105 95.115 180.905 ;
        RECT 95.285 180.275 95.615 181.075 ;
        RECT 96.450 181.195 97.660 181.715 ;
        RECT 97.830 181.365 99.040 181.885 ;
        RECT 96.450 180.105 99.040 181.195 ;
        RECT 99.210 180.105 99.500 181.270 ;
        RECT 101.725 180.540 102.075 181.790 ;
        RECT 103.555 181.280 103.895 182.110 ;
        RECT 107.245 180.540 107.595 181.790 ;
        RECT 109.075 181.280 109.415 182.110 ;
        RECT 111.170 181.905 112.380 182.655 ;
        RECT 111.170 181.195 111.690 181.735 ;
        RECT 111.860 181.365 112.380 181.905 ;
        RECT 100.135 180.105 105.480 180.540 ;
        RECT 105.655 180.105 111.000 180.540 ;
        RECT 111.170 180.105 112.380 181.195 ;
        RECT 18.165 179.935 112.465 180.105 ;
        RECT 18.250 178.845 19.460 179.935 ;
        RECT 20.110 179.135 20.390 179.935 ;
        RECT 20.590 178.965 20.920 179.765 ;
        RECT 21.120 179.135 21.290 179.935 ;
        RECT 21.460 178.965 21.790 179.765 ;
        RECT 18.250 178.135 18.770 178.675 ;
        RECT 18.940 178.305 19.460 178.845 ;
        RECT 20.090 178.295 20.330 178.965 ;
        RECT 20.510 178.795 21.790 178.965 ;
        RECT 21.960 178.795 22.220 179.935 ;
        RECT 22.505 179.305 22.790 179.765 ;
        RECT 22.960 179.475 23.230 179.935 ;
        RECT 22.505 179.085 23.460 179.305 ;
        RECT 18.250 177.385 19.460 178.135 ;
        RECT 20.510 178.125 20.680 178.795 ;
        RECT 20.850 178.295 21.160 178.625 ;
        RECT 21.330 178.295 21.710 178.625 ;
        RECT 21.910 178.295 22.195 178.625 ;
        RECT 22.390 178.355 23.080 178.915 ;
        RECT 20.955 178.125 21.160 178.295 ;
        RECT 20.090 177.555 20.785 178.125 ;
        RECT 20.955 177.600 21.305 178.125 ;
        RECT 21.495 177.600 21.710 178.295 ;
        RECT 23.250 178.185 23.460 179.085 ;
        RECT 21.880 177.385 22.215 178.125 ;
        RECT 22.505 178.015 23.460 178.185 ;
        RECT 23.630 178.915 24.030 179.765 ;
        RECT 24.220 179.305 24.500 179.765 ;
        RECT 25.020 179.475 25.345 179.935 ;
        RECT 24.220 179.085 25.345 179.305 ;
        RECT 23.630 178.355 24.725 178.915 ;
        RECT 24.895 178.625 25.345 179.085 ;
        RECT 25.515 178.795 25.900 179.765 ;
        RECT 22.505 177.555 22.790 178.015 ;
        RECT 22.960 177.385 23.230 177.845 ;
        RECT 23.630 177.555 24.030 178.355 ;
        RECT 24.895 178.295 25.450 178.625 ;
        RECT 24.895 178.185 25.345 178.295 ;
        RECT 24.220 178.015 25.345 178.185 ;
        RECT 25.620 178.125 25.900 178.795 ;
        RECT 26.070 178.845 27.740 179.935 ;
        RECT 27.910 179.425 28.210 179.935 ;
        RECT 28.380 179.255 28.710 179.765 ;
        RECT 28.880 179.425 29.510 179.935 ;
        RECT 30.090 179.425 30.470 179.595 ;
        RECT 30.640 179.425 30.940 179.935 ;
        RECT 30.300 179.255 30.470 179.425 ;
        RECT 27.910 179.085 30.130 179.255 ;
        RECT 26.070 178.325 26.820 178.845 ;
        RECT 26.990 178.155 27.740 178.675 ;
        RECT 24.220 177.555 24.500 178.015 ;
        RECT 25.020 177.385 25.345 177.845 ;
        RECT 25.515 177.555 25.900 178.125 ;
        RECT 26.070 177.385 27.740 178.155 ;
        RECT 27.910 178.125 28.080 179.085 ;
        RECT 28.250 178.745 29.790 178.915 ;
        RECT 28.250 178.295 28.495 178.745 ;
        RECT 28.755 178.375 29.450 178.575 ;
        RECT 29.620 178.545 29.790 178.745 ;
        RECT 29.960 178.885 30.130 179.085 ;
        RECT 30.300 179.055 30.960 179.255 ;
        RECT 29.960 178.715 30.620 178.885 ;
        RECT 29.620 178.375 30.220 178.545 ;
        RECT 30.450 178.295 30.620 178.715 ;
        RECT 27.910 177.580 28.375 178.125 ;
        RECT 28.880 177.385 29.050 178.205 ;
        RECT 29.220 178.125 30.130 178.205 ;
        RECT 30.790 178.125 30.960 179.055 ;
        RECT 29.220 178.035 30.470 178.125 ;
        RECT 29.220 177.555 29.550 178.035 ;
        RECT 29.960 177.955 30.470 178.035 ;
        RECT 29.720 177.385 30.070 177.775 ;
        RECT 30.240 177.555 30.470 177.955 ;
        RECT 30.640 177.645 30.960 178.125 ;
        RECT 31.590 178.125 31.850 179.750 ;
        RECT 33.600 179.485 33.930 179.935 ;
        RECT 32.030 179.095 34.640 179.305 ;
        RECT 32.030 178.295 32.250 179.095 ;
        RECT 32.490 178.295 32.790 178.915 ;
        RECT 32.960 178.295 33.290 178.915 ;
        RECT 33.460 178.295 33.780 178.915 ;
        RECT 33.950 178.295 34.300 178.915 ;
        RECT 34.470 178.125 34.640 179.095 ;
        RECT 34.810 178.770 35.100 179.935 ;
        RECT 31.590 177.955 33.430 178.125 ;
        RECT 31.860 177.385 32.190 177.780 ;
        RECT 32.360 177.600 32.560 177.955 ;
        RECT 32.730 177.385 33.060 177.785 ;
        RECT 33.230 177.610 33.430 177.955 ;
        RECT 33.600 177.385 33.930 178.125 ;
        RECT 34.165 177.955 34.640 178.125 ;
        RECT 36.190 178.125 36.450 179.750 ;
        RECT 38.200 179.485 38.530 179.935 ;
        RECT 39.410 179.435 39.670 179.765 ;
        RECT 39.980 179.555 40.310 179.935 ;
        RECT 36.630 179.095 39.240 179.305 ;
        RECT 36.630 178.295 36.850 179.095 ;
        RECT 37.090 178.295 37.390 178.915 ;
        RECT 37.560 178.295 37.890 178.915 ;
        RECT 38.060 178.295 38.380 178.915 ;
        RECT 38.550 178.295 38.900 178.915 ;
        RECT 39.070 178.125 39.240 179.095 ;
        RECT 34.165 177.705 34.335 177.955 ;
        RECT 34.810 177.385 35.100 178.110 ;
        RECT 36.190 177.955 38.030 178.125 ;
        RECT 36.460 177.385 36.790 177.780 ;
        RECT 36.960 177.600 37.160 177.955 ;
        RECT 37.330 177.385 37.660 177.785 ;
        RECT 37.830 177.610 38.030 177.955 ;
        RECT 38.200 177.385 38.530 178.125 ;
        RECT 38.765 177.955 39.240 178.125 ;
        RECT 39.410 178.755 39.580 179.435 ;
        RECT 40.550 179.385 40.740 179.765 ;
        RECT 40.990 179.555 41.320 179.935 ;
        RECT 41.530 179.385 41.700 179.765 ;
        RECT 41.895 179.555 42.225 179.935 ;
        RECT 42.485 179.385 42.655 179.765 ;
        RECT 43.080 179.555 43.410 179.935 ;
        RECT 39.750 178.925 40.100 179.255 ;
        RECT 40.550 179.215 41.290 179.385 ;
        RECT 40.370 178.875 40.950 179.045 ;
        RECT 40.370 178.755 40.540 178.875 ;
        RECT 39.410 178.585 40.540 178.755 ;
        RECT 41.120 178.705 41.290 179.215 ;
        RECT 38.765 177.705 38.935 177.955 ;
        RECT 39.410 177.885 39.580 178.585 ;
        RECT 40.720 178.535 41.290 178.705 ;
        RECT 41.460 179.215 43.410 179.385 ;
        RECT 39.930 178.245 40.550 178.415 ;
        RECT 39.930 178.065 40.140 178.245 ;
        RECT 40.720 178.055 40.890 178.535 ;
        RECT 41.460 178.225 41.630 179.215 ;
        RECT 42.220 178.625 42.405 178.935 ;
        RECT 42.675 178.625 42.870 178.935 ;
        RECT 39.410 177.555 39.670 177.885 ;
        RECT 39.980 177.385 40.310 177.765 ;
        RECT 40.490 177.725 40.890 178.055 ;
        RECT 41.080 177.895 41.630 178.225 ;
        RECT 41.800 177.725 41.970 178.625 ;
        RECT 40.490 177.555 41.970 177.725 ;
        RECT 42.220 178.295 42.450 178.625 ;
        RECT 42.675 178.295 42.930 178.625 ;
        RECT 43.240 178.295 43.410 179.215 ;
        RECT 42.220 177.715 42.405 178.295 ;
        RECT 42.675 177.720 42.870 178.295 ;
        RECT 43.080 177.385 43.410 177.765 ;
        RECT 43.580 177.555 43.840 179.765 ;
        RECT 44.010 178.845 45.680 179.935 ;
        RECT 44.010 178.325 44.760 178.845 ;
        RECT 45.910 178.795 46.120 179.935 ;
        RECT 46.290 178.785 46.620 179.765 ;
        RECT 46.790 178.795 47.020 179.935 ;
        RECT 44.930 178.155 45.680 178.675 ;
        RECT 44.010 177.385 45.680 178.155 ;
        RECT 45.910 177.385 46.120 178.205 ;
        RECT 46.290 178.185 46.540 178.785 ;
        RECT 47.235 178.745 47.490 179.625 ;
        RECT 47.660 178.795 47.965 179.935 ;
        RECT 48.305 179.555 48.635 179.935 ;
        RECT 48.815 179.385 48.985 179.675 ;
        RECT 49.155 179.475 49.405 179.935 ;
        RECT 48.185 179.215 48.985 179.385 ;
        RECT 49.575 179.425 50.445 179.765 ;
        RECT 46.710 178.375 47.040 178.625 ;
        RECT 46.290 177.555 46.620 178.185 ;
        RECT 46.790 177.385 47.020 178.205 ;
        RECT 47.235 178.095 47.445 178.745 ;
        RECT 48.185 178.625 48.355 179.215 ;
        RECT 49.575 179.045 49.745 179.425 ;
        RECT 50.680 179.305 50.850 179.765 ;
        RECT 51.020 179.475 51.390 179.935 ;
        RECT 51.685 179.335 51.855 179.675 ;
        RECT 52.025 179.505 52.355 179.935 ;
        RECT 52.590 179.335 52.760 179.675 ;
        RECT 48.525 178.875 49.745 179.045 ;
        RECT 49.915 178.965 50.375 179.255 ;
        RECT 50.680 179.135 51.240 179.305 ;
        RECT 51.685 179.165 52.760 179.335 ;
        RECT 52.930 179.435 53.610 179.765 ;
        RECT 53.825 179.435 54.075 179.765 ;
        RECT 54.245 179.475 54.495 179.935 ;
        RECT 51.070 178.995 51.240 179.135 ;
        RECT 49.915 178.955 50.880 178.965 ;
        RECT 49.575 178.785 49.745 178.875 ;
        RECT 50.205 178.795 50.880 178.955 ;
        RECT 47.615 178.595 48.355 178.625 ;
        RECT 47.615 178.295 48.530 178.595 ;
        RECT 48.205 178.120 48.530 178.295 ;
        RECT 47.235 177.565 47.490 178.095 ;
        RECT 47.660 177.385 47.965 177.845 ;
        RECT 48.210 177.765 48.530 178.120 ;
        RECT 48.700 178.335 49.240 178.705 ;
        RECT 49.575 178.615 49.980 178.785 ;
        RECT 48.700 177.935 48.940 178.335 ;
        RECT 49.420 178.165 49.640 178.445 ;
        RECT 49.110 177.995 49.640 178.165 ;
        RECT 49.110 177.765 49.280 177.995 ;
        RECT 49.810 177.835 49.980 178.615 ;
        RECT 50.150 178.005 50.500 178.625 ;
        RECT 50.670 178.005 50.880 178.795 ;
        RECT 51.070 178.825 52.570 178.995 ;
        RECT 51.070 178.135 51.240 178.825 ;
        RECT 52.930 178.655 53.100 179.435 ;
        RECT 53.905 179.305 54.075 179.435 ;
        RECT 51.410 178.485 53.100 178.655 ;
        RECT 53.270 178.875 53.735 179.265 ;
        RECT 53.905 179.135 54.300 179.305 ;
        RECT 51.410 178.305 51.580 178.485 ;
        RECT 48.210 177.595 49.280 177.765 ;
        RECT 49.450 177.385 49.640 177.825 ;
        RECT 49.810 177.555 50.760 177.835 ;
        RECT 51.070 177.745 51.330 178.135 ;
        RECT 51.750 178.065 52.540 178.315 ;
        RECT 50.980 177.575 51.330 177.745 ;
        RECT 51.540 177.385 51.870 177.845 ;
        RECT 52.745 177.775 52.915 178.485 ;
        RECT 53.270 178.285 53.440 178.875 ;
        RECT 53.085 178.065 53.440 178.285 ;
        RECT 53.610 178.065 53.960 178.685 ;
        RECT 54.130 177.775 54.300 179.135 ;
        RECT 54.665 178.965 54.990 179.750 ;
        RECT 54.470 177.915 54.930 178.965 ;
        RECT 52.745 177.605 53.600 177.775 ;
        RECT 53.805 177.605 54.300 177.775 ;
        RECT 54.470 177.385 54.800 177.745 ;
        RECT 55.160 177.645 55.330 179.765 ;
        RECT 55.500 179.435 55.830 179.935 ;
        RECT 56.000 179.265 56.255 179.765 ;
        RECT 55.505 179.095 56.255 179.265 ;
        RECT 55.505 178.105 55.735 179.095 ;
        RECT 56.635 178.965 56.965 179.765 ;
        RECT 57.135 179.135 57.465 179.935 ;
        RECT 57.765 178.965 58.095 179.765 ;
        RECT 58.740 179.135 58.990 179.935 ;
        RECT 55.905 178.275 56.255 178.925 ;
        RECT 56.635 178.795 59.070 178.965 ;
        RECT 59.260 178.795 59.430 179.935 ;
        RECT 59.600 178.795 59.940 179.765 ;
        RECT 56.430 178.375 56.780 178.625 ;
        RECT 56.965 178.165 57.135 178.795 ;
        RECT 57.305 178.375 57.635 178.575 ;
        RECT 57.805 178.375 58.135 178.575 ;
        RECT 58.305 178.375 58.725 178.575 ;
        RECT 58.900 178.545 59.070 178.795 ;
        RECT 58.900 178.375 59.595 178.545 ;
        RECT 55.505 177.935 56.255 178.105 ;
        RECT 55.500 177.385 55.830 177.765 ;
        RECT 56.000 177.645 56.255 177.935 ;
        RECT 56.635 177.555 57.135 178.165 ;
        RECT 57.765 178.035 58.990 178.205 ;
        RECT 59.765 178.185 59.940 178.795 ;
        RECT 60.570 178.770 60.860 179.935 ;
        RECT 61.070 178.795 61.300 179.935 ;
        RECT 61.470 178.785 61.800 179.765 ;
        RECT 61.970 178.795 62.180 179.935 ;
        RECT 62.410 179.175 62.925 179.585 ;
        RECT 63.160 179.175 63.330 179.935 ;
        RECT 63.500 179.595 65.530 179.765 ;
        RECT 61.050 178.375 61.380 178.625 ;
        RECT 57.765 177.555 58.095 178.035 ;
        RECT 58.265 177.385 58.490 177.845 ;
        RECT 58.660 177.555 58.990 178.035 ;
        RECT 59.180 177.385 59.430 178.185 ;
        RECT 59.600 177.555 59.940 178.185 ;
        RECT 60.570 177.385 60.860 178.110 ;
        RECT 61.070 177.385 61.300 178.205 ;
        RECT 61.550 178.185 61.800 178.785 ;
        RECT 62.410 178.365 62.750 179.175 ;
        RECT 63.500 178.930 63.670 179.595 ;
        RECT 64.065 179.255 65.190 179.425 ;
        RECT 62.920 178.740 63.670 178.930 ;
        RECT 63.840 178.915 64.850 179.085 ;
        RECT 61.470 177.555 61.800 178.185 ;
        RECT 61.970 177.385 62.180 178.205 ;
        RECT 62.410 178.195 63.640 178.365 ;
        RECT 62.685 177.590 62.930 178.195 ;
        RECT 63.150 177.385 63.660 177.920 ;
        RECT 63.840 177.555 64.030 178.915 ;
        RECT 64.200 178.575 64.475 178.715 ;
        RECT 64.200 178.405 64.480 178.575 ;
        RECT 64.200 177.555 64.475 178.405 ;
        RECT 64.680 178.115 64.850 178.915 ;
        RECT 65.020 178.125 65.190 179.255 ;
        RECT 65.360 178.625 65.530 179.595 ;
        RECT 65.700 178.795 65.870 179.935 ;
        RECT 66.040 178.795 66.375 179.765 ;
        RECT 66.665 179.305 66.950 179.765 ;
        RECT 67.120 179.475 67.390 179.935 ;
        RECT 66.665 179.085 67.620 179.305 ;
        RECT 65.360 178.295 65.555 178.625 ;
        RECT 65.780 178.295 66.035 178.625 ;
        RECT 65.780 178.125 65.950 178.295 ;
        RECT 66.205 178.125 66.375 178.795 ;
        RECT 66.550 178.355 67.240 178.915 ;
        RECT 67.410 178.185 67.620 179.085 ;
        RECT 65.020 177.955 65.950 178.125 ;
        RECT 65.020 177.920 65.195 177.955 ;
        RECT 64.665 177.555 65.195 177.920 ;
        RECT 65.620 177.385 65.950 177.785 ;
        RECT 66.120 177.555 66.375 178.125 ;
        RECT 66.665 178.015 67.620 178.185 ;
        RECT 67.790 178.915 68.190 179.765 ;
        RECT 68.380 179.305 68.660 179.765 ;
        RECT 69.180 179.475 69.505 179.935 ;
        RECT 68.380 179.085 69.505 179.305 ;
        RECT 67.790 178.355 68.885 178.915 ;
        RECT 69.055 178.625 69.505 179.085 ;
        RECT 69.675 178.795 70.060 179.765 ;
        RECT 66.665 177.555 66.950 178.015 ;
        RECT 67.120 177.385 67.390 177.845 ;
        RECT 67.790 177.555 68.190 178.355 ;
        RECT 69.055 178.295 69.610 178.625 ;
        RECT 69.055 178.185 69.505 178.295 ;
        RECT 68.380 178.015 69.505 178.185 ;
        RECT 69.780 178.125 70.060 178.795 ;
        RECT 68.380 177.555 68.660 178.015 ;
        RECT 69.180 177.385 69.505 177.845 ;
        RECT 69.675 177.555 70.060 178.125 ;
        RECT 70.230 178.795 70.570 179.765 ;
        RECT 70.740 178.795 70.910 179.935 ;
        RECT 71.180 179.135 71.430 179.935 ;
        RECT 72.075 178.965 72.405 179.765 ;
        RECT 72.705 179.135 73.035 179.935 ;
        RECT 73.205 178.965 73.535 179.765 ;
        RECT 73.915 179.265 74.170 179.765 ;
        RECT 74.340 179.435 74.670 179.935 ;
        RECT 73.915 179.095 74.665 179.265 ;
        RECT 71.100 178.795 73.535 178.965 ;
        RECT 70.230 178.745 70.460 178.795 ;
        RECT 70.230 178.185 70.405 178.745 ;
        RECT 71.100 178.545 71.270 178.795 ;
        RECT 70.575 178.375 71.270 178.545 ;
        RECT 71.445 178.375 71.865 178.575 ;
        RECT 72.035 178.375 72.365 178.575 ;
        RECT 72.535 178.375 72.865 178.575 ;
        RECT 70.230 177.555 70.570 178.185 ;
        RECT 70.740 177.385 70.990 178.185 ;
        RECT 71.180 178.035 72.405 178.205 ;
        RECT 71.180 177.555 71.510 178.035 ;
        RECT 71.680 177.385 71.905 177.845 ;
        RECT 72.075 177.555 72.405 178.035 ;
        RECT 73.035 178.165 73.205 178.795 ;
        RECT 73.390 178.375 73.740 178.625 ;
        RECT 73.915 178.275 74.265 178.925 ;
        RECT 73.035 177.555 73.535 178.165 ;
        RECT 74.435 178.105 74.665 179.095 ;
        RECT 73.915 177.935 74.665 178.105 ;
        RECT 73.915 177.645 74.170 177.935 ;
        RECT 74.340 177.385 74.670 177.765 ;
        RECT 74.840 177.645 75.010 179.765 ;
        RECT 75.180 178.965 75.505 179.750 ;
        RECT 75.675 179.475 75.925 179.935 ;
        RECT 76.095 179.435 76.345 179.765 ;
        RECT 76.560 179.435 77.240 179.765 ;
        RECT 76.095 179.305 76.265 179.435 ;
        RECT 75.870 179.135 76.265 179.305 ;
        RECT 75.240 177.915 75.700 178.965 ;
        RECT 75.870 177.775 76.040 179.135 ;
        RECT 76.435 178.875 76.900 179.265 ;
        RECT 76.210 178.065 76.560 178.685 ;
        RECT 76.730 178.285 76.900 178.875 ;
        RECT 77.070 178.655 77.240 179.435 ;
        RECT 77.410 179.335 77.580 179.675 ;
        RECT 77.815 179.505 78.145 179.935 ;
        RECT 78.315 179.335 78.485 179.675 ;
        RECT 78.780 179.475 79.150 179.935 ;
        RECT 77.410 179.165 78.485 179.335 ;
        RECT 79.320 179.305 79.490 179.765 ;
        RECT 79.725 179.425 80.595 179.765 ;
        RECT 80.765 179.475 81.015 179.935 ;
        RECT 78.930 179.135 79.490 179.305 ;
        RECT 78.930 178.995 79.100 179.135 ;
        RECT 77.600 178.825 79.100 178.995 ;
        RECT 79.795 178.965 80.255 179.255 ;
        RECT 77.070 178.485 78.760 178.655 ;
        RECT 76.730 178.065 77.085 178.285 ;
        RECT 77.255 177.775 77.425 178.485 ;
        RECT 77.630 178.065 78.420 178.315 ;
        RECT 78.590 178.305 78.760 178.485 ;
        RECT 78.930 178.135 79.100 178.825 ;
        RECT 75.370 177.385 75.700 177.745 ;
        RECT 75.870 177.605 76.365 177.775 ;
        RECT 76.570 177.605 77.425 177.775 ;
        RECT 78.300 177.385 78.630 177.845 ;
        RECT 78.840 177.745 79.100 178.135 ;
        RECT 79.290 178.955 80.255 178.965 ;
        RECT 80.425 179.045 80.595 179.425 ;
        RECT 81.185 179.385 81.355 179.675 ;
        RECT 81.535 179.555 81.865 179.935 ;
        RECT 81.185 179.215 81.985 179.385 ;
        RECT 79.290 178.795 79.965 178.955 ;
        RECT 80.425 178.875 81.645 179.045 ;
        RECT 79.290 178.005 79.500 178.795 ;
        RECT 80.425 178.785 80.595 178.875 ;
        RECT 79.670 178.005 80.020 178.625 ;
        RECT 80.190 178.615 80.595 178.785 ;
        RECT 80.190 177.835 80.360 178.615 ;
        RECT 80.530 178.165 80.750 178.445 ;
        RECT 80.930 178.335 81.470 178.705 ;
        RECT 81.815 178.625 81.985 179.215 ;
        RECT 82.205 178.795 82.510 179.935 ;
        RECT 82.680 178.745 82.935 179.625 ;
        RECT 81.815 178.595 82.555 178.625 ;
        RECT 80.530 177.995 81.060 178.165 ;
        RECT 78.840 177.575 79.190 177.745 ;
        RECT 79.410 177.555 80.360 177.835 ;
        RECT 80.530 177.385 80.720 177.825 ;
        RECT 80.890 177.765 81.060 177.995 ;
        RECT 81.230 177.935 81.470 178.335 ;
        RECT 81.640 178.295 82.555 178.595 ;
        RECT 81.640 178.120 81.965 178.295 ;
        RECT 81.640 177.765 81.960 178.120 ;
        RECT 82.725 178.095 82.935 178.745 ;
        RECT 80.890 177.595 81.960 177.765 ;
        RECT 82.205 177.385 82.510 177.845 ;
        RECT 82.680 177.565 82.935 178.095 ;
        RECT 83.110 178.795 83.380 179.765 ;
        RECT 83.590 179.135 83.870 179.935 ;
        RECT 84.040 179.425 85.695 179.715 ;
        RECT 84.105 179.085 85.695 179.255 ;
        RECT 84.105 178.965 84.275 179.085 ;
        RECT 83.550 178.795 84.275 178.965 ;
        RECT 83.110 178.060 83.280 178.795 ;
        RECT 83.550 178.625 83.720 178.795 ;
        RECT 83.450 178.295 83.720 178.625 ;
        RECT 83.890 178.295 84.295 178.625 ;
        RECT 84.465 178.295 85.175 178.915 ;
        RECT 85.375 178.795 85.695 179.085 ;
        RECT 86.330 178.770 86.620 179.935 ;
        RECT 86.790 178.845 88.460 179.935 ;
        RECT 83.550 178.125 83.720 178.295 ;
        RECT 83.110 177.715 83.380 178.060 ;
        RECT 83.550 177.955 85.160 178.125 ;
        RECT 85.345 178.055 85.695 178.625 ;
        RECT 86.790 178.325 87.540 178.845 ;
        RECT 88.630 178.795 88.970 179.765 ;
        RECT 89.140 178.795 89.310 179.935 ;
        RECT 89.580 179.135 89.830 179.935 ;
        RECT 90.475 178.965 90.805 179.765 ;
        RECT 91.105 179.135 91.435 179.935 ;
        RECT 91.605 178.965 91.935 179.765 ;
        RECT 89.500 178.795 91.935 178.965 ;
        RECT 92.310 179.175 92.825 179.585 ;
        RECT 93.060 179.175 93.230 179.935 ;
        RECT 93.400 179.595 95.430 179.765 ;
        RECT 87.710 178.155 88.460 178.675 ;
        RECT 83.570 177.385 83.950 177.785 ;
        RECT 84.120 177.605 84.290 177.955 ;
        RECT 84.460 177.385 84.790 177.785 ;
        RECT 84.990 177.605 85.160 177.955 ;
        RECT 85.360 177.385 85.690 177.885 ;
        RECT 86.330 177.385 86.620 178.110 ;
        RECT 86.790 177.385 88.460 178.155 ;
        RECT 88.630 178.235 88.805 178.795 ;
        RECT 89.500 178.545 89.670 178.795 ;
        RECT 88.975 178.375 89.670 178.545 ;
        RECT 89.845 178.375 90.265 178.575 ;
        RECT 90.435 178.375 90.765 178.575 ;
        RECT 90.935 178.375 91.265 178.575 ;
        RECT 88.630 178.185 88.860 178.235 ;
        RECT 88.630 177.555 88.970 178.185 ;
        RECT 89.140 177.385 89.390 178.185 ;
        RECT 89.580 178.035 90.805 178.205 ;
        RECT 89.580 177.555 89.910 178.035 ;
        RECT 90.080 177.385 90.305 177.845 ;
        RECT 90.475 177.555 90.805 178.035 ;
        RECT 91.435 178.165 91.605 178.795 ;
        RECT 91.790 178.375 92.140 178.625 ;
        RECT 92.310 178.365 92.650 179.175 ;
        RECT 93.400 178.930 93.570 179.595 ;
        RECT 93.965 179.255 95.090 179.425 ;
        RECT 92.820 178.740 93.570 178.930 ;
        RECT 93.740 178.915 94.750 179.085 ;
        RECT 92.310 178.195 93.540 178.365 ;
        RECT 91.435 177.555 91.935 178.165 ;
        RECT 92.585 177.590 92.830 178.195 ;
        RECT 93.050 177.385 93.560 177.920 ;
        RECT 93.740 177.555 93.930 178.915 ;
        RECT 94.100 178.575 94.375 178.715 ;
        RECT 94.100 178.405 94.380 178.575 ;
        RECT 94.100 177.555 94.375 178.405 ;
        RECT 94.580 178.115 94.750 178.915 ;
        RECT 94.920 178.125 95.090 179.255 ;
        RECT 95.260 178.625 95.430 179.595 ;
        RECT 95.600 178.795 95.770 179.935 ;
        RECT 95.940 178.795 96.275 179.765 ;
        RECT 96.510 178.795 96.720 179.935 ;
        RECT 95.260 178.295 95.455 178.625 ;
        RECT 95.680 178.295 95.935 178.625 ;
        RECT 95.680 178.125 95.850 178.295 ;
        RECT 96.105 178.125 96.275 178.795 ;
        RECT 96.890 178.785 97.220 179.765 ;
        RECT 97.390 178.795 97.620 179.935 ;
        RECT 98.290 178.845 100.880 179.935 ;
        RECT 94.920 177.955 95.850 178.125 ;
        RECT 94.920 177.920 95.095 177.955 ;
        RECT 94.565 177.555 95.095 177.920 ;
        RECT 95.520 177.385 95.850 177.785 ;
        RECT 96.020 177.555 96.275 178.125 ;
        RECT 96.510 177.385 96.720 178.205 ;
        RECT 96.890 178.185 97.140 178.785 ;
        RECT 97.310 178.375 97.640 178.625 ;
        RECT 98.290 178.325 99.500 178.845 ;
        RECT 101.090 178.795 101.320 179.935 ;
        RECT 101.490 178.785 101.820 179.765 ;
        RECT 101.990 178.795 102.200 179.935 ;
        RECT 102.890 178.845 105.480 179.935 ;
        RECT 105.655 179.500 111.000 179.935 ;
        RECT 96.890 177.555 97.220 178.185 ;
        RECT 97.390 177.385 97.620 178.205 ;
        RECT 99.670 178.155 100.880 178.675 ;
        RECT 101.070 178.375 101.400 178.625 ;
        RECT 98.290 177.385 100.880 178.155 ;
        RECT 101.090 177.385 101.320 178.205 ;
        RECT 101.570 178.185 101.820 178.785 ;
        RECT 102.890 178.325 104.100 178.845 ;
        RECT 101.490 177.555 101.820 178.185 ;
        RECT 101.990 177.385 102.200 178.205 ;
        RECT 104.270 178.155 105.480 178.675 ;
        RECT 107.245 178.250 107.595 179.500 ;
        RECT 111.170 178.845 112.380 179.935 ;
        RECT 102.890 177.385 105.480 178.155 ;
        RECT 109.075 177.930 109.415 178.760 ;
        RECT 111.170 178.305 111.690 178.845 ;
        RECT 111.860 178.135 112.380 178.675 ;
        RECT 105.655 177.385 111.000 177.930 ;
        RECT 111.170 177.385 112.380 178.135 ;
        RECT 18.165 177.215 112.465 177.385 ;
        RECT 18.250 176.465 19.460 177.215 ;
        RECT 18.250 175.925 18.770 176.465 ;
        RECT 20.610 176.395 20.820 177.215 ;
        RECT 20.990 176.415 21.320 177.045 ;
        RECT 18.940 175.755 19.460 176.295 ;
        RECT 20.990 175.815 21.240 176.415 ;
        RECT 21.490 176.395 21.720 177.215 ;
        RECT 21.930 176.490 22.220 177.215 ;
        RECT 22.395 176.505 22.650 177.035 ;
        RECT 22.820 176.755 23.125 177.215 ;
        RECT 23.370 176.835 24.440 177.005 ;
        RECT 21.410 175.975 21.740 176.225 ;
        RECT 22.395 175.855 22.605 176.505 ;
        RECT 23.370 176.480 23.690 176.835 ;
        RECT 23.365 176.305 23.690 176.480 ;
        RECT 22.775 176.005 23.690 176.305 ;
        RECT 23.860 176.265 24.100 176.665 ;
        RECT 24.270 176.605 24.440 176.835 ;
        RECT 24.610 176.775 24.800 177.215 ;
        RECT 24.970 176.765 25.920 177.045 ;
        RECT 26.140 176.855 26.490 177.025 ;
        RECT 24.270 176.435 24.800 176.605 ;
        RECT 22.775 175.975 23.515 176.005 ;
        RECT 18.250 174.665 19.460 175.755 ;
        RECT 20.610 174.665 20.820 175.805 ;
        RECT 20.990 174.835 21.320 175.815 ;
        RECT 21.490 174.665 21.720 175.805 ;
        RECT 21.930 174.665 22.220 175.830 ;
        RECT 22.395 174.975 22.650 175.855 ;
        RECT 22.820 174.665 23.125 175.805 ;
        RECT 23.345 175.385 23.515 175.975 ;
        RECT 23.860 175.895 24.400 176.265 ;
        RECT 24.580 176.155 24.800 176.435 ;
        RECT 24.970 175.985 25.140 176.765 ;
        RECT 24.735 175.815 25.140 175.985 ;
        RECT 25.310 175.975 25.660 176.595 ;
        RECT 24.735 175.725 24.905 175.815 ;
        RECT 25.830 175.805 26.040 176.595 ;
        RECT 23.685 175.555 24.905 175.725 ;
        RECT 25.365 175.645 26.040 175.805 ;
        RECT 23.345 175.215 24.145 175.385 ;
        RECT 23.465 174.665 23.795 175.045 ;
        RECT 23.975 174.925 24.145 175.215 ;
        RECT 24.735 175.175 24.905 175.555 ;
        RECT 25.075 175.635 26.040 175.645 ;
        RECT 26.230 176.465 26.490 176.855 ;
        RECT 26.700 176.755 27.030 177.215 ;
        RECT 27.905 176.825 28.760 176.995 ;
        RECT 28.965 176.825 29.460 176.995 ;
        RECT 29.630 176.855 29.960 177.215 ;
        RECT 26.230 175.775 26.400 176.465 ;
        RECT 26.570 176.115 26.740 176.295 ;
        RECT 26.910 176.285 27.700 176.535 ;
        RECT 27.905 176.115 28.075 176.825 ;
        RECT 28.245 176.315 28.600 176.535 ;
        RECT 26.570 175.945 28.260 176.115 ;
        RECT 25.075 175.345 25.535 175.635 ;
        RECT 26.230 175.605 27.730 175.775 ;
        RECT 26.230 175.465 26.400 175.605 ;
        RECT 25.840 175.295 26.400 175.465 ;
        RECT 24.315 174.665 24.565 175.125 ;
        RECT 24.735 174.835 25.605 175.175 ;
        RECT 25.840 174.835 26.010 175.295 ;
        RECT 26.845 175.265 27.920 175.435 ;
        RECT 26.180 174.665 26.550 175.125 ;
        RECT 26.845 174.925 27.015 175.265 ;
        RECT 27.185 174.665 27.515 175.095 ;
        RECT 27.750 174.925 27.920 175.265 ;
        RECT 28.090 175.165 28.260 175.945 ;
        RECT 28.430 175.725 28.600 176.315 ;
        RECT 28.770 175.915 29.120 176.535 ;
        RECT 28.430 175.335 28.895 175.725 ;
        RECT 29.290 175.465 29.460 176.825 ;
        RECT 29.630 175.635 30.090 176.685 ;
        RECT 29.065 175.295 29.460 175.465 ;
        RECT 29.065 175.165 29.235 175.295 ;
        RECT 28.090 174.835 28.770 175.165 ;
        RECT 28.985 174.835 29.235 175.165 ;
        RECT 29.405 174.665 29.655 175.125 ;
        RECT 29.825 174.850 30.150 175.635 ;
        RECT 30.320 174.835 30.490 176.955 ;
        RECT 30.660 176.835 30.990 177.215 ;
        RECT 31.160 176.665 31.415 176.955 ;
        RECT 30.665 176.495 31.415 176.665 ;
        RECT 30.665 175.505 30.895 176.495 ;
        RECT 31.650 176.395 31.860 177.215 ;
        RECT 32.030 176.415 32.360 177.045 ;
        RECT 31.065 175.675 31.415 176.325 ;
        RECT 32.030 175.815 32.280 176.415 ;
        RECT 32.530 176.395 32.760 177.215 ;
        RECT 33.240 176.820 33.570 177.215 ;
        RECT 33.740 176.645 33.940 177.000 ;
        RECT 34.110 176.815 34.440 177.215 ;
        RECT 34.610 176.645 34.810 176.990 ;
        RECT 32.970 176.475 34.810 176.645 ;
        RECT 34.980 176.475 35.310 177.215 ;
        RECT 35.545 176.645 35.715 176.895 ;
        RECT 36.275 176.645 36.450 177.045 ;
        RECT 36.620 176.835 36.950 177.215 ;
        RECT 37.195 176.715 37.425 177.045 ;
        RECT 35.545 176.475 36.020 176.645 ;
        RECT 36.275 176.475 36.905 176.645 ;
        RECT 32.450 175.975 32.780 176.225 ;
        RECT 30.665 175.335 31.415 175.505 ;
        RECT 30.660 174.665 30.990 175.165 ;
        RECT 31.160 174.835 31.415 175.335 ;
        RECT 31.650 174.665 31.860 175.805 ;
        RECT 32.030 174.835 32.360 175.815 ;
        RECT 32.530 174.665 32.760 175.805 ;
        RECT 32.970 174.850 33.230 176.475 ;
        RECT 33.410 175.505 33.630 176.305 ;
        RECT 33.870 175.685 34.170 176.305 ;
        RECT 34.340 175.685 34.670 176.305 ;
        RECT 34.840 175.685 35.160 176.305 ;
        RECT 35.330 175.685 35.680 176.305 ;
        RECT 35.850 175.505 36.020 176.475 ;
        RECT 36.735 176.305 36.905 176.475 ;
        RECT 36.190 175.625 36.555 176.305 ;
        RECT 36.735 175.975 37.085 176.305 ;
        RECT 33.410 175.295 36.020 175.505 ;
        RECT 36.735 175.455 36.905 175.975 ;
        RECT 36.275 175.285 36.905 175.455 ;
        RECT 37.255 175.425 37.425 176.715 ;
        RECT 37.625 175.605 37.905 176.880 ;
        RECT 38.130 175.855 38.400 176.880 ;
        RECT 38.860 176.835 39.190 177.215 ;
        RECT 39.360 176.960 39.695 177.005 ;
        RECT 38.090 175.685 38.400 175.855 ;
        RECT 38.130 175.605 38.400 175.685 ;
        RECT 38.590 175.605 38.930 176.635 ;
        RECT 39.360 176.495 39.700 176.960 ;
        RECT 39.100 175.975 39.360 176.305 ;
        RECT 39.100 175.425 39.270 175.975 ;
        RECT 39.530 175.805 39.700 176.495 ;
        RECT 40.445 176.585 40.730 177.045 ;
        RECT 40.900 176.755 41.170 177.215 ;
        RECT 40.445 176.415 41.400 176.585 ;
        RECT 34.980 174.665 35.310 175.115 ;
        RECT 36.275 174.835 36.450 175.285 ;
        RECT 37.255 175.255 39.270 175.425 ;
        RECT 36.620 174.665 36.950 175.105 ;
        RECT 37.255 174.835 37.425 175.255 ;
        RECT 37.660 174.665 38.330 175.075 ;
        RECT 38.545 174.835 38.715 175.255 ;
        RECT 38.915 174.665 39.245 175.075 ;
        RECT 39.440 174.835 39.700 175.805 ;
        RECT 40.330 175.685 41.020 176.245 ;
        RECT 41.190 175.515 41.400 176.415 ;
        RECT 40.445 175.295 41.400 175.515 ;
        RECT 41.570 176.245 41.970 177.045 ;
        RECT 42.160 176.585 42.440 177.045 ;
        RECT 42.960 176.755 43.285 177.215 ;
        RECT 42.160 176.415 43.285 176.585 ;
        RECT 43.455 176.475 43.840 177.045 ;
        RECT 42.835 176.305 43.285 176.415 ;
        RECT 41.570 175.685 42.665 176.245 ;
        RECT 42.835 175.975 43.390 176.305 ;
        RECT 40.445 174.835 40.730 175.295 ;
        RECT 40.900 174.665 41.170 175.125 ;
        RECT 41.570 174.835 41.970 175.685 ;
        RECT 42.835 175.515 43.285 175.975 ;
        RECT 43.560 175.805 43.840 176.475 ;
        RECT 44.215 176.435 44.715 177.045 ;
        RECT 44.010 175.975 44.360 176.225 ;
        RECT 44.545 175.805 44.715 176.435 ;
        RECT 45.345 176.565 45.675 177.045 ;
        RECT 45.845 176.755 46.070 177.215 ;
        RECT 46.240 176.565 46.570 177.045 ;
        RECT 45.345 176.395 46.570 176.565 ;
        RECT 46.760 176.415 47.010 177.215 ;
        RECT 47.180 176.415 47.520 177.045 ;
        RECT 47.690 176.490 47.980 177.215 ;
        RECT 44.885 176.025 45.215 176.225 ;
        RECT 45.385 176.025 45.715 176.225 ;
        RECT 45.885 176.025 46.305 176.225 ;
        RECT 46.480 176.055 47.175 176.225 ;
        RECT 46.480 175.805 46.650 176.055 ;
        RECT 47.345 175.805 47.520 176.415 ;
        RECT 48.210 176.395 48.420 177.215 ;
        RECT 48.590 176.415 48.920 177.045 ;
        RECT 42.160 175.295 43.285 175.515 ;
        RECT 42.160 174.835 42.440 175.295 ;
        RECT 42.960 174.665 43.285 175.125 ;
        RECT 43.455 174.835 43.840 175.805 ;
        RECT 44.215 175.635 46.650 175.805 ;
        RECT 44.215 174.835 44.545 175.635 ;
        RECT 44.715 174.665 45.045 175.465 ;
        RECT 45.345 174.835 45.675 175.635 ;
        RECT 46.320 174.665 46.570 175.465 ;
        RECT 46.840 174.665 47.010 175.805 ;
        RECT 47.180 174.835 47.520 175.805 ;
        RECT 47.690 174.665 47.980 175.830 ;
        RECT 48.590 175.815 48.840 176.415 ;
        RECT 49.090 176.395 49.320 177.215 ;
        RECT 49.530 176.465 50.740 177.215 ;
        RECT 49.010 175.975 49.340 176.225 ;
        RECT 48.210 174.665 48.420 175.805 ;
        RECT 48.590 174.835 48.920 175.815 ;
        RECT 49.090 174.665 49.320 175.805 ;
        RECT 49.530 175.755 50.050 176.295 ;
        RECT 50.220 175.925 50.740 176.465 ;
        RECT 51.025 176.585 51.310 177.045 ;
        RECT 51.480 176.755 51.750 177.215 ;
        RECT 51.025 176.415 51.980 176.585 ;
        RECT 49.530 174.665 50.740 175.755 ;
        RECT 50.910 175.685 51.600 176.245 ;
        RECT 51.770 175.515 51.980 176.415 ;
        RECT 51.025 175.295 51.980 175.515 ;
        RECT 52.150 176.245 52.550 177.045 ;
        RECT 52.740 176.585 53.020 177.045 ;
        RECT 53.540 176.755 53.865 177.215 ;
        RECT 52.740 176.415 53.865 176.585 ;
        RECT 54.035 176.475 54.420 177.045 ;
        RECT 53.415 176.305 53.865 176.415 ;
        RECT 52.150 175.685 53.245 176.245 ;
        RECT 53.415 175.975 53.970 176.305 ;
        RECT 51.025 174.835 51.310 175.295 ;
        RECT 51.480 174.665 51.750 175.125 ;
        RECT 52.150 174.835 52.550 175.685 ;
        RECT 53.415 175.515 53.865 175.975 ;
        RECT 54.140 175.805 54.420 176.475 ;
        RECT 52.740 175.295 53.865 175.515 ;
        RECT 52.740 174.835 53.020 175.295 ;
        RECT 53.540 174.665 53.865 175.125 ;
        RECT 54.035 174.835 54.420 175.805 ;
        RECT 54.590 176.415 54.930 177.045 ;
        RECT 55.100 176.415 55.350 177.215 ;
        RECT 55.540 176.565 55.870 177.045 ;
        RECT 56.040 176.755 56.265 177.215 ;
        RECT 56.435 176.565 56.765 177.045 ;
        RECT 54.590 175.805 54.765 176.415 ;
        RECT 55.540 176.395 56.765 176.565 ;
        RECT 57.395 176.435 57.895 177.045 ;
        RECT 59.190 176.715 59.450 177.045 ;
        RECT 59.660 176.735 59.935 177.215 ;
        RECT 54.935 176.055 55.630 176.225 ;
        RECT 55.460 175.805 55.630 176.055 ;
        RECT 55.805 176.025 56.225 176.225 ;
        RECT 56.395 176.025 56.725 176.225 ;
        RECT 56.895 176.025 57.225 176.225 ;
        RECT 57.395 175.805 57.565 176.435 ;
        RECT 57.750 175.975 58.100 176.225 ;
        RECT 59.190 175.805 59.360 176.715 ;
        RECT 60.145 176.645 60.350 177.045 ;
        RECT 60.520 176.815 60.855 177.215 ;
        RECT 59.530 175.975 59.890 176.555 ;
        RECT 60.145 176.475 60.830 176.645 ;
        RECT 60.070 175.805 60.320 176.305 ;
        RECT 54.590 174.835 54.930 175.805 ;
        RECT 55.100 174.665 55.270 175.805 ;
        RECT 55.460 175.635 57.895 175.805 ;
        RECT 55.540 174.665 55.790 175.465 ;
        RECT 56.435 174.835 56.765 175.635 ;
        RECT 57.065 174.665 57.395 175.465 ;
        RECT 57.565 174.835 57.895 175.635 ;
        RECT 59.190 175.635 60.320 175.805 ;
        RECT 59.190 174.865 59.460 175.635 ;
        RECT 60.490 175.445 60.830 176.475 ;
        RECT 61.305 176.405 61.550 177.010 ;
        RECT 61.770 176.680 62.280 177.215 ;
        RECT 59.630 174.665 59.960 175.445 ;
        RECT 60.165 175.270 60.830 175.445 ;
        RECT 61.030 176.235 62.260 176.405 ;
        RECT 61.030 175.425 61.370 176.235 ;
        RECT 61.540 175.670 62.290 175.860 ;
        RECT 60.165 174.865 60.350 175.270 ;
        RECT 60.520 174.665 60.855 175.090 ;
        RECT 61.030 175.015 61.545 175.425 ;
        RECT 61.780 174.665 61.950 175.425 ;
        RECT 62.120 175.005 62.290 175.670 ;
        RECT 62.460 175.685 62.650 177.045 ;
        RECT 62.820 176.195 63.095 177.045 ;
        RECT 63.285 176.680 63.815 177.045 ;
        RECT 64.240 176.815 64.570 177.215 ;
        RECT 63.640 176.645 63.815 176.680 ;
        RECT 62.820 176.025 63.100 176.195 ;
        RECT 62.820 175.885 63.095 176.025 ;
        RECT 63.300 175.685 63.470 176.485 ;
        RECT 62.460 175.515 63.470 175.685 ;
        RECT 63.640 176.475 64.570 176.645 ;
        RECT 64.740 176.475 64.995 177.045 ;
        RECT 65.260 176.665 65.430 177.045 ;
        RECT 65.645 176.835 65.975 177.215 ;
        RECT 65.260 176.495 65.975 176.665 ;
        RECT 63.640 175.345 63.810 176.475 ;
        RECT 64.400 176.305 64.570 176.475 ;
        RECT 62.685 175.175 63.810 175.345 ;
        RECT 63.980 175.975 64.175 176.305 ;
        RECT 64.400 175.975 64.655 176.305 ;
        RECT 63.980 175.005 64.150 175.975 ;
        RECT 64.825 175.805 64.995 176.475 ;
        RECT 65.170 175.945 65.525 176.315 ;
        RECT 65.805 176.305 65.975 176.495 ;
        RECT 66.145 176.470 66.400 177.045 ;
        RECT 65.805 175.975 66.060 176.305 ;
        RECT 62.120 174.835 64.150 175.005 ;
        RECT 64.320 174.665 64.490 175.805 ;
        RECT 64.660 174.835 64.995 175.805 ;
        RECT 65.805 175.765 65.975 175.975 ;
        RECT 65.260 175.595 65.975 175.765 ;
        RECT 66.230 175.740 66.400 176.470 ;
        RECT 66.575 176.375 66.835 177.215 ;
        RECT 67.010 176.540 67.280 176.885 ;
        RECT 67.470 176.815 67.850 177.215 ;
        RECT 68.020 176.645 68.190 176.995 ;
        RECT 68.360 176.815 68.690 177.215 ;
        RECT 68.890 176.645 69.060 176.995 ;
        RECT 69.260 176.715 69.590 177.215 ;
        RECT 65.260 174.835 65.430 175.595 ;
        RECT 65.645 174.665 65.975 175.425 ;
        RECT 66.145 174.835 66.400 175.740 ;
        RECT 66.575 174.665 66.835 175.815 ;
        RECT 67.010 175.805 67.180 176.540 ;
        RECT 67.450 176.475 69.060 176.645 ;
        RECT 67.450 176.305 67.620 176.475 ;
        RECT 67.350 175.975 67.620 176.305 ;
        RECT 67.790 175.975 68.195 176.305 ;
        RECT 67.450 175.805 67.620 175.975 ;
        RECT 67.010 174.835 67.280 175.805 ;
        RECT 67.450 175.635 68.175 175.805 ;
        RECT 68.365 175.685 69.075 176.305 ;
        RECT 69.245 175.975 69.595 176.545 ;
        RECT 69.770 176.415 70.110 177.045 ;
        RECT 70.280 176.415 70.530 177.215 ;
        RECT 70.720 176.565 71.050 177.045 ;
        RECT 71.220 176.755 71.445 177.215 ;
        RECT 71.615 176.565 71.945 177.045 ;
        RECT 69.770 176.365 70.000 176.415 ;
        RECT 70.720 176.395 71.945 176.565 ;
        RECT 72.575 176.435 73.075 177.045 ;
        RECT 73.450 176.490 73.740 177.215 ;
        RECT 74.000 176.665 74.170 177.045 ;
        RECT 74.385 176.835 74.715 177.215 ;
        RECT 74.000 176.495 74.715 176.665 ;
        RECT 69.770 175.805 69.945 176.365 ;
        RECT 70.115 176.055 70.810 176.225 ;
        RECT 70.640 175.805 70.810 176.055 ;
        RECT 70.985 176.025 71.405 176.225 ;
        RECT 71.575 176.025 71.905 176.225 ;
        RECT 72.075 176.025 72.405 176.225 ;
        RECT 72.575 175.805 72.745 176.435 ;
        RECT 72.930 175.975 73.280 176.225 ;
        RECT 73.910 175.945 74.265 176.315 ;
        RECT 74.545 176.305 74.715 176.495 ;
        RECT 74.885 176.470 75.140 177.045 ;
        RECT 74.545 175.975 74.800 176.305 ;
        RECT 68.005 175.515 68.175 175.635 ;
        RECT 69.275 175.515 69.595 175.805 ;
        RECT 67.490 174.665 67.770 175.465 ;
        RECT 68.005 175.345 69.595 175.515 ;
        RECT 67.940 174.885 69.595 175.175 ;
        RECT 69.770 174.835 70.110 175.805 ;
        RECT 70.280 174.665 70.450 175.805 ;
        RECT 70.640 175.635 73.075 175.805 ;
        RECT 70.720 174.665 70.970 175.465 ;
        RECT 71.615 174.835 71.945 175.635 ;
        RECT 72.245 174.665 72.575 175.465 ;
        RECT 72.745 174.835 73.075 175.635 ;
        RECT 73.450 174.665 73.740 175.830 ;
        RECT 74.545 175.765 74.715 175.975 ;
        RECT 74.000 175.595 74.715 175.765 ;
        RECT 74.970 175.740 75.140 176.470 ;
        RECT 75.315 176.375 75.575 177.215 ;
        RECT 75.840 176.665 76.010 177.045 ;
        RECT 76.225 176.835 76.555 177.215 ;
        RECT 75.840 176.495 76.555 176.665 ;
        RECT 75.750 175.945 76.105 176.315 ;
        RECT 76.385 176.305 76.555 176.495 ;
        RECT 76.725 176.470 76.980 177.045 ;
        RECT 76.385 175.975 76.640 176.305 ;
        RECT 74.000 174.835 74.170 175.595 ;
        RECT 74.385 174.665 74.715 175.425 ;
        RECT 74.885 174.835 75.140 175.740 ;
        RECT 75.315 174.665 75.575 175.815 ;
        RECT 76.385 175.765 76.555 175.975 ;
        RECT 75.840 175.595 76.555 175.765 ;
        RECT 76.810 175.740 76.980 176.470 ;
        RECT 77.155 176.375 77.415 177.215 ;
        RECT 78.255 176.435 78.755 177.045 ;
        RECT 78.050 175.975 78.400 176.225 ;
        RECT 75.840 174.835 76.010 175.595 ;
        RECT 76.225 174.665 76.555 175.425 ;
        RECT 76.725 174.835 76.980 175.740 ;
        RECT 77.155 174.665 77.415 175.815 ;
        RECT 78.585 175.805 78.755 176.435 ;
        RECT 79.385 176.565 79.715 177.045 ;
        RECT 79.885 176.755 80.110 177.215 ;
        RECT 80.280 176.565 80.610 177.045 ;
        RECT 79.385 176.395 80.610 176.565 ;
        RECT 80.800 176.415 81.050 177.215 ;
        RECT 81.220 176.415 81.560 177.045 ;
        RECT 81.935 176.435 82.435 177.045 ;
        RECT 78.925 176.025 79.255 176.225 ;
        RECT 79.425 176.025 79.755 176.225 ;
        RECT 79.925 176.025 80.345 176.225 ;
        RECT 80.520 176.055 81.215 176.225 ;
        RECT 80.520 175.805 80.690 176.055 ;
        RECT 81.385 175.805 81.560 176.415 ;
        RECT 81.730 175.975 82.080 176.225 ;
        RECT 82.265 175.805 82.435 176.435 ;
        RECT 83.065 176.565 83.395 177.045 ;
        RECT 83.565 176.755 83.790 177.215 ;
        RECT 83.960 176.565 84.290 177.045 ;
        RECT 83.065 176.395 84.290 176.565 ;
        RECT 84.480 176.415 84.730 177.215 ;
        RECT 84.900 176.415 85.240 177.045 ;
        RECT 85.525 176.585 85.810 177.045 ;
        RECT 85.980 176.755 86.250 177.215 ;
        RECT 85.525 176.415 86.480 176.585 ;
        RECT 82.605 176.025 82.935 176.225 ;
        RECT 83.105 176.025 83.435 176.225 ;
        RECT 83.605 176.025 84.025 176.225 ;
        RECT 84.200 176.055 84.895 176.225 ;
        RECT 84.200 175.805 84.370 176.055 ;
        RECT 85.065 175.805 85.240 176.415 ;
        RECT 78.255 175.635 80.690 175.805 ;
        RECT 78.255 174.835 78.585 175.635 ;
        RECT 78.755 174.665 79.085 175.465 ;
        RECT 79.385 174.835 79.715 175.635 ;
        RECT 80.360 174.665 80.610 175.465 ;
        RECT 80.880 174.665 81.050 175.805 ;
        RECT 81.220 174.835 81.560 175.805 ;
        RECT 81.935 175.635 84.370 175.805 ;
        RECT 81.935 174.835 82.265 175.635 ;
        RECT 82.435 174.665 82.765 175.465 ;
        RECT 83.065 174.835 83.395 175.635 ;
        RECT 84.040 174.665 84.290 175.465 ;
        RECT 84.560 174.665 84.730 175.805 ;
        RECT 84.900 174.835 85.240 175.805 ;
        RECT 85.410 175.685 86.100 176.245 ;
        RECT 86.270 175.515 86.480 176.415 ;
        RECT 85.525 175.295 86.480 175.515 ;
        RECT 86.650 176.245 87.050 177.045 ;
        RECT 87.240 176.585 87.520 177.045 ;
        RECT 88.040 176.755 88.365 177.215 ;
        RECT 87.240 176.415 88.365 176.585 ;
        RECT 88.535 176.475 88.920 177.045 ;
        RECT 87.915 176.305 88.365 176.415 ;
        RECT 86.650 175.685 87.745 176.245 ;
        RECT 87.915 175.975 88.470 176.305 ;
        RECT 85.525 174.835 85.810 175.295 ;
        RECT 85.980 174.665 86.250 175.125 ;
        RECT 86.650 174.835 87.050 175.685 ;
        RECT 87.915 175.515 88.365 175.975 ;
        RECT 88.640 175.805 88.920 176.475 ;
        RECT 87.240 175.295 88.365 175.515 ;
        RECT 87.240 174.835 87.520 175.295 ;
        RECT 88.040 174.665 88.365 175.125 ;
        RECT 88.535 174.835 88.920 175.805 ;
        RECT 90.015 176.505 90.270 177.035 ;
        RECT 90.440 176.755 90.745 177.215 ;
        RECT 90.990 176.835 92.060 177.005 ;
        RECT 90.015 175.855 90.225 176.505 ;
        RECT 90.990 176.480 91.310 176.835 ;
        RECT 90.985 176.305 91.310 176.480 ;
        RECT 90.395 176.005 91.310 176.305 ;
        RECT 91.480 176.265 91.720 176.665 ;
        RECT 91.890 176.605 92.060 176.835 ;
        RECT 92.230 176.775 92.420 177.215 ;
        RECT 92.590 176.765 93.540 177.045 ;
        RECT 93.760 176.855 94.110 177.025 ;
        RECT 91.890 176.435 92.420 176.605 ;
        RECT 90.395 175.975 91.135 176.005 ;
        RECT 90.015 174.975 90.270 175.855 ;
        RECT 90.440 174.665 90.745 175.805 ;
        RECT 90.965 175.385 91.135 175.975 ;
        RECT 91.480 175.895 92.020 176.265 ;
        RECT 92.200 176.155 92.420 176.435 ;
        RECT 92.590 175.985 92.760 176.765 ;
        RECT 92.355 175.815 92.760 175.985 ;
        RECT 92.930 175.975 93.280 176.595 ;
        RECT 92.355 175.725 92.525 175.815 ;
        RECT 93.450 175.805 93.660 176.595 ;
        RECT 91.305 175.555 92.525 175.725 ;
        RECT 92.985 175.645 93.660 175.805 ;
        RECT 90.965 175.215 91.765 175.385 ;
        RECT 91.085 174.665 91.415 175.045 ;
        RECT 91.595 174.925 91.765 175.215 ;
        RECT 92.355 175.175 92.525 175.555 ;
        RECT 92.695 175.635 93.660 175.645 ;
        RECT 93.850 176.465 94.110 176.855 ;
        RECT 94.320 176.755 94.650 177.215 ;
        RECT 95.525 176.825 96.380 176.995 ;
        RECT 96.585 176.825 97.080 176.995 ;
        RECT 97.250 176.855 97.580 177.215 ;
        RECT 93.850 175.775 94.020 176.465 ;
        RECT 94.190 176.115 94.360 176.295 ;
        RECT 94.530 176.285 95.320 176.535 ;
        RECT 95.525 176.115 95.695 176.825 ;
        RECT 95.865 176.315 96.220 176.535 ;
        RECT 94.190 175.945 95.880 176.115 ;
        RECT 92.695 175.345 93.155 175.635 ;
        RECT 93.850 175.605 95.350 175.775 ;
        RECT 93.850 175.465 94.020 175.605 ;
        RECT 93.460 175.295 94.020 175.465 ;
        RECT 91.935 174.665 92.185 175.125 ;
        RECT 92.355 174.835 93.225 175.175 ;
        RECT 93.460 174.835 93.630 175.295 ;
        RECT 94.465 175.265 95.540 175.435 ;
        RECT 93.800 174.665 94.170 175.125 ;
        RECT 94.465 174.925 94.635 175.265 ;
        RECT 94.805 174.665 95.135 175.095 ;
        RECT 95.370 174.925 95.540 175.265 ;
        RECT 95.710 175.165 95.880 175.945 ;
        RECT 96.050 175.725 96.220 176.315 ;
        RECT 96.390 175.915 96.740 176.535 ;
        RECT 96.050 175.335 96.515 175.725 ;
        RECT 96.910 175.465 97.080 176.825 ;
        RECT 97.250 175.635 97.710 176.685 ;
        RECT 96.685 175.295 97.080 175.465 ;
        RECT 96.685 175.165 96.855 175.295 ;
        RECT 95.710 174.835 96.390 175.165 ;
        RECT 96.605 174.835 96.855 175.165 ;
        RECT 97.025 174.665 97.275 175.125 ;
        RECT 97.445 174.850 97.770 175.635 ;
        RECT 97.940 174.835 98.110 176.955 ;
        RECT 98.280 176.835 98.610 177.215 ;
        RECT 98.780 176.665 99.035 176.955 ;
        RECT 98.285 176.495 99.035 176.665 ;
        RECT 98.285 175.505 98.515 176.495 ;
        RECT 99.210 176.490 99.500 177.215 ;
        RECT 100.045 176.505 100.300 177.035 ;
        RECT 100.480 176.755 100.765 177.215 ;
        RECT 98.685 175.675 99.035 176.325 ;
        RECT 98.285 175.335 99.035 175.505 ;
        RECT 98.280 174.665 98.610 175.165 ;
        RECT 98.780 174.835 99.035 175.335 ;
        RECT 99.210 174.665 99.500 175.830 ;
        RECT 100.045 175.645 100.225 176.505 ;
        RECT 100.945 176.305 101.195 176.955 ;
        RECT 100.395 175.975 101.195 176.305 ;
        RECT 100.045 175.175 100.300 175.645 ;
        RECT 99.960 175.005 100.300 175.175 ;
        RECT 100.045 174.975 100.300 175.005 ;
        RECT 100.480 174.665 100.765 175.465 ;
        RECT 100.945 175.385 101.195 175.975 ;
        RECT 101.395 176.620 101.715 176.950 ;
        RECT 101.895 176.735 102.555 177.215 ;
        RECT 102.755 176.825 103.605 176.995 ;
        RECT 101.395 175.725 101.585 176.620 ;
        RECT 101.905 176.295 102.565 176.565 ;
        RECT 102.235 176.235 102.565 176.295 ;
        RECT 101.755 176.065 102.085 176.125 ;
        RECT 102.755 176.065 102.925 176.825 ;
        RECT 104.165 176.755 104.485 177.215 ;
        RECT 104.685 176.575 104.935 177.005 ;
        RECT 105.225 176.775 105.635 177.215 ;
        RECT 105.805 176.835 106.820 177.035 ;
        RECT 103.095 176.405 104.345 176.575 ;
        RECT 103.095 176.285 103.425 176.405 ;
        RECT 101.755 175.895 103.655 176.065 ;
        RECT 101.395 175.555 103.315 175.725 ;
        RECT 101.395 175.535 101.715 175.555 ;
        RECT 100.945 174.875 101.275 175.385 ;
        RECT 101.545 174.925 101.715 175.535 ;
        RECT 103.485 175.385 103.655 175.895 ;
        RECT 103.825 175.825 104.005 176.235 ;
        RECT 104.175 175.645 104.345 176.405 ;
        RECT 101.885 174.665 102.215 175.355 ;
        RECT 102.445 175.215 103.655 175.385 ;
        RECT 103.825 175.335 104.345 175.645 ;
        RECT 104.515 176.235 104.935 176.575 ;
        RECT 105.225 176.235 105.635 176.565 ;
        RECT 104.515 175.465 104.705 176.235 ;
        RECT 105.805 176.105 105.975 176.835 ;
        RECT 107.120 176.665 107.290 176.995 ;
        RECT 107.460 176.835 107.790 177.215 ;
        RECT 106.145 176.285 106.495 176.655 ;
        RECT 105.805 176.065 106.225 176.105 ;
        RECT 104.875 175.895 106.225 176.065 ;
        RECT 104.875 175.735 105.125 175.895 ;
        RECT 105.635 175.465 105.885 175.725 ;
        RECT 104.515 175.215 105.885 175.465 ;
        RECT 102.445 174.925 102.685 175.215 ;
        RECT 103.485 175.135 103.655 175.215 ;
        RECT 102.885 174.665 103.305 175.045 ;
        RECT 103.485 174.885 104.115 175.135 ;
        RECT 104.585 174.665 104.915 175.045 ;
        RECT 105.085 174.925 105.255 175.215 ;
        RECT 106.055 175.050 106.225 175.895 ;
        RECT 106.675 175.725 106.895 176.595 ;
        RECT 107.120 176.475 107.815 176.665 ;
        RECT 106.395 175.345 106.895 175.725 ;
        RECT 107.065 175.675 107.475 176.295 ;
        RECT 107.645 175.505 107.815 176.475 ;
        RECT 107.120 175.335 107.815 175.505 ;
        RECT 105.435 174.665 105.815 175.045 ;
        RECT 106.055 174.880 106.885 175.050 ;
        RECT 107.120 174.835 107.290 175.335 ;
        RECT 107.460 174.665 107.790 175.165 ;
        RECT 108.005 174.835 108.230 176.955 ;
        RECT 108.400 176.835 108.730 177.215 ;
        RECT 108.900 176.665 109.070 176.955 ;
        RECT 108.405 176.495 109.070 176.665 ;
        RECT 108.405 175.505 108.635 176.495 ;
        RECT 109.330 176.445 111.000 177.215 ;
        RECT 111.170 176.465 112.380 177.215 ;
        RECT 108.805 175.675 109.155 176.325 ;
        RECT 109.330 175.755 110.080 176.275 ;
        RECT 110.250 175.925 111.000 176.445 ;
        RECT 111.170 175.755 111.690 176.295 ;
        RECT 111.860 175.925 112.380 176.465 ;
        RECT 108.405 175.335 109.070 175.505 ;
        RECT 108.400 174.665 108.730 175.165 ;
        RECT 108.900 174.835 109.070 175.335 ;
        RECT 109.330 174.665 111.000 175.755 ;
        RECT 111.170 174.665 112.380 175.755 ;
        RECT 18.165 174.495 112.465 174.665 ;
        RECT 18.250 173.405 19.460 174.495 ;
        RECT 18.250 172.695 18.770 173.235 ;
        RECT 18.940 172.865 19.460 173.405 ;
        RECT 19.630 173.405 22.220 174.495 ;
        RECT 19.630 172.885 20.840 173.405 ;
        RECT 22.430 173.355 22.660 174.495 ;
        RECT 22.830 173.345 23.160 174.325 ;
        RECT 23.330 173.355 23.540 174.495 ;
        RECT 23.770 173.405 27.280 174.495 ;
        RECT 27.455 174.070 27.790 174.495 ;
        RECT 27.960 173.890 28.145 174.295 ;
        RECT 27.480 173.715 28.145 173.890 ;
        RECT 28.350 173.715 28.680 174.495 ;
        RECT 21.010 172.715 22.220 173.235 ;
        RECT 22.410 172.935 22.740 173.185 ;
        RECT 18.250 171.945 19.460 172.695 ;
        RECT 19.630 171.945 22.220 172.715 ;
        RECT 22.430 171.945 22.660 172.765 ;
        RECT 22.910 172.745 23.160 173.345 ;
        RECT 23.770 172.885 25.460 173.405 ;
        RECT 22.830 172.115 23.160 172.745 ;
        RECT 23.330 171.945 23.540 172.765 ;
        RECT 25.630 172.715 27.280 173.235 ;
        RECT 23.770 171.945 27.280 172.715 ;
        RECT 27.480 172.685 27.820 173.715 ;
        RECT 28.850 173.525 29.120 174.295 ;
        RECT 29.345 173.625 29.630 174.495 ;
        RECT 29.800 173.865 30.060 174.325 ;
        RECT 30.235 174.035 30.490 174.495 ;
        RECT 30.660 173.865 30.920 174.325 ;
        RECT 29.800 173.695 30.920 173.865 ;
        RECT 31.090 173.695 31.400 174.495 ;
        RECT 27.990 173.355 29.120 173.525 ;
        RECT 29.800 173.445 30.060 173.695 ;
        RECT 31.570 173.525 31.880 174.325 ;
        RECT 32.105 173.625 32.390 174.495 ;
        RECT 32.560 173.865 32.820 174.325 ;
        RECT 32.995 174.035 33.250 174.495 ;
        RECT 33.420 173.865 33.680 174.325 ;
        RECT 32.560 173.695 33.680 173.865 ;
        RECT 33.850 173.695 34.160 174.495 ;
        RECT 27.990 172.855 28.240 173.355 ;
        RECT 27.480 172.515 28.165 172.685 ;
        RECT 28.420 172.605 28.780 173.185 ;
        RECT 27.455 171.945 27.790 172.345 ;
        RECT 27.960 172.115 28.165 172.515 ;
        RECT 28.950 172.445 29.120 173.355 ;
        RECT 29.305 173.275 30.060 173.445 ;
        RECT 30.850 173.355 31.880 173.525 ;
        RECT 32.560 173.445 32.820 173.695 ;
        RECT 34.330 173.525 34.640 174.325 ;
        RECT 29.305 172.765 29.710 173.275 ;
        RECT 30.850 173.105 31.020 173.355 ;
        RECT 29.880 172.935 31.020 173.105 ;
        RECT 29.305 172.595 30.955 172.765 ;
        RECT 31.190 172.615 31.540 173.185 ;
        RECT 28.375 171.945 28.650 172.425 ;
        RECT 28.860 172.115 29.120 172.445 ;
        RECT 29.350 171.945 29.630 172.425 ;
        RECT 29.800 172.205 30.060 172.595 ;
        RECT 30.235 171.945 30.490 172.425 ;
        RECT 30.660 172.205 30.955 172.595 ;
        RECT 31.710 172.445 31.880 173.355 ;
        RECT 32.065 173.275 32.820 173.445 ;
        RECT 33.610 173.355 34.640 173.525 ;
        RECT 32.065 172.765 32.470 173.275 ;
        RECT 33.610 173.105 33.780 173.355 ;
        RECT 32.640 172.935 33.780 173.105 ;
        RECT 32.065 172.595 33.715 172.765 ;
        RECT 33.950 172.615 34.300 173.185 ;
        RECT 31.135 171.945 31.410 172.425 ;
        RECT 31.580 172.115 31.880 172.445 ;
        RECT 32.110 171.945 32.390 172.425 ;
        RECT 32.560 172.205 32.820 172.595 ;
        RECT 32.995 171.945 33.250 172.425 ;
        RECT 33.420 172.205 33.715 172.595 ;
        RECT 34.470 172.445 34.640 173.355 ;
        RECT 34.810 173.330 35.100 174.495 ;
        RECT 35.350 173.565 35.530 174.325 ;
        RECT 35.710 173.735 36.040 174.495 ;
        RECT 35.350 173.395 36.025 173.565 ;
        RECT 36.210 173.420 36.480 174.325 ;
        RECT 35.855 173.250 36.025 173.395 ;
        RECT 35.290 172.845 35.630 173.215 ;
        RECT 35.855 172.920 36.130 173.250 ;
        RECT 33.895 171.945 34.170 172.425 ;
        RECT 34.340 172.115 34.640 172.445 ;
        RECT 34.810 171.945 35.100 172.670 ;
        RECT 35.855 172.665 36.025 172.920 ;
        RECT 35.360 172.495 36.025 172.665 ;
        RECT 36.300 172.620 36.480 173.420 ;
        RECT 35.360 172.115 35.530 172.495 ;
        RECT 35.710 171.945 36.040 172.325 ;
        RECT 36.220 172.115 36.480 172.620 ;
        RECT 36.650 172.685 36.910 174.310 ;
        RECT 38.660 174.045 38.990 174.495 ;
        RECT 37.090 173.655 39.700 173.865 ;
        RECT 37.090 172.855 37.310 173.655 ;
        RECT 37.550 172.855 37.850 173.475 ;
        RECT 38.020 172.855 38.350 173.475 ;
        RECT 38.520 172.855 38.840 173.475 ;
        RECT 39.010 172.855 39.360 173.475 ;
        RECT 39.530 172.685 39.700 173.655 ;
        RECT 36.650 172.515 38.490 172.685 ;
        RECT 36.920 171.945 37.250 172.340 ;
        RECT 37.420 172.160 37.620 172.515 ;
        RECT 37.790 171.945 38.120 172.345 ;
        RECT 38.290 172.170 38.490 172.515 ;
        RECT 38.660 171.945 38.990 172.685 ;
        RECT 39.225 172.515 39.700 172.685 ;
        RECT 39.870 173.355 40.210 174.325 ;
        RECT 40.380 173.355 40.550 174.495 ;
        RECT 40.820 173.695 41.070 174.495 ;
        RECT 41.715 173.525 42.045 174.325 ;
        RECT 42.345 173.695 42.675 174.495 ;
        RECT 42.845 173.525 43.175 174.325 ;
        RECT 40.740 173.355 43.175 173.525 ;
        RECT 39.870 172.745 40.045 173.355 ;
        RECT 40.740 173.105 40.910 173.355 ;
        RECT 40.215 172.935 40.910 173.105 ;
        RECT 41.085 172.935 41.505 173.135 ;
        RECT 41.675 172.935 42.005 173.135 ;
        RECT 42.175 172.935 42.505 173.135 ;
        RECT 39.225 172.265 39.395 172.515 ;
        RECT 39.870 172.115 40.210 172.745 ;
        RECT 40.380 171.945 40.630 172.745 ;
        RECT 40.820 172.595 42.045 172.765 ;
        RECT 40.820 172.115 41.150 172.595 ;
        RECT 41.320 171.945 41.545 172.405 ;
        RECT 41.715 172.115 42.045 172.595 ;
        RECT 42.675 172.725 42.845 173.355 ;
        RECT 44.015 173.305 44.270 174.185 ;
        RECT 44.440 173.355 44.745 174.495 ;
        RECT 45.085 174.115 45.415 174.495 ;
        RECT 45.595 173.945 45.765 174.235 ;
        RECT 45.935 174.035 46.185 174.495 ;
        RECT 44.965 173.775 45.765 173.945 ;
        RECT 46.355 173.985 47.225 174.325 ;
        RECT 43.030 172.935 43.380 173.185 ;
        RECT 42.675 172.115 43.175 172.725 ;
        RECT 44.015 172.655 44.225 173.305 ;
        RECT 44.965 173.185 45.135 173.775 ;
        RECT 46.355 173.605 46.525 173.985 ;
        RECT 47.460 173.865 47.630 174.325 ;
        RECT 47.800 174.035 48.170 174.495 ;
        RECT 48.465 173.895 48.635 174.235 ;
        RECT 48.805 174.065 49.135 174.495 ;
        RECT 49.370 173.895 49.540 174.235 ;
        RECT 45.305 173.435 46.525 173.605 ;
        RECT 46.695 173.525 47.155 173.815 ;
        RECT 47.460 173.695 48.020 173.865 ;
        RECT 48.465 173.725 49.540 173.895 ;
        RECT 49.710 173.995 50.390 174.325 ;
        RECT 50.605 173.995 50.855 174.325 ;
        RECT 51.025 174.035 51.275 174.495 ;
        RECT 47.850 173.555 48.020 173.695 ;
        RECT 46.695 173.515 47.660 173.525 ;
        RECT 46.355 173.345 46.525 173.435 ;
        RECT 46.985 173.355 47.660 173.515 ;
        RECT 44.395 173.155 45.135 173.185 ;
        RECT 44.395 172.855 45.310 173.155 ;
        RECT 44.985 172.680 45.310 172.855 ;
        RECT 44.015 172.125 44.270 172.655 ;
        RECT 44.440 171.945 44.745 172.405 ;
        RECT 44.990 172.325 45.310 172.680 ;
        RECT 45.480 172.895 46.020 173.265 ;
        RECT 46.355 173.175 46.760 173.345 ;
        RECT 45.480 172.495 45.720 172.895 ;
        RECT 46.200 172.725 46.420 173.005 ;
        RECT 45.890 172.555 46.420 172.725 ;
        RECT 45.890 172.325 46.060 172.555 ;
        RECT 46.590 172.395 46.760 173.175 ;
        RECT 46.930 172.565 47.280 173.185 ;
        RECT 47.450 172.565 47.660 173.355 ;
        RECT 47.850 173.385 49.350 173.555 ;
        RECT 47.850 172.695 48.020 173.385 ;
        RECT 49.710 173.215 49.880 173.995 ;
        RECT 50.685 173.865 50.855 173.995 ;
        RECT 48.190 173.045 49.880 173.215 ;
        RECT 50.050 173.435 50.515 173.825 ;
        RECT 50.685 173.695 51.080 173.865 ;
        RECT 48.190 172.865 48.360 173.045 ;
        RECT 44.990 172.155 46.060 172.325 ;
        RECT 46.230 171.945 46.420 172.385 ;
        RECT 46.590 172.115 47.540 172.395 ;
        RECT 47.850 172.305 48.110 172.695 ;
        RECT 48.530 172.625 49.320 172.875 ;
        RECT 47.760 172.135 48.110 172.305 ;
        RECT 48.320 171.945 48.650 172.405 ;
        RECT 49.525 172.335 49.695 173.045 ;
        RECT 50.050 172.845 50.220 173.435 ;
        RECT 49.865 172.625 50.220 172.845 ;
        RECT 50.390 172.625 50.740 173.245 ;
        RECT 50.910 172.335 51.080 173.695 ;
        RECT 51.445 173.525 51.770 174.310 ;
        RECT 51.250 172.475 51.710 173.525 ;
        RECT 49.525 172.165 50.380 172.335 ;
        RECT 50.585 172.165 51.080 172.335 ;
        RECT 51.250 171.945 51.580 172.305 ;
        RECT 51.940 172.205 52.110 174.325 ;
        RECT 52.280 173.995 52.610 174.495 ;
        RECT 52.780 173.825 53.035 174.325 ;
        RECT 52.285 173.655 53.035 173.825 ;
        RECT 52.285 172.665 52.515 173.655 ;
        RECT 52.685 172.835 53.035 173.485 ;
        RECT 53.670 173.405 56.260 174.495 ;
        RECT 56.430 173.735 56.945 174.145 ;
        RECT 57.180 173.735 57.350 174.495 ;
        RECT 57.520 174.155 59.550 174.325 ;
        RECT 53.670 172.885 54.880 173.405 ;
        RECT 55.050 172.715 56.260 173.235 ;
        RECT 56.430 172.925 56.770 173.735 ;
        RECT 57.520 173.490 57.690 174.155 ;
        RECT 58.085 173.815 59.210 173.985 ;
        RECT 56.940 173.300 57.690 173.490 ;
        RECT 57.860 173.475 58.870 173.645 ;
        RECT 56.430 172.755 57.660 172.925 ;
        RECT 52.285 172.495 53.035 172.665 ;
        RECT 52.280 171.945 52.610 172.325 ;
        RECT 52.780 172.205 53.035 172.495 ;
        RECT 53.670 171.945 56.260 172.715 ;
        RECT 56.705 172.150 56.950 172.755 ;
        RECT 57.170 171.945 57.680 172.480 ;
        RECT 57.860 172.115 58.050 173.475 ;
        RECT 58.220 172.455 58.495 173.275 ;
        RECT 58.700 172.675 58.870 173.475 ;
        RECT 59.040 172.685 59.210 173.815 ;
        RECT 59.380 173.185 59.550 174.155 ;
        RECT 59.720 173.355 59.890 174.495 ;
        RECT 60.060 173.355 60.395 174.325 ;
        RECT 59.380 172.855 59.575 173.185 ;
        RECT 59.800 172.855 60.055 173.185 ;
        RECT 59.800 172.685 59.970 172.855 ;
        RECT 60.225 172.685 60.395 173.355 ;
        RECT 60.570 173.330 60.860 174.495 ;
        RECT 61.120 173.825 61.290 174.325 ;
        RECT 61.460 173.995 61.790 174.495 ;
        RECT 61.120 173.655 61.785 173.825 ;
        RECT 61.035 172.835 61.385 173.485 ;
        RECT 59.040 172.515 59.970 172.685 ;
        RECT 59.040 172.480 59.215 172.515 ;
        RECT 58.220 172.285 58.500 172.455 ;
        RECT 58.220 172.115 58.495 172.285 ;
        RECT 58.685 172.115 59.215 172.480 ;
        RECT 59.640 171.945 59.970 172.345 ;
        RECT 60.140 172.115 60.395 172.685 ;
        RECT 60.570 171.945 60.860 172.670 ;
        RECT 61.555 172.665 61.785 173.655 ;
        RECT 61.120 172.495 61.785 172.665 ;
        RECT 61.120 172.205 61.290 172.495 ;
        RECT 61.460 171.945 61.790 172.325 ;
        RECT 61.960 172.205 62.185 174.325 ;
        RECT 62.400 173.995 62.730 174.495 ;
        RECT 62.900 173.825 63.070 174.325 ;
        RECT 63.305 174.110 64.135 174.280 ;
        RECT 64.375 174.115 64.755 174.495 ;
        RECT 62.375 173.655 63.070 173.825 ;
        RECT 62.375 172.685 62.545 173.655 ;
        RECT 62.715 172.865 63.125 173.485 ;
        RECT 63.295 173.435 63.795 173.815 ;
        RECT 62.375 172.495 63.070 172.685 ;
        RECT 63.295 172.565 63.515 173.435 ;
        RECT 63.965 173.265 64.135 174.110 ;
        RECT 64.935 173.945 65.105 174.235 ;
        RECT 65.275 174.115 65.605 174.495 ;
        RECT 66.075 174.025 66.705 174.275 ;
        RECT 66.885 174.115 67.305 174.495 ;
        RECT 66.535 173.945 66.705 174.025 ;
        RECT 67.505 173.945 67.745 174.235 ;
        RECT 64.305 173.695 65.675 173.945 ;
        RECT 64.305 173.435 64.555 173.695 ;
        RECT 65.065 173.265 65.315 173.425 ;
        RECT 63.965 173.095 65.315 173.265 ;
        RECT 63.965 173.055 64.385 173.095 ;
        RECT 63.695 172.505 64.045 172.875 ;
        RECT 62.400 171.945 62.730 172.325 ;
        RECT 62.900 172.165 63.070 172.495 ;
        RECT 64.215 172.325 64.385 173.055 ;
        RECT 65.485 172.925 65.675 173.695 ;
        RECT 64.555 172.595 64.965 172.925 ;
        RECT 65.255 172.585 65.675 172.925 ;
        RECT 65.845 173.515 66.365 173.825 ;
        RECT 66.535 173.775 67.745 173.945 ;
        RECT 67.975 173.805 68.305 174.495 ;
        RECT 65.845 172.755 66.015 173.515 ;
        RECT 66.185 172.925 66.365 173.335 ;
        RECT 66.535 173.265 66.705 173.775 ;
        RECT 68.475 173.625 68.645 174.235 ;
        RECT 68.915 173.775 69.245 174.285 ;
        RECT 68.475 173.605 68.795 173.625 ;
        RECT 66.875 173.435 68.795 173.605 ;
        RECT 66.535 173.095 68.435 173.265 ;
        RECT 66.765 172.755 67.095 172.875 ;
        RECT 65.845 172.585 67.095 172.755 ;
        RECT 63.370 172.125 64.385 172.325 ;
        RECT 64.555 171.945 64.965 172.385 ;
        RECT 65.255 172.155 65.505 172.585 ;
        RECT 65.705 171.945 66.025 172.405 ;
        RECT 67.265 172.335 67.435 173.095 ;
        RECT 68.105 173.035 68.435 173.095 ;
        RECT 67.625 172.865 67.955 172.925 ;
        RECT 67.625 172.595 68.285 172.865 ;
        RECT 68.605 172.540 68.795 173.435 ;
        RECT 66.585 172.165 67.435 172.335 ;
        RECT 67.635 171.945 68.295 172.425 ;
        RECT 68.475 172.210 68.795 172.540 ;
        RECT 68.995 173.185 69.245 173.775 ;
        RECT 69.425 173.695 69.710 174.495 ;
        RECT 69.890 174.155 70.145 174.185 ;
        RECT 69.890 173.985 70.230 174.155 ;
        RECT 69.890 173.515 70.145 173.985 ;
        RECT 68.995 172.855 69.795 173.185 ;
        RECT 68.995 172.205 69.245 172.855 ;
        RECT 69.965 172.655 70.145 173.515 ;
        RECT 69.425 171.945 69.710 172.405 ;
        RECT 69.890 172.125 70.145 172.655 ;
        RECT 70.690 173.355 71.030 174.325 ;
        RECT 71.200 173.355 71.370 174.495 ;
        RECT 71.640 173.695 71.890 174.495 ;
        RECT 72.535 173.525 72.865 174.325 ;
        RECT 73.165 173.695 73.495 174.495 ;
        RECT 73.665 173.525 73.995 174.325 ;
        RECT 75.295 174.060 80.640 174.495 ;
        RECT 71.560 173.355 73.995 173.525 ;
        RECT 70.690 172.745 70.865 173.355 ;
        RECT 71.560 173.105 71.730 173.355 ;
        RECT 71.035 172.935 71.730 173.105 ;
        RECT 71.905 172.935 72.325 173.135 ;
        RECT 72.495 172.935 72.825 173.135 ;
        RECT 72.995 172.935 73.325 173.135 ;
        RECT 70.690 172.115 71.030 172.745 ;
        RECT 71.200 171.945 71.450 172.745 ;
        RECT 71.640 172.595 72.865 172.765 ;
        RECT 71.640 172.115 71.970 172.595 ;
        RECT 72.140 171.945 72.365 172.405 ;
        RECT 72.535 172.115 72.865 172.595 ;
        RECT 73.495 172.725 73.665 173.355 ;
        RECT 73.850 172.935 74.200 173.185 ;
        RECT 76.885 172.810 77.235 174.060 ;
        RECT 80.850 173.355 81.080 174.495 ;
        RECT 81.250 173.345 81.580 174.325 ;
        RECT 81.750 173.355 81.960 174.495 ;
        RECT 82.190 173.735 82.705 174.145 ;
        RECT 82.940 173.735 83.110 174.495 ;
        RECT 83.280 174.155 85.310 174.325 ;
        RECT 73.495 172.115 73.995 172.725 ;
        RECT 78.715 172.490 79.055 173.320 ;
        RECT 80.830 172.935 81.160 173.185 ;
        RECT 75.295 171.945 80.640 172.490 ;
        RECT 80.850 171.945 81.080 172.765 ;
        RECT 81.330 172.745 81.580 173.345 ;
        RECT 82.190 172.925 82.530 173.735 ;
        RECT 83.280 173.490 83.450 174.155 ;
        RECT 83.845 173.815 84.970 173.985 ;
        RECT 82.700 173.300 83.450 173.490 ;
        RECT 83.620 173.475 84.630 173.645 ;
        RECT 81.250 172.115 81.580 172.745 ;
        RECT 81.750 171.945 81.960 172.765 ;
        RECT 82.190 172.755 83.420 172.925 ;
        RECT 82.465 172.150 82.710 172.755 ;
        RECT 82.930 171.945 83.440 172.480 ;
        RECT 83.620 172.115 83.810 173.475 ;
        RECT 83.980 173.135 84.255 173.275 ;
        RECT 83.980 172.965 84.260 173.135 ;
        RECT 83.980 172.115 84.255 172.965 ;
        RECT 84.460 172.675 84.630 173.475 ;
        RECT 84.800 172.685 84.970 173.815 ;
        RECT 85.140 173.185 85.310 174.155 ;
        RECT 85.480 173.355 85.650 174.495 ;
        RECT 85.820 173.355 86.155 174.325 ;
        RECT 85.140 172.855 85.335 173.185 ;
        RECT 85.560 172.855 85.815 173.185 ;
        RECT 85.560 172.685 85.730 172.855 ;
        RECT 85.985 172.685 86.155 173.355 ;
        RECT 86.330 173.330 86.620 174.495 ;
        RECT 86.995 173.525 87.325 174.325 ;
        RECT 87.495 173.695 87.825 174.495 ;
        RECT 88.125 173.525 88.455 174.325 ;
        RECT 89.100 173.695 89.350 174.495 ;
        RECT 86.995 173.355 89.430 173.525 ;
        RECT 89.620 173.355 89.790 174.495 ;
        RECT 89.960 173.355 90.300 174.325 ;
        RECT 86.790 172.935 87.140 173.185 ;
        RECT 87.325 172.725 87.495 173.355 ;
        RECT 87.665 172.935 87.995 173.135 ;
        RECT 88.165 172.935 88.495 173.135 ;
        RECT 88.665 172.935 89.085 173.135 ;
        RECT 89.260 173.105 89.430 173.355 ;
        RECT 89.260 172.935 89.955 173.105 ;
        RECT 84.800 172.515 85.730 172.685 ;
        RECT 84.800 172.480 84.975 172.515 ;
        RECT 84.445 172.115 84.975 172.480 ;
        RECT 85.400 171.945 85.730 172.345 ;
        RECT 85.900 172.115 86.155 172.685 ;
        RECT 86.330 171.945 86.620 172.670 ;
        RECT 86.995 172.115 87.495 172.725 ;
        RECT 88.125 172.595 89.350 172.765 ;
        RECT 90.125 172.745 90.300 173.355 ;
        RECT 90.930 173.405 92.600 174.495 ;
        RECT 92.770 173.735 93.285 174.145 ;
        RECT 93.520 173.735 93.690 174.495 ;
        RECT 93.860 174.155 95.890 174.325 ;
        RECT 90.930 172.885 91.680 173.405 ;
        RECT 88.125 172.115 88.455 172.595 ;
        RECT 88.625 171.945 88.850 172.405 ;
        RECT 89.020 172.115 89.350 172.595 ;
        RECT 89.540 171.945 89.790 172.745 ;
        RECT 89.960 172.115 90.300 172.745 ;
        RECT 91.850 172.715 92.600 173.235 ;
        RECT 92.770 172.925 93.110 173.735 ;
        RECT 93.860 173.490 94.030 174.155 ;
        RECT 94.425 173.815 95.550 173.985 ;
        RECT 93.280 173.300 94.030 173.490 ;
        RECT 94.200 173.475 95.210 173.645 ;
        RECT 92.770 172.755 94.000 172.925 ;
        RECT 90.930 171.945 92.600 172.715 ;
        RECT 93.045 172.150 93.290 172.755 ;
        RECT 93.510 171.945 94.020 172.480 ;
        RECT 94.200 172.115 94.390 173.475 ;
        RECT 94.560 173.135 94.835 173.275 ;
        RECT 94.560 172.965 94.840 173.135 ;
        RECT 94.560 172.115 94.835 172.965 ;
        RECT 95.040 172.675 95.210 173.475 ;
        RECT 95.380 172.685 95.550 173.815 ;
        RECT 95.720 173.185 95.890 174.155 ;
        RECT 96.060 173.355 96.230 174.495 ;
        RECT 96.400 173.355 96.735 174.325 ;
        RECT 95.720 172.855 95.915 173.185 ;
        RECT 96.140 172.855 96.395 173.185 ;
        RECT 96.140 172.685 96.310 172.855 ;
        RECT 96.565 172.685 96.735 173.355 ;
        RECT 96.910 173.735 97.425 174.145 ;
        RECT 97.660 173.735 97.830 174.495 ;
        RECT 98.000 174.155 100.030 174.325 ;
        RECT 96.910 172.925 97.250 173.735 ;
        RECT 98.000 173.490 98.170 174.155 ;
        RECT 98.565 173.815 99.690 173.985 ;
        RECT 97.420 173.300 98.170 173.490 ;
        RECT 98.340 173.475 99.350 173.645 ;
        RECT 96.910 172.755 98.140 172.925 ;
        RECT 95.380 172.515 96.310 172.685 ;
        RECT 95.380 172.480 95.555 172.515 ;
        RECT 95.025 172.115 95.555 172.480 ;
        RECT 95.980 171.945 96.310 172.345 ;
        RECT 96.480 172.115 96.735 172.685 ;
        RECT 97.185 172.150 97.430 172.755 ;
        RECT 97.650 171.945 98.160 172.480 ;
        RECT 98.340 172.115 98.530 173.475 ;
        RECT 98.700 172.795 98.975 173.275 ;
        RECT 98.700 172.625 98.980 172.795 ;
        RECT 99.180 172.675 99.350 173.475 ;
        RECT 99.520 172.685 99.690 173.815 ;
        RECT 99.860 173.185 100.030 174.155 ;
        RECT 100.200 173.355 100.370 174.495 ;
        RECT 100.540 173.355 100.875 174.325 ;
        RECT 99.860 172.855 100.055 173.185 ;
        RECT 100.280 172.855 100.535 173.185 ;
        RECT 100.280 172.685 100.450 172.855 ;
        RECT 100.705 172.685 100.875 173.355 ;
        RECT 98.700 172.115 98.975 172.625 ;
        RECT 99.520 172.515 100.450 172.685 ;
        RECT 99.520 172.480 99.695 172.515 ;
        RECT 99.165 172.115 99.695 172.480 ;
        RECT 100.120 171.945 100.450 172.345 ;
        RECT 100.620 172.115 100.875 172.685 ;
        RECT 101.425 173.515 101.680 174.185 ;
        RECT 101.860 173.695 102.145 174.495 ;
        RECT 102.325 173.775 102.655 174.285 ;
        RECT 101.425 172.655 101.605 173.515 ;
        RECT 102.325 173.185 102.575 173.775 ;
        RECT 102.925 173.625 103.095 174.235 ;
        RECT 103.265 173.805 103.595 174.495 ;
        RECT 103.825 173.945 104.065 174.235 ;
        RECT 104.265 174.115 104.685 174.495 ;
        RECT 104.865 174.025 105.495 174.275 ;
        RECT 105.965 174.115 106.295 174.495 ;
        RECT 104.865 173.945 105.035 174.025 ;
        RECT 106.465 173.945 106.635 174.235 ;
        RECT 106.815 174.115 107.195 174.495 ;
        RECT 107.435 174.110 108.265 174.280 ;
        RECT 103.825 173.775 105.035 173.945 ;
        RECT 101.775 172.855 102.575 173.185 ;
        RECT 101.425 172.455 101.680 172.655 ;
        RECT 101.340 172.285 101.680 172.455 ;
        RECT 101.425 172.125 101.680 172.285 ;
        RECT 101.860 171.945 102.145 172.405 ;
        RECT 102.325 172.205 102.575 172.855 ;
        RECT 102.775 173.605 103.095 173.625 ;
        RECT 102.775 173.435 104.695 173.605 ;
        RECT 102.775 172.540 102.965 173.435 ;
        RECT 104.865 173.265 105.035 173.775 ;
        RECT 105.205 173.515 105.725 173.825 ;
        RECT 103.135 173.095 105.035 173.265 ;
        RECT 103.135 173.035 103.465 173.095 ;
        RECT 103.615 172.865 103.945 172.925 ;
        RECT 103.285 172.595 103.945 172.865 ;
        RECT 102.775 172.210 103.095 172.540 ;
        RECT 103.275 171.945 103.935 172.425 ;
        RECT 104.135 172.335 104.305 173.095 ;
        RECT 105.205 172.925 105.385 173.335 ;
        RECT 104.475 172.755 104.805 172.875 ;
        RECT 105.555 172.755 105.725 173.515 ;
        RECT 104.475 172.585 105.725 172.755 ;
        RECT 105.895 173.695 107.265 173.945 ;
        RECT 105.895 172.925 106.085 173.695 ;
        RECT 107.015 173.435 107.265 173.695 ;
        RECT 106.255 173.265 106.505 173.425 ;
        RECT 107.435 173.265 107.605 174.110 ;
        RECT 108.500 173.825 108.670 174.325 ;
        RECT 108.840 173.995 109.170 174.495 ;
        RECT 107.775 173.435 108.275 173.815 ;
        RECT 108.500 173.655 109.195 173.825 ;
        RECT 106.255 173.095 107.605 173.265 ;
        RECT 107.185 173.055 107.605 173.095 ;
        RECT 105.895 172.585 106.315 172.925 ;
        RECT 106.605 172.595 107.015 172.925 ;
        RECT 104.135 172.165 104.985 172.335 ;
        RECT 105.545 171.945 105.865 172.405 ;
        RECT 106.065 172.155 106.315 172.585 ;
        RECT 106.605 171.945 107.015 172.385 ;
        RECT 107.185 172.325 107.355 173.055 ;
        RECT 107.525 172.505 107.875 172.875 ;
        RECT 108.055 172.565 108.275 173.435 ;
        RECT 108.445 172.865 108.855 173.485 ;
        RECT 109.025 172.685 109.195 173.655 ;
        RECT 108.500 172.495 109.195 172.685 ;
        RECT 107.185 172.125 108.200 172.325 ;
        RECT 108.500 172.165 108.670 172.495 ;
        RECT 108.840 171.945 109.170 172.325 ;
        RECT 109.385 172.205 109.610 174.325 ;
        RECT 109.780 173.995 110.110 174.495 ;
        RECT 110.280 173.825 110.450 174.325 ;
        RECT 109.785 173.655 110.450 173.825 ;
        RECT 109.785 172.665 110.015 173.655 ;
        RECT 110.185 172.835 110.535 173.485 ;
        RECT 111.170 173.405 112.380 174.495 ;
        RECT 111.170 172.865 111.690 173.405 ;
        RECT 111.860 172.695 112.380 173.235 ;
        RECT 109.785 172.495 110.450 172.665 ;
        RECT 109.780 171.945 110.110 172.325 ;
        RECT 110.280 172.205 110.450 172.495 ;
        RECT 111.170 171.945 112.380 172.695 ;
        RECT 18.165 171.775 112.465 171.945 ;
        RECT 18.250 171.025 19.460 171.775 ;
        RECT 20.640 171.225 20.810 171.605 ;
        RECT 20.990 171.395 21.320 171.775 ;
        RECT 20.640 171.055 21.305 171.225 ;
        RECT 21.500 171.100 21.760 171.605 ;
        RECT 18.250 170.485 18.770 171.025 ;
        RECT 18.940 170.315 19.460 170.855 ;
        RECT 20.570 170.505 20.910 170.875 ;
        RECT 21.135 170.800 21.305 171.055 ;
        RECT 21.135 170.470 21.410 170.800 ;
        RECT 21.135 170.325 21.305 170.470 ;
        RECT 18.250 169.225 19.460 170.315 ;
        RECT 20.630 170.155 21.305 170.325 ;
        RECT 21.580 170.300 21.760 171.100 ;
        RECT 21.930 171.050 22.220 171.775 ;
        RECT 22.940 171.225 23.110 171.605 ;
        RECT 23.325 171.395 23.655 171.775 ;
        RECT 22.940 171.055 23.655 171.225 ;
        RECT 22.850 170.505 23.205 170.875 ;
        RECT 23.485 170.865 23.655 171.055 ;
        RECT 23.825 171.030 24.080 171.605 ;
        RECT 23.485 170.535 23.740 170.865 ;
        RECT 20.630 169.395 20.810 170.155 ;
        RECT 20.990 169.225 21.320 169.985 ;
        RECT 21.490 169.395 21.760 170.300 ;
        RECT 21.930 169.225 22.220 170.390 ;
        RECT 23.485 170.325 23.655 170.535 ;
        RECT 22.940 170.155 23.655 170.325 ;
        RECT 23.910 170.300 24.080 171.030 ;
        RECT 24.255 170.935 24.515 171.775 ;
        RECT 25.670 170.955 25.880 171.775 ;
        RECT 26.050 170.975 26.380 171.605 ;
        RECT 26.050 170.375 26.300 170.975 ;
        RECT 26.550 170.955 26.780 171.775 ;
        RECT 26.995 171.225 27.250 171.515 ;
        RECT 27.420 171.395 27.750 171.775 ;
        RECT 26.995 171.055 27.745 171.225 ;
        RECT 26.470 170.535 26.800 170.785 ;
        RECT 22.940 169.395 23.110 170.155 ;
        RECT 23.325 169.225 23.655 169.985 ;
        RECT 23.825 169.395 24.080 170.300 ;
        RECT 24.255 169.225 24.515 170.375 ;
        RECT 25.670 169.225 25.880 170.365 ;
        RECT 26.050 169.395 26.380 170.375 ;
        RECT 26.550 169.225 26.780 170.365 ;
        RECT 26.995 170.235 27.345 170.885 ;
        RECT 27.515 170.065 27.745 171.055 ;
        RECT 26.995 169.895 27.745 170.065 ;
        RECT 26.995 169.395 27.250 169.895 ;
        RECT 27.420 169.225 27.750 169.725 ;
        RECT 27.920 169.395 28.090 171.515 ;
        RECT 28.450 171.415 28.780 171.775 ;
        RECT 28.950 171.385 29.445 171.555 ;
        RECT 29.650 171.385 30.505 171.555 ;
        RECT 28.320 170.195 28.780 171.245 ;
        RECT 28.260 169.410 28.585 170.195 ;
        RECT 28.950 170.025 29.120 171.385 ;
        RECT 29.290 170.475 29.640 171.095 ;
        RECT 29.810 170.875 30.165 171.095 ;
        RECT 29.810 170.285 29.980 170.875 ;
        RECT 30.335 170.675 30.505 171.385 ;
        RECT 31.380 171.315 31.710 171.775 ;
        RECT 31.920 171.415 32.270 171.585 ;
        RECT 30.710 170.845 31.500 171.095 ;
        RECT 31.920 171.025 32.180 171.415 ;
        RECT 32.490 171.325 33.440 171.605 ;
        RECT 33.610 171.335 33.800 171.775 ;
        RECT 33.970 171.395 35.040 171.565 ;
        RECT 31.670 170.675 31.840 170.855 ;
        RECT 28.950 169.855 29.345 170.025 ;
        RECT 29.515 169.895 29.980 170.285 ;
        RECT 30.150 170.505 31.840 170.675 ;
        RECT 29.175 169.725 29.345 169.855 ;
        RECT 30.150 169.725 30.320 170.505 ;
        RECT 32.010 170.335 32.180 171.025 ;
        RECT 30.680 170.165 32.180 170.335 ;
        RECT 32.370 170.365 32.580 171.155 ;
        RECT 32.750 170.535 33.100 171.155 ;
        RECT 33.270 170.545 33.440 171.325 ;
        RECT 33.970 171.165 34.140 171.395 ;
        RECT 33.610 170.995 34.140 171.165 ;
        RECT 33.610 170.715 33.830 170.995 ;
        RECT 34.310 170.825 34.550 171.225 ;
        RECT 33.270 170.375 33.675 170.545 ;
        RECT 34.010 170.455 34.550 170.825 ;
        RECT 34.720 171.040 35.040 171.395 ;
        RECT 35.285 171.315 35.590 171.775 ;
        RECT 35.760 171.065 36.015 171.595 ;
        RECT 34.720 170.865 35.045 171.040 ;
        RECT 34.720 170.565 35.635 170.865 ;
        RECT 34.895 170.535 35.635 170.565 ;
        RECT 32.370 170.205 33.045 170.365 ;
        RECT 33.505 170.285 33.675 170.375 ;
        RECT 32.370 170.195 33.335 170.205 ;
        RECT 32.010 170.025 32.180 170.165 ;
        RECT 28.755 169.225 29.005 169.685 ;
        RECT 29.175 169.395 29.425 169.725 ;
        RECT 29.640 169.395 30.320 169.725 ;
        RECT 30.490 169.825 31.565 169.995 ;
        RECT 32.010 169.855 32.570 170.025 ;
        RECT 32.875 169.905 33.335 170.195 ;
        RECT 33.505 170.115 34.725 170.285 ;
        RECT 30.490 169.485 30.660 169.825 ;
        RECT 30.895 169.225 31.225 169.655 ;
        RECT 31.395 169.485 31.565 169.825 ;
        RECT 31.860 169.225 32.230 169.685 ;
        RECT 32.400 169.395 32.570 169.855 ;
        RECT 33.505 169.735 33.675 170.115 ;
        RECT 34.895 169.945 35.065 170.535 ;
        RECT 35.805 170.415 36.015 171.065 ;
        RECT 36.280 171.225 36.450 171.605 ;
        RECT 36.630 171.395 36.960 171.775 ;
        RECT 36.280 171.055 36.945 171.225 ;
        RECT 37.140 171.100 37.400 171.605 ;
        RECT 36.210 170.505 36.550 170.875 ;
        RECT 36.775 170.800 36.945 171.055 ;
        RECT 32.805 169.395 33.675 169.735 ;
        RECT 34.265 169.775 35.065 169.945 ;
        RECT 33.845 169.225 34.095 169.685 ;
        RECT 34.265 169.485 34.435 169.775 ;
        RECT 34.615 169.225 34.945 169.605 ;
        RECT 35.285 169.225 35.590 170.365 ;
        RECT 35.760 169.535 36.015 170.415 ;
        RECT 36.775 170.470 37.050 170.800 ;
        RECT 36.775 170.325 36.945 170.470 ;
        RECT 36.270 170.155 36.945 170.325 ;
        RECT 37.220 170.300 37.400 171.100 ;
        RECT 36.270 169.395 36.450 170.155 ;
        RECT 36.630 169.225 36.960 169.985 ;
        RECT 37.130 169.395 37.400 170.300 ;
        RECT 37.570 170.975 37.910 171.605 ;
        RECT 38.080 170.975 38.330 171.775 ;
        RECT 38.520 171.125 38.850 171.605 ;
        RECT 39.020 171.315 39.245 171.775 ;
        RECT 39.415 171.125 39.745 171.605 ;
        RECT 37.570 170.415 37.745 170.975 ;
        RECT 38.520 170.955 39.745 171.125 ;
        RECT 40.375 170.995 40.875 171.605 ;
        RECT 37.915 170.615 38.610 170.785 ;
        RECT 37.570 170.365 37.800 170.415 ;
        RECT 38.440 170.365 38.610 170.615 ;
        RECT 38.785 170.585 39.205 170.785 ;
        RECT 39.375 170.585 39.705 170.785 ;
        RECT 39.875 170.585 40.205 170.785 ;
        RECT 40.375 170.365 40.545 170.995 ;
        RECT 42.230 170.955 42.440 171.775 ;
        RECT 42.610 170.975 42.940 171.605 ;
        RECT 40.730 170.535 41.080 170.785 ;
        RECT 42.610 170.375 42.860 170.975 ;
        RECT 43.110 170.955 43.340 171.775 ;
        RECT 43.825 170.965 44.070 171.570 ;
        RECT 44.290 171.240 44.800 171.775 ;
        RECT 43.550 170.795 44.780 170.965 ;
        RECT 43.030 170.535 43.360 170.785 ;
        RECT 37.570 169.395 37.910 170.365 ;
        RECT 38.080 169.225 38.250 170.365 ;
        RECT 38.440 170.195 40.875 170.365 ;
        RECT 38.520 169.225 38.770 170.025 ;
        RECT 39.415 169.395 39.745 170.195 ;
        RECT 40.045 169.225 40.375 170.025 ;
        RECT 40.545 169.395 40.875 170.195 ;
        RECT 42.230 169.225 42.440 170.365 ;
        RECT 42.610 169.395 42.940 170.375 ;
        RECT 43.110 169.225 43.340 170.365 ;
        RECT 43.550 169.985 43.890 170.795 ;
        RECT 44.060 170.230 44.810 170.420 ;
        RECT 43.550 169.575 44.065 169.985 ;
        RECT 44.300 169.225 44.470 169.985 ;
        RECT 44.640 169.565 44.810 170.230 ;
        RECT 44.980 170.245 45.170 171.605 ;
        RECT 45.340 170.755 45.615 171.605 ;
        RECT 45.805 171.240 46.335 171.605 ;
        RECT 46.760 171.375 47.090 171.775 ;
        RECT 46.160 171.205 46.335 171.240 ;
        RECT 45.340 170.585 45.620 170.755 ;
        RECT 45.340 170.445 45.615 170.585 ;
        RECT 45.820 170.245 45.990 171.045 ;
        RECT 44.980 170.075 45.990 170.245 ;
        RECT 46.160 171.035 47.090 171.205 ;
        RECT 47.260 171.035 47.515 171.605 ;
        RECT 47.690 171.050 47.980 171.775 ;
        RECT 48.265 171.145 48.550 171.605 ;
        RECT 48.720 171.315 48.990 171.775 ;
        RECT 46.160 169.905 46.330 171.035 ;
        RECT 46.920 170.865 47.090 171.035 ;
        RECT 45.205 169.735 46.330 169.905 ;
        RECT 46.500 170.535 46.695 170.865 ;
        RECT 46.920 170.535 47.175 170.865 ;
        RECT 46.500 169.565 46.670 170.535 ;
        RECT 47.345 170.365 47.515 171.035 ;
        RECT 48.265 170.975 49.220 171.145 ;
        RECT 44.640 169.395 46.670 169.565 ;
        RECT 46.840 169.225 47.010 170.365 ;
        RECT 47.180 169.395 47.515 170.365 ;
        RECT 47.690 169.225 47.980 170.390 ;
        RECT 48.150 170.245 48.840 170.805 ;
        RECT 49.010 170.075 49.220 170.975 ;
        RECT 48.265 169.855 49.220 170.075 ;
        RECT 49.390 170.805 49.790 171.605 ;
        RECT 49.980 171.145 50.260 171.605 ;
        RECT 50.780 171.315 51.105 171.775 ;
        RECT 49.980 170.975 51.105 171.145 ;
        RECT 51.275 171.035 51.660 171.605 ;
        RECT 50.655 170.865 51.105 170.975 ;
        RECT 49.390 170.245 50.485 170.805 ;
        RECT 50.655 170.535 51.210 170.865 ;
        RECT 48.265 169.395 48.550 169.855 ;
        RECT 48.720 169.225 48.990 169.685 ;
        RECT 49.390 169.395 49.790 170.245 ;
        RECT 50.655 170.075 51.105 170.535 ;
        RECT 51.380 170.365 51.660 171.035 ;
        RECT 51.835 170.935 52.095 171.775 ;
        RECT 52.270 171.030 52.525 171.605 ;
        RECT 52.695 171.395 53.025 171.775 ;
        RECT 53.240 171.225 53.410 171.605 ;
        RECT 52.695 171.055 53.410 171.225 ;
        RECT 49.980 169.855 51.105 170.075 ;
        RECT 49.980 169.395 50.260 169.855 ;
        RECT 50.780 169.225 51.105 169.685 ;
        RECT 51.275 169.395 51.660 170.365 ;
        RECT 51.835 169.225 52.095 170.375 ;
        RECT 52.270 170.300 52.440 171.030 ;
        RECT 52.695 170.865 52.865 171.055 ;
        RECT 53.730 170.955 53.940 171.775 ;
        RECT 54.110 170.975 54.440 171.605 ;
        RECT 52.610 170.535 52.865 170.865 ;
        RECT 52.695 170.325 52.865 170.535 ;
        RECT 53.145 170.505 53.500 170.875 ;
        RECT 54.110 170.375 54.360 170.975 ;
        RECT 54.610 170.955 54.840 171.775 ;
        RECT 55.425 171.435 55.680 171.595 ;
        RECT 55.340 171.265 55.680 171.435 ;
        RECT 55.860 171.315 56.145 171.775 ;
        RECT 55.425 171.065 55.680 171.265 ;
        RECT 54.530 170.535 54.860 170.785 ;
        RECT 52.270 169.395 52.525 170.300 ;
        RECT 52.695 170.155 53.410 170.325 ;
        RECT 52.695 169.225 53.025 169.985 ;
        RECT 53.240 169.395 53.410 170.155 ;
        RECT 53.730 169.225 53.940 170.365 ;
        RECT 54.110 169.395 54.440 170.375 ;
        RECT 54.610 169.225 54.840 170.365 ;
        RECT 55.425 170.205 55.605 171.065 ;
        RECT 56.325 170.865 56.575 171.515 ;
        RECT 55.775 170.535 56.575 170.865 ;
        RECT 55.425 169.535 55.680 170.205 ;
        RECT 55.860 169.225 56.145 170.025 ;
        RECT 56.325 169.945 56.575 170.535 ;
        RECT 56.775 171.180 57.095 171.510 ;
        RECT 57.275 171.295 57.935 171.775 ;
        RECT 58.135 171.385 58.985 171.555 ;
        RECT 56.775 170.285 56.965 171.180 ;
        RECT 57.285 170.855 57.945 171.125 ;
        RECT 57.615 170.795 57.945 170.855 ;
        RECT 57.135 170.625 57.465 170.685 ;
        RECT 58.135 170.625 58.305 171.385 ;
        RECT 59.545 171.315 59.865 171.775 ;
        RECT 60.065 171.135 60.315 171.565 ;
        RECT 60.605 171.335 61.015 171.775 ;
        RECT 61.185 171.395 62.200 171.595 ;
        RECT 58.475 170.965 59.725 171.135 ;
        RECT 58.475 170.845 58.805 170.965 ;
        RECT 57.135 170.455 59.035 170.625 ;
        RECT 56.775 170.115 58.695 170.285 ;
        RECT 56.775 170.095 57.095 170.115 ;
        RECT 56.325 169.435 56.655 169.945 ;
        RECT 56.925 169.485 57.095 170.095 ;
        RECT 58.865 169.945 59.035 170.455 ;
        RECT 59.205 170.385 59.385 170.795 ;
        RECT 59.555 170.205 59.725 170.965 ;
        RECT 57.265 169.225 57.595 169.915 ;
        RECT 57.825 169.775 59.035 169.945 ;
        RECT 59.205 169.895 59.725 170.205 ;
        RECT 59.895 170.795 60.315 171.135 ;
        RECT 60.605 170.795 61.015 171.125 ;
        RECT 59.895 170.025 60.085 170.795 ;
        RECT 61.185 170.665 61.355 171.395 ;
        RECT 62.500 171.225 62.670 171.555 ;
        RECT 62.840 171.395 63.170 171.775 ;
        RECT 61.525 170.845 61.875 171.215 ;
        RECT 61.185 170.625 61.605 170.665 ;
        RECT 60.255 170.455 61.605 170.625 ;
        RECT 60.255 170.295 60.505 170.455 ;
        RECT 61.015 170.025 61.265 170.285 ;
        RECT 59.895 169.775 61.265 170.025 ;
        RECT 57.825 169.485 58.065 169.775 ;
        RECT 58.865 169.695 59.035 169.775 ;
        RECT 58.265 169.225 58.685 169.605 ;
        RECT 58.865 169.445 59.495 169.695 ;
        RECT 59.965 169.225 60.295 169.605 ;
        RECT 60.465 169.485 60.635 169.775 ;
        RECT 61.435 169.610 61.605 170.455 ;
        RECT 62.055 170.285 62.275 171.155 ;
        RECT 62.500 171.035 63.195 171.225 ;
        RECT 61.775 169.905 62.275 170.285 ;
        RECT 62.445 170.235 62.855 170.855 ;
        RECT 63.025 170.065 63.195 171.035 ;
        RECT 62.500 169.895 63.195 170.065 ;
        RECT 60.815 169.225 61.195 169.605 ;
        RECT 61.435 169.440 62.265 169.610 ;
        RECT 62.500 169.395 62.670 169.895 ;
        RECT 62.840 169.225 63.170 169.725 ;
        RECT 63.385 169.395 63.610 171.515 ;
        RECT 63.780 171.395 64.110 171.775 ;
        RECT 64.280 171.225 64.450 171.515 ;
        RECT 63.785 171.055 64.450 171.225 ;
        RECT 63.785 170.065 64.015 171.055 ;
        RECT 65.630 171.005 69.140 171.775 ;
        RECT 64.185 170.235 64.535 170.885 ;
        RECT 65.630 170.315 67.320 170.835 ;
        RECT 67.490 170.485 69.140 171.005 ;
        RECT 69.585 170.965 69.830 171.570 ;
        RECT 70.050 171.240 70.560 171.775 ;
        RECT 69.310 170.795 70.540 170.965 ;
        RECT 63.785 169.895 64.450 170.065 ;
        RECT 63.780 169.225 64.110 169.725 ;
        RECT 64.280 169.395 64.450 169.895 ;
        RECT 65.630 169.225 69.140 170.315 ;
        RECT 69.310 169.985 69.650 170.795 ;
        RECT 69.820 170.230 70.570 170.420 ;
        RECT 69.310 169.575 69.825 169.985 ;
        RECT 70.060 169.225 70.230 169.985 ;
        RECT 70.400 169.565 70.570 170.230 ;
        RECT 70.740 170.245 70.930 171.605 ;
        RECT 71.100 170.755 71.375 171.605 ;
        RECT 71.565 171.240 72.095 171.605 ;
        RECT 72.520 171.375 72.850 171.775 ;
        RECT 71.920 171.205 72.095 171.240 ;
        RECT 71.100 170.585 71.380 170.755 ;
        RECT 71.100 170.445 71.375 170.585 ;
        RECT 71.580 170.245 71.750 171.045 ;
        RECT 70.740 170.075 71.750 170.245 ;
        RECT 71.920 171.035 72.850 171.205 ;
        RECT 73.020 171.035 73.275 171.605 ;
        RECT 73.450 171.050 73.740 171.775 ;
        RECT 71.920 169.905 72.090 171.035 ;
        RECT 72.680 170.865 72.850 171.035 ;
        RECT 70.965 169.735 72.090 169.905 ;
        RECT 72.260 170.535 72.455 170.865 ;
        RECT 72.680 170.535 72.935 170.865 ;
        RECT 72.260 169.565 72.430 170.535 ;
        RECT 73.105 170.365 73.275 171.035 ;
        RECT 73.950 170.955 74.180 171.775 ;
        RECT 74.350 170.975 74.680 171.605 ;
        RECT 73.930 170.535 74.260 170.785 ;
        RECT 70.400 169.395 72.430 169.565 ;
        RECT 72.600 169.225 72.770 170.365 ;
        RECT 72.940 169.395 73.275 170.365 ;
        RECT 73.450 169.225 73.740 170.390 ;
        RECT 74.430 170.375 74.680 170.975 ;
        RECT 74.850 170.955 75.060 171.775 ;
        RECT 75.750 171.005 77.420 171.775 ;
        RECT 73.950 169.225 74.180 170.365 ;
        RECT 74.350 169.395 74.680 170.375 ;
        RECT 74.850 169.225 75.060 170.365 ;
        RECT 75.750 170.315 76.500 170.835 ;
        RECT 76.670 170.485 77.420 171.005 ;
        RECT 77.595 170.935 77.855 171.775 ;
        RECT 78.030 171.030 78.285 171.605 ;
        RECT 78.455 171.395 78.785 171.775 ;
        RECT 79.000 171.225 79.170 171.605 ;
        RECT 79.805 171.435 80.060 171.595 ;
        RECT 79.720 171.265 80.060 171.435 ;
        RECT 80.240 171.315 80.525 171.775 ;
        RECT 78.455 171.055 79.170 171.225 ;
        RECT 79.805 171.065 80.060 171.265 ;
        RECT 75.750 169.225 77.420 170.315 ;
        RECT 77.595 169.225 77.855 170.375 ;
        RECT 78.030 170.300 78.200 171.030 ;
        RECT 78.455 170.865 78.625 171.055 ;
        RECT 78.370 170.535 78.625 170.865 ;
        RECT 78.455 170.325 78.625 170.535 ;
        RECT 78.905 170.505 79.260 170.875 ;
        RECT 78.030 169.395 78.285 170.300 ;
        RECT 78.455 170.155 79.170 170.325 ;
        RECT 78.455 169.225 78.785 169.985 ;
        RECT 79.000 169.395 79.170 170.155 ;
        RECT 79.805 170.205 79.985 171.065 ;
        RECT 80.705 170.865 80.955 171.515 ;
        RECT 80.155 170.535 80.955 170.865 ;
        RECT 79.805 169.535 80.060 170.205 ;
        RECT 80.240 169.225 80.525 170.025 ;
        RECT 80.705 169.945 80.955 170.535 ;
        RECT 81.155 171.180 81.475 171.510 ;
        RECT 81.655 171.295 82.315 171.775 ;
        RECT 82.515 171.385 83.365 171.555 ;
        RECT 81.155 170.285 81.345 171.180 ;
        RECT 81.665 170.855 82.325 171.125 ;
        RECT 81.995 170.795 82.325 170.855 ;
        RECT 81.515 170.625 81.845 170.685 ;
        RECT 82.515 170.625 82.685 171.385 ;
        RECT 83.925 171.315 84.245 171.775 ;
        RECT 84.445 171.135 84.695 171.565 ;
        RECT 84.985 171.335 85.395 171.775 ;
        RECT 85.565 171.395 86.580 171.595 ;
        RECT 82.855 170.965 84.105 171.135 ;
        RECT 82.855 170.845 83.185 170.965 ;
        RECT 81.515 170.455 83.415 170.625 ;
        RECT 81.155 170.115 83.075 170.285 ;
        RECT 81.155 170.095 81.475 170.115 ;
        RECT 80.705 169.435 81.035 169.945 ;
        RECT 81.305 169.485 81.475 170.095 ;
        RECT 83.245 169.945 83.415 170.455 ;
        RECT 83.585 170.385 83.765 170.795 ;
        RECT 83.935 170.205 84.105 170.965 ;
        RECT 81.645 169.225 81.975 169.915 ;
        RECT 82.205 169.775 83.415 169.945 ;
        RECT 83.585 169.895 84.105 170.205 ;
        RECT 84.275 170.795 84.695 171.135 ;
        RECT 84.985 170.795 85.395 171.125 ;
        RECT 84.275 170.025 84.465 170.795 ;
        RECT 85.565 170.665 85.735 171.395 ;
        RECT 86.880 171.225 87.050 171.555 ;
        RECT 87.220 171.395 87.550 171.775 ;
        RECT 85.905 170.845 86.255 171.215 ;
        RECT 85.565 170.625 85.985 170.665 ;
        RECT 84.635 170.455 85.985 170.625 ;
        RECT 84.635 170.295 84.885 170.455 ;
        RECT 85.395 170.025 85.645 170.285 ;
        RECT 84.275 169.775 85.645 170.025 ;
        RECT 82.205 169.485 82.445 169.775 ;
        RECT 83.245 169.695 83.415 169.775 ;
        RECT 82.645 169.225 83.065 169.605 ;
        RECT 83.245 169.445 83.875 169.695 ;
        RECT 84.345 169.225 84.675 169.605 ;
        RECT 84.845 169.485 85.015 169.775 ;
        RECT 85.815 169.610 85.985 170.455 ;
        RECT 86.435 170.285 86.655 171.155 ;
        RECT 86.880 171.035 87.575 171.225 ;
        RECT 86.155 169.905 86.655 170.285 ;
        RECT 86.825 170.235 87.235 170.855 ;
        RECT 87.405 170.065 87.575 171.035 ;
        RECT 86.880 169.895 87.575 170.065 ;
        RECT 85.195 169.225 85.575 169.605 ;
        RECT 85.815 169.440 86.645 169.610 ;
        RECT 86.880 169.395 87.050 169.895 ;
        RECT 87.220 169.225 87.550 169.725 ;
        RECT 87.765 169.395 87.990 171.515 ;
        RECT 88.160 171.395 88.490 171.775 ;
        RECT 88.660 171.225 88.830 171.515 ;
        RECT 88.165 171.055 88.830 171.225 ;
        RECT 89.205 171.145 89.490 171.605 ;
        RECT 89.660 171.315 89.930 171.775 ;
        RECT 88.165 170.065 88.395 171.055 ;
        RECT 89.205 170.975 90.160 171.145 ;
        RECT 88.565 170.235 88.915 170.885 ;
        RECT 89.090 170.245 89.780 170.805 ;
        RECT 89.950 170.075 90.160 170.975 ;
        RECT 88.165 169.895 88.830 170.065 ;
        RECT 88.160 169.225 88.490 169.725 ;
        RECT 88.660 169.395 88.830 169.895 ;
        RECT 89.205 169.855 90.160 170.075 ;
        RECT 90.330 170.805 90.730 171.605 ;
        RECT 90.920 171.145 91.200 171.605 ;
        RECT 91.720 171.315 92.045 171.775 ;
        RECT 90.920 170.975 92.045 171.145 ;
        RECT 92.215 171.035 92.600 171.605 ;
        RECT 91.595 170.865 92.045 170.975 ;
        RECT 90.330 170.245 91.425 170.805 ;
        RECT 91.595 170.535 92.150 170.865 ;
        RECT 89.205 169.395 89.490 169.855 ;
        RECT 89.660 169.225 89.930 169.685 ;
        RECT 90.330 169.395 90.730 170.245 ;
        RECT 91.595 170.075 92.045 170.535 ;
        RECT 92.320 170.365 92.600 171.035 ;
        RECT 93.805 171.145 94.090 171.605 ;
        RECT 94.260 171.315 94.530 171.775 ;
        RECT 93.805 170.975 94.760 171.145 ;
        RECT 90.920 169.855 92.045 170.075 ;
        RECT 90.920 169.395 91.200 169.855 ;
        RECT 91.720 169.225 92.045 169.685 ;
        RECT 92.215 169.395 92.600 170.365 ;
        RECT 93.690 170.245 94.380 170.805 ;
        RECT 94.550 170.075 94.760 170.975 ;
        RECT 93.805 169.855 94.760 170.075 ;
        RECT 94.930 170.805 95.330 171.605 ;
        RECT 95.520 171.145 95.800 171.605 ;
        RECT 96.320 171.315 96.645 171.775 ;
        RECT 95.520 170.975 96.645 171.145 ;
        RECT 96.815 171.035 97.200 171.605 ;
        RECT 96.195 170.865 96.645 170.975 ;
        RECT 94.930 170.245 96.025 170.805 ;
        RECT 96.195 170.535 96.750 170.865 ;
        RECT 93.805 169.395 94.090 169.855 ;
        RECT 94.260 169.225 94.530 169.685 ;
        RECT 94.930 169.395 95.330 170.245 ;
        RECT 96.195 170.075 96.645 170.535 ;
        RECT 96.920 170.365 97.200 171.035 ;
        RECT 97.370 171.005 99.040 171.775 ;
        RECT 99.210 171.050 99.500 171.775 ;
        RECT 99.670 171.025 100.880 171.775 ;
        RECT 95.520 169.855 96.645 170.075 ;
        RECT 95.520 169.395 95.800 169.855 ;
        RECT 96.320 169.225 96.645 169.685 ;
        RECT 96.815 169.395 97.200 170.365 ;
        RECT 97.370 170.315 98.120 170.835 ;
        RECT 98.290 170.485 99.040 171.005 ;
        RECT 97.370 169.225 99.040 170.315 ;
        RECT 99.210 169.225 99.500 170.390 ;
        RECT 99.670 170.315 100.190 170.855 ;
        RECT 100.360 170.485 100.880 171.025 ;
        RECT 101.050 171.005 104.560 171.775 ;
        RECT 101.050 170.315 102.740 170.835 ;
        RECT 102.910 170.485 104.560 171.005 ;
        RECT 104.790 170.955 105.000 171.775 ;
        RECT 105.170 170.975 105.500 171.605 ;
        RECT 105.170 170.375 105.420 170.975 ;
        RECT 105.670 170.955 105.900 171.775 ;
        RECT 106.110 171.025 107.320 171.775 ;
        RECT 105.590 170.535 105.920 170.785 ;
        RECT 99.670 169.225 100.880 170.315 ;
        RECT 101.050 169.225 104.560 170.315 ;
        RECT 104.790 169.225 105.000 170.365 ;
        RECT 105.170 169.395 105.500 170.375 ;
        RECT 105.670 169.225 105.900 170.365 ;
        RECT 106.110 170.315 106.630 170.855 ;
        RECT 106.800 170.485 107.320 171.025 ;
        RECT 107.490 171.005 111.000 171.775 ;
        RECT 111.170 171.025 112.380 171.775 ;
        RECT 107.490 170.315 109.180 170.835 ;
        RECT 109.350 170.485 111.000 171.005 ;
        RECT 111.170 170.315 111.690 170.855 ;
        RECT 111.860 170.485 112.380 171.025 ;
        RECT 106.110 169.225 107.320 170.315 ;
        RECT 107.490 169.225 111.000 170.315 ;
        RECT 111.170 169.225 112.380 170.315 ;
        RECT 18.165 169.055 112.465 169.225 ;
        RECT 18.250 167.965 19.460 169.055 ;
        RECT 19.940 168.215 20.110 169.055 ;
        RECT 20.320 168.045 20.570 168.885 ;
        RECT 20.780 168.215 20.950 169.055 ;
        RECT 21.120 168.045 21.410 168.885 ;
        RECT 18.250 167.255 18.770 167.795 ;
        RECT 18.940 167.425 19.460 167.965 ;
        RECT 19.685 167.875 21.410 168.045 ;
        RECT 21.620 167.995 21.790 169.055 ;
        RECT 22.085 168.675 22.415 169.055 ;
        RECT 22.595 168.505 22.765 168.795 ;
        RECT 22.935 168.595 23.185 169.055 ;
        RECT 21.965 168.335 22.765 168.505 ;
        RECT 23.355 168.545 24.225 168.885 ;
        RECT 19.685 167.325 20.095 167.875 ;
        RECT 21.965 167.715 22.135 168.335 ;
        RECT 23.355 168.165 23.525 168.545 ;
        RECT 24.460 168.425 24.630 168.885 ;
        RECT 24.800 168.595 25.170 169.055 ;
        RECT 25.465 168.455 25.635 168.795 ;
        RECT 25.805 168.625 26.135 169.055 ;
        RECT 26.370 168.455 26.540 168.795 ;
        RECT 22.305 167.995 23.525 168.165 ;
        RECT 23.695 168.085 24.155 168.375 ;
        RECT 24.460 168.255 25.020 168.425 ;
        RECT 25.465 168.285 26.540 168.455 ;
        RECT 26.710 168.555 27.390 168.885 ;
        RECT 27.605 168.555 27.855 168.885 ;
        RECT 28.025 168.595 28.275 169.055 ;
        RECT 24.850 168.115 25.020 168.255 ;
        RECT 23.695 168.075 24.660 168.085 ;
        RECT 23.355 167.905 23.525 167.995 ;
        RECT 23.985 167.915 24.660 168.075 ;
        RECT 21.965 167.705 22.310 167.715 ;
        RECT 20.280 167.495 22.310 167.705 ;
        RECT 18.250 166.505 19.460 167.255 ;
        RECT 19.685 167.155 21.450 167.325 ;
        RECT 19.940 166.505 20.110 166.975 ;
        RECT 20.280 166.675 20.610 167.155 ;
        RECT 20.780 166.505 20.950 166.975 ;
        RECT 21.120 166.675 21.450 167.155 ;
        RECT 21.620 166.505 21.790 167.315 ;
        RECT 21.985 167.240 22.310 167.495 ;
        RECT 21.990 166.885 22.310 167.240 ;
        RECT 22.480 167.455 23.020 167.825 ;
        RECT 23.355 167.735 23.760 167.905 ;
        RECT 22.480 167.055 22.720 167.455 ;
        RECT 23.200 167.285 23.420 167.565 ;
        RECT 22.890 167.115 23.420 167.285 ;
        RECT 22.890 166.885 23.060 167.115 ;
        RECT 23.590 166.955 23.760 167.735 ;
        RECT 23.930 167.125 24.280 167.745 ;
        RECT 24.450 167.125 24.660 167.915 ;
        RECT 24.850 167.945 26.350 168.115 ;
        RECT 24.850 167.255 25.020 167.945 ;
        RECT 26.710 167.775 26.880 168.555 ;
        RECT 27.685 168.425 27.855 168.555 ;
        RECT 25.190 167.605 26.880 167.775 ;
        RECT 27.050 167.995 27.515 168.385 ;
        RECT 27.685 168.255 28.080 168.425 ;
        RECT 25.190 167.425 25.360 167.605 ;
        RECT 21.990 166.715 23.060 166.885 ;
        RECT 23.230 166.505 23.420 166.945 ;
        RECT 23.590 166.675 24.540 166.955 ;
        RECT 24.850 166.865 25.110 167.255 ;
        RECT 25.530 167.185 26.320 167.435 ;
        RECT 24.760 166.695 25.110 166.865 ;
        RECT 25.320 166.505 25.650 166.965 ;
        RECT 26.525 166.895 26.695 167.605 ;
        RECT 27.050 167.405 27.220 167.995 ;
        RECT 26.865 167.185 27.220 167.405 ;
        RECT 27.390 167.185 27.740 167.805 ;
        RECT 27.910 166.895 28.080 168.255 ;
        RECT 28.445 168.085 28.770 168.870 ;
        RECT 28.250 167.035 28.710 168.085 ;
        RECT 26.525 166.725 27.380 166.895 ;
        RECT 27.585 166.725 28.080 166.895 ;
        RECT 28.250 166.505 28.580 166.865 ;
        RECT 28.940 166.765 29.110 168.885 ;
        RECT 29.280 168.555 29.610 169.055 ;
        RECT 29.780 168.385 30.035 168.885 ;
        RECT 29.285 168.215 30.035 168.385 ;
        RECT 30.670 168.295 31.185 168.705 ;
        RECT 31.420 168.295 31.590 169.055 ;
        RECT 31.760 168.715 33.790 168.885 ;
        RECT 29.285 167.225 29.515 168.215 ;
        RECT 29.685 167.395 30.035 168.045 ;
        RECT 30.670 167.485 31.010 168.295 ;
        RECT 31.760 168.050 31.930 168.715 ;
        RECT 32.325 168.375 33.450 168.545 ;
        RECT 31.180 167.860 31.930 168.050 ;
        RECT 32.100 168.035 33.110 168.205 ;
        RECT 30.670 167.315 31.900 167.485 ;
        RECT 29.285 167.055 30.035 167.225 ;
        RECT 29.280 166.505 29.610 166.885 ;
        RECT 29.780 166.765 30.035 167.055 ;
        RECT 30.945 166.710 31.190 167.315 ;
        RECT 31.410 166.505 31.920 167.040 ;
        RECT 32.100 166.675 32.290 168.035 ;
        RECT 32.460 167.015 32.735 167.835 ;
        RECT 32.940 167.235 33.110 168.035 ;
        RECT 33.280 167.245 33.450 168.375 ;
        RECT 33.620 167.745 33.790 168.715 ;
        RECT 33.960 167.915 34.130 169.055 ;
        RECT 34.300 167.915 34.635 168.885 ;
        RECT 33.620 167.415 33.815 167.745 ;
        RECT 34.040 167.415 34.295 167.745 ;
        RECT 34.040 167.245 34.210 167.415 ;
        RECT 34.465 167.245 34.635 167.915 ;
        RECT 34.810 167.890 35.100 169.055 ;
        RECT 35.270 168.335 35.730 168.885 ;
        RECT 35.920 168.335 36.250 169.055 ;
        RECT 33.280 167.075 34.210 167.245 ;
        RECT 33.280 167.040 33.455 167.075 ;
        RECT 32.460 166.845 32.740 167.015 ;
        RECT 32.460 166.675 32.735 166.845 ;
        RECT 32.925 166.675 33.455 167.040 ;
        RECT 33.880 166.505 34.210 166.905 ;
        RECT 34.380 166.675 34.635 167.245 ;
        RECT 34.810 166.505 35.100 167.230 ;
        RECT 35.270 166.965 35.520 168.335 ;
        RECT 36.450 168.165 36.750 168.715 ;
        RECT 36.920 168.385 37.200 169.055 ;
        RECT 37.685 168.425 37.970 168.885 ;
        RECT 38.140 168.595 38.410 169.055 ;
        RECT 37.685 168.205 38.640 168.425 ;
        RECT 35.810 167.995 36.750 168.165 ;
        RECT 35.810 167.745 35.980 167.995 ;
        RECT 37.120 167.745 37.385 168.105 ;
        RECT 35.690 167.415 35.980 167.745 ;
        RECT 36.150 167.495 36.490 167.745 ;
        RECT 36.710 167.495 37.385 167.745 ;
        RECT 37.570 167.475 38.260 168.035 ;
        RECT 35.810 167.325 35.980 167.415 ;
        RECT 35.810 167.135 37.200 167.325 ;
        RECT 38.430 167.305 38.640 168.205 ;
        RECT 35.270 166.675 35.830 166.965 ;
        RECT 36.000 166.505 36.250 166.965 ;
        RECT 36.870 166.775 37.200 167.135 ;
        RECT 37.685 167.135 38.640 167.305 ;
        RECT 38.810 168.035 39.210 168.885 ;
        RECT 39.400 168.425 39.680 168.885 ;
        RECT 40.200 168.595 40.525 169.055 ;
        RECT 39.400 168.205 40.525 168.425 ;
        RECT 38.810 167.475 39.905 168.035 ;
        RECT 40.075 167.745 40.525 168.205 ;
        RECT 40.695 167.915 41.080 168.885 ;
        RECT 37.685 166.675 37.970 167.135 ;
        RECT 38.140 166.505 38.410 166.965 ;
        RECT 38.810 166.675 39.210 167.475 ;
        RECT 40.075 167.415 40.630 167.745 ;
        RECT 40.075 167.305 40.525 167.415 ;
        RECT 39.400 167.135 40.525 167.305 ;
        RECT 40.800 167.245 41.080 167.915 ;
        RECT 41.250 168.295 41.765 168.705 ;
        RECT 42.000 168.295 42.170 169.055 ;
        RECT 42.340 168.715 44.370 168.885 ;
        RECT 41.250 167.485 41.590 168.295 ;
        RECT 42.340 168.050 42.510 168.715 ;
        RECT 42.905 168.375 44.030 168.545 ;
        RECT 41.760 167.860 42.510 168.050 ;
        RECT 42.680 168.035 43.690 168.205 ;
        RECT 41.250 167.315 42.480 167.485 ;
        RECT 39.400 166.675 39.680 167.135 ;
        RECT 40.200 166.505 40.525 166.965 ;
        RECT 40.695 166.675 41.080 167.245 ;
        RECT 41.525 166.710 41.770 167.315 ;
        RECT 41.990 166.505 42.500 167.040 ;
        RECT 42.680 166.675 42.870 168.035 ;
        RECT 43.040 167.695 43.315 167.835 ;
        RECT 43.040 167.525 43.320 167.695 ;
        RECT 43.040 166.675 43.315 167.525 ;
        RECT 43.520 167.235 43.690 168.035 ;
        RECT 43.860 167.245 44.030 168.375 ;
        RECT 44.200 167.745 44.370 168.715 ;
        RECT 44.540 167.915 44.710 169.055 ;
        RECT 44.880 167.915 45.215 168.885 ;
        RECT 45.450 167.915 45.660 169.055 ;
        RECT 44.200 167.415 44.395 167.745 ;
        RECT 44.620 167.415 44.875 167.745 ;
        RECT 44.620 167.245 44.790 167.415 ;
        RECT 45.045 167.245 45.215 167.915 ;
        RECT 45.830 167.905 46.160 168.885 ;
        RECT 46.330 167.915 46.560 169.055 ;
        RECT 46.780 168.245 47.075 169.055 ;
        RECT 43.860 167.075 44.790 167.245 ;
        RECT 43.860 167.040 44.035 167.075 ;
        RECT 43.505 166.675 44.035 167.040 ;
        RECT 44.460 166.505 44.790 166.905 ;
        RECT 44.960 166.675 45.215 167.245 ;
        RECT 45.450 166.505 45.660 167.325 ;
        RECT 45.830 167.305 46.080 167.905 ;
        RECT 47.255 167.745 47.500 168.885 ;
        RECT 47.675 168.245 47.935 169.055 ;
        RECT 48.535 169.050 54.810 169.055 ;
        RECT 48.115 167.745 48.365 168.880 ;
        RECT 48.535 168.255 48.795 169.050 ;
        RECT 48.965 168.155 49.225 168.880 ;
        RECT 49.395 168.325 49.655 169.050 ;
        RECT 49.825 168.155 50.085 168.880 ;
        RECT 50.255 168.325 50.515 169.050 ;
        RECT 50.685 168.155 50.945 168.880 ;
        RECT 51.115 168.325 51.375 169.050 ;
        RECT 51.545 168.155 51.805 168.880 ;
        RECT 51.975 168.325 52.220 169.050 ;
        RECT 52.390 168.155 52.650 168.880 ;
        RECT 52.835 168.325 53.080 169.050 ;
        RECT 53.250 168.155 53.510 168.880 ;
        RECT 53.695 168.325 53.940 169.050 ;
        RECT 54.110 168.155 54.370 168.880 ;
        RECT 54.555 168.325 54.810 169.050 ;
        RECT 48.965 168.140 54.370 168.155 ;
        RECT 54.980 168.140 55.270 168.880 ;
        RECT 55.440 168.310 55.710 169.055 ;
        RECT 48.965 167.915 55.710 168.140 ;
        RECT 46.250 167.495 46.580 167.745 ;
        RECT 45.830 166.675 46.160 167.305 ;
        RECT 46.330 166.505 46.560 167.325 ;
        RECT 46.770 167.185 47.085 167.745 ;
        RECT 47.255 167.495 54.375 167.745 ;
        RECT 46.770 166.505 47.075 167.015 ;
        RECT 47.255 166.685 47.505 167.495 ;
        RECT 47.675 166.505 47.935 167.030 ;
        RECT 48.115 166.685 48.365 167.495 ;
        RECT 54.545 167.355 55.710 167.915 ;
        RECT 55.975 167.915 56.310 168.885 ;
        RECT 56.480 167.915 56.650 169.055 ;
        RECT 56.820 168.715 58.850 168.885 ;
        RECT 54.545 167.325 55.740 167.355 ;
        RECT 48.965 167.185 55.740 167.325 ;
        RECT 55.975 167.245 56.145 167.915 ;
        RECT 56.820 167.745 56.990 168.715 ;
        RECT 56.315 167.415 56.570 167.745 ;
        RECT 56.795 167.415 56.990 167.745 ;
        RECT 57.160 168.375 58.285 168.545 ;
        RECT 56.400 167.245 56.570 167.415 ;
        RECT 57.160 167.245 57.330 168.375 ;
        RECT 48.965 167.155 55.710 167.185 ;
        RECT 48.535 166.505 48.795 167.065 ;
        RECT 48.965 166.700 49.225 167.155 ;
        RECT 49.395 166.505 49.655 166.985 ;
        RECT 49.825 166.700 50.085 167.155 ;
        RECT 50.255 166.505 50.515 166.985 ;
        RECT 50.685 166.700 50.945 167.155 ;
        RECT 51.115 166.505 51.360 166.985 ;
        RECT 51.530 166.700 51.805 167.155 ;
        RECT 51.975 166.505 52.220 166.985 ;
        RECT 52.390 166.700 52.650 167.155 ;
        RECT 52.830 166.505 53.080 166.985 ;
        RECT 53.250 166.700 53.510 167.155 ;
        RECT 53.690 166.505 53.940 166.985 ;
        RECT 54.110 166.700 54.370 167.155 ;
        RECT 54.550 166.505 54.810 166.985 ;
        RECT 54.980 166.700 55.240 167.155 ;
        RECT 55.410 166.505 55.710 166.985 ;
        RECT 55.975 166.675 56.230 167.245 ;
        RECT 56.400 167.075 57.330 167.245 ;
        RECT 57.500 168.035 58.510 168.205 ;
        RECT 57.500 167.235 57.670 168.035 ;
        RECT 57.875 167.695 58.150 167.835 ;
        RECT 57.870 167.525 58.150 167.695 ;
        RECT 57.155 167.040 57.330 167.075 ;
        RECT 56.400 166.505 56.730 166.905 ;
        RECT 57.155 166.675 57.685 167.040 ;
        RECT 57.875 166.675 58.150 167.525 ;
        RECT 58.320 166.675 58.510 168.035 ;
        RECT 58.680 168.050 58.850 168.715 ;
        RECT 59.020 168.295 59.190 169.055 ;
        RECT 59.425 168.295 59.940 168.705 ;
        RECT 58.680 167.860 59.430 168.050 ;
        RECT 59.600 167.485 59.940 168.295 ;
        RECT 60.570 167.890 60.860 169.055 ;
        RECT 61.090 167.915 61.300 169.055 ;
        RECT 61.470 167.905 61.800 168.885 ;
        RECT 61.970 167.915 62.200 169.055 ;
        RECT 62.410 167.965 64.080 169.055 ;
        RECT 58.710 167.315 59.940 167.485 ;
        RECT 58.690 166.505 59.200 167.040 ;
        RECT 59.420 166.710 59.665 167.315 ;
        RECT 60.570 166.505 60.860 167.230 ;
        RECT 61.090 166.505 61.300 167.325 ;
        RECT 61.470 167.305 61.720 167.905 ;
        RECT 61.890 167.495 62.220 167.745 ;
        RECT 62.410 167.445 63.160 167.965 ;
        RECT 64.310 167.915 64.520 169.055 ;
        RECT 64.690 167.905 65.020 168.885 ;
        RECT 65.190 167.915 65.420 169.055 ;
        RECT 65.630 168.295 66.145 168.705 ;
        RECT 66.380 168.295 66.550 169.055 ;
        RECT 66.720 168.715 68.750 168.885 ;
        RECT 61.470 166.675 61.800 167.305 ;
        RECT 61.970 166.505 62.200 167.325 ;
        RECT 63.330 167.275 64.080 167.795 ;
        RECT 62.410 166.505 64.080 167.275 ;
        RECT 64.310 166.505 64.520 167.325 ;
        RECT 64.690 167.305 64.940 167.905 ;
        RECT 65.110 167.495 65.440 167.745 ;
        RECT 65.630 167.485 65.970 168.295 ;
        RECT 66.720 168.050 66.890 168.715 ;
        RECT 67.285 168.375 68.410 168.545 ;
        RECT 66.140 167.860 66.890 168.050 ;
        RECT 67.060 168.035 68.070 168.205 ;
        RECT 64.690 166.675 65.020 167.305 ;
        RECT 65.190 166.505 65.420 167.325 ;
        RECT 65.630 167.315 66.860 167.485 ;
        RECT 65.905 166.710 66.150 167.315 ;
        RECT 66.370 166.505 66.880 167.040 ;
        RECT 67.060 166.675 67.250 168.035 ;
        RECT 67.420 167.695 67.695 167.835 ;
        RECT 67.420 167.525 67.700 167.695 ;
        RECT 67.420 166.675 67.695 167.525 ;
        RECT 67.900 167.235 68.070 168.035 ;
        RECT 68.240 167.245 68.410 168.375 ;
        RECT 68.580 167.745 68.750 168.715 ;
        RECT 68.920 167.915 69.090 169.055 ;
        RECT 69.260 167.915 69.595 168.885 ;
        RECT 69.860 168.385 70.030 168.885 ;
        RECT 70.200 168.555 70.530 169.055 ;
        RECT 69.860 168.215 70.525 168.385 ;
        RECT 68.580 167.415 68.775 167.745 ;
        RECT 69.000 167.415 69.255 167.745 ;
        RECT 69.000 167.245 69.170 167.415 ;
        RECT 69.425 167.245 69.595 167.915 ;
        RECT 69.775 167.395 70.125 168.045 ;
        RECT 68.240 167.075 69.170 167.245 ;
        RECT 68.240 167.040 68.415 167.075 ;
        RECT 67.885 166.675 68.415 167.040 ;
        RECT 68.840 166.505 69.170 166.905 ;
        RECT 69.340 166.675 69.595 167.245 ;
        RECT 70.295 167.225 70.525 168.215 ;
        RECT 69.860 167.055 70.525 167.225 ;
        RECT 69.860 166.765 70.030 167.055 ;
        RECT 70.200 166.505 70.530 166.885 ;
        RECT 70.700 166.765 70.925 168.885 ;
        RECT 71.140 168.555 71.470 169.055 ;
        RECT 71.640 168.385 71.810 168.885 ;
        RECT 72.045 168.670 72.875 168.840 ;
        RECT 73.115 168.675 73.495 169.055 ;
        RECT 71.115 168.215 71.810 168.385 ;
        RECT 71.115 167.245 71.285 168.215 ;
        RECT 71.455 167.425 71.865 168.045 ;
        RECT 72.035 167.995 72.535 168.375 ;
        RECT 71.115 167.055 71.810 167.245 ;
        RECT 72.035 167.125 72.255 167.995 ;
        RECT 72.705 167.825 72.875 168.670 ;
        RECT 73.675 168.505 73.845 168.795 ;
        RECT 74.015 168.675 74.345 169.055 ;
        RECT 74.815 168.585 75.445 168.835 ;
        RECT 75.625 168.675 76.045 169.055 ;
        RECT 75.275 168.505 75.445 168.585 ;
        RECT 76.245 168.505 76.485 168.795 ;
        RECT 73.045 168.255 74.415 168.505 ;
        RECT 73.045 167.995 73.295 168.255 ;
        RECT 73.805 167.825 74.055 167.985 ;
        RECT 72.705 167.655 74.055 167.825 ;
        RECT 72.705 167.615 73.125 167.655 ;
        RECT 72.435 167.065 72.785 167.435 ;
        RECT 71.140 166.505 71.470 166.885 ;
        RECT 71.640 166.725 71.810 167.055 ;
        RECT 72.955 166.885 73.125 167.615 ;
        RECT 74.225 167.485 74.415 168.255 ;
        RECT 73.295 167.155 73.705 167.485 ;
        RECT 73.995 167.145 74.415 167.485 ;
        RECT 74.585 168.075 75.105 168.385 ;
        RECT 75.275 168.335 76.485 168.505 ;
        RECT 76.715 168.365 77.045 169.055 ;
        RECT 74.585 167.315 74.755 168.075 ;
        RECT 74.925 167.485 75.105 167.895 ;
        RECT 75.275 167.825 75.445 168.335 ;
        RECT 77.215 168.185 77.385 168.795 ;
        RECT 77.655 168.335 77.985 168.845 ;
        RECT 77.215 168.165 77.535 168.185 ;
        RECT 75.615 167.995 77.535 168.165 ;
        RECT 75.275 167.655 77.175 167.825 ;
        RECT 75.505 167.315 75.835 167.435 ;
        RECT 74.585 167.145 75.835 167.315 ;
        RECT 72.110 166.685 73.125 166.885 ;
        RECT 73.295 166.505 73.705 166.945 ;
        RECT 73.995 166.715 74.245 167.145 ;
        RECT 74.445 166.505 74.765 166.965 ;
        RECT 76.005 166.895 76.175 167.655 ;
        RECT 76.845 167.595 77.175 167.655 ;
        RECT 76.365 167.425 76.695 167.485 ;
        RECT 76.365 167.155 77.025 167.425 ;
        RECT 77.345 167.100 77.535 167.995 ;
        RECT 75.325 166.725 76.175 166.895 ;
        RECT 76.375 166.505 77.035 166.985 ;
        RECT 77.215 166.770 77.535 167.100 ;
        RECT 77.735 167.745 77.985 168.335 ;
        RECT 78.165 168.255 78.450 169.055 ;
        RECT 78.630 168.715 78.885 168.745 ;
        RECT 78.630 168.545 78.970 168.715 ;
        RECT 78.630 168.075 78.885 168.545 ;
        RECT 80.090 168.385 80.370 169.055 ;
        RECT 80.540 168.165 80.840 168.715 ;
        RECT 81.040 168.335 81.370 169.055 ;
        RECT 81.560 168.335 82.020 168.885 ;
        RECT 77.735 167.415 78.535 167.745 ;
        RECT 77.735 166.765 77.985 167.415 ;
        RECT 78.705 167.215 78.885 168.075 ;
        RECT 79.905 167.745 80.170 168.105 ;
        RECT 80.540 167.995 81.480 168.165 ;
        RECT 81.310 167.745 81.480 167.995 ;
        RECT 79.905 167.495 80.580 167.745 ;
        RECT 80.800 167.495 81.140 167.745 ;
        RECT 81.310 167.415 81.600 167.745 ;
        RECT 81.310 167.325 81.480 167.415 ;
        RECT 78.165 166.505 78.450 166.965 ;
        RECT 78.630 166.685 78.885 167.215 ;
        RECT 80.090 167.135 81.480 167.325 ;
        RECT 80.090 166.775 80.420 167.135 ;
        RECT 81.770 166.965 82.020 168.335 ;
        RECT 82.190 168.295 82.705 168.705 ;
        RECT 82.940 168.295 83.110 169.055 ;
        RECT 83.280 168.715 85.310 168.885 ;
        RECT 82.190 167.485 82.530 168.295 ;
        RECT 83.280 168.050 83.450 168.715 ;
        RECT 83.845 168.375 84.970 168.545 ;
        RECT 82.700 167.860 83.450 168.050 ;
        RECT 83.620 168.035 84.630 168.205 ;
        RECT 82.190 167.315 83.420 167.485 ;
        RECT 81.040 166.505 81.290 166.965 ;
        RECT 81.460 166.675 82.020 166.965 ;
        RECT 82.465 166.710 82.710 167.315 ;
        RECT 82.930 166.505 83.440 167.040 ;
        RECT 83.620 166.675 83.810 168.035 ;
        RECT 83.980 167.695 84.255 167.835 ;
        RECT 83.980 167.525 84.260 167.695 ;
        RECT 83.980 166.675 84.255 167.525 ;
        RECT 84.460 167.235 84.630 168.035 ;
        RECT 84.800 167.245 84.970 168.375 ;
        RECT 85.140 167.745 85.310 168.715 ;
        RECT 85.480 167.915 85.650 169.055 ;
        RECT 85.820 167.915 86.155 168.885 ;
        RECT 85.140 167.415 85.335 167.745 ;
        RECT 85.560 167.415 85.815 167.745 ;
        RECT 85.560 167.245 85.730 167.415 ;
        RECT 85.985 167.245 86.155 167.915 ;
        RECT 86.330 167.890 86.620 169.055 ;
        RECT 86.790 167.915 87.060 168.885 ;
        RECT 87.270 168.255 87.550 169.055 ;
        RECT 87.720 168.545 89.375 168.835 ;
        RECT 87.785 168.205 89.375 168.375 ;
        RECT 87.785 168.085 87.955 168.205 ;
        RECT 87.230 167.915 87.955 168.085 ;
        RECT 84.800 167.075 85.730 167.245 ;
        RECT 84.800 167.040 84.975 167.075 ;
        RECT 84.445 166.675 84.975 167.040 ;
        RECT 85.400 166.505 85.730 166.905 ;
        RECT 85.900 166.675 86.155 167.245 ;
        RECT 86.330 166.505 86.620 167.230 ;
        RECT 86.790 167.180 86.960 167.915 ;
        RECT 87.230 167.745 87.400 167.915 ;
        RECT 88.145 167.865 88.860 168.035 ;
        RECT 89.055 167.915 89.375 168.205 ;
        RECT 89.550 167.915 89.890 168.885 ;
        RECT 90.060 167.915 90.230 169.055 ;
        RECT 90.500 168.255 90.750 169.055 ;
        RECT 91.395 168.085 91.725 168.885 ;
        RECT 92.025 168.255 92.355 169.055 ;
        RECT 92.525 168.085 92.855 168.885 ;
        RECT 90.420 167.915 92.855 168.085 ;
        RECT 93.230 168.295 93.745 168.705 ;
        RECT 93.980 168.295 94.150 169.055 ;
        RECT 94.320 168.715 96.350 168.885 ;
        RECT 87.130 167.415 87.400 167.745 ;
        RECT 87.570 167.415 87.975 167.745 ;
        RECT 88.145 167.415 88.855 167.865 ;
        RECT 87.230 167.245 87.400 167.415 ;
        RECT 86.790 166.835 87.060 167.180 ;
        RECT 87.230 167.075 88.840 167.245 ;
        RECT 89.025 167.175 89.375 167.745 ;
        RECT 89.550 167.355 89.725 167.915 ;
        RECT 90.420 167.665 90.590 167.915 ;
        RECT 89.895 167.495 90.590 167.665 ;
        RECT 90.765 167.495 91.185 167.695 ;
        RECT 91.355 167.495 91.685 167.695 ;
        RECT 91.855 167.495 92.185 167.695 ;
        RECT 89.550 167.305 89.780 167.355 ;
        RECT 87.250 166.505 87.630 166.905 ;
        RECT 87.800 166.725 87.970 167.075 ;
        RECT 88.140 166.505 88.470 166.905 ;
        RECT 88.670 166.725 88.840 167.075 ;
        RECT 89.040 166.505 89.370 167.005 ;
        RECT 89.550 166.675 89.890 167.305 ;
        RECT 90.060 166.505 90.310 167.305 ;
        RECT 90.500 167.155 91.725 167.325 ;
        RECT 90.500 166.675 90.830 167.155 ;
        RECT 91.000 166.505 91.225 166.965 ;
        RECT 91.395 166.675 91.725 167.155 ;
        RECT 92.355 167.285 92.525 167.915 ;
        RECT 92.710 167.495 93.060 167.745 ;
        RECT 93.230 167.485 93.570 168.295 ;
        RECT 94.320 168.050 94.490 168.715 ;
        RECT 94.885 168.375 96.010 168.545 ;
        RECT 93.740 167.860 94.490 168.050 ;
        RECT 94.660 168.035 95.670 168.205 ;
        RECT 93.230 167.315 94.460 167.485 ;
        RECT 92.355 166.675 92.855 167.285 ;
        RECT 93.505 166.710 93.750 167.315 ;
        RECT 93.970 166.505 94.480 167.040 ;
        RECT 94.660 166.675 94.850 168.035 ;
        RECT 95.020 167.695 95.295 167.835 ;
        RECT 95.020 167.525 95.300 167.695 ;
        RECT 95.020 166.675 95.295 167.525 ;
        RECT 95.500 167.235 95.670 168.035 ;
        RECT 95.840 167.245 96.010 168.375 ;
        RECT 96.180 167.745 96.350 168.715 ;
        RECT 96.520 167.915 96.690 169.055 ;
        RECT 96.860 167.915 97.195 168.885 ;
        RECT 96.180 167.415 96.375 167.745 ;
        RECT 96.600 167.415 96.855 167.745 ;
        RECT 96.600 167.245 96.770 167.415 ;
        RECT 97.025 167.245 97.195 167.915 ;
        RECT 97.370 167.965 99.960 169.055 ;
        RECT 100.130 168.295 100.645 168.705 ;
        RECT 100.880 168.295 101.050 169.055 ;
        RECT 101.220 168.715 103.250 168.885 ;
        RECT 97.370 167.445 98.580 167.965 ;
        RECT 98.750 167.275 99.960 167.795 ;
        RECT 100.130 167.485 100.470 168.295 ;
        RECT 101.220 168.050 101.390 168.715 ;
        RECT 101.785 168.375 102.910 168.545 ;
        RECT 100.640 167.860 101.390 168.050 ;
        RECT 101.560 168.035 102.570 168.205 ;
        RECT 100.130 167.315 101.360 167.485 ;
        RECT 95.840 167.075 96.770 167.245 ;
        RECT 95.840 167.040 96.015 167.075 ;
        RECT 95.485 166.675 96.015 167.040 ;
        RECT 96.440 166.505 96.770 166.905 ;
        RECT 96.940 166.675 97.195 167.245 ;
        RECT 97.370 166.505 99.960 167.275 ;
        RECT 100.405 166.710 100.650 167.315 ;
        RECT 100.870 166.505 101.380 167.040 ;
        RECT 101.560 166.675 101.750 168.035 ;
        RECT 101.920 167.695 102.195 167.835 ;
        RECT 101.920 167.525 102.200 167.695 ;
        RECT 101.920 166.675 102.195 167.525 ;
        RECT 102.400 167.235 102.570 168.035 ;
        RECT 102.740 167.245 102.910 168.375 ;
        RECT 103.080 167.745 103.250 168.715 ;
        RECT 103.420 167.915 103.590 169.055 ;
        RECT 103.760 167.915 104.095 168.885 ;
        RECT 104.790 167.915 105.000 169.055 ;
        RECT 103.080 167.415 103.275 167.745 ;
        RECT 103.500 167.415 103.755 167.745 ;
        RECT 103.500 167.245 103.670 167.415 ;
        RECT 103.925 167.245 104.095 167.915 ;
        RECT 105.170 167.905 105.500 168.885 ;
        RECT 105.670 167.915 105.900 169.055 ;
        RECT 106.110 167.965 107.320 169.055 ;
        RECT 107.490 167.965 111.000 169.055 ;
        RECT 111.170 167.965 112.380 169.055 ;
        RECT 102.740 167.075 103.670 167.245 ;
        RECT 102.740 167.040 102.915 167.075 ;
        RECT 102.385 166.675 102.915 167.040 ;
        RECT 103.340 166.505 103.670 166.905 ;
        RECT 103.840 166.675 104.095 167.245 ;
        RECT 104.790 166.505 105.000 167.325 ;
        RECT 105.170 167.305 105.420 167.905 ;
        RECT 105.590 167.495 105.920 167.745 ;
        RECT 106.110 167.425 106.630 167.965 ;
        RECT 105.170 166.675 105.500 167.305 ;
        RECT 105.670 166.505 105.900 167.325 ;
        RECT 106.800 167.255 107.320 167.795 ;
        RECT 107.490 167.445 109.180 167.965 ;
        RECT 109.350 167.275 111.000 167.795 ;
        RECT 111.170 167.425 111.690 167.965 ;
        RECT 106.110 166.505 107.320 167.255 ;
        RECT 107.490 166.505 111.000 167.275 ;
        RECT 111.860 167.255 112.380 167.795 ;
        RECT 111.170 166.505 112.380 167.255 ;
        RECT 18.165 166.335 112.465 166.505 ;
        RECT 18.250 165.585 19.460 166.335 ;
        RECT 20.090 165.835 20.350 166.165 ;
        RECT 20.560 165.855 20.835 166.335 ;
        RECT 18.250 165.045 18.770 165.585 ;
        RECT 18.940 164.875 19.460 165.415 ;
        RECT 18.250 163.785 19.460 164.875 ;
        RECT 20.090 164.925 20.260 165.835 ;
        RECT 21.045 165.765 21.250 166.165 ;
        RECT 21.420 165.935 21.755 166.335 ;
        RECT 20.430 165.095 20.790 165.675 ;
        RECT 21.045 165.595 21.730 165.765 ;
        RECT 21.930 165.610 22.220 166.335 ;
        RECT 22.940 165.785 23.110 166.165 ;
        RECT 23.325 165.955 23.655 166.335 ;
        RECT 22.940 165.615 23.655 165.785 ;
        RECT 20.970 164.925 21.220 165.425 ;
        RECT 20.090 164.755 21.220 164.925 ;
        RECT 20.090 163.985 20.360 164.755 ;
        RECT 21.390 164.565 21.730 165.595 ;
        RECT 22.850 165.065 23.205 165.435 ;
        RECT 23.485 165.425 23.655 165.615 ;
        RECT 23.825 165.590 24.080 166.165 ;
        RECT 23.485 165.095 23.740 165.425 ;
        RECT 20.530 163.785 20.860 164.565 ;
        RECT 21.065 164.390 21.730 164.565 ;
        RECT 21.065 163.985 21.250 164.390 ;
        RECT 21.420 163.785 21.755 164.210 ;
        RECT 21.930 163.785 22.220 164.950 ;
        RECT 23.485 164.885 23.655 165.095 ;
        RECT 22.940 164.715 23.655 164.885 ;
        RECT 23.910 164.860 24.080 165.590 ;
        RECT 24.255 165.495 24.515 166.335 ;
        RECT 24.690 165.835 24.990 166.165 ;
        RECT 25.160 165.855 25.435 166.335 ;
        RECT 22.940 163.955 23.110 164.715 ;
        RECT 23.325 163.785 23.655 164.545 ;
        RECT 23.825 163.955 24.080 164.860 ;
        RECT 24.255 163.785 24.515 164.935 ;
        RECT 24.690 164.925 24.860 165.835 ;
        RECT 25.615 165.685 25.910 166.075 ;
        RECT 26.080 165.855 26.335 166.335 ;
        RECT 26.510 165.685 26.770 166.075 ;
        RECT 26.940 165.855 27.220 166.335 ;
        RECT 25.030 165.095 25.380 165.665 ;
        RECT 25.615 165.515 27.265 165.685 ;
        RECT 25.550 165.175 26.690 165.345 ;
        RECT 25.550 164.925 25.720 165.175 ;
        RECT 26.860 165.005 27.265 165.515 ;
        RECT 24.690 164.755 25.720 164.925 ;
        RECT 26.510 164.835 27.265 165.005 ;
        RECT 27.450 165.660 27.720 166.005 ;
        RECT 27.910 165.935 28.290 166.335 ;
        RECT 28.460 165.765 28.630 166.115 ;
        RECT 28.800 165.935 29.130 166.335 ;
        RECT 29.330 165.765 29.500 166.115 ;
        RECT 29.700 165.835 30.030 166.335 ;
        RECT 27.450 164.925 27.620 165.660 ;
        RECT 27.890 165.595 29.500 165.765 ;
        RECT 27.890 165.425 28.060 165.595 ;
        RECT 27.790 165.095 28.060 165.425 ;
        RECT 28.230 165.095 28.635 165.425 ;
        RECT 27.890 164.925 28.060 165.095 ;
        RECT 28.805 164.975 29.515 165.425 ;
        RECT 29.685 165.095 30.035 165.665 ;
        RECT 30.210 165.595 30.595 166.165 ;
        RECT 30.765 165.875 31.090 166.335 ;
        RECT 31.610 165.705 31.890 166.165 ;
        RECT 24.690 163.955 25.000 164.755 ;
        RECT 26.510 164.585 26.770 164.835 ;
        RECT 25.170 163.785 25.480 164.585 ;
        RECT 25.650 164.415 26.770 164.585 ;
        RECT 25.650 163.955 25.910 164.415 ;
        RECT 26.080 163.785 26.335 164.245 ;
        RECT 26.510 163.955 26.770 164.415 ;
        RECT 26.940 163.785 27.225 164.655 ;
        RECT 27.450 163.955 27.720 164.925 ;
        RECT 27.890 164.755 28.615 164.925 ;
        RECT 28.805 164.805 29.520 164.975 ;
        RECT 30.210 164.925 30.490 165.595 ;
        RECT 30.765 165.535 31.890 165.705 ;
        RECT 30.765 165.425 31.215 165.535 ;
        RECT 30.660 165.095 31.215 165.425 ;
        RECT 32.080 165.365 32.480 166.165 ;
        RECT 32.880 165.875 33.150 166.335 ;
        RECT 33.320 165.705 33.605 166.165 ;
        RECT 28.445 164.635 28.615 164.755 ;
        RECT 29.715 164.635 30.035 164.925 ;
        RECT 27.930 163.785 28.210 164.585 ;
        RECT 28.445 164.465 30.035 164.635 ;
        RECT 28.380 164.005 30.035 164.295 ;
        RECT 30.210 163.955 30.595 164.925 ;
        RECT 30.765 164.635 31.215 165.095 ;
        RECT 31.385 164.805 32.480 165.365 ;
        RECT 30.765 164.415 31.890 164.635 ;
        RECT 30.765 163.785 31.090 164.245 ;
        RECT 31.610 163.955 31.890 164.415 ;
        RECT 32.080 163.955 32.480 164.805 ;
        RECT 32.650 165.535 33.605 165.705 ;
        RECT 33.890 165.535 34.230 166.165 ;
        RECT 34.400 165.535 34.650 166.335 ;
        RECT 34.840 165.685 35.170 166.165 ;
        RECT 35.340 165.875 35.565 166.335 ;
        RECT 35.735 165.685 36.065 166.165 ;
        RECT 32.650 164.635 32.860 165.535 ;
        RECT 33.890 165.485 34.120 165.535 ;
        RECT 34.840 165.515 36.065 165.685 ;
        RECT 36.695 165.555 37.195 166.165 ;
        RECT 37.945 165.995 38.200 166.155 ;
        RECT 37.860 165.825 38.200 165.995 ;
        RECT 38.380 165.875 38.665 166.335 ;
        RECT 37.945 165.625 38.200 165.825 ;
        RECT 33.030 164.805 33.720 165.365 ;
        RECT 33.890 164.925 34.065 165.485 ;
        RECT 34.235 165.175 34.930 165.345 ;
        RECT 34.760 164.925 34.930 165.175 ;
        RECT 35.105 165.145 35.525 165.345 ;
        RECT 35.695 165.145 36.025 165.345 ;
        RECT 36.195 165.145 36.525 165.345 ;
        RECT 36.695 164.925 36.865 165.555 ;
        RECT 37.050 165.095 37.400 165.345 ;
        RECT 32.650 164.415 33.605 164.635 ;
        RECT 32.880 163.785 33.150 164.245 ;
        RECT 33.320 163.955 33.605 164.415 ;
        RECT 33.890 163.955 34.230 164.925 ;
        RECT 34.400 163.785 34.570 164.925 ;
        RECT 34.760 164.755 37.195 164.925 ;
        RECT 34.840 163.785 35.090 164.585 ;
        RECT 35.735 163.955 36.065 164.755 ;
        RECT 36.365 163.785 36.695 164.585 ;
        RECT 36.865 163.955 37.195 164.755 ;
        RECT 37.945 164.765 38.125 165.625 ;
        RECT 38.845 165.425 39.095 166.075 ;
        RECT 38.295 165.095 39.095 165.425 ;
        RECT 37.945 164.095 38.200 164.765 ;
        RECT 38.380 163.785 38.665 164.585 ;
        RECT 38.845 164.505 39.095 165.095 ;
        RECT 39.295 165.740 39.615 166.070 ;
        RECT 39.795 165.855 40.455 166.335 ;
        RECT 40.655 165.945 41.505 166.115 ;
        RECT 39.295 164.845 39.485 165.740 ;
        RECT 39.805 165.415 40.465 165.685 ;
        RECT 40.135 165.355 40.465 165.415 ;
        RECT 39.655 165.185 39.985 165.245 ;
        RECT 40.655 165.185 40.825 165.945 ;
        RECT 42.065 165.875 42.385 166.335 ;
        RECT 42.585 165.695 42.835 166.125 ;
        RECT 43.125 165.895 43.535 166.335 ;
        RECT 43.705 165.955 44.720 166.155 ;
        RECT 40.995 165.525 42.245 165.695 ;
        RECT 40.995 165.405 41.325 165.525 ;
        RECT 39.655 165.015 41.555 165.185 ;
        RECT 39.295 164.675 41.215 164.845 ;
        RECT 39.295 164.655 39.615 164.675 ;
        RECT 38.845 163.995 39.175 164.505 ;
        RECT 39.445 164.045 39.615 164.655 ;
        RECT 41.385 164.505 41.555 165.015 ;
        RECT 41.725 164.945 41.905 165.355 ;
        RECT 42.075 164.765 42.245 165.525 ;
        RECT 39.785 163.785 40.115 164.475 ;
        RECT 40.345 164.335 41.555 164.505 ;
        RECT 41.725 164.455 42.245 164.765 ;
        RECT 42.415 165.355 42.835 165.695 ;
        RECT 43.125 165.355 43.535 165.685 ;
        RECT 42.415 164.585 42.605 165.355 ;
        RECT 43.705 165.225 43.875 165.955 ;
        RECT 45.020 165.785 45.190 166.115 ;
        RECT 45.360 165.955 45.690 166.335 ;
        RECT 44.045 165.405 44.395 165.775 ;
        RECT 43.705 165.185 44.125 165.225 ;
        RECT 42.775 165.015 44.125 165.185 ;
        RECT 42.775 164.855 43.025 165.015 ;
        RECT 43.535 164.585 43.785 164.845 ;
        RECT 42.415 164.335 43.785 164.585 ;
        RECT 40.345 164.045 40.585 164.335 ;
        RECT 41.385 164.255 41.555 164.335 ;
        RECT 40.785 163.785 41.205 164.165 ;
        RECT 41.385 164.005 42.015 164.255 ;
        RECT 42.485 163.785 42.815 164.165 ;
        RECT 42.985 164.045 43.155 164.335 ;
        RECT 43.955 164.170 44.125 165.015 ;
        RECT 44.575 164.845 44.795 165.715 ;
        RECT 45.020 165.595 45.715 165.785 ;
        RECT 44.295 164.465 44.795 164.845 ;
        RECT 44.965 164.795 45.375 165.415 ;
        RECT 45.545 164.625 45.715 165.595 ;
        RECT 45.020 164.455 45.715 164.625 ;
        RECT 43.335 163.785 43.715 164.165 ;
        RECT 43.955 164.000 44.785 164.170 ;
        RECT 45.020 163.955 45.190 164.455 ;
        RECT 45.360 163.785 45.690 164.285 ;
        RECT 45.905 163.955 46.130 166.075 ;
        RECT 46.300 165.955 46.630 166.335 ;
        RECT 46.800 165.785 46.970 166.075 ;
        RECT 46.305 165.615 46.970 165.785 ;
        RECT 46.305 164.625 46.535 165.615 ;
        RECT 47.690 165.610 47.980 166.335 ;
        RECT 48.190 165.515 48.420 166.335 ;
        RECT 48.590 165.535 48.920 166.165 ;
        RECT 46.705 164.795 47.055 165.445 ;
        RECT 48.170 165.095 48.500 165.345 ;
        RECT 46.305 164.455 46.970 164.625 ;
        RECT 46.300 163.785 46.630 164.285 ;
        RECT 46.800 163.955 46.970 164.455 ;
        RECT 47.690 163.785 47.980 164.950 ;
        RECT 48.670 164.935 48.920 165.535 ;
        RECT 49.090 165.515 49.300 166.335 ;
        RECT 49.905 165.995 50.160 166.155 ;
        RECT 49.820 165.825 50.160 165.995 ;
        RECT 50.340 165.875 50.625 166.335 ;
        RECT 49.905 165.625 50.160 165.825 ;
        RECT 48.190 163.785 48.420 164.925 ;
        RECT 48.590 163.955 48.920 164.935 ;
        RECT 49.090 163.785 49.300 164.925 ;
        RECT 49.905 164.765 50.085 165.625 ;
        RECT 50.805 165.425 51.055 166.075 ;
        RECT 50.255 165.095 51.055 165.425 ;
        RECT 49.905 164.095 50.160 164.765 ;
        RECT 50.340 163.785 50.625 164.585 ;
        RECT 50.805 164.505 51.055 165.095 ;
        RECT 51.255 165.740 51.575 166.070 ;
        RECT 51.755 165.855 52.415 166.335 ;
        RECT 52.615 165.945 53.465 166.115 ;
        RECT 51.255 164.845 51.445 165.740 ;
        RECT 51.765 165.415 52.425 165.685 ;
        RECT 52.095 165.355 52.425 165.415 ;
        RECT 51.615 165.185 51.945 165.245 ;
        RECT 52.615 165.185 52.785 165.945 ;
        RECT 54.025 165.875 54.345 166.335 ;
        RECT 54.545 165.695 54.795 166.125 ;
        RECT 55.085 165.895 55.495 166.335 ;
        RECT 55.665 165.955 56.680 166.155 ;
        RECT 52.955 165.525 54.205 165.695 ;
        RECT 52.955 165.405 53.285 165.525 ;
        RECT 51.615 165.015 53.515 165.185 ;
        RECT 51.255 164.675 53.175 164.845 ;
        RECT 51.255 164.655 51.575 164.675 ;
        RECT 50.805 163.995 51.135 164.505 ;
        RECT 51.405 164.045 51.575 164.655 ;
        RECT 53.345 164.505 53.515 165.015 ;
        RECT 53.685 164.945 53.865 165.355 ;
        RECT 54.035 164.765 54.205 165.525 ;
        RECT 51.745 163.785 52.075 164.475 ;
        RECT 52.305 164.335 53.515 164.505 ;
        RECT 53.685 164.455 54.205 164.765 ;
        RECT 54.375 165.355 54.795 165.695 ;
        RECT 55.085 165.355 55.495 165.685 ;
        RECT 54.375 164.585 54.565 165.355 ;
        RECT 55.665 165.225 55.835 165.955 ;
        RECT 56.980 165.785 57.150 166.115 ;
        RECT 57.320 165.955 57.650 166.335 ;
        RECT 56.005 165.405 56.355 165.775 ;
        RECT 55.665 165.185 56.085 165.225 ;
        RECT 54.735 165.015 56.085 165.185 ;
        RECT 54.735 164.855 54.985 165.015 ;
        RECT 55.495 164.585 55.745 164.845 ;
        RECT 54.375 164.335 55.745 164.585 ;
        RECT 52.305 164.045 52.545 164.335 ;
        RECT 53.345 164.255 53.515 164.335 ;
        RECT 52.745 163.785 53.165 164.165 ;
        RECT 53.345 164.005 53.975 164.255 ;
        RECT 54.445 163.785 54.775 164.165 ;
        RECT 54.945 164.045 55.115 164.335 ;
        RECT 55.915 164.170 56.085 165.015 ;
        RECT 56.535 164.845 56.755 165.715 ;
        RECT 56.980 165.595 57.675 165.785 ;
        RECT 56.255 164.465 56.755 164.845 ;
        RECT 56.925 164.795 57.335 165.415 ;
        RECT 57.505 164.625 57.675 165.595 ;
        RECT 56.980 164.455 57.675 164.625 ;
        RECT 55.295 163.785 55.675 164.165 ;
        RECT 55.915 164.000 56.745 164.170 ;
        RECT 56.980 163.955 57.150 164.455 ;
        RECT 57.320 163.785 57.650 164.285 ;
        RECT 57.865 163.955 58.090 166.075 ;
        RECT 58.260 165.955 58.590 166.335 ;
        RECT 58.760 165.785 58.930 166.075 ;
        RECT 58.265 165.615 58.930 165.785 ;
        RECT 58.265 164.625 58.495 165.615 ;
        RECT 59.190 165.585 60.400 166.335 ;
        RECT 58.665 164.795 59.015 165.445 ;
        RECT 59.190 164.875 59.710 165.415 ;
        RECT 59.880 165.045 60.400 165.585 ;
        RECT 60.685 165.705 60.970 166.165 ;
        RECT 61.140 165.875 61.410 166.335 ;
        RECT 60.685 165.535 61.640 165.705 ;
        RECT 58.265 164.455 58.930 164.625 ;
        RECT 58.260 163.785 58.590 164.285 ;
        RECT 58.760 163.955 58.930 164.455 ;
        RECT 59.190 163.785 60.400 164.875 ;
        RECT 60.570 164.805 61.260 165.365 ;
        RECT 61.430 164.635 61.640 165.535 ;
        RECT 60.685 164.415 61.640 164.635 ;
        RECT 61.810 165.365 62.210 166.165 ;
        RECT 62.400 165.705 62.680 166.165 ;
        RECT 63.200 165.875 63.525 166.335 ;
        RECT 62.400 165.535 63.525 165.705 ;
        RECT 63.695 165.595 64.080 166.165 ;
        RECT 63.075 165.425 63.525 165.535 ;
        RECT 61.810 164.805 62.905 165.365 ;
        RECT 63.075 165.095 63.630 165.425 ;
        RECT 60.685 163.955 60.970 164.415 ;
        RECT 61.140 163.785 61.410 164.245 ;
        RECT 61.810 163.955 62.210 164.805 ;
        RECT 63.075 164.635 63.525 165.095 ;
        RECT 63.800 164.925 64.080 165.595 ;
        RECT 62.400 164.415 63.525 164.635 ;
        RECT 62.400 163.955 62.680 164.415 ;
        RECT 63.200 163.785 63.525 164.245 ;
        RECT 63.695 163.955 64.080 164.925 ;
        RECT 64.255 165.625 64.510 166.155 ;
        RECT 64.680 165.875 64.985 166.335 ;
        RECT 65.230 165.955 66.300 166.125 ;
        RECT 64.255 164.975 64.465 165.625 ;
        RECT 65.230 165.600 65.550 165.955 ;
        RECT 65.225 165.425 65.550 165.600 ;
        RECT 64.635 165.125 65.550 165.425 ;
        RECT 65.720 165.385 65.960 165.785 ;
        RECT 66.130 165.725 66.300 165.955 ;
        RECT 66.470 165.895 66.660 166.335 ;
        RECT 66.830 165.885 67.780 166.165 ;
        RECT 68.000 165.975 68.350 166.145 ;
        RECT 66.130 165.555 66.660 165.725 ;
        RECT 64.635 165.095 65.375 165.125 ;
        RECT 64.255 164.095 64.510 164.975 ;
        RECT 64.680 163.785 64.985 164.925 ;
        RECT 65.205 164.505 65.375 165.095 ;
        RECT 65.720 165.015 66.260 165.385 ;
        RECT 66.440 165.275 66.660 165.555 ;
        RECT 66.830 165.105 67.000 165.885 ;
        RECT 66.595 164.935 67.000 165.105 ;
        RECT 67.170 165.095 67.520 165.715 ;
        RECT 66.595 164.845 66.765 164.935 ;
        RECT 67.690 164.925 67.900 165.715 ;
        RECT 65.545 164.675 66.765 164.845 ;
        RECT 67.225 164.765 67.900 164.925 ;
        RECT 65.205 164.335 66.005 164.505 ;
        RECT 65.325 163.785 65.655 164.165 ;
        RECT 65.835 164.045 66.005 164.335 ;
        RECT 66.595 164.295 66.765 164.675 ;
        RECT 66.935 164.755 67.900 164.765 ;
        RECT 68.090 165.585 68.350 165.975 ;
        RECT 68.560 165.875 68.890 166.335 ;
        RECT 69.765 165.945 70.620 166.115 ;
        RECT 70.825 165.945 71.320 166.115 ;
        RECT 71.490 165.975 71.820 166.335 ;
        RECT 68.090 164.895 68.260 165.585 ;
        RECT 68.430 165.235 68.600 165.415 ;
        RECT 68.770 165.405 69.560 165.655 ;
        RECT 69.765 165.235 69.935 165.945 ;
        RECT 70.105 165.435 70.460 165.655 ;
        RECT 68.430 165.065 70.120 165.235 ;
        RECT 66.935 164.465 67.395 164.755 ;
        RECT 68.090 164.725 69.590 164.895 ;
        RECT 68.090 164.585 68.260 164.725 ;
        RECT 67.700 164.415 68.260 164.585 ;
        RECT 66.175 163.785 66.425 164.245 ;
        RECT 66.595 163.955 67.465 164.295 ;
        RECT 67.700 163.955 67.870 164.415 ;
        RECT 68.705 164.385 69.780 164.555 ;
        RECT 68.040 163.785 68.410 164.245 ;
        RECT 68.705 164.045 68.875 164.385 ;
        RECT 69.045 163.785 69.375 164.215 ;
        RECT 69.610 164.045 69.780 164.385 ;
        RECT 69.950 164.285 70.120 165.065 ;
        RECT 70.290 164.845 70.460 165.435 ;
        RECT 70.630 165.035 70.980 165.655 ;
        RECT 70.290 164.455 70.755 164.845 ;
        RECT 71.150 164.585 71.320 165.945 ;
        RECT 71.490 164.755 71.950 165.805 ;
        RECT 70.925 164.415 71.320 164.585 ;
        RECT 70.925 164.285 71.095 164.415 ;
        RECT 69.950 163.955 70.630 164.285 ;
        RECT 70.845 163.955 71.095 164.285 ;
        RECT 71.265 163.785 71.515 164.245 ;
        RECT 71.685 163.970 72.010 164.755 ;
        RECT 72.180 163.955 72.350 166.075 ;
        RECT 72.520 165.955 72.850 166.335 ;
        RECT 73.020 165.785 73.275 166.075 ;
        RECT 72.525 165.615 73.275 165.785 ;
        RECT 72.525 164.625 72.755 165.615 ;
        RECT 73.450 165.610 73.740 166.335 ;
        RECT 74.870 165.515 75.100 166.335 ;
        RECT 75.270 165.535 75.600 166.165 ;
        RECT 72.925 164.795 73.275 165.445 ;
        RECT 74.850 165.095 75.180 165.345 ;
        RECT 72.525 164.455 73.275 164.625 ;
        RECT 72.520 163.785 72.850 164.285 ;
        RECT 73.020 163.955 73.275 164.455 ;
        RECT 73.450 163.785 73.740 164.950 ;
        RECT 75.350 164.935 75.600 165.535 ;
        RECT 75.770 165.515 75.980 166.335 ;
        RECT 76.270 165.855 76.550 166.335 ;
        RECT 76.720 165.685 76.980 166.075 ;
        RECT 77.155 165.855 77.410 166.335 ;
        RECT 77.580 165.685 77.875 166.075 ;
        RECT 78.055 165.855 78.330 166.335 ;
        RECT 78.500 165.835 78.800 166.165 ;
        RECT 76.225 165.515 77.875 165.685 ;
        RECT 74.870 163.785 75.100 164.925 ;
        RECT 75.270 163.955 75.600 164.935 ;
        RECT 76.225 165.005 76.630 165.515 ;
        RECT 76.800 165.175 77.940 165.345 ;
        RECT 75.770 163.785 75.980 164.925 ;
        RECT 76.225 164.835 76.980 165.005 ;
        RECT 76.265 163.785 76.550 164.655 ;
        RECT 76.720 164.585 76.980 164.835 ;
        RECT 77.770 164.925 77.940 165.175 ;
        RECT 78.110 165.095 78.460 165.665 ;
        RECT 78.630 164.925 78.800 165.835 ;
        RECT 77.770 164.755 78.800 164.925 ;
        RECT 76.720 164.415 77.840 164.585 ;
        RECT 76.720 163.955 76.980 164.415 ;
        RECT 77.155 163.785 77.410 164.245 ;
        RECT 77.580 163.955 77.840 164.415 ;
        RECT 78.010 163.785 78.320 164.585 ;
        RECT 78.490 163.955 78.800 164.755 ;
        RECT 79.345 165.625 79.600 166.155 ;
        RECT 79.780 165.875 80.065 166.335 ;
        RECT 79.345 164.765 79.525 165.625 ;
        RECT 80.245 165.425 80.495 166.075 ;
        RECT 79.695 165.095 80.495 165.425 ;
        RECT 79.345 164.295 79.600 164.765 ;
        RECT 79.260 164.125 79.600 164.295 ;
        RECT 79.345 164.095 79.600 164.125 ;
        RECT 79.780 163.785 80.065 164.585 ;
        RECT 80.245 164.505 80.495 165.095 ;
        RECT 80.695 165.740 81.015 166.070 ;
        RECT 81.195 165.855 81.855 166.335 ;
        RECT 82.055 165.945 82.905 166.115 ;
        RECT 80.695 164.845 80.885 165.740 ;
        RECT 81.205 165.415 81.865 165.685 ;
        RECT 81.535 165.355 81.865 165.415 ;
        RECT 81.055 165.185 81.385 165.245 ;
        RECT 82.055 165.185 82.225 165.945 ;
        RECT 83.465 165.875 83.785 166.335 ;
        RECT 83.985 165.695 84.235 166.125 ;
        RECT 84.525 165.895 84.935 166.335 ;
        RECT 85.105 165.955 86.120 166.155 ;
        RECT 82.395 165.525 83.645 165.695 ;
        RECT 82.395 165.405 82.725 165.525 ;
        RECT 81.055 165.015 82.955 165.185 ;
        RECT 80.695 164.675 82.615 164.845 ;
        RECT 80.695 164.655 81.015 164.675 ;
        RECT 80.245 163.995 80.575 164.505 ;
        RECT 80.845 164.045 81.015 164.655 ;
        RECT 82.785 164.505 82.955 165.015 ;
        RECT 83.125 164.945 83.305 165.355 ;
        RECT 83.475 164.765 83.645 165.525 ;
        RECT 81.185 163.785 81.515 164.475 ;
        RECT 81.745 164.335 82.955 164.505 ;
        RECT 83.125 164.455 83.645 164.765 ;
        RECT 83.815 165.355 84.235 165.695 ;
        RECT 84.525 165.355 84.935 165.685 ;
        RECT 83.815 164.585 84.005 165.355 ;
        RECT 85.105 165.225 85.275 165.955 ;
        RECT 86.420 165.785 86.590 166.115 ;
        RECT 86.760 165.955 87.090 166.335 ;
        RECT 85.445 165.405 85.795 165.775 ;
        RECT 85.105 165.185 85.525 165.225 ;
        RECT 84.175 165.015 85.525 165.185 ;
        RECT 84.175 164.855 84.425 165.015 ;
        RECT 84.935 164.585 85.185 164.845 ;
        RECT 83.815 164.335 85.185 164.585 ;
        RECT 81.745 164.045 81.985 164.335 ;
        RECT 82.785 164.255 82.955 164.335 ;
        RECT 82.185 163.785 82.605 164.165 ;
        RECT 82.785 164.005 83.415 164.255 ;
        RECT 83.885 163.785 84.215 164.165 ;
        RECT 84.385 164.045 84.555 164.335 ;
        RECT 85.355 164.170 85.525 165.015 ;
        RECT 85.975 164.845 86.195 165.715 ;
        RECT 86.420 165.595 87.115 165.785 ;
        RECT 85.695 164.465 86.195 164.845 ;
        RECT 86.365 164.795 86.775 165.415 ;
        RECT 86.945 164.625 87.115 165.595 ;
        RECT 86.420 164.455 87.115 164.625 ;
        RECT 84.735 163.785 85.115 164.165 ;
        RECT 85.355 164.000 86.185 164.170 ;
        RECT 86.420 163.955 86.590 164.455 ;
        RECT 86.760 163.785 87.090 164.285 ;
        RECT 87.305 163.955 87.530 166.075 ;
        RECT 87.700 165.955 88.030 166.335 ;
        RECT 88.200 165.785 88.370 166.075 ;
        RECT 87.705 165.615 88.370 165.785 ;
        RECT 87.705 164.625 87.935 165.615 ;
        RECT 88.690 165.515 88.900 166.335 ;
        RECT 89.070 165.535 89.400 166.165 ;
        RECT 88.105 164.795 88.455 165.445 ;
        RECT 89.070 164.935 89.320 165.535 ;
        RECT 89.570 165.515 89.800 166.335 ;
        RECT 90.015 165.625 90.270 166.155 ;
        RECT 90.440 165.875 90.745 166.335 ;
        RECT 90.990 165.955 92.060 166.125 ;
        RECT 89.490 165.095 89.820 165.345 ;
        RECT 90.015 164.975 90.225 165.625 ;
        RECT 90.990 165.600 91.310 165.955 ;
        RECT 90.985 165.425 91.310 165.600 ;
        RECT 90.395 165.125 91.310 165.425 ;
        RECT 91.480 165.385 91.720 165.785 ;
        RECT 91.890 165.725 92.060 165.955 ;
        RECT 92.230 165.895 92.420 166.335 ;
        RECT 92.590 165.885 93.540 166.165 ;
        RECT 93.760 165.975 94.110 166.145 ;
        RECT 91.890 165.555 92.420 165.725 ;
        RECT 90.395 165.095 91.135 165.125 ;
        RECT 87.705 164.455 88.370 164.625 ;
        RECT 87.700 163.785 88.030 164.285 ;
        RECT 88.200 163.955 88.370 164.455 ;
        RECT 88.690 163.785 88.900 164.925 ;
        RECT 89.070 163.955 89.400 164.935 ;
        RECT 89.570 163.785 89.800 164.925 ;
        RECT 90.015 164.095 90.270 164.975 ;
        RECT 90.440 163.785 90.745 164.925 ;
        RECT 90.965 164.505 91.135 165.095 ;
        RECT 91.480 165.015 92.020 165.385 ;
        RECT 92.200 165.275 92.420 165.555 ;
        RECT 92.590 165.105 92.760 165.885 ;
        RECT 92.355 164.935 92.760 165.105 ;
        RECT 92.930 165.095 93.280 165.715 ;
        RECT 92.355 164.845 92.525 164.935 ;
        RECT 93.450 164.925 93.660 165.715 ;
        RECT 91.305 164.675 92.525 164.845 ;
        RECT 92.985 164.765 93.660 164.925 ;
        RECT 90.965 164.335 91.765 164.505 ;
        RECT 91.085 163.785 91.415 164.165 ;
        RECT 91.595 164.045 91.765 164.335 ;
        RECT 92.355 164.295 92.525 164.675 ;
        RECT 92.695 164.755 93.660 164.765 ;
        RECT 93.850 165.585 94.110 165.975 ;
        RECT 94.320 165.875 94.650 166.335 ;
        RECT 95.525 165.945 96.380 166.115 ;
        RECT 96.585 165.945 97.080 166.115 ;
        RECT 97.250 165.975 97.580 166.335 ;
        RECT 93.850 164.895 94.020 165.585 ;
        RECT 94.190 165.235 94.360 165.415 ;
        RECT 94.530 165.405 95.320 165.655 ;
        RECT 95.525 165.235 95.695 165.945 ;
        RECT 95.865 165.435 96.220 165.655 ;
        RECT 94.190 165.065 95.880 165.235 ;
        RECT 92.695 164.465 93.155 164.755 ;
        RECT 93.850 164.725 95.350 164.895 ;
        RECT 93.850 164.585 94.020 164.725 ;
        RECT 93.460 164.415 94.020 164.585 ;
        RECT 91.935 163.785 92.185 164.245 ;
        RECT 92.355 163.955 93.225 164.295 ;
        RECT 93.460 163.955 93.630 164.415 ;
        RECT 94.465 164.385 95.540 164.555 ;
        RECT 93.800 163.785 94.170 164.245 ;
        RECT 94.465 164.045 94.635 164.385 ;
        RECT 94.805 163.785 95.135 164.215 ;
        RECT 95.370 164.045 95.540 164.385 ;
        RECT 95.710 164.285 95.880 165.065 ;
        RECT 96.050 164.845 96.220 165.435 ;
        RECT 96.390 165.035 96.740 165.655 ;
        RECT 96.050 164.455 96.515 164.845 ;
        RECT 96.910 164.585 97.080 165.945 ;
        RECT 97.250 164.755 97.710 165.805 ;
        RECT 96.685 164.415 97.080 164.585 ;
        RECT 96.685 164.285 96.855 164.415 ;
        RECT 95.710 163.955 96.390 164.285 ;
        RECT 96.605 163.955 96.855 164.285 ;
        RECT 97.025 163.785 97.275 164.245 ;
        RECT 97.445 163.970 97.770 164.755 ;
        RECT 97.940 163.955 98.110 166.075 ;
        RECT 98.280 165.955 98.610 166.335 ;
        RECT 98.780 165.785 99.035 166.075 ;
        RECT 98.285 165.615 99.035 165.785 ;
        RECT 98.285 164.625 98.515 165.615 ;
        RECT 99.210 165.610 99.500 166.335 ;
        RECT 99.670 165.585 100.880 166.335 ;
        RECT 101.425 165.655 101.680 166.155 ;
        RECT 101.860 165.875 102.145 166.335 ;
        RECT 98.685 164.795 99.035 165.445 ;
        RECT 98.285 164.455 99.035 164.625 ;
        RECT 98.280 163.785 98.610 164.285 ;
        RECT 98.780 163.955 99.035 164.455 ;
        RECT 99.210 163.785 99.500 164.950 ;
        RECT 99.670 164.875 100.190 165.415 ;
        RECT 100.360 165.045 100.880 165.585 ;
        RECT 101.340 165.625 101.680 165.655 ;
        RECT 101.340 165.485 101.605 165.625 ;
        RECT 99.670 163.785 100.880 164.875 ;
        RECT 101.425 164.765 101.605 165.485 ;
        RECT 102.325 165.425 102.575 166.075 ;
        RECT 101.775 165.095 102.575 165.425 ;
        RECT 101.425 164.095 101.680 164.765 ;
        RECT 101.860 163.785 102.145 164.585 ;
        RECT 102.325 164.505 102.575 165.095 ;
        RECT 102.775 165.740 103.095 166.070 ;
        RECT 103.275 165.855 103.935 166.335 ;
        RECT 104.135 165.945 104.985 166.115 ;
        RECT 102.775 164.845 102.965 165.740 ;
        RECT 103.285 165.415 103.945 165.685 ;
        RECT 103.615 165.355 103.945 165.415 ;
        RECT 103.135 165.185 103.465 165.245 ;
        RECT 104.135 165.185 104.305 165.945 ;
        RECT 105.545 165.875 105.865 166.335 ;
        RECT 106.065 165.695 106.315 166.125 ;
        RECT 106.605 165.895 107.015 166.335 ;
        RECT 107.185 165.955 108.200 166.155 ;
        RECT 104.475 165.525 105.725 165.695 ;
        RECT 104.475 165.405 104.805 165.525 ;
        RECT 103.135 165.015 105.035 165.185 ;
        RECT 102.775 164.675 104.695 164.845 ;
        RECT 102.775 164.655 103.095 164.675 ;
        RECT 102.325 163.995 102.655 164.505 ;
        RECT 102.925 164.045 103.095 164.655 ;
        RECT 104.865 164.505 105.035 165.015 ;
        RECT 105.205 164.945 105.385 165.355 ;
        RECT 105.555 164.765 105.725 165.525 ;
        RECT 103.265 163.785 103.595 164.475 ;
        RECT 103.825 164.335 105.035 164.505 ;
        RECT 105.205 164.455 105.725 164.765 ;
        RECT 105.895 165.355 106.315 165.695 ;
        RECT 106.605 165.355 107.015 165.685 ;
        RECT 105.895 164.585 106.085 165.355 ;
        RECT 107.185 165.225 107.355 165.955 ;
        RECT 108.500 165.785 108.670 166.115 ;
        RECT 108.840 165.955 109.170 166.335 ;
        RECT 107.525 165.405 107.875 165.775 ;
        RECT 107.185 165.185 107.605 165.225 ;
        RECT 106.255 165.015 107.605 165.185 ;
        RECT 106.255 164.855 106.505 165.015 ;
        RECT 107.015 164.585 107.265 164.845 ;
        RECT 105.895 164.335 107.265 164.585 ;
        RECT 103.825 164.045 104.065 164.335 ;
        RECT 104.865 164.255 105.035 164.335 ;
        RECT 104.265 163.785 104.685 164.165 ;
        RECT 104.865 164.005 105.495 164.255 ;
        RECT 105.965 163.785 106.295 164.165 ;
        RECT 106.465 164.045 106.635 164.335 ;
        RECT 107.435 164.170 107.605 165.015 ;
        RECT 108.055 164.845 108.275 165.715 ;
        RECT 108.500 165.595 109.195 165.785 ;
        RECT 107.775 164.465 108.275 164.845 ;
        RECT 108.445 164.795 108.855 165.415 ;
        RECT 109.025 164.625 109.195 165.595 ;
        RECT 108.500 164.455 109.195 164.625 ;
        RECT 106.815 163.785 107.195 164.165 ;
        RECT 107.435 164.000 108.265 164.170 ;
        RECT 108.500 163.955 108.670 164.455 ;
        RECT 108.840 163.785 109.170 164.285 ;
        RECT 109.385 163.955 109.610 166.075 ;
        RECT 109.780 165.955 110.110 166.335 ;
        RECT 110.280 165.785 110.450 166.075 ;
        RECT 109.785 165.615 110.450 165.785 ;
        RECT 109.785 164.625 110.015 165.615 ;
        RECT 111.170 165.585 112.380 166.335 ;
        RECT 110.185 164.795 110.535 165.445 ;
        RECT 111.170 164.875 111.690 165.415 ;
        RECT 111.860 165.045 112.380 165.585 ;
        RECT 109.785 164.455 110.450 164.625 ;
        RECT 109.780 163.785 110.110 164.285 ;
        RECT 110.280 163.955 110.450 164.455 ;
        RECT 111.170 163.785 112.380 164.875 ;
        RECT 18.165 163.615 112.465 163.785 ;
        RECT 18.250 162.525 19.460 163.615 ;
        RECT 18.250 161.815 18.770 162.355 ;
        RECT 18.940 161.985 19.460 162.525 ;
        RECT 20.095 162.465 20.355 163.615 ;
        RECT 20.530 162.540 20.785 163.445 ;
        RECT 20.955 162.855 21.285 163.615 ;
        RECT 21.500 162.685 21.670 163.445 ;
        RECT 22.045 162.985 22.330 163.445 ;
        RECT 22.500 163.155 22.770 163.615 ;
        RECT 22.045 162.765 23.000 162.985 ;
        RECT 18.250 161.065 19.460 161.815 ;
        RECT 20.095 161.065 20.355 161.905 ;
        RECT 20.530 161.810 20.700 162.540 ;
        RECT 20.955 162.515 21.670 162.685 ;
        RECT 20.955 162.305 21.125 162.515 ;
        RECT 20.870 161.975 21.125 162.305 ;
        RECT 20.530 161.235 20.785 161.810 ;
        RECT 20.955 161.785 21.125 161.975 ;
        RECT 21.405 161.965 21.760 162.335 ;
        RECT 21.930 162.035 22.620 162.595 ;
        RECT 22.790 161.865 23.000 162.765 ;
        RECT 20.955 161.615 21.670 161.785 ;
        RECT 20.955 161.065 21.285 161.445 ;
        RECT 21.500 161.235 21.670 161.615 ;
        RECT 22.045 161.695 23.000 161.865 ;
        RECT 23.170 162.595 23.570 163.445 ;
        RECT 23.760 162.985 24.040 163.445 ;
        RECT 24.560 163.155 24.885 163.615 ;
        RECT 23.760 162.765 24.885 162.985 ;
        RECT 23.170 162.035 24.265 162.595 ;
        RECT 24.435 162.305 24.885 162.765 ;
        RECT 25.055 162.475 25.440 163.445 ;
        RECT 22.045 161.235 22.330 161.695 ;
        RECT 22.500 161.065 22.770 161.525 ;
        RECT 23.170 161.235 23.570 162.035 ;
        RECT 24.435 161.975 24.990 162.305 ;
        RECT 24.435 161.865 24.885 161.975 ;
        RECT 23.760 161.695 24.885 161.865 ;
        RECT 25.160 161.805 25.440 162.475 ;
        RECT 23.760 161.235 24.040 161.695 ;
        RECT 24.560 161.065 24.885 161.525 ;
        RECT 25.055 161.235 25.440 161.805 ;
        RECT 25.615 162.425 25.870 163.305 ;
        RECT 26.040 162.475 26.345 163.615 ;
        RECT 26.685 163.235 27.015 163.615 ;
        RECT 27.195 163.065 27.365 163.355 ;
        RECT 27.535 163.155 27.785 163.615 ;
        RECT 26.565 162.895 27.365 163.065 ;
        RECT 27.955 163.105 28.825 163.445 ;
        RECT 25.615 161.775 25.825 162.425 ;
        RECT 26.565 162.305 26.735 162.895 ;
        RECT 27.955 162.725 28.125 163.105 ;
        RECT 29.060 162.985 29.230 163.445 ;
        RECT 29.400 163.155 29.770 163.615 ;
        RECT 30.065 163.015 30.235 163.355 ;
        RECT 30.405 163.185 30.735 163.615 ;
        RECT 30.970 163.015 31.140 163.355 ;
        RECT 26.905 162.555 28.125 162.725 ;
        RECT 28.295 162.645 28.755 162.935 ;
        RECT 29.060 162.815 29.620 162.985 ;
        RECT 30.065 162.845 31.140 163.015 ;
        RECT 31.310 163.115 31.990 163.445 ;
        RECT 32.205 163.115 32.455 163.445 ;
        RECT 32.625 163.155 32.875 163.615 ;
        RECT 29.450 162.675 29.620 162.815 ;
        RECT 28.295 162.635 29.260 162.645 ;
        RECT 27.955 162.465 28.125 162.555 ;
        RECT 28.585 162.475 29.260 162.635 ;
        RECT 25.995 162.275 26.735 162.305 ;
        RECT 25.995 161.975 26.910 162.275 ;
        RECT 26.585 161.800 26.910 161.975 ;
        RECT 25.615 161.245 25.870 161.775 ;
        RECT 26.040 161.065 26.345 161.525 ;
        RECT 26.590 161.445 26.910 161.800 ;
        RECT 27.080 162.015 27.620 162.385 ;
        RECT 27.955 162.295 28.360 162.465 ;
        RECT 27.080 161.615 27.320 162.015 ;
        RECT 27.800 161.845 28.020 162.125 ;
        RECT 27.490 161.675 28.020 161.845 ;
        RECT 27.490 161.445 27.660 161.675 ;
        RECT 28.190 161.515 28.360 162.295 ;
        RECT 28.530 161.685 28.880 162.305 ;
        RECT 29.050 161.685 29.260 162.475 ;
        RECT 29.450 162.505 30.950 162.675 ;
        RECT 29.450 161.815 29.620 162.505 ;
        RECT 31.310 162.335 31.480 163.115 ;
        RECT 32.285 162.985 32.455 163.115 ;
        RECT 29.790 162.165 31.480 162.335 ;
        RECT 31.650 162.555 32.115 162.945 ;
        RECT 32.285 162.815 32.680 162.985 ;
        RECT 29.790 161.985 29.960 162.165 ;
        RECT 26.590 161.275 27.660 161.445 ;
        RECT 27.830 161.065 28.020 161.505 ;
        RECT 28.190 161.235 29.140 161.515 ;
        RECT 29.450 161.425 29.710 161.815 ;
        RECT 30.130 161.745 30.920 161.995 ;
        RECT 29.360 161.255 29.710 161.425 ;
        RECT 29.920 161.065 30.250 161.525 ;
        RECT 31.125 161.455 31.295 162.165 ;
        RECT 31.650 161.965 31.820 162.555 ;
        RECT 31.465 161.745 31.820 161.965 ;
        RECT 31.990 161.745 32.340 162.365 ;
        RECT 32.510 161.455 32.680 162.815 ;
        RECT 33.045 162.645 33.370 163.430 ;
        RECT 32.850 161.595 33.310 162.645 ;
        RECT 31.125 161.285 31.980 161.455 ;
        RECT 32.185 161.285 32.680 161.455 ;
        RECT 32.850 161.065 33.180 161.425 ;
        RECT 33.540 161.325 33.710 163.445 ;
        RECT 33.880 163.115 34.210 163.615 ;
        RECT 34.380 162.945 34.635 163.445 ;
        RECT 33.885 162.775 34.635 162.945 ;
        RECT 33.885 161.785 34.115 162.775 ;
        RECT 34.285 161.955 34.635 162.605 ;
        RECT 34.810 162.450 35.100 163.615 ;
        RECT 35.360 162.870 35.630 163.615 ;
        RECT 36.260 163.610 42.535 163.615 ;
        RECT 35.800 162.700 36.090 163.440 ;
        RECT 36.260 162.885 36.515 163.610 ;
        RECT 36.700 162.715 36.960 163.440 ;
        RECT 37.130 162.885 37.375 163.610 ;
        RECT 37.560 162.715 37.820 163.440 ;
        RECT 37.990 162.885 38.235 163.610 ;
        RECT 38.420 162.715 38.680 163.440 ;
        RECT 38.850 162.885 39.095 163.610 ;
        RECT 39.265 162.715 39.525 163.440 ;
        RECT 39.695 162.885 39.955 163.610 ;
        RECT 40.125 162.715 40.385 163.440 ;
        RECT 40.555 162.885 40.815 163.610 ;
        RECT 40.985 162.715 41.245 163.440 ;
        RECT 41.415 162.885 41.675 163.610 ;
        RECT 41.845 162.715 42.105 163.440 ;
        RECT 42.275 162.815 42.535 163.610 ;
        RECT 36.700 162.700 42.105 162.715 ;
        RECT 35.360 162.475 42.105 162.700 ;
        RECT 35.360 161.885 36.525 162.475 ;
        RECT 42.705 162.305 42.955 163.440 ;
        RECT 43.135 162.805 43.395 163.615 ;
        RECT 43.570 162.305 43.815 163.445 ;
        RECT 43.995 162.805 44.290 163.615 ;
        RECT 45.045 162.985 45.330 163.445 ;
        RECT 45.500 163.155 45.770 163.615 ;
        RECT 45.045 162.765 46.000 162.985 ;
        RECT 36.695 162.055 43.815 162.305 ;
        RECT 33.885 161.615 34.635 161.785 ;
        RECT 33.880 161.065 34.210 161.445 ;
        RECT 34.380 161.325 34.635 161.615 ;
        RECT 34.810 161.065 35.100 161.790 ;
        RECT 35.360 161.715 42.105 161.885 ;
        RECT 35.360 161.065 35.660 161.545 ;
        RECT 35.830 161.260 36.090 161.715 ;
        RECT 36.260 161.065 36.520 161.545 ;
        RECT 36.700 161.260 36.960 161.715 ;
        RECT 37.130 161.065 37.380 161.545 ;
        RECT 37.560 161.260 37.820 161.715 ;
        RECT 37.990 161.065 38.240 161.545 ;
        RECT 38.420 161.260 38.680 161.715 ;
        RECT 38.850 161.065 39.095 161.545 ;
        RECT 39.265 161.260 39.540 161.715 ;
        RECT 39.710 161.065 39.955 161.545 ;
        RECT 40.125 161.260 40.385 161.715 ;
        RECT 40.555 161.065 40.815 161.545 ;
        RECT 40.985 161.260 41.245 161.715 ;
        RECT 41.415 161.065 41.675 161.545 ;
        RECT 41.845 161.260 42.105 161.715 ;
        RECT 42.275 161.065 42.535 161.625 ;
        RECT 42.705 161.245 42.955 162.055 ;
        RECT 43.135 161.065 43.395 161.590 ;
        RECT 43.565 161.245 43.815 162.055 ;
        RECT 43.985 161.745 44.300 162.305 ;
        RECT 44.930 162.035 45.620 162.595 ;
        RECT 45.790 161.865 46.000 162.765 ;
        RECT 45.045 161.695 46.000 161.865 ;
        RECT 46.170 162.595 46.570 163.445 ;
        RECT 46.760 162.985 47.040 163.445 ;
        RECT 47.560 163.155 47.885 163.615 ;
        RECT 46.760 162.765 47.885 162.985 ;
        RECT 46.170 162.035 47.265 162.595 ;
        RECT 47.435 162.305 47.885 162.765 ;
        RECT 48.055 162.475 48.440 163.445 ;
        RECT 48.725 162.985 49.010 163.445 ;
        RECT 49.180 163.155 49.450 163.615 ;
        RECT 48.725 162.765 49.680 162.985 ;
        RECT 43.995 161.065 44.300 161.575 ;
        RECT 45.045 161.235 45.330 161.695 ;
        RECT 45.500 161.065 45.770 161.525 ;
        RECT 46.170 161.235 46.570 162.035 ;
        RECT 47.435 161.975 47.990 162.305 ;
        RECT 47.435 161.865 47.885 161.975 ;
        RECT 46.760 161.695 47.885 161.865 ;
        RECT 48.160 161.805 48.440 162.475 ;
        RECT 48.610 162.035 49.300 162.595 ;
        RECT 49.470 161.865 49.680 162.765 ;
        RECT 46.760 161.235 47.040 161.695 ;
        RECT 47.560 161.065 47.885 161.525 ;
        RECT 48.055 161.235 48.440 161.805 ;
        RECT 48.725 161.695 49.680 161.865 ;
        RECT 49.850 162.595 50.250 163.445 ;
        RECT 50.440 162.985 50.720 163.445 ;
        RECT 51.240 163.155 51.565 163.615 ;
        RECT 50.440 162.765 51.565 162.985 ;
        RECT 49.850 162.035 50.945 162.595 ;
        RECT 51.115 162.305 51.565 162.765 ;
        RECT 51.735 162.475 52.120 163.445 ;
        RECT 48.725 161.235 49.010 161.695 ;
        RECT 49.180 161.065 49.450 161.525 ;
        RECT 49.850 161.235 50.250 162.035 ;
        RECT 51.115 161.975 51.670 162.305 ;
        RECT 51.115 161.865 51.565 161.975 ;
        RECT 50.440 161.695 51.565 161.865 ;
        RECT 51.840 161.805 52.120 162.475 ;
        RECT 52.290 162.855 52.805 163.265 ;
        RECT 53.040 162.855 53.210 163.615 ;
        RECT 53.380 163.275 55.410 163.445 ;
        RECT 52.290 162.045 52.630 162.855 ;
        RECT 53.380 162.610 53.550 163.275 ;
        RECT 53.945 162.935 55.070 163.105 ;
        RECT 52.800 162.420 53.550 162.610 ;
        RECT 53.720 162.595 54.730 162.765 ;
        RECT 52.290 161.875 53.520 162.045 ;
        RECT 50.440 161.235 50.720 161.695 ;
        RECT 51.240 161.065 51.565 161.525 ;
        RECT 51.735 161.235 52.120 161.805 ;
        RECT 52.565 161.270 52.810 161.875 ;
        RECT 53.030 161.065 53.540 161.600 ;
        RECT 53.720 161.235 53.910 162.595 ;
        RECT 54.080 162.255 54.355 162.395 ;
        RECT 54.080 162.085 54.360 162.255 ;
        RECT 54.080 161.235 54.355 162.085 ;
        RECT 54.560 161.795 54.730 162.595 ;
        RECT 54.900 161.805 55.070 162.935 ;
        RECT 55.240 162.305 55.410 163.275 ;
        RECT 55.580 162.475 55.750 163.615 ;
        RECT 55.920 162.475 56.255 163.445 ;
        RECT 55.240 161.975 55.435 162.305 ;
        RECT 55.660 161.975 55.915 162.305 ;
        RECT 55.660 161.805 55.830 161.975 ;
        RECT 56.085 161.805 56.255 162.475 ;
        RECT 56.560 162.445 56.890 163.615 ;
        RECT 57.090 162.275 57.420 163.445 ;
        RECT 57.620 162.445 57.950 163.615 ;
        RECT 58.150 162.275 58.510 163.445 ;
        RECT 58.680 162.475 59.010 163.615 ;
        RECT 59.230 162.475 59.460 163.615 ;
        RECT 59.630 162.465 59.960 163.445 ;
        RECT 60.130 162.475 60.340 163.615 ;
        RECT 57.090 161.995 58.510 162.275 ;
        RECT 54.900 161.635 55.830 161.805 ;
        RECT 54.900 161.600 55.075 161.635 ;
        RECT 54.545 161.235 55.075 161.600 ;
        RECT 55.500 161.065 55.830 161.465 ;
        RECT 56.000 161.235 56.255 161.805 ;
        RECT 57.100 161.065 57.430 161.755 ;
        RECT 58.150 161.660 58.510 161.995 ;
        RECT 58.680 161.725 59.020 162.305 ;
        RECT 59.210 162.055 59.540 162.305 ;
        RECT 57.890 161.235 58.510 161.660 ;
        RECT 58.680 161.065 59.010 161.555 ;
        RECT 59.230 161.065 59.460 161.885 ;
        RECT 59.710 161.865 59.960 162.465 ;
        RECT 60.570 162.450 60.860 163.615 ;
        RECT 61.490 162.855 62.005 163.265 ;
        RECT 62.240 162.855 62.410 163.615 ;
        RECT 62.580 163.275 64.610 163.445 ;
        RECT 61.490 162.045 61.830 162.855 ;
        RECT 62.580 162.610 62.750 163.275 ;
        RECT 63.145 162.935 64.270 163.105 ;
        RECT 62.000 162.420 62.750 162.610 ;
        RECT 62.920 162.595 63.930 162.765 ;
        RECT 59.630 161.235 59.960 161.865 ;
        RECT 60.130 161.065 60.340 161.885 ;
        RECT 61.490 161.875 62.720 162.045 ;
        RECT 60.570 161.065 60.860 161.790 ;
        RECT 61.765 161.270 62.010 161.875 ;
        RECT 62.230 161.065 62.740 161.600 ;
        RECT 62.920 161.235 63.110 162.595 ;
        RECT 63.280 161.575 63.555 162.395 ;
        RECT 63.760 161.795 63.930 162.595 ;
        RECT 64.100 161.805 64.270 162.935 ;
        RECT 64.440 162.305 64.610 163.275 ;
        RECT 64.780 162.475 64.950 163.615 ;
        RECT 65.120 162.475 65.455 163.445 ;
        RECT 64.440 161.975 64.635 162.305 ;
        RECT 64.860 161.975 65.115 162.305 ;
        RECT 64.860 161.805 65.030 161.975 ;
        RECT 65.285 161.805 65.455 162.475 ;
        RECT 65.630 162.525 66.840 163.615 ;
        RECT 67.125 162.985 67.410 163.445 ;
        RECT 67.580 163.155 67.850 163.615 ;
        RECT 67.125 162.765 68.080 162.985 ;
        RECT 65.630 161.985 66.150 162.525 ;
        RECT 66.320 161.815 66.840 162.355 ;
        RECT 67.010 162.035 67.700 162.595 ;
        RECT 67.870 161.865 68.080 162.765 ;
        RECT 64.100 161.635 65.030 161.805 ;
        RECT 64.100 161.600 64.275 161.635 ;
        RECT 63.280 161.405 63.560 161.575 ;
        RECT 63.280 161.235 63.555 161.405 ;
        RECT 63.745 161.235 64.275 161.600 ;
        RECT 64.700 161.065 65.030 161.465 ;
        RECT 65.200 161.235 65.455 161.805 ;
        RECT 65.630 161.065 66.840 161.815 ;
        RECT 67.125 161.695 68.080 161.865 ;
        RECT 68.250 162.595 68.650 163.445 ;
        RECT 68.840 162.985 69.120 163.445 ;
        RECT 69.640 163.155 69.965 163.615 ;
        RECT 68.840 162.765 69.965 162.985 ;
        RECT 68.250 162.035 69.345 162.595 ;
        RECT 69.515 162.305 69.965 162.765 ;
        RECT 70.135 162.475 70.520 163.445 ;
        RECT 71.240 162.870 71.510 163.615 ;
        RECT 72.140 163.610 78.415 163.615 ;
        RECT 71.680 162.700 71.970 163.440 ;
        RECT 72.140 162.885 72.395 163.610 ;
        RECT 72.580 162.715 72.840 163.440 ;
        RECT 73.010 162.885 73.255 163.610 ;
        RECT 73.440 162.715 73.700 163.440 ;
        RECT 73.870 162.885 74.115 163.610 ;
        RECT 74.300 162.715 74.560 163.440 ;
        RECT 74.730 162.885 74.975 163.610 ;
        RECT 75.145 162.715 75.405 163.440 ;
        RECT 75.575 162.885 75.835 163.610 ;
        RECT 76.005 162.715 76.265 163.440 ;
        RECT 76.435 162.885 76.695 163.610 ;
        RECT 76.865 162.715 77.125 163.440 ;
        RECT 77.295 162.885 77.555 163.610 ;
        RECT 77.725 162.715 77.985 163.440 ;
        RECT 78.155 162.815 78.415 163.610 ;
        RECT 72.580 162.700 77.985 162.715 ;
        RECT 67.125 161.235 67.410 161.695 ;
        RECT 67.580 161.065 67.850 161.525 ;
        RECT 68.250 161.235 68.650 162.035 ;
        RECT 69.515 161.975 70.070 162.305 ;
        RECT 69.515 161.865 69.965 161.975 ;
        RECT 68.840 161.695 69.965 161.865 ;
        RECT 70.240 161.805 70.520 162.475 ;
        RECT 68.840 161.235 69.120 161.695 ;
        RECT 69.640 161.065 69.965 161.525 ;
        RECT 70.135 161.235 70.520 161.805 ;
        RECT 71.240 162.475 77.985 162.700 ;
        RECT 71.240 161.885 72.405 162.475 ;
        RECT 78.585 162.305 78.835 163.440 ;
        RECT 79.015 162.805 79.275 163.615 ;
        RECT 79.450 162.305 79.695 163.445 ;
        RECT 79.875 162.805 80.170 163.615 ;
        RECT 80.355 162.475 80.690 163.445 ;
        RECT 80.860 162.475 81.030 163.615 ;
        RECT 81.200 163.275 83.230 163.445 ;
        RECT 72.575 162.055 79.695 162.305 ;
        RECT 71.240 161.715 77.985 161.885 ;
        RECT 71.240 161.065 71.540 161.545 ;
        RECT 71.710 161.260 71.970 161.715 ;
        RECT 72.140 161.065 72.400 161.545 ;
        RECT 72.580 161.260 72.840 161.715 ;
        RECT 73.010 161.065 73.260 161.545 ;
        RECT 73.440 161.260 73.700 161.715 ;
        RECT 73.870 161.065 74.120 161.545 ;
        RECT 74.300 161.260 74.560 161.715 ;
        RECT 74.730 161.065 74.975 161.545 ;
        RECT 75.145 161.260 75.420 161.715 ;
        RECT 75.590 161.065 75.835 161.545 ;
        RECT 76.005 161.260 76.265 161.715 ;
        RECT 76.435 161.065 76.695 161.545 ;
        RECT 76.865 161.260 77.125 161.715 ;
        RECT 77.295 161.065 77.555 161.545 ;
        RECT 77.725 161.260 77.985 161.715 ;
        RECT 78.155 161.065 78.415 161.625 ;
        RECT 78.585 161.245 78.835 162.055 ;
        RECT 79.015 161.065 79.275 161.590 ;
        RECT 79.445 161.245 79.695 162.055 ;
        RECT 79.865 161.745 80.180 162.305 ;
        RECT 80.355 161.805 80.525 162.475 ;
        RECT 81.200 162.305 81.370 163.275 ;
        RECT 80.695 161.975 80.950 162.305 ;
        RECT 81.175 161.975 81.370 162.305 ;
        RECT 81.540 162.935 82.665 163.105 ;
        RECT 80.780 161.805 80.950 161.975 ;
        RECT 81.540 161.805 81.710 162.935 ;
        RECT 79.875 161.065 80.180 161.575 ;
        RECT 80.355 161.235 80.610 161.805 ;
        RECT 80.780 161.635 81.710 161.805 ;
        RECT 81.880 162.595 82.890 162.765 ;
        RECT 81.880 161.795 82.050 162.595 ;
        RECT 81.535 161.600 81.710 161.635 ;
        RECT 80.780 161.065 81.110 161.465 ;
        RECT 81.535 161.235 82.065 161.600 ;
        RECT 82.255 161.575 82.530 162.395 ;
        RECT 82.250 161.405 82.530 161.575 ;
        RECT 82.255 161.235 82.530 161.405 ;
        RECT 82.700 161.235 82.890 162.595 ;
        RECT 83.060 162.610 83.230 163.275 ;
        RECT 83.400 162.855 83.570 163.615 ;
        RECT 83.805 162.855 84.320 163.265 ;
        RECT 83.060 162.420 83.810 162.610 ;
        RECT 83.980 162.045 84.320 162.855 ;
        RECT 84.550 162.780 84.805 163.615 ;
        RECT 84.975 162.610 85.235 163.415 ;
        RECT 85.405 162.780 85.665 163.615 ;
        RECT 85.835 162.610 86.090 163.415 ;
        RECT 83.090 161.875 84.320 162.045 ;
        RECT 84.490 162.440 86.090 162.610 ;
        RECT 86.330 162.450 86.620 163.615 ;
        RECT 86.800 162.805 87.095 163.615 ;
        RECT 84.490 161.875 84.770 162.440 ;
        RECT 87.275 162.305 87.520 163.445 ;
        RECT 87.695 162.805 87.955 163.615 ;
        RECT 88.555 163.610 94.830 163.615 ;
        RECT 88.135 162.305 88.385 163.440 ;
        RECT 88.555 162.815 88.815 163.610 ;
        RECT 88.985 162.715 89.245 163.440 ;
        RECT 89.415 162.885 89.675 163.610 ;
        RECT 89.845 162.715 90.105 163.440 ;
        RECT 90.275 162.885 90.535 163.610 ;
        RECT 90.705 162.715 90.965 163.440 ;
        RECT 91.135 162.885 91.395 163.610 ;
        RECT 91.565 162.715 91.825 163.440 ;
        RECT 91.995 162.885 92.240 163.610 ;
        RECT 92.410 162.715 92.670 163.440 ;
        RECT 92.855 162.885 93.100 163.610 ;
        RECT 93.270 162.715 93.530 163.440 ;
        RECT 93.715 162.885 93.960 163.610 ;
        RECT 94.130 162.715 94.390 163.440 ;
        RECT 94.575 162.885 94.830 163.610 ;
        RECT 88.985 162.700 94.390 162.715 ;
        RECT 95.000 162.700 95.290 163.440 ;
        RECT 95.460 162.870 95.730 163.615 ;
        RECT 95.990 162.855 96.505 163.265 ;
        RECT 96.740 162.855 96.910 163.615 ;
        RECT 97.080 163.275 99.110 163.445 ;
        RECT 88.985 162.475 95.730 162.700 ;
        RECT 84.940 162.045 86.160 162.270 ;
        RECT 83.070 161.065 83.580 161.600 ;
        RECT 83.800 161.270 84.045 161.875 ;
        RECT 84.490 161.705 85.220 161.875 ;
        RECT 84.495 161.065 84.825 161.535 ;
        RECT 84.995 161.260 85.220 161.705 ;
        RECT 85.390 161.065 85.685 161.590 ;
        RECT 86.330 161.065 86.620 161.790 ;
        RECT 86.790 161.745 87.105 162.305 ;
        RECT 87.275 162.055 94.395 162.305 ;
        RECT 94.565 162.255 95.730 162.475 ;
        RECT 94.565 162.085 95.760 162.255 ;
        RECT 86.790 161.065 87.095 161.575 ;
        RECT 87.275 161.245 87.525 162.055 ;
        RECT 87.695 161.065 87.955 161.590 ;
        RECT 88.135 161.245 88.385 162.055 ;
        RECT 94.565 161.885 95.730 162.085 ;
        RECT 88.985 161.715 95.730 161.885 ;
        RECT 95.990 162.045 96.330 162.855 ;
        RECT 97.080 162.610 97.250 163.275 ;
        RECT 97.645 162.935 98.770 163.105 ;
        RECT 96.500 162.420 97.250 162.610 ;
        RECT 97.420 162.595 98.430 162.765 ;
        RECT 95.990 161.875 97.220 162.045 ;
        RECT 88.555 161.065 88.815 161.625 ;
        RECT 88.985 161.260 89.245 161.715 ;
        RECT 89.415 161.065 89.675 161.545 ;
        RECT 89.845 161.260 90.105 161.715 ;
        RECT 90.275 161.065 90.535 161.545 ;
        RECT 90.705 161.260 90.965 161.715 ;
        RECT 91.135 161.065 91.380 161.545 ;
        RECT 91.550 161.260 91.825 161.715 ;
        RECT 91.995 161.065 92.240 161.545 ;
        RECT 92.410 161.260 92.670 161.715 ;
        RECT 92.850 161.065 93.100 161.545 ;
        RECT 93.270 161.260 93.530 161.715 ;
        RECT 93.710 161.065 93.960 161.545 ;
        RECT 94.130 161.260 94.390 161.715 ;
        RECT 94.570 161.065 94.830 161.545 ;
        RECT 95.000 161.260 95.260 161.715 ;
        RECT 95.430 161.065 95.730 161.545 ;
        RECT 96.265 161.270 96.510 161.875 ;
        RECT 96.730 161.065 97.240 161.600 ;
        RECT 97.420 161.235 97.610 162.595 ;
        RECT 97.780 161.915 98.055 162.395 ;
        RECT 97.780 161.745 98.060 161.915 ;
        RECT 98.260 161.795 98.430 162.595 ;
        RECT 98.600 161.805 98.770 162.935 ;
        RECT 98.940 162.305 99.110 163.275 ;
        RECT 99.280 162.475 99.450 163.615 ;
        RECT 99.620 162.475 99.955 163.445 ;
        RECT 98.940 161.975 99.135 162.305 ;
        RECT 99.360 161.975 99.615 162.305 ;
        RECT 99.360 161.805 99.530 161.975 ;
        RECT 99.785 161.805 99.955 162.475 ;
        RECT 97.780 161.235 98.055 161.745 ;
        RECT 98.600 161.635 99.530 161.805 ;
        RECT 98.600 161.600 98.775 161.635 ;
        RECT 98.245 161.235 98.775 161.600 ;
        RECT 99.200 161.065 99.530 161.465 ;
        RECT 99.700 161.235 99.955 161.805 ;
        RECT 100.505 162.635 100.760 163.305 ;
        RECT 100.940 162.815 101.225 163.615 ;
        RECT 101.405 162.895 101.735 163.405 ;
        RECT 100.505 161.775 100.685 162.635 ;
        RECT 101.405 162.305 101.655 162.895 ;
        RECT 102.005 162.745 102.175 163.355 ;
        RECT 102.345 162.925 102.675 163.615 ;
        RECT 102.905 163.065 103.145 163.355 ;
        RECT 103.345 163.235 103.765 163.615 ;
        RECT 103.945 163.145 104.575 163.395 ;
        RECT 105.045 163.235 105.375 163.615 ;
        RECT 103.945 163.065 104.115 163.145 ;
        RECT 105.545 163.065 105.715 163.355 ;
        RECT 105.895 163.235 106.275 163.615 ;
        RECT 106.515 163.230 107.345 163.400 ;
        RECT 102.905 162.895 104.115 163.065 ;
        RECT 100.855 161.975 101.655 162.305 ;
        RECT 100.505 161.575 100.760 161.775 ;
        RECT 100.420 161.405 100.760 161.575 ;
        RECT 100.505 161.245 100.760 161.405 ;
        RECT 100.940 161.065 101.225 161.525 ;
        RECT 101.405 161.325 101.655 161.975 ;
        RECT 101.855 162.725 102.175 162.745 ;
        RECT 101.855 162.555 103.775 162.725 ;
        RECT 101.855 161.660 102.045 162.555 ;
        RECT 103.945 162.385 104.115 162.895 ;
        RECT 104.285 162.635 104.805 162.945 ;
        RECT 102.215 162.215 104.115 162.385 ;
        RECT 102.215 162.155 102.545 162.215 ;
        RECT 102.695 161.985 103.025 162.045 ;
        RECT 102.365 161.715 103.025 161.985 ;
        RECT 101.855 161.330 102.175 161.660 ;
        RECT 102.355 161.065 103.015 161.545 ;
        RECT 103.215 161.455 103.385 162.215 ;
        RECT 104.285 162.045 104.465 162.455 ;
        RECT 103.555 161.875 103.885 161.995 ;
        RECT 104.635 161.875 104.805 162.635 ;
        RECT 103.555 161.705 104.805 161.875 ;
        RECT 104.975 162.815 106.345 163.065 ;
        RECT 104.975 162.045 105.165 162.815 ;
        RECT 106.095 162.555 106.345 162.815 ;
        RECT 105.335 162.385 105.585 162.545 ;
        RECT 106.515 162.385 106.685 163.230 ;
        RECT 107.580 162.945 107.750 163.445 ;
        RECT 107.920 163.115 108.250 163.615 ;
        RECT 106.855 162.555 107.355 162.935 ;
        RECT 107.580 162.775 108.275 162.945 ;
        RECT 105.335 162.215 106.685 162.385 ;
        RECT 106.265 162.175 106.685 162.215 ;
        RECT 104.975 161.705 105.395 162.045 ;
        RECT 105.685 161.715 106.095 162.045 ;
        RECT 103.215 161.285 104.065 161.455 ;
        RECT 104.625 161.065 104.945 161.525 ;
        RECT 105.145 161.275 105.395 161.705 ;
        RECT 105.685 161.065 106.095 161.505 ;
        RECT 106.265 161.445 106.435 162.175 ;
        RECT 106.605 161.625 106.955 161.995 ;
        RECT 107.135 161.685 107.355 162.555 ;
        RECT 107.525 161.985 107.935 162.605 ;
        RECT 108.105 161.805 108.275 162.775 ;
        RECT 107.580 161.615 108.275 161.805 ;
        RECT 106.265 161.245 107.280 161.445 ;
        RECT 107.580 161.285 107.750 161.615 ;
        RECT 107.920 161.065 108.250 161.445 ;
        RECT 108.465 161.325 108.690 163.445 ;
        RECT 108.860 163.115 109.190 163.615 ;
        RECT 109.360 162.945 109.530 163.445 ;
        RECT 108.865 162.775 109.530 162.945 ;
        RECT 108.865 161.785 109.095 162.775 ;
        RECT 109.265 161.955 109.615 162.605 ;
        RECT 109.790 162.525 111.000 163.615 ;
        RECT 111.170 162.525 112.380 163.615 ;
        RECT 109.790 161.985 110.310 162.525 ;
        RECT 110.480 161.815 111.000 162.355 ;
        RECT 111.170 161.985 111.690 162.525 ;
        RECT 111.860 161.815 112.380 162.355 ;
        RECT 108.865 161.615 109.530 161.785 ;
        RECT 108.860 161.065 109.190 161.445 ;
        RECT 109.360 161.325 109.530 161.615 ;
        RECT 109.790 161.065 111.000 161.815 ;
        RECT 111.170 161.065 112.380 161.815 ;
        RECT 18.165 160.895 112.465 161.065 ;
        RECT 18.250 160.145 19.460 160.895 ;
        RECT 18.250 159.605 18.770 160.145 ;
        RECT 20.610 160.075 20.820 160.895 ;
        RECT 20.990 160.095 21.320 160.725 ;
        RECT 18.940 159.435 19.460 159.975 ;
        RECT 20.990 159.495 21.240 160.095 ;
        RECT 21.490 160.075 21.720 160.895 ;
        RECT 21.930 160.170 22.220 160.895 ;
        RECT 22.700 160.425 22.870 160.895 ;
        RECT 23.040 160.245 23.370 160.725 ;
        RECT 23.540 160.425 23.710 160.895 ;
        RECT 23.880 160.245 24.210 160.725 ;
        RECT 22.445 160.075 24.210 160.245 ;
        RECT 24.380 160.085 24.550 160.895 ;
        RECT 24.750 160.515 25.820 160.685 ;
        RECT 24.750 160.160 25.070 160.515 ;
        RECT 21.410 159.655 21.740 159.905 ;
        RECT 22.445 159.525 22.855 160.075 ;
        RECT 24.745 159.905 25.070 160.160 ;
        RECT 23.040 159.695 25.070 159.905 ;
        RECT 24.725 159.685 25.070 159.695 ;
        RECT 25.240 159.945 25.480 160.345 ;
        RECT 25.650 160.285 25.820 160.515 ;
        RECT 25.990 160.455 26.180 160.895 ;
        RECT 26.350 160.445 27.300 160.725 ;
        RECT 27.520 160.535 27.870 160.705 ;
        RECT 25.650 160.115 26.180 160.285 ;
        RECT 18.250 158.345 19.460 159.435 ;
        RECT 20.610 158.345 20.820 159.485 ;
        RECT 20.990 158.515 21.320 159.495 ;
        RECT 21.490 158.345 21.720 159.485 ;
        RECT 21.930 158.345 22.220 159.510 ;
        RECT 22.445 159.355 24.170 159.525 ;
        RECT 22.700 158.345 22.870 159.185 ;
        RECT 23.080 158.515 23.330 159.355 ;
        RECT 23.540 158.345 23.710 159.185 ;
        RECT 23.880 158.515 24.170 159.355 ;
        RECT 24.380 158.345 24.550 159.405 ;
        RECT 24.725 159.065 24.895 159.685 ;
        RECT 25.240 159.575 25.780 159.945 ;
        RECT 25.960 159.835 26.180 160.115 ;
        RECT 26.350 159.665 26.520 160.445 ;
        RECT 26.115 159.495 26.520 159.665 ;
        RECT 26.690 159.655 27.040 160.275 ;
        RECT 26.115 159.405 26.285 159.495 ;
        RECT 27.210 159.485 27.420 160.275 ;
        RECT 25.065 159.235 26.285 159.405 ;
        RECT 26.745 159.325 27.420 159.485 ;
        RECT 24.725 158.895 25.525 159.065 ;
        RECT 24.845 158.345 25.175 158.725 ;
        RECT 25.355 158.605 25.525 158.895 ;
        RECT 26.115 158.855 26.285 159.235 ;
        RECT 26.455 159.315 27.420 159.325 ;
        RECT 27.610 160.145 27.870 160.535 ;
        RECT 28.080 160.435 28.410 160.895 ;
        RECT 29.285 160.505 30.140 160.675 ;
        RECT 30.345 160.505 30.840 160.675 ;
        RECT 31.010 160.535 31.340 160.895 ;
        RECT 27.610 159.455 27.780 160.145 ;
        RECT 27.950 159.795 28.120 159.975 ;
        RECT 28.290 159.965 29.080 160.215 ;
        RECT 29.285 159.795 29.455 160.505 ;
        RECT 29.625 159.995 29.980 160.215 ;
        RECT 27.950 159.625 29.640 159.795 ;
        RECT 26.455 159.025 26.915 159.315 ;
        RECT 27.610 159.285 29.110 159.455 ;
        RECT 27.610 159.145 27.780 159.285 ;
        RECT 27.220 158.975 27.780 159.145 ;
        RECT 25.695 158.345 25.945 158.805 ;
        RECT 26.115 158.515 26.985 158.855 ;
        RECT 27.220 158.515 27.390 158.975 ;
        RECT 28.225 158.945 29.300 159.115 ;
        RECT 27.560 158.345 27.930 158.805 ;
        RECT 28.225 158.605 28.395 158.945 ;
        RECT 28.565 158.345 28.895 158.775 ;
        RECT 29.130 158.605 29.300 158.945 ;
        RECT 29.470 158.845 29.640 159.625 ;
        RECT 29.810 159.405 29.980 159.995 ;
        RECT 30.150 159.595 30.500 160.215 ;
        RECT 29.810 159.015 30.275 159.405 ;
        RECT 30.670 159.145 30.840 160.505 ;
        RECT 31.010 159.315 31.470 160.365 ;
        RECT 30.445 158.975 30.840 159.145 ;
        RECT 30.445 158.845 30.615 158.975 ;
        RECT 29.470 158.515 30.150 158.845 ;
        RECT 30.365 158.515 30.615 158.845 ;
        RECT 30.785 158.345 31.035 158.805 ;
        RECT 31.205 158.530 31.530 159.315 ;
        RECT 31.700 158.515 31.870 160.635 ;
        RECT 32.040 160.515 32.370 160.895 ;
        RECT 32.540 160.345 32.795 160.635 ;
        RECT 32.045 160.175 32.795 160.345 ;
        RECT 32.045 159.185 32.275 160.175 ;
        RECT 32.975 160.155 33.230 160.725 ;
        RECT 33.400 160.495 33.730 160.895 ;
        RECT 34.155 160.360 34.685 160.725 ;
        RECT 34.875 160.555 35.150 160.725 ;
        RECT 34.870 160.385 35.150 160.555 ;
        RECT 34.155 160.325 34.330 160.360 ;
        RECT 33.400 160.155 34.330 160.325 ;
        RECT 32.445 159.355 32.795 160.005 ;
        RECT 32.975 159.485 33.145 160.155 ;
        RECT 33.400 159.985 33.570 160.155 ;
        RECT 33.315 159.655 33.570 159.985 ;
        RECT 33.795 159.655 33.990 159.985 ;
        RECT 32.045 159.015 32.795 159.185 ;
        RECT 32.040 158.345 32.370 158.845 ;
        RECT 32.540 158.515 32.795 159.015 ;
        RECT 32.975 158.515 33.310 159.485 ;
        RECT 33.480 158.345 33.650 159.485 ;
        RECT 33.820 158.685 33.990 159.655 ;
        RECT 34.160 159.025 34.330 160.155 ;
        RECT 34.500 159.365 34.670 160.165 ;
        RECT 34.875 159.565 35.150 160.385 ;
        RECT 35.320 159.365 35.510 160.725 ;
        RECT 35.690 160.360 36.200 160.895 ;
        RECT 36.420 160.085 36.665 160.690 ;
        RECT 37.110 160.220 37.380 160.565 ;
        RECT 37.570 160.495 37.950 160.895 ;
        RECT 38.120 160.325 38.290 160.675 ;
        RECT 38.460 160.495 38.790 160.895 ;
        RECT 38.990 160.325 39.160 160.675 ;
        RECT 39.360 160.395 39.690 160.895 ;
        RECT 35.710 159.915 36.940 160.085 ;
        RECT 34.500 159.195 35.510 159.365 ;
        RECT 35.680 159.350 36.430 159.540 ;
        RECT 34.160 158.855 35.285 159.025 ;
        RECT 35.680 158.685 35.850 159.350 ;
        RECT 36.600 159.105 36.940 159.915 ;
        RECT 33.820 158.515 35.850 158.685 ;
        RECT 36.020 158.345 36.190 159.105 ;
        RECT 36.425 158.695 36.940 159.105 ;
        RECT 37.110 159.485 37.280 160.220 ;
        RECT 37.550 160.155 39.160 160.325 ;
        RECT 37.550 159.985 37.720 160.155 ;
        RECT 37.450 159.655 37.720 159.985 ;
        RECT 37.890 159.655 38.295 159.985 ;
        RECT 37.550 159.485 37.720 159.655 ;
        RECT 38.465 159.535 39.175 159.985 ;
        RECT 39.345 159.655 39.695 160.225 ;
        RECT 39.870 160.095 40.210 160.725 ;
        RECT 40.380 160.095 40.630 160.895 ;
        RECT 40.820 160.245 41.150 160.725 ;
        RECT 41.320 160.435 41.545 160.895 ;
        RECT 41.715 160.245 42.045 160.725 ;
        RECT 39.870 159.535 40.045 160.095 ;
        RECT 40.820 160.075 42.045 160.245 ;
        RECT 42.675 160.115 43.175 160.725 ;
        RECT 40.215 159.735 40.910 159.905 ;
        RECT 37.110 158.515 37.380 159.485 ;
        RECT 37.550 159.315 38.275 159.485 ;
        RECT 38.465 159.365 39.180 159.535 ;
        RECT 39.870 159.485 40.100 159.535 ;
        RECT 40.740 159.485 40.910 159.735 ;
        RECT 41.085 159.705 41.505 159.905 ;
        RECT 41.675 159.705 42.005 159.905 ;
        RECT 42.175 159.705 42.505 159.905 ;
        RECT 42.675 159.485 42.845 160.115 ;
        RECT 43.825 160.085 44.070 160.690 ;
        RECT 44.290 160.360 44.800 160.895 ;
        RECT 43.550 159.915 44.780 160.085 ;
        RECT 43.030 159.655 43.380 159.905 ;
        RECT 38.105 159.195 38.275 159.315 ;
        RECT 39.375 159.195 39.695 159.485 ;
        RECT 37.590 158.345 37.870 159.145 ;
        RECT 38.105 159.025 39.695 159.195 ;
        RECT 38.040 158.565 39.695 158.855 ;
        RECT 39.870 158.515 40.210 159.485 ;
        RECT 40.380 158.345 40.550 159.485 ;
        RECT 40.740 159.315 43.175 159.485 ;
        RECT 40.820 158.345 41.070 159.145 ;
        RECT 41.715 158.515 42.045 159.315 ;
        RECT 42.345 158.345 42.675 159.145 ;
        RECT 42.845 158.515 43.175 159.315 ;
        RECT 43.550 159.105 43.890 159.915 ;
        RECT 44.060 159.350 44.810 159.540 ;
        RECT 43.550 158.695 44.065 159.105 ;
        RECT 44.300 158.345 44.470 159.105 ;
        RECT 44.640 158.685 44.810 159.350 ;
        RECT 44.980 159.365 45.170 160.725 ;
        RECT 45.340 160.215 45.615 160.725 ;
        RECT 45.805 160.360 46.335 160.725 ;
        RECT 46.760 160.495 47.090 160.895 ;
        RECT 46.160 160.325 46.335 160.360 ;
        RECT 45.340 160.045 45.620 160.215 ;
        RECT 45.340 159.565 45.615 160.045 ;
        RECT 45.820 159.365 45.990 160.165 ;
        RECT 44.980 159.195 45.990 159.365 ;
        RECT 46.160 160.155 47.090 160.325 ;
        RECT 47.260 160.155 47.515 160.725 ;
        RECT 47.690 160.170 47.980 160.895 ;
        RECT 48.615 160.185 48.870 160.715 ;
        RECT 49.040 160.435 49.345 160.895 ;
        RECT 49.590 160.515 50.660 160.685 ;
        RECT 46.160 159.025 46.330 160.155 ;
        RECT 46.920 159.985 47.090 160.155 ;
        RECT 45.205 158.855 46.330 159.025 ;
        RECT 46.500 159.655 46.695 159.985 ;
        RECT 46.920 159.655 47.175 159.985 ;
        RECT 46.500 158.685 46.670 159.655 ;
        RECT 47.345 159.485 47.515 160.155 ;
        RECT 48.615 159.535 48.825 160.185 ;
        RECT 49.590 160.160 49.910 160.515 ;
        RECT 49.585 159.985 49.910 160.160 ;
        RECT 48.995 159.685 49.910 159.985 ;
        RECT 50.080 159.945 50.320 160.345 ;
        RECT 50.490 160.285 50.660 160.515 ;
        RECT 50.830 160.455 51.020 160.895 ;
        RECT 51.190 160.445 52.140 160.725 ;
        RECT 52.360 160.535 52.710 160.705 ;
        RECT 50.490 160.115 51.020 160.285 ;
        RECT 48.995 159.655 49.735 159.685 ;
        RECT 44.640 158.515 46.670 158.685 ;
        RECT 46.840 158.345 47.010 159.485 ;
        RECT 47.180 158.515 47.515 159.485 ;
        RECT 47.690 158.345 47.980 159.510 ;
        RECT 48.615 158.655 48.870 159.535 ;
        RECT 49.040 158.345 49.345 159.485 ;
        RECT 49.565 159.065 49.735 159.655 ;
        RECT 50.080 159.575 50.620 159.945 ;
        RECT 50.800 159.835 51.020 160.115 ;
        RECT 51.190 159.665 51.360 160.445 ;
        RECT 50.955 159.495 51.360 159.665 ;
        RECT 51.530 159.655 51.880 160.275 ;
        RECT 50.955 159.405 51.125 159.495 ;
        RECT 52.050 159.485 52.260 160.275 ;
        RECT 49.905 159.235 51.125 159.405 ;
        RECT 51.585 159.325 52.260 159.485 ;
        RECT 49.565 158.895 50.365 159.065 ;
        RECT 49.685 158.345 50.015 158.725 ;
        RECT 50.195 158.605 50.365 158.895 ;
        RECT 50.955 158.855 51.125 159.235 ;
        RECT 51.295 159.315 52.260 159.325 ;
        RECT 52.450 160.145 52.710 160.535 ;
        RECT 52.920 160.435 53.250 160.895 ;
        RECT 54.125 160.505 54.980 160.675 ;
        RECT 55.185 160.505 55.680 160.675 ;
        RECT 55.850 160.535 56.180 160.895 ;
        RECT 52.450 159.455 52.620 160.145 ;
        RECT 52.790 159.795 52.960 159.975 ;
        RECT 53.130 159.965 53.920 160.215 ;
        RECT 54.125 159.795 54.295 160.505 ;
        RECT 54.465 159.995 54.820 160.215 ;
        RECT 52.790 159.625 54.480 159.795 ;
        RECT 51.295 159.025 51.755 159.315 ;
        RECT 52.450 159.285 53.950 159.455 ;
        RECT 52.450 159.145 52.620 159.285 ;
        RECT 52.060 158.975 52.620 159.145 ;
        RECT 50.535 158.345 50.785 158.805 ;
        RECT 50.955 158.515 51.825 158.855 ;
        RECT 52.060 158.515 52.230 158.975 ;
        RECT 53.065 158.945 54.140 159.115 ;
        RECT 52.400 158.345 52.770 158.805 ;
        RECT 53.065 158.605 53.235 158.945 ;
        RECT 53.405 158.345 53.735 158.775 ;
        RECT 53.970 158.605 54.140 158.945 ;
        RECT 54.310 158.845 54.480 159.625 ;
        RECT 54.650 159.405 54.820 159.995 ;
        RECT 54.990 159.595 55.340 160.215 ;
        RECT 54.650 159.015 55.115 159.405 ;
        RECT 55.510 159.145 55.680 160.505 ;
        RECT 55.850 159.315 56.310 160.365 ;
        RECT 55.285 158.975 55.680 159.145 ;
        RECT 55.285 158.845 55.455 158.975 ;
        RECT 54.310 158.515 54.990 158.845 ;
        RECT 55.205 158.515 55.455 158.845 ;
        RECT 55.625 158.345 55.875 158.805 ;
        RECT 56.045 158.530 56.370 159.315 ;
        RECT 56.540 158.515 56.710 160.635 ;
        RECT 56.880 160.515 57.210 160.895 ;
        RECT 57.380 160.345 57.635 160.635 ;
        RECT 56.885 160.175 57.635 160.345 ;
        RECT 58.735 160.185 58.990 160.715 ;
        RECT 59.160 160.435 59.465 160.895 ;
        RECT 59.710 160.515 60.780 160.685 ;
        RECT 56.885 159.185 57.115 160.175 ;
        RECT 57.285 159.355 57.635 160.005 ;
        RECT 58.735 159.535 58.945 160.185 ;
        RECT 59.710 160.160 60.030 160.515 ;
        RECT 59.705 159.985 60.030 160.160 ;
        RECT 59.115 159.685 60.030 159.985 ;
        RECT 60.200 159.945 60.440 160.345 ;
        RECT 60.610 160.285 60.780 160.515 ;
        RECT 60.950 160.455 61.140 160.895 ;
        RECT 61.310 160.445 62.260 160.725 ;
        RECT 62.480 160.535 62.830 160.705 ;
        RECT 60.610 160.115 61.140 160.285 ;
        RECT 59.115 159.655 59.855 159.685 ;
        RECT 56.885 159.015 57.635 159.185 ;
        RECT 56.880 158.345 57.210 158.845 ;
        RECT 57.380 158.515 57.635 159.015 ;
        RECT 58.735 158.655 58.990 159.535 ;
        RECT 59.160 158.345 59.465 159.485 ;
        RECT 59.685 159.065 59.855 159.655 ;
        RECT 60.200 159.575 60.740 159.945 ;
        RECT 60.920 159.835 61.140 160.115 ;
        RECT 61.310 159.665 61.480 160.445 ;
        RECT 61.075 159.495 61.480 159.665 ;
        RECT 61.650 159.655 62.000 160.275 ;
        RECT 61.075 159.405 61.245 159.495 ;
        RECT 62.170 159.485 62.380 160.275 ;
        RECT 60.025 159.235 61.245 159.405 ;
        RECT 61.705 159.325 62.380 159.485 ;
        RECT 59.685 158.895 60.485 159.065 ;
        RECT 59.805 158.345 60.135 158.725 ;
        RECT 60.315 158.605 60.485 158.895 ;
        RECT 61.075 158.855 61.245 159.235 ;
        RECT 61.415 159.315 62.380 159.325 ;
        RECT 62.570 160.145 62.830 160.535 ;
        RECT 63.040 160.435 63.370 160.895 ;
        RECT 64.245 160.505 65.100 160.675 ;
        RECT 65.305 160.505 65.800 160.675 ;
        RECT 65.970 160.535 66.300 160.895 ;
        RECT 62.570 159.455 62.740 160.145 ;
        RECT 62.910 159.795 63.080 159.975 ;
        RECT 63.250 159.965 64.040 160.215 ;
        RECT 64.245 159.795 64.415 160.505 ;
        RECT 64.585 159.995 64.940 160.215 ;
        RECT 62.910 159.625 64.600 159.795 ;
        RECT 61.415 159.025 61.875 159.315 ;
        RECT 62.570 159.285 64.070 159.455 ;
        RECT 62.570 159.145 62.740 159.285 ;
        RECT 62.180 158.975 62.740 159.145 ;
        RECT 60.655 158.345 60.905 158.805 ;
        RECT 61.075 158.515 61.945 158.855 ;
        RECT 62.180 158.515 62.350 158.975 ;
        RECT 63.185 158.945 64.260 159.115 ;
        RECT 62.520 158.345 62.890 158.805 ;
        RECT 63.185 158.605 63.355 158.945 ;
        RECT 63.525 158.345 63.855 158.775 ;
        RECT 64.090 158.605 64.260 158.945 ;
        RECT 64.430 158.845 64.600 159.625 ;
        RECT 64.770 159.405 64.940 159.995 ;
        RECT 65.110 159.595 65.460 160.215 ;
        RECT 64.770 159.015 65.235 159.405 ;
        RECT 65.630 159.145 65.800 160.505 ;
        RECT 65.970 159.315 66.430 160.365 ;
        RECT 65.405 158.975 65.800 159.145 ;
        RECT 65.405 158.845 65.575 158.975 ;
        RECT 64.430 158.515 65.110 158.845 ;
        RECT 65.325 158.515 65.575 158.845 ;
        RECT 65.745 158.345 65.995 158.805 ;
        RECT 66.165 158.530 66.490 159.315 ;
        RECT 66.660 158.515 66.830 160.635 ;
        RECT 67.000 160.515 67.330 160.895 ;
        RECT 67.500 160.345 67.755 160.635 ;
        RECT 67.005 160.175 67.755 160.345 ;
        RECT 67.005 159.185 67.235 160.175 ;
        RECT 67.970 160.075 68.200 160.895 ;
        RECT 68.370 160.095 68.700 160.725 ;
        RECT 67.405 159.355 67.755 160.005 ;
        RECT 67.950 159.655 68.280 159.905 ;
        RECT 68.450 159.495 68.700 160.095 ;
        RECT 68.870 160.075 69.080 160.895 ;
        RECT 69.585 160.085 69.830 160.690 ;
        RECT 70.050 160.360 70.560 160.895 ;
        RECT 67.005 159.015 67.755 159.185 ;
        RECT 67.000 158.345 67.330 158.845 ;
        RECT 67.500 158.515 67.755 159.015 ;
        RECT 67.970 158.345 68.200 159.485 ;
        RECT 68.370 158.515 68.700 159.495 ;
        RECT 69.310 159.915 70.540 160.085 ;
        RECT 68.870 158.345 69.080 159.485 ;
        RECT 69.310 159.105 69.650 159.915 ;
        RECT 69.820 159.350 70.570 159.540 ;
        RECT 69.310 158.695 69.825 159.105 ;
        RECT 70.060 158.345 70.230 159.105 ;
        RECT 70.400 158.685 70.570 159.350 ;
        RECT 70.740 159.365 70.930 160.725 ;
        RECT 71.100 160.555 71.375 160.725 ;
        RECT 71.100 160.385 71.380 160.555 ;
        RECT 71.100 159.565 71.375 160.385 ;
        RECT 71.565 160.360 72.095 160.725 ;
        RECT 72.520 160.495 72.850 160.895 ;
        RECT 71.920 160.325 72.095 160.360 ;
        RECT 71.580 159.365 71.750 160.165 ;
        RECT 70.740 159.195 71.750 159.365 ;
        RECT 71.920 160.155 72.850 160.325 ;
        RECT 73.020 160.155 73.275 160.725 ;
        RECT 73.450 160.170 73.740 160.895 ;
        RECT 74.285 160.555 74.540 160.715 ;
        RECT 74.200 160.385 74.540 160.555 ;
        RECT 74.720 160.435 75.005 160.895 ;
        RECT 74.285 160.185 74.540 160.385 ;
        RECT 71.920 159.025 72.090 160.155 ;
        RECT 72.680 159.985 72.850 160.155 ;
        RECT 70.965 158.855 72.090 159.025 ;
        RECT 72.260 159.655 72.455 159.985 ;
        RECT 72.680 159.655 72.935 159.985 ;
        RECT 72.260 158.685 72.430 159.655 ;
        RECT 73.105 159.485 73.275 160.155 ;
        RECT 70.400 158.515 72.430 158.685 ;
        RECT 72.600 158.345 72.770 159.485 ;
        RECT 72.940 158.515 73.275 159.485 ;
        RECT 73.450 158.345 73.740 159.510 ;
        RECT 74.285 159.325 74.465 160.185 ;
        RECT 75.185 159.985 75.435 160.635 ;
        RECT 74.635 159.655 75.435 159.985 ;
        RECT 74.285 158.655 74.540 159.325 ;
        RECT 74.720 158.345 75.005 159.145 ;
        RECT 75.185 159.065 75.435 159.655 ;
        RECT 75.635 160.300 75.955 160.630 ;
        RECT 76.135 160.415 76.795 160.895 ;
        RECT 76.995 160.505 77.845 160.675 ;
        RECT 75.635 159.405 75.825 160.300 ;
        RECT 76.145 159.975 76.805 160.245 ;
        RECT 76.475 159.915 76.805 159.975 ;
        RECT 75.995 159.745 76.325 159.805 ;
        RECT 76.995 159.745 77.165 160.505 ;
        RECT 78.405 160.435 78.725 160.895 ;
        RECT 78.925 160.255 79.175 160.685 ;
        RECT 79.465 160.455 79.875 160.895 ;
        RECT 80.045 160.515 81.060 160.715 ;
        RECT 77.335 160.085 78.585 160.255 ;
        RECT 77.335 159.965 77.665 160.085 ;
        RECT 75.995 159.575 77.895 159.745 ;
        RECT 75.635 159.235 77.555 159.405 ;
        RECT 75.635 159.215 75.955 159.235 ;
        RECT 75.185 158.555 75.515 159.065 ;
        RECT 75.785 158.605 75.955 159.215 ;
        RECT 77.725 159.065 77.895 159.575 ;
        RECT 78.065 159.505 78.245 159.915 ;
        RECT 78.415 159.325 78.585 160.085 ;
        RECT 76.125 158.345 76.455 159.035 ;
        RECT 76.685 158.895 77.895 159.065 ;
        RECT 78.065 159.015 78.585 159.325 ;
        RECT 78.755 159.915 79.175 160.255 ;
        RECT 79.465 159.915 79.875 160.245 ;
        RECT 78.755 159.145 78.945 159.915 ;
        RECT 80.045 159.785 80.215 160.515 ;
        RECT 81.360 160.345 81.530 160.675 ;
        RECT 81.700 160.515 82.030 160.895 ;
        RECT 80.385 159.965 80.735 160.335 ;
        RECT 80.045 159.745 80.465 159.785 ;
        RECT 79.115 159.575 80.465 159.745 ;
        RECT 79.115 159.415 79.365 159.575 ;
        RECT 79.875 159.145 80.125 159.405 ;
        RECT 78.755 158.895 80.125 159.145 ;
        RECT 76.685 158.605 76.925 158.895 ;
        RECT 77.725 158.815 77.895 158.895 ;
        RECT 77.125 158.345 77.545 158.725 ;
        RECT 77.725 158.565 78.355 158.815 ;
        RECT 78.825 158.345 79.155 158.725 ;
        RECT 79.325 158.605 79.495 158.895 ;
        RECT 80.295 158.730 80.465 159.575 ;
        RECT 80.915 159.405 81.135 160.275 ;
        RECT 81.360 160.155 82.055 160.345 ;
        RECT 80.635 159.025 81.135 159.405 ;
        RECT 81.305 159.355 81.715 159.975 ;
        RECT 81.885 159.185 82.055 160.155 ;
        RECT 81.360 159.015 82.055 159.185 ;
        RECT 79.675 158.345 80.055 158.725 ;
        RECT 80.295 158.560 81.125 158.730 ;
        RECT 81.360 158.515 81.530 159.015 ;
        RECT 81.700 158.345 82.030 158.845 ;
        RECT 82.245 158.515 82.470 160.635 ;
        RECT 82.640 160.515 82.970 160.895 ;
        RECT 83.140 160.345 83.310 160.635 ;
        RECT 82.645 160.175 83.310 160.345 ;
        RECT 82.645 159.185 82.875 160.175 ;
        RECT 83.775 160.115 84.275 160.725 ;
        RECT 83.045 159.355 83.395 160.005 ;
        RECT 83.570 159.655 83.920 159.905 ;
        RECT 84.105 159.485 84.275 160.115 ;
        RECT 84.905 160.245 85.235 160.725 ;
        RECT 85.405 160.435 85.630 160.895 ;
        RECT 85.800 160.245 86.130 160.725 ;
        RECT 84.905 160.075 86.130 160.245 ;
        RECT 86.320 160.095 86.570 160.895 ;
        RECT 86.740 160.095 87.080 160.725 ;
        RECT 84.445 159.705 84.775 159.905 ;
        RECT 84.945 159.705 85.275 159.905 ;
        RECT 85.445 159.705 85.865 159.905 ;
        RECT 86.040 159.735 86.735 159.905 ;
        RECT 86.040 159.485 86.210 159.735 ;
        RECT 86.905 159.485 87.080 160.095 ;
        RECT 83.775 159.315 86.210 159.485 ;
        RECT 82.645 159.015 83.310 159.185 ;
        RECT 82.640 158.345 82.970 158.845 ;
        RECT 83.140 158.515 83.310 159.015 ;
        RECT 83.775 158.515 84.105 159.315 ;
        RECT 84.275 158.345 84.605 159.145 ;
        RECT 84.905 158.515 85.235 159.315 ;
        RECT 85.880 158.345 86.130 159.145 ;
        RECT 86.400 158.345 86.570 159.485 ;
        RECT 86.740 158.515 87.080 159.485 ;
        RECT 87.710 160.095 88.050 160.725 ;
        RECT 88.220 160.095 88.470 160.895 ;
        RECT 88.660 160.245 88.990 160.725 ;
        RECT 89.160 160.435 89.385 160.895 ;
        RECT 89.555 160.245 89.885 160.725 ;
        RECT 87.710 159.485 87.885 160.095 ;
        RECT 88.660 160.075 89.885 160.245 ;
        RECT 90.515 160.115 91.015 160.725 ;
        RECT 91.505 160.265 91.790 160.725 ;
        RECT 91.960 160.435 92.230 160.895 ;
        RECT 88.055 159.735 88.750 159.905 ;
        RECT 88.580 159.485 88.750 159.735 ;
        RECT 88.925 159.705 89.345 159.905 ;
        RECT 89.515 159.705 89.845 159.905 ;
        RECT 90.015 159.705 90.345 159.905 ;
        RECT 90.515 159.485 90.685 160.115 ;
        RECT 91.505 160.095 92.460 160.265 ;
        RECT 90.870 159.655 91.220 159.905 ;
        RECT 87.710 158.515 88.050 159.485 ;
        RECT 88.220 158.345 88.390 159.485 ;
        RECT 88.580 159.315 91.015 159.485 ;
        RECT 91.390 159.365 92.080 159.925 ;
        RECT 88.660 158.345 88.910 159.145 ;
        RECT 89.555 158.515 89.885 159.315 ;
        RECT 90.185 158.345 90.515 159.145 ;
        RECT 90.685 158.515 91.015 159.315 ;
        RECT 92.250 159.195 92.460 160.095 ;
        RECT 91.505 158.975 92.460 159.195 ;
        RECT 92.630 159.925 93.030 160.725 ;
        RECT 93.220 160.265 93.500 160.725 ;
        RECT 94.020 160.435 94.345 160.895 ;
        RECT 93.220 160.095 94.345 160.265 ;
        RECT 94.515 160.155 94.900 160.725 ;
        RECT 93.895 159.985 94.345 160.095 ;
        RECT 92.630 159.365 93.725 159.925 ;
        RECT 93.895 159.655 94.450 159.985 ;
        RECT 91.505 158.515 91.790 158.975 ;
        RECT 91.960 158.345 92.230 158.805 ;
        RECT 92.630 158.515 93.030 159.365 ;
        RECT 93.895 159.195 94.345 159.655 ;
        RECT 94.620 159.485 94.900 160.155 ;
        RECT 95.345 160.085 95.590 160.690 ;
        RECT 95.810 160.360 96.320 160.895 ;
        RECT 93.220 158.975 94.345 159.195 ;
        RECT 93.220 158.515 93.500 158.975 ;
        RECT 94.020 158.345 94.345 158.805 ;
        RECT 94.515 158.515 94.900 159.485 ;
        RECT 95.070 159.915 96.300 160.085 ;
        RECT 95.070 159.105 95.410 159.915 ;
        RECT 95.580 159.350 96.330 159.540 ;
        RECT 95.070 158.695 95.585 159.105 ;
        RECT 95.820 158.345 95.990 159.105 ;
        RECT 96.160 158.685 96.330 159.350 ;
        RECT 96.500 159.365 96.690 160.725 ;
        RECT 96.860 159.875 97.135 160.725 ;
        RECT 97.325 160.360 97.855 160.725 ;
        RECT 98.280 160.495 98.610 160.895 ;
        RECT 97.680 160.325 97.855 160.360 ;
        RECT 96.860 159.705 97.140 159.875 ;
        RECT 96.860 159.565 97.135 159.705 ;
        RECT 97.340 159.365 97.510 160.165 ;
        RECT 96.500 159.195 97.510 159.365 ;
        RECT 97.680 160.155 98.610 160.325 ;
        RECT 98.780 160.155 99.035 160.725 ;
        RECT 99.210 160.170 99.500 160.895 ;
        RECT 97.680 159.025 97.850 160.155 ;
        RECT 98.440 159.985 98.610 160.155 ;
        RECT 96.725 158.855 97.850 159.025 ;
        RECT 98.020 159.655 98.215 159.985 ;
        RECT 98.440 159.655 98.695 159.985 ;
        RECT 98.020 158.685 98.190 159.655 ;
        RECT 98.865 159.485 99.035 160.155 ;
        RECT 99.875 160.115 100.375 160.725 ;
        RECT 99.670 159.655 100.020 159.905 ;
        RECT 96.160 158.515 98.190 158.685 ;
        RECT 98.360 158.345 98.530 159.485 ;
        RECT 98.700 158.515 99.035 159.485 ;
        RECT 99.210 158.345 99.500 159.510 ;
        RECT 100.205 159.485 100.375 160.115 ;
        RECT 101.005 160.245 101.335 160.725 ;
        RECT 101.505 160.435 101.730 160.895 ;
        RECT 101.900 160.245 102.230 160.725 ;
        RECT 101.005 160.075 102.230 160.245 ;
        RECT 102.420 160.095 102.670 160.895 ;
        RECT 102.840 160.095 103.180 160.725 ;
        RECT 100.545 159.705 100.875 159.905 ;
        RECT 101.045 159.705 101.375 159.905 ;
        RECT 101.545 159.705 101.965 159.905 ;
        RECT 102.140 159.735 102.835 159.905 ;
        RECT 102.140 159.485 102.310 159.735 ;
        RECT 103.005 159.485 103.180 160.095 ;
        RECT 103.390 160.075 103.620 160.895 ;
        RECT 103.790 160.095 104.120 160.725 ;
        RECT 103.370 159.655 103.700 159.905 ;
        RECT 103.870 159.495 104.120 160.095 ;
        RECT 104.290 160.075 104.500 160.895 ;
        RECT 104.790 160.075 105.000 160.895 ;
        RECT 105.170 160.095 105.500 160.725 ;
        RECT 99.875 159.315 102.310 159.485 ;
        RECT 99.875 158.515 100.205 159.315 ;
        RECT 100.375 158.345 100.705 159.145 ;
        RECT 101.005 158.515 101.335 159.315 ;
        RECT 101.980 158.345 102.230 159.145 ;
        RECT 102.500 158.345 102.670 159.485 ;
        RECT 102.840 158.515 103.180 159.485 ;
        RECT 103.390 158.345 103.620 159.485 ;
        RECT 103.790 158.515 104.120 159.495 ;
        RECT 105.170 159.495 105.420 160.095 ;
        RECT 105.670 160.075 105.900 160.895 ;
        RECT 106.110 160.145 107.320 160.895 ;
        RECT 105.590 159.655 105.920 159.905 ;
        RECT 104.290 158.345 104.500 159.485 ;
        RECT 104.790 158.345 105.000 159.485 ;
        RECT 105.170 158.515 105.500 159.495 ;
        RECT 105.670 158.345 105.900 159.485 ;
        RECT 106.110 159.435 106.630 159.975 ;
        RECT 106.800 159.605 107.320 160.145 ;
        RECT 107.490 160.125 111.000 160.895 ;
        RECT 111.170 160.145 112.380 160.895 ;
        RECT 107.490 159.435 109.180 159.955 ;
        RECT 109.350 159.605 111.000 160.125 ;
        RECT 111.170 159.435 111.690 159.975 ;
        RECT 111.860 159.605 112.380 160.145 ;
        RECT 106.110 158.345 107.320 159.435 ;
        RECT 107.490 158.345 111.000 159.435 ;
        RECT 111.170 158.345 112.380 159.435 ;
        RECT 18.165 158.175 112.465 158.345 ;
        RECT 18.250 157.085 19.460 158.175 ;
        RECT 18.250 156.375 18.770 156.915 ;
        RECT 18.940 156.545 19.460 157.085 ;
        RECT 19.630 157.085 22.220 158.175 ;
        RECT 22.470 157.245 22.650 158.005 ;
        RECT 22.830 157.415 23.160 158.175 ;
        RECT 19.630 156.565 20.840 157.085 ;
        RECT 22.470 157.075 23.145 157.245 ;
        RECT 23.330 157.100 23.600 158.005 ;
        RECT 24.235 157.740 29.580 158.175 ;
        RECT 22.975 156.930 23.145 157.075 ;
        RECT 21.010 156.395 22.220 156.915 ;
        RECT 22.410 156.525 22.750 156.895 ;
        RECT 22.975 156.600 23.250 156.930 ;
        RECT 18.250 155.625 19.460 156.375 ;
        RECT 19.630 155.625 22.220 156.395 ;
        RECT 22.975 156.345 23.145 156.600 ;
        RECT 22.480 156.175 23.145 156.345 ;
        RECT 23.420 156.300 23.600 157.100 ;
        RECT 25.825 156.490 26.175 157.740 ;
        RECT 29.810 157.035 30.020 158.175 ;
        RECT 30.190 157.025 30.520 158.005 ;
        RECT 30.690 157.035 30.920 158.175 ;
        RECT 31.335 157.205 31.665 158.005 ;
        RECT 31.835 157.375 32.165 158.175 ;
        RECT 32.465 157.205 32.795 158.005 ;
        RECT 33.440 157.375 33.690 158.175 ;
        RECT 31.335 157.035 33.770 157.205 ;
        RECT 33.960 157.035 34.130 158.175 ;
        RECT 34.300 157.035 34.640 158.005 ;
        RECT 22.480 155.795 22.650 156.175 ;
        RECT 22.830 155.625 23.160 156.005 ;
        RECT 23.340 155.795 23.600 156.300 ;
        RECT 27.655 156.170 27.995 157.000 ;
        RECT 24.235 155.625 29.580 156.170 ;
        RECT 29.810 155.625 30.020 156.445 ;
        RECT 30.190 156.425 30.440 157.025 ;
        RECT 30.610 156.615 30.940 156.865 ;
        RECT 31.130 156.615 31.480 156.865 ;
        RECT 30.190 155.795 30.520 156.425 ;
        RECT 30.690 155.625 30.920 156.445 ;
        RECT 31.665 156.405 31.835 157.035 ;
        RECT 32.005 156.615 32.335 156.815 ;
        RECT 32.505 156.615 32.835 156.815 ;
        RECT 33.005 156.615 33.425 156.815 ;
        RECT 33.600 156.785 33.770 157.035 ;
        RECT 33.600 156.615 34.295 156.785 ;
        RECT 31.335 155.795 31.835 156.405 ;
        RECT 32.465 156.275 33.690 156.445 ;
        RECT 34.465 156.425 34.640 157.035 ;
        RECT 34.810 157.010 35.100 158.175 ;
        RECT 35.275 157.025 35.535 158.175 ;
        RECT 35.710 157.100 35.965 158.005 ;
        RECT 36.135 157.415 36.465 158.175 ;
        RECT 36.680 157.245 36.850 158.005 ;
        RECT 32.465 155.795 32.795 156.275 ;
        RECT 32.965 155.625 33.190 156.085 ;
        RECT 33.360 155.795 33.690 156.275 ;
        RECT 33.880 155.625 34.130 156.425 ;
        RECT 34.300 155.795 34.640 156.425 ;
        RECT 34.810 155.625 35.100 156.350 ;
        RECT 35.275 155.625 35.535 156.465 ;
        RECT 35.710 156.370 35.880 157.100 ;
        RECT 36.135 157.075 36.850 157.245 ;
        RECT 37.110 157.455 37.570 158.005 ;
        RECT 37.760 157.455 38.090 158.175 ;
        RECT 36.135 156.865 36.305 157.075 ;
        RECT 36.050 156.535 36.305 156.865 ;
        RECT 35.710 155.795 35.965 156.370 ;
        RECT 36.135 156.345 36.305 156.535 ;
        RECT 36.585 156.525 36.940 156.895 ;
        RECT 36.135 156.175 36.850 156.345 ;
        RECT 36.135 155.625 36.465 156.005 ;
        RECT 36.680 155.795 36.850 156.175 ;
        RECT 37.110 156.085 37.360 157.455 ;
        RECT 38.290 157.285 38.590 157.835 ;
        RECT 38.760 157.505 39.040 158.175 ;
        RECT 37.650 157.115 38.590 157.285 ;
        RECT 37.650 156.865 37.820 157.115 ;
        RECT 38.960 156.865 39.225 157.225 ;
        RECT 37.530 156.535 37.820 156.865 ;
        RECT 37.990 156.615 38.330 156.865 ;
        RECT 38.550 156.615 39.225 156.865 ;
        RECT 39.410 157.035 39.750 158.005 ;
        RECT 39.920 157.035 40.090 158.175 ;
        RECT 40.360 157.375 40.610 158.175 ;
        RECT 41.255 157.205 41.585 158.005 ;
        RECT 41.885 157.375 42.215 158.175 ;
        RECT 42.385 157.205 42.715 158.005 ;
        RECT 40.280 157.035 42.715 157.205 ;
        RECT 37.650 156.445 37.820 156.535 ;
        RECT 37.650 156.255 39.040 156.445 ;
        RECT 37.110 155.795 37.670 156.085 ;
        RECT 37.840 155.625 38.090 156.085 ;
        RECT 38.710 155.895 39.040 156.255 ;
        RECT 39.410 156.425 39.585 157.035 ;
        RECT 40.280 156.785 40.450 157.035 ;
        RECT 39.755 156.615 40.450 156.785 ;
        RECT 40.625 156.615 41.045 156.815 ;
        RECT 41.215 156.615 41.545 156.815 ;
        RECT 41.715 156.615 42.045 156.815 ;
        RECT 39.410 155.795 39.750 156.425 ;
        RECT 39.920 155.625 40.170 156.425 ;
        RECT 40.360 156.275 41.585 156.445 ;
        RECT 40.360 155.795 40.690 156.275 ;
        RECT 40.860 155.625 41.085 156.085 ;
        RECT 41.255 155.795 41.585 156.275 ;
        RECT 42.215 156.405 42.385 157.035 ;
        RECT 43.095 156.985 43.350 157.865 ;
        RECT 43.520 157.035 43.825 158.175 ;
        RECT 44.165 157.795 44.495 158.175 ;
        RECT 44.675 157.625 44.845 157.915 ;
        RECT 45.015 157.715 45.265 158.175 ;
        RECT 44.045 157.455 44.845 157.625 ;
        RECT 45.435 157.665 46.305 158.005 ;
        RECT 42.570 156.615 42.920 156.865 ;
        RECT 42.215 155.795 42.715 156.405 ;
        RECT 43.095 156.335 43.305 156.985 ;
        RECT 44.045 156.865 44.215 157.455 ;
        RECT 45.435 157.285 45.605 157.665 ;
        RECT 46.540 157.545 46.710 158.005 ;
        RECT 46.880 157.715 47.250 158.175 ;
        RECT 47.545 157.575 47.715 157.915 ;
        RECT 47.885 157.745 48.215 158.175 ;
        RECT 48.450 157.575 48.620 157.915 ;
        RECT 44.385 157.115 45.605 157.285 ;
        RECT 45.775 157.205 46.235 157.495 ;
        RECT 46.540 157.375 47.100 157.545 ;
        RECT 47.545 157.405 48.620 157.575 ;
        RECT 48.790 157.675 49.470 158.005 ;
        RECT 49.685 157.675 49.935 158.005 ;
        RECT 50.105 157.715 50.355 158.175 ;
        RECT 46.930 157.235 47.100 157.375 ;
        RECT 45.775 157.195 46.740 157.205 ;
        RECT 45.435 157.025 45.605 157.115 ;
        RECT 46.065 157.035 46.740 157.195 ;
        RECT 43.475 156.835 44.215 156.865 ;
        RECT 43.475 156.535 44.390 156.835 ;
        RECT 44.065 156.360 44.390 156.535 ;
        RECT 43.095 155.805 43.350 156.335 ;
        RECT 43.520 155.625 43.825 156.085 ;
        RECT 44.070 156.005 44.390 156.360 ;
        RECT 44.560 156.575 45.100 156.945 ;
        RECT 45.435 156.855 45.840 157.025 ;
        RECT 44.560 156.175 44.800 156.575 ;
        RECT 45.280 156.405 45.500 156.685 ;
        RECT 44.970 156.235 45.500 156.405 ;
        RECT 44.970 156.005 45.140 156.235 ;
        RECT 45.670 156.075 45.840 156.855 ;
        RECT 46.010 156.245 46.360 156.865 ;
        RECT 46.530 156.245 46.740 157.035 ;
        RECT 46.930 157.065 48.430 157.235 ;
        RECT 46.930 156.375 47.100 157.065 ;
        RECT 48.790 156.895 48.960 157.675 ;
        RECT 49.765 157.545 49.935 157.675 ;
        RECT 47.270 156.725 48.960 156.895 ;
        RECT 49.130 157.115 49.595 157.505 ;
        RECT 49.765 157.375 50.160 157.545 ;
        RECT 47.270 156.545 47.440 156.725 ;
        RECT 44.070 155.835 45.140 156.005 ;
        RECT 45.310 155.625 45.500 156.065 ;
        RECT 45.670 155.795 46.620 156.075 ;
        RECT 46.930 155.985 47.190 156.375 ;
        RECT 47.610 156.305 48.400 156.555 ;
        RECT 46.840 155.815 47.190 155.985 ;
        RECT 47.400 155.625 47.730 156.085 ;
        RECT 48.605 156.015 48.775 156.725 ;
        RECT 49.130 156.525 49.300 157.115 ;
        RECT 48.945 156.305 49.300 156.525 ;
        RECT 49.470 156.305 49.820 156.925 ;
        RECT 49.990 156.015 50.160 157.375 ;
        RECT 50.525 157.205 50.850 157.990 ;
        RECT 50.330 156.155 50.790 157.205 ;
        RECT 48.605 155.845 49.460 156.015 ;
        RECT 49.665 155.845 50.160 156.015 ;
        RECT 50.330 155.625 50.660 155.985 ;
        RECT 51.020 155.885 51.190 158.005 ;
        RECT 51.360 157.675 51.690 158.175 ;
        RECT 51.860 157.505 52.115 158.005 ;
        RECT 51.365 157.335 52.115 157.505 ;
        RECT 52.405 157.545 52.690 158.005 ;
        RECT 52.860 157.715 53.130 158.175 ;
        RECT 51.365 156.345 51.595 157.335 ;
        RECT 52.405 157.325 53.360 157.545 ;
        RECT 51.765 156.515 52.115 157.165 ;
        RECT 52.290 156.595 52.980 157.155 ;
        RECT 53.150 156.425 53.360 157.325 ;
        RECT 51.365 156.175 52.115 156.345 ;
        RECT 51.360 155.625 51.690 156.005 ;
        RECT 51.860 155.885 52.115 156.175 ;
        RECT 52.405 156.255 53.360 156.425 ;
        RECT 53.530 157.155 53.930 158.005 ;
        RECT 54.120 157.545 54.400 158.005 ;
        RECT 54.920 157.715 55.245 158.175 ;
        RECT 54.120 157.325 55.245 157.545 ;
        RECT 53.530 156.595 54.625 157.155 ;
        RECT 54.795 156.865 55.245 157.325 ;
        RECT 55.415 157.035 55.800 158.005 ;
        RECT 52.405 155.795 52.690 156.255 ;
        RECT 52.860 155.625 53.130 156.085 ;
        RECT 53.530 155.795 53.930 156.595 ;
        RECT 54.795 156.535 55.350 156.865 ;
        RECT 54.795 156.425 55.245 156.535 ;
        RECT 54.120 156.255 55.245 156.425 ;
        RECT 55.520 156.365 55.800 157.035 ;
        RECT 54.120 155.795 54.400 156.255 ;
        RECT 54.920 155.625 55.245 156.085 ;
        RECT 55.415 155.795 55.800 156.365 ;
        RECT 56.890 157.035 57.230 158.005 ;
        RECT 57.400 157.035 57.570 158.175 ;
        RECT 57.840 157.375 58.090 158.175 ;
        RECT 58.735 157.205 59.065 158.005 ;
        RECT 59.365 157.375 59.695 158.175 ;
        RECT 59.865 157.205 60.195 158.005 ;
        RECT 57.760 157.035 60.195 157.205 ;
        RECT 56.890 156.425 57.065 157.035 ;
        RECT 57.760 156.785 57.930 157.035 ;
        RECT 57.235 156.615 57.930 156.785 ;
        RECT 58.105 156.615 58.525 156.815 ;
        RECT 58.695 156.615 59.025 156.815 ;
        RECT 59.195 156.615 59.525 156.815 ;
        RECT 56.890 155.795 57.230 156.425 ;
        RECT 57.400 155.625 57.650 156.425 ;
        RECT 57.840 156.275 59.065 156.445 ;
        RECT 57.840 155.795 58.170 156.275 ;
        RECT 58.340 155.625 58.565 156.085 ;
        RECT 58.735 155.795 59.065 156.275 ;
        RECT 59.695 156.405 59.865 157.035 ;
        RECT 60.570 157.010 60.860 158.175 ;
        RECT 61.490 157.035 61.830 158.005 ;
        RECT 62.000 157.035 62.170 158.175 ;
        RECT 62.440 157.375 62.690 158.175 ;
        RECT 63.335 157.205 63.665 158.005 ;
        RECT 63.965 157.375 64.295 158.175 ;
        RECT 64.465 157.205 64.795 158.005 ;
        RECT 62.360 157.035 64.795 157.205 ;
        RECT 65.170 157.085 66.380 158.175 ;
        RECT 66.925 157.195 67.180 157.865 ;
        RECT 67.360 157.375 67.645 158.175 ;
        RECT 67.825 157.455 68.155 157.965 ;
        RECT 60.050 156.615 60.400 156.865 ;
        RECT 61.490 156.425 61.665 157.035 ;
        RECT 62.360 156.785 62.530 157.035 ;
        RECT 61.835 156.615 62.530 156.785 ;
        RECT 62.705 156.615 63.125 156.815 ;
        RECT 63.295 156.615 63.625 156.815 ;
        RECT 63.795 156.615 64.125 156.815 ;
        RECT 59.695 155.795 60.195 156.405 ;
        RECT 60.570 155.625 60.860 156.350 ;
        RECT 61.490 155.795 61.830 156.425 ;
        RECT 62.000 155.625 62.250 156.425 ;
        RECT 62.440 156.275 63.665 156.445 ;
        RECT 62.440 155.795 62.770 156.275 ;
        RECT 62.940 155.625 63.165 156.085 ;
        RECT 63.335 155.795 63.665 156.275 ;
        RECT 64.295 156.405 64.465 157.035 ;
        RECT 64.650 156.615 65.000 156.865 ;
        RECT 65.170 156.545 65.690 157.085 ;
        RECT 64.295 155.795 64.795 156.405 ;
        RECT 65.860 156.375 66.380 156.915 ;
        RECT 65.170 155.625 66.380 156.375 ;
        RECT 66.925 156.335 67.105 157.195 ;
        RECT 67.825 156.865 68.075 157.455 ;
        RECT 68.425 157.305 68.595 157.915 ;
        RECT 68.765 157.485 69.095 158.175 ;
        RECT 69.325 157.625 69.565 157.915 ;
        RECT 69.765 157.795 70.185 158.175 ;
        RECT 70.365 157.705 70.995 157.955 ;
        RECT 71.465 157.795 71.795 158.175 ;
        RECT 70.365 157.625 70.535 157.705 ;
        RECT 71.965 157.625 72.135 157.915 ;
        RECT 72.315 157.795 72.695 158.175 ;
        RECT 72.935 157.790 73.765 157.960 ;
        RECT 69.325 157.455 70.535 157.625 ;
        RECT 67.275 156.535 68.075 156.865 ;
        RECT 66.925 156.135 67.180 156.335 ;
        RECT 66.840 155.965 67.180 156.135 ;
        RECT 66.925 155.805 67.180 155.965 ;
        RECT 67.360 155.625 67.645 156.085 ;
        RECT 67.825 155.885 68.075 156.535 ;
        RECT 68.275 157.285 68.595 157.305 ;
        RECT 68.275 157.115 70.195 157.285 ;
        RECT 68.275 156.220 68.465 157.115 ;
        RECT 70.365 156.945 70.535 157.455 ;
        RECT 70.705 157.195 71.225 157.505 ;
        RECT 68.635 156.775 70.535 156.945 ;
        RECT 68.635 156.715 68.965 156.775 ;
        RECT 69.115 156.545 69.445 156.605 ;
        RECT 68.785 156.275 69.445 156.545 ;
        RECT 68.275 155.890 68.595 156.220 ;
        RECT 68.775 155.625 69.435 156.105 ;
        RECT 69.635 156.015 69.805 156.775 ;
        RECT 70.705 156.605 70.885 157.015 ;
        RECT 69.975 156.435 70.305 156.555 ;
        RECT 71.055 156.435 71.225 157.195 ;
        RECT 69.975 156.265 71.225 156.435 ;
        RECT 71.395 157.375 72.765 157.625 ;
        RECT 71.395 156.605 71.585 157.375 ;
        RECT 72.515 157.115 72.765 157.375 ;
        RECT 71.755 156.945 72.005 157.105 ;
        RECT 72.935 156.945 73.105 157.790 ;
        RECT 74.000 157.505 74.170 158.005 ;
        RECT 74.340 157.675 74.670 158.175 ;
        RECT 73.275 157.115 73.775 157.495 ;
        RECT 74.000 157.335 74.695 157.505 ;
        RECT 71.755 156.775 73.105 156.945 ;
        RECT 72.685 156.735 73.105 156.775 ;
        RECT 71.395 156.265 71.815 156.605 ;
        RECT 72.105 156.275 72.515 156.605 ;
        RECT 69.635 155.845 70.485 156.015 ;
        RECT 71.045 155.625 71.365 156.085 ;
        RECT 71.565 155.835 71.815 156.265 ;
        RECT 72.105 155.625 72.515 156.065 ;
        RECT 72.685 156.005 72.855 156.735 ;
        RECT 73.025 156.185 73.375 156.555 ;
        RECT 73.555 156.245 73.775 157.115 ;
        RECT 73.945 156.545 74.355 157.165 ;
        RECT 74.525 156.365 74.695 157.335 ;
        RECT 74.000 156.175 74.695 156.365 ;
        RECT 72.685 155.805 73.700 156.005 ;
        RECT 74.000 155.845 74.170 156.175 ;
        RECT 74.340 155.625 74.670 156.005 ;
        RECT 74.885 155.885 75.110 158.005 ;
        RECT 75.280 157.675 75.610 158.175 ;
        RECT 75.780 157.505 75.950 158.005 ;
        RECT 75.285 157.335 75.950 157.505 ;
        RECT 75.285 156.345 75.515 157.335 ;
        RECT 75.685 156.515 76.035 157.165 ;
        RECT 76.710 157.035 76.940 158.175 ;
        RECT 77.110 157.025 77.440 158.005 ;
        RECT 77.610 157.035 77.820 158.175 ;
        RECT 78.510 157.085 81.100 158.175 ;
        RECT 76.690 156.615 77.020 156.865 ;
        RECT 75.285 156.175 75.950 156.345 ;
        RECT 75.280 155.625 75.610 156.005 ;
        RECT 75.780 155.885 75.950 156.175 ;
        RECT 76.710 155.625 76.940 156.445 ;
        RECT 77.190 156.425 77.440 157.025 ;
        RECT 78.510 156.565 79.720 157.085 ;
        RECT 81.310 157.035 81.540 158.175 ;
        RECT 81.710 157.025 82.040 158.005 ;
        RECT 82.210 157.035 82.420 158.175 ;
        RECT 82.855 157.205 83.185 158.005 ;
        RECT 83.355 157.375 83.685 158.175 ;
        RECT 83.985 157.205 84.315 158.005 ;
        RECT 84.960 157.375 85.210 158.175 ;
        RECT 82.855 157.035 85.290 157.205 ;
        RECT 85.480 157.035 85.650 158.175 ;
        RECT 85.820 157.035 86.160 158.005 ;
        RECT 77.110 155.795 77.440 156.425 ;
        RECT 77.610 155.625 77.820 156.445 ;
        RECT 79.890 156.395 81.100 156.915 ;
        RECT 81.290 156.615 81.620 156.865 ;
        RECT 78.510 155.625 81.100 156.395 ;
        RECT 81.310 155.625 81.540 156.445 ;
        RECT 81.790 156.425 82.040 157.025 ;
        RECT 82.650 156.615 83.000 156.865 ;
        RECT 81.710 155.795 82.040 156.425 ;
        RECT 82.210 155.625 82.420 156.445 ;
        RECT 83.185 156.405 83.355 157.035 ;
        RECT 83.525 156.615 83.855 156.815 ;
        RECT 84.025 156.615 84.355 156.815 ;
        RECT 84.525 156.615 84.945 156.815 ;
        RECT 85.120 156.785 85.290 157.035 ;
        RECT 85.120 156.615 85.815 156.785 ;
        RECT 82.855 155.795 83.355 156.405 ;
        RECT 83.985 156.275 85.210 156.445 ;
        RECT 85.985 156.425 86.160 157.035 ;
        RECT 86.330 157.010 86.620 158.175 ;
        RECT 86.990 157.505 87.270 158.175 ;
        RECT 87.440 157.285 87.740 157.835 ;
        RECT 87.940 157.455 88.270 158.175 ;
        RECT 88.460 157.455 88.920 158.005 ;
        RECT 86.805 156.865 87.070 157.225 ;
        RECT 87.440 157.115 88.380 157.285 ;
        RECT 88.210 156.865 88.380 157.115 ;
        RECT 86.805 156.615 87.480 156.865 ;
        RECT 87.700 156.615 88.040 156.865 ;
        RECT 88.210 156.535 88.500 156.865 ;
        RECT 88.210 156.445 88.380 156.535 ;
        RECT 83.985 155.795 84.315 156.275 ;
        RECT 84.485 155.625 84.710 156.085 ;
        RECT 84.880 155.795 85.210 156.275 ;
        RECT 85.400 155.625 85.650 156.425 ;
        RECT 85.820 155.795 86.160 156.425 ;
        RECT 86.330 155.625 86.620 156.350 ;
        RECT 86.990 156.255 88.380 156.445 ;
        RECT 86.990 155.895 87.320 156.255 ;
        RECT 88.670 156.085 88.920 157.455 ;
        RECT 87.940 155.625 88.190 156.085 ;
        RECT 88.360 155.795 88.920 156.085 ;
        RECT 89.090 157.035 89.430 158.005 ;
        RECT 89.600 157.035 89.770 158.175 ;
        RECT 90.040 157.375 90.290 158.175 ;
        RECT 90.935 157.205 91.265 158.005 ;
        RECT 91.565 157.375 91.895 158.175 ;
        RECT 92.065 157.205 92.395 158.005 ;
        RECT 89.960 157.035 92.395 157.205 ;
        RECT 92.770 157.415 93.285 157.825 ;
        RECT 93.520 157.415 93.690 158.175 ;
        RECT 93.860 157.835 95.890 158.005 ;
        RECT 89.090 156.425 89.265 157.035 ;
        RECT 89.960 156.785 90.130 157.035 ;
        RECT 89.435 156.615 90.130 156.785 ;
        RECT 90.305 156.615 90.725 156.815 ;
        RECT 90.895 156.615 91.225 156.815 ;
        RECT 91.395 156.615 91.725 156.815 ;
        RECT 89.090 155.795 89.430 156.425 ;
        RECT 89.600 155.625 89.850 156.425 ;
        RECT 90.040 156.275 91.265 156.445 ;
        RECT 90.040 155.795 90.370 156.275 ;
        RECT 90.540 155.625 90.765 156.085 ;
        RECT 90.935 155.795 91.265 156.275 ;
        RECT 91.895 156.405 92.065 157.035 ;
        RECT 92.250 156.615 92.600 156.865 ;
        RECT 92.770 156.605 93.110 157.415 ;
        RECT 93.860 157.170 94.030 157.835 ;
        RECT 94.425 157.495 95.550 157.665 ;
        RECT 93.280 156.980 94.030 157.170 ;
        RECT 94.200 157.155 95.210 157.325 ;
        RECT 92.770 156.435 94.000 156.605 ;
        RECT 91.895 155.795 92.395 156.405 ;
        RECT 93.045 155.830 93.290 156.435 ;
        RECT 93.510 155.625 94.020 156.160 ;
        RECT 94.200 155.795 94.390 157.155 ;
        RECT 94.560 156.815 94.835 156.955 ;
        RECT 94.560 156.645 94.840 156.815 ;
        RECT 94.560 155.795 94.835 156.645 ;
        RECT 95.040 156.355 95.210 157.155 ;
        RECT 95.380 156.365 95.550 157.495 ;
        RECT 95.720 156.865 95.890 157.835 ;
        RECT 96.060 157.035 96.230 158.175 ;
        RECT 96.400 157.035 96.735 158.005 ;
        RECT 95.720 156.535 95.915 156.865 ;
        RECT 96.140 156.535 96.395 156.865 ;
        RECT 96.140 156.365 96.310 156.535 ;
        RECT 96.565 156.365 96.735 157.035 ;
        RECT 96.910 157.085 98.120 158.175 ;
        RECT 98.665 157.835 98.920 157.865 ;
        RECT 98.580 157.665 98.920 157.835 ;
        RECT 98.665 157.195 98.920 157.665 ;
        RECT 99.100 157.375 99.385 158.175 ;
        RECT 99.565 157.455 99.895 157.965 ;
        RECT 96.910 156.545 97.430 157.085 ;
        RECT 97.600 156.375 98.120 156.915 ;
        RECT 95.380 156.195 96.310 156.365 ;
        RECT 95.380 156.160 95.555 156.195 ;
        RECT 95.025 155.795 95.555 156.160 ;
        RECT 95.980 155.625 96.310 156.025 ;
        RECT 96.480 155.795 96.735 156.365 ;
        RECT 96.910 155.625 98.120 156.375 ;
        RECT 98.665 156.335 98.845 157.195 ;
        RECT 99.565 156.865 99.815 157.455 ;
        RECT 100.165 157.305 100.335 157.915 ;
        RECT 100.505 157.485 100.835 158.175 ;
        RECT 101.065 157.625 101.305 157.915 ;
        RECT 101.505 157.795 101.925 158.175 ;
        RECT 102.105 157.705 102.735 157.955 ;
        RECT 103.205 157.795 103.535 158.175 ;
        RECT 102.105 157.625 102.275 157.705 ;
        RECT 103.705 157.625 103.875 157.915 ;
        RECT 104.055 157.795 104.435 158.175 ;
        RECT 104.675 157.790 105.505 157.960 ;
        RECT 101.065 157.455 102.275 157.625 ;
        RECT 99.015 156.535 99.815 156.865 ;
        RECT 98.665 155.805 98.920 156.335 ;
        RECT 99.100 155.625 99.385 156.085 ;
        RECT 99.565 155.885 99.815 156.535 ;
        RECT 100.015 157.285 100.335 157.305 ;
        RECT 100.015 157.115 101.935 157.285 ;
        RECT 100.015 156.220 100.205 157.115 ;
        RECT 102.105 156.945 102.275 157.455 ;
        RECT 102.445 157.195 102.965 157.505 ;
        RECT 100.375 156.775 102.275 156.945 ;
        RECT 100.375 156.715 100.705 156.775 ;
        RECT 100.855 156.545 101.185 156.605 ;
        RECT 100.525 156.275 101.185 156.545 ;
        RECT 100.015 155.890 100.335 156.220 ;
        RECT 100.515 155.625 101.175 156.105 ;
        RECT 101.375 156.015 101.545 156.775 ;
        RECT 102.445 156.605 102.625 157.015 ;
        RECT 101.715 156.435 102.045 156.555 ;
        RECT 102.795 156.435 102.965 157.195 ;
        RECT 101.715 156.265 102.965 156.435 ;
        RECT 103.135 157.375 104.505 157.625 ;
        RECT 103.135 156.605 103.325 157.375 ;
        RECT 104.255 157.115 104.505 157.375 ;
        RECT 103.495 156.945 103.745 157.105 ;
        RECT 104.675 156.945 104.845 157.790 ;
        RECT 105.740 157.505 105.910 158.005 ;
        RECT 106.080 157.675 106.410 158.175 ;
        RECT 105.015 157.115 105.515 157.495 ;
        RECT 105.740 157.335 106.435 157.505 ;
        RECT 103.495 156.775 104.845 156.945 ;
        RECT 104.425 156.735 104.845 156.775 ;
        RECT 103.135 156.265 103.555 156.605 ;
        RECT 103.845 156.275 104.255 156.605 ;
        RECT 101.375 155.845 102.225 156.015 ;
        RECT 102.785 155.625 103.105 156.085 ;
        RECT 103.305 155.835 103.555 156.265 ;
        RECT 103.845 155.625 104.255 156.065 ;
        RECT 104.425 156.005 104.595 156.735 ;
        RECT 104.765 156.185 105.115 156.555 ;
        RECT 105.295 156.245 105.515 157.115 ;
        RECT 105.685 156.545 106.095 157.165 ;
        RECT 106.265 156.365 106.435 157.335 ;
        RECT 105.740 156.175 106.435 156.365 ;
        RECT 104.425 155.805 105.440 156.005 ;
        RECT 105.740 155.845 105.910 156.175 ;
        RECT 106.080 155.625 106.410 156.005 ;
        RECT 106.625 155.885 106.850 158.005 ;
        RECT 107.020 157.675 107.350 158.175 ;
        RECT 107.520 157.505 107.690 158.005 ;
        RECT 107.025 157.335 107.690 157.505 ;
        RECT 107.025 156.345 107.255 157.335 ;
        RECT 107.425 156.515 107.775 157.165 ;
        RECT 108.410 157.085 111.000 158.175 ;
        RECT 111.170 157.085 112.380 158.175 ;
        RECT 108.410 156.565 109.620 157.085 ;
        RECT 109.790 156.395 111.000 156.915 ;
        RECT 111.170 156.545 111.690 157.085 ;
        RECT 107.025 156.175 107.690 156.345 ;
        RECT 107.020 155.625 107.350 156.005 ;
        RECT 107.520 155.885 107.690 156.175 ;
        RECT 108.410 155.625 111.000 156.395 ;
        RECT 111.860 156.375 112.380 156.915 ;
        RECT 111.170 155.625 112.380 156.375 ;
        RECT 18.165 155.455 112.465 155.625 ;
        RECT 18.250 154.705 19.460 155.455 ;
        RECT 18.250 154.165 18.770 154.705 ;
        RECT 20.610 154.635 20.820 155.455 ;
        RECT 20.990 154.655 21.320 155.285 ;
        RECT 18.940 153.995 19.460 154.535 ;
        RECT 20.990 154.055 21.240 154.655 ;
        RECT 21.490 154.635 21.720 155.455 ;
        RECT 21.930 154.730 22.220 155.455 ;
        RECT 22.700 154.985 22.870 155.455 ;
        RECT 23.040 154.805 23.370 155.285 ;
        RECT 23.540 154.985 23.710 155.455 ;
        RECT 23.880 154.805 24.210 155.285 ;
        RECT 22.445 154.635 24.210 154.805 ;
        RECT 24.380 154.645 24.550 155.455 ;
        RECT 24.750 155.075 25.820 155.245 ;
        RECT 24.750 154.720 25.070 155.075 ;
        RECT 21.410 154.215 21.740 154.465 ;
        RECT 22.445 154.085 22.855 154.635 ;
        RECT 24.745 154.465 25.070 154.720 ;
        RECT 23.040 154.255 25.070 154.465 ;
        RECT 24.725 154.245 25.070 154.255 ;
        RECT 25.240 154.505 25.480 154.905 ;
        RECT 25.650 154.845 25.820 155.075 ;
        RECT 25.990 155.015 26.180 155.455 ;
        RECT 26.350 155.005 27.300 155.285 ;
        RECT 27.520 155.095 27.870 155.265 ;
        RECT 25.650 154.675 26.180 154.845 ;
        RECT 18.250 152.905 19.460 153.995 ;
        RECT 20.610 152.905 20.820 154.045 ;
        RECT 20.990 153.075 21.320 154.055 ;
        RECT 21.490 152.905 21.720 154.045 ;
        RECT 21.930 152.905 22.220 154.070 ;
        RECT 22.445 153.915 24.170 154.085 ;
        RECT 22.700 152.905 22.870 153.745 ;
        RECT 23.080 153.075 23.330 153.915 ;
        RECT 23.540 152.905 23.710 153.745 ;
        RECT 23.880 153.075 24.170 153.915 ;
        RECT 24.380 152.905 24.550 153.965 ;
        RECT 24.725 153.625 24.895 154.245 ;
        RECT 25.240 154.135 25.780 154.505 ;
        RECT 25.960 154.395 26.180 154.675 ;
        RECT 26.350 154.225 26.520 155.005 ;
        RECT 26.115 154.055 26.520 154.225 ;
        RECT 26.690 154.215 27.040 154.835 ;
        RECT 26.115 153.965 26.285 154.055 ;
        RECT 27.210 154.045 27.420 154.835 ;
        RECT 25.065 153.795 26.285 153.965 ;
        RECT 26.745 153.885 27.420 154.045 ;
        RECT 24.725 153.455 25.525 153.625 ;
        RECT 24.845 152.905 25.175 153.285 ;
        RECT 25.355 153.165 25.525 153.455 ;
        RECT 26.115 153.415 26.285 153.795 ;
        RECT 26.455 153.875 27.420 153.885 ;
        RECT 27.610 154.705 27.870 155.095 ;
        RECT 28.080 154.995 28.410 155.455 ;
        RECT 29.285 155.065 30.140 155.235 ;
        RECT 30.345 155.065 30.840 155.235 ;
        RECT 31.010 155.095 31.340 155.455 ;
        RECT 27.610 154.015 27.780 154.705 ;
        RECT 27.950 154.355 28.120 154.535 ;
        RECT 28.290 154.525 29.080 154.775 ;
        RECT 29.285 154.355 29.455 155.065 ;
        RECT 29.625 154.555 29.980 154.775 ;
        RECT 27.950 154.185 29.640 154.355 ;
        RECT 26.455 153.585 26.915 153.875 ;
        RECT 27.610 153.845 29.110 154.015 ;
        RECT 27.610 153.705 27.780 153.845 ;
        RECT 27.220 153.535 27.780 153.705 ;
        RECT 25.695 152.905 25.945 153.365 ;
        RECT 26.115 153.075 26.985 153.415 ;
        RECT 27.220 153.075 27.390 153.535 ;
        RECT 28.225 153.505 29.300 153.675 ;
        RECT 27.560 152.905 27.930 153.365 ;
        RECT 28.225 153.165 28.395 153.505 ;
        RECT 28.565 152.905 28.895 153.335 ;
        RECT 29.130 153.165 29.300 153.505 ;
        RECT 29.470 153.405 29.640 154.185 ;
        RECT 29.810 153.965 29.980 154.555 ;
        RECT 30.150 154.155 30.500 154.775 ;
        RECT 29.810 153.575 30.275 153.965 ;
        RECT 30.670 153.705 30.840 155.065 ;
        RECT 31.010 153.875 31.470 154.925 ;
        RECT 30.445 153.535 30.840 153.705 ;
        RECT 30.445 153.405 30.615 153.535 ;
        RECT 29.470 153.075 30.150 153.405 ;
        RECT 30.365 153.075 30.615 153.405 ;
        RECT 30.785 152.905 31.035 153.365 ;
        RECT 31.205 153.090 31.530 153.875 ;
        RECT 31.700 153.075 31.870 155.195 ;
        RECT 32.040 155.075 32.370 155.455 ;
        RECT 32.540 154.905 32.795 155.195 ;
        RECT 32.045 154.735 32.795 154.905 ;
        RECT 32.045 153.745 32.275 154.735 ;
        RECT 33.930 154.635 34.160 155.455 ;
        RECT 34.330 154.655 34.660 155.285 ;
        RECT 32.445 153.915 32.795 154.565 ;
        RECT 33.910 154.215 34.240 154.465 ;
        RECT 34.410 154.055 34.660 154.655 ;
        RECT 34.830 154.635 35.040 155.455 ;
        RECT 35.360 154.905 35.530 155.285 ;
        RECT 35.710 155.075 36.040 155.455 ;
        RECT 35.360 154.735 36.025 154.905 ;
        RECT 36.220 154.780 36.480 155.285 ;
        RECT 35.290 154.185 35.630 154.555 ;
        RECT 35.855 154.480 36.025 154.735 ;
        RECT 32.045 153.575 32.795 153.745 ;
        RECT 32.040 152.905 32.370 153.405 ;
        RECT 32.540 153.075 32.795 153.575 ;
        RECT 33.930 152.905 34.160 154.045 ;
        RECT 34.330 153.075 34.660 154.055 ;
        RECT 35.855 154.150 36.130 154.480 ;
        RECT 34.830 152.905 35.040 154.045 ;
        RECT 35.855 154.005 36.025 154.150 ;
        RECT 35.350 153.835 36.025 154.005 ;
        RECT 36.300 153.980 36.480 154.780 ;
        RECT 36.650 154.705 37.860 155.455 ;
        RECT 38.120 154.905 38.290 155.285 ;
        RECT 38.505 155.075 38.835 155.455 ;
        RECT 38.120 154.735 38.835 154.905 ;
        RECT 35.350 153.075 35.530 153.835 ;
        RECT 35.710 152.905 36.040 153.665 ;
        RECT 36.210 153.075 36.480 153.980 ;
        RECT 36.650 153.995 37.170 154.535 ;
        RECT 37.340 154.165 37.860 154.705 ;
        RECT 38.030 154.185 38.385 154.555 ;
        RECT 38.665 154.545 38.835 154.735 ;
        RECT 39.005 154.710 39.260 155.285 ;
        RECT 38.665 154.215 38.920 154.545 ;
        RECT 38.665 154.005 38.835 154.215 ;
        RECT 36.650 152.905 37.860 153.995 ;
        RECT 38.120 153.835 38.835 154.005 ;
        RECT 39.090 153.980 39.260 154.710 ;
        RECT 39.435 154.615 39.695 155.455 ;
        RECT 39.870 154.780 40.140 155.125 ;
        RECT 40.330 155.055 40.710 155.455 ;
        RECT 40.880 154.885 41.050 155.235 ;
        RECT 41.220 155.055 41.550 155.455 ;
        RECT 41.750 154.885 41.920 155.235 ;
        RECT 42.120 154.955 42.450 155.455 ;
        RECT 38.120 153.075 38.290 153.835 ;
        RECT 38.505 152.905 38.835 153.665 ;
        RECT 39.005 153.075 39.260 153.980 ;
        RECT 39.435 152.905 39.695 154.055 ;
        RECT 39.870 154.045 40.040 154.780 ;
        RECT 40.310 154.715 41.920 154.885 ;
        RECT 40.310 154.545 40.480 154.715 ;
        RECT 40.210 154.215 40.480 154.545 ;
        RECT 40.650 154.215 41.055 154.545 ;
        RECT 40.310 154.045 40.480 154.215 ;
        RECT 41.225 154.095 41.935 154.545 ;
        RECT 42.105 154.215 42.455 154.785 ;
        RECT 42.905 154.645 43.150 155.250 ;
        RECT 43.370 154.920 43.880 155.455 ;
        RECT 42.630 154.475 43.860 154.645 ;
        RECT 39.870 153.075 40.140 154.045 ;
        RECT 40.310 153.875 41.035 154.045 ;
        RECT 41.225 153.925 41.940 154.095 ;
        RECT 40.865 153.755 41.035 153.875 ;
        RECT 42.135 153.755 42.455 154.045 ;
        RECT 40.350 152.905 40.630 153.705 ;
        RECT 40.865 153.585 42.455 153.755 ;
        RECT 42.630 153.665 42.970 154.475 ;
        RECT 43.140 153.910 43.890 154.100 ;
        RECT 40.800 153.125 42.455 153.415 ;
        RECT 42.630 153.255 43.145 153.665 ;
        RECT 43.380 152.905 43.550 153.665 ;
        RECT 43.720 153.245 43.890 153.910 ;
        RECT 44.060 153.925 44.250 155.285 ;
        RECT 44.420 155.115 44.695 155.285 ;
        RECT 44.420 154.945 44.700 155.115 ;
        RECT 44.420 154.125 44.695 154.945 ;
        RECT 44.885 154.920 45.415 155.285 ;
        RECT 45.840 155.055 46.170 155.455 ;
        RECT 45.240 154.885 45.415 154.920 ;
        RECT 44.900 153.925 45.070 154.725 ;
        RECT 44.060 153.755 45.070 153.925 ;
        RECT 45.240 154.715 46.170 154.885 ;
        RECT 46.340 154.715 46.595 155.285 ;
        RECT 47.690 154.730 47.980 155.455 ;
        RECT 45.240 153.585 45.410 154.715 ;
        RECT 46.000 154.545 46.170 154.715 ;
        RECT 44.285 153.415 45.410 153.585 ;
        RECT 45.580 154.215 45.775 154.545 ;
        RECT 46.000 154.215 46.255 154.545 ;
        RECT 45.580 153.245 45.750 154.215 ;
        RECT 46.425 154.045 46.595 154.715 ;
        RECT 48.150 154.655 48.490 155.285 ;
        RECT 48.660 154.655 48.910 155.455 ;
        RECT 49.100 154.805 49.430 155.285 ;
        RECT 49.600 154.995 49.825 155.455 ;
        RECT 49.995 154.805 50.325 155.285 ;
        RECT 48.150 154.605 48.380 154.655 ;
        RECT 49.100 154.635 50.325 154.805 ;
        RECT 50.955 154.675 51.455 155.285 ;
        RECT 52.865 154.825 53.150 155.285 ;
        RECT 53.320 154.995 53.590 155.455 ;
        RECT 43.720 153.075 45.750 153.245 ;
        RECT 45.920 152.905 46.090 154.045 ;
        RECT 46.260 153.075 46.595 154.045 ;
        RECT 47.690 152.905 47.980 154.070 ;
        RECT 48.150 154.045 48.325 154.605 ;
        RECT 48.495 154.295 49.190 154.465 ;
        RECT 49.020 154.045 49.190 154.295 ;
        RECT 49.365 154.265 49.785 154.465 ;
        RECT 49.955 154.265 50.285 154.465 ;
        RECT 50.455 154.265 50.785 154.465 ;
        RECT 50.955 154.045 51.125 154.675 ;
        RECT 52.865 154.655 53.820 154.825 ;
        RECT 51.310 154.215 51.660 154.465 ;
        RECT 48.150 153.075 48.490 154.045 ;
        RECT 48.660 152.905 48.830 154.045 ;
        RECT 49.020 153.875 51.455 154.045 ;
        RECT 52.750 153.925 53.440 154.485 ;
        RECT 49.100 152.905 49.350 153.705 ;
        RECT 49.995 153.075 50.325 153.875 ;
        RECT 50.625 152.905 50.955 153.705 ;
        RECT 51.125 153.075 51.455 153.875 ;
        RECT 53.610 153.755 53.820 154.655 ;
        RECT 52.865 153.535 53.820 153.755 ;
        RECT 53.990 154.485 54.390 155.285 ;
        RECT 54.580 154.825 54.860 155.285 ;
        RECT 55.380 154.995 55.705 155.455 ;
        RECT 54.580 154.655 55.705 154.825 ;
        RECT 55.875 154.715 56.260 155.285 ;
        RECT 55.255 154.545 55.705 154.655 ;
        RECT 53.990 153.925 55.085 154.485 ;
        RECT 55.255 154.215 55.810 154.545 ;
        RECT 52.865 153.075 53.150 153.535 ;
        RECT 53.320 152.905 53.590 153.365 ;
        RECT 53.990 153.075 54.390 153.925 ;
        RECT 55.255 153.755 55.705 154.215 ;
        RECT 55.980 154.045 56.260 154.715 ;
        RECT 54.580 153.535 55.705 153.755 ;
        RECT 54.580 153.075 54.860 153.535 ;
        RECT 55.380 152.905 55.705 153.365 ;
        RECT 55.875 153.075 56.260 154.045 ;
        RECT 57.350 154.655 57.690 155.285 ;
        RECT 57.860 154.655 58.110 155.455 ;
        RECT 58.300 154.805 58.630 155.285 ;
        RECT 58.800 154.995 59.025 155.455 ;
        RECT 59.195 154.805 59.525 155.285 ;
        RECT 57.350 154.045 57.525 154.655 ;
        RECT 58.300 154.635 59.525 154.805 ;
        RECT 60.155 154.675 60.655 155.285 ;
        RECT 61.035 154.745 61.290 155.275 ;
        RECT 61.460 154.995 61.765 155.455 ;
        RECT 62.010 155.075 63.080 155.245 ;
        RECT 57.695 154.295 58.390 154.465 ;
        RECT 58.220 154.045 58.390 154.295 ;
        RECT 58.565 154.265 58.985 154.465 ;
        RECT 59.155 154.265 59.485 154.465 ;
        RECT 59.655 154.265 59.985 154.465 ;
        RECT 60.155 154.045 60.325 154.675 ;
        RECT 60.510 154.215 60.860 154.465 ;
        RECT 61.035 154.095 61.245 154.745 ;
        RECT 62.010 154.720 62.330 155.075 ;
        RECT 62.005 154.545 62.330 154.720 ;
        RECT 61.415 154.245 62.330 154.545 ;
        RECT 62.500 154.505 62.740 154.905 ;
        RECT 62.910 154.845 63.080 155.075 ;
        RECT 63.250 155.015 63.440 155.455 ;
        RECT 63.610 155.005 64.560 155.285 ;
        RECT 64.780 155.095 65.130 155.265 ;
        RECT 62.910 154.675 63.440 154.845 ;
        RECT 61.415 154.215 62.155 154.245 ;
        RECT 57.350 153.075 57.690 154.045 ;
        RECT 57.860 152.905 58.030 154.045 ;
        RECT 58.220 153.875 60.655 154.045 ;
        RECT 58.300 152.905 58.550 153.705 ;
        RECT 59.195 153.075 59.525 153.875 ;
        RECT 59.825 152.905 60.155 153.705 ;
        RECT 60.325 153.075 60.655 153.875 ;
        RECT 61.035 153.215 61.290 154.095 ;
        RECT 61.460 152.905 61.765 154.045 ;
        RECT 61.985 153.625 62.155 154.215 ;
        RECT 62.500 154.135 63.040 154.505 ;
        RECT 63.220 154.395 63.440 154.675 ;
        RECT 63.610 154.225 63.780 155.005 ;
        RECT 63.375 154.055 63.780 154.225 ;
        RECT 63.950 154.215 64.300 154.835 ;
        RECT 63.375 153.965 63.545 154.055 ;
        RECT 64.470 154.045 64.680 154.835 ;
        RECT 62.325 153.795 63.545 153.965 ;
        RECT 64.005 153.885 64.680 154.045 ;
        RECT 61.985 153.455 62.785 153.625 ;
        RECT 62.105 152.905 62.435 153.285 ;
        RECT 62.615 153.165 62.785 153.455 ;
        RECT 63.375 153.415 63.545 153.795 ;
        RECT 63.715 153.875 64.680 153.885 ;
        RECT 64.870 154.705 65.130 155.095 ;
        RECT 65.340 154.995 65.670 155.455 ;
        RECT 66.545 155.065 67.400 155.235 ;
        RECT 67.605 155.065 68.100 155.235 ;
        RECT 68.270 155.095 68.600 155.455 ;
        RECT 64.870 154.015 65.040 154.705 ;
        RECT 65.210 154.355 65.380 154.535 ;
        RECT 65.550 154.525 66.340 154.775 ;
        RECT 66.545 154.355 66.715 155.065 ;
        RECT 66.885 154.555 67.240 154.775 ;
        RECT 65.210 154.185 66.900 154.355 ;
        RECT 63.715 153.585 64.175 153.875 ;
        RECT 64.870 153.845 66.370 154.015 ;
        RECT 64.870 153.705 65.040 153.845 ;
        RECT 64.480 153.535 65.040 153.705 ;
        RECT 62.955 152.905 63.205 153.365 ;
        RECT 63.375 153.075 64.245 153.415 ;
        RECT 64.480 153.075 64.650 153.535 ;
        RECT 65.485 153.505 66.560 153.675 ;
        RECT 64.820 152.905 65.190 153.365 ;
        RECT 65.485 153.165 65.655 153.505 ;
        RECT 65.825 152.905 66.155 153.335 ;
        RECT 66.390 153.165 66.560 153.505 ;
        RECT 66.730 153.405 66.900 154.185 ;
        RECT 67.070 153.965 67.240 154.555 ;
        RECT 67.410 154.155 67.760 154.775 ;
        RECT 67.070 153.575 67.535 153.965 ;
        RECT 67.930 153.705 68.100 155.065 ;
        RECT 68.270 153.875 68.730 154.925 ;
        RECT 67.705 153.535 68.100 153.705 ;
        RECT 67.705 153.405 67.875 153.535 ;
        RECT 66.730 153.075 67.410 153.405 ;
        RECT 67.625 153.075 67.875 153.405 ;
        RECT 68.045 152.905 68.295 153.365 ;
        RECT 68.465 153.090 68.790 153.875 ;
        RECT 68.960 153.075 69.130 155.195 ;
        RECT 69.300 155.075 69.630 155.455 ;
        RECT 69.800 154.905 70.055 155.195 ;
        RECT 69.305 154.735 70.055 154.905 ;
        RECT 69.305 153.745 69.535 154.735 ;
        RECT 70.690 154.685 73.280 155.455 ;
        RECT 73.450 154.730 73.740 155.455 ;
        RECT 75.205 154.745 75.460 155.275 ;
        RECT 75.640 154.995 75.925 155.455 ;
        RECT 69.705 153.915 70.055 154.565 ;
        RECT 70.690 153.995 71.900 154.515 ;
        RECT 72.070 154.165 73.280 154.685 ;
        RECT 69.305 153.575 70.055 153.745 ;
        RECT 69.300 152.905 69.630 153.405 ;
        RECT 69.800 153.075 70.055 153.575 ;
        RECT 70.690 152.905 73.280 153.995 ;
        RECT 73.450 152.905 73.740 154.070 ;
        RECT 75.205 153.885 75.385 154.745 ;
        RECT 76.105 154.545 76.355 155.195 ;
        RECT 75.555 154.215 76.355 154.545 ;
        RECT 75.205 153.415 75.460 153.885 ;
        RECT 75.120 153.245 75.460 153.415 ;
        RECT 75.205 153.215 75.460 153.245 ;
        RECT 75.640 152.905 75.925 153.705 ;
        RECT 76.105 153.625 76.355 154.215 ;
        RECT 76.555 154.860 76.875 155.190 ;
        RECT 77.055 154.975 77.715 155.455 ;
        RECT 77.915 155.065 78.765 155.235 ;
        RECT 76.555 153.965 76.745 154.860 ;
        RECT 77.065 154.535 77.725 154.805 ;
        RECT 77.395 154.475 77.725 154.535 ;
        RECT 76.915 154.305 77.245 154.365 ;
        RECT 77.915 154.305 78.085 155.065 ;
        RECT 79.325 154.995 79.645 155.455 ;
        RECT 79.845 154.815 80.095 155.245 ;
        RECT 80.385 155.015 80.795 155.455 ;
        RECT 80.965 155.075 81.980 155.275 ;
        RECT 78.255 154.645 79.505 154.815 ;
        RECT 78.255 154.525 78.585 154.645 ;
        RECT 76.915 154.135 78.815 154.305 ;
        RECT 76.555 153.795 78.475 153.965 ;
        RECT 76.555 153.775 76.875 153.795 ;
        RECT 76.105 153.115 76.435 153.625 ;
        RECT 76.705 153.165 76.875 153.775 ;
        RECT 78.645 153.625 78.815 154.135 ;
        RECT 78.985 154.065 79.165 154.475 ;
        RECT 79.335 153.885 79.505 154.645 ;
        RECT 77.045 152.905 77.375 153.595 ;
        RECT 77.605 153.455 78.815 153.625 ;
        RECT 78.985 153.575 79.505 153.885 ;
        RECT 79.675 154.475 80.095 154.815 ;
        RECT 80.385 154.475 80.795 154.805 ;
        RECT 79.675 153.705 79.865 154.475 ;
        RECT 80.965 154.345 81.135 155.075 ;
        RECT 82.280 154.905 82.450 155.235 ;
        RECT 82.620 155.075 82.950 155.455 ;
        RECT 81.305 154.525 81.655 154.895 ;
        RECT 80.965 154.305 81.385 154.345 ;
        RECT 80.035 154.135 81.385 154.305 ;
        RECT 80.035 153.975 80.285 154.135 ;
        RECT 80.795 153.705 81.045 153.965 ;
        RECT 79.675 153.455 81.045 153.705 ;
        RECT 77.605 153.165 77.845 153.455 ;
        RECT 78.645 153.375 78.815 153.455 ;
        RECT 78.045 152.905 78.465 153.285 ;
        RECT 78.645 153.125 79.275 153.375 ;
        RECT 79.745 152.905 80.075 153.285 ;
        RECT 80.245 153.165 80.415 153.455 ;
        RECT 81.215 153.290 81.385 154.135 ;
        RECT 81.835 153.965 82.055 154.835 ;
        RECT 82.280 154.715 82.975 154.905 ;
        RECT 81.555 153.585 82.055 153.965 ;
        RECT 82.225 153.915 82.635 154.535 ;
        RECT 82.805 153.745 82.975 154.715 ;
        RECT 82.280 153.575 82.975 153.745 ;
        RECT 80.595 152.905 80.975 153.285 ;
        RECT 81.215 153.120 82.045 153.290 ;
        RECT 82.280 153.075 82.450 153.575 ;
        RECT 82.620 152.905 82.950 153.405 ;
        RECT 83.165 153.075 83.390 155.195 ;
        RECT 83.560 155.075 83.890 155.455 ;
        RECT 84.060 154.905 84.230 155.195 ;
        RECT 83.565 154.735 84.230 154.905 ;
        RECT 83.565 153.745 83.795 154.735 ;
        RECT 85.685 154.645 85.930 155.250 ;
        RECT 86.150 154.920 86.660 155.455 ;
        RECT 83.965 153.915 84.315 154.565 ;
        RECT 85.410 154.475 86.640 154.645 ;
        RECT 83.565 153.575 84.230 153.745 ;
        RECT 83.560 152.905 83.890 153.405 ;
        RECT 84.060 153.075 84.230 153.575 ;
        RECT 85.410 153.665 85.750 154.475 ;
        RECT 85.920 153.910 86.670 154.100 ;
        RECT 85.410 153.255 85.925 153.665 ;
        RECT 86.160 152.905 86.330 153.665 ;
        RECT 86.500 153.245 86.670 153.910 ;
        RECT 86.840 153.925 87.030 155.285 ;
        RECT 87.200 154.435 87.475 155.285 ;
        RECT 87.665 154.920 88.195 155.285 ;
        RECT 88.620 155.055 88.950 155.455 ;
        RECT 88.020 154.885 88.195 154.920 ;
        RECT 87.200 154.265 87.480 154.435 ;
        RECT 87.200 154.125 87.475 154.265 ;
        RECT 87.680 153.925 87.850 154.725 ;
        RECT 86.840 153.755 87.850 153.925 ;
        RECT 88.020 154.715 88.950 154.885 ;
        RECT 89.120 154.715 89.375 155.285 ;
        RECT 88.020 153.585 88.190 154.715 ;
        RECT 88.780 154.545 88.950 154.715 ;
        RECT 87.065 153.415 88.190 153.585 ;
        RECT 88.360 154.215 88.555 154.545 ;
        RECT 88.780 154.215 89.035 154.545 ;
        RECT 88.360 153.245 88.530 154.215 ;
        RECT 89.205 154.045 89.375 154.715 ;
        RECT 89.925 154.745 90.180 155.275 ;
        RECT 90.360 154.995 90.645 155.455 ;
        RECT 89.925 154.095 90.105 154.745 ;
        RECT 90.825 154.545 91.075 155.195 ;
        RECT 90.275 154.215 91.075 154.545 ;
        RECT 86.500 153.075 88.530 153.245 ;
        RECT 88.700 152.905 88.870 154.045 ;
        RECT 89.040 153.075 89.375 154.045 ;
        RECT 89.840 153.925 90.105 154.095 ;
        RECT 89.925 153.885 90.105 153.925 ;
        RECT 89.925 153.215 90.180 153.885 ;
        RECT 90.360 152.905 90.645 153.705 ;
        RECT 90.825 153.625 91.075 154.215 ;
        RECT 91.275 154.860 91.595 155.190 ;
        RECT 91.775 154.975 92.435 155.455 ;
        RECT 92.635 155.065 93.485 155.235 ;
        RECT 91.275 153.965 91.465 154.860 ;
        RECT 91.785 154.535 92.445 154.805 ;
        RECT 92.115 154.475 92.445 154.535 ;
        RECT 91.635 154.305 91.965 154.365 ;
        RECT 92.635 154.305 92.805 155.065 ;
        RECT 94.045 154.995 94.365 155.455 ;
        RECT 94.565 154.815 94.815 155.245 ;
        RECT 95.105 155.015 95.515 155.455 ;
        RECT 95.685 155.075 96.700 155.275 ;
        RECT 92.975 154.645 94.225 154.815 ;
        RECT 92.975 154.525 93.305 154.645 ;
        RECT 91.635 154.135 93.535 154.305 ;
        RECT 91.275 153.795 93.195 153.965 ;
        RECT 91.275 153.775 91.595 153.795 ;
        RECT 90.825 153.115 91.155 153.625 ;
        RECT 91.425 153.165 91.595 153.775 ;
        RECT 93.365 153.625 93.535 154.135 ;
        RECT 93.705 154.065 93.885 154.475 ;
        RECT 94.055 153.885 94.225 154.645 ;
        RECT 91.765 152.905 92.095 153.595 ;
        RECT 92.325 153.455 93.535 153.625 ;
        RECT 93.705 153.575 94.225 153.885 ;
        RECT 94.395 154.475 94.815 154.815 ;
        RECT 95.105 154.475 95.515 154.805 ;
        RECT 94.395 153.705 94.585 154.475 ;
        RECT 95.685 154.345 95.855 155.075 ;
        RECT 97.000 154.905 97.170 155.235 ;
        RECT 97.340 155.075 97.670 155.455 ;
        RECT 96.025 154.525 96.375 154.895 ;
        RECT 95.685 154.305 96.105 154.345 ;
        RECT 94.755 154.135 96.105 154.305 ;
        RECT 94.755 153.975 95.005 154.135 ;
        RECT 95.515 153.705 95.765 153.965 ;
        RECT 94.395 153.455 95.765 153.705 ;
        RECT 92.325 153.165 92.565 153.455 ;
        RECT 93.365 153.375 93.535 153.455 ;
        RECT 92.765 152.905 93.185 153.285 ;
        RECT 93.365 153.125 93.995 153.375 ;
        RECT 94.465 152.905 94.795 153.285 ;
        RECT 94.965 153.165 95.135 153.455 ;
        RECT 95.935 153.290 96.105 154.135 ;
        RECT 96.555 153.965 96.775 154.835 ;
        RECT 97.000 154.715 97.695 154.905 ;
        RECT 96.275 153.585 96.775 153.965 ;
        RECT 96.945 153.915 97.355 154.535 ;
        RECT 97.525 153.745 97.695 154.715 ;
        RECT 97.000 153.575 97.695 153.745 ;
        RECT 95.315 152.905 95.695 153.285 ;
        RECT 95.935 153.120 96.765 153.290 ;
        RECT 97.000 153.075 97.170 153.575 ;
        RECT 97.340 152.905 97.670 153.405 ;
        RECT 97.885 153.075 98.110 155.195 ;
        RECT 98.280 155.075 98.610 155.455 ;
        RECT 98.780 154.905 98.950 155.195 ;
        RECT 98.285 154.735 98.950 154.905 ;
        RECT 98.285 153.745 98.515 154.735 ;
        RECT 99.210 154.730 99.500 155.455 ;
        RECT 100.595 154.905 100.850 155.195 ;
        RECT 101.020 155.075 101.350 155.455 ;
        RECT 100.595 154.735 101.345 154.905 ;
        RECT 98.685 153.915 99.035 154.565 ;
        RECT 98.285 153.575 98.950 153.745 ;
        RECT 98.280 152.905 98.610 153.405 ;
        RECT 98.780 153.075 98.950 153.575 ;
        RECT 99.210 152.905 99.500 154.070 ;
        RECT 100.595 153.915 100.945 154.565 ;
        RECT 101.115 153.745 101.345 154.735 ;
        RECT 100.595 153.575 101.345 153.745 ;
        RECT 100.595 153.075 100.850 153.575 ;
        RECT 101.020 152.905 101.350 153.405 ;
        RECT 101.520 153.075 101.690 155.195 ;
        RECT 102.050 155.095 102.380 155.455 ;
        RECT 102.550 155.065 103.045 155.235 ;
        RECT 103.250 155.065 104.105 155.235 ;
        RECT 101.920 153.875 102.380 154.925 ;
        RECT 101.860 153.090 102.185 153.875 ;
        RECT 102.550 153.705 102.720 155.065 ;
        RECT 102.890 154.155 103.240 154.775 ;
        RECT 103.410 154.555 103.765 154.775 ;
        RECT 103.410 153.965 103.580 154.555 ;
        RECT 103.935 154.355 104.105 155.065 ;
        RECT 104.980 154.995 105.310 155.455 ;
        RECT 105.520 155.095 105.870 155.265 ;
        RECT 104.310 154.525 105.100 154.775 ;
        RECT 105.520 154.705 105.780 155.095 ;
        RECT 106.090 155.005 107.040 155.285 ;
        RECT 107.210 155.015 107.400 155.455 ;
        RECT 107.570 155.075 108.640 155.245 ;
        RECT 105.270 154.355 105.440 154.535 ;
        RECT 102.550 153.535 102.945 153.705 ;
        RECT 103.115 153.575 103.580 153.965 ;
        RECT 103.750 154.185 105.440 154.355 ;
        RECT 102.775 153.405 102.945 153.535 ;
        RECT 103.750 153.405 103.920 154.185 ;
        RECT 105.610 154.015 105.780 154.705 ;
        RECT 104.280 153.845 105.780 154.015 ;
        RECT 105.970 154.045 106.180 154.835 ;
        RECT 106.350 154.215 106.700 154.835 ;
        RECT 106.870 154.225 107.040 155.005 ;
        RECT 107.570 154.845 107.740 155.075 ;
        RECT 107.210 154.675 107.740 154.845 ;
        RECT 107.210 154.395 107.430 154.675 ;
        RECT 107.910 154.505 108.150 154.905 ;
        RECT 106.870 154.055 107.275 154.225 ;
        RECT 107.610 154.135 108.150 154.505 ;
        RECT 108.320 154.720 108.640 155.075 ;
        RECT 108.320 154.465 108.645 154.720 ;
        RECT 108.840 154.645 109.010 155.455 ;
        RECT 109.180 154.805 109.510 155.285 ;
        RECT 109.680 154.985 109.850 155.455 ;
        RECT 110.020 154.805 110.350 155.285 ;
        RECT 110.520 154.985 110.690 155.455 ;
        RECT 109.180 154.635 110.945 154.805 ;
        RECT 111.170 154.705 112.380 155.455 ;
        RECT 108.320 154.255 110.350 154.465 ;
        RECT 108.320 154.245 108.665 154.255 ;
        RECT 105.970 153.885 106.645 154.045 ;
        RECT 107.105 153.965 107.275 154.055 ;
        RECT 105.970 153.875 106.935 153.885 ;
        RECT 105.610 153.705 105.780 153.845 ;
        RECT 102.355 152.905 102.605 153.365 ;
        RECT 102.775 153.075 103.025 153.405 ;
        RECT 103.240 153.075 103.920 153.405 ;
        RECT 104.090 153.505 105.165 153.675 ;
        RECT 105.610 153.535 106.170 153.705 ;
        RECT 106.475 153.585 106.935 153.875 ;
        RECT 107.105 153.795 108.325 153.965 ;
        RECT 104.090 153.165 104.260 153.505 ;
        RECT 104.495 152.905 104.825 153.335 ;
        RECT 104.995 153.165 105.165 153.505 ;
        RECT 105.460 152.905 105.830 153.365 ;
        RECT 106.000 153.075 106.170 153.535 ;
        RECT 107.105 153.415 107.275 153.795 ;
        RECT 108.495 153.625 108.665 154.245 ;
        RECT 110.535 154.085 110.945 154.635 ;
        RECT 106.405 153.075 107.275 153.415 ;
        RECT 107.865 153.455 108.665 153.625 ;
        RECT 107.445 152.905 107.695 153.365 ;
        RECT 107.865 153.165 108.035 153.455 ;
        RECT 108.215 152.905 108.545 153.285 ;
        RECT 108.840 152.905 109.010 153.965 ;
        RECT 109.220 153.915 110.945 154.085 ;
        RECT 111.170 153.995 111.690 154.535 ;
        RECT 111.860 154.165 112.380 154.705 ;
        RECT 109.220 153.075 109.510 153.915 ;
        RECT 109.680 152.905 109.850 153.745 ;
        RECT 110.060 153.075 110.310 153.915 ;
        RECT 110.520 152.905 110.690 153.745 ;
        RECT 111.170 152.905 112.380 153.995 ;
        RECT 18.165 152.735 112.465 152.905 ;
        RECT 18.250 151.645 19.460 152.735 ;
        RECT 20.095 152.300 25.440 152.735 ;
        RECT 18.250 150.935 18.770 151.475 ;
        RECT 18.940 151.105 19.460 151.645 ;
        RECT 21.685 151.050 22.035 152.300 ;
        RECT 18.250 150.185 19.460 150.935 ;
        RECT 23.515 150.730 23.855 151.560 ;
        RECT 25.615 151.545 25.870 152.425 ;
        RECT 26.040 151.595 26.345 152.735 ;
        RECT 26.685 152.355 27.015 152.735 ;
        RECT 27.195 152.185 27.365 152.475 ;
        RECT 27.535 152.275 27.785 152.735 ;
        RECT 26.565 152.015 27.365 152.185 ;
        RECT 27.955 152.225 28.825 152.565 ;
        RECT 25.615 150.895 25.825 151.545 ;
        RECT 26.565 151.425 26.735 152.015 ;
        RECT 27.955 151.845 28.125 152.225 ;
        RECT 29.060 152.105 29.230 152.565 ;
        RECT 29.400 152.275 29.770 152.735 ;
        RECT 30.065 152.135 30.235 152.475 ;
        RECT 30.405 152.305 30.735 152.735 ;
        RECT 30.970 152.135 31.140 152.475 ;
        RECT 26.905 151.675 28.125 151.845 ;
        RECT 28.295 151.765 28.755 152.055 ;
        RECT 29.060 151.935 29.620 152.105 ;
        RECT 30.065 151.965 31.140 152.135 ;
        RECT 31.310 152.235 31.990 152.565 ;
        RECT 32.205 152.235 32.455 152.565 ;
        RECT 32.625 152.275 32.875 152.735 ;
        RECT 29.450 151.795 29.620 151.935 ;
        RECT 28.295 151.755 29.260 151.765 ;
        RECT 27.955 151.585 28.125 151.675 ;
        RECT 28.585 151.595 29.260 151.755 ;
        RECT 25.995 151.395 26.735 151.425 ;
        RECT 25.995 151.095 26.910 151.395 ;
        RECT 26.585 150.920 26.910 151.095 ;
        RECT 20.095 150.185 25.440 150.730 ;
        RECT 25.615 150.365 25.870 150.895 ;
        RECT 26.040 150.185 26.345 150.645 ;
        RECT 26.590 150.565 26.910 150.920 ;
        RECT 27.080 151.135 27.620 151.505 ;
        RECT 27.955 151.415 28.360 151.585 ;
        RECT 27.080 150.735 27.320 151.135 ;
        RECT 27.800 150.965 28.020 151.245 ;
        RECT 27.490 150.795 28.020 150.965 ;
        RECT 27.490 150.565 27.660 150.795 ;
        RECT 28.190 150.635 28.360 151.415 ;
        RECT 28.530 150.805 28.880 151.425 ;
        RECT 29.050 150.805 29.260 151.595 ;
        RECT 29.450 151.625 30.950 151.795 ;
        RECT 29.450 150.935 29.620 151.625 ;
        RECT 31.310 151.455 31.480 152.235 ;
        RECT 32.285 152.105 32.455 152.235 ;
        RECT 29.790 151.285 31.480 151.455 ;
        RECT 31.650 151.675 32.115 152.065 ;
        RECT 32.285 151.935 32.680 152.105 ;
        RECT 29.790 151.105 29.960 151.285 ;
        RECT 26.590 150.395 27.660 150.565 ;
        RECT 27.830 150.185 28.020 150.625 ;
        RECT 28.190 150.355 29.140 150.635 ;
        RECT 29.450 150.545 29.710 150.935 ;
        RECT 30.130 150.865 30.920 151.115 ;
        RECT 29.360 150.375 29.710 150.545 ;
        RECT 29.920 150.185 30.250 150.645 ;
        RECT 31.125 150.575 31.295 151.285 ;
        RECT 31.650 151.085 31.820 151.675 ;
        RECT 31.465 150.865 31.820 151.085 ;
        RECT 31.990 150.865 32.340 151.485 ;
        RECT 32.510 150.575 32.680 151.935 ;
        RECT 33.045 151.765 33.370 152.550 ;
        RECT 32.850 150.715 33.310 151.765 ;
        RECT 31.125 150.405 31.980 150.575 ;
        RECT 32.185 150.405 32.680 150.575 ;
        RECT 32.850 150.185 33.180 150.545 ;
        RECT 33.540 150.445 33.710 152.565 ;
        RECT 33.880 152.235 34.210 152.735 ;
        RECT 34.380 152.065 34.635 152.565 ;
        RECT 33.885 151.895 34.635 152.065 ;
        RECT 33.885 150.905 34.115 151.895 ;
        RECT 34.285 151.075 34.635 151.725 ;
        RECT 34.810 151.570 35.100 152.735 ;
        RECT 35.935 151.765 36.265 152.565 ;
        RECT 36.435 151.935 36.765 152.735 ;
        RECT 37.065 151.765 37.395 152.565 ;
        RECT 38.040 151.935 38.290 152.735 ;
        RECT 35.935 151.595 38.370 151.765 ;
        RECT 38.560 151.595 38.730 152.735 ;
        RECT 38.900 151.595 39.240 152.565 ;
        RECT 39.785 152.055 40.040 152.425 ;
        RECT 39.700 151.885 40.040 152.055 ;
        RECT 40.220 151.935 40.505 152.735 ;
        RECT 40.685 152.015 41.015 152.525 ;
        RECT 35.730 151.175 36.080 151.425 ;
        RECT 36.265 150.965 36.435 151.595 ;
        RECT 36.605 151.175 36.935 151.375 ;
        RECT 37.105 151.175 37.435 151.375 ;
        RECT 37.605 151.175 38.025 151.375 ;
        RECT 38.200 151.345 38.370 151.595 ;
        RECT 38.200 151.175 38.895 151.345 ;
        RECT 33.885 150.735 34.635 150.905 ;
        RECT 33.880 150.185 34.210 150.565 ;
        RECT 34.380 150.445 34.635 150.735 ;
        RECT 34.810 150.185 35.100 150.910 ;
        RECT 35.935 150.355 36.435 150.965 ;
        RECT 37.065 150.835 38.290 151.005 ;
        RECT 39.065 150.985 39.240 151.595 ;
        RECT 37.065 150.355 37.395 150.835 ;
        RECT 37.565 150.185 37.790 150.645 ;
        RECT 37.960 150.355 38.290 150.835 ;
        RECT 38.480 150.185 38.730 150.985 ;
        RECT 38.900 150.355 39.240 150.985 ;
        RECT 39.785 151.755 40.040 151.885 ;
        RECT 39.785 150.895 39.965 151.755 ;
        RECT 40.685 151.425 40.935 152.015 ;
        RECT 41.285 151.865 41.455 152.475 ;
        RECT 41.625 152.045 41.955 152.735 ;
        RECT 42.185 152.185 42.425 152.475 ;
        RECT 42.625 152.355 43.045 152.735 ;
        RECT 43.225 152.265 43.855 152.515 ;
        RECT 44.325 152.355 44.655 152.735 ;
        RECT 43.225 152.185 43.395 152.265 ;
        RECT 44.825 152.185 44.995 152.475 ;
        RECT 45.175 152.355 45.555 152.735 ;
        RECT 45.795 152.350 46.625 152.520 ;
        RECT 42.185 152.015 43.395 152.185 ;
        RECT 40.135 151.095 40.935 151.425 ;
        RECT 39.785 150.365 40.040 150.895 ;
        RECT 40.220 150.185 40.505 150.645 ;
        RECT 40.685 150.445 40.935 151.095 ;
        RECT 41.135 151.845 41.455 151.865 ;
        RECT 41.135 151.675 43.055 151.845 ;
        RECT 41.135 150.780 41.325 151.675 ;
        RECT 43.225 151.505 43.395 152.015 ;
        RECT 43.565 151.755 44.085 152.065 ;
        RECT 41.495 151.335 43.395 151.505 ;
        RECT 41.495 151.275 41.825 151.335 ;
        RECT 41.975 151.105 42.305 151.165 ;
        RECT 41.645 150.835 42.305 151.105 ;
        RECT 41.135 150.450 41.455 150.780 ;
        RECT 41.635 150.185 42.295 150.665 ;
        RECT 42.495 150.575 42.665 151.335 ;
        RECT 43.565 151.165 43.745 151.575 ;
        RECT 42.835 150.995 43.165 151.115 ;
        RECT 43.915 150.995 44.085 151.755 ;
        RECT 42.835 150.825 44.085 150.995 ;
        RECT 44.255 151.935 45.625 152.185 ;
        RECT 44.255 151.165 44.445 151.935 ;
        RECT 45.375 151.675 45.625 151.935 ;
        RECT 44.615 151.505 44.865 151.665 ;
        RECT 45.795 151.505 45.965 152.350 ;
        RECT 46.860 152.065 47.030 152.565 ;
        RECT 47.200 152.235 47.530 152.735 ;
        RECT 46.135 151.675 46.635 152.055 ;
        RECT 46.860 151.895 47.555 152.065 ;
        RECT 44.615 151.335 45.965 151.505 ;
        RECT 45.545 151.295 45.965 151.335 ;
        RECT 44.255 150.825 44.675 151.165 ;
        RECT 44.965 150.835 45.375 151.165 ;
        RECT 42.495 150.405 43.345 150.575 ;
        RECT 43.905 150.185 44.225 150.645 ;
        RECT 44.425 150.395 44.675 150.825 ;
        RECT 44.965 150.185 45.375 150.625 ;
        RECT 45.545 150.565 45.715 151.295 ;
        RECT 45.885 150.745 46.235 151.115 ;
        RECT 46.415 150.805 46.635 151.675 ;
        RECT 46.805 151.105 47.215 151.725 ;
        RECT 47.385 150.925 47.555 151.895 ;
        RECT 46.860 150.735 47.555 150.925 ;
        RECT 45.545 150.365 46.560 150.565 ;
        RECT 46.860 150.405 47.030 150.735 ;
        RECT 47.200 150.185 47.530 150.565 ;
        RECT 47.745 150.445 47.970 152.565 ;
        RECT 48.140 152.235 48.470 152.735 ;
        RECT 48.640 152.065 48.810 152.565 ;
        RECT 48.145 151.895 48.810 152.065 ;
        RECT 48.145 150.905 48.375 151.895 ;
        RECT 48.545 151.075 48.895 151.725 ;
        RECT 49.530 151.645 53.040 152.735 ;
        RECT 49.530 151.125 51.220 151.645 ;
        RECT 53.210 151.595 53.480 152.565 ;
        RECT 53.690 151.935 53.970 152.735 ;
        RECT 54.140 152.225 55.795 152.515 ;
        RECT 54.205 151.885 55.795 152.055 ;
        RECT 54.205 151.765 54.375 151.885 ;
        RECT 53.650 151.595 54.375 151.765 ;
        RECT 51.390 150.955 53.040 151.475 ;
        RECT 48.145 150.735 48.810 150.905 ;
        RECT 48.140 150.185 48.470 150.565 ;
        RECT 48.640 150.445 48.810 150.735 ;
        RECT 49.530 150.185 53.040 150.955 ;
        RECT 53.210 150.860 53.380 151.595 ;
        RECT 53.650 151.425 53.820 151.595 ;
        RECT 54.565 151.545 55.280 151.715 ;
        RECT 55.475 151.595 55.795 151.885 ;
        RECT 55.970 151.975 56.485 152.385 ;
        RECT 56.720 151.975 56.890 152.735 ;
        RECT 57.060 152.395 59.090 152.565 ;
        RECT 53.550 151.095 53.820 151.425 ;
        RECT 53.990 151.095 54.395 151.425 ;
        RECT 54.565 151.095 55.275 151.545 ;
        RECT 53.650 150.925 53.820 151.095 ;
        RECT 53.210 150.515 53.480 150.860 ;
        RECT 53.650 150.755 55.260 150.925 ;
        RECT 55.445 150.855 55.795 151.425 ;
        RECT 55.970 151.165 56.310 151.975 ;
        RECT 57.060 151.730 57.230 152.395 ;
        RECT 57.625 152.055 58.750 152.225 ;
        RECT 56.480 151.540 57.230 151.730 ;
        RECT 57.400 151.715 58.410 151.885 ;
        RECT 55.970 150.995 57.200 151.165 ;
        RECT 53.670 150.185 54.050 150.585 ;
        RECT 54.220 150.405 54.390 150.755 ;
        RECT 54.560 150.185 54.890 150.585 ;
        RECT 55.090 150.405 55.260 150.755 ;
        RECT 55.460 150.185 55.790 150.685 ;
        RECT 56.245 150.390 56.490 150.995 ;
        RECT 56.710 150.185 57.220 150.720 ;
        RECT 57.400 150.355 57.590 151.715 ;
        RECT 57.760 150.695 58.035 151.515 ;
        RECT 58.240 150.915 58.410 151.715 ;
        RECT 58.580 150.925 58.750 152.055 ;
        RECT 58.920 151.425 59.090 152.395 ;
        RECT 59.260 151.595 59.430 152.735 ;
        RECT 59.600 151.595 59.935 152.565 ;
        RECT 58.920 151.095 59.115 151.425 ;
        RECT 59.340 151.095 59.595 151.425 ;
        RECT 59.340 150.925 59.510 151.095 ;
        RECT 59.765 150.925 59.935 151.595 ;
        RECT 60.570 151.570 60.860 152.735 ;
        RECT 61.030 152.015 61.490 152.565 ;
        RECT 61.680 152.015 62.010 152.735 ;
        RECT 58.580 150.755 59.510 150.925 ;
        RECT 58.580 150.720 58.755 150.755 ;
        RECT 57.760 150.525 58.040 150.695 ;
        RECT 57.760 150.355 58.035 150.525 ;
        RECT 58.225 150.355 58.755 150.720 ;
        RECT 59.180 150.185 59.510 150.585 ;
        RECT 59.680 150.355 59.935 150.925 ;
        RECT 60.570 150.185 60.860 150.910 ;
        RECT 61.030 150.645 61.280 152.015 ;
        RECT 62.210 151.845 62.510 152.395 ;
        RECT 62.680 152.065 62.960 152.735 ;
        RECT 61.570 151.675 62.510 151.845 ;
        RECT 63.330 151.975 63.845 152.385 ;
        RECT 64.080 151.975 64.250 152.735 ;
        RECT 64.420 152.395 66.450 152.565 ;
        RECT 61.570 151.425 61.740 151.675 ;
        RECT 62.880 151.425 63.145 151.785 ;
        RECT 61.450 151.095 61.740 151.425 ;
        RECT 61.910 151.175 62.250 151.425 ;
        RECT 62.470 151.175 63.145 151.425 ;
        RECT 61.570 151.005 61.740 151.095 ;
        RECT 63.330 151.165 63.670 151.975 ;
        RECT 64.420 151.730 64.590 152.395 ;
        RECT 64.985 152.055 66.110 152.225 ;
        RECT 63.840 151.540 64.590 151.730 ;
        RECT 64.760 151.715 65.770 151.885 ;
        RECT 61.570 150.815 62.960 151.005 ;
        RECT 63.330 150.995 64.560 151.165 ;
        RECT 61.030 150.355 61.590 150.645 ;
        RECT 61.760 150.185 62.010 150.645 ;
        RECT 62.630 150.455 62.960 150.815 ;
        RECT 63.605 150.390 63.850 150.995 ;
        RECT 64.070 150.185 64.580 150.720 ;
        RECT 64.760 150.355 64.950 151.715 ;
        RECT 65.120 151.375 65.395 151.515 ;
        RECT 65.120 151.205 65.400 151.375 ;
        RECT 65.120 150.355 65.395 151.205 ;
        RECT 65.600 150.915 65.770 151.715 ;
        RECT 65.940 150.925 66.110 152.055 ;
        RECT 66.280 151.425 66.450 152.395 ;
        RECT 66.620 151.595 66.790 152.735 ;
        RECT 66.960 151.595 67.295 152.565 ;
        RECT 66.280 151.095 66.475 151.425 ;
        RECT 66.700 151.095 66.955 151.425 ;
        RECT 66.700 150.925 66.870 151.095 ;
        RECT 67.125 150.925 67.295 151.595 ;
        RECT 67.470 151.645 69.140 152.735 ;
        RECT 69.685 152.055 69.940 152.425 ;
        RECT 69.600 151.885 69.940 152.055 ;
        RECT 70.120 151.935 70.405 152.735 ;
        RECT 70.585 152.015 70.915 152.525 ;
        RECT 69.685 151.755 69.940 151.885 ;
        RECT 67.470 151.125 68.220 151.645 ;
        RECT 68.390 150.955 69.140 151.475 ;
        RECT 65.940 150.755 66.870 150.925 ;
        RECT 65.940 150.720 66.115 150.755 ;
        RECT 65.585 150.355 66.115 150.720 ;
        RECT 66.540 150.185 66.870 150.585 ;
        RECT 67.040 150.355 67.295 150.925 ;
        RECT 67.470 150.185 69.140 150.955 ;
        RECT 69.685 150.895 69.865 151.755 ;
        RECT 70.585 151.425 70.835 152.015 ;
        RECT 71.185 151.865 71.355 152.475 ;
        RECT 71.525 152.045 71.855 152.735 ;
        RECT 72.085 152.185 72.325 152.475 ;
        RECT 72.525 152.355 72.945 152.735 ;
        RECT 73.125 152.265 73.755 152.515 ;
        RECT 74.225 152.355 74.555 152.735 ;
        RECT 73.125 152.185 73.295 152.265 ;
        RECT 74.725 152.185 74.895 152.475 ;
        RECT 75.075 152.355 75.455 152.735 ;
        RECT 75.695 152.350 76.525 152.520 ;
        RECT 72.085 152.015 73.295 152.185 ;
        RECT 70.035 151.095 70.835 151.425 ;
        RECT 69.685 150.365 69.940 150.895 ;
        RECT 70.120 150.185 70.405 150.645 ;
        RECT 70.585 150.445 70.835 151.095 ;
        RECT 71.035 151.845 71.355 151.865 ;
        RECT 71.035 151.675 72.955 151.845 ;
        RECT 71.035 150.780 71.225 151.675 ;
        RECT 73.125 151.505 73.295 152.015 ;
        RECT 73.465 151.755 73.985 152.065 ;
        RECT 71.395 151.335 73.295 151.505 ;
        RECT 71.395 151.275 71.725 151.335 ;
        RECT 71.875 151.105 72.205 151.165 ;
        RECT 71.545 150.835 72.205 151.105 ;
        RECT 71.035 150.450 71.355 150.780 ;
        RECT 71.535 150.185 72.195 150.665 ;
        RECT 72.395 150.575 72.565 151.335 ;
        RECT 73.465 151.165 73.645 151.575 ;
        RECT 72.735 150.995 73.065 151.115 ;
        RECT 73.815 150.995 73.985 151.755 ;
        RECT 72.735 150.825 73.985 150.995 ;
        RECT 74.155 151.935 75.525 152.185 ;
        RECT 74.155 151.165 74.345 151.935 ;
        RECT 75.275 151.675 75.525 151.935 ;
        RECT 74.515 151.505 74.765 151.665 ;
        RECT 75.695 151.505 75.865 152.350 ;
        RECT 76.760 152.065 76.930 152.565 ;
        RECT 77.100 152.235 77.430 152.735 ;
        RECT 76.035 151.675 76.535 152.055 ;
        RECT 76.760 151.895 77.455 152.065 ;
        RECT 74.515 151.335 75.865 151.505 ;
        RECT 75.445 151.295 75.865 151.335 ;
        RECT 74.155 150.825 74.575 151.165 ;
        RECT 74.865 150.835 75.275 151.165 ;
        RECT 72.395 150.405 73.245 150.575 ;
        RECT 73.805 150.185 74.125 150.645 ;
        RECT 74.325 150.395 74.575 150.825 ;
        RECT 74.865 150.185 75.275 150.625 ;
        RECT 75.445 150.565 75.615 151.295 ;
        RECT 75.785 150.745 76.135 151.115 ;
        RECT 76.315 150.805 76.535 151.675 ;
        RECT 76.705 151.105 77.115 151.725 ;
        RECT 77.285 150.925 77.455 151.895 ;
        RECT 76.760 150.735 77.455 150.925 ;
        RECT 75.445 150.365 76.460 150.565 ;
        RECT 76.760 150.405 76.930 150.735 ;
        RECT 77.100 150.185 77.430 150.565 ;
        RECT 77.645 150.445 77.870 152.565 ;
        RECT 78.040 152.235 78.370 152.735 ;
        RECT 78.540 152.065 78.710 152.565 ;
        RECT 78.045 151.895 78.710 152.065 ;
        RECT 78.970 151.975 79.485 152.385 ;
        RECT 79.720 151.975 79.890 152.735 ;
        RECT 80.060 152.395 82.090 152.565 ;
        RECT 78.045 150.905 78.275 151.895 ;
        RECT 78.445 151.075 78.795 151.725 ;
        RECT 78.970 151.165 79.310 151.975 ;
        RECT 80.060 151.730 80.230 152.395 ;
        RECT 80.625 152.055 81.750 152.225 ;
        RECT 79.480 151.540 80.230 151.730 ;
        RECT 80.400 151.715 81.410 151.885 ;
        RECT 78.970 150.995 80.200 151.165 ;
        RECT 78.045 150.735 78.710 150.905 ;
        RECT 78.040 150.185 78.370 150.565 ;
        RECT 78.540 150.445 78.710 150.735 ;
        RECT 79.245 150.390 79.490 150.995 ;
        RECT 79.710 150.185 80.220 150.720 ;
        RECT 80.400 150.355 80.590 151.715 ;
        RECT 80.760 151.375 81.035 151.515 ;
        RECT 80.760 151.205 81.040 151.375 ;
        RECT 80.760 150.355 81.035 151.205 ;
        RECT 81.240 150.915 81.410 151.715 ;
        RECT 81.580 150.925 81.750 152.055 ;
        RECT 81.920 151.425 82.090 152.395 ;
        RECT 82.260 151.595 82.430 152.735 ;
        RECT 82.600 151.595 82.935 152.565 ;
        RECT 83.625 151.865 83.910 152.735 ;
        RECT 84.080 152.105 84.340 152.565 ;
        RECT 84.515 152.275 84.770 152.735 ;
        RECT 84.940 152.105 85.200 152.565 ;
        RECT 84.080 151.935 85.200 152.105 ;
        RECT 85.370 151.935 85.680 152.735 ;
        RECT 84.080 151.685 84.340 151.935 ;
        RECT 85.850 151.765 86.160 152.565 ;
        RECT 81.920 151.095 82.115 151.425 ;
        RECT 82.340 151.095 82.595 151.425 ;
        RECT 82.340 150.925 82.510 151.095 ;
        RECT 82.765 150.925 82.935 151.595 ;
        RECT 81.580 150.755 82.510 150.925 ;
        RECT 81.580 150.720 81.755 150.755 ;
        RECT 81.225 150.355 81.755 150.720 ;
        RECT 82.180 150.185 82.510 150.585 ;
        RECT 82.680 150.355 82.935 150.925 ;
        RECT 83.585 151.515 84.340 151.685 ;
        RECT 85.130 151.595 86.160 151.765 ;
        RECT 83.585 151.005 83.990 151.515 ;
        RECT 85.130 151.345 85.300 151.595 ;
        RECT 84.160 151.175 85.300 151.345 ;
        RECT 83.585 150.835 85.235 151.005 ;
        RECT 85.470 150.855 85.820 151.425 ;
        RECT 83.630 150.185 83.910 150.665 ;
        RECT 84.080 150.445 84.340 150.835 ;
        RECT 84.515 150.185 84.770 150.665 ;
        RECT 84.940 150.445 85.235 150.835 ;
        RECT 85.990 150.685 86.160 151.595 ;
        RECT 86.330 151.570 86.620 152.735 ;
        RECT 86.790 151.645 88.000 152.735 ;
        RECT 88.175 152.225 89.830 152.515 ;
        RECT 88.175 151.885 89.765 152.055 ;
        RECT 90.000 151.935 90.280 152.735 ;
        RECT 86.790 151.105 87.310 151.645 ;
        RECT 88.175 151.595 88.495 151.885 ;
        RECT 89.595 151.765 89.765 151.885 ;
        RECT 87.480 150.935 88.000 151.475 ;
        RECT 85.415 150.185 85.690 150.665 ;
        RECT 85.860 150.355 86.160 150.685 ;
        RECT 86.330 150.185 86.620 150.910 ;
        RECT 86.790 150.185 88.000 150.935 ;
        RECT 88.175 150.855 88.525 151.425 ;
        RECT 88.695 151.095 89.405 151.715 ;
        RECT 89.595 151.595 90.320 151.765 ;
        RECT 90.490 151.595 90.760 152.565 ;
        RECT 90.150 151.425 90.320 151.595 ;
        RECT 89.575 151.095 89.980 151.425 ;
        RECT 90.150 151.095 90.420 151.425 ;
        RECT 90.150 150.925 90.320 151.095 ;
        RECT 88.710 150.755 90.320 150.925 ;
        RECT 90.590 150.860 90.760 151.595 ;
        RECT 88.180 150.185 88.510 150.685 ;
        RECT 88.710 150.405 88.880 150.755 ;
        RECT 89.080 150.185 89.410 150.585 ;
        RECT 89.580 150.405 89.750 150.755 ;
        RECT 89.920 150.185 90.300 150.585 ;
        RECT 90.490 150.515 90.760 150.860 ;
        RECT 91.850 151.765 92.160 152.565 ;
        RECT 92.330 151.935 92.640 152.735 ;
        RECT 92.810 152.105 93.070 152.565 ;
        RECT 93.240 152.275 93.495 152.735 ;
        RECT 93.670 152.105 93.930 152.565 ;
        RECT 92.810 151.935 93.930 152.105 ;
        RECT 91.850 151.595 92.880 151.765 ;
        RECT 91.850 150.685 92.020 151.595 ;
        RECT 92.190 150.855 92.540 151.425 ;
        RECT 92.710 151.345 92.880 151.595 ;
        RECT 93.670 151.685 93.930 151.935 ;
        RECT 94.100 151.865 94.385 152.735 ;
        RECT 93.670 151.515 94.425 151.685 ;
        RECT 95.130 151.595 95.340 152.735 ;
        RECT 92.710 151.175 93.850 151.345 ;
        RECT 94.020 151.005 94.425 151.515 ;
        RECT 95.510 151.585 95.840 152.565 ;
        RECT 96.010 151.595 96.240 152.735 ;
        RECT 96.910 151.645 100.420 152.735 ;
        RECT 100.595 152.300 105.940 152.735 ;
        RECT 92.775 150.835 94.425 151.005 ;
        RECT 91.850 150.355 92.150 150.685 ;
        RECT 92.320 150.185 92.595 150.665 ;
        RECT 92.775 150.445 93.070 150.835 ;
        RECT 93.240 150.185 93.495 150.665 ;
        RECT 93.670 150.445 93.930 150.835 ;
        RECT 94.100 150.185 94.380 150.665 ;
        RECT 95.130 150.185 95.340 151.005 ;
        RECT 95.510 150.985 95.760 151.585 ;
        RECT 95.930 151.175 96.260 151.425 ;
        RECT 96.910 151.125 98.600 151.645 ;
        RECT 95.510 150.355 95.840 150.985 ;
        RECT 96.010 150.185 96.240 151.005 ;
        RECT 98.770 150.955 100.420 151.475 ;
        RECT 102.185 151.050 102.535 152.300 ;
        RECT 106.150 151.595 106.380 152.735 ;
        RECT 106.550 151.585 106.880 152.565 ;
        RECT 107.050 151.595 107.260 152.735 ;
        RECT 107.490 151.645 111.000 152.735 ;
        RECT 111.170 151.645 112.380 152.735 ;
        RECT 96.910 150.185 100.420 150.955 ;
        RECT 104.015 150.730 104.355 151.560 ;
        RECT 106.130 151.175 106.460 151.425 ;
        RECT 100.595 150.185 105.940 150.730 ;
        RECT 106.150 150.185 106.380 151.005 ;
        RECT 106.630 150.985 106.880 151.585 ;
        RECT 107.490 151.125 109.180 151.645 ;
        RECT 106.550 150.355 106.880 150.985 ;
        RECT 107.050 150.185 107.260 151.005 ;
        RECT 109.350 150.955 111.000 151.475 ;
        RECT 111.170 151.105 111.690 151.645 ;
        RECT 107.490 150.185 111.000 150.955 ;
        RECT 111.860 150.935 112.380 151.475 ;
        RECT 111.170 150.185 112.380 150.935 ;
        RECT 18.165 150.015 112.465 150.185 ;
        RECT 18.250 149.265 19.460 150.015 ;
        RECT 18.250 148.725 18.770 149.265 ;
        RECT 20.610 149.195 20.820 150.015 ;
        RECT 20.990 149.215 21.320 149.845 ;
        RECT 18.940 148.555 19.460 149.095 ;
        RECT 20.990 148.615 21.240 149.215 ;
        RECT 21.490 149.195 21.720 150.015 ;
        RECT 21.930 149.290 22.220 150.015 ;
        RECT 22.700 149.545 22.870 150.015 ;
        RECT 23.040 149.365 23.370 149.845 ;
        RECT 23.540 149.545 23.710 150.015 ;
        RECT 23.880 149.365 24.210 149.845 ;
        RECT 22.445 149.195 24.210 149.365 ;
        RECT 24.380 149.205 24.550 150.015 ;
        RECT 24.750 149.635 25.820 149.805 ;
        RECT 24.750 149.280 25.070 149.635 ;
        RECT 21.410 148.775 21.740 149.025 ;
        RECT 22.445 148.645 22.855 149.195 ;
        RECT 24.745 149.025 25.070 149.280 ;
        RECT 23.040 148.815 25.070 149.025 ;
        RECT 24.725 148.805 25.070 148.815 ;
        RECT 25.240 149.065 25.480 149.465 ;
        RECT 25.650 149.405 25.820 149.635 ;
        RECT 25.990 149.575 26.180 150.015 ;
        RECT 26.350 149.565 27.300 149.845 ;
        RECT 27.520 149.655 27.870 149.825 ;
        RECT 25.650 149.235 26.180 149.405 ;
        RECT 18.250 147.465 19.460 148.555 ;
        RECT 20.610 147.465 20.820 148.605 ;
        RECT 20.990 147.635 21.320 148.615 ;
        RECT 21.490 147.465 21.720 148.605 ;
        RECT 21.930 147.465 22.220 148.630 ;
        RECT 22.445 148.475 24.170 148.645 ;
        RECT 22.700 147.465 22.870 148.305 ;
        RECT 23.080 147.635 23.330 148.475 ;
        RECT 23.540 147.465 23.710 148.305 ;
        RECT 23.880 147.635 24.170 148.475 ;
        RECT 24.380 147.465 24.550 148.525 ;
        RECT 24.725 148.185 24.895 148.805 ;
        RECT 25.240 148.695 25.780 149.065 ;
        RECT 25.960 148.955 26.180 149.235 ;
        RECT 26.350 148.785 26.520 149.565 ;
        RECT 26.115 148.615 26.520 148.785 ;
        RECT 26.690 148.775 27.040 149.395 ;
        RECT 26.115 148.525 26.285 148.615 ;
        RECT 27.210 148.605 27.420 149.395 ;
        RECT 25.065 148.355 26.285 148.525 ;
        RECT 26.745 148.445 27.420 148.605 ;
        RECT 24.725 148.015 25.525 148.185 ;
        RECT 24.845 147.465 25.175 147.845 ;
        RECT 25.355 147.725 25.525 148.015 ;
        RECT 26.115 147.975 26.285 148.355 ;
        RECT 26.455 148.435 27.420 148.445 ;
        RECT 27.610 149.265 27.870 149.655 ;
        RECT 28.080 149.555 28.410 150.015 ;
        RECT 29.285 149.625 30.140 149.795 ;
        RECT 30.345 149.625 30.840 149.795 ;
        RECT 31.010 149.655 31.340 150.015 ;
        RECT 27.610 148.575 27.780 149.265 ;
        RECT 27.950 148.915 28.120 149.095 ;
        RECT 28.290 149.085 29.080 149.335 ;
        RECT 29.285 148.915 29.455 149.625 ;
        RECT 29.625 149.115 29.980 149.335 ;
        RECT 27.950 148.745 29.640 148.915 ;
        RECT 26.455 148.145 26.915 148.435 ;
        RECT 27.610 148.405 29.110 148.575 ;
        RECT 27.610 148.265 27.780 148.405 ;
        RECT 27.220 148.095 27.780 148.265 ;
        RECT 25.695 147.465 25.945 147.925 ;
        RECT 26.115 147.635 26.985 147.975 ;
        RECT 27.220 147.635 27.390 148.095 ;
        RECT 28.225 148.065 29.300 148.235 ;
        RECT 27.560 147.465 27.930 147.925 ;
        RECT 28.225 147.725 28.395 148.065 ;
        RECT 28.565 147.465 28.895 147.895 ;
        RECT 29.130 147.725 29.300 148.065 ;
        RECT 29.470 147.965 29.640 148.745 ;
        RECT 29.810 148.525 29.980 149.115 ;
        RECT 30.150 148.715 30.500 149.335 ;
        RECT 29.810 148.135 30.275 148.525 ;
        RECT 30.670 148.265 30.840 149.625 ;
        RECT 31.010 148.435 31.470 149.485 ;
        RECT 30.445 148.095 30.840 148.265 ;
        RECT 30.445 147.965 30.615 148.095 ;
        RECT 29.470 147.635 30.150 147.965 ;
        RECT 30.365 147.635 30.615 147.965 ;
        RECT 30.785 147.465 31.035 147.925 ;
        RECT 31.205 147.650 31.530 148.435 ;
        RECT 31.700 147.635 31.870 149.755 ;
        RECT 32.040 149.635 32.370 150.015 ;
        RECT 32.540 149.465 32.795 149.755 ;
        RECT 32.045 149.295 32.795 149.465 ;
        RECT 32.975 149.305 33.230 149.835 ;
        RECT 33.400 149.555 33.705 150.015 ;
        RECT 33.950 149.635 35.020 149.805 ;
        RECT 32.045 148.305 32.275 149.295 ;
        RECT 32.445 148.475 32.795 149.125 ;
        RECT 32.975 148.655 33.185 149.305 ;
        RECT 33.950 149.280 34.270 149.635 ;
        RECT 33.945 149.105 34.270 149.280 ;
        RECT 33.355 148.805 34.270 149.105 ;
        RECT 34.440 149.065 34.680 149.465 ;
        RECT 34.850 149.405 35.020 149.635 ;
        RECT 35.190 149.575 35.380 150.015 ;
        RECT 35.550 149.565 36.500 149.845 ;
        RECT 36.720 149.655 37.070 149.825 ;
        RECT 34.850 149.235 35.380 149.405 ;
        RECT 33.355 148.775 34.095 148.805 ;
        RECT 32.045 148.135 32.795 148.305 ;
        RECT 32.040 147.465 32.370 147.965 ;
        RECT 32.540 147.635 32.795 148.135 ;
        RECT 32.975 147.775 33.230 148.655 ;
        RECT 33.400 147.465 33.705 148.605 ;
        RECT 33.925 148.185 34.095 148.775 ;
        RECT 34.440 148.695 34.980 149.065 ;
        RECT 35.160 148.955 35.380 149.235 ;
        RECT 35.550 148.785 35.720 149.565 ;
        RECT 35.315 148.615 35.720 148.785 ;
        RECT 35.890 148.775 36.240 149.395 ;
        RECT 35.315 148.525 35.485 148.615 ;
        RECT 36.410 148.605 36.620 149.395 ;
        RECT 34.265 148.355 35.485 148.525 ;
        RECT 35.945 148.445 36.620 148.605 ;
        RECT 33.925 148.015 34.725 148.185 ;
        RECT 34.045 147.465 34.375 147.845 ;
        RECT 34.555 147.725 34.725 148.015 ;
        RECT 35.315 147.975 35.485 148.355 ;
        RECT 35.655 148.435 36.620 148.445 ;
        RECT 36.810 149.265 37.070 149.655 ;
        RECT 37.280 149.555 37.610 150.015 ;
        RECT 38.485 149.625 39.340 149.795 ;
        RECT 39.545 149.625 40.040 149.795 ;
        RECT 40.210 149.655 40.540 150.015 ;
        RECT 36.810 148.575 36.980 149.265 ;
        RECT 37.150 148.915 37.320 149.095 ;
        RECT 37.490 149.085 38.280 149.335 ;
        RECT 38.485 148.915 38.655 149.625 ;
        RECT 38.825 149.115 39.180 149.335 ;
        RECT 37.150 148.745 38.840 148.915 ;
        RECT 35.655 148.145 36.115 148.435 ;
        RECT 36.810 148.405 38.310 148.575 ;
        RECT 36.810 148.265 36.980 148.405 ;
        RECT 36.420 148.095 36.980 148.265 ;
        RECT 34.895 147.465 35.145 147.925 ;
        RECT 35.315 147.635 36.185 147.975 ;
        RECT 36.420 147.635 36.590 148.095 ;
        RECT 37.425 148.065 38.500 148.235 ;
        RECT 36.760 147.465 37.130 147.925 ;
        RECT 37.425 147.725 37.595 148.065 ;
        RECT 37.765 147.465 38.095 147.895 ;
        RECT 38.330 147.725 38.500 148.065 ;
        RECT 38.670 147.965 38.840 148.745 ;
        RECT 39.010 148.525 39.180 149.115 ;
        RECT 39.350 148.715 39.700 149.335 ;
        RECT 39.010 148.135 39.475 148.525 ;
        RECT 39.870 148.265 40.040 149.625 ;
        RECT 40.210 148.435 40.670 149.485 ;
        RECT 39.645 148.095 40.040 148.265 ;
        RECT 39.645 147.965 39.815 148.095 ;
        RECT 38.670 147.635 39.350 147.965 ;
        RECT 39.565 147.635 39.815 147.965 ;
        RECT 39.985 147.465 40.235 147.925 ;
        RECT 40.405 147.650 40.730 148.435 ;
        RECT 40.900 147.635 41.070 149.755 ;
        RECT 41.240 149.635 41.570 150.015 ;
        RECT 41.740 149.465 41.995 149.755 ;
        RECT 41.245 149.295 41.995 149.465 ;
        RECT 41.245 148.305 41.475 149.295 ;
        RECT 42.670 149.195 42.900 150.015 ;
        RECT 43.070 149.215 43.400 149.845 ;
        RECT 41.645 148.475 41.995 149.125 ;
        RECT 42.650 148.775 42.980 149.025 ;
        RECT 43.150 148.615 43.400 149.215 ;
        RECT 43.570 149.195 43.780 150.015 ;
        RECT 44.010 149.215 44.350 149.845 ;
        RECT 44.520 149.215 44.770 150.015 ;
        RECT 44.960 149.365 45.290 149.845 ;
        RECT 45.460 149.555 45.685 150.015 ;
        RECT 45.855 149.365 46.185 149.845 ;
        RECT 41.245 148.135 41.995 148.305 ;
        RECT 41.240 147.465 41.570 147.965 ;
        RECT 41.740 147.635 41.995 148.135 ;
        RECT 42.670 147.465 42.900 148.605 ;
        RECT 43.070 147.635 43.400 148.615 ;
        RECT 44.010 148.605 44.185 149.215 ;
        RECT 44.960 149.195 46.185 149.365 ;
        RECT 46.815 149.235 47.315 149.845 ;
        RECT 47.690 149.290 47.980 150.015 ;
        RECT 48.610 149.245 52.120 150.015 ;
        RECT 52.665 149.675 52.920 149.835 ;
        RECT 52.580 149.505 52.920 149.675 ;
        RECT 53.100 149.555 53.385 150.015 ;
        RECT 44.355 148.855 45.050 149.025 ;
        RECT 44.880 148.605 45.050 148.855 ;
        RECT 45.225 148.825 45.645 149.025 ;
        RECT 45.815 148.825 46.145 149.025 ;
        RECT 46.315 148.825 46.645 149.025 ;
        RECT 46.815 148.605 46.985 149.235 ;
        RECT 47.170 148.775 47.520 149.025 ;
        RECT 43.570 147.465 43.780 148.605 ;
        RECT 44.010 147.635 44.350 148.605 ;
        RECT 44.520 147.465 44.690 148.605 ;
        RECT 44.880 148.435 47.315 148.605 ;
        RECT 44.960 147.465 45.210 148.265 ;
        RECT 45.855 147.635 46.185 148.435 ;
        RECT 46.485 147.465 46.815 148.265 ;
        RECT 46.985 147.635 47.315 148.435 ;
        RECT 47.690 147.465 47.980 148.630 ;
        RECT 48.610 148.555 50.300 149.075 ;
        RECT 50.470 148.725 52.120 149.245 ;
        RECT 52.665 149.305 52.920 149.505 ;
        RECT 48.610 147.465 52.120 148.555 ;
        RECT 52.665 148.445 52.845 149.305 ;
        RECT 53.565 149.105 53.815 149.755 ;
        RECT 53.015 148.775 53.815 149.105 ;
        RECT 52.665 147.775 52.920 148.445 ;
        RECT 53.100 147.465 53.385 148.265 ;
        RECT 53.565 148.185 53.815 148.775 ;
        RECT 54.015 149.420 54.335 149.750 ;
        RECT 54.515 149.535 55.175 150.015 ;
        RECT 55.375 149.625 56.225 149.795 ;
        RECT 54.015 148.525 54.205 149.420 ;
        RECT 54.525 149.095 55.185 149.365 ;
        RECT 54.855 149.035 55.185 149.095 ;
        RECT 54.375 148.865 54.705 148.925 ;
        RECT 55.375 148.865 55.545 149.625 ;
        RECT 56.785 149.555 57.105 150.015 ;
        RECT 57.305 149.375 57.555 149.805 ;
        RECT 57.845 149.575 58.255 150.015 ;
        RECT 58.425 149.635 59.440 149.835 ;
        RECT 55.715 149.205 56.965 149.375 ;
        RECT 55.715 149.085 56.045 149.205 ;
        RECT 54.375 148.695 56.275 148.865 ;
        RECT 54.015 148.355 55.935 148.525 ;
        RECT 54.015 148.335 54.335 148.355 ;
        RECT 53.565 147.675 53.895 148.185 ;
        RECT 54.165 147.725 54.335 148.335 ;
        RECT 56.105 148.185 56.275 148.695 ;
        RECT 56.445 148.625 56.625 149.035 ;
        RECT 56.795 148.445 56.965 149.205 ;
        RECT 54.505 147.465 54.835 148.155 ;
        RECT 55.065 148.015 56.275 148.185 ;
        RECT 56.445 148.135 56.965 148.445 ;
        RECT 57.135 149.035 57.555 149.375 ;
        RECT 57.845 149.035 58.255 149.365 ;
        RECT 57.135 148.265 57.325 149.035 ;
        RECT 58.425 148.905 58.595 149.635 ;
        RECT 59.740 149.465 59.910 149.795 ;
        RECT 60.080 149.635 60.410 150.015 ;
        RECT 58.765 149.085 59.115 149.455 ;
        RECT 58.425 148.865 58.845 148.905 ;
        RECT 57.495 148.695 58.845 148.865 ;
        RECT 57.495 148.535 57.745 148.695 ;
        RECT 58.255 148.265 58.505 148.525 ;
        RECT 57.135 148.015 58.505 148.265 ;
        RECT 55.065 147.725 55.305 148.015 ;
        RECT 56.105 147.935 56.275 148.015 ;
        RECT 55.505 147.465 55.925 147.845 ;
        RECT 56.105 147.685 56.735 147.935 ;
        RECT 57.205 147.465 57.535 147.845 ;
        RECT 57.705 147.725 57.875 148.015 ;
        RECT 58.675 147.850 58.845 148.695 ;
        RECT 59.295 148.525 59.515 149.395 ;
        RECT 59.740 149.275 60.435 149.465 ;
        RECT 59.015 148.145 59.515 148.525 ;
        RECT 59.685 148.475 60.095 149.095 ;
        RECT 60.265 148.305 60.435 149.275 ;
        RECT 59.740 148.135 60.435 148.305 ;
        RECT 58.055 147.465 58.435 147.845 ;
        RECT 58.675 147.680 59.505 147.850 ;
        RECT 59.740 147.635 59.910 148.135 ;
        RECT 60.080 147.465 60.410 147.965 ;
        RECT 60.625 147.635 60.850 149.755 ;
        RECT 61.020 149.635 61.350 150.015 ;
        RECT 61.520 149.465 61.690 149.755 ;
        RECT 61.025 149.295 61.690 149.465 ;
        RECT 61.025 148.305 61.255 149.295 ;
        RECT 61.950 149.245 63.620 150.015 ;
        RECT 61.425 148.475 61.775 149.125 ;
        RECT 61.950 148.555 62.700 149.075 ;
        RECT 62.870 148.725 63.620 149.245 ;
        RECT 63.830 149.195 64.060 150.015 ;
        RECT 64.230 149.215 64.560 149.845 ;
        RECT 63.810 148.775 64.140 149.025 ;
        RECT 64.310 148.615 64.560 149.215 ;
        RECT 64.730 149.195 64.940 150.015 ;
        RECT 65.630 149.245 69.140 150.015 ;
        RECT 61.025 148.135 61.690 148.305 ;
        RECT 61.020 147.465 61.350 147.965 ;
        RECT 61.520 147.635 61.690 148.135 ;
        RECT 61.950 147.465 63.620 148.555 ;
        RECT 63.830 147.465 64.060 148.605 ;
        RECT 64.230 147.635 64.560 148.615 ;
        RECT 64.730 147.465 64.940 148.605 ;
        RECT 65.630 148.555 67.320 149.075 ;
        RECT 67.490 148.725 69.140 149.245 ;
        RECT 69.585 149.205 69.830 149.810 ;
        RECT 70.050 149.480 70.560 150.015 ;
        RECT 69.310 149.035 70.540 149.205 ;
        RECT 65.630 147.465 69.140 148.555 ;
        RECT 69.310 148.225 69.650 149.035 ;
        RECT 69.820 148.470 70.570 148.660 ;
        RECT 69.310 147.815 69.825 148.225 ;
        RECT 70.060 147.465 70.230 148.225 ;
        RECT 70.400 147.805 70.570 148.470 ;
        RECT 70.740 148.485 70.930 149.845 ;
        RECT 71.100 149.675 71.375 149.845 ;
        RECT 71.100 149.505 71.380 149.675 ;
        RECT 71.100 148.685 71.375 149.505 ;
        RECT 71.565 149.480 72.095 149.845 ;
        RECT 72.520 149.615 72.850 150.015 ;
        RECT 71.920 149.445 72.095 149.480 ;
        RECT 71.580 148.485 71.750 149.285 ;
        RECT 70.740 148.315 71.750 148.485 ;
        RECT 71.920 149.275 72.850 149.445 ;
        RECT 73.020 149.275 73.275 149.845 ;
        RECT 73.450 149.290 73.740 150.015 ;
        RECT 71.920 148.145 72.090 149.275 ;
        RECT 72.680 149.105 72.850 149.275 ;
        RECT 70.965 147.975 72.090 148.145 ;
        RECT 72.260 148.775 72.455 149.105 ;
        RECT 72.680 148.775 72.935 149.105 ;
        RECT 72.260 147.805 72.430 148.775 ;
        RECT 73.105 148.605 73.275 149.275 ;
        RECT 73.970 149.195 74.180 150.015 ;
        RECT 74.350 149.215 74.680 149.845 ;
        RECT 70.400 147.635 72.430 147.805 ;
        RECT 72.600 147.465 72.770 148.605 ;
        RECT 72.940 147.635 73.275 148.605 ;
        RECT 73.450 147.465 73.740 148.630 ;
        RECT 74.350 148.615 74.600 149.215 ;
        RECT 74.850 149.195 75.080 150.015 ;
        RECT 75.750 149.245 78.340 150.015 ;
        RECT 74.770 148.775 75.100 149.025 ;
        RECT 73.970 147.465 74.180 148.605 ;
        RECT 74.350 147.635 74.680 148.615 ;
        RECT 74.850 147.465 75.080 148.605 ;
        RECT 75.750 148.555 76.960 149.075 ;
        RECT 77.130 148.725 78.340 149.245 ;
        RECT 78.570 149.195 78.780 150.015 ;
        RECT 78.950 149.215 79.280 149.845 ;
        RECT 78.950 148.615 79.200 149.215 ;
        RECT 79.450 149.195 79.680 150.015 ;
        RECT 80.350 149.245 82.020 150.015 ;
        RECT 79.370 148.775 79.700 149.025 ;
        RECT 75.750 147.465 78.340 148.555 ;
        RECT 78.570 147.465 78.780 148.605 ;
        RECT 78.950 147.635 79.280 148.615 ;
        RECT 79.450 147.465 79.680 148.605 ;
        RECT 80.350 148.555 81.100 149.075 ;
        RECT 81.270 148.725 82.020 149.245 ;
        RECT 82.565 149.305 82.820 149.835 ;
        RECT 83.000 149.555 83.285 150.015 ;
        RECT 82.565 148.655 82.745 149.305 ;
        RECT 83.465 149.105 83.715 149.755 ;
        RECT 82.915 148.775 83.715 149.105 ;
        RECT 80.350 147.465 82.020 148.555 ;
        RECT 82.480 148.485 82.745 148.655 ;
        RECT 82.565 148.445 82.745 148.485 ;
        RECT 82.565 147.775 82.820 148.445 ;
        RECT 83.000 147.465 83.285 148.265 ;
        RECT 83.465 148.185 83.715 148.775 ;
        RECT 83.915 149.420 84.235 149.750 ;
        RECT 84.415 149.535 85.075 150.015 ;
        RECT 85.275 149.625 86.125 149.795 ;
        RECT 83.915 148.525 84.105 149.420 ;
        RECT 84.425 149.095 85.085 149.365 ;
        RECT 84.755 149.035 85.085 149.095 ;
        RECT 84.275 148.865 84.605 148.925 ;
        RECT 85.275 148.865 85.445 149.625 ;
        RECT 86.685 149.555 87.005 150.015 ;
        RECT 87.205 149.375 87.455 149.805 ;
        RECT 87.745 149.575 88.155 150.015 ;
        RECT 88.325 149.635 89.340 149.835 ;
        RECT 85.615 149.205 86.865 149.375 ;
        RECT 85.615 149.085 85.945 149.205 ;
        RECT 84.275 148.695 86.175 148.865 ;
        RECT 83.915 148.355 85.835 148.525 ;
        RECT 83.915 148.335 84.235 148.355 ;
        RECT 83.465 147.675 83.795 148.185 ;
        RECT 84.065 147.725 84.235 148.335 ;
        RECT 86.005 148.185 86.175 148.695 ;
        RECT 86.345 148.625 86.525 149.035 ;
        RECT 86.695 148.445 86.865 149.205 ;
        RECT 84.405 147.465 84.735 148.155 ;
        RECT 84.965 148.015 86.175 148.185 ;
        RECT 86.345 148.135 86.865 148.445 ;
        RECT 87.035 149.035 87.455 149.375 ;
        RECT 87.745 149.035 88.155 149.365 ;
        RECT 87.035 148.265 87.225 149.035 ;
        RECT 88.325 148.905 88.495 149.635 ;
        RECT 89.640 149.465 89.810 149.795 ;
        RECT 89.980 149.635 90.310 150.015 ;
        RECT 88.665 149.085 89.015 149.455 ;
        RECT 88.325 148.865 88.745 148.905 ;
        RECT 87.395 148.695 88.745 148.865 ;
        RECT 87.395 148.535 87.645 148.695 ;
        RECT 88.155 148.265 88.405 148.525 ;
        RECT 87.035 148.015 88.405 148.265 ;
        RECT 84.965 147.725 85.205 148.015 ;
        RECT 86.005 147.935 86.175 148.015 ;
        RECT 85.405 147.465 85.825 147.845 ;
        RECT 86.005 147.685 86.635 147.935 ;
        RECT 87.105 147.465 87.435 147.845 ;
        RECT 87.605 147.725 87.775 148.015 ;
        RECT 88.575 147.850 88.745 148.695 ;
        RECT 89.195 148.525 89.415 149.395 ;
        RECT 89.640 149.275 90.335 149.465 ;
        RECT 88.915 148.145 89.415 148.525 ;
        RECT 89.585 148.475 89.995 149.095 ;
        RECT 90.165 148.305 90.335 149.275 ;
        RECT 89.640 148.135 90.335 148.305 ;
        RECT 87.955 147.465 88.335 147.845 ;
        RECT 88.575 147.680 89.405 147.850 ;
        RECT 89.640 147.635 89.810 148.135 ;
        RECT 89.980 147.465 90.310 147.965 ;
        RECT 90.525 147.635 90.750 149.755 ;
        RECT 90.920 149.635 91.250 150.015 ;
        RECT 91.420 149.465 91.590 149.755 ;
        RECT 90.925 149.295 91.590 149.465 ;
        RECT 90.925 148.305 91.155 149.295 ;
        RECT 91.850 149.245 93.520 150.015 ;
        RECT 93.695 149.470 99.040 150.015 ;
        RECT 91.325 148.475 91.675 149.125 ;
        RECT 91.850 148.555 92.600 149.075 ;
        RECT 92.770 148.725 93.520 149.245 ;
        RECT 90.925 148.135 91.590 148.305 ;
        RECT 90.920 147.465 91.250 147.965 ;
        RECT 91.420 147.635 91.590 148.135 ;
        RECT 91.850 147.465 93.520 148.555 ;
        RECT 95.285 147.900 95.635 149.150 ;
        RECT 97.115 148.640 97.455 149.470 ;
        RECT 99.210 149.290 99.500 150.015 ;
        RECT 100.190 149.195 100.400 150.015 ;
        RECT 100.570 149.215 100.900 149.845 ;
        RECT 93.695 147.465 99.040 147.900 ;
        RECT 99.210 147.465 99.500 148.630 ;
        RECT 100.570 148.615 100.820 149.215 ;
        RECT 101.070 149.195 101.300 150.015 ;
        RECT 101.600 149.365 101.770 149.845 ;
        RECT 101.950 149.535 102.190 150.015 ;
        RECT 102.440 149.365 102.610 149.845 ;
        RECT 102.780 149.535 103.110 150.015 ;
        RECT 103.280 149.365 103.450 149.845 ;
        RECT 101.600 149.195 102.235 149.365 ;
        RECT 102.440 149.195 103.450 149.365 ;
        RECT 103.620 149.215 103.950 150.015 ;
        RECT 104.270 149.265 105.480 150.015 ;
        RECT 105.655 149.470 111.000 150.015 ;
        RECT 102.065 149.025 102.235 149.195 ;
        RECT 100.990 148.775 101.320 149.025 ;
        RECT 101.515 148.785 101.895 149.025 ;
        RECT 102.065 148.855 102.565 149.025 ;
        RECT 102.065 148.615 102.235 148.855 ;
        RECT 102.955 148.655 103.450 149.195 ;
        RECT 100.190 147.465 100.400 148.605 ;
        RECT 100.570 147.635 100.900 148.615 ;
        RECT 101.070 147.465 101.300 148.605 ;
        RECT 101.520 148.445 102.235 148.615 ;
        RECT 102.440 148.485 103.450 148.655 ;
        RECT 101.520 147.635 101.850 148.445 ;
        RECT 102.020 147.465 102.260 148.265 ;
        RECT 102.440 147.635 102.610 148.485 ;
        RECT 102.780 147.465 103.110 148.265 ;
        RECT 103.280 147.635 103.450 148.485 ;
        RECT 103.620 147.465 103.950 148.615 ;
        RECT 104.270 148.555 104.790 149.095 ;
        RECT 104.960 148.725 105.480 149.265 ;
        RECT 104.270 147.465 105.480 148.555 ;
        RECT 107.245 147.900 107.595 149.150 ;
        RECT 109.075 148.640 109.415 149.470 ;
        RECT 111.170 149.265 112.380 150.015 ;
        RECT 111.170 148.555 111.690 149.095 ;
        RECT 111.860 148.725 112.380 149.265 ;
        RECT 105.655 147.465 111.000 147.900 ;
        RECT 111.170 147.465 112.380 148.555 ;
        RECT 18.165 147.295 112.465 147.465 ;
        RECT 18.250 146.205 19.460 147.295 ;
        RECT 20.095 146.860 25.440 147.295 ;
        RECT 18.250 145.495 18.770 146.035 ;
        RECT 18.940 145.665 19.460 146.205 ;
        RECT 21.685 145.610 22.035 146.860 ;
        RECT 25.725 146.665 26.010 147.125 ;
        RECT 26.180 146.835 26.450 147.295 ;
        RECT 25.725 146.445 26.680 146.665 ;
        RECT 18.250 144.745 19.460 145.495 ;
        RECT 23.515 145.290 23.855 146.120 ;
        RECT 25.610 145.715 26.300 146.275 ;
        RECT 26.470 145.545 26.680 146.445 ;
        RECT 25.725 145.375 26.680 145.545 ;
        RECT 26.850 146.275 27.250 147.125 ;
        RECT 27.440 146.665 27.720 147.125 ;
        RECT 28.240 146.835 28.565 147.295 ;
        RECT 27.440 146.445 28.565 146.665 ;
        RECT 26.850 145.715 27.945 146.275 ;
        RECT 28.115 145.985 28.565 146.445 ;
        RECT 28.735 146.155 29.120 147.125 ;
        RECT 29.350 146.155 29.560 147.295 ;
        RECT 20.095 144.745 25.440 145.290 ;
        RECT 25.725 144.915 26.010 145.375 ;
        RECT 26.180 144.745 26.450 145.205 ;
        RECT 26.850 144.915 27.250 145.715 ;
        RECT 28.115 145.655 28.670 145.985 ;
        RECT 28.115 145.545 28.565 145.655 ;
        RECT 27.440 145.375 28.565 145.545 ;
        RECT 28.840 145.485 29.120 146.155 ;
        RECT 29.730 146.145 30.060 147.125 ;
        RECT 30.230 146.155 30.460 147.295 ;
        RECT 30.670 146.535 31.185 146.945 ;
        RECT 31.420 146.535 31.590 147.295 ;
        RECT 31.760 146.955 33.790 147.125 ;
        RECT 27.440 144.915 27.720 145.375 ;
        RECT 28.240 144.745 28.565 145.205 ;
        RECT 28.735 144.915 29.120 145.485 ;
        RECT 29.350 144.745 29.560 145.565 ;
        RECT 29.730 145.545 29.980 146.145 ;
        RECT 30.150 145.735 30.480 145.985 ;
        RECT 30.670 145.725 31.010 146.535 ;
        RECT 31.760 146.290 31.930 146.955 ;
        RECT 32.325 146.615 33.450 146.785 ;
        RECT 31.180 146.100 31.930 146.290 ;
        RECT 32.100 146.275 33.110 146.445 ;
        RECT 29.730 144.915 30.060 145.545 ;
        RECT 30.230 144.745 30.460 145.565 ;
        RECT 30.670 145.555 31.900 145.725 ;
        RECT 30.945 144.950 31.190 145.555 ;
        RECT 31.410 144.745 31.920 145.280 ;
        RECT 32.100 144.915 32.290 146.275 ;
        RECT 32.460 145.255 32.735 146.075 ;
        RECT 32.940 145.475 33.110 146.275 ;
        RECT 33.280 145.485 33.450 146.615 ;
        RECT 33.620 145.985 33.790 146.955 ;
        RECT 33.960 146.155 34.130 147.295 ;
        RECT 34.300 146.155 34.635 147.125 ;
        RECT 33.620 145.655 33.815 145.985 ;
        RECT 34.040 145.655 34.295 145.985 ;
        RECT 34.040 145.485 34.210 145.655 ;
        RECT 34.465 145.485 34.635 146.155 ;
        RECT 34.810 146.130 35.100 147.295 ;
        RECT 35.730 146.535 36.245 146.945 ;
        RECT 36.480 146.535 36.650 147.295 ;
        RECT 36.820 146.955 38.850 147.125 ;
        RECT 35.730 145.725 36.070 146.535 ;
        RECT 36.820 146.290 36.990 146.955 ;
        RECT 37.385 146.615 38.510 146.785 ;
        RECT 36.240 146.100 36.990 146.290 ;
        RECT 37.160 146.275 38.170 146.445 ;
        RECT 35.730 145.555 36.960 145.725 ;
        RECT 33.280 145.315 34.210 145.485 ;
        RECT 33.280 145.280 33.455 145.315 ;
        RECT 32.460 145.085 32.740 145.255 ;
        RECT 32.460 144.915 32.735 145.085 ;
        RECT 32.925 144.915 33.455 145.280 ;
        RECT 33.880 144.745 34.210 145.145 ;
        RECT 34.380 144.915 34.635 145.485 ;
        RECT 34.810 144.745 35.100 145.470 ;
        RECT 36.005 144.950 36.250 145.555 ;
        RECT 36.470 144.745 36.980 145.280 ;
        RECT 37.160 144.915 37.350 146.275 ;
        RECT 37.520 145.935 37.795 146.075 ;
        RECT 37.520 145.765 37.800 145.935 ;
        RECT 37.520 144.915 37.795 145.765 ;
        RECT 38.000 145.475 38.170 146.275 ;
        RECT 38.340 145.485 38.510 146.615 ;
        RECT 38.680 145.985 38.850 146.955 ;
        RECT 39.020 146.155 39.190 147.295 ;
        RECT 39.360 146.155 39.695 147.125 ;
        RECT 38.680 145.655 38.875 145.985 ;
        RECT 39.100 145.655 39.355 145.985 ;
        RECT 39.100 145.485 39.270 145.655 ;
        RECT 39.525 145.485 39.695 146.155 ;
        RECT 40.330 146.205 42.920 147.295 ;
        RECT 43.090 146.575 43.550 147.125 ;
        RECT 43.740 146.575 44.070 147.295 ;
        RECT 40.330 145.685 41.540 146.205 ;
        RECT 41.710 145.515 42.920 146.035 ;
        RECT 38.340 145.315 39.270 145.485 ;
        RECT 38.340 145.280 38.515 145.315 ;
        RECT 37.985 144.915 38.515 145.280 ;
        RECT 38.940 144.745 39.270 145.145 ;
        RECT 39.440 144.915 39.695 145.485 ;
        RECT 40.330 144.745 42.920 145.515 ;
        RECT 43.090 145.205 43.340 146.575 ;
        RECT 44.270 146.405 44.570 146.955 ;
        RECT 44.740 146.625 45.020 147.295 ;
        RECT 43.630 146.235 44.570 146.405 ;
        RECT 43.630 145.985 43.800 146.235 ;
        RECT 44.940 145.985 45.205 146.345 ;
        RECT 43.510 145.655 43.800 145.985 ;
        RECT 43.970 145.735 44.310 145.985 ;
        RECT 44.530 145.735 45.205 145.985 ;
        RECT 46.310 146.205 49.820 147.295 ;
        RECT 49.990 146.535 50.505 146.945 ;
        RECT 50.740 146.535 50.910 147.295 ;
        RECT 51.080 146.955 53.110 147.125 ;
        RECT 46.310 145.685 48.000 146.205 ;
        RECT 43.630 145.565 43.800 145.655 ;
        RECT 43.630 145.375 45.020 145.565 ;
        RECT 48.170 145.515 49.820 146.035 ;
        RECT 49.990 145.725 50.330 146.535 ;
        RECT 51.080 146.290 51.250 146.955 ;
        RECT 51.645 146.615 52.770 146.785 ;
        RECT 50.500 146.100 51.250 146.290 ;
        RECT 51.420 146.275 52.430 146.445 ;
        RECT 49.990 145.555 51.220 145.725 ;
        RECT 43.090 144.915 43.650 145.205 ;
        RECT 43.820 144.745 44.070 145.205 ;
        RECT 44.690 145.015 45.020 145.375 ;
        RECT 46.310 144.745 49.820 145.515 ;
        RECT 50.265 144.950 50.510 145.555 ;
        RECT 50.730 144.745 51.240 145.280 ;
        RECT 51.420 144.915 51.610 146.275 ;
        RECT 51.780 145.255 52.055 146.075 ;
        RECT 52.260 145.475 52.430 146.275 ;
        RECT 52.600 145.485 52.770 146.615 ;
        RECT 52.940 145.985 53.110 146.955 ;
        RECT 53.280 146.155 53.450 147.295 ;
        RECT 53.620 146.155 53.955 147.125 ;
        RECT 52.940 145.655 53.135 145.985 ;
        RECT 53.360 145.655 53.615 145.985 ;
        RECT 53.360 145.485 53.530 145.655 ;
        RECT 53.785 145.485 53.955 146.155 ;
        RECT 54.130 146.205 55.340 147.295 ;
        RECT 54.130 145.665 54.650 146.205 ;
        RECT 55.550 146.155 55.780 147.295 ;
        RECT 55.950 146.145 56.280 147.125 ;
        RECT 56.450 146.155 56.660 147.295 ;
        RECT 56.890 146.205 60.400 147.295 ;
        RECT 54.820 145.495 55.340 146.035 ;
        RECT 55.530 145.735 55.860 145.985 ;
        RECT 52.600 145.315 53.530 145.485 ;
        RECT 52.600 145.280 52.775 145.315 ;
        RECT 51.780 145.085 52.060 145.255 ;
        RECT 51.780 144.915 52.055 145.085 ;
        RECT 52.245 144.915 52.775 145.280 ;
        RECT 53.200 144.745 53.530 145.145 ;
        RECT 53.700 144.915 53.955 145.485 ;
        RECT 54.130 144.745 55.340 145.495 ;
        RECT 55.550 144.745 55.780 145.565 ;
        RECT 56.030 145.545 56.280 146.145 ;
        RECT 56.890 145.685 58.580 146.205 ;
        RECT 60.570 146.130 60.860 147.295 ;
        RECT 61.120 146.550 61.390 147.295 ;
        RECT 62.020 147.290 68.295 147.295 ;
        RECT 61.560 146.380 61.850 147.120 ;
        RECT 62.020 146.565 62.275 147.290 ;
        RECT 62.460 146.395 62.720 147.120 ;
        RECT 62.890 146.565 63.135 147.290 ;
        RECT 63.320 146.395 63.580 147.120 ;
        RECT 63.750 146.565 63.995 147.290 ;
        RECT 64.180 146.395 64.440 147.120 ;
        RECT 64.610 146.565 64.855 147.290 ;
        RECT 65.025 146.395 65.285 147.120 ;
        RECT 65.455 146.565 65.715 147.290 ;
        RECT 65.885 146.395 66.145 147.120 ;
        RECT 66.315 146.565 66.575 147.290 ;
        RECT 66.745 146.395 67.005 147.120 ;
        RECT 67.175 146.565 67.435 147.290 ;
        RECT 67.605 146.395 67.865 147.120 ;
        RECT 68.035 146.495 68.295 147.290 ;
        RECT 62.460 146.380 67.865 146.395 ;
        RECT 61.120 146.155 67.865 146.380 ;
        RECT 55.950 144.915 56.280 145.545 ;
        RECT 56.450 144.745 56.660 145.565 ;
        RECT 58.750 145.515 60.400 146.035 ;
        RECT 61.120 145.595 62.285 146.155 ;
        RECT 68.465 145.985 68.715 147.120 ;
        RECT 68.895 146.485 69.155 147.295 ;
        RECT 69.330 145.985 69.575 147.125 ;
        RECT 69.755 146.485 70.050 147.295 ;
        RECT 70.690 146.205 73.280 147.295 ;
        RECT 73.455 146.860 78.800 147.295 ;
        RECT 62.455 145.735 69.575 145.985 ;
        RECT 56.890 144.745 60.400 145.515 ;
        RECT 61.090 145.565 62.285 145.595 ;
        RECT 60.570 144.745 60.860 145.470 ;
        RECT 61.090 145.425 67.865 145.565 ;
        RECT 61.120 145.395 67.865 145.425 ;
        RECT 61.120 144.745 61.420 145.225 ;
        RECT 61.590 144.940 61.850 145.395 ;
        RECT 62.020 144.745 62.280 145.225 ;
        RECT 62.460 144.940 62.720 145.395 ;
        RECT 62.890 144.745 63.140 145.225 ;
        RECT 63.320 144.940 63.580 145.395 ;
        RECT 63.750 144.745 64.000 145.225 ;
        RECT 64.180 144.940 64.440 145.395 ;
        RECT 64.610 144.745 64.855 145.225 ;
        RECT 65.025 144.940 65.300 145.395 ;
        RECT 65.470 144.745 65.715 145.225 ;
        RECT 65.885 144.940 66.145 145.395 ;
        RECT 66.315 144.745 66.575 145.225 ;
        RECT 66.745 144.940 67.005 145.395 ;
        RECT 67.175 144.745 67.435 145.225 ;
        RECT 67.605 144.940 67.865 145.395 ;
        RECT 68.035 144.745 68.295 145.305 ;
        RECT 68.465 144.925 68.715 145.735 ;
        RECT 68.895 144.745 69.155 145.270 ;
        RECT 69.325 144.925 69.575 145.735 ;
        RECT 69.745 145.425 70.060 145.985 ;
        RECT 70.690 145.685 71.900 146.205 ;
        RECT 72.070 145.515 73.280 146.035 ;
        RECT 75.045 145.610 75.395 146.860 ;
        RECT 79.010 146.155 79.240 147.295 ;
        RECT 79.410 146.145 79.740 147.125 ;
        RECT 79.910 146.155 80.120 147.295 ;
        RECT 80.360 146.315 80.690 147.125 ;
        RECT 80.860 146.495 81.100 147.295 ;
        RECT 80.360 146.145 81.075 146.315 ;
        RECT 69.755 144.745 70.060 145.255 ;
        RECT 70.690 144.745 73.280 145.515 ;
        RECT 76.875 145.290 77.215 146.120 ;
        RECT 78.990 145.735 79.320 145.985 ;
        RECT 73.455 144.745 78.800 145.290 ;
        RECT 79.010 144.745 79.240 145.565 ;
        RECT 79.490 145.545 79.740 146.145 ;
        RECT 80.355 145.735 80.735 145.975 ;
        RECT 80.905 145.905 81.075 146.145 ;
        RECT 81.280 146.275 81.450 147.125 ;
        RECT 81.620 146.495 81.950 147.295 ;
        RECT 82.120 146.275 82.290 147.125 ;
        RECT 81.280 146.105 82.290 146.275 ;
        RECT 82.460 146.145 82.790 147.295 ;
        RECT 83.570 146.205 86.160 147.295 ;
        RECT 81.795 145.935 82.290 146.105 ;
        RECT 80.905 145.735 81.405 145.905 ;
        RECT 81.790 145.765 82.290 145.935 ;
        RECT 80.905 145.565 81.075 145.735 ;
        RECT 81.795 145.565 82.290 145.765 ;
        RECT 83.570 145.685 84.780 146.205 ;
        RECT 86.330 146.130 86.620 147.295 ;
        RECT 86.790 146.205 88.000 147.295 ;
        RECT 88.240 146.355 88.500 147.125 ;
        RECT 88.670 146.525 89.000 147.295 ;
        RECT 89.170 146.955 90.290 147.125 ;
        RECT 89.170 146.355 89.360 146.955 ;
        RECT 79.410 144.915 79.740 145.545 ;
        RECT 79.910 144.745 80.120 145.565 ;
        RECT 80.440 145.395 81.075 145.565 ;
        RECT 81.280 145.395 82.290 145.565 ;
        RECT 80.440 144.915 80.610 145.395 ;
        RECT 80.790 144.745 81.030 145.225 ;
        RECT 81.280 144.915 81.450 145.395 ;
        RECT 81.620 144.745 81.950 145.225 ;
        RECT 82.120 144.915 82.290 145.395 ;
        RECT 82.460 144.745 82.790 145.545 ;
        RECT 84.950 145.515 86.160 146.035 ;
        RECT 86.790 145.665 87.310 146.205 ;
        RECT 88.240 146.185 89.360 146.355 ;
        RECT 89.530 146.370 89.860 146.785 ;
        RECT 90.030 146.760 90.290 146.955 ;
        RECT 90.520 146.575 90.850 147.295 ;
        RECT 91.020 146.370 91.210 147.125 ;
        RECT 91.380 146.575 91.710 147.295 ;
        RECT 91.880 146.370 92.140 147.125 ;
        RECT 92.310 146.835 92.570 147.295 ;
        RECT 89.530 146.200 92.140 146.370 ;
        RECT 83.570 144.745 86.160 145.515 ;
        RECT 87.480 145.495 88.000 146.035 ;
        RECT 86.330 144.745 86.620 145.470 ;
        RECT 86.790 144.745 88.000 145.495 ;
        RECT 88.230 145.905 89.125 145.955 ;
        RECT 88.230 145.735 89.180 145.905 ;
        RECT 89.350 145.735 90.320 146.015 ;
        RECT 90.780 145.735 91.640 146.025 ;
        RECT 88.230 145.425 88.570 145.735 ;
        RECT 88.740 145.295 91.280 145.505 ;
        RECT 88.740 145.175 88.930 145.295 ;
        RECT 91.450 145.125 91.640 145.550 ;
        RECT 91.810 145.330 92.140 146.200 ;
        RECT 92.310 145.655 92.600 146.630 ;
        RECT 92.770 146.205 96.280 147.295 ;
        RECT 96.825 146.315 97.080 146.985 ;
        RECT 97.260 146.495 97.545 147.295 ;
        RECT 97.725 146.575 98.055 147.085 ;
        RECT 92.770 145.685 94.460 146.205 ;
        RECT 94.630 145.515 96.280 146.035 ;
        RECT 90.520 145.105 91.640 145.125 ;
        RECT 88.240 144.745 88.570 145.105 ;
        RECT 89.100 144.745 89.430 145.105 ;
        RECT 89.960 144.745 90.290 145.105 ;
        RECT 90.520 144.915 92.590 145.105 ;
        RECT 92.770 144.745 96.280 145.515 ;
        RECT 96.825 145.455 97.005 146.315 ;
        RECT 97.725 145.985 97.975 146.575 ;
        RECT 98.325 146.425 98.495 147.035 ;
        RECT 98.665 146.605 98.995 147.295 ;
        RECT 99.225 146.745 99.465 147.035 ;
        RECT 99.665 146.915 100.085 147.295 ;
        RECT 100.265 146.825 100.895 147.075 ;
        RECT 101.365 146.915 101.695 147.295 ;
        RECT 100.265 146.745 100.435 146.825 ;
        RECT 101.865 146.745 102.035 147.035 ;
        RECT 102.215 146.915 102.595 147.295 ;
        RECT 102.835 146.910 103.665 147.080 ;
        RECT 99.225 146.575 100.435 146.745 ;
        RECT 97.175 145.655 97.975 145.985 ;
        RECT 96.825 145.255 97.080 145.455 ;
        RECT 96.740 145.085 97.080 145.255 ;
        RECT 96.825 144.925 97.080 145.085 ;
        RECT 97.260 144.745 97.545 145.205 ;
        RECT 97.725 145.005 97.975 145.655 ;
        RECT 98.175 146.405 98.495 146.425 ;
        RECT 98.175 146.235 100.095 146.405 ;
        RECT 98.175 145.340 98.365 146.235 ;
        RECT 100.265 146.065 100.435 146.575 ;
        RECT 100.605 146.315 101.125 146.625 ;
        RECT 98.535 145.895 100.435 146.065 ;
        RECT 98.535 145.835 98.865 145.895 ;
        RECT 99.015 145.665 99.345 145.725 ;
        RECT 98.685 145.395 99.345 145.665 ;
        RECT 98.175 145.010 98.495 145.340 ;
        RECT 98.675 144.745 99.335 145.225 ;
        RECT 99.535 145.135 99.705 145.895 ;
        RECT 100.605 145.725 100.785 146.135 ;
        RECT 99.875 145.555 100.205 145.675 ;
        RECT 100.955 145.555 101.125 146.315 ;
        RECT 99.875 145.385 101.125 145.555 ;
        RECT 101.295 146.495 102.665 146.745 ;
        RECT 101.295 145.725 101.485 146.495 ;
        RECT 102.415 146.235 102.665 146.495 ;
        RECT 101.655 146.065 101.905 146.225 ;
        RECT 102.835 146.065 103.005 146.910 ;
        RECT 103.900 146.625 104.070 147.125 ;
        RECT 104.240 146.795 104.570 147.295 ;
        RECT 103.175 146.235 103.675 146.615 ;
        RECT 103.900 146.455 104.595 146.625 ;
        RECT 101.655 145.895 103.005 146.065 ;
        RECT 102.585 145.855 103.005 145.895 ;
        RECT 101.295 145.385 101.715 145.725 ;
        RECT 102.005 145.395 102.415 145.725 ;
        RECT 99.535 144.965 100.385 145.135 ;
        RECT 100.945 144.745 101.265 145.205 ;
        RECT 101.465 144.955 101.715 145.385 ;
        RECT 102.005 144.745 102.415 145.185 ;
        RECT 102.585 145.125 102.755 145.855 ;
        RECT 102.925 145.305 103.275 145.675 ;
        RECT 103.455 145.365 103.675 146.235 ;
        RECT 103.845 145.665 104.255 146.285 ;
        RECT 104.425 145.485 104.595 146.455 ;
        RECT 103.900 145.295 104.595 145.485 ;
        RECT 102.585 144.925 103.600 145.125 ;
        RECT 103.900 144.965 104.070 145.295 ;
        RECT 104.240 144.745 104.570 145.125 ;
        RECT 104.785 145.005 105.010 147.125 ;
        RECT 105.180 146.795 105.510 147.295 ;
        RECT 105.680 146.625 105.850 147.125 ;
        RECT 105.185 146.455 105.850 146.625 ;
        RECT 105.185 145.465 105.415 146.455 ;
        RECT 105.585 145.635 105.935 146.285 ;
        RECT 106.170 146.155 106.380 147.295 ;
        RECT 106.550 146.145 106.880 147.125 ;
        RECT 107.050 146.155 107.280 147.295 ;
        RECT 107.490 146.205 111.000 147.295 ;
        RECT 111.170 146.205 112.380 147.295 ;
        RECT 105.185 145.295 105.850 145.465 ;
        RECT 105.180 144.745 105.510 145.125 ;
        RECT 105.680 145.005 105.850 145.295 ;
        RECT 106.170 144.745 106.380 145.565 ;
        RECT 106.550 145.545 106.800 146.145 ;
        RECT 106.970 145.735 107.300 145.985 ;
        RECT 107.490 145.685 109.180 146.205 ;
        RECT 106.550 144.915 106.880 145.545 ;
        RECT 107.050 144.745 107.280 145.565 ;
        RECT 109.350 145.515 111.000 146.035 ;
        RECT 111.170 145.665 111.690 146.205 ;
        RECT 107.490 144.745 111.000 145.515 ;
        RECT 111.860 145.495 112.380 146.035 ;
        RECT 111.170 144.745 112.380 145.495 ;
        RECT 18.165 144.575 112.465 144.745 ;
        RECT 18.250 143.825 19.460 144.575 ;
        RECT 18.250 143.285 18.770 143.825 ;
        RECT 20.090 143.805 21.760 144.575 ;
        RECT 21.930 143.850 22.220 144.575 ;
        RECT 22.390 143.805 25.900 144.575 ;
        RECT 26.075 144.030 31.420 144.575 ;
        RECT 18.940 143.115 19.460 143.655 ;
        RECT 18.250 142.025 19.460 143.115 ;
        RECT 20.090 143.115 20.840 143.635 ;
        RECT 21.010 143.285 21.760 143.805 ;
        RECT 20.090 142.025 21.760 143.115 ;
        RECT 21.930 142.025 22.220 143.190 ;
        RECT 22.390 143.115 24.080 143.635 ;
        RECT 24.250 143.285 25.900 143.805 ;
        RECT 22.390 142.025 25.900 143.115 ;
        RECT 27.665 142.460 28.015 143.710 ;
        RECT 29.495 143.200 29.835 144.030 ;
        RECT 31.590 143.835 31.975 144.405 ;
        RECT 32.145 144.115 32.470 144.575 ;
        RECT 32.990 143.945 33.270 144.405 ;
        RECT 31.590 143.165 31.870 143.835 ;
        RECT 32.145 143.775 33.270 143.945 ;
        RECT 32.145 143.665 32.595 143.775 ;
        RECT 32.040 143.335 32.595 143.665 ;
        RECT 33.460 143.605 33.860 144.405 ;
        RECT 34.260 144.115 34.530 144.575 ;
        RECT 34.700 143.945 34.985 144.405 ;
        RECT 26.075 142.025 31.420 142.460 ;
        RECT 31.590 142.195 31.975 143.165 ;
        RECT 32.145 142.875 32.595 143.335 ;
        RECT 32.765 143.045 33.860 143.605 ;
        RECT 32.145 142.655 33.270 142.875 ;
        RECT 32.145 142.025 32.470 142.485 ;
        RECT 32.990 142.195 33.270 142.655 ;
        RECT 33.460 142.195 33.860 143.045 ;
        RECT 34.030 143.775 34.985 143.945 ;
        RECT 35.730 143.805 39.240 144.575 ;
        RECT 39.415 144.030 44.760 144.575 ;
        RECT 34.030 142.875 34.240 143.775 ;
        RECT 34.410 143.045 35.100 143.605 ;
        RECT 35.730 143.115 37.420 143.635 ;
        RECT 37.590 143.285 39.240 143.805 ;
        RECT 34.030 142.655 34.985 142.875 ;
        RECT 34.260 142.025 34.530 142.485 ;
        RECT 34.700 142.195 34.985 142.655 ;
        RECT 35.730 142.025 39.240 143.115 ;
        RECT 41.005 142.460 41.355 143.710 ;
        RECT 42.835 143.200 43.175 144.030 ;
        RECT 44.970 143.755 45.200 144.575 ;
        RECT 45.370 143.775 45.700 144.405 ;
        RECT 44.950 143.335 45.280 143.585 ;
        RECT 45.450 143.175 45.700 143.775 ;
        RECT 45.870 143.755 46.080 144.575 ;
        RECT 46.350 143.755 46.580 144.575 ;
        RECT 46.750 143.775 47.080 144.405 ;
        RECT 46.330 143.335 46.660 143.585 ;
        RECT 46.830 143.175 47.080 143.775 ;
        RECT 47.250 143.755 47.460 144.575 ;
        RECT 47.690 143.850 47.980 144.575 ;
        RECT 48.985 144.235 49.240 144.395 ;
        RECT 48.900 144.065 49.240 144.235 ;
        RECT 49.420 144.115 49.705 144.575 ;
        RECT 48.985 143.865 49.240 144.065 ;
        RECT 39.415 142.025 44.760 142.460 ;
        RECT 44.970 142.025 45.200 143.165 ;
        RECT 45.370 142.195 45.700 143.175 ;
        RECT 45.870 142.025 46.080 143.165 ;
        RECT 46.350 142.025 46.580 143.165 ;
        RECT 46.750 142.195 47.080 143.175 ;
        RECT 47.250 142.025 47.460 143.165 ;
        RECT 47.690 142.025 47.980 143.190 ;
        RECT 48.985 143.005 49.165 143.865 ;
        RECT 49.885 143.665 50.135 144.315 ;
        RECT 49.335 143.335 50.135 143.665 ;
        RECT 48.985 142.335 49.240 143.005 ;
        RECT 49.420 142.025 49.705 142.825 ;
        RECT 49.885 142.745 50.135 143.335 ;
        RECT 50.335 143.980 50.655 144.310 ;
        RECT 50.835 144.095 51.495 144.575 ;
        RECT 51.695 144.185 52.545 144.355 ;
        RECT 50.335 143.085 50.525 143.980 ;
        RECT 50.845 143.655 51.505 143.925 ;
        RECT 51.175 143.595 51.505 143.655 ;
        RECT 50.695 143.425 51.025 143.485 ;
        RECT 51.695 143.425 51.865 144.185 ;
        RECT 53.105 144.115 53.425 144.575 ;
        RECT 53.625 143.935 53.875 144.365 ;
        RECT 54.165 144.135 54.575 144.575 ;
        RECT 54.745 144.195 55.760 144.395 ;
        RECT 52.035 143.765 53.285 143.935 ;
        RECT 52.035 143.645 52.365 143.765 ;
        RECT 50.695 143.255 52.595 143.425 ;
        RECT 50.335 142.915 52.255 143.085 ;
        RECT 50.335 142.895 50.655 142.915 ;
        RECT 49.885 142.235 50.215 142.745 ;
        RECT 50.485 142.285 50.655 142.895 ;
        RECT 52.425 142.745 52.595 143.255 ;
        RECT 52.765 143.185 52.945 143.595 ;
        RECT 53.115 143.005 53.285 143.765 ;
        RECT 50.825 142.025 51.155 142.715 ;
        RECT 51.385 142.575 52.595 142.745 ;
        RECT 52.765 142.695 53.285 143.005 ;
        RECT 53.455 143.595 53.875 143.935 ;
        RECT 54.165 143.595 54.575 143.925 ;
        RECT 53.455 142.825 53.645 143.595 ;
        RECT 54.745 143.465 54.915 144.195 ;
        RECT 56.060 144.025 56.230 144.355 ;
        RECT 56.400 144.195 56.730 144.575 ;
        RECT 55.085 143.645 55.435 144.015 ;
        RECT 54.745 143.425 55.165 143.465 ;
        RECT 53.815 143.255 55.165 143.425 ;
        RECT 53.815 143.095 54.065 143.255 ;
        RECT 54.575 142.825 54.825 143.085 ;
        RECT 53.455 142.575 54.825 142.825 ;
        RECT 51.385 142.285 51.625 142.575 ;
        RECT 52.425 142.495 52.595 142.575 ;
        RECT 51.825 142.025 52.245 142.405 ;
        RECT 52.425 142.245 53.055 142.495 ;
        RECT 53.525 142.025 53.855 142.405 ;
        RECT 54.025 142.285 54.195 142.575 ;
        RECT 54.995 142.410 55.165 143.255 ;
        RECT 55.615 143.085 55.835 143.955 ;
        RECT 56.060 143.835 56.755 144.025 ;
        RECT 55.335 142.705 55.835 143.085 ;
        RECT 56.005 143.035 56.415 143.655 ;
        RECT 56.585 142.865 56.755 143.835 ;
        RECT 56.060 142.695 56.755 142.865 ;
        RECT 54.375 142.025 54.755 142.405 ;
        RECT 54.995 142.240 55.825 142.410 ;
        RECT 56.060 142.195 56.230 142.695 ;
        RECT 56.400 142.025 56.730 142.525 ;
        RECT 56.945 142.195 57.170 144.315 ;
        RECT 57.340 144.195 57.670 144.575 ;
        RECT 57.840 144.025 58.010 144.315 ;
        RECT 57.345 143.855 58.010 144.025 ;
        RECT 57.345 142.865 57.575 143.855 ;
        RECT 58.270 143.825 59.480 144.575 ;
        RECT 57.745 143.035 58.095 143.685 ;
        RECT 58.270 143.115 58.790 143.655 ;
        RECT 58.960 143.285 59.480 143.825 ;
        RECT 59.655 143.865 59.910 144.395 ;
        RECT 60.080 144.115 60.385 144.575 ;
        RECT 60.630 144.195 61.700 144.365 ;
        RECT 59.655 143.215 59.865 143.865 ;
        RECT 60.630 143.840 60.950 144.195 ;
        RECT 60.625 143.665 60.950 143.840 ;
        RECT 60.035 143.365 60.950 143.665 ;
        RECT 61.120 143.625 61.360 144.025 ;
        RECT 61.530 143.965 61.700 144.195 ;
        RECT 61.870 144.135 62.060 144.575 ;
        RECT 62.230 144.125 63.180 144.405 ;
        RECT 63.400 144.215 63.750 144.385 ;
        RECT 61.530 143.795 62.060 143.965 ;
        RECT 60.035 143.335 60.775 143.365 ;
        RECT 57.345 142.695 58.010 142.865 ;
        RECT 57.340 142.025 57.670 142.525 ;
        RECT 57.840 142.195 58.010 142.695 ;
        RECT 58.270 142.025 59.480 143.115 ;
        RECT 59.655 142.335 59.910 143.215 ;
        RECT 60.080 142.025 60.385 143.165 ;
        RECT 60.605 142.745 60.775 143.335 ;
        RECT 61.120 143.255 61.660 143.625 ;
        RECT 61.840 143.515 62.060 143.795 ;
        RECT 62.230 143.345 62.400 144.125 ;
        RECT 61.995 143.175 62.400 143.345 ;
        RECT 62.570 143.335 62.920 143.955 ;
        RECT 61.995 143.085 62.165 143.175 ;
        RECT 63.090 143.165 63.300 143.955 ;
        RECT 60.945 142.915 62.165 143.085 ;
        RECT 62.625 143.005 63.300 143.165 ;
        RECT 60.605 142.575 61.405 142.745 ;
        RECT 60.725 142.025 61.055 142.405 ;
        RECT 61.235 142.285 61.405 142.575 ;
        RECT 61.995 142.535 62.165 142.915 ;
        RECT 62.335 142.995 63.300 143.005 ;
        RECT 63.490 143.825 63.750 144.215 ;
        RECT 63.960 144.115 64.290 144.575 ;
        RECT 65.165 144.185 66.020 144.355 ;
        RECT 66.225 144.185 66.720 144.355 ;
        RECT 66.890 144.215 67.220 144.575 ;
        RECT 63.490 143.135 63.660 143.825 ;
        RECT 63.830 143.475 64.000 143.655 ;
        RECT 64.170 143.645 64.960 143.895 ;
        RECT 65.165 143.475 65.335 144.185 ;
        RECT 65.505 143.675 65.860 143.895 ;
        RECT 63.830 143.305 65.520 143.475 ;
        RECT 62.335 142.705 62.795 142.995 ;
        RECT 63.490 142.965 64.990 143.135 ;
        RECT 63.490 142.825 63.660 142.965 ;
        RECT 63.100 142.655 63.660 142.825 ;
        RECT 61.575 142.025 61.825 142.485 ;
        RECT 61.995 142.195 62.865 142.535 ;
        RECT 63.100 142.195 63.270 142.655 ;
        RECT 64.105 142.625 65.180 142.795 ;
        RECT 63.440 142.025 63.810 142.485 ;
        RECT 64.105 142.285 64.275 142.625 ;
        RECT 64.445 142.025 64.775 142.455 ;
        RECT 65.010 142.285 65.180 142.625 ;
        RECT 65.350 142.525 65.520 143.305 ;
        RECT 65.690 143.085 65.860 143.675 ;
        RECT 66.030 143.275 66.380 143.895 ;
        RECT 65.690 142.695 66.155 143.085 ;
        RECT 66.550 142.825 66.720 144.185 ;
        RECT 66.890 142.995 67.350 144.045 ;
        RECT 66.325 142.655 66.720 142.825 ;
        RECT 66.325 142.525 66.495 142.655 ;
        RECT 65.350 142.195 66.030 142.525 ;
        RECT 66.245 142.195 66.495 142.525 ;
        RECT 66.665 142.025 66.915 142.485 ;
        RECT 67.085 142.210 67.410 142.995 ;
        RECT 67.580 142.195 67.750 144.315 ;
        RECT 67.920 144.195 68.250 144.575 ;
        RECT 68.420 144.025 68.675 144.315 ;
        RECT 67.925 143.855 68.675 144.025 ;
        RECT 67.925 142.865 68.155 143.855 ;
        RECT 69.585 143.765 69.830 144.370 ;
        RECT 70.050 144.040 70.560 144.575 ;
        RECT 68.325 143.035 68.675 143.685 ;
        RECT 69.310 143.595 70.540 143.765 ;
        RECT 67.925 142.695 68.675 142.865 ;
        RECT 67.920 142.025 68.250 142.525 ;
        RECT 68.420 142.195 68.675 142.695 ;
        RECT 69.310 142.785 69.650 143.595 ;
        RECT 69.820 143.030 70.570 143.220 ;
        RECT 69.310 142.375 69.825 142.785 ;
        RECT 70.060 142.025 70.230 142.785 ;
        RECT 70.400 142.365 70.570 143.030 ;
        RECT 70.740 143.045 70.930 144.405 ;
        RECT 71.100 144.235 71.375 144.405 ;
        RECT 71.100 144.065 71.380 144.235 ;
        RECT 71.100 143.245 71.375 144.065 ;
        RECT 71.565 144.040 72.095 144.405 ;
        RECT 72.520 144.175 72.850 144.575 ;
        RECT 71.920 144.005 72.095 144.040 ;
        RECT 71.580 143.045 71.750 143.845 ;
        RECT 70.740 142.875 71.750 143.045 ;
        RECT 71.920 143.835 72.850 144.005 ;
        RECT 73.020 143.835 73.275 144.405 ;
        RECT 73.450 143.850 73.740 144.575 ;
        RECT 74.000 144.025 74.170 144.315 ;
        RECT 74.340 144.195 74.670 144.575 ;
        RECT 74.000 143.855 74.665 144.025 ;
        RECT 71.920 142.705 72.090 143.835 ;
        RECT 72.680 143.665 72.850 143.835 ;
        RECT 70.965 142.535 72.090 142.705 ;
        RECT 72.260 143.335 72.455 143.665 ;
        RECT 72.680 143.335 72.935 143.665 ;
        RECT 72.260 142.365 72.430 143.335 ;
        RECT 73.105 143.165 73.275 143.835 ;
        RECT 70.400 142.195 72.430 142.365 ;
        RECT 72.600 142.025 72.770 143.165 ;
        RECT 72.940 142.195 73.275 143.165 ;
        RECT 73.450 142.025 73.740 143.190 ;
        RECT 73.915 143.035 74.265 143.685 ;
        RECT 74.435 142.865 74.665 143.855 ;
        RECT 74.000 142.695 74.665 142.865 ;
        RECT 74.000 142.195 74.170 142.695 ;
        RECT 74.340 142.025 74.670 142.525 ;
        RECT 74.840 142.195 75.065 144.315 ;
        RECT 75.280 144.195 75.610 144.575 ;
        RECT 75.780 144.025 75.950 144.355 ;
        RECT 76.250 144.195 77.265 144.395 ;
        RECT 75.255 143.835 75.950 144.025 ;
        RECT 75.255 142.865 75.425 143.835 ;
        RECT 75.595 143.035 76.005 143.655 ;
        RECT 76.175 143.085 76.395 143.955 ;
        RECT 76.575 143.645 76.925 144.015 ;
        RECT 77.095 143.465 77.265 144.195 ;
        RECT 77.435 144.135 77.845 144.575 ;
        RECT 78.135 143.935 78.385 144.365 ;
        RECT 78.585 144.115 78.905 144.575 ;
        RECT 79.465 144.185 80.315 144.355 ;
        RECT 77.435 143.595 77.845 143.925 ;
        RECT 78.135 143.595 78.555 143.935 ;
        RECT 76.845 143.425 77.265 143.465 ;
        RECT 76.845 143.255 78.195 143.425 ;
        RECT 75.255 142.695 75.950 142.865 ;
        RECT 76.175 142.705 76.675 143.085 ;
        RECT 75.280 142.025 75.610 142.525 ;
        RECT 75.780 142.195 75.950 142.695 ;
        RECT 76.845 142.410 77.015 143.255 ;
        RECT 77.945 143.095 78.195 143.255 ;
        RECT 77.185 142.825 77.435 143.085 ;
        RECT 78.365 142.825 78.555 143.595 ;
        RECT 77.185 142.575 78.555 142.825 ;
        RECT 78.725 143.765 79.975 143.935 ;
        RECT 78.725 143.005 78.895 143.765 ;
        RECT 79.645 143.645 79.975 143.765 ;
        RECT 79.065 143.185 79.245 143.595 ;
        RECT 80.145 143.425 80.315 144.185 ;
        RECT 80.515 144.095 81.175 144.575 ;
        RECT 81.355 143.980 81.675 144.310 ;
        RECT 80.505 143.655 81.165 143.925 ;
        RECT 80.505 143.595 80.835 143.655 ;
        RECT 80.985 143.425 81.315 143.485 ;
        RECT 79.415 143.255 81.315 143.425 ;
        RECT 78.725 142.695 79.245 143.005 ;
        RECT 79.415 142.745 79.585 143.255 ;
        RECT 81.485 143.085 81.675 143.980 ;
        RECT 79.755 142.915 81.675 143.085 ;
        RECT 81.355 142.895 81.675 142.915 ;
        RECT 81.875 143.665 82.125 144.315 ;
        RECT 82.305 144.115 82.590 144.575 ;
        RECT 82.770 143.865 83.025 144.395 ;
        RECT 84.500 144.215 86.570 144.405 ;
        RECT 86.800 144.215 87.130 144.575 ;
        RECT 87.660 144.215 87.990 144.575 ;
        RECT 88.520 144.215 88.850 144.575 ;
        RECT 89.100 144.215 91.170 144.405 ;
        RECT 91.400 144.215 91.730 144.575 ;
        RECT 92.260 144.215 92.590 144.575 ;
        RECT 93.120 144.215 93.450 144.575 ;
        RECT 85.450 144.195 86.570 144.215 ;
        RECT 90.050 144.195 91.170 144.215 ;
        RECT 81.875 143.335 82.675 143.665 ;
        RECT 79.415 142.575 80.625 142.745 ;
        RECT 76.185 142.240 77.015 142.410 ;
        RECT 77.255 142.025 77.635 142.405 ;
        RECT 77.815 142.285 77.985 142.575 ;
        RECT 79.415 142.495 79.585 142.575 ;
        RECT 78.155 142.025 78.485 142.405 ;
        RECT 78.955 142.245 79.585 142.495 ;
        RECT 79.765 142.025 80.185 142.405 ;
        RECT 80.385 142.285 80.625 142.575 ;
        RECT 80.855 142.025 81.185 142.715 ;
        RECT 81.355 142.285 81.525 142.895 ;
        RECT 81.875 142.745 82.125 143.335 ;
        RECT 82.845 143.005 83.025 143.865 ;
        RECT 81.795 142.235 82.125 142.745 ;
        RECT 82.305 142.025 82.590 142.825 ;
        RECT 82.770 142.535 83.025 143.005 ;
        RECT 84.490 142.690 84.780 143.665 ;
        RECT 84.950 143.120 85.280 143.990 ;
        RECT 85.450 143.770 85.640 144.195 ;
        RECT 88.160 144.025 88.350 144.145 ;
        RECT 85.810 143.815 88.350 144.025 ;
        RECT 88.520 143.585 88.860 143.895 ;
        RECT 85.450 143.295 86.310 143.585 ;
        RECT 86.770 143.305 87.740 143.585 ;
        RECT 87.910 143.415 88.860 143.585 ;
        RECT 87.965 143.365 88.860 143.415 ;
        RECT 84.950 142.950 87.560 143.120 ;
        RECT 82.770 142.365 83.110 142.535 ;
        RECT 82.770 142.335 83.025 142.365 ;
        RECT 84.520 142.025 84.780 142.485 ;
        RECT 84.950 142.195 85.210 142.950 ;
        RECT 85.380 142.025 85.710 142.745 ;
        RECT 85.880 142.195 86.070 142.950 ;
        RECT 86.240 142.025 86.570 142.745 ;
        RECT 86.800 142.365 87.060 142.560 ;
        RECT 87.230 142.535 87.560 142.950 ;
        RECT 87.730 142.965 88.850 143.135 ;
        RECT 87.730 142.365 87.920 142.965 ;
        RECT 86.800 142.195 87.920 142.365 ;
        RECT 88.090 142.025 88.420 142.795 ;
        RECT 88.590 142.195 88.850 142.965 ;
        RECT 89.090 142.690 89.380 143.665 ;
        RECT 89.550 143.120 89.880 143.990 ;
        RECT 90.050 143.770 90.240 144.195 ;
        RECT 92.760 144.025 92.950 144.145 ;
        RECT 90.410 143.815 92.950 144.025 ;
        RECT 93.120 143.585 93.460 143.895 ;
        RECT 93.750 143.755 93.960 144.575 ;
        RECT 94.130 143.775 94.460 144.405 ;
        RECT 90.050 143.295 90.910 143.585 ;
        RECT 91.370 143.305 92.340 143.585 ;
        RECT 92.510 143.415 93.460 143.585 ;
        RECT 92.565 143.365 93.460 143.415 ;
        RECT 94.130 143.175 94.380 143.775 ;
        RECT 94.630 143.755 94.860 144.575 ;
        RECT 95.345 143.765 95.590 144.370 ;
        RECT 95.810 144.040 96.320 144.575 ;
        RECT 95.070 143.595 96.300 143.765 ;
        RECT 94.550 143.335 94.880 143.585 ;
        RECT 89.550 142.950 92.160 143.120 ;
        RECT 89.120 142.025 89.380 142.485 ;
        RECT 89.550 142.195 89.810 142.950 ;
        RECT 89.980 142.025 90.310 142.745 ;
        RECT 90.480 142.195 90.670 142.950 ;
        RECT 90.840 142.025 91.170 142.745 ;
        RECT 91.400 142.365 91.660 142.560 ;
        RECT 91.830 142.535 92.160 142.950 ;
        RECT 92.330 142.965 93.450 143.135 ;
        RECT 92.330 142.365 92.520 142.965 ;
        RECT 91.400 142.195 92.520 142.365 ;
        RECT 92.690 142.025 93.020 142.795 ;
        RECT 93.190 142.195 93.450 142.965 ;
        RECT 93.750 142.025 93.960 143.165 ;
        RECT 94.130 142.195 94.460 143.175 ;
        RECT 94.630 142.025 94.860 143.165 ;
        RECT 95.070 142.785 95.410 143.595 ;
        RECT 95.580 143.030 96.330 143.220 ;
        RECT 95.070 142.375 95.585 142.785 ;
        RECT 95.820 142.025 95.990 142.785 ;
        RECT 96.160 142.365 96.330 143.030 ;
        RECT 96.500 143.045 96.690 144.405 ;
        RECT 96.860 144.235 97.135 144.405 ;
        RECT 96.860 144.065 97.140 144.235 ;
        RECT 96.860 143.245 97.135 144.065 ;
        RECT 97.325 144.040 97.855 144.405 ;
        RECT 98.280 144.175 98.610 144.575 ;
        RECT 97.680 144.005 97.855 144.040 ;
        RECT 97.340 143.045 97.510 143.845 ;
        RECT 96.500 142.875 97.510 143.045 ;
        RECT 97.680 143.835 98.610 144.005 ;
        RECT 98.780 143.835 99.035 144.405 ;
        RECT 99.210 143.850 99.500 144.575 ;
        RECT 99.760 144.025 99.930 144.315 ;
        RECT 100.100 144.195 100.430 144.575 ;
        RECT 99.760 143.855 100.425 144.025 ;
        RECT 97.680 142.705 97.850 143.835 ;
        RECT 98.440 143.665 98.610 143.835 ;
        RECT 96.725 142.535 97.850 142.705 ;
        RECT 98.020 143.335 98.215 143.665 ;
        RECT 98.440 143.335 98.695 143.665 ;
        RECT 98.020 142.365 98.190 143.335 ;
        RECT 98.865 143.165 99.035 143.835 ;
        RECT 96.160 142.195 98.190 142.365 ;
        RECT 98.360 142.025 98.530 143.165 ;
        RECT 98.700 142.195 99.035 143.165 ;
        RECT 99.210 142.025 99.500 143.190 ;
        RECT 99.675 143.035 100.025 143.685 ;
        RECT 100.195 142.865 100.425 143.855 ;
        RECT 99.760 142.695 100.425 142.865 ;
        RECT 99.760 142.195 99.930 142.695 ;
        RECT 100.100 142.025 100.430 142.525 ;
        RECT 100.600 142.195 100.825 144.315 ;
        RECT 101.040 144.195 101.370 144.575 ;
        RECT 101.540 144.025 101.710 144.355 ;
        RECT 102.010 144.195 103.025 144.395 ;
        RECT 101.015 143.835 101.710 144.025 ;
        RECT 101.015 142.865 101.185 143.835 ;
        RECT 101.355 143.035 101.765 143.655 ;
        RECT 101.935 143.085 102.155 143.955 ;
        RECT 102.335 143.645 102.685 144.015 ;
        RECT 102.855 143.465 103.025 144.195 ;
        RECT 103.195 144.135 103.605 144.575 ;
        RECT 103.895 143.935 104.145 144.365 ;
        RECT 104.345 144.115 104.665 144.575 ;
        RECT 105.225 144.185 106.075 144.355 ;
        RECT 103.195 143.595 103.605 143.925 ;
        RECT 103.895 143.595 104.315 143.935 ;
        RECT 102.605 143.425 103.025 143.465 ;
        RECT 102.605 143.255 103.955 143.425 ;
        RECT 101.015 142.695 101.710 142.865 ;
        RECT 101.935 142.705 102.435 143.085 ;
        RECT 101.040 142.025 101.370 142.525 ;
        RECT 101.540 142.195 101.710 142.695 ;
        RECT 102.605 142.410 102.775 143.255 ;
        RECT 103.705 143.095 103.955 143.255 ;
        RECT 102.945 142.825 103.195 143.085 ;
        RECT 104.125 142.825 104.315 143.595 ;
        RECT 102.945 142.575 104.315 142.825 ;
        RECT 104.485 143.765 105.735 143.935 ;
        RECT 104.485 143.005 104.655 143.765 ;
        RECT 105.405 143.645 105.735 143.765 ;
        RECT 104.825 143.185 105.005 143.595 ;
        RECT 105.905 143.425 106.075 144.185 ;
        RECT 106.275 144.095 106.935 144.575 ;
        RECT 107.115 143.980 107.435 144.310 ;
        RECT 106.265 143.655 106.925 143.925 ;
        RECT 106.265 143.595 106.595 143.655 ;
        RECT 106.745 143.425 107.075 143.485 ;
        RECT 105.175 143.255 107.075 143.425 ;
        RECT 104.485 142.695 105.005 143.005 ;
        RECT 105.175 142.745 105.345 143.255 ;
        RECT 107.245 143.085 107.435 143.980 ;
        RECT 105.515 142.915 107.435 143.085 ;
        RECT 107.115 142.895 107.435 142.915 ;
        RECT 107.635 143.665 107.885 144.315 ;
        RECT 108.065 144.115 108.350 144.575 ;
        RECT 108.530 144.235 108.785 144.395 ;
        RECT 108.530 144.065 108.870 144.235 ;
        RECT 108.530 143.865 108.785 144.065 ;
        RECT 107.635 143.335 108.435 143.665 ;
        RECT 105.175 142.575 106.385 142.745 ;
        RECT 101.945 142.240 102.775 142.410 ;
        RECT 103.015 142.025 103.395 142.405 ;
        RECT 103.575 142.285 103.745 142.575 ;
        RECT 105.175 142.495 105.345 142.575 ;
        RECT 103.915 142.025 104.245 142.405 ;
        RECT 104.715 142.245 105.345 142.495 ;
        RECT 105.525 142.025 105.945 142.405 ;
        RECT 106.145 142.285 106.385 142.575 ;
        RECT 106.615 142.025 106.945 142.715 ;
        RECT 107.115 142.285 107.285 142.895 ;
        RECT 107.635 142.745 107.885 143.335 ;
        RECT 108.605 143.005 108.785 143.865 ;
        RECT 107.555 142.235 107.885 142.745 ;
        RECT 108.065 142.025 108.350 142.825 ;
        RECT 108.530 142.335 108.785 143.005 ;
        RECT 109.790 143.900 110.050 144.405 ;
        RECT 110.230 144.195 110.560 144.575 ;
        RECT 110.740 144.025 110.910 144.405 ;
        RECT 109.790 143.100 109.960 143.900 ;
        RECT 110.245 143.855 110.910 144.025 ;
        RECT 110.245 143.600 110.415 143.855 ;
        RECT 111.170 143.825 112.380 144.575 ;
        RECT 110.130 143.270 110.415 143.600 ;
        RECT 110.650 143.305 110.980 143.675 ;
        RECT 110.245 143.125 110.415 143.270 ;
        RECT 109.790 142.195 110.060 143.100 ;
        RECT 110.245 142.955 110.910 143.125 ;
        RECT 110.230 142.025 110.560 142.785 ;
        RECT 110.740 142.195 110.910 142.955 ;
        RECT 111.170 143.115 111.690 143.655 ;
        RECT 111.860 143.285 112.380 143.825 ;
        RECT 111.170 142.025 112.380 143.115 ;
        RECT 18.165 141.855 112.465 142.025 ;
        RECT 18.250 140.765 19.460 141.855 ;
        RECT 18.250 140.055 18.770 140.595 ;
        RECT 18.940 140.225 19.460 140.765 ;
        RECT 20.550 140.765 24.060 141.855 ;
        RECT 24.235 141.420 29.580 141.855 ;
        RECT 20.550 140.245 22.240 140.765 ;
        RECT 22.410 140.075 24.060 140.595 ;
        RECT 25.825 140.170 26.175 141.420 ;
        RECT 29.810 140.715 30.020 141.855 ;
        RECT 30.190 140.705 30.520 141.685 ;
        RECT 30.690 140.715 30.920 141.855 ;
        RECT 31.130 140.765 34.640 141.855 ;
        RECT 18.250 139.305 19.460 140.055 ;
        RECT 20.550 139.305 24.060 140.075 ;
        RECT 27.655 139.850 27.995 140.680 ;
        RECT 24.235 139.305 29.580 139.850 ;
        RECT 29.810 139.305 30.020 140.125 ;
        RECT 30.190 140.105 30.440 140.705 ;
        RECT 30.610 140.295 30.940 140.545 ;
        RECT 31.130 140.245 32.820 140.765 ;
        RECT 34.810 140.690 35.100 141.855 ;
        RECT 35.790 140.715 36.000 141.855 ;
        RECT 36.170 140.705 36.500 141.685 ;
        RECT 36.670 140.715 36.900 141.855 ;
        RECT 37.570 140.715 37.910 141.685 ;
        RECT 38.080 140.715 38.250 141.855 ;
        RECT 38.520 141.055 38.770 141.855 ;
        RECT 39.415 140.885 39.745 141.685 ;
        RECT 40.045 141.055 40.375 141.855 ;
        RECT 40.545 140.885 40.875 141.685 ;
        RECT 38.440 140.715 40.875 140.885 ;
        RECT 41.250 140.715 41.590 141.685 ;
        RECT 41.760 140.715 41.930 141.855 ;
        RECT 42.200 141.055 42.450 141.855 ;
        RECT 43.095 140.885 43.425 141.685 ;
        RECT 43.725 141.055 44.055 141.855 ;
        RECT 44.225 140.885 44.555 141.685 ;
        RECT 42.120 140.715 44.555 140.885 ;
        RECT 45.305 140.875 45.560 141.545 ;
        RECT 45.740 141.055 46.025 141.855 ;
        RECT 46.205 141.135 46.535 141.645 ;
        RECT 30.190 139.475 30.520 140.105 ;
        RECT 30.690 139.305 30.920 140.125 ;
        RECT 32.990 140.075 34.640 140.595 ;
        RECT 31.130 139.305 34.640 140.075 ;
        RECT 34.810 139.305 35.100 140.030 ;
        RECT 35.790 139.305 36.000 140.125 ;
        RECT 36.170 140.105 36.420 140.705 ;
        RECT 36.590 140.295 36.920 140.545 ;
        RECT 37.570 140.155 37.745 140.715 ;
        RECT 38.440 140.465 38.610 140.715 ;
        RECT 37.915 140.295 38.610 140.465 ;
        RECT 38.785 140.295 39.205 140.495 ;
        RECT 39.375 140.295 39.705 140.495 ;
        RECT 39.875 140.295 40.205 140.495 ;
        RECT 36.170 139.475 36.500 140.105 ;
        RECT 36.670 139.305 36.900 140.125 ;
        RECT 37.570 140.105 37.800 140.155 ;
        RECT 37.570 139.475 37.910 140.105 ;
        RECT 38.080 139.305 38.330 140.105 ;
        RECT 38.520 139.955 39.745 140.125 ;
        RECT 38.520 139.475 38.850 139.955 ;
        RECT 39.020 139.305 39.245 139.765 ;
        RECT 39.415 139.475 39.745 139.955 ;
        RECT 40.375 140.085 40.545 140.715 ;
        RECT 40.730 140.295 41.080 140.545 ;
        RECT 41.250 140.105 41.425 140.715 ;
        RECT 42.120 140.465 42.290 140.715 ;
        RECT 41.595 140.295 42.290 140.465 ;
        RECT 42.465 140.295 42.885 140.495 ;
        RECT 43.055 140.295 43.385 140.495 ;
        RECT 43.555 140.295 43.885 140.495 ;
        RECT 40.375 139.475 40.875 140.085 ;
        RECT 41.250 139.475 41.590 140.105 ;
        RECT 41.760 139.305 42.010 140.105 ;
        RECT 42.200 139.955 43.425 140.125 ;
        RECT 42.200 139.475 42.530 139.955 ;
        RECT 42.700 139.305 42.925 139.765 ;
        RECT 43.095 139.475 43.425 139.955 ;
        RECT 44.055 140.085 44.225 140.715 ;
        RECT 44.410 140.295 44.760 140.545 ;
        RECT 45.305 140.155 45.485 140.875 ;
        RECT 46.205 140.545 46.455 141.135 ;
        RECT 46.805 140.985 46.975 141.595 ;
        RECT 47.145 141.165 47.475 141.855 ;
        RECT 47.705 141.305 47.945 141.595 ;
        RECT 48.145 141.475 48.565 141.855 ;
        RECT 48.745 141.385 49.375 141.635 ;
        RECT 49.845 141.475 50.175 141.855 ;
        RECT 48.745 141.305 48.915 141.385 ;
        RECT 50.345 141.305 50.515 141.595 ;
        RECT 50.695 141.475 51.075 141.855 ;
        RECT 51.315 141.470 52.145 141.640 ;
        RECT 47.705 141.135 48.915 141.305 ;
        RECT 45.655 140.215 46.455 140.545 ;
        RECT 44.055 139.475 44.555 140.085 ;
        RECT 45.220 140.015 45.485 140.155 ;
        RECT 45.220 139.985 45.560 140.015 ;
        RECT 45.305 139.485 45.560 139.985 ;
        RECT 45.740 139.305 46.025 139.765 ;
        RECT 46.205 139.565 46.455 140.215 ;
        RECT 46.655 140.965 46.975 140.985 ;
        RECT 46.655 140.795 48.575 140.965 ;
        RECT 46.655 139.900 46.845 140.795 ;
        RECT 48.745 140.625 48.915 141.135 ;
        RECT 49.085 140.875 49.605 141.185 ;
        RECT 47.015 140.455 48.915 140.625 ;
        RECT 47.015 140.395 47.345 140.455 ;
        RECT 47.495 140.225 47.825 140.285 ;
        RECT 47.165 139.955 47.825 140.225 ;
        RECT 46.655 139.570 46.975 139.900 ;
        RECT 47.155 139.305 47.815 139.785 ;
        RECT 48.015 139.695 48.185 140.455 ;
        RECT 49.085 140.285 49.265 140.695 ;
        RECT 48.355 140.115 48.685 140.235 ;
        RECT 49.435 140.115 49.605 140.875 ;
        RECT 48.355 139.945 49.605 140.115 ;
        RECT 49.775 141.055 51.145 141.305 ;
        RECT 49.775 140.285 49.965 141.055 ;
        RECT 50.895 140.795 51.145 141.055 ;
        RECT 50.135 140.625 50.385 140.785 ;
        RECT 51.315 140.625 51.485 141.470 ;
        RECT 52.380 141.185 52.550 141.685 ;
        RECT 52.720 141.355 53.050 141.855 ;
        RECT 51.655 140.795 52.155 141.175 ;
        RECT 52.380 141.015 53.075 141.185 ;
        RECT 50.135 140.455 51.485 140.625 ;
        RECT 51.065 140.415 51.485 140.455 ;
        RECT 49.775 139.945 50.195 140.285 ;
        RECT 50.485 139.955 50.895 140.285 ;
        RECT 48.015 139.525 48.865 139.695 ;
        RECT 49.425 139.305 49.745 139.765 ;
        RECT 49.945 139.515 50.195 139.945 ;
        RECT 50.485 139.305 50.895 139.745 ;
        RECT 51.065 139.685 51.235 140.415 ;
        RECT 51.405 139.865 51.755 140.235 ;
        RECT 51.935 139.925 52.155 140.795 ;
        RECT 52.325 140.225 52.735 140.845 ;
        RECT 52.905 140.045 53.075 141.015 ;
        RECT 52.380 139.855 53.075 140.045 ;
        RECT 51.065 139.485 52.080 139.685 ;
        RECT 52.380 139.525 52.550 139.855 ;
        RECT 52.720 139.305 53.050 139.685 ;
        RECT 53.265 139.565 53.490 141.685 ;
        RECT 53.660 141.355 53.990 141.855 ;
        RECT 54.160 141.185 54.330 141.685 ;
        RECT 53.665 141.015 54.330 141.185 ;
        RECT 53.665 140.025 53.895 141.015 ;
        RECT 54.065 140.195 54.415 140.845 ;
        RECT 54.595 140.715 54.930 141.685 ;
        RECT 55.100 140.715 55.270 141.855 ;
        RECT 55.440 141.515 57.470 141.685 ;
        RECT 54.595 140.045 54.765 140.715 ;
        RECT 55.440 140.545 55.610 141.515 ;
        RECT 54.935 140.215 55.190 140.545 ;
        RECT 55.415 140.215 55.610 140.545 ;
        RECT 55.780 141.175 56.905 141.345 ;
        RECT 55.020 140.045 55.190 140.215 ;
        RECT 55.780 140.045 55.950 141.175 ;
        RECT 53.665 139.855 54.330 140.025 ;
        RECT 53.660 139.305 53.990 139.685 ;
        RECT 54.160 139.565 54.330 139.855 ;
        RECT 54.595 139.475 54.850 140.045 ;
        RECT 55.020 139.875 55.950 140.045 ;
        RECT 56.120 140.835 57.130 141.005 ;
        RECT 56.120 140.035 56.290 140.835 ;
        RECT 55.775 139.840 55.950 139.875 ;
        RECT 55.020 139.305 55.350 139.705 ;
        RECT 55.775 139.475 56.305 139.840 ;
        RECT 56.495 139.815 56.770 140.635 ;
        RECT 56.490 139.645 56.770 139.815 ;
        RECT 56.495 139.475 56.770 139.645 ;
        RECT 56.940 139.475 57.130 140.835 ;
        RECT 57.300 140.850 57.470 141.515 ;
        RECT 57.640 141.095 57.810 141.855 ;
        RECT 58.045 141.095 58.560 141.505 ;
        RECT 57.300 140.660 58.050 140.850 ;
        RECT 58.220 140.285 58.560 141.095 ;
        RECT 58.790 140.715 59.000 141.855 ;
        RECT 57.330 140.115 58.560 140.285 ;
        RECT 59.170 140.705 59.500 141.685 ;
        RECT 59.670 140.715 59.900 141.855 ;
        RECT 57.310 139.305 57.820 139.840 ;
        RECT 58.040 139.510 58.285 140.115 ;
        RECT 58.790 139.305 59.000 140.125 ;
        RECT 59.170 140.105 59.420 140.705 ;
        RECT 60.570 140.690 60.860 141.855 ;
        RECT 61.070 140.715 61.300 141.855 ;
        RECT 61.470 140.705 61.800 141.685 ;
        RECT 61.970 140.715 62.180 141.855 ;
        RECT 62.410 141.095 62.925 141.505 ;
        RECT 63.160 141.095 63.330 141.855 ;
        RECT 63.500 141.515 65.530 141.685 ;
        RECT 59.590 140.295 59.920 140.545 ;
        RECT 61.050 140.295 61.380 140.545 ;
        RECT 59.170 139.475 59.500 140.105 ;
        RECT 59.670 139.305 59.900 140.125 ;
        RECT 60.570 139.305 60.860 140.030 ;
        RECT 61.070 139.305 61.300 140.125 ;
        RECT 61.550 140.105 61.800 140.705 ;
        RECT 62.410 140.285 62.750 141.095 ;
        RECT 63.500 140.850 63.670 141.515 ;
        RECT 64.065 141.175 65.190 141.345 ;
        RECT 62.920 140.660 63.670 140.850 ;
        RECT 63.840 140.835 64.850 141.005 ;
        RECT 61.470 139.475 61.800 140.105 ;
        RECT 61.970 139.305 62.180 140.125 ;
        RECT 62.410 140.115 63.640 140.285 ;
        RECT 62.685 139.510 62.930 140.115 ;
        RECT 63.150 139.305 63.660 139.840 ;
        RECT 63.840 139.475 64.030 140.835 ;
        RECT 64.200 139.815 64.475 140.635 ;
        RECT 64.680 140.035 64.850 140.835 ;
        RECT 65.020 140.045 65.190 141.175 ;
        RECT 65.360 140.545 65.530 141.515 ;
        RECT 65.700 140.715 65.870 141.855 ;
        RECT 66.040 140.715 66.375 141.685 ;
        RECT 65.360 140.215 65.555 140.545 ;
        RECT 65.780 140.215 66.035 140.545 ;
        RECT 65.780 140.045 65.950 140.215 ;
        RECT 66.205 140.045 66.375 140.715 ;
        RECT 66.550 140.765 67.760 141.855 ;
        RECT 68.305 140.875 68.560 141.545 ;
        RECT 68.740 141.055 69.025 141.855 ;
        RECT 69.205 141.135 69.535 141.645 ;
        RECT 68.305 140.835 68.485 140.875 ;
        RECT 66.550 140.225 67.070 140.765 ;
        RECT 68.220 140.665 68.485 140.835 ;
        RECT 67.240 140.055 67.760 140.595 ;
        RECT 65.020 139.875 65.950 140.045 ;
        RECT 65.020 139.840 65.195 139.875 ;
        RECT 64.200 139.645 64.480 139.815 ;
        RECT 64.200 139.475 64.475 139.645 ;
        RECT 64.665 139.475 65.195 139.840 ;
        RECT 65.620 139.305 65.950 139.705 ;
        RECT 66.120 139.475 66.375 140.045 ;
        RECT 66.550 139.305 67.760 140.055 ;
        RECT 68.305 140.015 68.485 140.665 ;
        RECT 69.205 140.545 69.455 141.135 ;
        RECT 69.805 140.985 69.975 141.595 ;
        RECT 70.145 141.165 70.475 141.855 ;
        RECT 70.705 141.305 70.945 141.595 ;
        RECT 71.145 141.475 71.565 141.855 ;
        RECT 71.745 141.385 72.375 141.635 ;
        RECT 72.845 141.475 73.175 141.855 ;
        RECT 71.745 141.305 71.915 141.385 ;
        RECT 73.345 141.305 73.515 141.595 ;
        RECT 73.695 141.475 74.075 141.855 ;
        RECT 74.315 141.470 75.145 141.640 ;
        RECT 70.705 141.135 71.915 141.305 ;
        RECT 68.655 140.215 69.455 140.545 ;
        RECT 68.305 139.485 68.560 140.015 ;
        RECT 68.740 139.305 69.025 139.765 ;
        RECT 69.205 139.565 69.455 140.215 ;
        RECT 69.655 140.965 69.975 140.985 ;
        RECT 69.655 140.795 71.575 140.965 ;
        RECT 69.655 139.900 69.845 140.795 ;
        RECT 71.745 140.625 71.915 141.135 ;
        RECT 72.085 140.875 72.605 141.185 ;
        RECT 70.015 140.455 71.915 140.625 ;
        RECT 70.015 140.395 70.345 140.455 ;
        RECT 70.495 140.225 70.825 140.285 ;
        RECT 70.165 139.955 70.825 140.225 ;
        RECT 69.655 139.570 69.975 139.900 ;
        RECT 70.155 139.305 70.815 139.785 ;
        RECT 71.015 139.695 71.185 140.455 ;
        RECT 72.085 140.285 72.265 140.695 ;
        RECT 71.355 140.115 71.685 140.235 ;
        RECT 72.435 140.115 72.605 140.875 ;
        RECT 71.355 139.945 72.605 140.115 ;
        RECT 72.775 141.055 74.145 141.305 ;
        RECT 72.775 140.285 72.965 141.055 ;
        RECT 73.895 140.795 74.145 141.055 ;
        RECT 73.135 140.625 73.385 140.785 ;
        RECT 74.315 140.625 74.485 141.470 ;
        RECT 75.380 141.185 75.550 141.685 ;
        RECT 75.720 141.355 76.050 141.855 ;
        RECT 74.655 140.795 75.155 141.175 ;
        RECT 75.380 141.015 76.075 141.185 ;
        RECT 73.135 140.455 74.485 140.625 ;
        RECT 74.065 140.415 74.485 140.455 ;
        RECT 72.775 139.945 73.195 140.285 ;
        RECT 73.485 139.955 73.895 140.285 ;
        RECT 71.015 139.525 71.865 139.695 ;
        RECT 72.425 139.305 72.745 139.765 ;
        RECT 72.945 139.515 73.195 139.945 ;
        RECT 73.485 139.305 73.895 139.745 ;
        RECT 74.065 139.685 74.235 140.415 ;
        RECT 74.405 139.865 74.755 140.235 ;
        RECT 74.935 139.925 75.155 140.795 ;
        RECT 75.325 140.225 75.735 140.845 ;
        RECT 75.905 140.045 76.075 141.015 ;
        RECT 75.380 139.855 76.075 140.045 ;
        RECT 74.065 139.485 75.080 139.685 ;
        RECT 75.380 139.525 75.550 139.855 ;
        RECT 75.720 139.305 76.050 139.685 ;
        RECT 76.265 139.565 76.490 141.685 ;
        RECT 76.660 141.355 76.990 141.855 ;
        RECT 77.160 141.185 77.330 141.685 ;
        RECT 76.665 141.015 77.330 141.185 ;
        RECT 78.165 141.225 78.450 141.685 ;
        RECT 78.620 141.395 78.890 141.855 ;
        RECT 76.665 140.025 76.895 141.015 ;
        RECT 78.165 141.005 79.120 141.225 ;
        RECT 77.065 140.195 77.415 140.845 ;
        RECT 78.050 140.275 78.740 140.835 ;
        RECT 78.910 140.105 79.120 141.005 ;
        RECT 76.665 139.855 77.330 140.025 ;
        RECT 76.660 139.305 76.990 139.685 ;
        RECT 77.160 139.565 77.330 139.855 ;
        RECT 78.165 139.935 79.120 140.105 ;
        RECT 79.290 140.835 79.690 141.685 ;
        RECT 79.880 141.225 80.160 141.685 ;
        RECT 80.680 141.395 81.005 141.855 ;
        RECT 79.880 141.005 81.005 141.225 ;
        RECT 79.290 140.275 80.385 140.835 ;
        RECT 80.555 140.545 81.005 141.005 ;
        RECT 81.175 140.715 81.560 141.685 ;
        RECT 81.790 140.715 82.000 141.855 ;
        RECT 78.165 139.475 78.450 139.935 ;
        RECT 78.620 139.305 78.890 139.765 ;
        RECT 79.290 139.475 79.690 140.275 ;
        RECT 80.555 140.215 81.110 140.545 ;
        RECT 80.555 140.105 81.005 140.215 ;
        RECT 79.880 139.935 81.005 140.105 ;
        RECT 81.280 140.045 81.560 140.715 ;
        RECT 82.170 140.705 82.500 141.685 ;
        RECT 82.670 140.715 82.900 141.855 ;
        RECT 83.115 141.465 83.450 141.685 ;
        RECT 84.455 141.475 84.810 141.855 ;
        RECT 83.115 140.845 83.370 141.465 ;
        RECT 83.620 141.305 83.850 141.345 ;
        RECT 84.980 141.305 85.230 141.685 ;
        RECT 83.620 141.105 85.230 141.305 ;
        RECT 83.620 141.015 83.805 141.105 ;
        RECT 84.395 141.095 85.230 141.105 ;
        RECT 85.480 141.075 85.730 141.855 ;
        RECT 85.900 141.005 86.160 141.685 ;
        RECT 83.960 140.905 84.290 140.935 ;
        RECT 83.960 140.845 85.760 140.905 ;
        RECT 83.115 140.735 85.820 140.845 ;
        RECT 79.880 139.475 80.160 139.935 ;
        RECT 80.680 139.305 81.005 139.765 ;
        RECT 81.175 139.475 81.560 140.045 ;
        RECT 81.790 139.305 82.000 140.125 ;
        RECT 82.170 140.105 82.420 140.705 ;
        RECT 83.115 140.675 84.290 140.735 ;
        RECT 85.620 140.700 85.820 140.735 ;
        RECT 82.590 140.295 82.920 140.545 ;
        RECT 83.110 140.295 83.600 140.495 ;
        RECT 83.790 140.295 84.265 140.505 ;
        RECT 82.170 139.475 82.500 140.105 ;
        RECT 82.670 139.305 82.900 140.125 ;
        RECT 83.115 139.305 83.570 140.070 ;
        RECT 84.045 139.895 84.265 140.295 ;
        RECT 84.510 140.295 84.840 140.505 ;
        RECT 84.510 139.895 84.720 140.295 ;
        RECT 85.010 140.260 85.420 140.565 ;
        RECT 85.650 140.125 85.820 140.700 ;
        RECT 85.550 140.005 85.820 140.125 ;
        RECT 84.975 139.960 85.820 140.005 ;
        RECT 84.975 139.835 85.730 139.960 ;
        RECT 84.975 139.685 85.145 139.835 ;
        RECT 85.990 139.815 86.160 141.005 ;
        RECT 86.330 140.690 86.620 141.855 ;
        RECT 86.990 141.185 87.270 141.855 ;
        RECT 87.440 140.965 87.740 141.515 ;
        RECT 87.940 141.135 88.270 141.855 ;
        RECT 88.460 141.135 88.920 141.685 ;
        RECT 86.805 140.545 87.070 140.905 ;
        RECT 87.440 140.795 88.380 140.965 ;
        RECT 88.210 140.545 88.380 140.795 ;
        RECT 86.805 140.295 87.480 140.545 ;
        RECT 87.700 140.295 88.040 140.545 ;
        RECT 88.210 140.215 88.500 140.545 ;
        RECT 88.210 140.125 88.380 140.215 ;
        RECT 85.930 139.805 86.160 139.815 ;
        RECT 83.845 139.475 85.145 139.685 ;
        RECT 85.400 139.305 85.730 139.665 ;
        RECT 85.900 139.475 86.160 139.805 ;
        RECT 86.330 139.305 86.620 140.030 ;
        RECT 86.990 139.935 88.380 140.125 ;
        RECT 86.990 139.575 87.320 139.935 ;
        RECT 88.670 139.765 88.920 141.135 ;
        RECT 87.940 139.305 88.190 139.765 ;
        RECT 88.360 139.475 88.920 139.765 ;
        RECT 89.090 140.715 89.430 141.685 ;
        RECT 89.600 140.715 89.770 141.855 ;
        RECT 90.040 141.055 90.290 141.855 ;
        RECT 90.935 140.885 91.265 141.685 ;
        RECT 91.565 141.055 91.895 141.855 ;
        RECT 92.065 140.885 92.395 141.685 ;
        RECT 89.960 140.715 92.395 140.885 ;
        RECT 92.770 141.095 93.285 141.505 ;
        RECT 93.520 141.095 93.690 141.855 ;
        RECT 93.860 141.515 95.890 141.685 ;
        RECT 89.090 140.105 89.265 140.715 ;
        RECT 89.960 140.465 90.130 140.715 ;
        RECT 89.435 140.295 90.130 140.465 ;
        RECT 90.305 140.295 90.725 140.495 ;
        RECT 90.895 140.295 91.225 140.495 ;
        RECT 91.395 140.295 91.725 140.495 ;
        RECT 89.090 139.475 89.430 140.105 ;
        RECT 89.600 139.305 89.850 140.105 ;
        RECT 90.040 139.955 91.265 140.125 ;
        RECT 90.040 139.475 90.370 139.955 ;
        RECT 90.540 139.305 90.765 139.765 ;
        RECT 90.935 139.475 91.265 139.955 ;
        RECT 91.895 140.085 92.065 140.715 ;
        RECT 92.250 140.295 92.600 140.545 ;
        RECT 92.770 140.285 93.110 141.095 ;
        RECT 93.860 140.850 94.030 141.515 ;
        RECT 94.425 141.175 95.550 141.345 ;
        RECT 93.280 140.660 94.030 140.850 ;
        RECT 94.200 140.835 95.210 141.005 ;
        RECT 92.770 140.115 94.000 140.285 ;
        RECT 91.895 139.475 92.395 140.085 ;
        RECT 93.045 139.510 93.290 140.115 ;
        RECT 93.510 139.305 94.020 139.840 ;
        RECT 94.200 139.475 94.390 140.835 ;
        RECT 94.560 139.815 94.835 140.635 ;
        RECT 95.040 140.035 95.210 140.835 ;
        RECT 95.380 140.045 95.550 141.175 ;
        RECT 95.720 140.545 95.890 141.515 ;
        RECT 96.060 140.715 96.230 141.855 ;
        RECT 96.400 140.715 96.735 141.685 ;
        RECT 95.720 140.215 95.915 140.545 ;
        RECT 96.140 140.215 96.395 140.545 ;
        RECT 96.140 140.045 96.310 140.215 ;
        RECT 96.565 140.045 96.735 140.715 ;
        RECT 95.380 139.875 96.310 140.045 ;
        RECT 95.380 139.840 95.555 139.875 ;
        RECT 94.560 139.645 94.840 139.815 ;
        RECT 94.560 139.475 94.835 139.645 ;
        RECT 95.025 139.475 95.555 139.840 ;
        RECT 95.980 139.305 96.310 139.705 ;
        RECT 96.480 139.475 96.735 140.045 ;
        RECT 97.285 140.875 97.540 141.545 ;
        RECT 97.720 141.055 98.005 141.855 ;
        RECT 98.185 141.135 98.515 141.645 ;
        RECT 97.285 140.015 97.465 140.875 ;
        RECT 98.185 140.545 98.435 141.135 ;
        RECT 98.785 140.985 98.955 141.595 ;
        RECT 99.125 141.165 99.455 141.855 ;
        RECT 99.685 141.305 99.925 141.595 ;
        RECT 100.125 141.475 100.545 141.855 ;
        RECT 100.725 141.385 101.355 141.635 ;
        RECT 101.825 141.475 102.155 141.855 ;
        RECT 100.725 141.305 100.895 141.385 ;
        RECT 102.325 141.305 102.495 141.595 ;
        RECT 102.675 141.475 103.055 141.855 ;
        RECT 103.295 141.470 104.125 141.640 ;
        RECT 99.685 141.135 100.895 141.305 ;
        RECT 97.635 140.215 98.435 140.545 ;
        RECT 97.285 139.815 97.540 140.015 ;
        RECT 97.200 139.645 97.540 139.815 ;
        RECT 97.285 139.485 97.540 139.645 ;
        RECT 97.720 139.305 98.005 139.765 ;
        RECT 98.185 139.565 98.435 140.215 ;
        RECT 98.635 140.965 98.955 140.985 ;
        RECT 98.635 140.795 100.555 140.965 ;
        RECT 98.635 139.900 98.825 140.795 ;
        RECT 100.725 140.625 100.895 141.135 ;
        RECT 101.065 140.875 101.585 141.185 ;
        RECT 98.995 140.455 100.895 140.625 ;
        RECT 98.995 140.395 99.325 140.455 ;
        RECT 99.475 140.225 99.805 140.285 ;
        RECT 99.145 139.955 99.805 140.225 ;
        RECT 98.635 139.570 98.955 139.900 ;
        RECT 99.135 139.305 99.795 139.785 ;
        RECT 99.995 139.695 100.165 140.455 ;
        RECT 101.065 140.285 101.245 140.695 ;
        RECT 100.335 140.115 100.665 140.235 ;
        RECT 101.415 140.115 101.585 140.875 ;
        RECT 100.335 139.945 101.585 140.115 ;
        RECT 101.755 141.055 103.125 141.305 ;
        RECT 101.755 140.285 101.945 141.055 ;
        RECT 102.875 140.795 103.125 141.055 ;
        RECT 102.115 140.625 102.365 140.785 ;
        RECT 103.295 140.625 103.465 141.470 ;
        RECT 104.360 141.185 104.530 141.685 ;
        RECT 104.700 141.355 105.030 141.855 ;
        RECT 103.635 140.795 104.135 141.175 ;
        RECT 104.360 141.015 105.055 141.185 ;
        RECT 102.115 140.455 103.465 140.625 ;
        RECT 103.045 140.415 103.465 140.455 ;
        RECT 101.755 139.945 102.175 140.285 ;
        RECT 102.465 139.955 102.875 140.285 ;
        RECT 99.995 139.525 100.845 139.695 ;
        RECT 101.405 139.305 101.725 139.765 ;
        RECT 101.925 139.515 102.175 139.945 ;
        RECT 102.465 139.305 102.875 139.745 ;
        RECT 103.045 139.685 103.215 140.415 ;
        RECT 103.385 139.865 103.735 140.235 ;
        RECT 103.915 139.925 104.135 140.795 ;
        RECT 104.305 140.225 104.715 140.845 ;
        RECT 104.885 140.045 105.055 141.015 ;
        RECT 104.360 139.855 105.055 140.045 ;
        RECT 103.045 139.485 104.060 139.685 ;
        RECT 104.360 139.525 104.530 139.855 ;
        RECT 104.700 139.305 105.030 139.685 ;
        RECT 105.245 139.565 105.470 141.685 ;
        RECT 105.640 141.355 105.970 141.855 ;
        RECT 106.140 141.185 106.310 141.685 ;
        RECT 105.645 141.015 106.310 141.185 ;
        RECT 105.645 140.025 105.875 141.015 ;
        RECT 106.045 140.195 106.395 140.845 ;
        RECT 107.490 140.765 111.000 141.855 ;
        RECT 111.170 140.765 112.380 141.855 ;
        RECT 107.490 140.245 109.180 140.765 ;
        RECT 109.350 140.075 111.000 140.595 ;
        RECT 111.170 140.225 111.690 140.765 ;
        RECT 105.645 139.855 106.310 140.025 ;
        RECT 105.640 139.305 105.970 139.685 ;
        RECT 106.140 139.565 106.310 139.855 ;
        RECT 107.490 139.305 111.000 140.075 ;
        RECT 111.860 140.055 112.380 140.595 ;
        RECT 111.170 139.305 112.380 140.055 ;
        RECT 18.165 139.135 112.465 139.305 ;
        RECT 18.250 138.385 19.460 139.135 ;
        RECT 18.250 137.845 18.770 138.385 ;
        RECT 20.610 138.315 20.820 139.135 ;
        RECT 20.990 138.335 21.320 138.965 ;
        RECT 18.940 137.675 19.460 138.215 ;
        RECT 20.990 137.735 21.240 138.335 ;
        RECT 21.490 138.315 21.720 139.135 ;
        RECT 21.930 138.410 22.220 139.135 ;
        RECT 22.390 138.385 23.600 139.135 ;
        RECT 23.775 138.585 24.030 138.875 ;
        RECT 24.200 138.755 24.530 139.135 ;
        RECT 23.775 138.415 24.525 138.585 ;
        RECT 21.410 137.895 21.740 138.145 ;
        RECT 18.250 136.585 19.460 137.675 ;
        RECT 20.610 136.585 20.820 137.725 ;
        RECT 20.990 136.755 21.320 137.735 ;
        RECT 21.490 136.585 21.720 137.725 ;
        RECT 21.930 136.585 22.220 137.750 ;
        RECT 22.390 137.675 22.910 138.215 ;
        RECT 23.080 137.845 23.600 138.385 ;
        RECT 22.390 136.585 23.600 137.675 ;
        RECT 23.775 137.595 24.125 138.245 ;
        RECT 24.295 137.425 24.525 138.415 ;
        RECT 23.775 137.255 24.525 137.425 ;
        RECT 23.775 136.755 24.030 137.255 ;
        RECT 24.200 136.585 24.530 137.085 ;
        RECT 24.700 136.755 24.870 138.875 ;
        RECT 25.230 138.775 25.560 139.135 ;
        RECT 25.730 138.745 26.225 138.915 ;
        RECT 26.430 138.745 27.285 138.915 ;
        RECT 25.100 137.555 25.560 138.605 ;
        RECT 25.040 136.770 25.365 137.555 ;
        RECT 25.730 137.385 25.900 138.745 ;
        RECT 26.070 137.835 26.420 138.455 ;
        RECT 26.590 138.235 26.945 138.455 ;
        RECT 26.590 137.645 26.760 138.235 ;
        RECT 27.115 138.035 27.285 138.745 ;
        RECT 28.160 138.675 28.490 139.135 ;
        RECT 28.700 138.775 29.050 138.945 ;
        RECT 27.490 138.205 28.280 138.455 ;
        RECT 28.700 138.385 28.960 138.775 ;
        RECT 29.270 138.685 30.220 138.965 ;
        RECT 30.390 138.695 30.580 139.135 ;
        RECT 30.750 138.755 31.820 138.925 ;
        RECT 28.450 138.035 28.620 138.215 ;
        RECT 25.730 137.215 26.125 137.385 ;
        RECT 26.295 137.255 26.760 137.645 ;
        RECT 26.930 137.865 28.620 138.035 ;
        RECT 25.955 137.085 26.125 137.215 ;
        RECT 26.930 137.085 27.100 137.865 ;
        RECT 28.790 137.695 28.960 138.385 ;
        RECT 27.460 137.525 28.960 137.695 ;
        RECT 29.150 137.725 29.360 138.515 ;
        RECT 29.530 137.895 29.880 138.515 ;
        RECT 30.050 137.905 30.220 138.685 ;
        RECT 30.750 138.525 30.920 138.755 ;
        RECT 30.390 138.355 30.920 138.525 ;
        RECT 30.390 138.075 30.610 138.355 ;
        RECT 31.090 138.185 31.330 138.585 ;
        RECT 30.050 137.735 30.455 137.905 ;
        RECT 30.790 137.815 31.330 138.185 ;
        RECT 31.500 138.400 31.820 138.755 ;
        RECT 32.065 138.675 32.370 139.135 ;
        RECT 32.540 138.425 32.795 138.955 ;
        RECT 31.500 138.225 31.825 138.400 ;
        RECT 31.500 137.925 32.415 138.225 ;
        RECT 31.675 137.895 32.415 137.925 ;
        RECT 29.150 137.565 29.825 137.725 ;
        RECT 30.285 137.645 30.455 137.735 ;
        RECT 29.150 137.555 30.115 137.565 ;
        RECT 28.790 137.385 28.960 137.525 ;
        RECT 25.535 136.585 25.785 137.045 ;
        RECT 25.955 136.755 26.205 137.085 ;
        RECT 26.420 136.755 27.100 137.085 ;
        RECT 27.270 137.185 28.345 137.355 ;
        RECT 28.790 137.215 29.350 137.385 ;
        RECT 29.655 137.265 30.115 137.555 ;
        RECT 30.285 137.475 31.505 137.645 ;
        RECT 27.270 136.845 27.440 137.185 ;
        RECT 27.675 136.585 28.005 137.015 ;
        RECT 28.175 136.845 28.345 137.185 ;
        RECT 28.640 136.585 29.010 137.045 ;
        RECT 29.180 136.755 29.350 137.215 ;
        RECT 30.285 137.095 30.455 137.475 ;
        RECT 31.675 137.305 31.845 137.895 ;
        RECT 32.585 137.775 32.795 138.425 ;
        RECT 29.585 136.755 30.455 137.095 ;
        RECT 31.045 137.135 31.845 137.305 ;
        RECT 30.625 136.585 30.875 137.045 ;
        RECT 31.045 136.845 31.215 137.135 ;
        RECT 31.395 136.585 31.725 136.965 ;
        RECT 32.065 136.585 32.370 137.725 ;
        RECT 32.540 136.895 32.795 137.775 ;
        RECT 32.975 138.425 33.230 138.955 ;
        RECT 33.400 138.675 33.705 139.135 ;
        RECT 33.950 138.755 35.020 138.925 ;
        RECT 32.975 137.775 33.185 138.425 ;
        RECT 33.950 138.400 34.270 138.755 ;
        RECT 33.945 138.225 34.270 138.400 ;
        RECT 33.355 137.925 34.270 138.225 ;
        RECT 34.440 138.185 34.680 138.585 ;
        RECT 34.850 138.525 35.020 138.755 ;
        RECT 35.190 138.695 35.380 139.135 ;
        RECT 35.550 138.685 36.500 138.965 ;
        RECT 36.720 138.775 37.070 138.945 ;
        RECT 34.850 138.355 35.380 138.525 ;
        RECT 33.355 137.895 34.095 137.925 ;
        RECT 32.975 136.895 33.230 137.775 ;
        RECT 33.400 136.585 33.705 137.725 ;
        RECT 33.925 137.305 34.095 137.895 ;
        RECT 34.440 137.815 34.980 138.185 ;
        RECT 35.160 138.075 35.380 138.355 ;
        RECT 35.550 137.905 35.720 138.685 ;
        RECT 35.315 137.735 35.720 137.905 ;
        RECT 35.890 137.895 36.240 138.515 ;
        RECT 35.315 137.645 35.485 137.735 ;
        RECT 36.410 137.725 36.620 138.515 ;
        RECT 34.265 137.475 35.485 137.645 ;
        RECT 35.945 137.565 36.620 137.725 ;
        RECT 33.925 137.135 34.725 137.305 ;
        RECT 34.045 136.585 34.375 136.965 ;
        RECT 34.555 136.845 34.725 137.135 ;
        RECT 35.315 137.095 35.485 137.475 ;
        RECT 35.655 137.555 36.620 137.565 ;
        RECT 36.810 138.385 37.070 138.775 ;
        RECT 37.280 138.675 37.610 139.135 ;
        RECT 38.485 138.745 39.340 138.915 ;
        RECT 39.545 138.745 40.040 138.915 ;
        RECT 40.210 138.775 40.540 139.135 ;
        RECT 36.810 137.695 36.980 138.385 ;
        RECT 37.150 138.035 37.320 138.215 ;
        RECT 37.490 138.205 38.280 138.455 ;
        RECT 38.485 138.035 38.655 138.745 ;
        RECT 38.825 138.235 39.180 138.455 ;
        RECT 37.150 137.865 38.840 138.035 ;
        RECT 35.655 137.265 36.115 137.555 ;
        RECT 36.810 137.525 38.310 137.695 ;
        RECT 36.810 137.385 36.980 137.525 ;
        RECT 36.420 137.215 36.980 137.385 ;
        RECT 34.895 136.585 35.145 137.045 ;
        RECT 35.315 136.755 36.185 137.095 ;
        RECT 36.420 136.755 36.590 137.215 ;
        RECT 37.425 137.185 38.500 137.355 ;
        RECT 36.760 136.585 37.130 137.045 ;
        RECT 37.425 136.845 37.595 137.185 ;
        RECT 37.765 136.585 38.095 137.015 ;
        RECT 38.330 136.845 38.500 137.185 ;
        RECT 38.670 137.085 38.840 137.865 ;
        RECT 39.010 137.645 39.180 138.235 ;
        RECT 39.350 137.835 39.700 138.455 ;
        RECT 39.010 137.255 39.475 137.645 ;
        RECT 39.870 137.385 40.040 138.745 ;
        RECT 40.210 137.555 40.670 138.605 ;
        RECT 39.645 137.215 40.040 137.385 ;
        RECT 39.645 137.085 39.815 137.215 ;
        RECT 38.670 136.755 39.350 137.085 ;
        RECT 39.565 136.755 39.815 137.085 ;
        RECT 39.985 136.585 40.235 137.045 ;
        RECT 40.405 136.770 40.730 137.555 ;
        RECT 40.900 136.755 41.070 138.875 ;
        RECT 41.240 138.755 41.570 139.135 ;
        RECT 41.740 138.585 41.995 138.875 ;
        RECT 41.245 138.415 41.995 138.585 ;
        RECT 41.245 137.425 41.475 138.415 ;
        RECT 42.175 138.295 42.435 139.135 ;
        RECT 42.610 138.390 42.865 138.965 ;
        RECT 43.035 138.755 43.365 139.135 ;
        RECT 43.580 138.585 43.750 138.965 ;
        RECT 43.035 138.415 43.750 138.585 ;
        RECT 41.645 137.595 41.995 138.245 ;
        RECT 41.245 137.255 41.995 137.425 ;
        RECT 41.240 136.585 41.570 137.085 ;
        RECT 41.740 136.755 41.995 137.255 ;
        RECT 42.175 136.585 42.435 137.735 ;
        RECT 42.610 137.660 42.780 138.390 ;
        RECT 43.035 138.225 43.205 138.415 ;
        RECT 44.010 138.335 44.350 138.965 ;
        RECT 44.520 138.335 44.770 139.135 ;
        RECT 44.960 138.485 45.290 138.965 ;
        RECT 45.460 138.675 45.685 139.135 ;
        RECT 45.855 138.485 46.185 138.965 ;
        RECT 42.950 137.895 43.205 138.225 ;
        RECT 43.035 137.685 43.205 137.895 ;
        RECT 43.485 137.865 43.840 138.235 ;
        RECT 44.010 137.725 44.185 138.335 ;
        RECT 44.960 138.315 46.185 138.485 ;
        RECT 46.815 138.355 47.315 138.965 ;
        RECT 47.690 138.410 47.980 139.135 ;
        RECT 49.445 138.795 49.700 138.955 ;
        RECT 49.360 138.625 49.700 138.795 ;
        RECT 49.880 138.675 50.165 139.135 ;
        RECT 49.445 138.425 49.700 138.625 ;
        RECT 44.355 137.975 45.050 138.145 ;
        RECT 44.880 137.725 45.050 137.975 ;
        RECT 45.225 137.945 45.645 138.145 ;
        RECT 45.815 137.945 46.145 138.145 ;
        RECT 46.315 137.945 46.645 138.145 ;
        RECT 46.815 137.725 46.985 138.355 ;
        RECT 47.170 137.895 47.520 138.145 ;
        RECT 42.610 136.755 42.865 137.660 ;
        RECT 43.035 137.515 43.750 137.685 ;
        RECT 43.035 136.585 43.365 137.345 ;
        RECT 43.580 136.755 43.750 137.515 ;
        RECT 44.010 136.755 44.350 137.725 ;
        RECT 44.520 136.585 44.690 137.725 ;
        RECT 44.880 137.555 47.315 137.725 ;
        RECT 44.960 136.585 45.210 137.385 ;
        RECT 45.855 136.755 46.185 137.555 ;
        RECT 46.485 136.585 46.815 137.385 ;
        RECT 46.985 136.755 47.315 137.555 ;
        RECT 47.690 136.585 47.980 137.750 ;
        RECT 49.445 137.565 49.625 138.425 ;
        RECT 50.345 138.225 50.595 138.875 ;
        RECT 49.795 137.895 50.595 138.225 ;
        RECT 49.445 136.895 49.700 137.565 ;
        RECT 49.880 136.585 50.165 137.385 ;
        RECT 50.345 137.305 50.595 137.895 ;
        RECT 50.795 138.540 51.115 138.870 ;
        RECT 51.295 138.655 51.955 139.135 ;
        RECT 52.155 138.745 53.005 138.915 ;
        RECT 50.795 137.645 50.985 138.540 ;
        RECT 51.305 138.215 51.965 138.485 ;
        RECT 51.635 138.155 51.965 138.215 ;
        RECT 51.155 137.985 51.485 138.045 ;
        RECT 52.155 137.985 52.325 138.745 ;
        RECT 53.565 138.675 53.885 139.135 ;
        RECT 54.085 138.495 54.335 138.925 ;
        RECT 54.625 138.695 55.035 139.135 ;
        RECT 55.205 138.755 56.220 138.955 ;
        RECT 52.495 138.325 53.745 138.495 ;
        RECT 52.495 138.205 52.825 138.325 ;
        RECT 51.155 137.815 53.055 137.985 ;
        RECT 50.795 137.475 52.715 137.645 ;
        RECT 50.795 137.455 51.115 137.475 ;
        RECT 50.345 136.795 50.675 137.305 ;
        RECT 50.945 136.845 51.115 137.455 ;
        RECT 52.885 137.305 53.055 137.815 ;
        RECT 53.225 137.745 53.405 138.155 ;
        RECT 53.575 137.565 53.745 138.325 ;
        RECT 51.285 136.585 51.615 137.275 ;
        RECT 51.845 137.135 53.055 137.305 ;
        RECT 53.225 137.255 53.745 137.565 ;
        RECT 53.915 138.155 54.335 138.495 ;
        RECT 54.625 138.155 55.035 138.485 ;
        RECT 53.915 137.385 54.105 138.155 ;
        RECT 55.205 138.025 55.375 138.755 ;
        RECT 56.520 138.585 56.690 138.915 ;
        RECT 56.860 138.755 57.190 139.135 ;
        RECT 55.545 138.205 55.895 138.575 ;
        RECT 55.205 137.985 55.625 138.025 ;
        RECT 54.275 137.815 55.625 137.985 ;
        RECT 54.275 137.655 54.525 137.815 ;
        RECT 55.035 137.385 55.285 137.645 ;
        RECT 53.915 137.135 55.285 137.385 ;
        RECT 51.845 136.845 52.085 137.135 ;
        RECT 52.885 137.055 53.055 137.135 ;
        RECT 52.285 136.585 52.705 136.965 ;
        RECT 52.885 136.805 53.515 137.055 ;
        RECT 53.985 136.585 54.315 136.965 ;
        RECT 54.485 136.845 54.655 137.135 ;
        RECT 55.455 136.970 55.625 137.815 ;
        RECT 56.075 137.645 56.295 138.515 ;
        RECT 56.520 138.395 57.215 138.585 ;
        RECT 55.795 137.265 56.295 137.645 ;
        RECT 56.465 137.595 56.875 138.215 ;
        RECT 57.045 137.425 57.215 138.395 ;
        RECT 56.520 137.255 57.215 137.425 ;
        RECT 54.835 136.585 55.215 136.965 ;
        RECT 55.455 136.800 56.285 136.970 ;
        RECT 56.520 136.755 56.690 137.255 ;
        RECT 56.860 136.585 57.190 137.085 ;
        RECT 57.405 136.755 57.630 138.875 ;
        RECT 57.800 138.755 58.130 139.135 ;
        RECT 58.300 138.585 58.470 138.875 ;
        RECT 57.805 138.415 58.470 138.585 ;
        RECT 58.845 138.505 59.130 138.965 ;
        RECT 59.300 138.675 59.570 139.135 ;
        RECT 57.805 137.425 58.035 138.415 ;
        RECT 58.845 138.335 59.800 138.505 ;
        RECT 58.205 137.595 58.555 138.245 ;
        RECT 58.730 137.605 59.420 138.165 ;
        RECT 59.590 137.435 59.800 138.335 ;
        RECT 57.805 137.255 58.470 137.425 ;
        RECT 57.800 136.585 58.130 137.085 ;
        RECT 58.300 136.755 58.470 137.255 ;
        RECT 58.845 137.215 59.800 137.435 ;
        RECT 59.970 138.165 60.370 138.965 ;
        RECT 60.560 138.505 60.840 138.965 ;
        RECT 61.360 138.675 61.685 139.135 ;
        RECT 60.560 138.335 61.685 138.505 ;
        RECT 61.855 138.395 62.240 138.965 ;
        RECT 61.235 138.225 61.685 138.335 ;
        RECT 59.970 137.605 61.065 138.165 ;
        RECT 61.235 137.895 61.790 138.225 ;
        RECT 58.845 136.755 59.130 137.215 ;
        RECT 59.300 136.585 59.570 137.045 ;
        RECT 59.970 136.755 60.370 137.605 ;
        RECT 61.235 137.435 61.685 137.895 ;
        RECT 61.960 137.725 62.240 138.395 ;
        RECT 60.560 137.215 61.685 137.435 ;
        RECT 60.560 136.755 60.840 137.215 ;
        RECT 61.360 136.585 61.685 137.045 ;
        RECT 61.855 136.755 62.240 137.725 ;
        RECT 62.410 138.335 62.750 138.965 ;
        RECT 62.920 138.335 63.170 139.135 ;
        RECT 63.360 138.485 63.690 138.965 ;
        RECT 63.860 138.675 64.085 139.135 ;
        RECT 64.255 138.485 64.585 138.965 ;
        RECT 62.410 137.725 62.585 138.335 ;
        RECT 63.360 138.315 64.585 138.485 ;
        RECT 65.215 138.355 65.715 138.965 ;
        RECT 66.090 138.365 67.760 139.135 ;
        RECT 62.755 137.975 63.450 138.145 ;
        RECT 63.280 137.725 63.450 137.975 ;
        RECT 63.625 137.945 64.045 138.145 ;
        RECT 64.215 137.945 64.545 138.145 ;
        RECT 64.715 137.945 65.045 138.145 ;
        RECT 65.215 137.725 65.385 138.355 ;
        RECT 65.570 137.895 65.920 138.145 ;
        RECT 62.410 136.755 62.750 137.725 ;
        RECT 62.920 136.585 63.090 137.725 ;
        RECT 63.280 137.555 65.715 137.725 ;
        RECT 63.360 136.585 63.610 137.385 ;
        RECT 64.255 136.755 64.585 137.555 ;
        RECT 64.885 136.585 65.215 137.385 ;
        RECT 65.385 136.755 65.715 137.555 ;
        RECT 66.090 137.675 66.840 138.195 ;
        RECT 67.010 137.845 67.760 138.365 ;
        RECT 67.930 138.335 68.270 138.965 ;
        RECT 68.440 138.335 68.690 139.135 ;
        RECT 68.880 138.485 69.210 138.965 ;
        RECT 69.380 138.675 69.605 139.135 ;
        RECT 69.775 138.485 70.105 138.965 ;
        RECT 67.930 137.725 68.105 138.335 ;
        RECT 68.880 138.315 70.105 138.485 ;
        RECT 70.735 138.355 71.235 138.965 ;
        RECT 68.275 137.975 68.970 138.145 ;
        RECT 68.800 137.725 68.970 137.975 ;
        RECT 69.145 137.945 69.565 138.145 ;
        RECT 69.735 137.945 70.065 138.145 ;
        RECT 70.235 137.945 70.565 138.145 ;
        RECT 70.735 137.725 70.905 138.355 ;
        RECT 71.670 138.315 71.880 139.135 ;
        RECT 72.050 138.335 72.380 138.965 ;
        RECT 71.090 137.895 71.440 138.145 ;
        RECT 72.050 137.735 72.300 138.335 ;
        RECT 72.550 138.315 72.780 139.135 ;
        RECT 73.450 138.410 73.740 139.135 ;
        RECT 74.185 138.325 74.430 138.930 ;
        RECT 74.650 138.600 75.160 139.135 ;
        RECT 73.910 138.155 75.140 138.325 ;
        RECT 72.470 137.895 72.800 138.145 ;
        RECT 66.090 136.585 67.760 137.675 ;
        RECT 67.930 136.755 68.270 137.725 ;
        RECT 68.440 136.585 68.610 137.725 ;
        RECT 68.800 137.555 71.235 137.725 ;
        RECT 68.880 136.585 69.130 137.385 ;
        RECT 69.775 136.755 70.105 137.555 ;
        RECT 70.405 136.585 70.735 137.385 ;
        RECT 70.905 136.755 71.235 137.555 ;
        RECT 71.670 136.585 71.880 137.725 ;
        RECT 72.050 136.755 72.380 137.735 ;
        RECT 72.550 136.585 72.780 137.725 ;
        RECT 73.450 136.585 73.740 137.750 ;
        RECT 73.910 137.345 74.250 138.155 ;
        RECT 74.420 137.590 75.170 137.780 ;
        RECT 73.910 136.935 74.425 137.345 ;
        RECT 74.660 136.585 74.830 137.345 ;
        RECT 75.000 136.925 75.170 137.590 ;
        RECT 75.340 137.605 75.530 138.965 ;
        RECT 75.700 138.455 75.975 138.965 ;
        RECT 76.165 138.600 76.695 138.965 ;
        RECT 77.120 138.735 77.450 139.135 ;
        RECT 76.520 138.565 76.695 138.600 ;
        RECT 75.700 138.285 75.980 138.455 ;
        RECT 75.700 137.805 75.975 138.285 ;
        RECT 76.180 137.605 76.350 138.405 ;
        RECT 75.340 137.435 76.350 137.605 ;
        RECT 76.520 138.395 77.450 138.565 ;
        RECT 77.620 138.395 77.875 138.965 ;
        RECT 76.520 137.265 76.690 138.395 ;
        RECT 77.280 138.225 77.450 138.395 ;
        RECT 75.565 137.095 76.690 137.265 ;
        RECT 76.860 137.895 77.055 138.225 ;
        RECT 77.280 137.895 77.535 138.225 ;
        RECT 76.860 136.925 77.030 137.895 ;
        RECT 77.705 137.725 77.875 138.395 ;
        RECT 78.050 138.385 79.260 139.135 ;
        RECT 79.805 138.795 80.060 138.955 ;
        RECT 79.720 138.625 80.060 138.795 ;
        RECT 80.240 138.675 80.525 139.135 ;
        RECT 75.000 136.755 77.030 136.925 ;
        RECT 77.200 136.585 77.370 137.725 ;
        RECT 77.540 136.755 77.875 137.725 ;
        RECT 78.050 137.675 78.570 138.215 ;
        RECT 78.740 137.845 79.260 138.385 ;
        RECT 79.805 138.425 80.060 138.625 ;
        RECT 78.050 136.585 79.260 137.675 ;
        RECT 79.805 137.565 79.985 138.425 ;
        RECT 80.705 138.225 80.955 138.875 ;
        RECT 80.155 137.895 80.955 138.225 ;
        RECT 79.805 136.895 80.060 137.565 ;
        RECT 80.240 136.585 80.525 137.385 ;
        RECT 80.705 137.305 80.955 137.895 ;
        RECT 81.155 138.540 81.475 138.870 ;
        RECT 81.655 138.655 82.315 139.135 ;
        RECT 82.515 138.745 83.365 138.915 ;
        RECT 81.155 137.645 81.345 138.540 ;
        RECT 81.665 138.215 82.325 138.485 ;
        RECT 81.995 138.155 82.325 138.215 ;
        RECT 81.515 137.985 81.845 138.045 ;
        RECT 82.515 137.985 82.685 138.745 ;
        RECT 83.925 138.675 84.245 139.135 ;
        RECT 84.445 138.495 84.695 138.925 ;
        RECT 84.985 138.695 85.395 139.135 ;
        RECT 85.565 138.755 86.580 138.955 ;
        RECT 82.855 138.325 84.105 138.495 ;
        RECT 82.855 138.205 83.185 138.325 ;
        RECT 81.515 137.815 83.415 137.985 ;
        RECT 81.155 137.475 83.075 137.645 ;
        RECT 81.155 137.455 81.475 137.475 ;
        RECT 80.705 136.795 81.035 137.305 ;
        RECT 81.305 136.845 81.475 137.455 ;
        RECT 83.245 137.305 83.415 137.815 ;
        RECT 83.585 137.745 83.765 138.155 ;
        RECT 83.935 137.565 84.105 138.325 ;
        RECT 81.645 136.585 81.975 137.275 ;
        RECT 82.205 137.135 83.415 137.305 ;
        RECT 83.585 137.255 84.105 137.565 ;
        RECT 84.275 138.155 84.695 138.495 ;
        RECT 84.985 138.155 85.395 138.485 ;
        RECT 84.275 137.385 84.465 138.155 ;
        RECT 85.565 138.025 85.735 138.755 ;
        RECT 86.880 138.585 87.050 138.915 ;
        RECT 87.220 138.755 87.550 139.135 ;
        RECT 85.905 138.205 86.255 138.575 ;
        RECT 85.565 137.985 85.985 138.025 ;
        RECT 84.635 137.815 85.985 137.985 ;
        RECT 84.635 137.655 84.885 137.815 ;
        RECT 85.395 137.385 85.645 137.645 ;
        RECT 84.275 137.135 85.645 137.385 ;
        RECT 82.205 136.845 82.445 137.135 ;
        RECT 83.245 137.055 83.415 137.135 ;
        RECT 82.645 136.585 83.065 136.965 ;
        RECT 83.245 136.805 83.875 137.055 ;
        RECT 84.345 136.585 84.675 136.965 ;
        RECT 84.845 136.845 85.015 137.135 ;
        RECT 85.815 136.970 85.985 137.815 ;
        RECT 86.435 137.645 86.655 138.515 ;
        RECT 86.880 138.395 87.575 138.585 ;
        RECT 86.155 137.265 86.655 137.645 ;
        RECT 86.825 137.595 87.235 138.215 ;
        RECT 87.405 137.425 87.575 138.395 ;
        RECT 86.880 137.255 87.575 137.425 ;
        RECT 85.195 136.585 85.575 136.965 ;
        RECT 85.815 136.800 86.645 136.970 ;
        RECT 86.880 136.755 87.050 137.255 ;
        RECT 87.220 136.585 87.550 137.085 ;
        RECT 87.765 136.755 87.990 138.875 ;
        RECT 88.160 138.755 88.490 139.135 ;
        RECT 88.660 138.585 88.830 138.875 ;
        RECT 88.165 138.415 88.830 138.585 ;
        RECT 88.165 137.425 88.395 138.415 ;
        RECT 89.090 138.335 89.430 138.965 ;
        RECT 89.600 138.335 89.850 139.135 ;
        RECT 90.040 138.485 90.370 138.965 ;
        RECT 90.540 138.675 90.765 139.135 ;
        RECT 90.935 138.485 91.265 138.965 ;
        RECT 88.565 137.595 88.915 138.245 ;
        RECT 89.090 137.725 89.265 138.335 ;
        RECT 90.040 138.315 91.265 138.485 ;
        RECT 91.895 138.355 92.395 138.965 ;
        RECT 93.230 138.365 94.900 139.135 ;
        RECT 89.435 137.975 90.130 138.145 ;
        RECT 89.960 137.725 90.130 137.975 ;
        RECT 90.305 137.945 90.725 138.145 ;
        RECT 90.895 137.945 91.225 138.145 ;
        RECT 91.395 137.945 91.725 138.145 ;
        RECT 91.895 137.725 92.065 138.355 ;
        RECT 92.250 137.895 92.600 138.145 ;
        RECT 88.165 137.255 88.830 137.425 ;
        RECT 88.160 136.585 88.490 137.085 ;
        RECT 88.660 136.755 88.830 137.255 ;
        RECT 89.090 136.755 89.430 137.725 ;
        RECT 89.600 136.585 89.770 137.725 ;
        RECT 89.960 137.555 92.395 137.725 ;
        RECT 90.040 136.585 90.290 137.385 ;
        RECT 90.935 136.755 91.265 137.555 ;
        RECT 91.565 136.585 91.895 137.385 ;
        RECT 92.065 136.755 92.395 137.555 ;
        RECT 93.230 137.675 93.980 138.195 ;
        RECT 94.150 137.845 94.900 138.365 ;
        RECT 95.345 138.325 95.590 138.930 ;
        RECT 95.810 138.600 96.320 139.135 ;
        RECT 95.070 138.155 96.300 138.325 ;
        RECT 93.230 136.585 94.900 137.675 ;
        RECT 95.070 137.345 95.410 138.155 ;
        RECT 95.580 137.590 96.330 137.780 ;
        RECT 95.070 136.935 95.585 137.345 ;
        RECT 95.820 136.585 95.990 137.345 ;
        RECT 96.160 136.925 96.330 137.590 ;
        RECT 96.500 137.605 96.690 138.965 ;
        RECT 96.860 138.455 97.135 138.965 ;
        RECT 97.325 138.600 97.855 138.965 ;
        RECT 98.280 138.735 98.610 139.135 ;
        RECT 97.680 138.565 97.855 138.600 ;
        RECT 96.860 138.285 97.140 138.455 ;
        RECT 96.860 137.805 97.135 138.285 ;
        RECT 97.340 137.605 97.510 138.405 ;
        RECT 96.500 137.435 97.510 137.605 ;
        RECT 97.680 138.395 98.610 138.565 ;
        RECT 98.780 138.395 99.035 138.965 ;
        RECT 99.210 138.410 99.500 139.135 ;
        RECT 100.595 138.585 100.850 138.875 ;
        RECT 101.020 138.755 101.350 139.135 ;
        RECT 100.595 138.415 101.345 138.585 ;
        RECT 97.680 137.265 97.850 138.395 ;
        RECT 98.440 138.225 98.610 138.395 ;
        RECT 96.725 137.095 97.850 137.265 ;
        RECT 98.020 137.895 98.215 138.225 ;
        RECT 98.440 137.895 98.695 138.225 ;
        RECT 98.020 136.925 98.190 137.895 ;
        RECT 98.865 137.725 99.035 138.395 ;
        RECT 96.160 136.755 98.190 136.925 ;
        RECT 98.360 136.585 98.530 137.725 ;
        RECT 98.700 136.755 99.035 137.725 ;
        RECT 99.210 136.585 99.500 137.750 ;
        RECT 100.595 137.595 100.945 138.245 ;
        RECT 101.115 137.425 101.345 138.415 ;
        RECT 100.595 137.255 101.345 137.425 ;
        RECT 100.595 136.755 100.850 137.255 ;
        RECT 101.020 136.585 101.350 137.085 ;
        RECT 101.520 136.755 101.690 138.875 ;
        RECT 102.050 138.775 102.380 139.135 ;
        RECT 102.550 138.745 103.045 138.915 ;
        RECT 103.250 138.745 104.105 138.915 ;
        RECT 101.920 137.555 102.380 138.605 ;
        RECT 101.860 136.770 102.185 137.555 ;
        RECT 102.550 137.385 102.720 138.745 ;
        RECT 102.890 137.835 103.240 138.455 ;
        RECT 103.410 138.235 103.765 138.455 ;
        RECT 103.410 137.645 103.580 138.235 ;
        RECT 103.935 138.035 104.105 138.745 ;
        RECT 104.980 138.675 105.310 139.135 ;
        RECT 105.520 138.775 105.870 138.945 ;
        RECT 104.310 138.205 105.100 138.455 ;
        RECT 105.520 138.385 105.780 138.775 ;
        RECT 106.090 138.685 107.040 138.965 ;
        RECT 107.210 138.695 107.400 139.135 ;
        RECT 107.570 138.755 108.640 138.925 ;
        RECT 105.270 138.035 105.440 138.215 ;
        RECT 102.550 137.215 102.945 137.385 ;
        RECT 103.115 137.255 103.580 137.645 ;
        RECT 103.750 137.865 105.440 138.035 ;
        RECT 102.775 137.085 102.945 137.215 ;
        RECT 103.750 137.085 103.920 137.865 ;
        RECT 105.610 137.695 105.780 138.385 ;
        RECT 104.280 137.525 105.780 137.695 ;
        RECT 105.970 137.725 106.180 138.515 ;
        RECT 106.350 137.895 106.700 138.515 ;
        RECT 106.870 137.905 107.040 138.685 ;
        RECT 107.570 138.525 107.740 138.755 ;
        RECT 107.210 138.355 107.740 138.525 ;
        RECT 107.210 138.075 107.430 138.355 ;
        RECT 107.910 138.185 108.150 138.585 ;
        RECT 106.870 137.735 107.275 137.905 ;
        RECT 107.610 137.815 108.150 138.185 ;
        RECT 108.320 138.400 108.640 138.755 ;
        RECT 108.320 138.145 108.645 138.400 ;
        RECT 108.840 138.325 109.010 139.135 ;
        RECT 109.180 138.485 109.510 138.965 ;
        RECT 109.680 138.665 109.850 139.135 ;
        RECT 110.020 138.485 110.350 138.965 ;
        RECT 110.520 138.665 110.690 139.135 ;
        RECT 109.180 138.315 110.945 138.485 ;
        RECT 111.170 138.385 112.380 139.135 ;
        RECT 108.320 137.935 110.350 138.145 ;
        RECT 108.320 137.925 108.665 137.935 ;
        RECT 105.970 137.565 106.645 137.725 ;
        RECT 107.105 137.645 107.275 137.735 ;
        RECT 105.970 137.555 106.935 137.565 ;
        RECT 105.610 137.385 105.780 137.525 ;
        RECT 102.355 136.585 102.605 137.045 ;
        RECT 102.775 136.755 103.025 137.085 ;
        RECT 103.240 136.755 103.920 137.085 ;
        RECT 104.090 137.185 105.165 137.355 ;
        RECT 105.610 137.215 106.170 137.385 ;
        RECT 106.475 137.265 106.935 137.555 ;
        RECT 107.105 137.475 108.325 137.645 ;
        RECT 104.090 136.845 104.260 137.185 ;
        RECT 104.495 136.585 104.825 137.015 ;
        RECT 104.995 136.845 105.165 137.185 ;
        RECT 105.460 136.585 105.830 137.045 ;
        RECT 106.000 136.755 106.170 137.215 ;
        RECT 107.105 137.095 107.275 137.475 ;
        RECT 108.495 137.305 108.665 137.925 ;
        RECT 110.535 137.765 110.945 138.315 ;
        RECT 106.405 136.755 107.275 137.095 ;
        RECT 107.865 137.135 108.665 137.305 ;
        RECT 107.445 136.585 107.695 137.045 ;
        RECT 107.865 136.845 108.035 137.135 ;
        RECT 108.215 136.585 108.545 136.965 ;
        RECT 108.840 136.585 109.010 137.645 ;
        RECT 109.220 137.595 110.945 137.765 ;
        RECT 111.170 137.675 111.690 138.215 ;
        RECT 111.860 137.845 112.380 138.385 ;
        RECT 109.220 136.755 109.510 137.595 ;
        RECT 109.680 136.585 109.850 137.425 ;
        RECT 110.060 136.755 110.310 137.595 ;
        RECT 110.520 136.585 110.690 137.425 ;
        RECT 111.170 136.585 112.380 137.675 ;
        RECT 18.165 136.415 112.465 136.585 ;
        RECT 18.250 135.325 19.460 136.415 ;
        RECT 20.605 135.545 20.890 136.415 ;
        RECT 21.060 135.785 21.320 136.245 ;
        RECT 21.495 135.955 21.750 136.415 ;
        RECT 21.920 135.785 22.180 136.245 ;
        RECT 21.060 135.615 22.180 135.785 ;
        RECT 22.350 135.615 22.660 136.415 ;
        RECT 21.060 135.365 21.320 135.615 ;
        RECT 22.830 135.445 23.140 136.245 ;
        RECT 18.250 134.615 18.770 135.155 ;
        RECT 18.940 134.785 19.460 135.325 ;
        RECT 20.565 135.195 21.320 135.365 ;
        RECT 22.110 135.275 23.140 135.445 ;
        RECT 20.565 134.685 20.970 135.195 ;
        RECT 22.110 135.025 22.280 135.275 ;
        RECT 21.140 134.855 22.280 135.025 ;
        RECT 18.250 133.865 19.460 134.615 ;
        RECT 20.565 134.515 22.215 134.685 ;
        RECT 22.450 134.535 22.800 135.105 ;
        RECT 20.610 133.865 20.890 134.345 ;
        RECT 21.060 134.125 21.320 134.515 ;
        RECT 21.495 133.865 21.750 134.345 ;
        RECT 21.920 134.125 22.215 134.515 ;
        RECT 22.970 134.365 23.140 135.275 ;
        RECT 22.395 133.865 22.670 134.345 ;
        RECT 22.840 134.035 23.140 134.365 ;
        RECT 23.310 135.275 23.695 136.245 ;
        RECT 23.865 135.955 24.190 136.415 ;
        RECT 24.710 135.785 24.990 136.245 ;
        RECT 23.865 135.565 24.990 135.785 ;
        RECT 23.310 134.605 23.590 135.275 ;
        RECT 23.865 135.105 24.315 135.565 ;
        RECT 25.180 135.395 25.580 136.245 ;
        RECT 25.980 135.955 26.250 136.415 ;
        RECT 26.420 135.785 26.705 136.245 ;
        RECT 23.760 134.775 24.315 135.105 ;
        RECT 24.485 134.835 25.580 135.395 ;
        RECT 23.865 134.665 24.315 134.775 ;
        RECT 23.310 134.035 23.695 134.605 ;
        RECT 23.865 134.495 24.990 134.665 ;
        RECT 23.865 133.865 24.190 134.325 ;
        RECT 24.710 134.035 24.990 134.495 ;
        RECT 25.180 134.035 25.580 134.835 ;
        RECT 25.750 135.565 26.705 135.785 ;
        RECT 27.105 135.785 27.390 136.245 ;
        RECT 27.560 135.955 27.830 136.415 ;
        RECT 27.105 135.565 28.060 135.785 ;
        RECT 25.750 134.665 25.960 135.565 ;
        RECT 26.130 134.835 26.820 135.395 ;
        RECT 26.990 134.835 27.680 135.395 ;
        RECT 27.850 134.665 28.060 135.565 ;
        RECT 25.750 134.495 26.705 134.665 ;
        RECT 25.980 133.865 26.250 134.325 ;
        RECT 26.420 134.035 26.705 134.495 ;
        RECT 27.105 134.495 28.060 134.665 ;
        RECT 28.230 135.395 28.630 136.245 ;
        RECT 28.820 135.785 29.100 136.245 ;
        RECT 29.620 135.955 29.945 136.415 ;
        RECT 28.820 135.565 29.945 135.785 ;
        RECT 28.230 134.835 29.325 135.395 ;
        RECT 29.495 135.105 29.945 135.565 ;
        RECT 30.115 135.275 30.500 136.245 ;
        RECT 27.105 134.035 27.390 134.495 ;
        RECT 27.560 133.865 27.830 134.325 ;
        RECT 28.230 134.035 28.630 134.835 ;
        RECT 29.495 134.775 30.050 135.105 ;
        RECT 29.495 134.665 29.945 134.775 ;
        RECT 28.820 134.495 29.945 134.665 ;
        RECT 30.220 134.605 30.500 135.275 ;
        RECT 28.820 134.035 29.100 134.495 ;
        RECT 29.620 133.865 29.945 134.325 ;
        RECT 30.115 134.035 30.500 134.605 ;
        RECT 30.675 135.275 31.010 136.245 ;
        RECT 31.180 135.275 31.350 136.415 ;
        RECT 31.520 136.075 33.550 136.245 ;
        RECT 30.675 134.605 30.845 135.275 ;
        RECT 31.520 135.105 31.690 136.075 ;
        RECT 31.015 134.775 31.270 135.105 ;
        RECT 31.495 134.775 31.690 135.105 ;
        RECT 31.860 135.735 32.985 135.905 ;
        RECT 31.100 134.605 31.270 134.775 ;
        RECT 31.860 134.605 32.030 135.735 ;
        RECT 30.675 134.035 30.930 134.605 ;
        RECT 31.100 134.435 32.030 134.605 ;
        RECT 32.200 135.395 33.210 135.565 ;
        RECT 32.200 134.595 32.370 135.395 ;
        RECT 32.575 134.715 32.850 135.195 ;
        RECT 32.570 134.545 32.850 134.715 ;
        RECT 31.855 134.400 32.030 134.435 ;
        RECT 31.100 133.865 31.430 134.265 ;
        RECT 31.855 134.035 32.385 134.400 ;
        RECT 32.575 134.035 32.850 134.545 ;
        RECT 33.020 134.035 33.210 135.395 ;
        RECT 33.380 135.410 33.550 136.075 ;
        RECT 33.720 135.655 33.890 136.415 ;
        RECT 34.125 135.655 34.640 136.065 ;
        RECT 33.380 135.220 34.130 135.410 ;
        RECT 34.300 134.845 34.640 135.655 ;
        RECT 34.810 135.250 35.100 136.415 ;
        RECT 35.735 135.265 35.995 136.415 ;
        RECT 36.170 135.340 36.425 136.245 ;
        RECT 36.595 135.655 36.925 136.415 ;
        RECT 37.140 135.485 37.310 136.245 ;
        RECT 33.410 134.675 34.640 134.845 ;
        RECT 33.390 133.865 33.900 134.400 ;
        RECT 34.120 134.070 34.365 134.675 ;
        RECT 34.810 133.865 35.100 134.590 ;
        RECT 35.735 133.865 35.995 134.705 ;
        RECT 36.170 134.610 36.340 135.340 ;
        RECT 36.595 135.315 37.310 135.485 ;
        RECT 37.570 135.655 38.085 136.065 ;
        RECT 38.320 135.655 38.490 136.415 ;
        RECT 38.660 136.075 40.690 136.245 ;
        RECT 36.595 135.105 36.765 135.315 ;
        RECT 36.510 134.775 36.765 135.105 ;
        RECT 36.170 134.035 36.425 134.610 ;
        RECT 36.595 134.585 36.765 134.775 ;
        RECT 37.045 134.765 37.400 135.135 ;
        RECT 37.570 134.845 37.910 135.655 ;
        RECT 38.660 135.410 38.830 136.075 ;
        RECT 39.225 135.735 40.350 135.905 ;
        RECT 38.080 135.220 38.830 135.410 ;
        RECT 39.000 135.395 40.010 135.565 ;
        RECT 37.570 134.675 38.800 134.845 ;
        RECT 36.595 134.415 37.310 134.585 ;
        RECT 36.595 133.865 36.925 134.245 ;
        RECT 37.140 134.035 37.310 134.415 ;
        RECT 37.845 134.070 38.090 134.675 ;
        RECT 38.310 133.865 38.820 134.400 ;
        RECT 39.000 134.035 39.190 135.395 ;
        RECT 39.360 134.375 39.635 135.195 ;
        RECT 39.840 134.595 40.010 135.395 ;
        RECT 40.180 134.605 40.350 135.735 ;
        RECT 40.520 135.105 40.690 136.075 ;
        RECT 40.860 135.275 41.030 136.415 ;
        RECT 41.200 135.275 41.535 136.245 ;
        RECT 40.520 134.775 40.715 135.105 ;
        RECT 40.940 134.775 41.195 135.105 ;
        RECT 40.940 134.605 41.110 134.775 ;
        RECT 41.365 134.605 41.535 135.275 ;
        RECT 40.180 134.435 41.110 134.605 ;
        RECT 40.180 134.400 40.355 134.435 ;
        RECT 39.360 134.205 39.640 134.375 ;
        RECT 39.360 134.035 39.635 134.205 ;
        RECT 39.825 134.035 40.355 134.400 ;
        RECT 40.780 133.865 41.110 134.265 ;
        RECT 41.280 134.035 41.535 134.605 ;
        RECT 42.170 135.275 42.510 136.245 ;
        RECT 42.680 135.275 42.850 136.415 ;
        RECT 43.120 135.615 43.370 136.415 ;
        RECT 44.015 135.445 44.345 136.245 ;
        RECT 44.645 135.615 44.975 136.415 ;
        RECT 45.145 135.445 45.475 136.245 ;
        RECT 46.315 135.980 51.660 136.415 ;
        RECT 43.040 135.275 45.475 135.445 ;
        RECT 42.170 134.665 42.345 135.275 ;
        RECT 43.040 135.025 43.210 135.275 ;
        RECT 42.515 134.855 43.210 135.025 ;
        RECT 43.385 134.855 43.805 135.055 ;
        RECT 43.975 134.855 44.305 135.055 ;
        RECT 44.475 134.855 44.805 135.055 ;
        RECT 42.170 134.035 42.510 134.665 ;
        RECT 42.680 133.865 42.930 134.665 ;
        RECT 43.120 134.515 44.345 134.685 ;
        RECT 43.120 134.035 43.450 134.515 ;
        RECT 43.620 133.865 43.845 134.325 ;
        RECT 44.015 134.035 44.345 134.515 ;
        RECT 44.975 134.645 45.145 135.275 ;
        RECT 45.330 134.855 45.680 135.105 ;
        RECT 47.905 134.730 48.255 135.980 ;
        RECT 51.830 135.655 52.345 136.065 ;
        RECT 52.580 135.655 52.750 136.415 ;
        RECT 52.920 136.075 54.950 136.245 ;
        RECT 44.975 134.035 45.475 134.645 ;
        RECT 49.735 134.410 50.075 135.240 ;
        RECT 51.830 134.845 52.170 135.655 ;
        RECT 52.920 135.410 53.090 136.075 ;
        RECT 53.485 135.735 54.610 135.905 ;
        RECT 52.340 135.220 53.090 135.410 ;
        RECT 53.260 135.395 54.270 135.565 ;
        RECT 51.830 134.675 53.060 134.845 ;
        RECT 46.315 133.865 51.660 134.410 ;
        RECT 52.105 134.070 52.350 134.675 ;
        RECT 52.570 133.865 53.080 134.400 ;
        RECT 53.260 134.035 53.450 135.395 ;
        RECT 53.620 135.055 53.895 135.195 ;
        RECT 53.620 134.885 53.900 135.055 ;
        RECT 53.620 134.035 53.895 134.885 ;
        RECT 54.100 134.595 54.270 135.395 ;
        RECT 54.440 134.605 54.610 135.735 ;
        RECT 54.780 135.105 54.950 136.075 ;
        RECT 55.120 135.275 55.290 136.415 ;
        RECT 55.460 135.275 55.795 136.245 ;
        RECT 56.470 135.275 56.700 136.415 ;
        RECT 54.780 134.775 54.975 135.105 ;
        RECT 55.200 134.775 55.455 135.105 ;
        RECT 55.200 134.605 55.370 134.775 ;
        RECT 55.625 134.605 55.795 135.275 ;
        RECT 56.870 135.265 57.200 136.245 ;
        RECT 57.370 135.275 57.580 136.415 ;
        RECT 57.960 135.265 58.290 136.415 ;
        RECT 58.460 135.395 58.630 136.245 ;
        RECT 58.800 135.615 59.130 136.415 ;
        RECT 59.300 135.395 59.470 136.245 ;
        RECT 59.650 135.615 59.890 136.415 ;
        RECT 60.060 135.435 60.390 136.245 ;
        RECT 56.450 134.855 56.780 135.105 ;
        RECT 54.440 134.435 55.370 134.605 ;
        RECT 54.440 134.400 54.615 134.435 ;
        RECT 54.085 134.035 54.615 134.400 ;
        RECT 55.040 133.865 55.370 134.265 ;
        RECT 55.540 134.035 55.795 134.605 ;
        RECT 56.470 133.865 56.700 134.685 ;
        RECT 56.950 134.665 57.200 135.265 ;
        RECT 58.460 135.225 59.470 135.395 ;
        RECT 59.675 135.265 60.390 135.435 ;
        RECT 58.460 134.685 58.955 135.225 ;
        RECT 59.675 135.025 59.845 135.265 ;
        RECT 60.570 135.250 60.860 136.415 ;
        RECT 61.180 135.265 61.510 136.415 ;
        RECT 61.680 135.395 61.850 136.245 ;
        RECT 62.020 135.615 62.350 136.415 ;
        RECT 62.520 135.395 62.690 136.245 ;
        RECT 62.870 135.615 63.110 136.415 ;
        RECT 63.280 135.435 63.610 136.245 ;
        RECT 61.680 135.225 62.690 135.395 ;
        RECT 62.895 135.265 63.610 135.435 ;
        RECT 63.790 135.655 64.305 136.065 ;
        RECT 64.540 135.655 64.710 136.415 ;
        RECT 64.880 136.075 66.910 136.245 ;
        RECT 59.345 134.855 59.845 135.025 ;
        RECT 60.015 134.855 60.395 135.095 ;
        RECT 59.675 134.685 59.845 134.855 ;
        RECT 61.680 134.715 62.175 135.225 ;
        RECT 62.895 135.025 63.065 135.265 ;
        RECT 62.565 134.855 63.065 135.025 ;
        RECT 63.235 134.855 63.615 135.095 ;
        RECT 61.680 134.685 62.180 134.715 ;
        RECT 62.895 134.685 63.065 134.855 ;
        RECT 63.790 134.845 64.130 135.655 ;
        RECT 64.880 135.410 65.050 136.075 ;
        RECT 65.445 135.735 66.570 135.905 ;
        RECT 64.300 135.220 65.050 135.410 ;
        RECT 65.220 135.395 66.230 135.565 ;
        RECT 56.870 134.035 57.200 134.665 ;
        RECT 57.370 133.865 57.580 134.685 ;
        RECT 57.960 133.865 58.290 134.665 ;
        RECT 58.460 134.515 59.470 134.685 ;
        RECT 59.675 134.515 60.310 134.685 ;
        RECT 58.460 134.035 58.630 134.515 ;
        RECT 58.800 133.865 59.130 134.345 ;
        RECT 59.300 134.035 59.470 134.515 ;
        RECT 59.720 133.865 59.960 134.345 ;
        RECT 60.140 134.035 60.310 134.515 ;
        RECT 60.570 133.865 60.860 134.590 ;
        RECT 61.180 133.865 61.510 134.665 ;
        RECT 61.680 134.515 62.690 134.685 ;
        RECT 62.895 134.515 63.530 134.685 ;
        RECT 63.790 134.675 65.020 134.845 ;
        RECT 61.680 134.035 61.850 134.515 ;
        RECT 62.020 133.865 62.350 134.345 ;
        RECT 62.520 134.035 62.690 134.515 ;
        RECT 62.940 133.865 63.180 134.345 ;
        RECT 63.360 134.035 63.530 134.515 ;
        RECT 64.065 134.070 64.310 134.675 ;
        RECT 64.530 133.865 65.040 134.400 ;
        RECT 65.220 134.035 65.410 135.395 ;
        RECT 65.580 134.715 65.855 135.195 ;
        RECT 65.580 134.545 65.860 134.715 ;
        RECT 66.060 134.595 66.230 135.395 ;
        RECT 66.400 134.605 66.570 135.735 ;
        RECT 66.740 135.105 66.910 136.075 ;
        RECT 67.080 135.275 67.250 136.415 ;
        RECT 67.420 135.275 67.755 136.245 ;
        RECT 66.740 134.775 66.935 135.105 ;
        RECT 67.160 134.775 67.415 135.105 ;
        RECT 67.160 134.605 67.330 134.775 ;
        RECT 67.585 134.605 67.755 135.275 ;
        RECT 65.580 134.035 65.855 134.545 ;
        RECT 66.400 134.435 67.330 134.605 ;
        RECT 66.400 134.400 66.575 134.435 ;
        RECT 66.045 134.035 66.575 134.400 ;
        RECT 67.000 133.865 67.330 134.265 ;
        RECT 67.500 134.035 67.755 134.605 ;
        RECT 67.930 135.445 68.240 136.245 ;
        RECT 68.410 135.615 68.720 136.415 ;
        RECT 68.890 135.785 69.150 136.245 ;
        RECT 69.320 135.955 69.575 136.415 ;
        RECT 69.750 135.785 70.010 136.245 ;
        RECT 68.890 135.615 70.010 135.785 ;
        RECT 67.930 135.275 68.960 135.445 ;
        RECT 67.930 134.365 68.100 135.275 ;
        RECT 68.270 134.535 68.620 135.105 ;
        RECT 68.790 135.025 68.960 135.275 ;
        RECT 69.750 135.365 70.010 135.615 ;
        RECT 70.180 135.545 70.465 136.415 ;
        RECT 70.745 135.545 71.030 136.415 ;
        RECT 71.200 135.785 71.460 136.245 ;
        RECT 71.635 135.955 71.890 136.415 ;
        RECT 72.060 135.785 72.320 136.245 ;
        RECT 71.200 135.615 72.320 135.785 ;
        RECT 72.490 135.615 72.800 136.415 ;
        RECT 71.200 135.365 71.460 135.615 ;
        RECT 72.970 135.445 73.280 136.245 ;
        RECT 69.750 135.195 70.505 135.365 ;
        RECT 68.790 134.855 69.930 135.025 ;
        RECT 70.100 134.685 70.505 135.195 ;
        RECT 68.855 134.515 70.505 134.685 ;
        RECT 70.705 135.195 71.460 135.365 ;
        RECT 72.250 135.275 73.280 135.445 ;
        RECT 73.655 135.445 73.985 136.245 ;
        RECT 74.155 135.615 74.485 136.415 ;
        RECT 74.785 135.445 75.115 136.245 ;
        RECT 75.760 135.615 76.010 136.415 ;
        RECT 73.655 135.275 76.090 135.445 ;
        RECT 76.280 135.275 76.450 136.415 ;
        RECT 76.620 135.275 76.960 136.245 ;
        RECT 70.705 134.685 71.110 135.195 ;
        RECT 72.250 135.025 72.420 135.275 ;
        RECT 71.280 134.855 72.420 135.025 ;
        RECT 70.705 134.515 72.355 134.685 ;
        RECT 72.590 134.535 72.940 135.105 ;
        RECT 67.930 134.035 68.230 134.365 ;
        RECT 68.400 133.865 68.675 134.345 ;
        RECT 68.855 134.125 69.150 134.515 ;
        RECT 69.320 133.865 69.575 134.345 ;
        RECT 69.750 134.125 70.010 134.515 ;
        RECT 70.180 133.865 70.460 134.345 ;
        RECT 70.750 133.865 71.030 134.345 ;
        RECT 71.200 134.125 71.460 134.515 ;
        RECT 71.635 133.865 71.890 134.345 ;
        RECT 72.060 134.125 72.355 134.515 ;
        RECT 73.110 134.365 73.280 135.275 ;
        RECT 73.450 134.855 73.800 135.105 ;
        RECT 73.985 134.645 74.155 135.275 ;
        RECT 74.325 134.855 74.655 135.055 ;
        RECT 74.825 134.855 75.155 135.055 ;
        RECT 75.325 134.855 75.745 135.055 ;
        RECT 75.920 135.025 76.090 135.275 ;
        RECT 75.920 134.855 76.615 135.025 ;
        RECT 72.535 133.865 72.810 134.345 ;
        RECT 72.980 134.035 73.280 134.365 ;
        RECT 73.655 134.035 74.155 134.645 ;
        RECT 74.785 134.515 76.010 134.685 ;
        RECT 76.785 134.665 76.960 135.275 ;
        RECT 77.130 135.655 77.645 136.065 ;
        RECT 77.880 135.655 78.050 136.415 ;
        RECT 78.220 136.075 80.250 136.245 ;
        RECT 77.130 134.845 77.470 135.655 ;
        RECT 78.220 135.410 78.390 136.075 ;
        RECT 78.785 135.735 79.910 135.905 ;
        RECT 77.640 135.220 78.390 135.410 ;
        RECT 78.560 135.395 79.570 135.565 ;
        RECT 77.130 134.675 78.360 134.845 ;
        RECT 74.785 134.035 75.115 134.515 ;
        RECT 75.285 133.865 75.510 134.325 ;
        RECT 75.680 134.035 76.010 134.515 ;
        RECT 76.200 133.865 76.450 134.665 ;
        RECT 76.620 134.035 76.960 134.665 ;
        RECT 77.405 134.070 77.650 134.675 ;
        RECT 77.870 133.865 78.380 134.400 ;
        RECT 78.560 134.035 78.750 135.395 ;
        RECT 78.920 135.055 79.195 135.195 ;
        RECT 78.920 134.885 79.200 135.055 ;
        RECT 78.920 134.035 79.195 134.885 ;
        RECT 79.400 134.595 79.570 135.395 ;
        RECT 79.740 134.605 79.910 135.735 ;
        RECT 80.080 135.105 80.250 136.075 ;
        RECT 80.420 135.275 80.590 136.415 ;
        RECT 80.760 135.275 81.095 136.245 ;
        RECT 80.080 134.775 80.275 135.105 ;
        RECT 80.500 134.775 80.755 135.105 ;
        RECT 80.500 134.605 80.670 134.775 ;
        RECT 80.925 134.605 81.095 135.275 ;
        RECT 82.190 135.655 82.705 136.065 ;
        RECT 82.940 135.655 83.110 136.415 ;
        RECT 83.280 136.075 85.310 136.245 ;
        RECT 82.190 134.845 82.530 135.655 ;
        RECT 83.280 135.410 83.450 136.075 ;
        RECT 83.845 135.735 84.970 135.905 ;
        RECT 82.700 135.220 83.450 135.410 ;
        RECT 83.620 135.395 84.630 135.565 ;
        RECT 82.190 134.675 83.420 134.845 ;
        RECT 79.740 134.435 80.670 134.605 ;
        RECT 79.740 134.400 79.915 134.435 ;
        RECT 79.385 134.035 79.915 134.400 ;
        RECT 80.340 133.865 80.670 134.265 ;
        RECT 80.840 134.035 81.095 134.605 ;
        RECT 82.465 134.070 82.710 134.675 ;
        RECT 82.930 133.865 83.440 134.400 ;
        RECT 83.620 134.035 83.810 135.395 ;
        RECT 83.980 134.375 84.255 135.195 ;
        RECT 84.460 134.595 84.630 135.395 ;
        RECT 84.800 134.605 84.970 135.735 ;
        RECT 85.140 135.105 85.310 136.075 ;
        RECT 85.480 135.275 85.650 136.415 ;
        RECT 85.820 135.275 86.155 136.245 ;
        RECT 85.140 134.775 85.335 135.105 ;
        RECT 85.560 134.775 85.815 135.105 ;
        RECT 85.560 134.605 85.730 134.775 ;
        RECT 85.985 134.605 86.155 135.275 ;
        RECT 86.330 135.250 86.620 136.415 ;
        RECT 86.790 135.445 87.100 136.245 ;
        RECT 87.270 135.615 87.580 136.415 ;
        RECT 87.750 135.785 88.010 136.245 ;
        RECT 88.180 135.955 88.435 136.415 ;
        RECT 88.610 135.785 88.870 136.245 ;
        RECT 87.750 135.615 88.870 135.785 ;
        RECT 86.790 135.275 87.820 135.445 ;
        RECT 84.800 134.435 85.730 134.605 ;
        RECT 84.800 134.400 84.975 134.435 ;
        RECT 83.980 134.205 84.260 134.375 ;
        RECT 83.980 134.035 84.255 134.205 ;
        RECT 84.445 134.035 84.975 134.400 ;
        RECT 85.400 133.865 85.730 134.265 ;
        RECT 85.900 134.035 86.155 134.605 ;
        RECT 86.330 133.865 86.620 134.590 ;
        RECT 86.790 134.365 86.960 135.275 ;
        RECT 87.130 134.535 87.480 135.105 ;
        RECT 87.650 135.025 87.820 135.275 ;
        RECT 88.610 135.365 88.870 135.615 ;
        RECT 89.040 135.545 89.325 136.415 ;
        RECT 88.610 135.195 89.365 135.365 ;
        RECT 87.650 134.855 88.790 135.025 ;
        RECT 88.960 134.685 89.365 135.195 ;
        RECT 87.715 134.515 89.365 134.685 ;
        RECT 89.550 135.275 89.890 136.245 ;
        RECT 90.060 135.275 90.230 136.415 ;
        RECT 90.500 135.615 90.750 136.415 ;
        RECT 91.395 135.445 91.725 136.245 ;
        RECT 92.025 135.615 92.355 136.415 ;
        RECT 92.525 135.445 92.855 136.245 ;
        RECT 90.420 135.275 92.855 135.445 ;
        RECT 93.435 135.445 93.765 136.245 ;
        RECT 93.935 135.615 94.265 136.415 ;
        RECT 94.565 135.445 94.895 136.245 ;
        RECT 95.540 135.615 95.790 136.415 ;
        RECT 93.435 135.275 95.870 135.445 ;
        RECT 96.060 135.275 96.230 136.415 ;
        RECT 96.400 135.275 96.740 136.245 ;
        RECT 89.550 134.665 89.725 135.275 ;
        RECT 90.420 135.025 90.590 135.275 ;
        RECT 89.895 134.855 90.590 135.025 ;
        RECT 90.765 134.855 91.185 135.055 ;
        RECT 91.355 134.855 91.685 135.055 ;
        RECT 91.855 134.855 92.185 135.055 ;
        RECT 86.790 134.035 87.090 134.365 ;
        RECT 87.260 133.865 87.535 134.345 ;
        RECT 87.715 134.125 88.010 134.515 ;
        RECT 88.180 133.865 88.435 134.345 ;
        RECT 88.610 134.125 88.870 134.515 ;
        RECT 89.040 133.865 89.320 134.345 ;
        RECT 89.550 134.035 89.890 134.665 ;
        RECT 90.060 133.865 90.310 134.665 ;
        RECT 90.500 134.515 91.725 134.685 ;
        RECT 90.500 134.035 90.830 134.515 ;
        RECT 91.000 133.865 91.225 134.325 ;
        RECT 91.395 134.035 91.725 134.515 ;
        RECT 92.355 134.645 92.525 135.275 ;
        RECT 92.710 134.855 93.060 135.105 ;
        RECT 93.230 134.855 93.580 135.105 ;
        RECT 93.765 134.645 93.935 135.275 ;
        RECT 94.105 134.855 94.435 135.055 ;
        RECT 94.605 134.855 94.935 135.055 ;
        RECT 95.105 134.855 95.525 135.055 ;
        RECT 95.700 135.025 95.870 135.275 ;
        RECT 95.700 134.855 96.395 135.025 ;
        RECT 92.355 134.035 92.855 134.645 ;
        RECT 93.435 134.035 93.935 134.645 ;
        RECT 94.565 134.515 95.790 134.685 ;
        RECT 96.565 134.665 96.740 135.275 ;
        RECT 96.910 135.325 99.500 136.415 ;
        RECT 96.910 134.805 98.120 135.325 ;
        RECT 99.710 135.275 99.940 136.415 ;
        RECT 100.110 135.265 100.440 136.245 ;
        RECT 100.610 135.275 100.820 136.415 ;
        RECT 101.050 135.445 101.360 136.245 ;
        RECT 101.530 135.615 101.840 136.415 ;
        RECT 102.010 135.785 102.270 136.245 ;
        RECT 102.440 135.955 102.695 136.415 ;
        RECT 102.870 135.785 103.130 136.245 ;
        RECT 102.010 135.615 103.130 135.785 ;
        RECT 101.050 135.275 102.080 135.445 ;
        RECT 94.565 134.035 94.895 134.515 ;
        RECT 95.065 133.865 95.290 134.325 ;
        RECT 95.460 134.035 95.790 134.515 ;
        RECT 95.980 133.865 96.230 134.665 ;
        RECT 96.400 134.035 96.740 134.665 ;
        RECT 98.290 134.635 99.500 135.155 ;
        RECT 99.690 134.855 100.020 135.105 ;
        RECT 96.910 133.865 99.500 134.635 ;
        RECT 99.710 133.865 99.940 134.685 ;
        RECT 100.190 134.665 100.440 135.265 ;
        RECT 100.110 134.035 100.440 134.665 ;
        RECT 100.610 133.865 100.820 134.685 ;
        RECT 101.050 134.365 101.220 135.275 ;
        RECT 101.390 134.535 101.740 135.105 ;
        RECT 101.910 135.025 102.080 135.275 ;
        RECT 102.870 135.365 103.130 135.615 ;
        RECT 103.300 135.545 103.585 136.415 ;
        RECT 102.870 135.195 103.625 135.365 ;
        RECT 101.910 134.855 103.050 135.025 ;
        RECT 103.220 134.685 103.625 135.195 ;
        RECT 104.270 135.325 105.940 136.415 ;
        RECT 104.270 134.805 105.020 135.325 ;
        RECT 106.170 135.275 106.380 136.415 ;
        RECT 106.550 135.265 106.880 136.245 ;
        RECT 107.050 135.275 107.280 136.415 ;
        RECT 107.490 135.325 111.000 136.415 ;
        RECT 111.170 135.325 112.380 136.415 ;
        RECT 101.975 134.515 103.625 134.685 ;
        RECT 105.190 134.635 105.940 135.155 ;
        RECT 101.050 134.035 101.350 134.365 ;
        RECT 101.520 133.865 101.795 134.345 ;
        RECT 101.975 134.125 102.270 134.515 ;
        RECT 102.440 133.865 102.695 134.345 ;
        RECT 102.870 134.125 103.130 134.515 ;
        RECT 103.300 133.865 103.580 134.345 ;
        RECT 104.270 133.865 105.940 134.635 ;
        RECT 106.170 133.865 106.380 134.685 ;
        RECT 106.550 134.665 106.800 135.265 ;
        RECT 106.970 134.855 107.300 135.105 ;
        RECT 107.490 134.805 109.180 135.325 ;
        RECT 106.550 134.035 106.880 134.665 ;
        RECT 107.050 133.865 107.280 134.685 ;
        RECT 109.350 134.635 111.000 135.155 ;
        RECT 111.170 134.785 111.690 135.325 ;
        RECT 107.490 133.865 111.000 134.635 ;
        RECT 111.860 134.615 112.380 135.155 ;
        RECT 111.170 133.865 112.380 134.615 ;
        RECT 18.165 133.695 112.465 133.865 ;
        RECT 18.250 132.945 19.460 133.695 ;
        RECT 18.250 132.405 18.770 132.945 ;
        RECT 20.610 132.875 20.820 133.695 ;
        RECT 20.990 132.895 21.320 133.525 ;
        RECT 18.940 132.235 19.460 132.775 ;
        RECT 20.990 132.295 21.240 132.895 ;
        RECT 21.490 132.875 21.720 133.695 ;
        RECT 21.930 132.970 22.220 133.695 ;
        RECT 22.505 133.065 22.790 133.525 ;
        RECT 22.960 133.235 23.230 133.695 ;
        RECT 22.505 132.895 23.460 133.065 ;
        RECT 21.410 132.455 21.740 132.705 ;
        RECT 18.250 131.145 19.460 132.235 ;
        RECT 20.610 131.145 20.820 132.285 ;
        RECT 20.990 131.315 21.320 132.295 ;
        RECT 21.490 131.145 21.720 132.285 ;
        RECT 21.930 131.145 22.220 132.310 ;
        RECT 22.390 132.165 23.080 132.725 ;
        RECT 23.250 131.995 23.460 132.895 ;
        RECT 22.505 131.775 23.460 131.995 ;
        RECT 23.630 132.725 24.030 133.525 ;
        RECT 24.220 133.065 24.500 133.525 ;
        RECT 25.020 133.235 25.345 133.695 ;
        RECT 24.220 132.895 25.345 133.065 ;
        RECT 25.515 132.955 25.900 133.525 ;
        RECT 24.895 132.785 25.345 132.895 ;
        RECT 23.630 132.165 24.725 132.725 ;
        RECT 24.895 132.455 25.450 132.785 ;
        RECT 22.505 131.315 22.790 131.775 ;
        RECT 22.960 131.145 23.230 131.605 ;
        RECT 23.630 131.315 24.030 132.165 ;
        RECT 24.895 131.995 25.345 132.455 ;
        RECT 25.620 132.285 25.900 132.955 ;
        RECT 24.220 131.775 25.345 131.995 ;
        RECT 24.220 131.315 24.500 131.775 ;
        RECT 25.020 131.145 25.345 131.605 ;
        RECT 25.515 131.315 25.900 132.285 ;
        RECT 26.075 132.985 26.330 133.515 ;
        RECT 26.500 133.235 26.805 133.695 ;
        RECT 27.050 133.315 28.120 133.485 ;
        RECT 26.075 132.335 26.285 132.985 ;
        RECT 27.050 132.960 27.370 133.315 ;
        RECT 27.045 132.785 27.370 132.960 ;
        RECT 26.455 132.485 27.370 132.785 ;
        RECT 27.540 132.745 27.780 133.145 ;
        RECT 27.950 133.085 28.120 133.315 ;
        RECT 28.290 133.255 28.480 133.695 ;
        RECT 28.650 133.245 29.600 133.525 ;
        RECT 29.820 133.335 30.170 133.505 ;
        RECT 27.950 132.915 28.480 133.085 ;
        RECT 26.455 132.455 27.195 132.485 ;
        RECT 26.075 131.455 26.330 132.335 ;
        RECT 26.500 131.145 26.805 132.285 ;
        RECT 27.025 131.865 27.195 132.455 ;
        RECT 27.540 132.375 28.080 132.745 ;
        RECT 28.260 132.635 28.480 132.915 ;
        RECT 28.650 132.465 28.820 133.245 ;
        RECT 28.415 132.295 28.820 132.465 ;
        RECT 28.990 132.455 29.340 133.075 ;
        RECT 28.415 132.205 28.585 132.295 ;
        RECT 29.510 132.285 29.720 133.075 ;
        RECT 27.365 132.035 28.585 132.205 ;
        RECT 29.045 132.125 29.720 132.285 ;
        RECT 27.025 131.695 27.825 131.865 ;
        RECT 27.145 131.145 27.475 131.525 ;
        RECT 27.655 131.405 27.825 131.695 ;
        RECT 28.415 131.655 28.585 132.035 ;
        RECT 28.755 132.115 29.720 132.125 ;
        RECT 29.910 132.945 30.170 133.335 ;
        RECT 30.380 133.235 30.710 133.695 ;
        RECT 31.585 133.305 32.440 133.475 ;
        RECT 32.645 133.305 33.140 133.475 ;
        RECT 33.310 133.335 33.640 133.695 ;
        RECT 29.910 132.255 30.080 132.945 ;
        RECT 30.250 132.595 30.420 132.775 ;
        RECT 30.590 132.765 31.380 133.015 ;
        RECT 31.585 132.595 31.755 133.305 ;
        RECT 31.925 132.795 32.280 133.015 ;
        RECT 30.250 132.425 31.940 132.595 ;
        RECT 28.755 131.825 29.215 132.115 ;
        RECT 29.910 132.085 31.410 132.255 ;
        RECT 29.910 131.945 30.080 132.085 ;
        RECT 29.520 131.775 30.080 131.945 ;
        RECT 27.995 131.145 28.245 131.605 ;
        RECT 28.415 131.315 29.285 131.655 ;
        RECT 29.520 131.315 29.690 131.775 ;
        RECT 30.525 131.745 31.600 131.915 ;
        RECT 29.860 131.145 30.230 131.605 ;
        RECT 30.525 131.405 30.695 131.745 ;
        RECT 30.865 131.145 31.195 131.575 ;
        RECT 31.430 131.405 31.600 131.745 ;
        RECT 31.770 131.645 31.940 132.425 ;
        RECT 32.110 132.205 32.280 132.795 ;
        RECT 32.450 132.395 32.800 133.015 ;
        RECT 32.110 131.815 32.575 132.205 ;
        RECT 32.970 131.945 33.140 133.305 ;
        RECT 33.310 132.115 33.770 133.165 ;
        RECT 32.745 131.775 33.140 131.945 ;
        RECT 32.745 131.645 32.915 131.775 ;
        RECT 31.770 131.315 32.450 131.645 ;
        RECT 32.665 131.315 32.915 131.645 ;
        RECT 33.085 131.145 33.335 131.605 ;
        RECT 33.505 131.330 33.830 132.115 ;
        RECT 34.000 131.315 34.170 133.435 ;
        RECT 34.340 133.315 34.670 133.695 ;
        RECT 34.840 133.145 35.095 133.435 ;
        RECT 34.345 132.975 35.095 133.145 ;
        RECT 34.345 131.985 34.575 132.975 ;
        RECT 35.330 132.875 35.540 133.695 ;
        RECT 35.710 132.895 36.040 133.525 ;
        RECT 34.745 132.155 35.095 132.805 ;
        RECT 35.710 132.295 35.960 132.895 ;
        RECT 36.210 132.875 36.440 133.695 ;
        RECT 36.650 132.895 36.990 133.525 ;
        RECT 37.160 132.895 37.410 133.695 ;
        RECT 37.600 133.045 37.930 133.525 ;
        RECT 38.100 133.235 38.325 133.695 ;
        RECT 38.495 133.045 38.825 133.525 ;
        RECT 36.130 132.455 36.460 132.705 ;
        RECT 34.345 131.815 35.095 131.985 ;
        RECT 34.340 131.145 34.670 131.645 ;
        RECT 34.840 131.315 35.095 131.815 ;
        RECT 35.330 131.145 35.540 132.285 ;
        RECT 35.710 131.315 36.040 132.295 ;
        RECT 36.650 132.285 36.825 132.895 ;
        RECT 37.600 132.875 38.825 133.045 ;
        RECT 39.455 132.915 39.955 133.525 ;
        RECT 40.445 133.065 40.730 133.525 ;
        RECT 40.900 133.235 41.170 133.695 ;
        RECT 36.995 132.535 37.690 132.705 ;
        RECT 37.520 132.285 37.690 132.535 ;
        RECT 37.865 132.505 38.285 132.705 ;
        RECT 38.455 132.505 38.785 132.705 ;
        RECT 38.955 132.505 39.285 132.705 ;
        RECT 39.455 132.285 39.625 132.915 ;
        RECT 40.445 132.895 41.400 133.065 ;
        RECT 39.810 132.455 40.160 132.705 ;
        RECT 36.210 131.145 36.440 132.285 ;
        RECT 36.650 131.315 36.990 132.285 ;
        RECT 37.160 131.145 37.330 132.285 ;
        RECT 37.520 132.115 39.955 132.285 ;
        RECT 40.330 132.165 41.020 132.725 ;
        RECT 37.600 131.145 37.850 131.945 ;
        RECT 38.495 131.315 38.825 132.115 ;
        RECT 39.125 131.145 39.455 131.945 ;
        RECT 39.625 131.315 39.955 132.115 ;
        RECT 41.190 131.995 41.400 132.895 ;
        RECT 40.445 131.775 41.400 131.995 ;
        RECT 41.570 132.725 41.970 133.525 ;
        RECT 42.160 133.065 42.440 133.525 ;
        RECT 42.960 133.235 43.285 133.695 ;
        RECT 42.160 132.895 43.285 133.065 ;
        RECT 43.455 132.955 43.840 133.525 ;
        RECT 42.835 132.785 43.285 132.895 ;
        RECT 41.570 132.165 42.665 132.725 ;
        RECT 42.835 132.455 43.390 132.785 ;
        RECT 40.445 131.315 40.730 131.775 ;
        RECT 40.900 131.145 41.170 131.605 ;
        RECT 41.570 131.315 41.970 132.165 ;
        RECT 42.835 131.995 43.285 132.455 ;
        RECT 43.560 132.285 43.840 132.955 ;
        RECT 42.160 131.775 43.285 131.995 ;
        RECT 42.160 131.315 42.440 131.775 ;
        RECT 42.960 131.145 43.285 131.605 ;
        RECT 43.455 131.315 43.840 132.285 ;
        RECT 44.010 132.895 44.350 133.525 ;
        RECT 44.520 132.895 44.770 133.695 ;
        RECT 44.960 133.045 45.290 133.525 ;
        RECT 45.460 133.235 45.685 133.695 ;
        RECT 45.855 133.045 46.185 133.525 ;
        RECT 44.010 132.285 44.185 132.895 ;
        RECT 44.960 132.875 46.185 133.045 ;
        RECT 46.815 132.915 47.315 133.525 ;
        RECT 47.690 132.970 47.980 133.695 ;
        RECT 48.150 132.945 49.360 133.695 ;
        RECT 44.355 132.535 45.050 132.705 ;
        RECT 44.880 132.285 45.050 132.535 ;
        RECT 45.225 132.505 45.645 132.705 ;
        RECT 45.815 132.505 46.145 132.705 ;
        RECT 46.315 132.505 46.645 132.705 ;
        RECT 46.815 132.285 46.985 132.915 ;
        RECT 47.170 132.455 47.520 132.705 ;
        RECT 44.010 131.315 44.350 132.285 ;
        RECT 44.520 131.145 44.690 132.285 ;
        RECT 44.880 132.115 47.315 132.285 ;
        RECT 44.960 131.145 45.210 131.945 ;
        RECT 45.855 131.315 46.185 132.115 ;
        RECT 46.485 131.145 46.815 131.945 ;
        RECT 46.985 131.315 47.315 132.115 ;
        RECT 47.690 131.145 47.980 132.310 ;
        RECT 48.150 132.235 48.670 132.775 ;
        RECT 48.840 132.405 49.360 132.945 ;
        RECT 49.535 132.985 49.790 133.515 ;
        RECT 49.960 133.235 50.265 133.695 ;
        RECT 50.510 133.315 51.580 133.485 ;
        RECT 49.535 132.335 49.745 132.985 ;
        RECT 50.510 132.960 50.830 133.315 ;
        RECT 50.505 132.785 50.830 132.960 ;
        RECT 49.915 132.485 50.830 132.785 ;
        RECT 51.000 132.745 51.240 133.145 ;
        RECT 51.410 133.085 51.580 133.315 ;
        RECT 51.750 133.255 51.940 133.695 ;
        RECT 52.110 133.245 53.060 133.525 ;
        RECT 53.280 133.335 53.630 133.505 ;
        RECT 51.410 132.915 51.940 133.085 ;
        RECT 49.915 132.455 50.655 132.485 ;
        RECT 48.150 131.145 49.360 132.235 ;
        RECT 49.535 131.455 49.790 132.335 ;
        RECT 49.960 131.145 50.265 132.285 ;
        RECT 50.485 131.865 50.655 132.455 ;
        RECT 51.000 132.375 51.540 132.745 ;
        RECT 51.720 132.635 51.940 132.915 ;
        RECT 52.110 132.465 52.280 133.245 ;
        RECT 51.875 132.295 52.280 132.465 ;
        RECT 52.450 132.455 52.800 133.075 ;
        RECT 51.875 132.205 52.045 132.295 ;
        RECT 52.970 132.285 53.180 133.075 ;
        RECT 50.825 132.035 52.045 132.205 ;
        RECT 52.505 132.125 53.180 132.285 ;
        RECT 50.485 131.695 51.285 131.865 ;
        RECT 50.605 131.145 50.935 131.525 ;
        RECT 51.115 131.405 51.285 131.695 ;
        RECT 51.875 131.655 52.045 132.035 ;
        RECT 52.215 132.115 53.180 132.125 ;
        RECT 53.370 132.945 53.630 133.335 ;
        RECT 53.840 133.235 54.170 133.695 ;
        RECT 55.045 133.305 55.900 133.475 ;
        RECT 56.105 133.305 56.600 133.475 ;
        RECT 56.770 133.335 57.100 133.695 ;
        RECT 53.370 132.255 53.540 132.945 ;
        RECT 53.710 132.595 53.880 132.775 ;
        RECT 54.050 132.765 54.840 133.015 ;
        RECT 55.045 132.595 55.215 133.305 ;
        RECT 55.385 132.795 55.740 133.015 ;
        RECT 53.710 132.425 55.400 132.595 ;
        RECT 52.215 131.825 52.675 132.115 ;
        RECT 53.370 132.085 54.870 132.255 ;
        RECT 53.370 131.945 53.540 132.085 ;
        RECT 52.980 131.775 53.540 131.945 ;
        RECT 51.455 131.145 51.705 131.605 ;
        RECT 51.875 131.315 52.745 131.655 ;
        RECT 52.980 131.315 53.150 131.775 ;
        RECT 53.985 131.745 55.060 131.915 ;
        RECT 53.320 131.145 53.690 131.605 ;
        RECT 53.985 131.405 54.155 131.745 ;
        RECT 54.325 131.145 54.655 131.575 ;
        RECT 54.890 131.405 55.060 131.745 ;
        RECT 55.230 131.645 55.400 132.425 ;
        RECT 55.570 132.205 55.740 132.795 ;
        RECT 55.910 132.395 56.260 133.015 ;
        RECT 55.570 131.815 56.035 132.205 ;
        RECT 56.430 131.945 56.600 133.305 ;
        RECT 56.770 132.115 57.230 133.165 ;
        RECT 56.205 131.775 56.600 131.945 ;
        RECT 56.205 131.645 56.375 131.775 ;
        RECT 55.230 131.315 55.910 131.645 ;
        RECT 56.125 131.315 56.375 131.645 ;
        RECT 56.545 131.145 56.795 131.605 ;
        RECT 56.965 131.330 57.290 132.115 ;
        RECT 57.460 131.315 57.630 133.435 ;
        RECT 57.800 133.315 58.130 133.695 ;
        RECT 58.300 133.145 58.555 133.435 ;
        RECT 57.805 132.975 58.555 133.145 ;
        RECT 57.805 131.985 58.035 132.975 ;
        RECT 58.730 132.945 59.940 133.695 ;
        RECT 60.485 133.355 60.740 133.515 ;
        RECT 60.400 133.185 60.740 133.355 ;
        RECT 60.920 133.235 61.205 133.695 ;
        RECT 58.205 132.155 58.555 132.805 ;
        RECT 58.730 132.235 59.250 132.775 ;
        RECT 59.420 132.405 59.940 132.945 ;
        RECT 60.485 132.985 60.740 133.185 ;
        RECT 57.805 131.815 58.555 131.985 ;
        RECT 57.800 131.145 58.130 131.645 ;
        RECT 58.300 131.315 58.555 131.815 ;
        RECT 58.730 131.145 59.940 132.235 ;
        RECT 60.485 132.125 60.665 132.985 ;
        RECT 61.385 132.785 61.635 133.435 ;
        RECT 60.835 132.455 61.635 132.785 ;
        RECT 60.485 131.455 60.740 132.125 ;
        RECT 60.920 131.145 61.205 131.945 ;
        RECT 61.385 131.865 61.635 132.455 ;
        RECT 61.835 133.100 62.155 133.430 ;
        RECT 62.335 133.215 62.995 133.695 ;
        RECT 63.195 133.305 64.045 133.475 ;
        RECT 61.835 132.205 62.025 133.100 ;
        RECT 62.345 132.775 63.005 133.045 ;
        RECT 62.675 132.715 63.005 132.775 ;
        RECT 62.195 132.545 62.525 132.605 ;
        RECT 63.195 132.545 63.365 133.305 ;
        RECT 64.605 133.235 64.925 133.695 ;
        RECT 65.125 133.055 65.375 133.485 ;
        RECT 65.665 133.255 66.075 133.695 ;
        RECT 66.245 133.315 67.260 133.515 ;
        RECT 63.535 132.885 64.785 133.055 ;
        RECT 63.535 132.765 63.865 132.885 ;
        RECT 62.195 132.375 64.095 132.545 ;
        RECT 61.835 132.035 63.755 132.205 ;
        RECT 61.835 132.015 62.155 132.035 ;
        RECT 61.385 131.355 61.715 131.865 ;
        RECT 61.985 131.405 62.155 132.015 ;
        RECT 63.925 131.865 64.095 132.375 ;
        RECT 64.265 132.305 64.445 132.715 ;
        RECT 64.615 132.125 64.785 132.885 ;
        RECT 62.325 131.145 62.655 131.835 ;
        RECT 62.885 131.695 64.095 131.865 ;
        RECT 64.265 131.815 64.785 132.125 ;
        RECT 64.955 132.715 65.375 133.055 ;
        RECT 65.665 132.715 66.075 133.045 ;
        RECT 64.955 131.945 65.145 132.715 ;
        RECT 66.245 132.585 66.415 133.315 ;
        RECT 67.560 133.145 67.730 133.475 ;
        RECT 67.900 133.315 68.230 133.695 ;
        RECT 66.585 132.765 66.935 133.135 ;
        RECT 66.245 132.545 66.665 132.585 ;
        RECT 65.315 132.375 66.665 132.545 ;
        RECT 65.315 132.215 65.565 132.375 ;
        RECT 66.075 131.945 66.325 132.205 ;
        RECT 64.955 131.695 66.325 131.945 ;
        RECT 62.885 131.405 63.125 131.695 ;
        RECT 63.925 131.615 64.095 131.695 ;
        RECT 63.325 131.145 63.745 131.525 ;
        RECT 63.925 131.365 64.555 131.615 ;
        RECT 65.025 131.145 65.355 131.525 ;
        RECT 65.525 131.405 65.695 131.695 ;
        RECT 66.495 131.530 66.665 132.375 ;
        RECT 67.115 132.205 67.335 133.075 ;
        RECT 67.560 132.955 68.255 133.145 ;
        RECT 66.835 131.825 67.335 132.205 ;
        RECT 67.505 132.155 67.915 132.775 ;
        RECT 68.085 131.985 68.255 132.955 ;
        RECT 67.560 131.815 68.255 131.985 ;
        RECT 65.875 131.145 66.255 131.525 ;
        RECT 66.495 131.360 67.325 131.530 ;
        RECT 67.560 131.315 67.730 131.815 ;
        RECT 67.900 131.145 68.230 131.645 ;
        RECT 68.445 131.315 68.670 133.435 ;
        RECT 68.840 133.315 69.170 133.695 ;
        RECT 69.340 133.145 69.510 133.435 ;
        RECT 68.845 132.975 69.510 133.145 ;
        RECT 68.845 131.985 69.075 132.975 ;
        RECT 70.230 132.925 71.900 133.695 ;
        RECT 69.245 132.155 69.595 132.805 ;
        RECT 70.230 132.235 70.980 132.755 ;
        RECT 71.150 132.405 71.900 132.925 ;
        RECT 72.110 132.875 72.340 133.695 ;
        RECT 72.510 132.895 72.840 133.525 ;
        RECT 72.090 132.455 72.420 132.705 ;
        RECT 72.590 132.295 72.840 132.895 ;
        RECT 73.010 132.875 73.220 133.695 ;
        RECT 73.450 132.970 73.740 133.695 ;
        RECT 74.285 132.985 74.540 133.515 ;
        RECT 74.720 133.235 75.005 133.695 ;
        RECT 68.845 131.815 69.510 131.985 ;
        RECT 68.840 131.145 69.170 131.645 ;
        RECT 69.340 131.315 69.510 131.815 ;
        RECT 70.230 131.145 71.900 132.235 ;
        RECT 72.110 131.145 72.340 132.285 ;
        RECT 72.510 131.315 72.840 132.295 ;
        RECT 73.010 131.145 73.220 132.285 ;
        RECT 73.450 131.145 73.740 132.310 ;
        RECT 74.285 132.125 74.465 132.985 ;
        RECT 75.185 132.785 75.435 133.435 ;
        RECT 74.635 132.455 75.435 132.785 ;
        RECT 74.285 131.655 74.540 132.125 ;
        RECT 74.200 131.485 74.540 131.655 ;
        RECT 74.285 131.455 74.540 131.485 ;
        RECT 74.720 131.145 75.005 131.945 ;
        RECT 75.185 131.865 75.435 132.455 ;
        RECT 75.635 133.100 75.955 133.430 ;
        RECT 76.135 133.215 76.795 133.695 ;
        RECT 76.995 133.305 77.845 133.475 ;
        RECT 75.635 132.205 75.825 133.100 ;
        RECT 76.145 132.775 76.805 133.045 ;
        RECT 76.475 132.715 76.805 132.775 ;
        RECT 75.995 132.545 76.325 132.605 ;
        RECT 76.995 132.545 77.165 133.305 ;
        RECT 78.405 133.235 78.725 133.695 ;
        RECT 78.925 133.055 79.175 133.485 ;
        RECT 79.465 133.255 79.875 133.695 ;
        RECT 80.045 133.315 81.060 133.515 ;
        RECT 77.335 132.885 78.585 133.055 ;
        RECT 77.335 132.765 77.665 132.885 ;
        RECT 75.995 132.375 77.895 132.545 ;
        RECT 75.635 132.035 77.555 132.205 ;
        RECT 75.635 132.015 75.955 132.035 ;
        RECT 75.185 131.355 75.515 131.865 ;
        RECT 75.785 131.405 75.955 132.015 ;
        RECT 77.725 131.865 77.895 132.375 ;
        RECT 78.065 132.305 78.245 132.715 ;
        RECT 78.415 132.125 78.585 132.885 ;
        RECT 76.125 131.145 76.455 131.835 ;
        RECT 76.685 131.695 77.895 131.865 ;
        RECT 78.065 131.815 78.585 132.125 ;
        RECT 78.755 132.715 79.175 133.055 ;
        RECT 79.465 132.715 79.875 133.045 ;
        RECT 78.755 131.945 78.945 132.715 ;
        RECT 80.045 132.585 80.215 133.315 ;
        RECT 81.360 133.145 81.530 133.475 ;
        RECT 81.700 133.315 82.030 133.695 ;
        RECT 80.385 132.765 80.735 133.135 ;
        RECT 80.045 132.545 80.465 132.585 ;
        RECT 79.115 132.375 80.465 132.545 ;
        RECT 79.115 132.215 79.365 132.375 ;
        RECT 79.875 131.945 80.125 132.205 ;
        RECT 78.755 131.695 80.125 131.945 ;
        RECT 76.685 131.405 76.925 131.695 ;
        RECT 77.725 131.615 77.895 131.695 ;
        RECT 77.125 131.145 77.545 131.525 ;
        RECT 77.725 131.365 78.355 131.615 ;
        RECT 78.825 131.145 79.155 131.525 ;
        RECT 79.325 131.405 79.495 131.695 ;
        RECT 80.295 131.530 80.465 132.375 ;
        RECT 80.915 132.205 81.135 133.075 ;
        RECT 81.360 132.955 82.055 133.145 ;
        RECT 80.635 131.825 81.135 132.205 ;
        RECT 81.305 132.155 81.715 132.775 ;
        RECT 81.885 131.985 82.055 132.955 ;
        RECT 81.360 131.815 82.055 131.985 ;
        RECT 79.675 131.145 80.055 131.525 ;
        RECT 80.295 131.360 81.125 131.530 ;
        RECT 81.360 131.315 81.530 131.815 ;
        RECT 81.700 131.145 82.030 131.645 ;
        RECT 82.245 131.315 82.470 133.435 ;
        RECT 82.640 133.315 82.970 133.695 ;
        RECT 83.140 133.145 83.310 133.435 ;
        RECT 83.570 133.185 83.875 133.695 ;
        RECT 82.645 132.975 83.310 133.145 ;
        RECT 82.645 131.985 82.875 132.975 ;
        RECT 83.045 132.155 83.395 132.805 ;
        RECT 83.570 132.455 83.885 133.015 ;
        RECT 84.055 132.705 84.305 133.515 ;
        RECT 84.475 133.170 84.735 133.695 ;
        RECT 84.915 132.705 85.165 133.515 ;
        RECT 85.335 133.135 85.595 133.695 ;
        RECT 85.765 133.045 86.025 133.500 ;
        RECT 86.195 133.215 86.455 133.695 ;
        RECT 86.625 133.045 86.885 133.500 ;
        RECT 87.055 133.215 87.315 133.695 ;
        RECT 87.485 133.045 87.745 133.500 ;
        RECT 87.915 133.215 88.160 133.695 ;
        RECT 88.330 133.045 88.605 133.500 ;
        RECT 88.775 133.215 89.020 133.695 ;
        RECT 89.190 133.045 89.450 133.500 ;
        RECT 89.630 133.215 89.880 133.695 ;
        RECT 90.050 133.045 90.310 133.500 ;
        RECT 90.490 133.215 90.740 133.695 ;
        RECT 90.910 133.045 91.170 133.500 ;
        RECT 91.350 133.215 91.610 133.695 ;
        RECT 91.780 133.045 92.040 133.500 ;
        RECT 92.210 133.215 92.510 133.695 ;
        RECT 85.765 132.875 92.510 133.045 ;
        RECT 93.230 132.925 94.900 133.695 ;
        RECT 84.055 132.455 91.175 132.705 ;
        RECT 91.345 132.675 92.510 132.875 ;
        RECT 91.345 132.505 92.540 132.675 ;
        RECT 82.645 131.815 83.310 131.985 ;
        RECT 82.640 131.145 82.970 131.645 ;
        RECT 83.140 131.315 83.310 131.815 ;
        RECT 83.580 131.145 83.875 131.955 ;
        RECT 84.055 131.315 84.300 132.455 ;
        RECT 84.475 131.145 84.735 131.955 ;
        RECT 84.915 131.320 85.165 132.455 ;
        RECT 91.345 132.285 92.510 132.505 ;
        RECT 85.765 132.060 92.510 132.285 ;
        RECT 93.230 132.235 93.980 132.755 ;
        RECT 94.150 132.405 94.900 132.925 ;
        RECT 95.345 132.885 95.590 133.490 ;
        RECT 95.810 133.160 96.320 133.695 ;
        RECT 95.070 132.715 96.300 132.885 ;
        RECT 85.765 132.045 91.170 132.060 ;
        RECT 85.335 131.150 85.595 131.945 ;
        RECT 85.765 131.320 86.025 132.045 ;
        RECT 86.195 131.150 86.455 131.875 ;
        RECT 86.625 131.320 86.885 132.045 ;
        RECT 87.055 131.150 87.315 131.875 ;
        RECT 87.485 131.320 87.745 132.045 ;
        RECT 87.915 131.150 88.175 131.875 ;
        RECT 88.345 131.320 88.605 132.045 ;
        RECT 88.775 131.150 89.020 131.875 ;
        RECT 89.190 131.320 89.450 132.045 ;
        RECT 89.635 131.150 89.880 131.875 ;
        RECT 90.050 131.320 90.310 132.045 ;
        RECT 90.495 131.150 90.740 131.875 ;
        RECT 90.910 131.320 91.170 132.045 ;
        RECT 91.355 131.150 91.610 131.875 ;
        RECT 91.780 131.320 92.070 132.060 ;
        RECT 85.335 131.145 91.610 131.150 ;
        RECT 92.240 131.145 92.510 131.890 ;
        RECT 93.230 131.145 94.900 132.235 ;
        RECT 95.070 131.905 95.410 132.715 ;
        RECT 95.580 132.150 96.330 132.340 ;
        RECT 95.070 131.495 95.585 131.905 ;
        RECT 95.820 131.145 95.990 131.905 ;
        RECT 96.160 131.485 96.330 132.150 ;
        RECT 96.500 132.165 96.690 133.525 ;
        RECT 96.860 133.015 97.135 133.525 ;
        RECT 97.325 133.160 97.855 133.525 ;
        RECT 98.280 133.295 98.610 133.695 ;
        RECT 97.680 133.125 97.855 133.160 ;
        RECT 96.860 132.845 97.140 133.015 ;
        RECT 96.860 132.365 97.135 132.845 ;
        RECT 97.340 132.165 97.510 132.965 ;
        RECT 96.500 131.995 97.510 132.165 ;
        RECT 97.680 132.955 98.610 133.125 ;
        RECT 98.780 132.955 99.035 133.525 ;
        RECT 99.210 132.970 99.500 133.695 ;
        RECT 100.595 133.145 100.850 133.435 ;
        RECT 101.020 133.315 101.350 133.695 ;
        RECT 100.595 132.975 101.345 133.145 ;
        RECT 97.680 131.825 97.850 132.955 ;
        RECT 98.440 132.785 98.610 132.955 ;
        RECT 96.725 131.655 97.850 131.825 ;
        RECT 98.020 132.455 98.215 132.785 ;
        RECT 98.440 132.455 98.695 132.785 ;
        RECT 98.020 131.485 98.190 132.455 ;
        RECT 98.865 132.285 99.035 132.955 ;
        RECT 96.160 131.315 98.190 131.485 ;
        RECT 98.360 131.145 98.530 132.285 ;
        RECT 98.700 131.315 99.035 132.285 ;
        RECT 99.210 131.145 99.500 132.310 ;
        RECT 100.595 132.155 100.945 132.805 ;
        RECT 101.115 131.985 101.345 132.975 ;
        RECT 100.595 131.815 101.345 131.985 ;
        RECT 100.595 131.315 100.850 131.815 ;
        RECT 101.020 131.145 101.350 131.645 ;
        RECT 101.520 131.315 101.690 133.435 ;
        RECT 102.050 133.335 102.380 133.695 ;
        RECT 102.550 133.305 103.045 133.475 ;
        RECT 103.250 133.305 104.105 133.475 ;
        RECT 101.920 132.115 102.380 133.165 ;
        RECT 101.860 131.330 102.185 132.115 ;
        RECT 102.550 131.945 102.720 133.305 ;
        RECT 102.890 132.395 103.240 133.015 ;
        RECT 103.410 132.795 103.765 133.015 ;
        RECT 103.410 132.205 103.580 132.795 ;
        RECT 103.935 132.595 104.105 133.305 ;
        RECT 104.980 133.235 105.310 133.695 ;
        RECT 105.520 133.335 105.870 133.505 ;
        RECT 104.310 132.765 105.100 133.015 ;
        RECT 105.520 132.945 105.780 133.335 ;
        RECT 106.090 133.245 107.040 133.525 ;
        RECT 107.210 133.255 107.400 133.695 ;
        RECT 107.570 133.315 108.640 133.485 ;
        RECT 105.270 132.595 105.440 132.775 ;
        RECT 102.550 131.775 102.945 131.945 ;
        RECT 103.115 131.815 103.580 132.205 ;
        RECT 103.750 132.425 105.440 132.595 ;
        RECT 102.775 131.645 102.945 131.775 ;
        RECT 103.750 131.645 103.920 132.425 ;
        RECT 105.610 132.255 105.780 132.945 ;
        RECT 104.280 132.085 105.780 132.255 ;
        RECT 105.970 132.285 106.180 133.075 ;
        RECT 106.350 132.455 106.700 133.075 ;
        RECT 106.870 132.465 107.040 133.245 ;
        RECT 107.570 133.085 107.740 133.315 ;
        RECT 107.210 132.915 107.740 133.085 ;
        RECT 107.210 132.635 107.430 132.915 ;
        RECT 107.910 132.745 108.150 133.145 ;
        RECT 106.870 132.295 107.275 132.465 ;
        RECT 107.610 132.375 108.150 132.745 ;
        RECT 108.320 132.960 108.640 133.315 ;
        RECT 108.320 132.705 108.645 132.960 ;
        RECT 108.840 132.885 109.010 133.695 ;
        RECT 109.180 133.045 109.510 133.525 ;
        RECT 109.680 133.225 109.850 133.695 ;
        RECT 110.020 133.045 110.350 133.525 ;
        RECT 110.520 133.225 110.690 133.695 ;
        RECT 109.180 132.875 110.945 133.045 ;
        RECT 111.170 132.945 112.380 133.695 ;
        RECT 108.320 132.495 110.350 132.705 ;
        RECT 108.320 132.485 108.665 132.495 ;
        RECT 105.970 132.125 106.645 132.285 ;
        RECT 107.105 132.205 107.275 132.295 ;
        RECT 105.970 132.115 106.935 132.125 ;
        RECT 105.610 131.945 105.780 132.085 ;
        RECT 102.355 131.145 102.605 131.605 ;
        RECT 102.775 131.315 103.025 131.645 ;
        RECT 103.240 131.315 103.920 131.645 ;
        RECT 104.090 131.745 105.165 131.915 ;
        RECT 105.610 131.775 106.170 131.945 ;
        RECT 106.475 131.825 106.935 132.115 ;
        RECT 107.105 132.035 108.325 132.205 ;
        RECT 104.090 131.405 104.260 131.745 ;
        RECT 104.495 131.145 104.825 131.575 ;
        RECT 104.995 131.405 105.165 131.745 ;
        RECT 105.460 131.145 105.830 131.605 ;
        RECT 106.000 131.315 106.170 131.775 ;
        RECT 107.105 131.655 107.275 132.035 ;
        RECT 108.495 131.865 108.665 132.485 ;
        RECT 110.535 132.325 110.945 132.875 ;
        RECT 106.405 131.315 107.275 131.655 ;
        RECT 107.865 131.695 108.665 131.865 ;
        RECT 107.445 131.145 107.695 131.605 ;
        RECT 107.865 131.405 108.035 131.695 ;
        RECT 108.215 131.145 108.545 131.525 ;
        RECT 108.840 131.145 109.010 132.205 ;
        RECT 109.220 132.155 110.945 132.325 ;
        RECT 111.170 132.235 111.690 132.775 ;
        RECT 111.860 132.405 112.380 132.945 ;
        RECT 109.220 131.315 109.510 132.155 ;
        RECT 109.680 131.145 109.850 131.985 ;
        RECT 110.060 131.315 110.310 132.155 ;
        RECT 110.520 131.145 110.690 131.985 ;
        RECT 111.170 131.145 112.380 132.235 ;
        RECT 18.165 130.975 112.465 131.145 ;
        RECT 18.250 129.885 19.460 130.975 ;
        RECT 19.940 130.135 20.110 130.975 ;
        RECT 20.320 129.965 20.570 130.805 ;
        RECT 20.780 130.135 20.950 130.975 ;
        RECT 21.120 129.965 21.410 130.805 ;
        RECT 18.250 129.175 18.770 129.715 ;
        RECT 18.940 129.345 19.460 129.885 ;
        RECT 19.685 129.795 21.410 129.965 ;
        RECT 21.620 129.915 21.790 130.975 ;
        RECT 22.085 130.595 22.415 130.975 ;
        RECT 22.595 130.425 22.765 130.715 ;
        RECT 22.935 130.515 23.185 130.975 ;
        RECT 21.965 130.255 22.765 130.425 ;
        RECT 23.355 130.465 24.225 130.805 ;
        RECT 19.685 129.245 20.095 129.795 ;
        RECT 21.965 129.635 22.135 130.255 ;
        RECT 23.355 130.085 23.525 130.465 ;
        RECT 24.460 130.345 24.630 130.805 ;
        RECT 24.800 130.515 25.170 130.975 ;
        RECT 25.465 130.375 25.635 130.715 ;
        RECT 25.805 130.545 26.135 130.975 ;
        RECT 26.370 130.375 26.540 130.715 ;
        RECT 22.305 129.915 23.525 130.085 ;
        RECT 23.695 130.005 24.155 130.295 ;
        RECT 24.460 130.175 25.020 130.345 ;
        RECT 25.465 130.205 26.540 130.375 ;
        RECT 26.710 130.475 27.390 130.805 ;
        RECT 27.605 130.475 27.855 130.805 ;
        RECT 28.025 130.515 28.275 130.975 ;
        RECT 24.850 130.035 25.020 130.175 ;
        RECT 23.695 129.995 24.660 130.005 ;
        RECT 23.355 129.825 23.525 129.915 ;
        RECT 23.985 129.835 24.660 129.995 ;
        RECT 21.965 129.625 22.310 129.635 ;
        RECT 20.280 129.415 22.310 129.625 ;
        RECT 18.250 128.425 19.460 129.175 ;
        RECT 19.685 129.075 21.450 129.245 ;
        RECT 19.940 128.425 20.110 128.895 ;
        RECT 20.280 128.595 20.610 129.075 ;
        RECT 20.780 128.425 20.950 128.895 ;
        RECT 21.120 128.595 21.450 129.075 ;
        RECT 21.620 128.425 21.790 129.235 ;
        RECT 21.985 129.160 22.310 129.415 ;
        RECT 21.990 128.805 22.310 129.160 ;
        RECT 22.480 129.375 23.020 129.745 ;
        RECT 23.355 129.655 23.760 129.825 ;
        RECT 22.480 128.975 22.720 129.375 ;
        RECT 23.200 129.205 23.420 129.485 ;
        RECT 22.890 129.035 23.420 129.205 ;
        RECT 22.890 128.805 23.060 129.035 ;
        RECT 23.590 128.875 23.760 129.655 ;
        RECT 23.930 129.045 24.280 129.665 ;
        RECT 24.450 129.045 24.660 129.835 ;
        RECT 24.850 129.865 26.350 130.035 ;
        RECT 24.850 129.175 25.020 129.865 ;
        RECT 26.710 129.695 26.880 130.475 ;
        RECT 27.685 130.345 27.855 130.475 ;
        RECT 25.190 129.525 26.880 129.695 ;
        RECT 27.050 129.915 27.515 130.305 ;
        RECT 27.685 130.175 28.080 130.345 ;
        RECT 25.190 129.345 25.360 129.525 ;
        RECT 21.990 128.635 23.060 128.805 ;
        RECT 23.230 128.425 23.420 128.865 ;
        RECT 23.590 128.595 24.540 128.875 ;
        RECT 24.850 128.785 25.110 129.175 ;
        RECT 25.530 129.105 26.320 129.355 ;
        RECT 24.760 128.615 25.110 128.785 ;
        RECT 25.320 128.425 25.650 128.885 ;
        RECT 26.525 128.815 26.695 129.525 ;
        RECT 27.050 129.325 27.220 129.915 ;
        RECT 26.865 129.105 27.220 129.325 ;
        RECT 27.390 129.105 27.740 129.725 ;
        RECT 27.910 128.815 28.080 130.175 ;
        RECT 28.445 130.005 28.770 130.790 ;
        RECT 28.250 128.955 28.710 130.005 ;
        RECT 26.525 128.645 27.380 128.815 ;
        RECT 27.585 128.645 28.080 128.815 ;
        RECT 28.250 128.425 28.580 128.785 ;
        RECT 28.940 128.685 29.110 130.805 ;
        RECT 29.280 130.475 29.610 130.975 ;
        RECT 29.780 130.305 30.035 130.805 ;
        RECT 29.285 130.135 30.035 130.305 ;
        RECT 30.210 130.215 30.725 130.625 ;
        RECT 30.960 130.215 31.130 130.975 ;
        RECT 31.300 130.635 33.330 130.805 ;
        RECT 29.285 129.145 29.515 130.135 ;
        RECT 29.685 129.315 30.035 129.965 ;
        RECT 30.210 129.405 30.550 130.215 ;
        RECT 31.300 129.970 31.470 130.635 ;
        RECT 31.865 130.295 32.990 130.465 ;
        RECT 30.720 129.780 31.470 129.970 ;
        RECT 31.640 129.955 32.650 130.125 ;
        RECT 30.210 129.235 31.440 129.405 ;
        RECT 29.285 128.975 30.035 129.145 ;
        RECT 29.280 128.425 29.610 128.805 ;
        RECT 29.780 128.685 30.035 128.975 ;
        RECT 30.485 128.630 30.730 129.235 ;
        RECT 30.950 128.425 31.460 128.960 ;
        RECT 31.640 128.595 31.830 129.955 ;
        RECT 32.000 129.615 32.275 129.755 ;
        RECT 32.000 129.445 32.280 129.615 ;
        RECT 32.000 128.595 32.275 129.445 ;
        RECT 32.480 129.155 32.650 129.955 ;
        RECT 32.820 129.165 32.990 130.295 ;
        RECT 33.160 129.665 33.330 130.635 ;
        RECT 33.500 129.835 33.670 130.975 ;
        RECT 33.840 129.835 34.175 130.805 ;
        RECT 33.160 129.335 33.355 129.665 ;
        RECT 33.580 129.335 33.835 129.665 ;
        RECT 33.580 129.165 33.750 129.335 ;
        RECT 34.005 129.165 34.175 129.835 ;
        RECT 34.810 129.810 35.100 130.975 ;
        RECT 35.820 130.230 36.090 130.975 ;
        RECT 36.720 130.970 42.995 130.975 ;
        RECT 36.260 130.060 36.550 130.800 ;
        RECT 36.720 130.245 36.975 130.970 ;
        RECT 37.160 130.075 37.420 130.800 ;
        RECT 37.590 130.245 37.835 130.970 ;
        RECT 38.020 130.075 38.280 130.800 ;
        RECT 38.450 130.245 38.695 130.970 ;
        RECT 38.880 130.075 39.140 130.800 ;
        RECT 39.310 130.245 39.555 130.970 ;
        RECT 39.725 130.075 39.985 130.800 ;
        RECT 40.155 130.245 40.415 130.970 ;
        RECT 40.585 130.075 40.845 130.800 ;
        RECT 41.015 130.245 41.275 130.970 ;
        RECT 41.445 130.075 41.705 130.800 ;
        RECT 41.875 130.245 42.135 130.970 ;
        RECT 42.305 130.075 42.565 130.800 ;
        RECT 42.735 130.175 42.995 130.970 ;
        RECT 37.160 130.060 42.565 130.075 ;
        RECT 35.820 129.835 42.565 130.060 ;
        RECT 35.820 129.275 36.985 129.835 ;
        RECT 43.165 129.665 43.415 130.800 ;
        RECT 43.595 130.165 43.855 130.975 ;
        RECT 44.030 129.665 44.275 130.805 ;
        RECT 44.455 130.165 44.750 130.975 ;
        RECT 45.500 130.175 45.670 130.975 ;
        RECT 45.840 129.955 46.170 130.805 ;
        RECT 46.340 130.175 46.510 130.975 ;
        RECT 46.680 129.955 47.010 130.805 ;
        RECT 47.180 130.175 47.350 130.975 ;
        RECT 47.520 129.955 47.850 130.805 ;
        RECT 48.020 130.175 48.190 130.975 ;
        RECT 48.360 129.955 48.690 130.805 ;
        RECT 48.860 130.175 49.030 130.975 ;
        RECT 49.200 129.955 49.530 130.805 ;
        RECT 49.700 130.175 49.870 130.975 ;
        RECT 50.040 129.955 50.370 130.805 ;
        RECT 50.540 130.175 50.710 130.975 ;
        RECT 50.880 129.955 51.210 130.805 ;
        RECT 51.380 130.175 51.550 130.975 ;
        RECT 51.720 129.955 52.050 130.805 ;
        RECT 52.220 130.175 52.390 130.975 ;
        RECT 52.560 129.955 52.890 130.805 ;
        RECT 53.060 130.175 53.230 130.975 ;
        RECT 53.400 129.955 53.730 130.805 ;
        RECT 53.900 130.175 54.070 130.975 ;
        RECT 54.240 129.955 54.570 130.805 ;
        RECT 54.740 130.125 54.910 130.975 ;
        RECT 55.080 129.955 55.410 130.805 ;
        RECT 55.580 130.125 55.750 130.975 ;
        RECT 55.920 129.955 56.250 130.805 ;
        RECT 45.390 129.785 52.050 129.955 ;
        RECT 52.220 129.785 54.570 129.955 ;
        RECT 54.740 129.785 56.250 129.955 ;
        RECT 56.430 129.885 59.020 130.975 ;
        RECT 37.155 129.415 44.275 129.665 ;
        RECT 32.820 128.995 33.750 129.165 ;
        RECT 32.820 128.960 32.995 128.995 ;
        RECT 32.465 128.595 32.995 128.960 ;
        RECT 33.420 128.425 33.750 128.825 ;
        RECT 33.920 128.595 34.175 129.165 ;
        RECT 35.790 129.245 36.985 129.275 ;
        RECT 34.810 128.425 35.100 129.150 ;
        RECT 35.790 129.105 42.565 129.245 ;
        RECT 35.820 129.075 42.565 129.105 ;
        RECT 35.820 128.425 36.120 128.905 ;
        RECT 36.290 128.620 36.550 129.075 ;
        RECT 36.720 128.425 36.980 128.905 ;
        RECT 37.160 128.620 37.420 129.075 ;
        RECT 37.590 128.425 37.840 128.905 ;
        RECT 38.020 128.620 38.280 129.075 ;
        RECT 38.450 128.425 38.700 128.905 ;
        RECT 38.880 128.620 39.140 129.075 ;
        RECT 39.310 128.425 39.555 128.905 ;
        RECT 39.725 128.620 40.000 129.075 ;
        RECT 40.170 128.425 40.415 128.905 ;
        RECT 40.585 128.620 40.845 129.075 ;
        RECT 41.015 128.425 41.275 128.905 ;
        RECT 41.445 128.620 41.705 129.075 ;
        RECT 41.875 128.425 42.135 128.905 ;
        RECT 42.305 128.620 42.565 129.075 ;
        RECT 42.735 128.425 42.995 128.985 ;
        RECT 43.165 128.605 43.415 129.415 ;
        RECT 43.595 128.425 43.855 128.950 ;
        RECT 44.025 128.605 44.275 129.415 ;
        RECT 44.445 129.105 44.760 129.665 ;
        RECT 45.390 129.245 45.665 129.785 ;
        RECT 52.220 129.615 52.395 129.785 ;
        RECT 54.740 129.615 54.910 129.785 ;
        RECT 45.835 129.415 52.395 129.615 ;
        RECT 52.600 129.415 54.910 129.615 ;
        RECT 55.080 129.415 56.255 129.615 ;
        RECT 52.220 129.245 52.395 129.415 ;
        RECT 54.740 129.245 54.910 129.415 ;
        RECT 56.430 129.365 57.640 129.885 ;
        RECT 59.230 129.835 59.460 130.975 ;
        RECT 59.630 129.825 59.960 130.805 ;
        RECT 60.130 129.835 60.340 130.975 ;
        RECT 45.390 129.075 52.050 129.245 ;
        RECT 52.220 129.075 54.570 129.245 ;
        RECT 54.740 129.075 56.250 129.245 ;
        RECT 57.810 129.195 59.020 129.715 ;
        RECT 59.210 129.415 59.540 129.665 ;
        RECT 44.455 128.425 44.760 128.935 ;
        RECT 45.500 128.425 45.670 128.905 ;
        RECT 45.840 128.600 46.170 129.075 ;
        RECT 46.340 128.425 46.510 128.905 ;
        RECT 46.680 128.600 47.010 129.075 ;
        RECT 47.180 128.425 47.350 128.905 ;
        RECT 47.520 128.600 47.850 129.075 ;
        RECT 48.020 128.425 48.190 128.905 ;
        RECT 48.360 128.600 48.690 129.075 ;
        RECT 48.860 128.425 49.030 128.905 ;
        RECT 49.200 128.600 49.530 129.075 ;
        RECT 49.700 128.425 49.870 128.905 ;
        RECT 50.040 128.600 50.370 129.075 ;
        RECT 50.120 128.595 50.290 128.600 ;
        RECT 50.540 128.425 50.710 128.905 ;
        RECT 50.880 128.600 51.210 129.075 ;
        RECT 50.960 128.595 51.130 128.600 ;
        RECT 51.380 128.425 51.550 128.905 ;
        RECT 51.720 128.600 52.050 129.075 ;
        RECT 51.800 128.595 52.050 128.600 ;
        RECT 52.220 128.425 52.390 128.905 ;
        RECT 52.560 128.600 52.890 129.075 ;
        RECT 53.060 128.425 53.230 128.905 ;
        RECT 53.400 128.600 53.730 129.075 ;
        RECT 53.900 128.425 54.070 128.905 ;
        RECT 54.240 128.600 54.570 129.075 ;
        RECT 54.740 128.425 54.910 128.905 ;
        RECT 55.080 128.600 55.410 129.075 ;
        RECT 55.580 128.425 55.750 128.905 ;
        RECT 55.920 128.600 56.250 129.075 ;
        RECT 56.430 128.425 59.020 129.195 ;
        RECT 59.230 128.425 59.460 129.245 ;
        RECT 59.710 129.225 59.960 129.825 ;
        RECT 60.570 129.810 60.860 130.975 ;
        RECT 61.030 130.215 61.545 130.625 ;
        RECT 61.780 130.215 61.950 130.975 ;
        RECT 62.120 130.635 64.150 130.805 ;
        RECT 61.030 129.405 61.370 130.215 ;
        RECT 62.120 129.970 62.290 130.635 ;
        RECT 62.685 130.295 63.810 130.465 ;
        RECT 61.540 129.780 62.290 129.970 ;
        RECT 62.460 129.955 63.470 130.125 ;
        RECT 59.630 128.595 59.960 129.225 ;
        RECT 60.130 128.425 60.340 129.245 ;
        RECT 61.030 129.235 62.260 129.405 ;
        RECT 60.570 128.425 60.860 129.150 ;
        RECT 61.305 128.630 61.550 129.235 ;
        RECT 61.770 128.425 62.280 128.960 ;
        RECT 62.460 128.595 62.650 129.955 ;
        RECT 62.820 129.275 63.095 129.755 ;
        RECT 62.820 129.105 63.100 129.275 ;
        RECT 63.300 129.155 63.470 129.955 ;
        RECT 63.640 129.165 63.810 130.295 ;
        RECT 63.980 129.665 64.150 130.635 ;
        RECT 64.320 129.835 64.490 130.975 ;
        RECT 64.660 129.835 64.995 130.805 ;
        RECT 63.980 129.335 64.175 129.665 ;
        RECT 64.400 129.335 64.655 129.665 ;
        RECT 64.400 129.165 64.570 129.335 ;
        RECT 64.825 129.165 64.995 129.835 ;
        RECT 65.170 129.885 66.840 130.975 ;
        RECT 65.170 129.365 65.920 129.885 ;
        RECT 67.015 129.785 67.270 130.665 ;
        RECT 67.440 129.835 67.745 130.975 ;
        RECT 68.085 130.595 68.415 130.975 ;
        RECT 68.595 130.425 68.765 130.715 ;
        RECT 68.935 130.515 69.185 130.975 ;
        RECT 67.965 130.255 68.765 130.425 ;
        RECT 69.355 130.465 70.225 130.805 ;
        RECT 66.090 129.195 66.840 129.715 ;
        RECT 62.820 128.595 63.095 129.105 ;
        RECT 63.640 128.995 64.570 129.165 ;
        RECT 63.640 128.960 63.815 128.995 ;
        RECT 63.285 128.595 63.815 128.960 ;
        RECT 64.240 128.425 64.570 128.825 ;
        RECT 64.740 128.595 64.995 129.165 ;
        RECT 65.170 128.425 66.840 129.195 ;
        RECT 67.015 129.135 67.225 129.785 ;
        RECT 67.965 129.665 68.135 130.255 ;
        RECT 69.355 130.085 69.525 130.465 ;
        RECT 70.460 130.345 70.630 130.805 ;
        RECT 70.800 130.515 71.170 130.975 ;
        RECT 71.465 130.375 71.635 130.715 ;
        RECT 71.805 130.545 72.135 130.975 ;
        RECT 72.370 130.375 72.540 130.715 ;
        RECT 68.305 129.915 69.525 130.085 ;
        RECT 69.695 130.005 70.155 130.295 ;
        RECT 70.460 130.175 71.020 130.345 ;
        RECT 71.465 130.205 72.540 130.375 ;
        RECT 72.710 130.475 73.390 130.805 ;
        RECT 73.605 130.475 73.855 130.805 ;
        RECT 74.025 130.515 74.275 130.975 ;
        RECT 70.850 130.035 71.020 130.175 ;
        RECT 69.695 129.995 70.660 130.005 ;
        RECT 69.355 129.825 69.525 129.915 ;
        RECT 69.985 129.835 70.660 129.995 ;
        RECT 67.395 129.635 68.135 129.665 ;
        RECT 67.395 129.335 68.310 129.635 ;
        RECT 67.985 129.160 68.310 129.335 ;
        RECT 67.015 128.605 67.270 129.135 ;
        RECT 67.440 128.425 67.745 128.885 ;
        RECT 67.990 128.805 68.310 129.160 ;
        RECT 68.480 129.375 69.020 129.745 ;
        RECT 69.355 129.655 69.760 129.825 ;
        RECT 68.480 128.975 68.720 129.375 ;
        RECT 69.200 129.205 69.420 129.485 ;
        RECT 68.890 129.035 69.420 129.205 ;
        RECT 68.890 128.805 69.060 129.035 ;
        RECT 69.590 128.875 69.760 129.655 ;
        RECT 69.930 129.045 70.280 129.665 ;
        RECT 70.450 129.045 70.660 129.835 ;
        RECT 70.850 129.865 72.350 130.035 ;
        RECT 70.850 129.175 71.020 129.865 ;
        RECT 72.710 129.695 72.880 130.475 ;
        RECT 73.685 130.345 73.855 130.475 ;
        RECT 71.190 129.525 72.880 129.695 ;
        RECT 73.050 129.915 73.515 130.305 ;
        RECT 73.685 130.175 74.080 130.345 ;
        RECT 71.190 129.345 71.360 129.525 ;
        RECT 67.990 128.635 69.060 128.805 ;
        RECT 69.230 128.425 69.420 128.865 ;
        RECT 69.590 128.595 70.540 128.875 ;
        RECT 70.850 128.785 71.110 129.175 ;
        RECT 71.530 129.105 72.320 129.355 ;
        RECT 70.760 128.615 71.110 128.785 ;
        RECT 71.320 128.425 71.650 128.885 ;
        RECT 72.525 128.815 72.695 129.525 ;
        RECT 73.050 129.325 73.220 129.915 ;
        RECT 72.865 129.105 73.220 129.325 ;
        RECT 73.390 129.105 73.740 129.725 ;
        RECT 73.910 128.815 74.080 130.175 ;
        RECT 74.445 130.005 74.770 130.790 ;
        RECT 74.250 128.955 74.710 130.005 ;
        RECT 72.525 128.645 73.380 128.815 ;
        RECT 73.585 128.645 74.080 128.815 ;
        RECT 74.250 128.425 74.580 128.785 ;
        RECT 74.940 128.685 75.110 130.805 ;
        RECT 75.280 130.475 75.610 130.975 ;
        RECT 75.780 130.305 76.035 130.805 ;
        RECT 75.285 130.135 76.035 130.305 ;
        RECT 75.285 129.145 75.515 130.135 ;
        RECT 77.045 129.995 77.300 130.665 ;
        RECT 77.480 130.175 77.765 130.975 ;
        RECT 77.945 130.255 78.275 130.765 ;
        RECT 75.685 129.315 76.035 129.965 ;
        RECT 75.285 128.975 76.035 129.145 ;
        RECT 75.280 128.425 75.610 128.805 ;
        RECT 75.780 128.685 76.035 128.975 ;
        RECT 77.045 129.135 77.225 129.995 ;
        RECT 77.945 129.665 78.195 130.255 ;
        RECT 78.545 130.105 78.715 130.715 ;
        RECT 78.885 130.285 79.215 130.975 ;
        RECT 79.445 130.425 79.685 130.715 ;
        RECT 79.885 130.595 80.305 130.975 ;
        RECT 80.485 130.505 81.115 130.755 ;
        RECT 81.585 130.595 81.915 130.975 ;
        RECT 80.485 130.425 80.655 130.505 ;
        RECT 82.085 130.425 82.255 130.715 ;
        RECT 82.435 130.595 82.815 130.975 ;
        RECT 83.055 130.590 83.885 130.760 ;
        RECT 79.445 130.255 80.655 130.425 ;
        RECT 77.395 129.335 78.195 129.665 ;
        RECT 77.045 128.935 77.300 129.135 ;
        RECT 76.960 128.765 77.300 128.935 ;
        RECT 77.045 128.605 77.300 128.765 ;
        RECT 77.480 128.425 77.765 128.885 ;
        RECT 77.945 128.685 78.195 129.335 ;
        RECT 78.395 130.085 78.715 130.105 ;
        RECT 78.395 129.915 80.315 130.085 ;
        RECT 78.395 129.020 78.585 129.915 ;
        RECT 80.485 129.745 80.655 130.255 ;
        RECT 80.825 129.995 81.345 130.305 ;
        RECT 78.755 129.575 80.655 129.745 ;
        RECT 78.755 129.515 79.085 129.575 ;
        RECT 79.235 129.345 79.565 129.405 ;
        RECT 78.905 129.075 79.565 129.345 ;
        RECT 78.395 128.690 78.715 129.020 ;
        RECT 78.895 128.425 79.555 128.905 ;
        RECT 79.755 128.815 79.925 129.575 ;
        RECT 80.825 129.405 81.005 129.815 ;
        RECT 80.095 129.235 80.425 129.355 ;
        RECT 81.175 129.235 81.345 129.995 ;
        RECT 80.095 129.065 81.345 129.235 ;
        RECT 81.515 130.175 82.885 130.425 ;
        RECT 81.515 129.405 81.705 130.175 ;
        RECT 82.635 129.915 82.885 130.175 ;
        RECT 81.875 129.745 82.125 129.905 ;
        RECT 83.055 129.745 83.225 130.590 ;
        RECT 84.120 130.305 84.290 130.805 ;
        RECT 84.460 130.475 84.790 130.975 ;
        RECT 83.395 129.915 83.895 130.295 ;
        RECT 84.120 130.135 84.815 130.305 ;
        RECT 81.875 129.575 83.225 129.745 ;
        RECT 82.805 129.535 83.225 129.575 ;
        RECT 81.515 129.065 81.935 129.405 ;
        RECT 82.225 129.075 82.635 129.405 ;
        RECT 79.755 128.645 80.605 128.815 ;
        RECT 81.165 128.425 81.485 128.885 ;
        RECT 81.685 128.635 81.935 129.065 ;
        RECT 82.225 128.425 82.635 128.865 ;
        RECT 82.805 128.805 82.975 129.535 ;
        RECT 83.145 128.985 83.495 129.355 ;
        RECT 83.675 129.045 83.895 129.915 ;
        RECT 84.065 129.345 84.475 129.965 ;
        RECT 84.645 129.165 84.815 130.135 ;
        RECT 84.120 128.975 84.815 129.165 ;
        RECT 82.805 128.605 83.820 128.805 ;
        RECT 84.120 128.645 84.290 128.975 ;
        RECT 84.460 128.425 84.790 128.805 ;
        RECT 85.005 128.685 85.230 130.805 ;
        RECT 85.400 130.475 85.730 130.975 ;
        RECT 85.900 130.305 86.070 130.805 ;
        RECT 85.405 130.135 86.070 130.305 ;
        RECT 85.405 129.145 85.635 130.135 ;
        RECT 85.805 129.315 86.155 129.965 ;
        RECT 86.330 129.810 86.620 130.975 ;
        RECT 87.960 130.245 88.255 130.975 ;
        RECT 88.425 130.075 88.685 130.800 ;
        RECT 88.855 130.245 89.115 130.975 ;
        RECT 89.285 130.075 89.545 130.800 ;
        RECT 89.715 130.245 89.975 130.975 ;
        RECT 90.145 130.075 90.405 130.800 ;
        RECT 90.575 130.245 90.835 130.975 ;
        RECT 91.005 130.075 91.265 130.800 ;
        RECT 87.955 129.835 91.265 130.075 ;
        RECT 91.435 129.865 91.695 130.975 ;
        RECT 87.955 129.245 88.925 129.835 ;
        RECT 91.865 129.665 92.115 130.800 ;
        RECT 92.295 129.865 92.590 130.975 ;
        RECT 92.810 129.835 93.040 130.975 ;
        RECT 93.210 129.825 93.540 130.805 ;
        RECT 93.710 129.835 93.920 130.975 ;
        RECT 89.095 129.415 92.115 129.665 ;
        RECT 85.405 128.975 86.070 129.145 ;
        RECT 85.400 128.425 85.730 128.805 ;
        RECT 85.900 128.685 86.070 128.975 ;
        RECT 86.330 128.425 86.620 129.150 ;
        RECT 87.955 129.075 91.265 129.245 ;
        RECT 87.955 128.425 88.255 128.905 ;
        RECT 88.425 128.620 88.685 129.075 ;
        RECT 88.855 128.425 89.115 128.905 ;
        RECT 89.285 128.620 89.545 129.075 ;
        RECT 89.715 128.425 89.975 128.905 ;
        RECT 90.145 128.620 90.405 129.075 ;
        RECT 90.575 128.425 90.835 128.905 ;
        RECT 91.005 128.620 91.265 129.075 ;
        RECT 91.435 128.425 91.695 128.950 ;
        RECT 91.865 128.605 92.115 129.415 ;
        RECT 92.285 129.055 92.600 129.665 ;
        RECT 92.790 129.415 93.120 129.665 ;
        RECT 92.295 128.425 92.540 128.885 ;
        RECT 92.810 128.425 93.040 129.245 ;
        RECT 93.290 129.225 93.540 129.825 ;
        RECT 95.075 129.785 95.330 130.665 ;
        RECT 95.500 129.835 95.805 130.975 ;
        RECT 96.145 130.595 96.475 130.975 ;
        RECT 96.655 130.425 96.825 130.715 ;
        RECT 96.995 130.515 97.245 130.975 ;
        RECT 96.025 130.255 96.825 130.425 ;
        RECT 97.415 130.465 98.285 130.805 ;
        RECT 93.210 128.595 93.540 129.225 ;
        RECT 93.710 128.425 93.920 129.245 ;
        RECT 95.075 129.135 95.285 129.785 ;
        RECT 96.025 129.665 96.195 130.255 ;
        RECT 97.415 130.085 97.585 130.465 ;
        RECT 98.520 130.345 98.690 130.805 ;
        RECT 98.860 130.515 99.230 130.975 ;
        RECT 99.525 130.375 99.695 130.715 ;
        RECT 99.865 130.545 100.195 130.975 ;
        RECT 100.430 130.375 100.600 130.715 ;
        RECT 96.365 129.915 97.585 130.085 ;
        RECT 97.755 130.005 98.215 130.295 ;
        RECT 98.520 130.175 99.080 130.345 ;
        RECT 99.525 130.205 100.600 130.375 ;
        RECT 100.770 130.475 101.450 130.805 ;
        RECT 101.665 130.475 101.915 130.805 ;
        RECT 102.085 130.515 102.335 130.975 ;
        RECT 98.910 130.035 99.080 130.175 ;
        RECT 97.755 129.995 98.720 130.005 ;
        RECT 97.415 129.825 97.585 129.915 ;
        RECT 98.045 129.835 98.720 129.995 ;
        RECT 95.455 129.635 96.195 129.665 ;
        RECT 95.455 129.335 96.370 129.635 ;
        RECT 96.045 129.160 96.370 129.335 ;
        RECT 95.075 128.605 95.330 129.135 ;
        RECT 95.500 128.425 95.805 128.885 ;
        RECT 96.050 128.805 96.370 129.160 ;
        RECT 96.540 129.375 97.080 129.745 ;
        RECT 97.415 129.655 97.820 129.825 ;
        RECT 96.540 128.975 96.780 129.375 ;
        RECT 97.260 129.205 97.480 129.485 ;
        RECT 96.950 129.035 97.480 129.205 ;
        RECT 96.950 128.805 97.120 129.035 ;
        RECT 97.650 128.875 97.820 129.655 ;
        RECT 97.990 129.045 98.340 129.665 ;
        RECT 98.510 129.045 98.720 129.835 ;
        RECT 98.910 129.865 100.410 130.035 ;
        RECT 98.910 129.175 99.080 129.865 ;
        RECT 100.770 129.695 100.940 130.475 ;
        RECT 101.745 130.345 101.915 130.475 ;
        RECT 99.250 129.525 100.940 129.695 ;
        RECT 101.110 129.915 101.575 130.305 ;
        RECT 101.745 130.175 102.140 130.345 ;
        RECT 99.250 129.345 99.420 129.525 ;
        RECT 96.050 128.635 97.120 128.805 ;
        RECT 97.290 128.425 97.480 128.865 ;
        RECT 97.650 128.595 98.600 128.875 ;
        RECT 98.910 128.785 99.170 129.175 ;
        RECT 99.590 129.105 100.380 129.355 ;
        RECT 98.820 128.615 99.170 128.785 ;
        RECT 99.380 128.425 99.710 128.885 ;
        RECT 100.585 128.815 100.755 129.525 ;
        RECT 101.110 129.325 101.280 129.915 ;
        RECT 100.925 129.105 101.280 129.325 ;
        RECT 101.450 129.105 101.800 129.725 ;
        RECT 101.970 128.815 102.140 130.175 ;
        RECT 102.505 130.005 102.830 130.790 ;
        RECT 102.310 128.955 102.770 130.005 ;
        RECT 100.585 128.645 101.440 128.815 ;
        RECT 101.645 128.645 102.140 128.815 ;
        RECT 102.310 128.425 102.640 128.785 ;
        RECT 103.000 128.685 103.170 130.805 ;
        RECT 103.340 130.475 103.670 130.975 ;
        RECT 103.840 130.305 104.095 130.805 ;
        RECT 103.345 130.135 104.095 130.305 ;
        RECT 103.345 129.145 103.575 130.135 ;
        RECT 103.745 129.315 104.095 129.965 ;
        RECT 104.270 129.885 105.480 130.975 ;
        RECT 104.270 129.345 104.790 129.885 ;
        RECT 105.690 129.835 105.920 130.975 ;
        RECT 106.090 129.825 106.420 130.805 ;
        RECT 106.590 129.835 106.800 130.975 ;
        RECT 107.490 129.885 111.000 130.975 ;
        RECT 111.170 129.885 112.380 130.975 ;
        RECT 104.960 129.175 105.480 129.715 ;
        RECT 105.670 129.415 106.000 129.665 ;
        RECT 103.345 128.975 104.095 129.145 ;
        RECT 103.340 128.425 103.670 128.805 ;
        RECT 103.840 128.685 104.095 128.975 ;
        RECT 104.270 128.425 105.480 129.175 ;
        RECT 105.690 128.425 105.920 129.245 ;
        RECT 106.170 129.225 106.420 129.825 ;
        RECT 107.490 129.365 109.180 129.885 ;
        RECT 106.090 128.595 106.420 129.225 ;
        RECT 106.590 128.425 106.800 129.245 ;
        RECT 109.350 129.195 111.000 129.715 ;
        RECT 111.170 129.345 111.690 129.885 ;
        RECT 107.490 128.425 111.000 129.195 ;
        RECT 111.860 129.175 112.380 129.715 ;
        RECT 111.170 128.425 112.380 129.175 ;
        RECT 18.165 128.255 112.465 128.425 ;
        RECT 18.250 127.505 19.460 128.255 ;
        RECT 18.250 126.965 18.770 127.505 ;
        RECT 20.610 127.435 20.820 128.255 ;
        RECT 20.990 127.455 21.320 128.085 ;
        RECT 18.940 126.795 19.460 127.335 ;
        RECT 20.990 126.855 21.240 127.455 ;
        RECT 21.490 127.435 21.720 128.255 ;
        RECT 21.930 127.530 22.220 128.255 ;
        RECT 22.700 127.785 22.870 128.255 ;
        RECT 23.040 127.605 23.370 128.085 ;
        RECT 23.540 127.785 23.710 128.255 ;
        RECT 23.880 127.605 24.210 128.085 ;
        RECT 22.445 127.435 24.210 127.605 ;
        RECT 24.380 127.445 24.550 128.255 ;
        RECT 24.750 127.875 25.820 128.045 ;
        RECT 24.750 127.520 25.070 127.875 ;
        RECT 21.410 127.015 21.740 127.265 ;
        RECT 22.445 126.885 22.855 127.435 ;
        RECT 24.745 127.265 25.070 127.520 ;
        RECT 23.040 127.055 25.070 127.265 ;
        RECT 24.725 127.045 25.070 127.055 ;
        RECT 25.240 127.305 25.480 127.705 ;
        RECT 25.650 127.645 25.820 127.875 ;
        RECT 25.990 127.815 26.180 128.255 ;
        RECT 26.350 127.805 27.300 128.085 ;
        RECT 27.520 127.895 27.870 128.065 ;
        RECT 25.650 127.475 26.180 127.645 ;
        RECT 18.250 125.705 19.460 126.795 ;
        RECT 20.610 125.705 20.820 126.845 ;
        RECT 20.990 125.875 21.320 126.855 ;
        RECT 21.490 125.705 21.720 126.845 ;
        RECT 21.930 125.705 22.220 126.870 ;
        RECT 22.445 126.715 24.170 126.885 ;
        RECT 22.700 125.705 22.870 126.545 ;
        RECT 23.080 125.875 23.330 126.715 ;
        RECT 23.540 125.705 23.710 126.545 ;
        RECT 23.880 125.875 24.170 126.715 ;
        RECT 24.380 125.705 24.550 126.765 ;
        RECT 24.725 126.425 24.895 127.045 ;
        RECT 25.240 126.935 25.780 127.305 ;
        RECT 25.960 127.195 26.180 127.475 ;
        RECT 26.350 127.025 26.520 127.805 ;
        RECT 26.115 126.855 26.520 127.025 ;
        RECT 26.690 127.015 27.040 127.635 ;
        RECT 26.115 126.765 26.285 126.855 ;
        RECT 27.210 126.845 27.420 127.635 ;
        RECT 25.065 126.595 26.285 126.765 ;
        RECT 26.745 126.685 27.420 126.845 ;
        RECT 24.725 126.255 25.525 126.425 ;
        RECT 24.845 125.705 25.175 126.085 ;
        RECT 25.355 125.965 25.525 126.255 ;
        RECT 26.115 126.215 26.285 126.595 ;
        RECT 26.455 126.675 27.420 126.685 ;
        RECT 27.610 127.505 27.870 127.895 ;
        RECT 28.080 127.795 28.410 128.255 ;
        RECT 29.285 127.865 30.140 128.035 ;
        RECT 30.345 127.865 30.840 128.035 ;
        RECT 31.010 127.895 31.340 128.255 ;
        RECT 27.610 126.815 27.780 127.505 ;
        RECT 27.950 127.155 28.120 127.335 ;
        RECT 28.290 127.325 29.080 127.575 ;
        RECT 29.285 127.155 29.455 127.865 ;
        RECT 29.625 127.355 29.980 127.575 ;
        RECT 27.950 126.985 29.640 127.155 ;
        RECT 26.455 126.385 26.915 126.675 ;
        RECT 27.610 126.645 29.110 126.815 ;
        RECT 27.610 126.505 27.780 126.645 ;
        RECT 27.220 126.335 27.780 126.505 ;
        RECT 25.695 125.705 25.945 126.165 ;
        RECT 26.115 125.875 26.985 126.215 ;
        RECT 27.220 125.875 27.390 126.335 ;
        RECT 28.225 126.305 29.300 126.475 ;
        RECT 27.560 125.705 27.930 126.165 ;
        RECT 28.225 125.965 28.395 126.305 ;
        RECT 28.565 125.705 28.895 126.135 ;
        RECT 29.130 125.965 29.300 126.305 ;
        RECT 29.470 126.205 29.640 126.985 ;
        RECT 29.810 126.765 29.980 127.355 ;
        RECT 30.150 126.955 30.500 127.575 ;
        RECT 29.810 126.375 30.275 126.765 ;
        RECT 30.670 126.505 30.840 127.865 ;
        RECT 31.010 126.675 31.470 127.725 ;
        RECT 30.445 126.335 30.840 126.505 ;
        RECT 30.445 126.205 30.615 126.335 ;
        RECT 29.470 125.875 30.150 126.205 ;
        RECT 30.365 125.875 30.615 126.205 ;
        RECT 30.785 125.705 31.035 126.165 ;
        RECT 31.205 125.890 31.530 126.675 ;
        RECT 31.700 125.875 31.870 127.995 ;
        RECT 32.040 127.875 32.370 128.255 ;
        RECT 32.540 127.705 32.795 127.995 ;
        RECT 32.045 127.535 32.795 127.705 ;
        RECT 33.980 127.705 34.150 128.085 ;
        RECT 34.330 127.875 34.660 128.255 ;
        RECT 33.980 127.535 34.645 127.705 ;
        RECT 34.840 127.580 35.100 128.085 ;
        RECT 32.045 126.545 32.275 127.535 ;
        RECT 32.445 126.715 32.795 127.365 ;
        RECT 33.910 126.985 34.250 127.355 ;
        RECT 34.475 127.280 34.645 127.535 ;
        RECT 34.475 126.950 34.750 127.280 ;
        RECT 34.475 126.805 34.645 126.950 ;
        RECT 33.970 126.635 34.645 126.805 ;
        RECT 34.920 126.780 35.100 127.580 ;
        RECT 32.045 126.375 32.795 126.545 ;
        RECT 32.040 125.705 32.370 126.205 ;
        RECT 32.540 125.875 32.795 126.375 ;
        RECT 33.970 125.875 34.150 126.635 ;
        RECT 34.330 125.705 34.660 126.465 ;
        RECT 34.830 125.875 35.100 126.780 ;
        RECT 35.270 127.455 35.610 128.085 ;
        RECT 35.780 127.455 36.030 128.255 ;
        RECT 36.220 127.605 36.550 128.085 ;
        RECT 36.720 127.795 36.945 128.255 ;
        RECT 37.115 127.605 37.445 128.085 ;
        RECT 35.270 126.845 35.445 127.455 ;
        RECT 36.220 127.435 37.445 127.605 ;
        RECT 38.075 127.475 38.575 128.085 ;
        RECT 35.615 127.095 36.310 127.265 ;
        RECT 36.140 126.845 36.310 127.095 ;
        RECT 36.485 127.065 36.905 127.265 ;
        RECT 37.075 127.065 37.405 127.265 ;
        RECT 37.575 127.065 37.905 127.265 ;
        RECT 38.075 126.845 38.245 127.475 ;
        RECT 39.870 127.455 40.210 128.085 ;
        RECT 40.380 127.455 40.630 128.255 ;
        RECT 40.820 127.605 41.150 128.085 ;
        RECT 41.320 127.795 41.545 128.255 ;
        RECT 41.715 127.605 42.045 128.085 ;
        RECT 39.870 127.405 40.100 127.455 ;
        RECT 40.820 127.435 42.045 127.605 ;
        RECT 42.675 127.475 43.175 128.085 ;
        RECT 38.430 127.015 38.780 127.265 ;
        RECT 39.870 126.845 40.045 127.405 ;
        RECT 40.215 127.095 40.910 127.265 ;
        RECT 40.740 126.845 40.910 127.095 ;
        RECT 41.085 127.065 41.505 127.265 ;
        RECT 41.675 127.065 42.005 127.265 ;
        RECT 42.175 127.065 42.505 127.265 ;
        RECT 42.675 126.845 42.845 127.475 ;
        RECT 43.825 127.445 44.070 128.050 ;
        RECT 44.290 127.720 44.800 128.255 ;
        RECT 43.550 127.275 44.780 127.445 ;
        RECT 43.030 127.015 43.380 127.265 ;
        RECT 35.270 125.875 35.610 126.845 ;
        RECT 35.780 125.705 35.950 126.845 ;
        RECT 36.140 126.675 38.575 126.845 ;
        RECT 36.220 125.705 36.470 126.505 ;
        RECT 37.115 125.875 37.445 126.675 ;
        RECT 37.745 125.705 38.075 126.505 ;
        RECT 38.245 125.875 38.575 126.675 ;
        RECT 39.870 125.875 40.210 126.845 ;
        RECT 40.380 125.705 40.550 126.845 ;
        RECT 40.740 126.675 43.175 126.845 ;
        RECT 40.820 125.705 41.070 126.505 ;
        RECT 41.715 125.875 42.045 126.675 ;
        RECT 42.345 125.705 42.675 126.505 ;
        RECT 42.845 125.875 43.175 126.675 ;
        RECT 43.550 126.465 43.890 127.275 ;
        RECT 44.060 126.710 44.810 126.900 ;
        RECT 43.550 126.055 44.065 126.465 ;
        RECT 44.300 125.705 44.470 126.465 ;
        RECT 44.640 126.045 44.810 126.710 ;
        RECT 44.980 126.725 45.170 128.085 ;
        RECT 45.340 127.575 45.615 128.085 ;
        RECT 45.805 127.720 46.335 128.085 ;
        RECT 46.760 127.855 47.090 128.255 ;
        RECT 46.160 127.685 46.335 127.720 ;
        RECT 45.340 127.405 45.620 127.575 ;
        RECT 45.340 126.925 45.615 127.405 ;
        RECT 45.820 126.725 45.990 127.525 ;
        RECT 44.980 126.555 45.990 126.725 ;
        RECT 46.160 127.515 47.090 127.685 ;
        RECT 47.260 127.515 47.515 128.085 ;
        RECT 47.690 127.530 47.980 128.255 ;
        RECT 48.195 127.795 48.460 128.255 ;
        RECT 48.630 127.615 48.960 128.085 ;
        RECT 49.130 127.795 49.300 128.255 ;
        RECT 49.470 127.615 49.800 128.085 ;
        RECT 49.970 127.790 50.220 128.255 ;
        RECT 46.160 126.385 46.330 127.515 ;
        RECT 46.920 127.345 47.090 127.515 ;
        RECT 45.205 126.215 46.330 126.385 ;
        RECT 46.500 127.015 46.695 127.345 ;
        RECT 46.920 127.015 47.175 127.345 ;
        RECT 46.500 126.045 46.670 127.015 ;
        RECT 47.345 126.845 47.515 127.515 ;
        RECT 48.630 127.435 50.235 127.615 ;
        RECT 51.410 127.435 51.640 128.255 ;
        RECT 51.810 127.455 52.140 128.085 ;
        RECT 48.170 127.015 49.800 127.265 ;
        RECT 44.640 125.875 46.670 126.045 ;
        RECT 46.840 125.705 47.010 126.845 ;
        RECT 47.180 125.875 47.515 126.845 ;
        RECT 47.690 125.705 47.980 126.870 ;
        RECT 49.970 126.845 50.235 127.435 ;
        RECT 51.390 127.015 51.720 127.265 ;
        RECT 51.890 126.855 52.140 127.455 ;
        RECT 52.310 127.435 52.520 128.255 ;
        RECT 53.025 127.445 53.270 128.050 ;
        RECT 53.490 127.720 54.000 128.255 ;
        RECT 48.195 125.705 48.460 126.845 ;
        RECT 48.630 126.675 50.235 126.845 ;
        RECT 48.630 125.875 48.960 126.675 ;
        RECT 49.470 126.655 50.235 126.675 ;
        RECT 49.130 125.705 49.300 126.505 ;
        RECT 49.470 125.875 49.800 126.655 ;
        RECT 49.970 125.705 50.180 126.165 ;
        RECT 51.410 125.705 51.640 126.845 ;
        RECT 51.810 125.875 52.140 126.855 ;
        RECT 52.750 127.275 53.980 127.445 ;
        RECT 52.310 125.705 52.520 126.845 ;
        RECT 52.750 126.465 53.090 127.275 ;
        RECT 53.260 126.710 54.010 126.900 ;
        RECT 52.750 126.055 53.265 126.465 ;
        RECT 53.500 125.705 53.670 126.465 ;
        RECT 53.840 126.045 54.010 126.710 ;
        RECT 54.180 126.725 54.370 128.085 ;
        RECT 54.540 127.235 54.815 128.085 ;
        RECT 55.005 127.720 55.535 128.085 ;
        RECT 55.960 127.855 56.290 128.255 ;
        RECT 55.360 127.685 55.535 127.720 ;
        RECT 54.540 127.065 54.820 127.235 ;
        RECT 54.540 126.925 54.815 127.065 ;
        RECT 55.020 126.725 55.190 127.525 ;
        RECT 54.180 126.555 55.190 126.725 ;
        RECT 55.360 127.515 56.290 127.685 ;
        RECT 56.460 127.515 56.715 128.085 ;
        RECT 55.360 126.385 55.530 127.515 ;
        RECT 56.120 127.345 56.290 127.515 ;
        RECT 54.405 126.215 55.530 126.385 ;
        RECT 55.700 127.015 55.895 127.345 ;
        RECT 56.120 127.015 56.375 127.345 ;
        RECT 55.700 126.045 55.870 127.015 ;
        RECT 56.545 126.845 56.715 127.515 ;
        RECT 57.265 127.545 57.520 128.075 ;
        RECT 57.700 127.795 57.985 128.255 ;
        RECT 57.265 126.895 57.445 127.545 ;
        RECT 58.165 127.345 58.415 127.995 ;
        RECT 57.615 127.015 58.415 127.345 ;
        RECT 53.840 125.875 55.870 126.045 ;
        RECT 56.040 125.705 56.210 126.845 ;
        RECT 56.380 125.875 56.715 126.845 ;
        RECT 57.180 126.725 57.445 126.895 ;
        RECT 57.265 126.685 57.445 126.725 ;
        RECT 57.265 126.015 57.520 126.685 ;
        RECT 57.700 125.705 57.985 126.505 ;
        RECT 58.165 126.425 58.415 127.015 ;
        RECT 58.615 127.660 58.935 127.990 ;
        RECT 59.115 127.775 59.775 128.255 ;
        RECT 59.975 127.865 60.825 128.035 ;
        RECT 58.615 126.765 58.805 127.660 ;
        RECT 59.125 127.335 59.785 127.605 ;
        RECT 59.455 127.275 59.785 127.335 ;
        RECT 58.975 127.105 59.305 127.165 ;
        RECT 59.975 127.105 60.145 127.865 ;
        RECT 61.385 127.795 61.705 128.255 ;
        RECT 61.905 127.615 62.155 128.045 ;
        RECT 62.445 127.815 62.855 128.255 ;
        RECT 63.025 127.875 64.040 128.075 ;
        RECT 60.315 127.445 61.565 127.615 ;
        RECT 60.315 127.325 60.645 127.445 ;
        RECT 58.975 126.935 60.875 127.105 ;
        RECT 58.615 126.595 60.535 126.765 ;
        RECT 58.615 126.575 58.935 126.595 ;
        RECT 58.165 125.915 58.495 126.425 ;
        RECT 58.765 125.965 58.935 126.575 ;
        RECT 60.705 126.425 60.875 126.935 ;
        RECT 61.045 126.865 61.225 127.275 ;
        RECT 61.395 126.685 61.565 127.445 ;
        RECT 59.105 125.705 59.435 126.395 ;
        RECT 59.665 126.255 60.875 126.425 ;
        RECT 61.045 126.375 61.565 126.685 ;
        RECT 61.735 127.275 62.155 127.615 ;
        RECT 62.445 127.275 62.855 127.605 ;
        RECT 61.735 126.505 61.925 127.275 ;
        RECT 63.025 127.145 63.195 127.875 ;
        RECT 64.340 127.705 64.510 128.035 ;
        RECT 64.680 127.875 65.010 128.255 ;
        RECT 63.365 127.325 63.715 127.695 ;
        RECT 63.025 127.105 63.445 127.145 ;
        RECT 62.095 126.935 63.445 127.105 ;
        RECT 62.095 126.775 62.345 126.935 ;
        RECT 62.855 126.505 63.105 126.765 ;
        RECT 61.735 126.255 63.105 126.505 ;
        RECT 59.665 125.965 59.905 126.255 ;
        RECT 60.705 126.175 60.875 126.255 ;
        RECT 60.105 125.705 60.525 126.085 ;
        RECT 60.705 125.925 61.335 126.175 ;
        RECT 61.805 125.705 62.135 126.085 ;
        RECT 62.305 125.965 62.475 126.255 ;
        RECT 63.275 126.090 63.445 126.935 ;
        RECT 63.895 126.765 64.115 127.635 ;
        RECT 64.340 127.515 65.035 127.705 ;
        RECT 63.615 126.385 64.115 126.765 ;
        RECT 64.285 126.715 64.695 127.335 ;
        RECT 64.865 126.545 65.035 127.515 ;
        RECT 64.340 126.375 65.035 126.545 ;
        RECT 62.655 125.705 63.035 126.085 ;
        RECT 63.275 125.920 64.105 126.090 ;
        RECT 64.340 125.875 64.510 126.375 ;
        RECT 64.680 125.705 65.010 126.205 ;
        RECT 65.225 125.875 65.450 127.995 ;
        RECT 65.620 127.875 65.950 128.255 ;
        RECT 66.120 127.705 66.290 127.995 ;
        RECT 65.625 127.535 66.290 127.705 ;
        RECT 65.625 126.545 65.855 127.535 ;
        RECT 66.550 127.505 67.760 128.255 ;
        RECT 66.025 126.715 66.375 127.365 ;
        RECT 66.550 126.795 67.070 127.335 ;
        RECT 67.240 126.965 67.760 127.505 ;
        RECT 67.990 127.435 68.200 128.255 ;
        RECT 68.370 127.455 68.700 128.085 ;
        RECT 68.370 126.855 68.620 127.455 ;
        RECT 68.870 127.435 69.100 128.255 ;
        RECT 69.585 127.445 69.830 128.050 ;
        RECT 70.050 127.720 70.560 128.255 ;
        RECT 69.310 127.275 70.540 127.445 ;
        RECT 68.790 127.015 69.120 127.265 ;
        RECT 65.625 126.375 66.290 126.545 ;
        RECT 65.620 125.705 65.950 126.205 ;
        RECT 66.120 125.875 66.290 126.375 ;
        RECT 66.550 125.705 67.760 126.795 ;
        RECT 67.990 125.705 68.200 126.845 ;
        RECT 68.370 125.875 68.700 126.855 ;
        RECT 68.870 125.705 69.100 126.845 ;
        RECT 69.310 126.465 69.650 127.275 ;
        RECT 69.820 126.710 70.570 126.900 ;
        RECT 69.310 126.055 69.825 126.465 ;
        RECT 70.060 125.705 70.230 126.465 ;
        RECT 70.400 126.045 70.570 126.710 ;
        RECT 70.740 126.725 70.930 128.085 ;
        RECT 71.100 127.235 71.375 128.085 ;
        RECT 71.565 127.720 72.095 128.085 ;
        RECT 72.520 127.855 72.850 128.255 ;
        RECT 71.920 127.685 72.095 127.720 ;
        RECT 71.100 127.065 71.380 127.235 ;
        RECT 71.100 126.925 71.375 127.065 ;
        RECT 71.580 126.725 71.750 127.525 ;
        RECT 70.740 126.555 71.750 126.725 ;
        RECT 71.920 127.515 72.850 127.685 ;
        RECT 73.020 127.515 73.275 128.085 ;
        RECT 73.450 127.530 73.740 128.255 ;
        RECT 74.000 127.775 74.300 128.255 ;
        RECT 74.470 127.605 74.730 128.060 ;
        RECT 74.900 127.775 75.160 128.255 ;
        RECT 75.340 127.605 75.600 128.060 ;
        RECT 75.770 127.775 76.020 128.255 ;
        RECT 76.200 127.605 76.460 128.060 ;
        RECT 76.630 127.775 76.880 128.255 ;
        RECT 77.060 127.605 77.320 128.060 ;
        RECT 77.490 127.775 77.735 128.255 ;
        RECT 77.905 127.605 78.180 128.060 ;
        RECT 78.350 127.775 78.595 128.255 ;
        RECT 78.765 127.605 79.025 128.060 ;
        RECT 79.195 127.775 79.455 128.255 ;
        RECT 79.625 127.605 79.885 128.060 ;
        RECT 80.055 127.775 80.315 128.255 ;
        RECT 80.485 127.605 80.745 128.060 ;
        RECT 80.915 127.695 81.175 128.255 ;
        RECT 71.920 126.385 72.090 127.515 ;
        RECT 72.680 127.345 72.850 127.515 ;
        RECT 70.965 126.215 72.090 126.385 ;
        RECT 72.260 127.015 72.455 127.345 ;
        RECT 72.680 127.015 72.935 127.345 ;
        RECT 72.260 126.045 72.430 127.015 ;
        RECT 73.105 126.845 73.275 127.515 ;
        RECT 74.000 127.435 80.745 127.605 ;
        RECT 70.400 125.875 72.430 126.045 ;
        RECT 72.600 125.705 72.770 126.845 ;
        RECT 72.940 125.875 73.275 126.845 ;
        RECT 73.450 125.705 73.740 126.870 ;
        RECT 74.000 126.845 75.165 127.435 ;
        RECT 81.345 127.265 81.595 128.075 ;
        RECT 81.775 127.730 82.035 128.255 ;
        RECT 82.205 127.265 82.455 128.075 ;
        RECT 82.635 127.745 82.940 128.255 ;
        RECT 75.335 127.015 82.455 127.265 ;
        RECT 82.625 127.015 82.940 127.575 ;
        RECT 83.945 127.545 84.200 128.075 ;
        RECT 84.380 127.795 84.665 128.255 ;
        RECT 83.945 127.235 84.125 127.545 ;
        RECT 84.845 127.345 85.095 127.995 ;
        RECT 83.860 127.065 84.125 127.235 ;
        RECT 74.000 126.620 80.745 126.845 ;
        RECT 74.000 125.705 74.270 126.450 ;
        RECT 74.440 125.880 74.730 126.620 ;
        RECT 75.340 126.605 80.745 126.620 ;
        RECT 74.900 125.710 75.155 126.435 ;
        RECT 75.340 125.880 75.600 126.605 ;
        RECT 75.770 125.710 76.015 126.435 ;
        RECT 76.200 125.880 76.460 126.605 ;
        RECT 76.630 125.710 76.875 126.435 ;
        RECT 77.060 125.880 77.320 126.605 ;
        RECT 77.490 125.710 77.735 126.435 ;
        RECT 77.905 125.880 78.165 126.605 ;
        RECT 78.335 125.710 78.595 126.435 ;
        RECT 78.765 125.880 79.025 126.605 ;
        RECT 79.195 125.710 79.455 126.435 ;
        RECT 79.625 125.880 79.885 126.605 ;
        RECT 80.055 125.710 80.315 126.435 ;
        RECT 80.485 125.880 80.745 126.605 ;
        RECT 80.915 125.710 81.175 126.505 ;
        RECT 81.345 125.880 81.595 127.015 ;
        RECT 74.900 125.705 81.175 125.710 ;
        RECT 81.775 125.705 82.035 126.515 ;
        RECT 82.210 125.875 82.455 127.015 ;
        RECT 83.945 126.685 84.125 127.065 ;
        RECT 84.295 127.015 85.095 127.345 ;
        RECT 82.635 125.705 82.930 126.515 ;
        RECT 83.945 126.015 84.200 126.685 ;
        RECT 84.380 125.705 84.665 126.505 ;
        RECT 84.845 126.425 85.095 127.015 ;
        RECT 85.295 127.660 85.615 127.990 ;
        RECT 85.795 127.775 86.455 128.255 ;
        RECT 86.655 127.865 87.505 128.035 ;
        RECT 85.295 126.765 85.485 127.660 ;
        RECT 85.805 127.335 86.465 127.605 ;
        RECT 86.135 127.275 86.465 127.335 ;
        RECT 85.655 127.105 85.985 127.165 ;
        RECT 86.655 127.105 86.825 127.865 ;
        RECT 88.065 127.795 88.385 128.255 ;
        RECT 88.585 127.615 88.835 128.045 ;
        RECT 89.125 127.815 89.535 128.255 ;
        RECT 89.705 127.875 90.720 128.075 ;
        RECT 86.995 127.445 88.245 127.615 ;
        RECT 86.995 127.325 87.325 127.445 ;
        RECT 85.655 126.935 87.555 127.105 ;
        RECT 85.295 126.595 87.215 126.765 ;
        RECT 85.295 126.575 85.615 126.595 ;
        RECT 84.845 125.915 85.175 126.425 ;
        RECT 85.445 125.965 85.615 126.575 ;
        RECT 87.385 126.425 87.555 126.935 ;
        RECT 87.725 126.865 87.905 127.275 ;
        RECT 88.075 126.685 88.245 127.445 ;
        RECT 85.785 125.705 86.115 126.395 ;
        RECT 86.345 126.255 87.555 126.425 ;
        RECT 87.725 126.375 88.245 126.685 ;
        RECT 88.415 127.275 88.835 127.615 ;
        RECT 89.125 127.275 89.535 127.605 ;
        RECT 88.415 126.505 88.605 127.275 ;
        RECT 89.705 127.145 89.875 127.875 ;
        RECT 91.020 127.705 91.190 128.035 ;
        RECT 91.360 127.875 91.690 128.255 ;
        RECT 90.045 127.325 90.395 127.695 ;
        RECT 89.705 127.105 90.125 127.145 ;
        RECT 88.775 126.935 90.125 127.105 ;
        RECT 88.775 126.775 89.025 126.935 ;
        RECT 89.535 126.505 89.785 126.765 ;
        RECT 88.415 126.255 89.785 126.505 ;
        RECT 86.345 125.965 86.585 126.255 ;
        RECT 87.385 126.175 87.555 126.255 ;
        RECT 86.785 125.705 87.205 126.085 ;
        RECT 87.385 125.925 88.015 126.175 ;
        RECT 88.485 125.705 88.815 126.085 ;
        RECT 88.985 125.965 89.155 126.255 ;
        RECT 89.955 126.090 90.125 126.935 ;
        RECT 90.575 126.765 90.795 127.635 ;
        RECT 91.020 127.515 91.715 127.705 ;
        RECT 90.295 126.385 90.795 126.765 ;
        RECT 90.965 126.715 91.375 127.335 ;
        RECT 91.545 126.545 91.715 127.515 ;
        RECT 91.020 126.375 91.715 126.545 ;
        RECT 89.335 125.705 89.715 126.085 ;
        RECT 89.955 125.920 90.785 126.090 ;
        RECT 91.020 125.875 91.190 126.375 ;
        RECT 91.360 125.705 91.690 126.205 ;
        RECT 91.905 125.875 92.130 127.995 ;
        RECT 92.300 127.875 92.630 128.255 ;
        RECT 92.800 127.705 92.970 127.995 ;
        RECT 92.305 127.535 92.970 127.705 ;
        RECT 92.305 126.545 92.535 127.535 ;
        RECT 93.230 127.455 93.570 128.085 ;
        RECT 93.740 127.455 93.990 128.255 ;
        RECT 94.180 127.605 94.510 128.085 ;
        RECT 94.680 127.795 94.905 128.255 ;
        RECT 95.075 127.605 95.405 128.085 ;
        RECT 92.705 126.715 93.055 127.365 ;
        RECT 93.230 126.845 93.405 127.455 ;
        RECT 94.180 127.435 95.405 127.605 ;
        RECT 96.035 127.475 96.535 128.085 ;
        RECT 93.575 127.095 94.270 127.265 ;
        RECT 94.100 126.845 94.270 127.095 ;
        RECT 94.445 127.065 94.865 127.265 ;
        RECT 95.035 127.065 95.365 127.265 ;
        RECT 95.535 127.065 95.865 127.265 ;
        RECT 96.035 126.845 96.205 127.475 ;
        RECT 97.890 127.435 98.100 128.255 ;
        RECT 98.270 127.455 98.600 128.085 ;
        RECT 96.390 127.015 96.740 127.265 ;
        RECT 98.270 126.855 98.520 127.455 ;
        RECT 98.770 127.435 99.000 128.255 ;
        RECT 99.210 127.530 99.500 128.255 ;
        RECT 99.785 127.625 100.070 128.085 ;
        RECT 100.240 127.795 100.510 128.255 ;
        RECT 99.785 127.455 100.740 127.625 ;
        RECT 98.690 127.015 99.020 127.265 ;
        RECT 92.305 126.375 92.970 126.545 ;
        RECT 92.300 125.705 92.630 126.205 ;
        RECT 92.800 125.875 92.970 126.375 ;
        RECT 93.230 125.875 93.570 126.845 ;
        RECT 93.740 125.705 93.910 126.845 ;
        RECT 94.100 126.675 96.535 126.845 ;
        RECT 94.180 125.705 94.430 126.505 ;
        RECT 95.075 125.875 95.405 126.675 ;
        RECT 95.705 125.705 96.035 126.505 ;
        RECT 96.205 125.875 96.535 126.675 ;
        RECT 97.890 125.705 98.100 126.845 ;
        RECT 98.270 125.875 98.600 126.855 ;
        RECT 98.770 125.705 99.000 126.845 ;
        RECT 99.210 125.705 99.500 126.870 ;
        RECT 99.670 126.725 100.360 127.285 ;
        RECT 100.530 126.555 100.740 127.455 ;
        RECT 99.785 126.335 100.740 126.555 ;
        RECT 100.910 127.285 101.310 128.085 ;
        RECT 101.500 127.625 101.780 128.085 ;
        RECT 102.300 127.795 102.625 128.255 ;
        RECT 101.500 127.455 102.625 127.625 ;
        RECT 102.795 127.515 103.180 128.085 ;
        RECT 102.175 127.345 102.625 127.455 ;
        RECT 100.910 126.725 102.005 127.285 ;
        RECT 102.175 127.015 102.730 127.345 ;
        RECT 99.785 125.875 100.070 126.335 ;
        RECT 100.240 125.705 100.510 126.165 ;
        RECT 100.910 125.875 101.310 126.725 ;
        RECT 102.175 126.555 102.625 127.015 ;
        RECT 102.900 126.845 103.180 127.515 ;
        RECT 101.500 126.335 102.625 126.555 ;
        RECT 101.500 125.875 101.780 126.335 ;
        RECT 102.300 125.705 102.625 126.165 ;
        RECT 102.795 125.875 103.180 126.845 ;
        RECT 103.350 127.755 103.650 128.085 ;
        RECT 103.820 127.775 104.095 128.255 ;
        RECT 103.350 126.845 103.520 127.755 ;
        RECT 104.275 127.605 104.570 127.995 ;
        RECT 104.740 127.775 104.995 128.255 ;
        RECT 105.170 127.605 105.430 127.995 ;
        RECT 105.600 127.775 105.880 128.255 ;
        RECT 103.690 127.015 104.040 127.585 ;
        RECT 104.275 127.435 105.925 127.605 ;
        RECT 106.110 127.505 107.320 128.255 ;
        RECT 104.210 127.095 105.350 127.265 ;
        RECT 104.210 126.845 104.380 127.095 ;
        RECT 105.520 126.925 105.925 127.435 ;
        RECT 103.350 126.675 104.380 126.845 ;
        RECT 105.170 126.755 105.925 126.925 ;
        RECT 106.110 126.795 106.630 127.335 ;
        RECT 106.800 126.965 107.320 127.505 ;
        RECT 107.490 127.485 111.000 128.255 ;
        RECT 111.170 127.505 112.380 128.255 ;
        RECT 107.490 126.795 109.180 127.315 ;
        RECT 109.350 126.965 111.000 127.485 ;
        RECT 111.170 126.795 111.690 127.335 ;
        RECT 111.860 126.965 112.380 127.505 ;
        RECT 103.350 125.875 103.660 126.675 ;
        RECT 105.170 126.505 105.430 126.755 ;
        RECT 103.830 125.705 104.140 126.505 ;
        RECT 104.310 126.335 105.430 126.505 ;
        RECT 104.310 125.875 104.570 126.335 ;
        RECT 104.740 125.705 104.995 126.165 ;
        RECT 105.170 125.875 105.430 126.335 ;
        RECT 105.600 125.705 105.885 126.575 ;
        RECT 106.110 125.705 107.320 126.795 ;
        RECT 107.490 125.705 111.000 126.795 ;
        RECT 111.170 125.705 112.380 126.795 ;
        RECT 18.165 125.535 112.465 125.705 ;
        RECT 18.250 124.445 19.460 125.535 ;
        RECT 18.250 123.735 18.770 124.275 ;
        RECT 18.940 123.905 19.460 124.445 ;
        RECT 19.630 124.445 21.300 125.535 ;
        RECT 19.630 123.925 20.380 124.445 ;
        RECT 21.510 124.395 21.740 125.535 ;
        RECT 21.910 124.385 22.240 125.365 ;
        RECT 22.410 124.395 22.620 125.535 ;
        RECT 22.905 124.665 23.190 125.535 ;
        RECT 23.360 124.905 23.620 125.365 ;
        RECT 23.795 125.075 24.050 125.535 ;
        RECT 24.220 124.905 24.480 125.365 ;
        RECT 23.360 124.735 24.480 124.905 ;
        RECT 24.650 124.735 24.960 125.535 ;
        RECT 23.360 124.485 23.620 124.735 ;
        RECT 25.130 124.565 25.440 125.365 ;
        RECT 25.725 124.905 26.010 125.365 ;
        RECT 26.180 125.075 26.450 125.535 ;
        RECT 25.725 124.685 26.680 124.905 ;
        RECT 20.550 123.755 21.300 124.275 ;
        RECT 21.490 123.975 21.820 124.225 ;
        RECT 18.250 122.985 19.460 123.735 ;
        RECT 19.630 122.985 21.300 123.755 ;
        RECT 21.510 122.985 21.740 123.805 ;
        RECT 21.990 123.785 22.240 124.385 ;
        RECT 22.865 124.315 23.620 124.485 ;
        RECT 24.410 124.395 25.440 124.565 ;
        RECT 22.865 123.805 23.270 124.315 ;
        RECT 24.410 124.145 24.580 124.395 ;
        RECT 23.440 123.975 24.580 124.145 ;
        RECT 21.910 123.155 22.240 123.785 ;
        RECT 22.410 122.985 22.620 123.805 ;
        RECT 22.865 123.635 24.515 123.805 ;
        RECT 24.750 123.655 25.100 124.225 ;
        RECT 22.910 122.985 23.190 123.465 ;
        RECT 23.360 123.245 23.620 123.635 ;
        RECT 23.795 122.985 24.050 123.465 ;
        RECT 24.220 123.245 24.515 123.635 ;
        RECT 25.270 123.485 25.440 124.395 ;
        RECT 25.610 123.955 26.300 124.515 ;
        RECT 26.470 123.785 26.680 124.685 ;
        RECT 24.695 122.985 24.970 123.465 ;
        RECT 25.140 123.155 25.440 123.485 ;
        RECT 25.725 123.615 26.680 123.785 ;
        RECT 26.850 124.515 27.250 125.365 ;
        RECT 27.440 124.905 27.720 125.365 ;
        RECT 28.240 125.075 28.565 125.535 ;
        RECT 27.440 124.685 28.565 124.905 ;
        RECT 26.850 123.955 27.945 124.515 ;
        RECT 28.115 124.225 28.565 124.685 ;
        RECT 28.735 124.395 29.120 125.365 ;
        RECT 25.725 123.155 26.010 123.615 ;
        RECT 26.180 122.985 26.450 123.445 ;
        RECT 26.850 123.155 27.250 123.955 ;
        RECT 28.115 123.895 28.670 124.225 ;
        RECT 28.115 123.785 28.565 123.895 ;
        RECT 27.440 123.615 28.565 123.785 ;
        RECT 28.840 123.725 29.120 124.395 ;
        RECT 29.290 124.445 30.500 125.535 ;
        RECT 30.670 124.775 31.185 125.185 ;
        RECT 31.420 124.775 31.590 125.535 ;
        RECT 31.760 125.195 33.790 125.365 ;
        RECT 29.290 123.905 29.810 124.445 ;
        RECT 29.980 123.735 30.500 124.275 ;
        RECT 30.670 123.965 31.010 124.775 ;
        RECT 31.760 124.530 31.930 125.195 ;
        RECT 32.325 124.855 33.450 125.025 ;
        RECT 31.180 124.340 31.930 124.530 ;
        RECT 32.100 124.515 33.110 124.685 ;
        RECT 30.670 123.795 31.900 123.965 ;
        RECT 27.440 123.155 27.720 123.615 ;
        RECT 28.240 122.985 28.565 123.445 ;
        RECT 28.735 123.155 29.120 123.725 ;
        RECT 29.290 122.985 30.500 123.735 ;
        RECT 30.945 123.190 31.190 123.795 ;
        RECT 31.410 122.985 31.920 123.520 ;
        RECT 32.100 123.155 32.290 124.515 ;
        RECT 32.460 124.175 32.735 124.315 ;
        RECT 32.460 124.005 32.740 124.175 ;
        RECT 32.460 123.155 32.735 124.005 ;
        RECT 32.940 123.715 33.110 124.515 ;
        RECT 33.280 123.725 33.450 124.855 ;
        RECT 33.620 124.225 33.790 125.195 ;
        RECT 33.960 124.395 34.130 125.535 ;
        RECT 34.300 124.395 34.635 125.365 ;
        RECT 33.620 123.895 33.815 124.225 ;
        RECT 34.040 123.895 34.295 124.225 ;
        RECT 34.040 123.725 34.210 123.895 ;
        RECT 34.465 123.725 34.635 124.395 ;
        RECT 34.810 124.370 35.100 125.535 ;
        RECT 35.270 124.395 35.540 125.365 ;
        RECT 35.750 124.735 36.030 125.535 ;
        RECT 36.200 125.025 37.855 125.315 ;
        RECT 36.265 124.685 37.855 124.855 ;
        RECT 36.265 124.565 36.435 124.685 ;
        RECT 35.710 124.395 36.435 124.565 ;
        RECT 33.280 123.555 34.210 123.725 ;
        RECT 33.280 123.520 33.455 123.555 ;
        RECT 32.925 123.155 33.455 123.520 ;
        RECT 33.880 122.985 34.210 123.385 ;
        RECT 34.380 123.155 34.635 123.725 ;
        RECT 34.810 122.985 35.100 123.710 ;
        RECT 35.270 123.660 35.440 124.395 ;
        RECT 35.710 124.225 35.880 124.395 ;
        RECT 36.625 124.345 37.340 124.515 ;
        RECT 37.535 124.395 37.855 124.685 ;
        RECT 38.035 124.345 38.290 125.225 ;
        RECT 38.460 124.395 38.765 125.535 ;
        RECT 39.105 125.155 39.435 125.535 ;
        RECT 39.615 124.985 39.785 125.275 ;
        RECT 39.955 125.075 40.205 125.535 ;
        RECT 38.985 124.815 39.785 124.985 ;
        RECT 40.375 125.025 41.245 125.365 ;
        RECT 35.610 123.895 35.880 124.225 ;
        RECT 36.050 123.895 36.455 124.225 ;
        RECT 36.625 123.895 37.335 124.345 ;
        RECT 35.710 123.725 35.880 123.895 ;
        RECT 35.270 123.315 35.540 123.660 ;
        RECT 35.710 123.555 37.320 123.725 ;
        RECT 37.505 123.655 37.855 124.225 ;
        RECT 38.035 123.695 38.245 124.345 ;
        RECT 38.985 124.225 39.155 124.815 ;
        RECT 40.375 124.645 40.545 125.025 ;
        RECT 41.480 124.905 41.650 125.365 ;
        RECT 41.820 125.075 42.190 125.535 ;
        RECT 42.485 124.935 42.655 125.275 ;
        RECT 42.825 125.105 43.155 125.535 ;
        RECT 43.390 124.935 43.560 125.275 ;
        RECT 39.325 124.475 40.545 124.645 ;
        RECT 40.715 124.565 41.175 124.855 ;
        RECT 41.480 124.735 42.040 124.905 ;
        RECT 42.485 124.765 43.560 124.935 ;
        RECT 43.730 125.035 44.410 125.365 ;
        RECT 44.625 125.035 44.875 125.365 ;
        RECT 45.045 125.075 45.295 125.535 ;
        RECT 41.870 124.595 42.040 124.735 ;
        RECT 40.715 124.555 41.680 124.565 ;
        RECT 40.375 124.385 40.545 124.475 ;
        RECT 41.005 124.395 41.680 124.555 ;
        RECT 38.415 124.195 39.155 124.225 ;
        RECT 38.415 123.895 39.330 124.195 ;
        RECT 39.005 123.720 39.330 123.895 ;
        RECT 35.730 122.985 36.110 123.385 ;
        RECT 36.280 123.205 36.450 123.555 ;
        RECT 36.620 122.985 36.950 123.385 ;
        RECT 37.150 123.205 37.320 123.555 ;
        RECT 37.520 122.985 37.850 123.485 ;
        RECT 38.035 123.165 38.290 123.695 ;
        RECT 38.460 122.985 38.765 123.445 ;
        RECT 39.010 123.365 39.330 123.720 ;
        RECT 39.500 123.935 40.040 124.305 ;
        RECT 40.375 124.215 40.780 124.385 ;
        RECT 39.500 123.535 39.740 123.935 ;
        RECT 40.220 123.765 40.440 124.045 ;
        RECT 39.910 123.595 40.440 123.765 ;
        RECT 39.910 123.365 40.080 123.595 ;
        RECT 40.610 123.435 40.780 124.215 ;
        RECT 40.950 123.605 41.300 124.225 ;
        RECT 41.470 123.605 41.680 124.395 ;
        RECT 41.870 124.425 43.370 124.595 ;
        RECT 41.870 123.735 42.040 124.425 ;
        RECT 43.730 124.255 43.900 125.035 ;
        RECT 44.705 124.905 44.875 125.035 ;
        RECT 42.210 124.085 43.900 124.255 ;
        RECT 44.070 124.475 44.535 124.865 ;
        RECT 44.705 124.735 45.100 124.905 ;
        RECT 42.210 123.905 42.380 124.085 ;
        RECT 39.010 123.195 40.080 123.365 ;
        RECT 40.250 122.985 40.440 123.425 ;
        RECT 40.610 123.155 41.560 123.435 ;
        RECT 41.870 123.345 42.130 123.735 ;
        RECT 42.550 123.665 43.340 123.915 ;
        RECT 41.780 123.175 42.130 123.345 ;
        RECT 42.340 122.985 42.670 123.445 ;
        RECT 43.545 123.375 43.715 124.085 ;
        RECT 44.070 123.885 44.240 124.475 ;
        RECT 43.885 123.665 44.240 123.885 ;
        RECT 44.410 123.665 44.760 124.285 ;
        RECT 44.930 123.375 45.100 124.735 ;
        RECT 45.465 124.565 45.790 125.350 ;
        RECT 45.270 123.515 45.730 124.565 ;
        RECT 43.545 123.205 44.400 123.375 ;
        RECT 44.605 123.205 45.100 123.375 ;
        RECT 45.270 122.985 45.600 123.345 ;
        RECT 45.960 123.245 46.130 125.365 ;
        RECT 46.300 125.035 46.630 125.535 ;
        RECT 46.800 124.865 47.055 125.365 ;
        RECT 46.305 124.695 47.055 124.865 ;
        RECT 47.240 124.725 47.535 125.535 ;
        RECT 46.305 123.705 46.535 124.695 ;
        RECT 46.705 123.875 47.055 124.525 ;
        RECT 47.715 124.225 47.960 125.365 ;
        RECT 48.135 124.725 48.395 125.535 ;
        RECT 48.995 125.530 55.270 125.535 ;
        RECT 48.575 124.225 48.825 125.360 ;
        RECT 48.995 124.735 49.255 125.530 ;
        RECT 49.425 124.635 49.685 125.360 ;
        RECT 49.855 124.805 50.115 125.530 ;
        RECT 50.285 124.635 50.545 125.360 ;
        RECT 50.715 124.805 50.975 125.530 ;
        RECT 51.145 124.635 51.405 125.360 ;
        RECT 51.575 124.805 51.835 125.530 ;
        RECT 52.005 124.635 52.265 125.360 ;
        RECT 52.435 124.805 52.680 125.530 ;
        RECT 52.850 124.635 53.110 125.360 ;
        RECT 53.295 124.805 53.540 125.530 ;
        RECT 53.710 124.635 53.970 125.360 ;
        RECT 54.155 124.805 54.400 125.530 ;
        RECT 54.570 124.635 54.830 125.360 ;
        RECT 55.015 124.805 55.270 125.530 ;
        RECT 49.425 124.620 54.830 124.635 ;
        RECT 55.440 124.620 55.730 125.360 ;
        RECT 55.900 124.790 56.170 125.535 ;
        RECT 49.425 124.395 56.170 124.620 ;
        RECT 57.095 124.565 57.425 125.365 ;
        RECT 57.595 124.735 57.925 125.535 ;
        RECT 58.225 124.565 58.555 125.365 ;
        RECT 59.200 124.735 59.450 125.535 ;
        RECT 57.095 124.395 59.530 124.565 ;
        RECT 59.720 124.395 59.890 125.535 ;
        RECT 60.060 124.395 60.400 125.365 ;
        RECT 46.305 123.535 47.055 123.705 ;
        RECT 47.230 123.665 47.545 124.225 ;
        RECT 47.715 123.975 54.835 124.225 ;
        RECT 46.300 122.985 46.630 123.365 ;
        RECT 46.800 123.245 47.055 123.535 ;
        RECT 47.230 122.985 47.535 123.495 ;
        RECT 47.715 123.165 47.965 123.975 ;
        RECT 48.135 122.985 48.395 123.510 ;
        RECT 48.575 123.165 48.825 123.975 ;
        RECT 55.005 123.835 56.170 124.395 ;
        RECT 56.890 123.975 57.240 124.225 ;
        RECT 55.005 123.805 56.200 123.835 ;
        RECT 49.425 123.665 56.200 123.805 ;
        RECT 57.425 123.765 57.595 124.395 ;
        RECT 57.765 123.975 58.095 124.175 ;
        RECT 58.265 123.975 58.595 124.175 ;
        RECT 58.765 123.975 59.185 124.175 ;
        RECT 59.360 124.145 59.530 124.395 ;
        RECT 59.360 123.975 60.055 124.145 ;
        RECT 49.425 123.635 56.170 123.665 ;
        RECT 48.995 122.985 49.255 123.545 ;
        RECT 49.425 123.180 49.685 123.635 ;
        RECT 49.855 122.985 50.115 123.465 ;
        RECT 50.285 123.180 50.545 123.635 ;
        RECT 50.715 122.985 50.975 123.465 ;
        RECT 51.145 123.180 51.405 123.635 ;
        RECT 51.575 122.985 51.820 123.465 ;
        RECT 51.990 123.180 52.265 123.635 ;
        RECT 52.435 122.985 52.680 123.465 ;
        RECT 52.850 123.180 53.110 123.635 ;
        RECT 53.290 122.985 53.540 123.465 ;
        RECT 53.710 123.180 53.970 123.635 ;
        RECT 54.150 122.985 54.400 123.465 ;
        RECT 54.570 123.180 54.830 123.635 ;
        RECT 55.010 122.985 55.270 123.465 ;
        RECT 55.440 123.180 55.700 123.635 ;
        RECT 55.870 122.985 56.170 123.465 ;
        RECT 57.095 123.155 57.595 123.765 ;
        RECT 58.225 123.635 59.450 123.805 ;
        RECT 60.225 123.785 60.400 124.395 ;
        RECT 60.570 124.370 60.860 125.535 ;
        RECT 61.030 124.395 61.370 125.365 ;
        RECT 61.540 124.395 61.710 125.535 ;
        RECT 61.980 124.735 62.230 125.535 ;
        RECT 62.875 124.565 63.205 125.365 ;
        RECT 63.505 124.735 63.835 125.535 ;
        RECT 64.005 124.565 64.335 125.365 ;
        RECT 61.900 124.395 64.335 124.565 ;
        RECT 65.170 124.445 67.760 125.535 ;
        RECT 67.930 124.775 68.445 125.185 ;
        RECT 68.680 124.775 68.850 125.535 ;
        RECT 69.020 125.195 71.050 125.365 ;
        RECT 58.225 123.155 58.555 123.635 ;
        RECT 58.725 122.985 58.950 123.445 ;
        RECT 59.120 123.155 59.450 123.635 ;
        RECT 59.640 122.985 59.890 123.785 ;
        RECT 60.060 123.155 60.400 123.785 ;
        RECT 61.030 123.785 61.205 124.395 ;
        RECT 61.900 124.145 62.070 124.395 ;
        RECT 61.375 123.975 62.070 124.145 ;
        RECT 62.245 123.975 62.665 124.175 ;
        RECT 62.835 123.975 63.165 124.175 ;
        RECT 63.335 123.975 63.665 124.175 ;
        RECT 60.570 122.985 60.860 123.710 ;
        RECT 61.030 123.155 61.370 123.785 ;
        RECT 61.540 122.985 61.790 123.785 ;
        RECT 61.980 123.635 63.205 123.805 ;
        RECT 61.980 123.155 62.310 123.635 ;
        RECT 62.480 122.985 62.705 123.445 ;
        RECT 62.875 123.155 63.205 123.635 ;
        RECT 63.835 123.765 64.005 124.395 ;
        RECT 64.190 123.975 64.540 124.225 ;
        RECT 65.170 123.925 66.380 124.445 ;
        RECT 63.835 123.155 64.335 123.765 ;
        RECT 66.550 123.755 67.760 124.275 ;
        RECT 67.930 123.965 68.270 124.775 ;
        RECT 69.020 124.530 69.190 125.195 ;
        RECT 69.585 124.855 70.710 125.025 ;
        RECT 68.440 124.340 69.190 124.530 ;
        RECT 69.360 124.515 70.370 124.685 ;
        RECT 67.930 123.795 69.160 123.965 ;
        RECT 65.170 122.985 67.760 123.755 ;
        RECT 68.205 123.190 68.450 123.795 ;
        RECT 68.670 122.985 69.180 123.520 ;
        RECT 69.360 123.155 69.550 124.515 ;
        RECT 69.720 123.835 69.995 124.315 ;
        RECT 69.720 123.665 70.000 123.835 ;
        RECT 70.200 123.715 70.370 124.515 ;
        RECT 70.540 123.725 70.710 124.855 ;
        RECT 70.880 124.225 71.050 125.195 ;
        RECT 71.220 124.395 71.390 125.535 ;
        RECT 71.560 124.395 71.895 125.365 ;
        RECT 72.160 124.865 72.330 125.365 ;
        RECT 72.500 125.035 72.830 125.535 ;
        RECT 72.160 124.695 72.825 124.865 ;
        RECT 70.880 123.895 71.075 124.225 ;
        RECT 71.300 123.895 71.555 124.225 ;
        RECT 71.300 123.725 71.470 123.895 ;
        RECT 71.725 123.725 71.895 124.395 ;
        RECT 72.075 123.875 72.425 124.525 ;
        RECT 69.720 123.155 69.995 123.665 ;
        RECT 70.540 123.555 71.470 123.725 ;
        RECT 70.540 123.520 70.715 123.555 ;
        RECT 70.185 123.155 70.715 123.520 ;
        RECT 71.140 122.985 71.470 123.385 ;
        RECT 71.640 123.155 71.895 123.725 ;
        RECT 72.595 123.705 72.825 124.695 ;
        RECT 72.160 123.535 72.825 123.705 ;
        RECT 72.160 123.245 72.330 123.535 ;
        RECT 72.500 122.985 72.830 123.365 ;
        RECT 73.000 123.245 73.225 125.365 ;
        RECT 73.440 125.035 73.770 125.535 ;
        RECT 73.940 124.865 74.110 125.365 ;
        RECT 74.345 125.150 75.175 125.320 ;
        RECT 75.415 125.155 75.795 125.535 ;
        RECT 73.415 124.695 74.110 124.865 ;
        RECT 73.415 123.725 73.585 124.695 ;
        RECT 73.755 123.905 74.165 124.525 ;
        RECT 74.335 124.475 74.835 124.855 ;
        RECT 73.415 123.535 74.110 123.725 ;
        RECT 74.335 123.605 74.555 124.475 ;
        RECT 75.005 124.305 75.175 125.150 ;
        RECT 75.975 124.985 76.145 125.275 ;
        RECT 76.315 125.155 76.645 125.535 ;
        RECT 77.115 125.065 77.745 125.315 ;
        RECT 77.925 125.155 78.345 125.535 ;
        RECT 77.575 124.985 77.745 125.065 ;
        RECT 78.545 124.985 78.785 125.275 ;
        RECT 75.345 124.735 76.715 124.985 ;
        RECT 75.345 124.475 75.595 124.735 ;
        RECT 76.105 124.305 76.355 124.465 ;
        RECT 75.005 124.135 76.355 124.305 ;
        RECT 75.005 124.095 75.425 124.135 ;
        RECT 74.735 123.545 75.085 123.915 ;
        RECT 73.440 122.985 73.770 123.365 ;
        RECT 73.940 123.205 74.110 123.535 ;
        RECT 75.255 123.365 75.425 124.095 ;
        RECT 76.525 123.965 76.715 124.735 ;
        RECT 75.595 123.635 76.005 123.965 ;
        RECT 76.295 123.625 76.715 123.965 ;
        RECT 76.885 124.555 77.405 124.865 ;
        RECT 77.575 124.815 78.785 124.985 ;
        RECT 79.015 124.845 79.345 125.535 ;
        RECT 76.885 123.795 77.055 124.555 ;
        RECT 77.225 123.965 77.405 124.375 ;
        RECT 77.575 124.305 77.745 124.815 ;
        RECT 79.515 124.665 79.685 125.275 ;
        RECT 79.955 124.815 80.285 125.325 ;
        RECT 79.515 124.645 79.835 124.665 ;
        RECT 77.915 124.475 79.835 124.645 ;
        RECT 77.575 124.135 79.475 124.305 ;
        RECT 77.805 123.795 78.135 123.915 ;
        RECT 76.885 123.625 78.135 123.795 ;
        RECT 74.410 123.165 75.425 123.365 ;
        RECT 75.595 122.985 76.005 123.425 ;
        RECT 76.295 123.195 76.545 123.625 ;
        RECT 76.745 122.985 77.065 123.445 ;
        RECT 78.305 123.375 78.475 124.135 ;
        RECT 79.145 124.075 79.475 124.135 ;
        RECT 78.665 123.905 78.995 123.965 ;
        RECT 78.665 123.635 79.325 123.905 ;
        RECT 79.645 123.580 79.835 124.475 ;
        RECT 77.625 123.205 78.475 123.375 ;
        RECT 78.675 122.985 79.335 123.465 ;
        RECT 79.515 123.250 79.835 123.580 ;
        RECT 80.035 124.225 80.285 124.815 ;
        RECT 80.465 124.735 80.750 125.535 ;
        RECT 80.930 125.195 81.185 125.225 ;
        RECT 80.930 125.025 81.270 125.195 ;
        RECT 80.930 124.555 81.185 125.025 ;
        RECT 80.035 123.895 80.835 124.225 ;
        RECT 80.035 123.245 80.285 123.895 ;
        RECT 81.005 123.695 81.185 124.555 ;
        RECT 82.190 124.775 82.705 125.185 ;
        RECT 82.940 124.775 83.110 125.535 ;
        RECT 83.280 125.195 85.310 125.365 ;
        RECT 82.190 123.965 82.530 124.775 ;
        RECT 83.280 124.530 83.450 125.195 ;
        RECT 83.845 124.855 84.970 125.025 ;
        RECT 82.700 124.340 83.450 124.530 ;
        RECT 83.620 124.515 84.630 124.685 ;
        RECT 82.190 123.795 83.420 123.965 ;
        RECT 80.465 122.985 80.750 123.445 ;
        RECT 80.930 123.165 81.185 123.695 ;
        RECT 82.465 123.190 82.710 123.795 ;
        RECT 82.930 122.985 83.440 123.520 ;
        RECT 83.620 123.155 83.810 124.515 ;
        RECT 83.980 124.175 84.255 124.315 ;
        RECT 83.980 124.005 84.260 124.175 ;
        RECT 83.980 123.155 84.255 124.005 ;
        RECT 84.460 123.715 84.630 124.515 ;
        RECT 84.800 123.725 84.970 124.855 ;
        RECT 85.140 124.225 85.310 125.195 ;
        RECT 85.480 124.395 85.650 125.535 ;
        RECT 85.820 124.395 86.155 125.365 ;
        RECT 85.140 123.895 85.335 124.225 ;
        RECT 85.560 123.895 85.815 124.225 ;
        RECT 85.560 123.725 85.730 123.895 ;
        RECT 85.985 123.725 86.155 124.395 ;
        RECT 86.330 124.370 86.620 125.535 ;
        RECT 87.915 124.565 88.245 125.365 ;
        RECT 88.415 124.735 88.745 125.535 ;
        RECT 89.045 124.565 89.375 125.365 ;
        RECT 90.020 124.735 90.270 125.535 ;
        RECT 87.915 124.395 90.350 124.565 ;
        RECT 90.540 124.395 90.710 125.535 ;
        RECT 90.880 124.395 91.220 125.365 ;
        RECT 87.710 123.975 88.060 124.225 ;
        RECT 88.245 123.765 88.415 124.395 ;
        RECT 88.585 123.975 88.915 124.175 ;
        RECT 89.085 123.975 89.415 124.175 ;
        RECT 89.585 123.975 90.005 124.175 ;
        RECT 90.180 124.145 90.350 124.395 ;
        RECT 90.180 123.975 90.875 124.145 ;
        RECT 84.800 123.555 85.730 123.725 ;
        RECT 84.800 123.520 84.975 123.555 ;
        RECT 84.445 123.155 84.975 123.520 ;
        RECT 85.400 122.985 85.730 123.385 ;
        RECT 85.900 123.155 86.155 123.725 ;
        RECT 86.330 122.985 86.620 123.710 ;
        RECT 87.915 123.155 88.415 123.765 ;
        RECT 89.045 123.635 90.270 123.805 ;
        RECT 91.045 123.785 91.220 124.395 ;
        RECT 91.390 124.445 93.060 125.535 ;
        RECT 93.345 124.905 93.630 125.365 ;
        RECT 93.800 125.075 94.070 125.535 ;
        RECT 93.345 124.685 94.300 124.905 ;
        RECT 91.390 123.925 92.140 124.445 ;
        RECT 89.045 123.155 89.375 123.635 ;
        RECT 89.545 122.985 89.770 123.445 ;
        RECT 89.940 123.155 90.270 123.635 ;
        RECT 90.460 122.985 90.710 123.785 ;
        RECT 90.880 123.155 91.220 123.785 ;
        RECT 92.310 123.755 93.060 124.275 ;
        RECT 93.230 123.955 93.920 124.515 ;
        RECT 94.090 123.785 94.300 124.685 ;
        RECT 91.390 122.985 93.060 123.755 ;
        RECT 93.345 123.615 94.300 123.785 ;
        RECT 94.470 124.515 94.870 125.365 ;
        RECT 95.060 124.905 95.340 125.365 ;
        RECT 95.860 125.075 96.185 125.535 ;
        RECT 95.060 124.685 96.185 124.905 ;
        RECT 94.470 123.955 95.565 124.515 ;
        RECT 95.735 124.225 96.185 124.685 ;
        RECT 96.355 124.395 96.740 125.365 ;
        RECT 93.345 123.155 93.630 123.615 ;
        RECT 93.800 122.985 94.070 123.445 ;
        RECT 94.470 123.155 94.870 123.955 ;
        RECT 95.735 123.895 96.290 124.225 ;
        RECT 95.735 123.785 96.185 123.895 ;
        RECT 95.060 123.615 96.185 123.785 ;
        RECT 96.460 123.725 96.740 124.395 ;
        RECT 95.060 123.155 95.340 123.615 ;
        RECT 95.860 122.985 96.185 123.445 ;
        RECT 96.355 123.155 96.740 123.725 ;
        RECT 96.915 124.345 97.170 125.225 ;
        RECT 97.340 124.395 97.645 125.535 ;
        RECT 97.985 125.155 98.315 125.535 ;
        RECT 98.495 124.985 98.665 125.275 ;
        RECT 98.835 125.075 99.085 125.535 ;
        RECT 97.865 124.815 98.665 124.985 ;
        RECT 99.255 125.025 100.125 125.365 ;
        RECT 96.915 123.695 97.125 124.345 ;
        RECT 97.865 124.225 98.035 124.815 ;
        RECT 99.255 124.645 99.425 125.025 ;
        RECT 100.360 124.905 100.530 125.365 ;
        RECT 100.700 125.075 101.070 125.535 ;
        RECT 101.365 124.935 101.535 125.275 ;
        RECT 101.705 125.105 102.035 125.535 ;
        RECT 102.270 124.935 102.440 125.275 ;
        RECT 98.205 124.475 99.425 124.645 ;
        RECT 99.595 124.565 100.055 124.855 ;
        RECT 100.360 124.735 100.920 124.905 ;
        RECT 101.365 124.765 102.440 124.935 ;
        RECT 102.610 125.035 103.290 125.365 ;
        RECT 103.505 125.035 103.755 125.365 ;
        RECT 103.925 125.075 104.175 125.535 ;
        RECT 100.750 124.595 100.920 124.735 ;
        RECT 99.595 124.555 100.560 124.565 ;
        RECT 99.255 124.385 99.425 124.475 ;
        RECT 99.885 124.395 100.560 124.555 ;
        RECT 97.295 124.195 98.035 124.225 ;
        RECT 97.295 123.895 98.210 124.195 ;
        RECT 97.885 123.720 98.210 123.895 ;
        RECT 96.915 123.165 97.170 123.695 ;
        RECT 97.340 122.985 97.645 123.445 ;
        RECT 97.890 123.365 98.210 123.720 ;
        RECT 98.380 123.935 98.920 124.305 ;
        RECT 99.255 124.215 99.660 124.385 ;
        RECT 98.380 123.535 98.620 123.935 ;
        RECT 99.100 123.765 99.320 124.045 ;
        RECT 98.790 123.595 99.320 123.765 ;
        RECT 98.790 123.365 98.960 123.595 ;
        RECT 99.490 123.435 99.660 124.215 ;
        RECT 99.830 123.605 100.180 124.225 ;
        RECT 100.350 123.605 100.560 124.395 ;
        RECT 100.750 124.425 102.250 124.595 ;
        RECT 100.750 123.735 100.920 124.425 ;
        RECT 102.610 124.255 102.780 125.035 ;
        RECT 103.585 124.905 103.755 125.035 ;
        RECT 101.090 124.085 102.780 124.255 ;
        RECT 102.950 124.475 103.415 124.865 ;
        RECT 103.585 124.735 103.980 124.905 ;
        RECT 101.090 123.905 101.260 124.085 ;
        RECT 97.890 123.195 98.960 123.365 ;
        RECT 99.130 122.985 99.320 123.425 ;
        RECT 99.490 123.155 100.440 123.435 ;
        RECT 100.750 123.345 101.010 123.735 ;
        RECT 101.430 123.665 102.220 123.915 ;
        RECT 100.660 123.175 101.010 123.345 ;
        RECT 101.220 122.985 101.550 123.445 ;
        RECT 102.425 123.375 102.595 124.085 ;
        RECT 102.950 123.885 103.120 124.475 ;
        RECT 102.765 123.665 103.120 123.885 ;
        RECT 103.290 123.665 103.640 124.285 ;
        RECT 103.810 123.375 103.980 124.735 ;
        RECT 104.345 124.565 104.670 125.350 ;
        RECT 104.150 123.515 104.610 124.565 ;
        RECT 102.425 123.205 103.280 123.375 ;
        RECT 103.485 123.205 103.980 123.375 ;
        RECT 104.150 122.985 104.480 123.345 ;
        RECT 104.840 123.245 105.010 125.365 ;
        RECT 105.180 125.035 105.510 125.535 ;
        RECT 105.680 124.865 105.935 125.365 ;
        RECT 105.185 124.695 105.935 124.865 ;
        RECT 105.185 123.705 105.415 124.695 ;
        RECT 105.585 123.875 105.935 124.525 ;
        RECT 106.110 124.445 107.320 125.535 ;
        RECT 107.490 124.445 111.000 125.535 ;
        RECT 111.170 124.445 112.380 125.535 ;
        RECT 106.110 123.905 106.630 124.445 ;
        RECT 106.800 123.735 107.320 124.275 ;
        RECT 107.490 123.925 109.180 124.445 ;
        RECT 109.350 123.755 111.000 124.275 ;
        RECT 111.170 123.905 111.690 124.445 ;
        RECT 105.185 123.535 105.935 123.705 ;
        RECT 105.180 122.985 105.510 123.365 ;
        RECT 105.680 123.245 105.935 123.535 ;
        RECT 106.110 122.985 107.320 123.735 ;
        RECT 107.490 122.985 111.000 123.755 ;
        RECT 111.860 123.735 112.380 124.275 ;
        RECT 111.170 122.985 112.380 123.735 ;
        RECT 18.165 122.815 112.465 122.985 ;
        RECT 18.250 122.065 19.460 122.815 ;
        RECT 18.250 121.525 18.770 122.065 ;
        RECT 20.090 122.045 21.760 122.815 ;
        RECT 21.930 122.090 22.220 122.815 ;
        RECT 22.390 122.065 23.600 122.815 ;
        RECT 18.940 121.355 19.460 121.895 ;
        RECT 18.250 120.265 19.460 121.355 ;
        RECT 20.090 121.355 20.840 121.875 ;
        RECT 21.010 121.525 21.760 122.045 ;
        RECT 20.090 120.265 21.760 121.355 ;
        RECT 21.930 120.265 22.220 121.430 ;
        RECT 22.390 121.355 22.910 121.895 ;
        RECT 23.080 121.525 23.600 122.065 ;
        RECT 23.830 121.995 24.040 122.815 ;
        RECT 24.210 122.015 24.540 122.645 ;
        RECT 24.210 121.415 24.460 122.015 ;
        RECT 24.710 121.995 24.940 122.815 ;
        RECT 25.150 122.065 26.360 122.815 ;
        RECT 24.630 121.575 24.960 121.825 ;
        RECT 22.390 120.265 23.600 121.355 ;
        RECT 23.830 120.265 24.040 121.405 ;
        RECT 24.210 120.435 24.540 121.415 ;
        RECT 24.710 120.265 24.940 121.405 ;
        RECT 25.150 121.355 25.670 121.895 ;
        RECT 25.840 121.525 26.360 122.065 ;
        RECT 26.735 122.035 27.235 122.645 ;
        RECT 26.530 121.575 26.880 121.825 ;
        RECT 27.065 121.405 27.235 122.035 ;
        RECT 27.865 122.165 28.195 122.645 ;
        RECT 28.365 122.355 28.590 122.815 ;
        RECT 28.760 122.165 29.090 122.645 ;
        RECT 27.865 121.995 29.090 122.165 ;
        RECT 29.280 122.015 29.530 122.815 ;
        RECT 29.700 122.015 30.040 122.645 ;
        RECT 30.215 122.265 30.470 122.555 ;
        RECT 30.640 122.435 30.970 122.815 ;
        RECT 30.215 122.095 30.965 122.265 ;
        RECT 27.405 121.625 27.735 121.825 ;
        RECT 27.905 121.625 28.235 121.825 ;
        RECT 28.405 121.625 28.825 121.825 ;
        RECT 29.000 121.655 29.695 121.825 ;
        RECT 29.000 121.405 29.170 121.655 ;
        RECT 29.865 121.405 30.040 122.015 ;
        RECT 25.150 120.265 26.360 121.355 ;
        RECT 26.735 121.235 29.170 121.405 ;
        RECT 26.735 120.435 27.065 121.235 ;
        RECT 27.235 120.265 27.565 121.065 ;
        RECT 27.865 120.435 28.195 121.235 ;
        RECT 28.840 120.265 29.090 121.065 ;
        RECT 29.360 120.265 29.530 121.405 ;
        RECT 29.700 120.435 30.040 121.405 ;
        RECT 30.215 121.275 30.565 121.925 ;
        RECT 30.735 121.105 30.965 122.095 ;
        RECT 30.215 120.935 30.965 121.105 ;
        RECT 30.215 120.435 30.470 120.935 ;
        RECT 30.640 120.265 30.970 120.765 ;
        RECT 31.140 120.435 31.310 122.555 ;
        RECT 31.670 122.455 32.000 122.815 ;
        RECT 32.170 122.425 32.665 122.595 ;
        RECT 32.870 122.425 33.725 122.595 ;
        RECT 31.540 121.235 32.000 122.285 ;
        RECT 31.480 120.450 31.805 121.235 ;
        RECT 32.170 121.065 32.340 122.425 ;
        RECT 32.510 121.515 32.860 122.135 ;
        RECT 33.030 121.915 33.385 122.135 ;
        RECT 33.030 121.325 33.200 121.915 ;
        RECT 33.555 121.715 33.725 122.425 ;
        RECT 34.600 122.355 34.930 122.815 ;
        RECT 35.140 122.455 35.490 122.625 ;
        RECT 33.930 121.885 34.720 122.135 ;
        RECT 35.140 122.065 35.400 122.455 ;
        RECT 35.710 122.365 36.660 122.645 ;
        RECT 36.830 122.375 37.020 122.815 ;
        RECT 37.190 122.435 38.260 122.605 ;
        RECT 34.890 121.715 35.060 121.895 ;
        RECT 32.170 120.895 32.565 121.065 ;
        RECT 32.735 120.935 33.200 121.325 ;
        RECT 33.370 121.545 35.060 121.715 ;
        RECT 32.395 120.765 32.565 120.895 ;
        RECT 33.370 120.765 33.540 121.545 ;
        RECT 35.230 121.375 35.400 122.065 ;
        RECT 33.900 121.205 35.400 121.375 ;
        RECT 35.590 121.405 35.800 122.195 ;
        RECT 35.970 121.575 36.320 122.195 ;
        RECT 36.490 121.585 36.660 122.365 ;
        RECT 37.190 122.205 37.360 122.435 ;
        RECT 36.830 122.035 37.360 122.205 ;
        RECT 36.830 121.755 37.050 122.035 ;
        RECT 37.530 121.865 37.770 122.265 ;
        RECT 36.490 121.415 36.895 121.585 ;
        RECT 37.230 121.495 37.770 121.865 ;
        RECT 37.940 122.080 38.260 122.435 ;
        RECT 38.505 122.355 38.810 122.815 ;
        RECT 38.980 122.105 39.235 122.635 ;
        RECT 37.940 121.905 38.265 122.080 ;
        RECT 37.940 121.605 38.855 121.905 ;
        RECT 38.115 121.575 38.855 121.605 ;
        RECT 35.590 121.245 36.265 121.405 ;
        RECT 36.725 121.325 36.895 121.415 ;
        RECT 35.590 121.235 36.555 121.245 ;
        RECT 35.230 121.065 35.400 121.205 ;
        RECT 31.975 120.265 32.225 120.725 ;
        RECT 32.395 120.435 32.645 120.765 ;
        RECT 32.860 120.435 33.540 120.765 ;
        RECT 33.710 120.865 34.785 121.035 ;
        RECT 35.230 120.895 35.790 121.065 ;
        RECT 36.095 120.945 36.555 121.235 ;
        RECT 36.725 121.155 37.945 121.325 ;
        RECT 33.710 120.525 33.880 120.865 ;
        RECT 34.115 120.265 34.445 120.695 ;
        RECT 34.615 120.525 34.785 120.865 ;
        RECT 35.080 120.265 35.450 120.725 ;
        RECT 35.620 120.435 35.790 120.895 ;
        RECT 36.725 120.775 36.895 121.155 ;
        RECT 38.115 120.985 38.285 121.575 ;
        RECT 39.025 121.455 39.235 122.105 ;
        RECT 39.985 122.185 40.270 122.645 ;
        RECT 40.440 122.355 40.710 122.815 ;
        RECT 39.985 122.015 40.940 122.185 ;
        RECT 36.025 120.435 36.895 120.775 ;
        RECT 37.485 120.815 38.285 120.985 ;
        RECT 37.065 120.265 37.315 120.725 ;
        RECT 37.485 120.525 37.655 120.815 ;
        RECT 37.835 120.265 38.165 120.645 ;
        RECT 38.505 120.265 38.810 121.405 ;
        RECT 38.980 120.575 39.235 121.455 ;
        RECT 39.870 121.285 40.560 121.845 ;
        RECT 40.730 121.115 40.940 122.015 ;
        RECT 39.985 120.895 40.940 121.115 ;
        RECT 41.110 121.845 41.510 122.645 ;
        RECT 41.700 122.185 41.980 122.645 ;
        RECT 42.500 122.355 42.825 122.815 ;
        RECT 41.700 122.015 42.825 122.185 ;
        RECT 42.995 122.075 43.380 122.645 ;
        RECT 42.375 121.905 42.825 122.015 ;
        RECT 41.110 121.285 42.205 121.845 ;
        RECT 42.375 121.575 42.930 121.905 ;
        RECT 39.985 120.435 40.270 120.895 ;
        RECT 40.440 120.265 40.710 120.725 ;
        RECT 41.110 120.435 41.510 121.285 ;
        RECT 42.375 121.115 42.825 121.575 ;
        RECT 43.100 121.405 43.380 122.075 ;
        RECT 43.825 122.005 44.070 122.610 ;
        RECT 44.290 122.280 44.800 122.815 ;
        RECT 41.700 120.895 42.825 121.115 ;
        RECT 41.700 120.435 41.980 120.895 ;
        RECT 42.500 120.265 42.825 120.725 ;
        RECT 42.995 120.435 43.380 121.405 ;
        RECT 43.550 121.835 44.780 122.005 ;
        RECT 43.550 121.025 43.890 121.835 ;
        RECT 44.060 121.270 44.810 121.460 ;
        RECT 43.550 120.615 44.065 121.025 ;
        RECT 44.300 120.265 44.470 121.025 ;
        RECT 44.640 120.605 44.810 121.270 ;
        RECT 44.980 121.285 45.170 122.645 ;
        RECT 45.340 121.795 45.615 122.645 ;
        RECT 45.805 122.280 46.335 122.645 ;
        RECT 46.760 122.415 47.090 122.815 ;
        RECT 46.160 122.245 46.335 122.280 ;
        RECT 45.340 121.625 45.620 121.795 ;
        RECT 45.340 121.485 45.615 121.625 ;
        RECT 45.820 121.285 45.990 122.085 ;
        RECT 44.980 121.115 45.990 121.285 ;
        RECT 46.160 122.075 47.090 122.245 ;
        RECT 47.260 122.075 47.515 122.645 ;
        RECT 47.690 122.090 47.980 122.815 ;
        RECT 46.160 120.945 46.330 122.075 ;
        RECT 46.920 121.905 47.090 122.075 ;
        RECT 45.205 120.775 46.330 120.945 ;
        RECT 46.500 121.575 46.695 121.905 ;
        RECT 46.920 121.575 47.175 121.905 ;
        RECT 46.500 120.605 46.670 121.575 ;
        RECT 47.345 121.405 47.515 122.075 ;
        RECT 48.670 121.995 48.880 122.815 ;
        RECT 49.050 122.015 49.380 122.645 ;
        RECT 44.640 120.435 46.670 120.605 ;
        RECT 46.840 120.265 47.010 121.405 ;
        RECT 47.180 120.435 47.515 121.405 ;
        RECT 47.690 120.265 47.980 121.430 ;
        RECT 49.050 121.415 49.300 122.015 ;
        RECT 49.550 121.995 49.780 122.815 ;
        RECT 50.265 122.005 50.510 122.610 ;
        RECT 50.730 122.280 51.240 122.815 ;
        RECT 49.990 121.835 51.220 122.005 ;
        RECT 49.470 121.575 49.800 121.825 ;
        RECT 48.670 120.265 48.880 121.405 ;
        RECT 49.050 120.435 49.380 121.415 ;
        RECT 49.550 120.265 49.780 121.405 ;
        RECT 49.990 121.025 50.330 121.835 ;
        RECT 50.500 121.270 51.250 121.460 ;
        RECT 49.990 120.615 50.505 121.025 ;
        RECT 50.740 120.265 50.910 121.025 ;
        RECT 51.080 120.605 51.250 121.270 ;
        RECT 51.420 121.285 51.610 122.645 ;
        RECT 51.780 122.475 52.055 122.645 ;
        RECT 51.780 122.305 52.060 122.475 ;
        RECT 51.780 121.485 52.055 122.305 ;
        RECT 52.245 122.280 52.775 122.645 ;
        RECT 53.200 122.415 53.530 122.815 ;
        RECT 52.600 122.245 52.775 122.280 ;
        RECT 52.260 121.285 52.430 122.085 ;
        RECT 51.420 121.115 52.430 121.285 ;
        RECT 52.600 122.075 53.530 122.245 ;
        RECT 53.700 122.075 53.955 122.645 ;
        RECT 52.600 120.945 52.770 122.075 ;
        RECT 53.360 121.905 53.530 122.075 ;
        RECT 51.645 120.775 52.770 120.945 ;
        RECT 52.940 121.575 53.135 121.905 ;
        RECT 53.360 121.575 53.615 121.905 ;
        RECT 52.940 120.605 53.110 121.575 ;
        RECT 53.785 121.405 53.955 122.075 ;
        RECT 55.165 122.185 55.450 122.645 ;
        RECT 55.620 122.355 55.890 122.815 ;
        RECT 55.165 122.015 56.120 122.185 ;
        RECT 51.080 120.435 53.110 120.605 ;
        RECT 53.280 120.265 53.450 121.405 ;
        RECT 53.620 120.435 53.955 121.405 ;
        RECT 55.050 121.285 55.740 121.845 ;
        RECT 55.910 121.115 56.120 122.015 ;
        RECT 55.165 120.895 56.120 121.115 ;
        RECT 56.290 121.845 56.690 122.645 ;
        RECT 56.880 122.185 57.160 122.645 ;
        RECT 57.680 122.355 58.005 122.815 ;
        RECT 56.880 122.015 58.005 122.185 ;
        RECT 58.175 122.075 58.560 122.645 ;
        RECT 57.555 121.905 58.005 122.015 ;
        RECT 56.290 121.285 57.385 121.845 ;
        RECT 57.555 121.575 58.110 121.905 ;
        RECT 55.165 120.435 55.450 120.895 ;
        RECT 55.620 120.265 55.890 120.725 ;
        RECT 56.290 120.435 56.690 121.285 ;
        RECT 57.555 121.115 58.005 121.575 ;
        RECT 58.280 121.405 58.560 122.075 ;
        RECT 56.880 120.895 58.005 121.115 ;
        RECT 56.880 120.435 57.160 120.895 ;
        RECT 57.680 120.265 58.005 120.725 ;
        RECT 58.175 120.435 58.560 121.405 ;
        RECT 59.650 122.015 59.990 122.645 ;
        RECT 60.160 122.015 60.410 122.815 ;
        RECT 60.600 122.165 60.930 122.645 ;
        RECT 61.100 122.355 61.325 122.815 ;
        RECT 61.495 122.165 61.825 122.645 ;
        RECT 59.650 121.405 59.825 122.015 ;
        RECT 60.600 121.995 61.825 122.165 ;
        RECT 62.455 122.035 62.955 122.645 ;
        RECT 63.445 122.185 63.730 122.645 ;
        RECT 63.900 122.355 64.170 122.815 ;
        RECT 59.995 121.655 60.690 121.825 ;
        RECT 60.520 121.405 60.690 121.655 ;
        RECT 60.865 121.625 61.285 121.825 ;
        RECT 61.455 121.625 61.785 121.825 ;
        RECT 61.955 121.625 62.285 121.825 ;
        RECT 62.455 121.405 62.625 122.035 ;
        RECT 63.445 122.015 64.400 122.185 ;
        RECT 62.810 121.575 63.160 121.825 ;
        RECT 59.650 120.435 59.990 121.405 ;
        RECT 60.160 120.265 60.330 121.405 ;
        RECT 60.520 121.235 62.955 121.405 ;
        RECT 63.330 121.285 64.020 121.845 ;
        RECT 60.600 120.265 60.850 121.065 ;
        RECT 61.495 120.435 61.825 121.235 ;
        RECT 62.125 120.265 62.455 121.065 ;
        RECT 62.625 120.435 62.955 121.235 ;
        RECT 64.190 121.115 64.400 122.015 ;
        RECT 63.445 120.895 64.400 121.115 ;
        RECT 64.570 121.845 64.970 122.645 ;
        RECT 65.160 122.185 65.440 122.645 ;
        RECT 65.960 122.355 66.285 122.815 ;
        RECT 65.160 122.015 66.285 122.185 ;
        RECT 66.455 122.075 66.840 122.645 ;
        RECT 65.835 121.905 66.285 122.015 ;
        RECT 64.570 121.285 65.665 121.845 ;
        RECT 65.835 121.575 66.390 121.905 ;
        RECT 63.445 120.435 63.730 120.895 ;
        RECT 63.900 120.265 64.170 120.725 ;
        RECT 64.570 120.435 64.970 121.285 ;
        RECT 65.835 121.115 66.285 121.575 ;
        RECT 66.560 121.405 66.840 122.075 ;
        RECT 65.160 120.895 66.285 121.115 ;
        RECT 65.160 120.435 65.440 120.895 ;
        RECT 65.960 120.265 66.285 120.725 ;
        RECT 66.455 120.435 66.840 121.405 ;
        RECT 67.015 122.075 67.270 122.645 ;
        RECT 67.440 122.415 67.770 122.815 ;
        RECT 68.195 122.280 68.725 122.645 ;
        RECT 68.195 122.245 68.370 122.280 ;
        RECT 67.440 122.075 68.370 122.245 ;
        RECT 68.915 122.135 69.190 122.645 ;
        RECT 67.015 121.405 67.185 122.075 ;
        RECT 67.440 121.905 67.610 122.075 ;
        RECT 67.355 121.575 67.610 121.905 ;
        RECT 67.835 121.575 68.030 121.905 ;
        RECT 67.015 120.435 67.350 121.405 ;
        RECT 67.520 120.265 67.690 121.405 ;
        RECT 67.860 120.605 68.030 121.575 ;
        RECT 68.200 120.945 68.370 122.075 ;
        RECT 68.540 121.285 68.710 122.085 ;
        RECT 68.910 121.965 69.190 122.135 ;
        RECT 68.915 121.485 69.190 121.965 ;
        RECT 69.360 121.285 69.550 122.645 ;
        RECT 69.730 122.280 70.240 122.815 ;
        RECT 70.460 122.005 70.705 122.610 ;
        RECT 71.615 122.345 71.945 122.815 ;
        RECT 72.115 122.175 72.340 122.620 ;
        RECT 72.510 122.290 72.805 122.815 ;
        RECT 71.610 122.005 72.340 122.175 ;
        RECT 73.450 122.090 73.740 122.815 ;
        RECT 69.750 121.835 70.980 122.005 ;
        RECT 68.540 121.115 69.550 121.285 ;
        RECT 69.720 121.270 70.470 121.460 ;
        RECT 68.200 120.775 69.325 120.945 ;
        RECT 69.720 120.605 69.890 121.270 ;
        RECT 70.640 121.025 70.980 121.835 ;
        RECT 71.610 121.440 71.890 122.005 ;
        RECT 73.950 121.995 74.180 122.815 ;
        RECT 74.350 122.015 74.680 122.645 ;
        RECT 72.060 121.610 73.280 121.835 ;
        RECT 73.930 121.575 74.260 121.825 ;
        RECT 71.610 121.270 73.210 121.440 ;
        RECT 67.860 120.435 69.890 120.605 ;
        RECT 70.060 120.265 70.230 121.025 ;
        RECT 70.465 120.615 70.980 121.025 ;
        RECT 71.670 120.265 71.925 121.100 ;
        RECT 72.095 120.465 72.355 121.270 ;
        RECT 72.525 120.265 72.785 121.100 ;
        RECT 72.955 120.465 73.210 121.270 ;
        RECT 73.450 120.265 73.740 121.430 ;
        RECT 74.430 121.415 74.680 122.015 ;
        RECT 74.850 121.995 75.060 122.815 ;
        RECT 75.290 122.075 75.675 122.645 ;
        RECT 75.845 122.355 76.170 122.815 ;
        RECT 76.690 122.185 76.970 122.645 ;
        RECT 73.950 120.265 74.180 121.405 ;
        RECT 74.350 120.435 74.680 121.415 ;
        RECT 75.290 121.405 75.570 122.075 ;
        RECT 75.845 122.015 76.970 122.185 ;
        RECT 75.845 121.905 76.295 122.015 ;
        RECT 75.740 121.575 76.295 121.905 ;
        RECT 77.160 121.845 77.560 122.645 ;
        RECT 77.960 122.355 78.230 122.815 ;
        RECT 78.400 122.185 78.685 122.645 ;
        RECT 74.850 120.265 75.060 121.405 ;
        RECT 75.290 120.435 75.675 121.405 ;
        RECT 75.845 121.115 76.295 121.575 ;
        RECT 76.465 121.285 77.560 121.845 ;
        RECT 75.845 120.895 76.970 121.115 ;
        RECT 75.845 120.265 76.170 120.725 ;
        RECT 76.690 120.435 76.970 120.895 ;
        RECT 77.160 120.435 77.560 121.285 ;
        RECT 77.730 122.015 78.685 122.185 ;
        RECT 78.970 122.315 79.270 122.645 ;
        RECT 79.440 122.335 79.715 122.815 ;
        RECT 77.730 121.115 77.940 122.015 ;
        RECT 78.110 121.285 78.800 121.845 ;
        RECT 78.970 121.405 79.140 122.315 ;
        RECT 79.895 122.165 80.190 122.555 ;
        RECT 80.360 122.335 80.615 122.815 ;
        RECT 80.790 122.165 81.050 122.555 ;
        RECT 81.220 122.335 81.500 122.815 ;
        RECT 79.310 121.575 79.660 122.145 ;
        RECT 79.895 121.995 81.545 122.165 ;
        RECT 81.730 122.065 82.940 122.815 ;
        RECT 79.830 121.655 80.970 121.825 ;
        RECT 79.830 121.405 80.000 121.655 ;
        RECT 81.140 121.485 81.545 121.995 ;
        RECT 78.970 121.235 80.000 121.405 ;
        RECT 80.790 121.315 81.545 121.485 ;
        RECT 81.730 121.355 82.250 121.895 ;
        RECT 82.420 121.525 82.940 122.065 ;
        RECT 83.110 122.015 83.450 122.645 ;
        RECT 83.620 122.015 83.870 122.815 ;
        RECT 84.060 122.165 84.390 122.645 ;
        RECT 84.560 122.355 84.785 122.815 ;
        RECT 84.955 122.165 85.285 122.645 ;
        RECT 83.110 121.405 83.285 122.015 ;
        RECT 84.060 121.995 85.285 122.165 ;
        RECT 85.915 122.035 86.415 122.645 ;
        RECT 83.455 121.655 84.150 121.825 ;
        RECT 83.980 121.405 84.150 121.655 ;
        RECT 84.325 121.625 84.745 121.825 ;
        RECT 84.915 121.625 85.245 121.825 ;
        RECT 85.415 121.625 85.745 121.825 ;
        RECT 85.915 121.405 86.085 122.035 ;
        RECT 86.790 122.015 87.130 122.645 ;
        RECT 87.300 122.015 87.550 122.815 ;
        RECT 87.740 122.165 88.070 122.645 ;
        RECT 88.240 122.355 88.465 122.815 ;
        RECT 88.635 122.165 88.965 122.645 ;
        RECT 86.270 121.575 86.620 121.825 ;
        RECT 86.790 121.405 86.965 122.015 ;
        RECT 87.740 121.995 88.965 122.165 ;
        RECT 89.595 122.035 90.095 122.645 ;
        RECT 91.595 122.035 92.095 122.645 ;
        RECT 87.135 121.655 87.830 121.825 ;
        RECT 87.660 121.405 87.830 121.655 ;
        RECT 88.005 121.625 88.425 121.825 ;
        RECT 88.595 121.625 88.925 121.825 ;
        RECT 89.095 121.625 89.425 121.825 ;
        RECT 89.595 121.405 89.765 122.035 ;
        RECT 89.950 121.575 90.300 121.825 ;
        RECT 91.390 121.575 91.740 121.825 ;
        RECT 91.925 121.405 92.095 122.035 ;
        RECT 92.725 122.165 93.055 122.645 ;
        RECT 93.225 122.355 93.450 122.815 ;
        RECT 93.620 122.165 93.950 122.645 ;
        RECT 92.725 121.995 93.950 122.165 ;
        RECT 94.140 122.015 94.390 122.815 ;
        RECT 94.560 122.015 94.900 122.645 ;
        RECT 92.265 121.625 92.595 121.825 ;
        RECT 92.765 121.625 93.095 121.825 ;
        RECT 93.265 121.625 93.685 121.825 ;
        RECT 93.860 121.655 94.555 121.825 ;
        RECT 93.860 121.405 94.030 121.655 ;
        RECT 94.725 121.405 94.900 122.015 ;
        RECT 95.345 122.005 95.590 122.610 ;
        RECT 95.810 122.280 96.320 122.815 ;
        RECT 77.730 120.895 78.685 121.115 ;
        RECT 77.960 120.265 78.230 120.725 ;
        RECT 78.400 120.435 78.685 120.895 ;
        RECT 78.970 120.435 79.280 121.235 ;
        RECT 80.790 121.065 81.050 121.315 ;
        RECT 79.450 120.265 79.760 121.065 ;
        RECT 79.930 120.895 81.050 121.065 ;
        RECT 79.930 120.435 80.190 120.895 ;
        RECT 80.360 120.265 80.615 120.725 ;
        RECT 80.790 120.435 81.050 120.895 ;
        RECT 81.220 120.265 81.505 121.135 ;
        RECT 81.730 120.265 82.940 121.355 ;
        RECT 83.110 120.435 83.450 121.405 ;
        RECT 83.620 120.265 83.790 121.405 ;
        RECT 83.980 121.235 86.415 121.405 ;
        RECT 84.060 120.265 84.310 121.065 ;
        RECT 84.955 120.435 85.285 121.235 ;
        RECT 85.585 120.265 85.915 121.065 ;
        RECT 86.085 120.435 86.415 121.235 ;
        RECT 86.790 120.435 87.130 121.405 ;
        RECT 87.300 120.265 87.470 121.405 ;
        RECT 87.660 121.235 90.095 121.405 ;
        RECT 87.740 120.265 87.990 121.065 ;
        RECT 88.635 120.435 88.965 121.235 ;
        RECT 89.265 120.265 89.595 121.065 ;
        RECT 89.765 120.435 90.095 121.235 ;
        RECT 91.595 121.235 94.030 121.405 ;
        RECT 91.595 120.435 91.925 121.235 ;
        RECT 92.095 120.265 92.425 121.065 ;
        RECT 92.725 120.435 93.055 121.235 ;
        RECT 93.700 120.265 93.950 121.065 ;
        RECT 94.220 120.265 94.390 121.405 ;
        RECT 94.560 120.435 94.900 121.405 ;
        RECT 95.070 121.835 96.300 122.005 ;
        RECT 95.070 121.025 95.410 121.835 ;
        RECT 95.580 121.270 96.330 121.460 ;
        RECT 95.070 120.615 95.585 121.025 ;
        RECT 95.820 120.265 95.990 121.025 ;
        RECT 96.160 120.605 96.330 121.270 ;
        RECT 96.500 121.285 96.690 122.645 ;
        RECT 96.860 121.795 97.135 122.645 ;
        RECT 97.325 122.280 97.855 122.645 ;
        RECT 98.280 122.415 98.610 122.815 ;
        RECT 97.680 122.245 97.855 122.280 ;
        RECT 96.860 121.625 97.140 121.795 ;
        RECT 96.860 121.485 97.135 121.625 ;
        RECT 97.340 121.285 97.510 122.085 ;
        RECT 96.500 121.115 97.510 121.285 ;
        RECT 97.680 122.075 98.610 122.245 ;
        RECT 98.780 122.075 99.035 122.645 ;
        RECT 99.210 122.090 99.500 122.815 ;
        RECT 99.785 122.185 100.070 122.645 ;
        RECT 100.240 122.355 100.510 122.815 ;
        RECT 97.680 120.945 97.850 122.075 ;
        RECT 98.440 121.905 98.610 122.075 ;
        RECT 96.725 120.775 97.850 120.945 ;
        RECT 98.020 121.575 98.215 121.905 ;
        RECT 98.440 121.575 98.695 121.905 ;
        RECT 98.020 120.605 98.190 121.575 ;
        RECT 98.865 121.405 99.035 122.075 ;
        RECT 99.785 122.015 100.740 122.185 ;
        RECT 96.160 120.435 98.190 120.605 ;
        RECT 98.360 120.265 98.530 121.405 ;
        RECT 98.700 120.435 99.035 121.405 ;
        RECT 99.210 120.265 99.500 121.430 ;
        RECT 99.670 121.285 100.360 121.845 ;
        RECT 100.530 121.115 100.740 122.015 ;
        RECT 99.785 120.895 100.740 121.115 ;
        RECT 100.910 121.845 101.310 122.645 ;
        RECT 101.500 122.185 101.780 122.645 ;
        RECT 102.300 122.355 102.625 122.815 ;
        RECT 101.500 122.015 102.625 122.185 ;
        RECT 102.795 122.075 103.180 122.645 ;
        RECT 102.175 121.905 102.625 122.015 ;
        RECT 100.910 121.285 102.005 121.845 ;
        RECT 102.175 121.575 102.730 121.905 ;
        RECT 99.785 120.435 100.070 120.895 ;
        RECT 100.240 120.265 100.510 120.725 ;
        RECT 100.910 120.435 101.310 121.285 ;
        RECT 102.175 121.115 102.625 121.575 ;
        RECT 102.900 121.405 103.180 122.075 ;
        RECT 103.390 121.995 103.620 122.815 ;
        RECT 103.790 122.015 104.120 122.645 ;
        RECT 103.370 121.575 103.700 121.825 ;
        RECT 103.870 121.415 104.120 122.015 ;
        RECT 104.290 121.995 104.500 122.815 ;
        RECT 105.655 122.270 111.000 122.815 ;
        RECT 101.500 120.895 102.625 121.115 ;
        RECT 101.500 120.435 101.780 120.895 ;
        RECT 102.300 120.265 102.625 120.725 ;
        RECT 102.795 120.435 103.180 121.405 ;
        RECT 103.390 120.265 103.620 121.405 ;
        RECT 103.790 120.435 104.120 121.415 ;
        RECT 104.290 120.265 104.500 121.405 ;
        RECT 107.245 120.700 107.595 121.950 ;
        RECT 109.075 121.440 109.415 122.270 ;
        RECT 111.170 122.065 112.380 122.815 ;
        RECT 111.170 121.355 111.690 121.895 ;
        RECT 111.860 121.525 112.380 122.065 ;
        RECT 105.655 120.265 111.000 120.700 ;
        RECT 111.170 120.265 112.380 121.355 ;
        RECT 18.165 120.095 112.465 120.265 ;
        RECT 18.250 119.005 19.460 120.095 ;
        RECT 19.940 119.255 20.110 120.095 ;
        RECT 20.320 119.085 20.570 119.925 ;
        RECT 20.780 119.255 20.950 120.095 ;
        RECT 21.120 119.085 21.410 119.925 ;
        RECT 18.250 118.295 18.770 118.835 ;
        RECT 18.940 118.465 19.460 119.005 ;
        RECT 19.685 118.915 21.410 119.085 ;
        RECT 21.620 119.035 21.790 120.095 ;
        RECT 22.085 119.715 22.415 120.095 ;
        RECT 22.595 119.545 22.765 119.835 ;
        RECT 22.935 119.635 23.185 120.095 ;
        RECT 21.965 119.375 22.765 119.545 ;
        RECT 23.355 119.585 24.225 119.925 ;
        RECT 19.685 118.365 20.095 118.915 ;
        RECT 21.965 118.755 22.135 119.375 ;
        RECT 23.355 119.205 23.525 119.585 ;
        RECT 24.460 119.465 24.630 119.925 ;
        RECT 24.800 119.635 25.170 120.095 ;
        RECT 25.465 119.495 25.635 119.835 ;
        RECT 25.805 119.665 26.135 120.095 ;
        RECT 26.370 119.495 26.540 119.835 ;
        RECT 22.305 119.035 23.525 119.205 ;
        RECT 23.695 119.125 24.155 119.415 ;
        RECT 24.460 119.295 25.020 119.465 ;
        RECT 25.465 119.325 26.540 119.495 ;
        RECT 26.710 119.595 27.390 119.925 ;
        RECT 27.605 119.595 27.855 119.925 ;
        RECT 28.025 119.635 28.275 120.095 ;
        RECT 24.850 119.155 25.020 119.295 ;
        RECT 23.695 119.115 24.660 119.125 ;
        RECT 23.355 118.945 23.525 119.035 ;
        RECT 23.985 118.955 24.660 119.115 ;
        RECT 21.965 118.745 22.310 118.755 ;
        RECT 20.280 118.535 22.310 118.745 ;
        RECT 18.250 117.545 19.460 118.295 ;
        RECT 19.685 118.195 21.450 118.365 ;
        RECT 19.940 117.545 20.110 118.015 ;
        RECT 20.280 117.715 20.610 118.195 ;
        RECT 20.780 117.545 20.950 118.015 ;
        RECT 21.120 117.715 21.450 118.195 ;
        RECT 21.620 117.545 21.790 118.355 ;
        RECT 21.985 118.280 22.310 118.535 ;
        RECT 21.990 117.925 22.310 118.280 ;
        RECT 22.480 118.495 23.020 118.865 ;
        RECT 23.355 118.775 23.760 118.945 ;
        RECT 22.480 118.095 22.720 118.495 ;
        RECT 23.200 118.325 23.420 118.605 ;
        RECT 22.890 118.155 23.420 118.325 ;
        RECT 22.890 117.925 23.060 118.155 ;
        RECT 23.590 117.995 23.760 118.775 ;
        RECT 23.930 118.165 24.280 118.785 ;
        RECT 24.450 118.165 24.660 118.955 ;
        RECT 24.850 118.985 26.350 119.155 ;
        RECT 24.850 118.295 25.020 118.985 ;
        RECT 26.710 118.815 26.880 119.595 ;
        RECT 27.685 119.465 27.855 119.595 ;
        RECT 25.190 118.645 26.880 118.815 ;
        RECT 27.050 119.035 27.515 119.425 ;
        RECT 27.685 119.295 28.080 119.465 ;
        RECT 25.190 118.465 25.360 118.645 ;
        RECT 21.990 117.755 23.060 117.925 ;
        RECT 23.230 117.545 23.420 117.985 ;
        RECT 23.590 117.715 24.540 117.995 ;
        RECT 24.850 117.905 25.110 118.295 ;
        RECT 25.530 118.225 26.320 118.475 ;
        RECT 24.760 117.735 25.110 117.905 ;
        RECT 25.320 117.545 25.650 118.005 ;
        RECT 26.525 117.935 26.695 118.645 ;
        RECT 27.050 118.445 27.220 119.035 ;
        RECT 26.865 118.225 27.220 118.445 ;
        RECT 27.390 118.225 27.740 118.845 ;
        RECT 27.910 117.935 28.080 119.295 ;
        RECT 28.445 119.125 28.770 119.910 ;
        RECT 28.250 118.075 28.710 119.125 ;
        RECT 26.525 117.765 27.380 117.935 ;
        RECT 27.585 117.765 28.080 117.935 ;
        RECT 28.250 117.545 28.580 117.905 ;
        RECT 28.940 117.805 29.110 119.925 ;
        RECT 29.280 119.595 29.610 120.095 ;
        RECT 29.780 119.425 30.035 119.925 ;
        RECT 29.285 119.255 30.035 119.425 ;
        RECT 29.285 118.265 29.515 119.255 ;
        RECT 29.685 118.435 30.035 119.085 ;
        RECT 31.130 118.955 31.515 119.925 ;
        RECT 31.685 119.635 32.010 120.095 ;
        RECT 32.530 119.465 32.810 119.925 ;
        RECT 31.685 119.245 32.810 119.465 ;
        RECT 31.130 118.285 31.410 118.955 ;
        RECT 31.685 118.785 32.135 119.245 ;
        RECT 33.000 119.075 33.400 119.925 ;
        RECT 33.800 119.635 34.070 120.095 ;
        RECT 34.240 119.465 34.525 119.925 ;
        RECT 31.580 118.455 32.135 118.785 ;
        RECT 32.305 118.515 33.400 119.075 ;
        RECT 31.685 118.345 32.135 118.455 ;
        RECT 29.285 118.095 30.035 118.265 ;
        RECT 29.280 117.545 29.610 117.925 ;
        RECT 29.780 117.805 30.035 118.095 ;
        RECT 31.130 117.715 31.515 118.285 ;
        RECT 31.685 118.175 32.810 118.345 ;
        RECT 31.685 117.545 32.010 118.005 ;
        RECT 32.530 117.715 32.810 118.175 ;
        RECT 33.000 117.715 33.400 118.515 ;
        RECT 33.570 119.245 34.525 119.465 ;
        RECT 33.570 118.345 33.780 119.245 ;
        RECT 33.950 118.515 34.640 119.075 ;
        RECT 34.810 118.930 35.100 120.095 ;
        RECT 35.270 118.955 35.610 119.925 ;
        RECT 35.780 118.955 35.950 120.095 ;
        RECT 36.220 119.295 36.470 120.095 ;
        RECT 37.115 119.125 37.445 119.925 ;
        RECT 37.745 119.295 38.075 120.095 ;
        RECT 38.245 119.125 38.575 119.925 ;
        RECT 38.955 119.425 39.210 119.925 ;
        RECT 39.380 119.595 39.710 120.095 ;
        RECT 38.955 119.255 39.705 119.425 ;
        RECT 36.140 118.955 38.575 119.125 ;
        RECT 35.270 118.345 35.445 118.955 ;
        RECT 36.140 118.705 36.310 118.955 ;
        RECT 35.615 118.535 36.310 118.705 ;
        RECT 36.485 118.535 36.905 118.735 ;
        RECT 37.075 118.535 37.405 118.735 ;
        RECT 37.575 118.535 37.905 118.735 ;
        RECT 33.570 118.175 34.525 118.345 ;
        RECT 33.800 117.545 34.070 118.005 ;
        RECT 34.240 117.715 34.525 118.175 ;
        RECT 34.810 117.545 35.100 118.270 ;
        RECT 35.270 117.715 35.610 118.345 ;
        RECT 35.780 117.545 36.030 118.345 ;
        RECT 36.220 118.195 37.445 118.365 ;
        RECT 36.220 117.715 36.550 118.195 ;
        RECT 36.720 117.545 36.945 118.005 ;
        RECT 37.115 117.715 37.445 118.195 ;
        RECT 38.075 118.325 38.245 118.955 ;
        RECT 38.430 118.535 38.780 118.785 ;
        RECT 38.955 118.435 39.305 119.085 ;
        RECT 38.075 117.715 38.575 118.325 ;
        RECT 39.475 118.265 39.705 119.255 ;
        RECT 38.955 118.095 39.705 118.265 ;
        RECT 38.955 117.805 39.210 118.095 ;
        RECT 39.380 117.545 39.710 117.925 ;
        RECT 39.880 117.805 40.050 119.925 ;
        RECT 40.220 119.125 40.545 119.910 ;
        RECT 40.715 119.635 40.965 120.095 ;
        RECT 41.135 119.595 41.385 119.925 ;
        RECT 41.600 119.595 42.280 119.925 ;
        RECT 41.135 119.465 41.305 119.595 ;
        RECT 40.910 119.295 41.305 119.465 ;
        RECT 40.280 118.075 40.740 119.125 ;
        RECT 40.910 117.935 41.080 119.295 ;
        RECT 41.475 119.035 41.940 119.425 ;
        RECT 41.250 118.225 41.600 118.845 ;
        RECT 41.770 118.445 41.940 119.035 ;
        RECT 42.110 118.815 42.280 119.595 ;
        RECT 42.450 119.495 42.620 119.835 ;
        RECT 42.855 119.665 43.185 120.095 ;
        RECT 43.355 119.495 43.525 119.835 ;
        RECT 43.820 119.635 44.190 120.095 ;
        RECT 42.450 119.325 43.525 119.495 ;
        RECT 44.360 119.465 44.530 119.925 ;
        RECT 44.765 119.585 45.635 119.925 ;
        RECT 45.805 119.635 46.055 120.095 ;
        RECT 43.970 119.295 44.530 119.465 ;
        RECT 43.970 119.155 44.140 119.295 ;
        RECT 42.640 118.985 44.140 119.155 ;
        RECT 44.835 119.125 45.295 119.415 ;
        RECT 42.110 118.645 43.800 118.815 ;
        RECT 41.770 118.225 42.125 118.445 ;
        RECT 42.295 117.935 42.465 118.645 ;
        RECT 42.670 118.225 43.460 118.475 ;
        RECT 43.630 118.465 43.800 118.645 ;
        RECT 43.970 118.295 44.140 118.985 ;
        RECT 40.410 117.545 40.740 117.905 ;
        RECT 40.910 117.765 41.405 117.935 ;
        RECT 41.610 117.765 42.465 117.935 ;
        RECT 43.340 117.545 43.670 118.005 ;
        RECT 43.880 117.905 44.140 118.295 ;
        RECT 44.330 119.115 45.295 119.125 ;
        RECT 45.465 119.205 45.635 119.585 ;
        RECT 46.225 119.545 46.395 119.835 ;
        RECT 46.575 119.715 46.905 120.095 ;
        RECT 46.225 119.375 47.025 119.545 ;
        RECT 44.330 118.955 45.005 119.115 ;
        RECT 45.465 119.035 46.685 119.205 ;
        RECT 44.330 118.165 44.540 118.955 ;
        RECT 45.465 118.945 45.635 119.035 ;
        RECT 44.710 118.165 45.060 118.785 ;
        RECT 45.230 118.775 45.635 118.945 ;
        RECT 45.230 117.995 45.400 118.775 ;
        RECT 45.570 118.325 45.790 118.605 ;
        RECT 45.970 118.495 46.510 118.865 ;
        RECT 46.855 118.785 47.025 119.375 ;
        RECT 47.245 118.955 47.550 120.095 ;
        RECT 47.720 118.905 47.975 119.785 ;
        RECT 46.855 118.755 47.595 118.785 ;
        RECT 45.570 118.155 46.100 118.325 ;
        RECT 43.880 117.735 44.230 117.905 ;
        RECT 44.450 117.715 45.400 117.995 ;
        RECT 45.570 117.545 45.760 117.985 ;
        RECT 45.930 117.925 46.100 118.155 ;
        RECT 46.270 118.095 46.510 118.495 ;
        RECT 46.680 118.455 47.595 118.755 ;
        RECT 46.680 118.280 47.005 118.455 ;
        RECT 46.680 117.925 47.000 118.280 ;
        RECT 47.765 118.255 47.975 118.905 ;
        RECT 45.930 117.755 47.000 117.925 ;
        RECT 47.245 117.545 47.550 118.005 ;
        RECT 47.720 117.725 47.975 118.255 ;
        RECT 48.155 118.905 48.410 119.785 ;
        RECT 48.580 118.955 48.885 120.095 ;
        RECT 49.225 119.715 49.555 120.095 ;
        RECT 49.735 119.545 49.905 119.835 ;
        RECT 50.075 119.635 50.325 120.095 ;
        RECT 49.105 119.375 49.905 119.545 ;
        RECT 50.495 119.585 51.365 119.925 ;
        RECT 48.155 118.255 48.365 118.905 ;
        RECT 49.105 118.785 49.275 119.375 ;
        RECT 50.495 119.205 50.665 119.585 ;
        RECT 51.600 119.465 51.770 119.925 ;
        RECT 51.940 119.635 52.310 120.095 ;
        RECT 52.605 119.495 52.775 119.835 ;
        RECT 52.945 119.665 53.275 120.095 ;
        RECT 53.510 119.495 53.680 119.835 ;
        RECT 49.445 119.035 50.665 119.205 ;
        RECT 50.835 119.125 51.295 119.415 ;
        RECT 51.600 119.295 52.160 119.465 ;
        RECT 52.605 119.325 53.680 119.495 ;
        RECT 53.850 119.595 54.530 119.925 ;
        RECT 54.745 119.595 54.995 119.925 ;
        RECT 55.165 119.635 55.415 120.095 ;
        RECT 51.990 119.155 52.160 119.295 ;
        RECT 50.835 119.115 51.800 119.125 ;
        RECT 50.495 118.945 50.665 119.035 ;
        RECT 51.125 118.955 51.800 119.115 ;
        RECT 48.535 118.755 49.275 118.785 ;
        RECT 48.535 118.455 49.450 118.755 ;
        RECT 49.125 118.280 49.450 118.455 ;
        RECT 48.155 117.725 48.410 118.255 ;
        RECT 48.580 117.545 48.885 118.005 ;
        RECT 49.130 117.925 49.450 118.280 ;
        RECT 49.620 118.495 50.160 118.865 ;
        RECT 50.495 118.775 50.900 118.945 ;
        RECT 49.620 118.095 49.860 118.495 ;
        RECT 50.340 118.325 50.560 118.605 ;
        RECT 50.030 118.155 50.560 118.325 ;
        RECT 50.030 117.925 50.200 118.155 ;
        RECT 50.730 117.995 50.900 118.775 ;
        RECT 51.070 118.165 51.420 118.785 ;
        RECT 51.590 118.165 51.800 118.955 ;
        RECT 51.990 118.985 53.490 119.155 ;
        RECT 51.990 118.295 52.160 118.985 ;
        RECT 53.850 118.815 54.020 119.595 ;
        RECT 54.825 119.465 54.995 119.595 ;
        RECT 52.330 118.645 54.020 118.815 ;
        RECT 54.190 119.035 54.655 119.425 ;
        RECT 54.825 119.295 55.220 119.465 ;
        RECT 52.330 118.465 52.500 118.645 ;
        RECT 49.130 117.755 50.200 117.925 ;
        RECT 50.370 117.545 50.560 117.985 ;
        RECT 50.730 117.715 51.680 117.995 ;
        RECT 51.990 117.905 52.250 118.295 ;
        RECT 52.670 118.225 53.460 118.475 ;
        RECT 51.900 117.735 52.250 117.905 ;
        RECT 52.460 117.545 52.790 118.005 ;
        RECT 53.665 117.935 53.835 118.645 ;
        RECT 54.190 118.445 54.360 119.035 ;
        RECT 54.005 118.225 54.360 118.445 ;
        RECT 54.530 118.225 54.880 118.845 ;
        RECT 55.050 117.935 55.220 119.295 ;
        RECT 55.585 119.125 55.910 119.910 ;
        RECT 55.390 118.075 55.850 119.125 ;
        RECT 53.665 117.765 54.520 117.935 ;
        RECT 54.725 117.765 55.220 117.935 ;
        RECT 55.390 117.545 55.720 117.905 ;
        RECT 56.080 117.805 56.250 119.925 ;
        RECT 56.420 119.595 56.750 120.095 ;
        RECT 56.920 119.425 57.175 119.925 ;
        RECT 56.425 119.255 57.175 119.425 ;
        RECT 56.425 118.265 56.655 119.255 ;
        RECT 56.825 118.435 57.175 119.085 ;
        RECT 57.810 118.955 58.080 119.925 ;
        RECT 58.290 119.295 58.570 120.095 ;
        RECT 58.740 119.585 60.395 119.875 ;
        RECT 58.805 119.245 60.395 119.415 ;
        RECT 58.805 119.125 58.975 119.245 ;
        RECT 58.250 118.955 58.975 119.125 ;
        RECT 56.425 118.095 57.175 118.265 ;
        RECT 56.420 117.545 56.750 117.925 ;
        RECT 56.920 117.805 57.175 118.095 ;
        RECT 57.810 118.220 57.980 118.955 ;
        RECT 58.250 118.785 58.420 118.955 ;
        RECT 59.165 118.905 59.880 119.075 ;
        RECT 60.075 118.955 60.395 119.245 ;
        RECT 60.570 118.930 60.860 120.095 ;
        RECT 61.030 119.375 61.490 119.925 ;
        RECT 61.680 119.375 62.010 120.095 ;
        RECT 58.150 118.455 58.420 118.785 ;
        RECT 58.590 118.455 58.995 118.785 ;
        RECT 59.165 118.455 59.875 118.905 ;
        RECT 58.250 118.285 58.420 118.455 ;
        RECT 57.810 117.875 58.080 118.220 ;
        RECT 58.250 118.115 59.860 118.285 ;
        RECT 60.045 118.215 60.395 118.785 ;
        RECT 58.270 117.545 58.650 117.945 ;
        RECT 58.820 117.765 58.990 118.115 ;
        RECT 59.160 117.545 59.490 117.945 ;
        RECT 59.690 117.765 59.860 118.115 ;
        RECT 60.060 117.545 60.390 118.045 ;
        RECT 60.570 117.545 60.860 118.270 ;
        RECT 61.030 118.005 61.280 119.375 ;
        RECT 62.210 119.205 62.510 119.755 ;
        RECT 62.680 119.425 62.960 120.095 ;
        RECT 61.570 119.035 62.510 119.205 ;
        RECT 61.570 118.785 61.740 119.035 ;
        RECT 62.880 118.785 63.145 119.145 ;
        RECT 61.450 118.455 61.740 118.785 ;
        RECT 61.910 118.535 62.250 118.785 ;
        RECT 62.470 118.535 63.145 118.785 ;
        RECT 63.330 118.955 63.600 119.925 ;
        RECT 63.810 119.295 64.090 120.095 ;
        RECT 64.260 119.585 65.915 119.875 ;
        RECT 66.095 119.425 66.350 119.925 ;
        RECT 66.520 119.595 66.850 120.095 ;
        RECT 64.325 119.245 65.915 119.415 ;
        RECT 66.095 119.255 66.845 119.425 ;
        RECT 64.325 119.125 64.495 119.245 ;
        RECT 63.770 118.955 64.495 119.125 ;
        RECT 61.570 118.365 61.740 118.455 ;
        RECT 61.570 118.175 62.960 118.365 ;
        RECT 61.030 117.715 61.590 118.005 ;
        RECT 61.760 117.545 62.010 118.005 ;
        RECT 62.630 117.815 62.960 118.175 ;
        RECT 63.330 118.220 63.500 118.955 ;
        RECT 63.770 118.785 63.940 118.955 ;
        RECT 63.670 118.455 63.940 118.785 ;
        RECT 64.110 118.455 64.515 118.785 ;
        RECT 64.685 118.455 65.395 119.075 ;
        RECT 65.595 118.955 65.915 119.245 ;
        RECT 63.770 118.285 63.940 118.455 ;
        RECT 63.330 117.875 63.600 118.220 ;
        RECT 63.770 118.115 65.380 118.285 ;
        RECT 65.565 118.215 65.915 118.785 ;
        RECT 66.095 118.435 66.445 119.085 ;
        RECT 66.615 118.265 66.845 119.255 ;
        RECT 63.790 117.545 64.170 117.945 ;
        RECT 64.340 117.765 64.510 118.115 ;
        RECT 64.680 117.545 65.010 117.945 ;
        RECT 65.210 117.765 65.380 118.115 ;
        RECT 66.095 118.095 66.845 118.265 ;
        RECT 65.580 117.545 65.910 118.045 ;
        RECT 66.095 117.805 66.350 118.095 ;
        RECT 66.520 117.545 66.850 117.925 ;
        RECT 67.020 117.805 67.190 119.925 ;
        RECT 67.360 119.125 67.685 119.910 ;
        RECT 67.855 119.635 68.105 120.095 ;
        RECT 68.275 119.595 68.525 119.925 ;
        RECT 68.740 119.595 69.420 119.925 ;
        RECT 68.275 119.465 68.445 119.595 ;
        RECT 68.050 119.295 68.445 119.465 ;
        RECT 67.420 118.075 67.880 119.125 ;
        RECT 68.050 117.935 68.220 119.295 ;
        RECT 68.615 119.035 69.080 119.425 ;
        RECT 68.390 118.225 68.740 118.845 ;
        RECT 68.910 118.445 69.080 119.035 ;
        RECT 69.250 118.815 69.420 119.595 ;
        RECT 69.590 119.495 69.760 119.835 ;
        RECT 69.995 119.665 70.325 120.095 ;
        RECT 70.495 119.495 70.665 119.835 ;
        RECT 70.960 119.635 71.330 120.095 ;
        RECT 69.590 119.325 70.665 119.495 ;
        RECT 71.500 119.465 71.670 119.925 ;
        RECT 71.905 119.585 72.775 119.925 ;
        RECT 72.945 119.635 73.195 120.095 ;
        RECT 71.110 119.295 71.670 119.465 ;
        RECT 71.110 119.155 71.280 119.295 ;
        RECT 69.780 118.985 71.280 119.155 ;
        RECT 71.975 119.125 72.435 119.415 ;
        RECT 69.250 118.645 70.940 118.815 ;
        RECT 68.910 118.225 69.265 118.445 ;
        RECT 69.435 117.935 69.605 118.645 ;
        RECT 69.810 118.225 70.600 118.475 ;
        RECT 70.770 118.465 70.940 118.645 ;
        RECT 71.110 118.295 71.280 118.985 ;
        RECT 67.550 117.545 67.880 117.905 ;
        RECT 68.050 117.765 68.545 117.935 ;
        RECT 68.750 117.765 69.605 117.935 ;
        RECT 70.480 117.545 70.810 118.005 ;
        RECT 71.020 117.905 71.280 118.295 ;
        RECT 71.470 119.115 72.435 119.125 ;
        RECT 72.605 119.205 72.775 119.585 ;
        RECT 73.365 119.545 73.535 119.835 ;
        RECT 73.715 119.715 74.045 120.095 ;
        RECT 73.365 119.375 74.165 119.545 ;
        RECT 71.470 118.955 72.145 119.115 ;
        RECT 72.605 119.035 73.825 119.205 ;
        RECT 71.470 118.165 71.680 118.955 ;
        RECT 72.605 118.945 72.775 119.035 ;
        RECT 71.850 118.165 72.200 118.785 ;
        RECT 72.370 118.775 72.775 118.945 ;
        RECT 72.370 117.995 72.540 118.775 ;
        RECT 72.710 118.325 72.930 118.605 ;
        RECT 73.110 118.495 73.650 118.865 ;
        RECT 73.995 118.785 74.165 119.375 ;
        RECT 74.385 118.955 74.690 120.095 ;
        RECT 74.860 118.905 75.115 119.785 ;
        RECT 73.995 118.755 74.735 118.785 ;
        RECT 72.710 118.155 73.240 118.325 ;
        RECT 71.020 117.735 71.370 117.905 ;
        RECT 71.590 117.715 72.540 117.995 ;
        RECT 72.710 117.545 72.900 117.985 ;
        RECT 73.070 117.925 73.240 118.155 ;
        RECT 73.410 118.095 73.650 118.495 ;
        RECT 73.820 118.455 74.735 118.755 ;
        RECT 73.820 118.280 74.145 118.455 ;
        RECT 73.820 117.925 74.140 118.280 ;
        RECT 74.905 118.255 75.115 118.905 ;
        RECT 75.290 119.335 75.805 119.745 ;
        RECT 76.040 119.335 76.210 120.095 ;
        RECT 76.380 119.755 78.410 119.925 ;
        RECT 75.290 118.525 75.630 119.335 ;
        RECT 76.380 119.090 76.550 119.755 ;
        RECT 76.945 119.415 78.070 119.585 ;
        RECT 75.800 118.900 76.550 119.090 ;
        RECT 76.720 119.075 77.730 119.245 ;
        RECT 75.290 118.355 76.520 118.525 ;
        RECT 73.070 117.755 74.140 117.925 ;
        RECT 74.385 117.545 74.690 118.005 ;
        RECT 74.860 117.725 75.115 118.255 ;
        RECT 75.565 117.750 75.810 118.355 ;
        RECT 76.030 117.545 76.540 118.080 ;
        RECT 76.720 117.715 76.910 119.075 ;
        RECT 77.080 118.735 77.355 118.875 ;
        RECT 77.080 118.565 77.360 118.735 ;
        RECT 77.080 117.715 77.355 118.565 ;
        RECT 77.560 118.275 77.730 119.075 ;
        RECT 77.900 118.285 78.070 119.415 ;
        RECT 78.240 118.785 78.410 119.755 ;
        RECT 78.580 118.955 78.750 120.095 ;
        RECT 78.920 118.955 79.255 119.925 ;
        RECT 78.240 118.455 78.435 118.785 ;
        RECT 78.660 118.455 78.915 118.785 ;
        RECT 78.660 118.285 78.830 118.455 ;
        RECT 79.085 118.285 79.255 118.955 ;
        RECT 77.900 118.115 78.830 118.285 ;
        RECT 77.900 118.080 78.075 118.115 ;
        RECT 77.545 117.715 78.075 118.080 ;
        RECT 78.500 117.545 78.830 117.945 ;
        RECT 79.000 117.715 79.255 118.285 ;
        RECT 79.890 119.125 80.200 119.925 ;
        RECT 80.370 119.295 80.680 120.095 ;
        RECT 80.850 119.465 81.110 119.925 ;
        RECT 81.280 119.635 81.535 120.095 ;
        RECT 81.710 119.465 81.970 119.925 ;
        RECT 80.850 119.295 81.970 119.465 ;
        RECT 79.890 118.955 80.920 119.125 ;
        RECT 79.890 118.045 80.060 118.955 ;
        RECT 80.230 118.215 80.580 118.785 ;
        RECT 80.750 118.705 80.920 118.955 ;
        RECT 81.710 119.045 81.970 119.295 ;
        RECT 82.140 119.225 82.425 120.095 ;
        RECT 81.710 118.875 82.465 119.045 ;
        RECT 80.750 118.535 81.890 118.705 ;
        RECT 82.060 118.365 82.465 118.875 ;
        RECT 80.815 118.195 82.465 118.365 ;
        RECT 82.650 118.955 82.990 119.925 ;
        RECT 83.160 118.955 83.330 120.095 ;
        RECT 83.600 119.295 83.850 120.095 ;
        RECT 84.495 119.125 84.825 119.925 ;
        RECT 85.125 119.295 85.455 120.095 ;
        RECT 85.625 119.125 85.955 119.925 ;
        RECT 83.520 118.955 85.955 119.125 ;
        RECT 82.650 118.345 82.825 118.955 ;
        RECT 83.520 118.705 83.690 118.955 ;
        RECT 82.995 118.535 83.690 118.705 ;
        RECT 83.865 118.535 84.285 118.735 ;
        RECT 84.455 118.535 84.785 118.735 ;
        RECT 84.955 118.535 85.285 118.735 ;
        RECT 79.890 117.715 80.190 118.045 ;
        RECT 80.360 117.545 80.635 118.025 ;
        RECT 80.815 117.805 81.110 118.195 ;
        RECT 81.280 117.545 81.535 118.025 ;
        RECT 81.710 117.805 81.970 118.195 ;
        RECT 82.140 117.545 82.420 118.025 ;
        RECT 82.650 117.715 82.990 118.345 ;
        RECT 83.160 117.545 83.410 118.345 ;
        RECT 83.600 118.195 84.825 118.365 ;
        RECT 83.600 117.715 83.930 118.195 ;
        RECT 84.100 117.545 84.325 118.005 ;
        RECT 84.495 117.715 84.825 118.195 ;
        RECT 85.455 118.325 85.625 118.955 ;
        RECT 86.330 118.930 86.620 120.095 ;
        RECT 86.830 118.955 87.060 120.095 ;
        RECT 87.230 118.945 87.560 119.925 ;
        RECT 87.730 118.955 87.940 120.095 ;
        RECT 88.170 118.955 88.510 119.925 ;
        RECT 88.680 118.955 88.850 120.095 ;
        RECT 89.120 119.295 89.370 120.095 ;
        RECT 90.015 119.125 90.345 119.925 ;
        RECT 90.645 119.295 90.975 120.095 ;
        RECT 91.145 119.125 91.475 119.925 ;
        RECT 89.040 118.955 91.475 119.125 ;
        RECT 91.850 119.335 92.365 119.745 ;
        RECT 92.600 119.335 92.770 120.095 ;
        RECT 92.940 119.755 94.970 119.925 ;
        RECT 85.810 118.535 86.160 118.785 ;
        RECT 86.810 118.535 87.140 118.785 ;
        RECT 85.455 117.715 85.955 118.325 ;
        RECT 86.330 117.545 86.620 118.270 ;
        RECT 86.830 117.545 87.060 118.365 ;
        RECT 87.310 118.345 87.560 118.945 ;
        RECT 88.170 118.905 88.400 118.955 ;
        RECT 87.230 117.715 87.560 118.345 ;
        RECT 87.730 117.545 87.940 118.365 ;
        RECT 88.170 118.345 88.345 118.905 ;
        RECT 89.040 118.705 89.210 118.955 ;
        RECT 88.515 118.535 89.210 118.705 ;
        RECT 89.385 118.535 89.805 118.735 ;
        RECT 89.975 118.535 90.305 118.735 ;
        RECT 90.475 118.535 90.805 118.735 ;
        RECT 88.170 117.715 88.510 118.345 ;
        RECT 88.680 117.545 88.930 118.345 ;
        RECT 89.120 118.195 90.345 118.365 ;
        RECT 89.120 117.715 89.450 118.195 ;
        RECT 89.620 117.545 89.845 118.005 ;
        RECT 90.015 117.715 90.345 118.195 ;
        RECT 90.975 118.325 91.145 118.955 ;
        RECT 91.330 118.535 91.680 118.785 ;
        RECT 91.850 118.525 92.190 119.335 ;
        RECT 92.940 119.090 93.110 119.755 ;
        RECT 93.505 119.415 94.630 119.585 ;
        RECT 92.360 118.900 93.110 119.090 ;
        RECT 93.280 119.075 94.290 119.245 ;
        RECT 91.850 118.355 93.080 118.525 ;
        RECT 90.975 117.715 91.475 118.325 ;
        RECT 92.125 117.750 92.370 118.355 ;
        RECT 92.590 117.545 93.100 118.080 ;
        RECT 93.280 117.715 93.470 119.075 ;
        RECT 93.640 118.055 93.915 118.875 ;
        RECT 94.120 118.275 94.290 119.075 ;
        RECT 94.460 118.285 94.630 119.415 ;
        RECT 94.800 118.785 94.970 119.755 ;
        RECT 95.140 118.955 95.310 120.095 ;
        RECT 95.480 118.955 95.815 119.925 ;
        RECT 95.995 119.425 96.250 119.925 ;
        RECT 96.420 119.595 96.750 120.095 ;
        RECT 95.995 119.255 96.745 119.425 ;
        RECT 94.800 118.455 94.995 118.785 ;
        RECT 95.220 118.455 95.475 118.785 ;
        RECT 95.220 118.285 95.390 118.455 ;
        RECT 95.645 118.285 95.815 118.955 ;
        RECT 95.995 118.435 96.345 119.085 ;
        RECT 94.460 118.115 95.390 118.285 ;
        RECT 94.460 118.080 94.635 118.115 ;
        RECT 93.640 117.885 93.920 118.055 ;
        RECT 93.640 117.715 93.915 117.885 ;
        RECT 94.105 117.715 94.635 118.080 ;
        RECT 95.060 117.545 95.390 117.945 ;
        RECT 95.560 117.715 95.815 118.285 ;
        RECT 96.515 118.265 96.745 119.255 ;
        RECT 95.995 118.095 96.745 118.265 ;
        RECT 95.995 117.805 96.250 118.095 ;
        RECT 96.420 117.545 96.750 117.925 ;
        RECT 96.920 117.805 97.090 119.925 ;
        RECT 97.260 119.125 97.585 119.910 ;
        RECT 97.755 119.635 98.005 120.095 ;
        RECT 98.175 119.595 98.425 119.925 ;
        RECT 98.640 119.595 99.320 119.925 ;
        RECT 98.175 119.465 98.345 119.595 ;
        RECT 97.950 119.295 98.345 119.465 ;
        RECT 97.320 118.075 97.780 119.125 ;
        RECT 97.950 117.935 98.120 119.295 ;
        RECT 98.515 119.035 98.980 119.425 ;
        RECT 98.290 118.225 98.640 118.845 ;
        RECT 98.810 118.445 98.980 119.035 ;
        RECT 99.150 118.815 99.320 119.595 ;
        RECT 99.490 119.495 99.660 119.835 ;
        RECT 99.895 119.665 100.225 120.095 ;
        RECT 100.395 119.495 100.565 119.835 ;
        RECT 100.860 119.635 101.230 120.095 ;
        RECT 99.490 119.325 100.565 119.495 ;
        RECT 101.400 119.465 101.570 119.925 ;
        RECT 101.805 119.585 102.675 119.925 ;
        RECT 102.845 119.635 103.095 120.095 ;
        RECT 101.010 119.295 101.570 119.465 ;
        RECT 101.010 119.155 101.180 119.295 ;
        RECT 99.680 118.985 101.180 119.155 ;
        RECT 101.875 119.125 102.335 119.415 ;
        RECT 99.150 118.645 100.840 118.815 ;
        RECT 98.810 118.225 99.165 118.445 ;
        RECT 99.335 117.935 99.505 118.645 ;
        RECT 99.710 118.225 100.500 118.475 ;
        RECT 100.670 118.465 100.840 118.645 ;
        RECT 101.010 118.295 101.180 118.985 ;
        RECT 97.450 117.545 97.780 117.905 ;
        RECT 97.950 117.765 98.445 117.935 ;
        RECT 98.650 117.765 99.505 117.935 ;
        RECT 100.380 117.545 100.710 118.005 ;
        RECT 100.920 117.905 101.180 118.295 ;
        RECT 101.370 119.115 102.335 119.125 ;
        RECT 102.505 119.205 102.675 119.585 ;
        RECT 103.265 119.545 103.435 119.835 ;
        RECT 103.615 119.715 103.945 120.095 ;
        RECT 103.265 119.375 104.065 119.545 ;
        RECT 101.370 118.955 102.045 119.115 ;
        RECT 102.505 119.035 103.725 119.205 ;
        RECT 101.370 118.165 101.580 118.955 ;
        RECT 102.505 118.945 102.675 119.035 ;
        RECT 101.750 118.165 102.100 118.785 ;
        RECT 102.270 118.775 102.675 118.945 ;
        RECT 102.270 117.995 102.440 118.775 ;
        RECT 102.610 118.325 102.830 118.605 ;
        RECT 103.010 118.495 103.550 118.865 ;
        RECT 103.895 118.785 104.065 119.375 ;
        RECT 104.285 118.955 104.590 120.095 ;
        RECT 104.760 118.905 105.015 119.785 ;
        RECT 105.655 119.660 111.000 120.095 ;
        RECT 103.895 118.755 104.635 118.785 ;
        RECT 102.610 118.155 103.140 118.325 ;
        RECT 100.920 117.735 101.270 117.905 ;
        RECT 101.490 117.715 102.440 117.995 ;
        RECT 102.610 117.545 102.800 117.985 ;
        RECT 102.970 117.925 103.140 118.155 ;
        RECT 103.310 118.095 103.550 118.495 ;
        RECT 103.720 118.455 104.635 118.755 ;
        RECT 103.720 118.280 104.045 118.455 ;
        RECT 103.720 117.925 104.040 118.280 ;
        RECT 104.805 118.255 105.015 118.905 ;
        RECT 107.245 118.410 107.595 119.660 ;
        RECT 111.170 119.005 112.380 120.095 ;
        RECT 102.970 117.755 104.040 117.925 ;
        RECT 104.285 117.545 104.590 118.005 ;
        RECT 104.760 117.725 105.015 118.255 ;
        RECT 109.075 118.090 109.415 118.920 ;
        RECT 111.170 118.465 111.690 119.005 ;
        RECT 111.860 118.295 112.380 118.835 ;
        RECT 105.655 117.545 111.000 118.090 ;
        RECT 111.170 117.545 112.380 118.295 ;
        RECT 18.165 117.375 112.465 117.545 ;
        RECT 18.250 116.625 19.460 117.375 ;
        RECT 18.250 116.085 18.770 116.625 ;
        RECT 20.090 116.605 21.760 117.375 ;
        RECT 21.930 116.650 22.220 117.375 ;
        RECT 23.160 116.905 23.330 117.375 ;
        RECT 23.500 116.725 23.830 117.205 ;
        RECT 24.000 116.905 24.170 117.375 ;
        RECT 24.340 116.725 24.670 117.205 ;
        RECT 18.940 115.915 19.460 116.455 ;
        RECT 18.250 114.825 19.460 115.915 ;
        RECT 20.090 115.915 20.840 116.435 ;
        RECT 21.010 116.085 21.760 116.605 ;
        RECT 22.905 116.555 24.670 116.725 ;
        RECT 24.840 116.565 25.010 117.375 ;
        RECT 25.210 116.995 26.280 117.165 ;
        RECT 25.210 116.640 25.530 116.995 ;
        RECT 22.905 116.005 23.315 116.555 ;
        RECT 25.205 116.385 25.530 116.640 ;
        RECT 23.500 116.175 25.530 116.385 ;
        RECT 25.185 116.165 25.530 116.175 ;
        RECT 25.700 116.425 25.940 116.825 ;
        RECT 26.110 116.765 26.280 116.995 ;
        RECT 26.450 116.935 26.640 117.375 ;
        RECT 26.810 116.925 27.760 117.205 ;
        RECT 27.980 117.015 28.330 117.185 ;
        RECT 26.110 116.595 26.640 116.765 ;
        RECT 20.090 114.825 21.760 115.915 ;
        RECT 21.930 114.825 22.220 115.990 ;
        RECT 22.905 115.835 24.630 116.005 ;
        RECT 23.160 114.825 23.330 115.665 ;
        RECT 23.540 114.995 23.790 115.835 ;
        RECT 24.000 114.825 24.170 115.665 ;
        RECT 24.340 114.995 24.630 115.835 ;
        RECT 24.840 114.825 25.010 115.885 ;
        RECT 25.185 115.545 25.355 116.165 ;
        RECT 25.700 116.055 26.240 116.425 ;
        RECT 26.420 116.315 26.640 116.595 ;
        RECT 26.810 116.145 26.980 116.925 ;
        RECT 26.575 115.975 26.980 116.145 ;
        RECT 27.150 116.135 27.500 116.755 ;
        RECT 26.575 115.885 26.745 115.975 ;
        RECT 27.670 115.965 27.880 116.755 ;
        RECT 25.525 115.715 26.745 115.885 ;
        RECT 27.205 115.805 27.880 115.965 ;
        RECT 25.185 115.375 25.985 115.545 ;
        RECT 25.305 114.825 25.635 115.205 ;
        RECT 25.815 115.085 25.985 115.375 ;
        RECT 26.575 115.335 26.745 115.715 ;
        RECT 26.915 115.795 27.880 115.805 ;
        RECT 28.070 116.625 28.330 117.015 ;
        RECT 28.540 116.915 28.870 117.375 ;
        RECT 29.745 116.985 30.600 117.155 ;
        RECT 30.805 116.985 31.300 117.155 ;
        RECT 31.470 117.015 31.800 117.375 ;
        RECT 28.070 115.935 28.240 116.625 ;
        RECT 28.410 116.275 28.580 116.455 ;
        RECT 28.750 116.445 29.540 116.695 ;
        RECT 29.745 116.275 29.915 116.985 ;
        RECT 30.085 116.475 30.440 116.695 ;
        RECT 28.410 116.105 30.100 116.275 ;
        RECT 26.915 115.505 27.375 115.795 ;
        RECT 28.070 115.765 29.570 115.935 ;
        RECT 28.070 115.625 28.240 115.765 ;
        RECT 27.680 115.455 28.240 115.625 ;
        RECT 26.155 114.825 26.405 115.285 ;
        RECT 26.575 114.995 27.445 115.335 ;
        RECT 27.680 114.995 27.850 115.455 ;
        RECT 28.685 115.425 29.760 115.595 ;
        RECT 28.020 114.825 28.390 115.285 ;
        RECT 28.685 115.085 28.855 115.425 ;
        RECT 29.025 114.825 29.355 115.255 ;
        RECT 29.590 115.085 29.760 115.425 ;
        RECT 29.930 115.325 30.100 116.105 ;
        RECT 30.270 115.885 30.440 116.475 ;
        RECT 30.610 116.075 30.960 116.695 ;
        RECT 30.270 115.495 30.735 115.885 ;
        RECT 31.130 115.625 31.300 116.985 ;
        RECT 31.470 115.795 31.930 116.845 ;
        RECT 30.905 115.455 31.300 115.625 ;
        RECT 30.905 115.325 31.075 115.455 ;
        RECT 29.930 114.995 30.610 115.325 ;
        RECT 30.825 114.995 31.075 115.325 ;
        RECT 31.245 114.825 31.495 115.285 ;
        RECT 31.665 115.010 31.990 115.795 ;
        RECT 32.160 114.995 32.330 117.115 ;
        RECT 32.500 116.995 32.830 117.375 ;
        RECT 33.000 116.825 33.255 117.115 ;
        RECT 33.490 116.895 33.770 117.375 ;
        RECT 32.505 116.655 33.255 116.825 ;
        RECT 33.940 116.725 34.200 117.115 ;
        RECT 34.375 116.895 34.630 117.375 ;
        RECT 34.800 116.725 35.095 117.115 ;
        RECT 35.275 116.895 35.550 117.375 ;
        RECT 35.720 116.875 36.020 117.205 ;
        RECT 32.505 115.665 32.735 116.655 ;
        RECT 33.445 116.555 35.095 116.725 ;
        RECT 32.905 115.835 33.255 116.485 ;
        RECT 33.445 116.045 33.850 116.555 ;
        RECT 34.020 116.215 35.160 116.385 ;
        RECT 33.445 115.875 34.200 116.045 ;
        RECT 32.505 115.495 33.255 115.665 ;
        RECT 32.500 114.825 32.830 115.325 ;
        RECT 33.000 114.995 33.255 115.495 ;
        RECT 33.485 114.825 33.770 115.695 ;
        RECT 33.940 115.625 34.200 115.875 ;
        RECT 34.990 115.965 35.160 116.215 ;
        RECT 35.330 116.135 35.680 116.705 ;
        RECT 35.850 115.965 36.020 116.875 ;
        RECT 36.305 116.745 36.590 117.205 ;
        RECT 36.760 116.915 37.030 117.375 ;
        RECT 36.305 116.575 37.260 116.745 ;
        RECT 34.990 115.795 36.020 115.965 ;
        RECT 36.190 115.845 36.880 116.405 ;
        RECT 34.410 115.625 34.580 115.675 ;
        RECT 33.940 115.455 35.060 115.625 ;
        RECT 33.940 114.995 34.200 115.455 ;
        RECT 34.375 114.825 34.630 115.285 ;
        RECT 34.800 114.995 35.060 115.455 ;
        RECT 35.230 114.825 35.540 115.625 ;
        RECT 35.710 114.995 36.020 115.795 ;
        RECT 37.050 115.675 37.260 116.575 ;
        RECT 36.305 115.455 37.260 115.675 ;
        RECT 37.430 116.405 37.830 117.205 ;
        RECT 38.020 116.745 38.300 117.205 ;
        RECT 38.820 116.915 39.145 117.375 ;
        RECT 38.020 116.575 39.145 116.745 ;
        RECT 39.315 116.635 39.700 117.205 ;
        RECT 38.695 116.465 39.145 116.575 ;
        RECT 37.430 115.845 38.525 116.405 ;
        RECT 38.695 116.135 39.250 116.465 ;
        RECT 36.305 114.995 36.590 115.455 ;
        RECT 36.760 114.825 37.030 115.285 ;
        RECT 37.430 114.995 37.830 115.845 ;
        RECT 38.695 115.675 39.145 116.135 ;
        RECT 39.420 115.965 39.700 116.635 ;
        RECT 39.985 116.745 40.270 117.205 ;
        RECT 40.440 116.915 40.710 117.375 ;
        RECT 39.985 116.575 40.940 116.745 ;
        RECT 38.020 115.455 39.145 115.675 ;
        RECT 38.020 114.995 38.300 115.455 ;
        RECT 38.820 114.825 39.145 115.285 ;
        RECT 39.315 114.995 39.700 115.965 ;
        RECT 39.870 115.845 40.560 116.405 ;
        RECT 40.730 115.675 40.940 116.575 ;
        RECT 39.985 115.455 40.940 115.675 ;
        RECT 41.110 116.405 41.510 117.205 ;
        RECT 41.700 116.745 41.980 117.205 ;
        RECT 42.500 116.915 42.825 117.375 ;
        RECT 41.700 116.575 42.825 116.745 ;
        RECT 42.995 116.635 43.380 117.205 ;
        RECT 42.375 116.465 42.825 116.575 ;
        RECT 41.110 115.845 42.205 116.405 ;
        RECT 42.375 116.135 42.930 116.465 ;
        RECT 39.985 114.995 40.270 115.455 ;
        RECT 40.440 114.825 40.710 115.285 ;
        RECT 41.110 114.995 41.510 115.845 ;
        RECT 42.375 115.675 42.825 116.135 ;
        RECT 43.100 115.965 43.380 116.635 ;
        RECT 41.700 115.455 42.825 115.675 ;
        RECT 41.700 114.995 41.980 115.455 ;
        RECT 42.500 114.825 42.825 115.285 ;
        RECT 42.995 114.995 43.380 115.965 ;
        RECT 43.550 116.635 43.935 117.205 ;
        RECT 44.105 116.915 44.430 117.375 ;
        RECT 44.950 116.745 45.230 117.205 ;
        RECT 43.550 115.965 43.830 116.635 ;
        RECT 44.105 116.575 45.230 116.745 ;
        RECT 44.105 116.465 44.555 116.575 ;
        RECT 44.000 116.135 44.555 116.465 ;
        RECT 45.420 116.405 45.820 117.205 ;
        RECT 46.220 116.915 46.490 117.375 ;
        RECT 46.660 116.745 46.945 117.205 ;
        RECT 43.550 114.995 43.935 115.965 ;
        RECT 44.105 115.675 44.555 116.135 ;
        RECT 44.725 115.845 45.820 116.405 ;
        RECT 44.105 115.455 45.230 115.675 ;
        RECT 44.105 114.825 44.430 115.285 ;
        RECT 44.950 114.995 45.230 115.455 ;
        RECT 45.420 114.995 45.820 115.845 ;
        RECT 45.990 116.575 46.945 116.745 ;
        RECT 47.690 116.650 47.980 117.375 ;
        RECT 48.150 116.575 48.490 117.205 ;
        RECT 48.660 116.575 48.910 117.375 ;
        RECT 49.100 116.725 49.430 117.205 ;
        RECT 49.600 116.915 49.825 117.375 ;
        RECT 49.995 116.725 50.325 117.205 ;
        RECT 45.990 115.675 46.200 116.575 ;
        RECT 46.370 115.845 47.060 116.405 ;
        RECT 45.990 115.455 46.945 115.675 ;
        RECT 46.220 114.825 46.490 115.285 ;
        RECT 46.660 114.995 46.945 115.455 ;
        RECT 47.690 114.825 47.980 115.990 ;
        RECT 48.150 115.965 48.325 116.575 ;
        RECT 49.100 116.555 50.325 116.725 ;
        RECT 50.955 116.595 51.455 117.205 ;
        RECT 48.495 116.215 49.190 116.385 ;
        RECT 49.020 115.965 49.190 116.215 ;
        RECT 49.365 116.185 49.785 116.385 ;
        RECT 49.955 116.185 50.285 116.385 ;
        RECT 50.455 116.185 50.785 116.385 ;
        RECT 50.955 115.965 51.125 116.595 ;
        RECT 51.890 116.555 52.100 117.375 ;
        RECT 52.270 116.575 52.600 117.205 ;
        RECT 51.310 116.135 51.660 116.385 ;
        RECT 52.270 115.975 52.520 116.575 ;
        RECT 52.770 116.555 53.000 117.375 ;
        RECT 53.210 116.605 56.720 117.375 ;
        RECT 56.980 116.825 57.150 117.115 ;
        RECT 57.320 116.995 57.650 117.375 ;
        RECT 56.980 116.655 57.645 116.825 ;
        RECT 52.690 116.135 53.020 116.385 ;
        RECT 48.150 114.995 48.490 115.965 ;
        RECT 48.660 114.825 48.830 115.965 ;
        RECT 49.020 115.795 51.455 115.965 ;
        RECT 49.100 114.825 49.350 115.625 ;
        RECT 49.995 114.995 50.325 115.795 ;
        RECT 50.625 114.825 50.955 115.625 ;
        RECT 51.125 114.995 51.455 115.795 ;
        RECT 51.890 114.825 52.100 115.965 ;
        RECT 52.270 114.995 52.600 115.975 ;
        RECT 52.770 114.825 53.000 115.965 ;
        RECT 53.210 115.915 54.900 116.435 ;
        RECT 55.070 116.085 56.720 116.605 ;
        RECT 53.210 114.825 56.720 115.915 ;
        RECT 56.895 115.835 57.245 116.485 ;
        RECT 57.415 115.665 57.645 116.655 ;
        RECT 56.980 115.495 57.645 115.665 ;
        RECT 56.980 114.995 57.150 115.495 ;
        RECT 57.320 114.825 57.650 115.325 ;
        RECT 57.820 114.995 58.045 117.115 ;
        RECT 58.260 116.995 58.590 117.375 ;
        RECT 58.760 116.825 58.930 117.155 ;
        RECT 59.230 116.995 60.245 117.195 ;
        RECT 58.235 116.635 58.930 116.825 ;
        RECT 58.235 115.665 58.405 116.635 ;
        RECT 58.575 115.835 58.985 116.455 ;
        RECT 59.155 115.885 59.375 116.755 ;
        RECT 59.555 116.445 59.905 116.815 ;
        RECT 60.075 116.265 60.245 116.995 ;
        RECT 60.415 116.935 60.825 117.375 ;
        RECT 61.115 116.735 61.365 117.165 ;
        RECT 61.565 116.915 61.885 117.375 ;
        RECT 62.445 116.985 63.295 117.155 ;
        RECT 60.415 116.395 60.825 116.725 ;
        RECT 61.115 116.395 61.535 116.735 ;
        RECT 59.825 116.225 60.245 116.265 ;
        RECT 59.825 116.055 61.175 116.225 ;
        RECT 58.235 115.495 58.930 115.665 ;
        RECT 59.155 115.505 59.655 115.885 ;
        RECT 58.260 114.825 58.590 115.325 ;
        RECT 58.760 114.995 58.930 115.495 ;
        RECT 59.825 115.210 59.995 116.055 ;
        RECT 60.925 115.895 61.175 116.055 ;
        RECT 60.165 115.625 60.415 115.885 ;
        RECT 61.345 115.625 61.535 116.395 ;
        RECT 60.165 115.375 61.535 115.625 ;
        RECT 61.705 116.565 62.955 116.735 ;
        RECT 61.705 115.805 61.875 116.565 ;
        RECT 62.625 116.445 62.955 116.565 ;
        RECT 62.045 115.985 62.225 116.395 ;
        RECT 63.125 116.225 63.295 116.985 ;
        RECT 63.495 116.895 64.155 117.375 ;
        RECT 64.335 116.780 64.655 117.110 ;
        RECT 63.485 116.455 64.145 116.725 ;
        RECT 63.485 116.395 63.815 116.455 ;
        RECT 63.965 116.225 64.295 116.285 ;
        RECT 62.395 116.055 64.295 116.225 ;
        RECT 61.705 115.495 62.225 115.805 ;
        RECT 62.395 115.545 62.565 116.055 ;
        RECT 64.465 115.885 64.655 116.780 ;
        RECT 62.735 115.715 64.655 115.885 ;
        RECT 64.335 115.695 64.655 115.715 ;
        RECT 64.855 116.465 65.105 117.115 ;
        RECT 65.285 116.915 65.570 117.375 ;
        RECT 65.750 116.665 66.005 117.195 ;
        RECT 64.855 116.135 65.655 116.465 ;
        RECT 62.395 115.375 63.605 115.545 ;
        RECT 59.165 115.040 59.995 115.210 ;
        RECT 60.235 114.825 60.615 115.205 ;
        RECT 60.795 115.085 60.965 115.375 ;
        RECT 62.395 115.295 62.565 115.375 ;
        RECT 61.135 114.825 61.465 115.205 ;
        RECT 61.935 115.045 62.565 115.295 ;
        RECT 62.745 114.825 63.165 115.205 ;
        RECT 63.365 115.085 63.605 115.375 ;
        RECT 63.835 114.825 64.165 115.515 ;
        RECT 64.335 115.085 64.505 115.695 ;
        RECT 64.855 115.545 65.105 116.135 ;
        RECT 65.825 115.805 66.005 116.665 ;
        RECT 64.775 115.035 65.105 115.545 ;
        RECT 65.285 114.825 65.570 115.625 ;
        RECT 65.750 115.335 66.005 115.805 ;
        RECT 67.010 116.575 67.350 117.205 ;
        RECT 67.520 116.575 67.770 117.375 ;
        RECT 67.960 116.725 68.290 117.205 ;
        RECT 68.460 116.915 68.685 117.375 ;
        RECT 68.855 116.725 69.185 117.205 ;
        RECT 67.010 116.525 67.240 116.575 ;
        RECT 67.960 116.555 69.185 116.725 ;
        RECT 69.815 116.595 70.315 117.205 ;
        RECT 67.010 115.965 67.185 116.525 ;
        RECT 67.355 116.215 68.050 116.385 ;
        RECT 67.880 115.965 68.050 116.215 ;
        RECT 68.225 116.185 68.645 116.385 ;
        RECT 68.815 116.185 69.145 116.385 ;
        RECT 69.315 116.185 69.645 116.385 ;
        RECT 69.815 115.965 69.985 116.595 ;
        RECT 70.730 116.555 70.960 117.375 ;
        RECT 71.130 116.575 71.460 117.205 ;
        RECT 70.170 116.135 70.520 116.385 ;
        RECT 70.710 116.135 71.040 116.385 ;
        RECT 71.210 115.975 71.460 116.575 ;
        RECT 71.630 116.555 71.840 117.375 ;
        RECT 72.110 116.555 72.340 117.375 ;
        RECT 72.510 116.575 72.840 117.205 ;
        RECT 72.090 116.135 72.420 116.385 ;
        RECT 72.590 115.975 72.840 116.575 ;
        RECT 73.010 116.555 73.220 117.375 ;
        RECT 73.450 116.650 73.740 117.375 ;
        RECT 74.835 116.825 75.090 117.115 ;
        RECT 75.260 116.995 75.590 117.375 ;
        RECT 74.835 116.655 75.585 116.825 ;
        RECT 65.750 115.165 66.090 115.335 ;
        RECT 65.750 115.135 66.005 115.165 ;
        RECT 67.010 114.995 67.350 115.965 ;
        RECT 67.520 114.825 67.690 115.965 ;
        RECT 67.880 115.795 70.315 115.965 ;
        RECT 67.960 114.825 68.210 115.625 ;
        RECT 68.855 114.995 69.185 115.795 ;
        RECT 69.485 114.825 69.815 115.625 ;
        RECT 69.985 114.995 70.315 115.795 ;
        RECT 70.730 114.825 70.960 115.965 ;
        RECT 71.130 114.995 71.460 115.975 ;
        RECT 71.630 114.825 71.840 115.965 ;
        RECT 72.110 114.825 72.340 115.965 ;
        RECT 72.510 114.995 72.840 115.975 ;
        RECT 73.010 114.825 73.220 115.965 ;
        RECT 73.450 114.825 73.740 115.990 ;
        RECT 74.835 115.835 75.185 116.485 ;
        RECT 75.355 115.665 75.585 116.655 ;
        RECT 74.835 115.495 75.585 115.665 ;
        RECT 74.835 114.995 75.090 115.495 ;
        RECT 75.260 114.825 75.590 115.325 ;
        RECT 75.760 114.995 75.930 117.115 ;
        RECT 76.290 117.015 76.620 117.375 ;
        RECT 76.790 116.985 77.285 117.155 ;
        RECT 77.490 116.985 78.345 117.155 ;
        RECT 76.160 115.795 76.620 116.845 ;
        RECT 76.100 115.010 76.425 115.795 ;
        RECT 76.790 115.625 76.960 116.985 ;
        RECT 77.130 116.075 77.480 116.695 ;
        RECT 77.650 116.475 78.005 116.695 ;
        RECT 77.650 115.885 77.820 116.475 ;
        RECT 78.175 116.275 78.345 116.985 ;
        RECT 79.220 116.915 79.550 117.375 ;
        RECT 79.760 117.015 80.110 117.185 ;
        RECT 78.550 116.445 79.340 116.695 ;
        RECT 79.760 116.625 80.020 117.015 ;
        RECT 80.330 116.925 81.280 117.205 ;
        RECT 81.450 116.935 81.640 117.375 ;
        RECT 81.810 116.995 82.880 117.165 ;
        RECT 79.510 116.275 79.680 116.455 ;
        RECT 76.790 115.455 77.185 115.625 ;
        RECT 77.355 115.495 77.820 115.885 ;
        RECT 77.990 116.105 79.680 116.275 ;
        RECT 77.015 115.325 77.185 115.455 ;
        RECT 77.990 115.325 78.160 116.105 ;
        RECT 79.850 115.935 80.020 116.625 ;
        RECT 78.520 115.765 80.020 115.935 ;
        RECT 80.210 115.965 80.420 116.755 ;
        RECT 80.590 116.135 80.940 116.755 ;
        RECT 81.110 116.145 81.280 116.925 ;
        RECT 81.810 116.765 81.980 116.995 ;
        RECT 81.450 116.595 81.980 116.765 ;
        RECT 81.450 116.315 81.670 116.595 ;
        RECT 82.150 116.425 82.390 116.825 ;
        RECT 81.110 115.975 81.515 116.145 ;
        RECT 81.850 116.055 82.390 116.425 ;
        RECT 82.560 116.640 82.880 116.995 ;
        RECT 83.125 116.915 83.430 117.375 ;
        RECT 83.600 116.665 83.855 117.195 ;
        RECT 82.560 116.465 82.885 116.640 ;
        RECT 82.560 116.165 83.475 116.465 ;
        RECT 82.735 116.135 83.475 116.165 ;
        RECT 80.210 115.805 80.885 115.965 ;
        RECT 81.345 115.885 81.515 115.975 ;
        RECT 80.210 115.795 81.175 115.805 ;
        RECT 79.850 115.625 80.020 115.765 ;
        RECT 76.595 114.825 76.845 115.285 ;
        RECT 77.015 114.995 77.265 115.325 ;
        RECT 77.480 114.995 78.160 115.325 ;
        RECT 78.330 115.425 79.405 115.595 ;
        RECT 79.850 115.455 80.410 115.625 ;
        RECT 80.715 115.505 81.175 115.795 ;
        RECT 81.345 115.715 82.565 115.885 ;
        RECT 78.330 115.085 78.500 115.425 ;
        RECT 78.735 114.825 79.065 115.255 ;
        RECT 79.235 115.085 79.405 115.425 ;
        RECT 79.700 114.825 80.070 115.285 ;
        RECT 80.240 114.995 80.410 115.455 ;
        RECT 81.345 115.335 81.515 115.715 ;
        RECT 82.735 115.545 82.905 116.135 ;
        RECT 83.645 116.015 83.855 116.665 ;
        RECT 85.065 116.745 85.350 117.205 ;
        RECT 85.520 116.915 85.790 117.375 ;
        RECT 85.065 116.575 86.020 116.745 ;
        RECT 80.645 114.995 81.515 115.335 ;
        RECT 82.105 115.375 82.905 115.545 ;
        RECT 81.685 114.825 81.935 115.285 ;
        RECT 82.105 115.085 82.275 115.375 ;
        RECT 82.455 114.825 82.785 115.205 ;
        RECT 83.125 114.825 83.430 115.965 ;
        RECT 83.600 115.135 83.855 116.015 ;
        RECT 84.950 115.845 85.640 116.405 ;
        RECT 85.810 115.675 86.020 116.575 ;
        RECT 85.065 115.455 86.020 115.675 ;
        RECT 86.190 116.405 86.590 117.205 ;
        RECT 86.780 116.745 87.060 117.205 ;
        RECT 87.580 116.915 87.905 117.375 ;
        RECT 86.780 116.575 87.905 116.745 ;
        RECT 88.075 116.635 88.460 117.205 ;
        RECT 87.455 116.465 87.905 116.575 ;
        RECT 86.190 115.845 87.285 116.405 ;
        RECT 87.455 116.135 88.010 116.465 ;
        RECT 85.065 114.995 85.350 115.455 ;
        RECT 85.520 114.825 85.790 115.285 ;
        RECT 86.190 114.995 86.590 115.845 ;
        RECT 87.455 115.675 87.905 116.135 ;
        RECT 88.180 115.965 88.460 116.635 ;
        RECT 88.630 116.625 89.840 117.375 ;
        RECT 90.020 116.875 90.350 117.375 ;
        RECT 90.550 116.805 90.720 117.155 ;
        RECT 90.920 116.975 91.250 117.375 ;
        RECT 91.420 116.805 91.590 117.155 ;
        RECT 91.760 116.975 92.140 117.375 ;
        RECT 86.780 115.455 87.905 115.675 ;
        RECT 86.780 114.995 87.060 115.455 ;
        RECT 87.580 114.825 87.905 115.285 ;
        RECT 88.075 114.995 88.460 115.965 ;
        RECT 88.630 115.915 89.150 116.455 ;
        RECT 89.320 116.085 89.840 116.625 ;
        RECT 90.015 116.135 90.365 116.705 ;
        RECT 90.550 116.635 92.160 116.805 ;
        RECT 92.330 116.700 92.600 117.045 ;
        RECT 91.990 116.465 92.160 116.635 ;
        RECT 90.535 116.015 91.245 116.465 ;
        RECT 91.415 116.135 91.820 116.465 ;
        RECT 91.990 116.135 92.260 116.465 ;
        RECT 88.630 114.825 89.840 115.915 ;
        RECT 90.015 115.675 90.335 115.965 ;
        RECT 90.530 115.845 91.245 116.015 ;
        RECT 91.990 115.965 92.160 116.135 ;
        RECT 92.430 115.965 92.600 116.700 ;
        RECT 92.885 116.745 93.170 117.205 ;
        RECT 93.340 116.915 93.610 117.375 ;
        RECT 92.885 116.575 93.840 116.745 ;
        RECT 91.435 115.795 92.160 115.965 ;
        RECT 91.435 115.675 91.605 115.795 ;
        RECT 90.015 115.505 91.605 115.675 ;
        RECT 90.015 115.045 91.670 115.335 ;
        RECT 91.840 114.825 92.120 115.625 ;
        RECT 92.330 114.995 92.600 115.965 ;
        RECT 92.770 115.845 93.460 116.405 ;
        RECT 93.630 115.675 93.840 116.575 ;
        RECT 92.885 115.455 93.840 115.675 ;
        RECT 94.010 116.405 94.410 117.205 ;
        RECT 94.600 116.745 94.880 117.205 ;
        RECT 95.400 116.915 95.725 117.375 ;
        RECT 94.600 116.575 95.725 116.745 ;
        RECT 95.895 116.635 96.280 117.205 ;
        RECT 96.460 116.875 96.790 117.375 ;
        RECT 96.990 116.805 97.160 117.155 ;
        RECT 97.360 116.975 97.690 117.375 ;
        RECT 97.860 116.805 98.030 117.155 ;
        RECT 98.200 116.975 98.580 117.375 ;
        RECT 95.275 116.465 95.725 116.575 ;
        RECT 94.010 115.845 95.105 116.405 ;
        RECT 95.275 116.135 95.830 116.465 ;
        RECT 92.885 114.995 93.170 115.455 ;
        RECT 93.340 114.825 93.610 115.285 ;
        RECT 94.010 114.995 94.410 115.845 ;
        RECT 95.275 115.675 95.725 116.135 ;
        RECT 96.000 115.965 96.280 116.635 ;
        RECT 96.455 116.135 96.805 116.705 ;
        RECT 96.990 116.635 98.600 116.805 ;
        RECT 98.770 116.700 99.040 117.045 ;
        RECT 98.430 116.465 98.600 116.635 ;
        RECT 96.975 116.015 97.685 116.465 ;
        RECT 97.855 116.135 98.260 116.465 ;
        RECT 98.430 116.135 98.700 116.465 ;
        RECT 94.600 115.455 95.725 115.675 ;
        RECT 94.600 114.995 94.880 115.455 ;
        RECT 95.400 114.825 95.725 115.285 ;
        RECT 95.895 114.995 96.280 115.965 ;
        RECT 96.455 115.675 96.775 115.965 ;
        RECT 96.970 115.845 97.685 116.015 ;
        RECT 98.430 115.965 98.600 116.135 ;
        RECT 98.870 115.965 99.040 116.700 ;
        RECT 99.210 116.650 99.500 117.375 ;
        RECT 99.670 116.915 100.230 117.205 ;
        RECT 100.400 116.915 100.650 117.375 ;
        RECT 97.875 115.795 98.600 115.965 ;
        RECT 97.875 115.675 98.045 115.795 ;
        RECT 96.455 115.505 98.045 115.675 ;
        RECT 96.455 115.045 98.110 115.335 ;
        RECT 98.280 114.825 98.560 115.625 ;
        RECT 98.770 114.995 99.040 115.965 ;
        RECT 99.210 114.825 99.500 115.990 ;
        RECT 99.670 115.545 99.920 116.915 ;
        RECT 101.270 116.745 101.600 117.105 ;
        RECT 100.210 116.555 101.600 116.745 ;
        RECT 101.970 116.915 102.530 117.205 ;
        RECT 102.700 116.915 102.950 117.375 ;
        RECT 100.210 116.465 100.380 116.555 ;
        RECT 100.090 116.135 100.380 116.465 ;
        RECT 100.550 116.135 100.890 116.385 ;
        RECT 101.110 116.135 101.785 116.385 ;
        RECT 100.210 115.885 100.380 116.135 ;
        RECT 100.210 115.715 101.150 115.885 ;
        RECT 101.520 115.775 101.785 116.135 ;
        RECT 99.670 114.995 100.130 115.545 ;
        RECT 100.320 114.825 100.650 115.545 ;
        RECT 100.850 115.165 101.150 115.715 ;
        RECT 101.970 115.545 102.220 116.915 ;
        RECT 103.570 116.745 103.900 117.105 ;
        RECT 102.510 116.555 103.900 116.745 ;
        RECT 104.330 116.555 104.540 117.375 ;
        RECT 104.710 116.575 105.040 117.205 ;
        RECT 102.510 116.465 102.680 116.555 ;
        RECT 102.390 116.135 102.680 116.465 ;
        RECT 102.850 116.135 103.190 116.385 ;
        RECT 103.410 116.135 104.085 116.385 ;
        RECT 102.510 115.885 102.680 116.135 ;
        RECT 102.510 115.715 103.450 115.885 ;
        RECT 103.820 115.775 104.085 116.135 ;
        RECT 104.710 115.975 104.960 116.575 ;
        RECT 105.210 116.555 105.440 117.375 ;
        RECT 105.655 116.830 111.000 117.375 ;
        RECT 105.130 116.135 105.460 116.385 ;
        RECT 101.320 114.825 101.600 115.495 ;
        RECT 101.970 114.995 102.430 115.545 ;
        RECT 102.620 114.825 102.950 115.545 ;
        RECT 103.150 115.165 103.450 115.715 ;
        RECT 103.620 114.825 103.900 115.495 ;
        RECT 104.330 114.825 104.540 115.965 ;
        RECT 104.710 114.995 105.040 115.975 ;
        RECT 105.210 114.825 105.440 115.965 ;
        RECT 107.245 115.260 107.595 116.510 ;
        RECT 109.075 116.000 109.415 116.830 ;
        RECT 111.170 116.625 112.380 117.375 ;
        RECT 111.170 115.915 111.690 116.455 ;
        RECT 111.860 116.085 112.380 116.625 ;
        RECT 105.655 114.825 111.000 115.260 ;
        RECT 111.170 114.825 112.380 115.915 ;
        RECT 18.165 114.655 112.465 114.825 ;
        RECT 18.250 113.565 19.460 114.655 ;
        RECT 20.555 114.220 25.900 114.655 ;
        RECT 18.250 112.855 18.770 113.395 ;
        RECT 18.940 113.025 19.460 113.565 ;
        RECT 22.145 112.970 22.495 114.220 ;
        RECT 26.110 113.515 26.340 114.655 ;
        RECT 26.510 113.505 26.840 114.485 ;
        RECT 27.010 113.515 27.220 114.655 ;
        RECT 27.650 113.985 27.930 114.655 ;
        RECT 28.100 113.765 28.400 114.315 ;
        RECT 28.600 113.935 28.930 114.655 ;
        RECT 29.120 113.935 29.580 114.485 ;
        RECT 29.950 113.985 30.230 114.655 ;
        RECT 18.250 112.105 19.460 112.855 ;
        RECT 23.975 112.650 24.315 113.480 ;
        RECT 26.090 113.095 26.420 113.345 ;
        RECT 20.555 112.105 25.900 112.650 ;
        RECT 26.110 112.105 26.340 112.925 ;
        RECT 26.590 112.905 26.840 113.505 ;
        RECT 27.465 113.345 27.730 113.705 ;
        RECT 28.100 113.595 29.040 113.765 ;
        RECT 28.870 113.345 29.040 113.595 ;
        RECT 27.465 113.095 28.140 113.345 ;
        RECT 28.360 113.095 28.700 113.345 ;
        RECT 28.870 113.015 29.160 113.345 ;
        RECT 28.870 112.925 29.040 113.015 ;
        RECT 26.510 112.275 26.840 112.905 ;
        RECT 27.010 112.105 27.220 112.925 ;
        RECT 27.650 112.735 29.040 112.925 ;
        RECT 27.650 112.375 27.980 112.735 ;
        RECT 29.330 112.565 29.580 113.935 ;
        RECT 30.400 113.765 30.700 114.315 ;
        RECT 30.900 113.935 31.230 114.655 ;
        RECT 31.420 113.935 31.880 114.485 ;
        RECT 29.765 113.345 30.030 113.705 ;
        RECT 30.400 113.595 31.340 113.765 ;
        RECT 31.170 113.345 31.340 113.595 ;
        RECT 29.765 113.095 30.440 113.345 ;
        RECT 30.660 113.095 31.000 113.345 ;
        RECT 31.170 113.015 31.460 113.345 ;
        RECT 31.170 112.925 31.340 113.015 ;
        RECT 28.600 112.105 28.850 112.565 ;
        RECT 29.020 112.275 29.580 112.565 ;
        RECT 29.950 112.735 31.340 112.925 ;
        RECT 29.950 112.375 30.280 112.735 ;
        RECT 31.630 112.565 31.880 113.935 ;
        RECT 30.900 112.105 31.150 112.565 ;
        RECT 31.320 112.275 31.880 112.565 ;
        RECT 32.050 113.515 32.320 114.485 ;
        RECT 32.530 113.855 32.810 114.655 ;
        RECT 32.980 114.145 34.635 114.435 ;
        RECT 33.045 113.805 34.635 113.975 ;
        RECT 33.045 113.685 33.215 113.805 ;
        RECT 32.490 113.515 33.215 113.685 ;
        RECT 32.050 112.780 32.220 113.515 ;
        RECT 32.490 113.345 32.660 113.515 ;
        RECT 33.405 113.465 34.120 113.635 ;
        RECT 34.315 113.515 34.635 113.805 ;
        RECT 34.810 113.490 35.100 114.655 ;
        RECT 35.270 113.685 35.540 114.455 ;
        RECT 35.710 113.875 36.040 114.655 ;
        RECT 36.245 114.050 36.430 114.455 ;
        RECT 36.600 114.230 36.935 114.655 ;
        RECT 36.245 113.875 36.910 114.050 ;
        RECT 35.270 113.515 36.400 113.685 ;
        RECT 32.390 113.015 32.660 113.345 ;
        RECT 32.830 113.015 33.235 113.345 ;
        RECT 33.405 113.015 34.115 113.465 ;
        RECT 32.490 112.845 32.660 113.015 ;
        RECT 32.050 112.435 32.320 112.780 ;
        RECT 32.490 112.675 34.100 112.845 ;
        RECT 34.285 112.775 34.635 113.345 ;
        RECT 32.510 112.105 32.890 112.505 ;
        RECT 33.060 112.325 33.230 112.675 ;
        RECT 33.400 112.105 33.730 112.505 ;
        RECT 33.930 112.325 34.100 112.675 ;
        RECT 34.300 112.105 34.630 112.605 ;
        RECT 34.810 112.105 35.100 112.830 ;
        RECT 35.270 112.605 35.440 113.515 ;
        RECT 35.610 112.765 35.970 113.345 ;
        RECT 36.150 113.015 36.400 113.515 ;
        RECT 36.570 112.845 36.910 113.875 ;
        RECT 36.225 112.675 36.910 112.845 ;
        RECT 37.110 113.515 37.450 114.485 ;
        RECT 37.620 113.515 37.790 114.655 ;
        RECT 38.060 113.855 38.310 114.655 ;
        RECT 38.955 113.685 39.285 114.485 ;
        RECT 39.585 113.855 39.915 114.655 ;
        RECT 40.085 113.685 40.415 114.485 ;
        RECT 37.980 113.515 40.415 113.685 ;
        RECT 40.790 113.895 41.305 114.305 ;
        RECT 41.540 113.895 41.710 114.655 ;
        RECT 41.880 114.315 43.910 114.485 ;
        RECT 37.110 112.905 37.285 113.515 ;
        RECT 37.980 113.265 38.150 113.515 ;
        RECT 37.455 113.095 38.150 113.265 ;
        RECT 38.325 113.095 38.745 113.295 ;
        RECT 38.915 113.095 39.245 113.295 ;
        RECT 39.415 113.095 39.745 113.295 ;
        RECT 35.270 112.275 35.530 112.605 ;
        RECT 35.740 112.105 36.015 112.585 ;
        RECT 36.225 112.275 36.430 112.675 ;
        RECT 36.600 112.105 36.935 112.505 ;
        RECT 37.110 112.275 37.450 112.905 ;
        RECT 37.620 112.105 37.870 112.905 ;
        RECT 38.060 112.755 39.285 112.925 ;
        RECT 38.060 112.275 38.390 112.755 ;
        RECT 38.560 112.105 38.785 112.565 ;
        RECT 38.955 112.275 39.285 112.755 ;
        RECT 39.915 112.885 40.085 113.515 ;
        RECT 40.270 113.095 40.620 113.345 ;
        RECT 40.790 113.085 41.130 113.895 ;
        RECT 41.880 113.650 42.050 114.315 ;
        RECT 42.445 113.975 43.570 114.145 ;
        RECT 41.300 113.460 42.050 113.650 ;
        RECT 42.220 113.635 43.230 113.805 ;
        RECT 40.790 112.915 42.020 113.085 ;
        RECT 39.915 112.275 40.415 112.885 ;
        RECT 41.065 112.310 41.310 112.915 ;
        RECT 41.530 112.105 42.040 112.640 ;
        RECT 42.220 112.275 42.410 113.635 ;
        RECT 42.580 112.615 42.855 113.435 ;
        RECT 43.060 112.835 43.230 113.635 ;
        RECT 43.400 112.845 43.570 113.975 ;
        RECT 43.740 113.345 43.910 114.315 ;
        RECT 44.080 113.515 44.250 114.655 ;
        RECT 44.420 113.515 44.755 114.485 ;
        RECT 43.740 113.015 43.935 113.345 ;
        RECT 44.160 113.015 44.415 113.345 ;
        RECT 44.160 112.845 44.330 113.015 ;
        RECT 44.585 112.845 44.755 113.515 ;
        RECT 43.400 112.675 44.330 112.845 ;
        RECT 43.400 112.640 43.575 112.675 ;
        RECT 42.580 112.445 42.860 112.615 ;
        RECT 42.580 112.275 42.855 112.445 ;
        RECT 43.045 112.275 43.575 112.640 ;
        RECT 44.000 112.105 44.330 112.505 ;
        RECT 44.500 112.275 44.755 112.845 ;
        RECT 45.390 113.935 45.850 114.485 ;
        RECT 46.040 113.935 46.370 114.655 ;
        RECT 45.390 112.565 45.640 113.935 ;
        RECT 46.570 113.765 46.870 114.315 ;
        RECT 47.040 113.985 47.320 114.655 ;
        RECT 45.930 113.595 46.870 113.765 ;
        RECT 45.930 113.345 46.100 113.595 ;
        RECT 47.240 113.345 47.505 113.705 ;
        RECT 45.810 113.015 46.100 113.345 ;
        RECT 46.270 113.095 46.610 113.345 ;
        RECT 46.830 113.095 47.505 113.345 ;
        RECT 47.690 113.565 49.360 114.655 ;
        RECT 49.535 114.220 54.880 114.655 ;
        RECT 47.690 113.045 48.440 113.565 ;
        RECT 45.930 112.925 46.100 113.015 ;
        RECT 45.930 112.735 47.320 112.925 ;
        RECT 48.610 112.875 49.360 113.395 ;
        RECT 51.125 112.970 51.475 114.220 ;
        RECT 55.090 113.515 55.320 114.655 ;
        RECT 55.490 113.505 55.820 114.485 ;
        RECT 55.990 113.515 56.200 114.655 ;
        RECT 56.430 113.895 56.945 114.305 ;
        RECT 57.180 113.895 57.350 114.655 ;
        RECT 57.520 114.315 59.550 114.485 ;
        RECT 45.390 112.275 45.950 112.565 ;
        RECT 46.120 112.105 46.370 112.565 ;
        RECT 46.990 112.375 47.320 112.735 ;
        RECT 47.690 112.105 49.360 112.875 ;
        RECT 52.955 112.650 53.295 113.480 ;
        RECT 55.070 113.095 55.400 113.345 ;
        RECT 49.535 112.105 54.880 112.650 ;
        RECT 55.090 112.105 55.320 112.925 ;
        RECT 55.570 112.905 55.820 113.505 ;
        RECT 56.430 113.085 56.770 113.895 ;
        RECT 57.520 113.650 57.690 114.315 ;
        RECT 58.085 113.975 59.210 114.145 ;
        RECT 56.940 113.460 57.690 113.650 ;
        RECT 57.860 113.635 58.870 113.805 ;
        RECT 55.490 112.275 55.820 112.905 ;
        RECT 55.990 112.105 56.200 112.925 ;
        RECT 56.430 112.915 57.660 113.085 ;
        RECT 56.705 112.310 56.950 112.915 ;
        RECT 57.170 112.105 57.680 112.640 ;
        RECT 57.860 112.275 58.050 113.635 ;
        RECT 58.220 112.615 58.495 113.435 ;
        RECT 58.700 112.835 58.870 113.635 ;
        RECT 59.040 112.845 59.210 113.975 ;
        RECT 59.380 113.345 59.550 114.315 ;
        RECT 59.720 113.515 59.890 114.655 ;
        RECT 60.060 113.515 60.395 114.485 ;
        RECT 59.380 113.015 59.575 113.345 ;
        RECT 59.800 113.015 60.055 113.345 ;
        RECT 59.800 112.845 59.970 113.015 ;
        RECT 60.225 112.845 60.395 113.515 ;
        RECT 60.570 113.490 60.860 114.655 ;
        RECT 61.490 113.685 61.760 114.455 ;
        RECT 61.930 113.875 62.260 114.655 ;
        RECT 62.465 114.050 62.650 114.455 ;
        RECT 62.820 114.230 63.155 114.655 ;
        RECT 62.465 113.875 63.130 114.050 ;
        RECT 61.490 113.515 62.620 113.685 ;
        RECT 59.040 112.675 59.970 112.845 ;
        RECT 59.040 112.640 59.215 112.675 ;
        RECT 58.220 112.445 58.500 112.615 ;
        RECT 58.220 112.275 58.495 112.445 ;
        RECT 58.685 112.275 59.215 112.640 ;
        RECT 59.640 112.105 59.970 112.505 ;
        RECT 60.140 112.275 60.395 112.845 ;
        RECT 60.570 112.105 60.860 112.830 ;
        RECT 61.490 112.605 61.660 113.515 ;
        RECT 61.830 112.765 62.190 113.345 ;
        RECT 62.370 113.015 62.620 113.515 ;
        RECT 62.790 112.845 63.130 113.875 ;
        RECT 63.790 113.565 67.300 114.655 ;
        RECT 67.470 113.935 67.930 114.485 ;
        RECT 68.120 113.935 68.450 114.655 ;
        RECT 63.790 113.045 65.480 113.565 ;
        RECT 65.650 112.875 67.300 113.395 ;
        RECT 62.445 112.675 63.130 112.845 ;
        RECT 61.490 112.275 61.750 112.605 ;
        RECT 61.960 112.105 62.235 112.585 ;
        RECT 62.445 112.275 62.650 112.675 ;
        RECT 62.820 112.105 63.155 112.505 ;
        RECT 63.790 112.105 67.300 112.875 ;
        RECT 67.470 112.565 67.720 113.935 ;
        RECT 68.650 113.765 68.950 114.315 ;
        RECT 69.120 113.985 69.400 114.655 ;
        RECT 70.430 113.985 70.710 114.655 ;
        RECT 68.010 113.595 68.950 113.765 ;
        RECT 70.880 113.765 71.180 114.315 ;
        RECT 71.380 113.935 71.710 114.655 ;
        RECT 71.900 113.935 72.360 114.485 ;
        RECT 68.010 113.345 68.180 113.595 ;
        RECT 69.320 113.345 69.585 113.705 ;
        RECT 67.890 113.015 68.180 113.345 ;
        RECT 68.350 113.095 68.690 113.345 ;
        RECT 68.910 113.095 69.585 113.345 ;
        RECT 70.245 113.345 70.510 113.705 ;
        RECT 70.880 113.595 71.820 113.765 ;
        RECT 71.650 113.345 71.820 113.595 ;
        RECT 70.245 113.095 70.920 113.345 ;
        RECT 71.140 113.095 71.480 113.345 ;
        RECT 68.010 112.925 68.180 113.015 ;
        RECT 71.650 113.015 71.940 113.345 ;
        RECT 71.650 112.925 71.820 113.015 ;
        RECT 68.010 112.735 69.400 112.925 ;
        RECT 67.470 112.275 68.030 112.565 ;
        RECT 68.200 112.105 68.450 112.565 ;
        RECT 69.070 112.375 69.400 112.735 ;
        RECT 70.430 112.735 71.820 112.925 ;
        RECT 70.430 112.375 70.760 112.735 ;
        RECT 72.110 112.565 72.360 113.935 ;
        RECT 72.645 114.025 72.930 114.485 ;
        RECT 73.100 114.195 73.370 114.655 ;
        RECT 72.645 113.805 73.600 114.025 ;
        RECT 72.530 113.075 73.220 113.635 ;
        RECT 73.390 112.905 73.600 113.805 ;
        RECT 71.380 112.105 71.630 112.565 ;
        RECT 71.800 112.275 72.360 112.565 ;
        RECT 72.645 112.735 73.600 112.905 ;
        RECT 73.770 113.635 74.170 114.485 ;
        RECT 74.360 114.025 74.640 114.485 ;
        RECT 75.160 114.195 75.485 114.655 ;
        RECT 74.360 113.805 75.485 114.025 ;
        RECT 73.770 113.075 74.865 113.635 ;
        RECT 75.035 113.345 75.485 113.805 ;
        RECT 75.655 113.515 76.040 114.485 ;
        RECT 72.645 112.275 72.930 112.735 ;
        RECT 73.100 112.105 73.370 112.565 ;
        RECT 73.770 112.275 74.170 113.075 ;
        RECT 75.035 113.015 75.590 113.345 ;
        RECT 75.035 112.905 75.485 113.015 ;
        RECT 74.360 112.735 75.485 112.905 ;
        RECT 75.760 112.845 76.040 113.515 ;
        RECT 74.360 112.275 74.640 112.735 ;
        RECT 75.160 112.105 75.485 112.565 ;
        RECT 75.655 112.275 76.040 112.845 ;
        RECT 76.210 113.515 76.595 114.485 ;
        RECT 76.765 114.195 77.090 114.655 ;
        RECT 77.610 114.025 77.890 114.485 ;
        RECT 76.765 113.805 77.890 114.025 ;
        RECT 76.210 112.845 76.490 113.515 ;
        RECT 76.765 113.345 77.215 113.805 ;
        RECT 78.080 113.635 78.480 114.485 ;
        RECT 78.880 114.195 79.150 114.655 ;
        RECT 79.320 114.025 79.605 114.485 ;
        RECT 79.895 114.145 81.550 114.435 ;
        RECT 76.660 113.015 77.215 113.345 ;
        RECT 77.385 113.075 78.480 113.635 ;
        RECT 76.765 112.905 77.215 113.015 ;
        RECT 76.210 112.275 76.595 112.845 ;
        RECT 76.765 112.735 77.890 112.905 ;
        RECT 76.765 112.105 77.090 112.565 ;
        RECT 77.610 112.275 77.890 112.735 ;
        RECT 78.080 112.275 78.480 113.075 ;
        RECT 78.650 113.805 79.605 114.025 ;
        RECT 79.895 113.805 81.485 113.975 ;
        RECT 81.720 113.855 82.000 114.655 ;
        RECT 78.650 112.905 78.860 113.805 ;
        RECT 79.030 113.075 79.720 113.635 ;
        RECT 79.895 113.515 80.215 113.805 ;
        RECT 81.315 113.685 81.485 113.805 ;
        RECT 78.650 112.735 79.605 112.905 ;
        RECT 79.895 112.775 80.245 113.345 ;
        RECT 80.415 113.015 81.125 113.635 ;
        RECT 81.315 113.515 82.040 113.685 ;
        RECT 82.210 113.515 82.480 114.485 ;
        RECT 81.870 113.345 82.040 113.515 ;
        RECT 81.295 113.015 81.700 113.345 ;
        RECT 81.870 113.015 82.140 113.345 ;
        RECT 81.870 112.845 82.040 113.015 ;
        RECT 78.880 112.105 79.150 112.565 ;
        RECT 79.320 112.275 79.605 112.735 ;
        RECT 80.430 112.675 82.040 112.845 ;
        RECT 82.310 112.780 82.480 113.515 ;
        RECT 79.900 112.105 80.230 112.605 ;
        RECT 80.430 112.325 80.600 112.675 ;
        RECT 80.800 112.105 81.130 112.505 ;
        RECT 81.300 112.325 81.470 112.675 ;
        RECT 81.640 112.105 82.020 112.505 ;
        RECT 82.210 112.435 82.480 112.780 ;
        RECT 83.570 113.515 83.840 114.485 ;
        RECT 84.050 113.855 84.330 114.655 ;
        RECT 84.500 114.145 86.155 114.435 ;
        RECT 84.565 113.805 86.155 113.975 ;
        RECT 84.565 113.685 84.735 113.805 ;
        RECT 84.010 113.515 84.735 113.685 ;
        RECT 83.570 112.780 83.740 113.515 ;
        RECT 84.010 113.345 84.180 113.515 ;
        RECT 84.925 113.465 85.640 113.635 ;
        RECT 85.835 113.515 86.155 113.805 ;
        RECT 86.330 113.490 86.620 114.655 ;
        RECT 86.850 113.515 87.060 114.655 ;
        RECT 87.230 113.505 87.560 114.485 ;
        RECT 87.730 113.515 87.960 114.655 ;
        RECT 88.170 113.895 88.685 114.305 ;
        RECT 88.920 113.895 89.090 114.655 ;
        RECT 89.260 114.315 91.290 114.485 ;
        RECT 83.910 113.015 84.180 113.345 ;
        RECT 84.350 113.015 84.755 113.345 ;
        RECT 84.925 113.015 85.635 113.465 ;
        RECT 84.010 112.845 84.180 113.015 ;
        RECT 83.570 112.435 83.840 112.780 ;
        RECT 84.010 112.675 85.620 112.845 ;
        RECT 85.805 112.775 86.155 113.345 ;
        RECT 84.030 112.105 84.410 112.505 ;
        RECT 84.580 112.325 84.750 112.675 ;
        RECT 84.920 112.105 85.250 112.505 ;
        RECT 85.450 112.325 85.620 112.675 ;
        RECT 85.820 112.105 86.150 112.605 ;
        RECT 86.330 112.105 86.620 112.830 ;
        RECT 86.850 112.105 87.060 112.925 ;
        RECT 87.230 112.905 87.480 113.505 ;
        RECT 87.650 113.095 87.980 113.345 ;
        RECT 88.170 113.085 88.510 113.895 ;
        RECT 89.260 113.650 89.430 114.315 ;
        RECT 89.825 113.975 90.950 114.145 ;
        RECT 88.680 113.460 89.430 113.650 ;
        RECT 89.600 113.635 90.610 113.805 ;
        RECT 87.230 112.275 87.560 112.905 ;
        RECT 87.730 112.105 87.960 112.925 ;
        RECT 88.170 112.915 89.400 113.085 ;
        RECT 88.445 112.310 88.690 112.915 ;
        RECT 88.910 112.105 89.420 112.640 ;
        RECT 89.600 112.275 89.790 113.635 ;
        RECT 89.960 113.295 90.235 113.435 ;
        RECT 89.960 113.125 90.240 113.295 ;
        RECT 89.960 112.275 90.235 113.125 ;
        RECT 90.440 112.835 90.610 113.635 ;
        RECT 90.780 112.845 90.950 113.975 ;
        RECT 91.120 113.345 91.290 114.315 ;
        RECT 91.460 113.515 91.630 114.655 ;
        RECT 91.800 113.515 92.135 114.485 ;
        RECT 91.120 113.015 91.315 113.345 ;
        RECT 91.540 113.015 91.795 113.345 ;
        RECT 91.540 112.845 91.710 113.015 ;
        RECT 91.965 112.845 92.135 113.515 ;
        RECT 92.685 113.675 92.940 114.345 ;
        RECT 93.120 113.855 93.405 114.655 ;
        RECT 93.585 113.935 93.915 114.445 ;
        RECT 92.685 112.955 92.865 113.675 ;
        RECT 93.585 113.345 93.835 113.935 ;
        RECT 94.185 113.785 94.355 114.395 ;
        RECT 94.525 113.965 94.855 114.655 ;
        RECT 95.085 114.105 95.325 114.395 ;
        RECT 95.525 114.275 95.945 114.655 ;
        RECT 96.125 114.185 96.755 114.435 ;
        RECT 97.225 114.275 97.555 114.655 ;
        RECT 96.125 114.105 96.295 114.185 ;
        RECT 97.725 114.105 97.895 114.395 ;
        RECT 98.075 114.275 98.455 114.655 ;
        RECT 98.695 114.270 99.525 114.440 ;
        RECT 95.085 113.935 96.295 114.105 ;
        RECT 93.035 113.015 93.835 113.345 ;
        RECT 90.780 112.675 91.710 112.845 ;
        RECT 90.780 112.640 90.955 112.675 ;
        RECT 90.425 112.275 90.955 112.640 ;
        RECT 91.380 112.105 91.710 112.505 ;
        RECT 91.880 112.275 92.135 112.845 ;
        RECT 92.600 112.815 92.865 112.955 ;
        RECT 92.600 112.785 92.940 112.815 ;
        RECT 92.685 112.285 92.940 112.785 ;
        RECT 93.120 112.105 93.405 112.565 ;
        RECT 93.585 112.365 93.835 113.015 ;
        RECT 94.035 113.765 94.355 113.785 ;
        RECT 94.035 113.595 95.955 113.765 ;
        RECT 94.035 112.700 94.225 113.595 ;
        RECT 96.125 113.425 96.295 113.935 ;
        RECT 96.465 113.675 96.985 113.985 ;
        RECT 94.395 113.255 96.295 113.425 ;
        RECT 94.395 113.195 94.725 113.255 ;
        RECT 94.875 113.025 95.205 113.085 ;
        RECT 94.545 112.755 95.205 113.025 ;
        RECT 94.035 112.370 94.355 112.700 ;
        RECT 94.535 112.105 95.195 112.585 ;
        RECT 95.395 112.495 95.565 113.255 ;
        RECT 96.465 113.085 96.645 113.495 ;
        RECT 95.735 112.915 96.065 113.035 ;
        RECT 96.815 112.915 96.985 113.675 ;
        RECT 95.735 112.745 96.985 112.915 ;
        RECT 97.155 113.855 98.525 114.105 ;
        RECT 97.155 113.085 97.345 113.855 ;
        RECT 98.275 113.595 98.525 113.855 ;
        RECT 97.515 113.425 97.765 113.585 ;
        RECT 98.695 113.425 98.865 114.270 ;
        RECT 99.760 113.985 99.930 114.485 ;
        RECT 100.100 114.155 100.430 114.655 ;
        RECT 99.035 113.595 99.535 113.975 ;
        RECT 99.760 113.815 100.455 113.985 ;
        RECT 97.515 113.255 98.865 113.425 ;
        RECT 98.445 113.215 98.865 113.255 ;
        RECT 97.155 112.745 97.575 113.085 ;
        RECT 97.865 112.755 98.275 113.085 ;
        RECT 95.395 112.325 96.245 112.495 ;
        RECT 96.805 112.105 97.125 112.565 ;
        RECT 97.325 112.315 97.575 112.745 ;
        RECT 97.865 112.105 98.275 112.545 ;
        RECT 98.445 112.485 98.615 113.215 ;
        RECT 98.785 112.665 99.135 113.035 ;
        RECT 99.315 112.725 99.535 113.595 ;
        RECT 99.705 113.025 100.115 113.645 ;
        RECT 100.285 112.845 100.455 113.815 ;
        RECT 99.760 112.655 100.455 112.845 ;
        RECT 98.445 112.285 99.460 112.485 ;
        RECT 99.760 112.325 99.930 112.655 ;
        RECT 100.100 112.105 100.430 112.485 ;
        RECT 100.645 112.365 100.870 114.485 ;
        RECT 101.040 114.155 101.370 114.655 ;
        RECT 101.540 113.985 101.710 114.485 ;
        RECT 101.045 113.815 101.710 113.985 ;
        RECT 101.045 112.825 101.275 113.815 ;
        RECT 101.445 112.995 101.795 113.645 ;
        RECT 101.970 113.565 105.480 114.655 ;
        RECT 105.655 114.220 111.000 114.655 ;
        RECT 101.970 113.045 103.660 113.565 ;
        RECT 103.830 112.875 105.480 113.395 ;
        RECT 107.245 112.970 107.595 114.220 ;
        RECT 111.170 113.565 112.380 114.655 ;
        RECT 101.045 112.655 101.710 112.825 ;
        RECT 101.040 112.105 101.370 112.485 ;
        RECT 101.540 112.365 101.710 112.655 ;
        RECT 101.970 112.105 105.480 112.875 ;
        RECT 109.075 112.650 109.415 113.480 ;
        RECT 111.170 113.025 111.690 113.565 ;
        RECT 111.860 112.855 112.380 113.395 ;
        RECT 105.655 112.105 111.000 112.650 ;
        RECT 111.170 112.105 112.380 112.855 ;
        RECT 18.165 111.935 112.465 112.105 ;
        RECT 18.250 111.185 19.460 111.935 ;
        RECT 18.250 110.645 18.770 111.185 ;
        RECT 20.090 111.165 21.760 111.935 ;
        RECT 21.930 111.210 22.220 111.935 ;
        RECT 22.390 111.165 24.980 111.935 ;
        RECT 25.155 111.390 30.500 111.935 ;
        RECT 18.940 110.475 19.460 111.015 ;
        RECT 18.250 109.385 19.460 110.475 ;
        RECT 20.090 110.475 20.840 110.995 ;
        RECT 21.010 110.645 21.760 111.165 ;
        RECT 20.090 109.385 21.760 110.475 ;
        RECT 21.930 109.385 22.220 110.550 ;
        RECT 22.390 110.475 23.600 110.995 ;
        RECT 23.770 110.645 24.980 111.165 ;
        RECT 22.390 109.385 24.980 110.475 ;
        RECT 26.745 109.820 27.095 111.070 ;
        RECT 28.575 110.560 28.915 111.390 ;
        RECT 30.710 111.115 30.940 111.935 ;
        RECT 31.110 111.135 31.440 111.765 ;
        RECT 30.690 110.695 31.020 110.945 ;
        RECT 31.190 110.535 31.440 111.135 ;
        RECT 31.610 111.115 31.820 111.935 ;
        RECT 32.050 111.260 32.320 111.605 ;
        RECT 32.510 111.535 32.890 111.935 ;
        RECT 33.060 111.365 33.230 111.715 ;
        RECT 33.400 111.535 33.730 111.935 ;
        RECT 33.930 111.365 34.100 111.715 ;
        RECT 34.300 111.435 34.630 111.935 ;
        RECT 25.155 109.385 30.500 109.820 ;
        RECT 30.710 109.385 30.940 110.525 ;
        RECT 31.110 109.555 31.440 110.535 ;
        RECT 32.050 110.525 32.220 111.260 ;
        RECT 32.490 111.195 34.100 111.365 ;
        RECT 32.490 111.025 32.660 111.195 ;
        RECT 32.390 110.695 32.660 111.025 ;
        RECT 32.830 110.695 33.235 111.025 ;
        RECT 32.490 110.525 32.660 110.695 ;
        RECT 31.610 109.385 31.820 110.525 ;
        RECT 32.050 109.555 32.320 110.525 ;
        RECT 32.490 110.355 33.215 110.525 ;
        RECT 33.405 110.405 34.115 111.025 ;
        RECT 34.285 110.695 34.635 111.265 ;
        RECT 34.810 111.260 35.080 111.605 ;
        RECT 35.270 111.535 35.650 111.935 ;
        RECT 35.820 111.365 35.990 111.715 ;
        RECT 36.160 111.535 36.490 111.935 ;
        RECT 36.690 111.365 36.860 111.715 ;
        RECT 37.060 111.435 37.390 111.935 ;
        RECT 34.810 110.525 34.980 111.260 ;
        RECT 35.250 111.195 36.860 111.365 ;
        RECT 35.250 111.025 35.420 111.195 ;
        RECT 35.150 110.695 35.420 111.025 ;
        RECT 35.590 110.695 35.995 111.025 ;
        RECT 35.250 110.525 35.420 110.695 ;
        RECT 33.045 110.235 33.215 110.355 ;
        RECT 34.315 110.235 34.635 110.525 ;
        RECT 32.530 109.385 32.810 110.185 ;
        RECT 33.045 110.065 34.635 110.235 ;
        RECT 32.980 109.605 34.635 109.895 ;
        RECT 34.810 109.555 35.080 110.525 ;
        RECT 35.250 110.355 35.975 110.525 ;
        RECT 36.165 110.405 36.875 111.025 ;
        RECT 37.045 110.695 37.395 111.265 ;
        RECT 37.945 111.225 38.200 111.755 ;
        RECT 38.380 111.475 38.665 111.935 ;
        RECT 37.945 110.575 38.125 111.225 ;
        RECT 38.845 111.025 39.095 111.675 ;
        RECT 38.295 110.695 39.095 111.025 ;
        RECT 35.805 110.235 35.975 110.355 ;
        RECT 37.075 110.235 37.395 110.525 ;
        RECT 37.860 110.405 38.125 110.575 ;
        RECT 35.290 109.385 35.570 110.185 ;
        RECT 35.805 110.065 37.395 110.235 ;
        RECT 37.945 110.365 38.125 110.405 ;
        RECT 35.740 109.605 37.395 109.895 ;
        RECT 37.945 109.695 38.200 110.365 ;
        RECT 38.380 109.385 38.665 110.185 ;
        RECT 38.845 110.105 39.095 110.695 ;
        RECT 39.295 111.340 39.615 111.670 ;
        RECT 39.795 111.455 40.455 111.935 ;
        RECT 40.655 111.545 41.505 111.715 ;
        RECT 39.295 110.445 39.485 111.340 ;
        RECT 39.805 111.015 40.465 111.285 ;
        RECT 40.135 110.955 40.465 111.015 ;
        RECT 39.655 110.785 39.985 110.845 ;
        RECT 40.655 110.785 40.825 111.545 ;
        RECT 42.065 111.475 42.385 111.935 ;
        RECT 42.585 111.295 42.835 111.725 ;
        RECT 43.125 111.495 43.535 111.935 ;
        RECT 43.705 111.555 44.720 111.755 ;
        RECT 40.995 111.125 42.245 111.295 ;
        RECT 40.995 111.005 41.325 111.125 ;
        RECT 39.655 110.615 41.555 110.785 ;
        RECT 39.295 110.275 41.215 110.445 ;
        RECT 39.295 110.255 39.615 110.275 ;
        RECT 38.845 109.595 39.175 110.105 ;
        RECT 39.445 109.645 39.615 110.255 ;
        RECT 41.385 110.105 41.555 110.615 ;
        RECT 41.725 110.545 41.905 110.955 ;
        RECT 42.075 110.365 42.245 111.125 ;
        RECT 39.785 109.385 40.115 110.075 ;
        RECT 40.345 109.935 41.555 110.105 ;
        RECT 41.725 110.055 42.245 110.365 ;
        RECT 42.415 110.955 42.835 111.295 ;
        RECT 43.125 110.955 43.535 111.285 ;
        RECT 42.415 110.185 42.605 110.955 ;
        RECT 43.705 110.825 43.875 111.555 ;
        RECT 45.020 111.385 45.190 111.715 ;
        RECT 45.360 111.555 45.690 111.935 ;
        RECT 44.045 111.005 44.395 111.375 ;
        RECT 43.705 110.785 44.125 110.825 ;
        RECT 42.775 110.615 44.125 110.785 ;
        RECT 42.775 110.455 43.025 110.615 ;
        RECT 43.535 110.185 43.785 110.445 ;
        RECT 42.415 109.935 43.785 110.185 ;
        RECT 40.345 109.645 40.585 109.935 ;
        RECT 41.385 109.855 41.555 109.935 ;
        RECT 40.785 109.385 41.205 109.765 ;
        RECT 41.385 109.605 42.015 109.855 ;
        RECT 42.485 109.385 42.815 109.765 ;
        RECT 42.985 109.645 43.155 109.935 ;
        RECT 43.955 109.770 44.125 110.615 ;
        RECT 44.575 110.445 44.795 111.315 ;
        RECT 45.020 111.195 45.715 111.385 ;
        RECT 44.295 110.065 44.795 110.445 ;
        RECT 44.965 110.395 45.375 111.015 ;
        RECT 45.545 110.225 45.715 111.195 ;
        RECT 45.020 110.055 45.715 110.225 ;
        RECT 43.335 109.385 43.715 109.765 ;
        RECT 43.955 109.600 44.785 109.770 ;
        RECT 45.020 109.555 45.190 110.055 ;
        RECT 45.360 109.385 45.690 109.885 ;
        RECT 45.905 109.555 46.130 111.675 ;
        RECT 46.300 111.555 46.630 111.935 ;
        RECT 46.800 111.385 46.970 111.675 ;
        RECT 46.305 111.215 46.970 111.385 ;
        RECT 46.305 110.225 46.535 111.215 ;
        RECT 47.690 111.210 47.980 111.935 ;
        RECT 48.210 111.115 48.420 111.935 ;
        RECT 48.590 111.135 48.920 111.765 ;
        RECT 46.705 110.395 47.055 111.045 ;
        RECT 46.305 110.055 46.970 110.225 ;
        RECT 46.300 109.385 46.630 109.885 ;
        RECT 46.800 109.555 46.970 110.055 ;
        RECT 47.690 109.385 47.980 110.550 ;
        RECT 48.590 110.535 48.840 111.135 ;
        RECT 49.090 111.115 49.320 111.935 ;
        RECT 49.990 111.165 53.500 111.935 ;
        RECT 54.045 111.595 54.300 111.755 ;
        RECT 53.960 111.425 54.300 111.595 ;
        RECT 54.480 111.475 54.765 111.935 ;
        RECT 49.010 110.695 49.340 110.945 ;
        RECT 48.210 109.385 48.420 110.525 ;
        RECT 48.590 109.555 48.920 110.535 ;
        RECT 49.090 109.385 49.320 110.525 ;
        RECT 49.990 110.475 51.680 110.995 ;
        RECT 51.850 110.645 53.500 111.165 ;
        RECT 54.045 111.225 54.300 111.425 ;
        RECT 49.990 109.385 53.500 110.475 ;
        RECT 54.045 110.365 54.225 111.225 ;
        RECT 54.945 111.025 55.195 111.675 ;
        RECT 54.395 110.695 55.195 111.025 ;
        RECT 54.045 109.695 54.300 110.365 ;
        RECT 54.480 109.385 54.765 110.185 ;
        RECT 54.945 110.105 55.195 110.695 ;
        RECT 55.395 111.340 55.715 111.670 ;
        RECT 55.895 111.455 56.555 111.935 ;
        RECT 56.755 111.545 57.605 111.715 ;
        RECT 55.395 110.445 55.585 111.340 ;
        RECT 55.905 111.015 56.565 111.285 ;
        RECT 56.235 110.955 56.565 111.015 ;
        RECT 55.755 110.785 56.085 110.845 ;
        RECT 56.755 110.785 56.925 111.545 ;
        RECT 58.165 111.475 58.485 111.935 ;
        RECT 58.685 111.295 58.935 111.725 ;
        RECT 59.225 111.495 59.635 111.935 ;
        RECT 59.805 111.555 60.820 111.755 ;
        RECT 57.095 111.125 58.345 111.295 ;
        RECT 57.095 111.005 57.425 111.125 ;
        RECT 55.755 110.615 57.655 110.785 ;
        RECT 55.395 110.275 57.315 110.445 ;
        RECT 55.395 110.255 55.715 110.275 ;
        RECT 54.945 109.595 55.275 110.105 ;
        RECT 55.545 109.645 55.715 110.255 ;
        RECT 57.485 110.105 57.655 110.615 ;
        RECT 57.825 110.545 58.005 110.955 ;
        RECT 58.175 110.365 58.345 111.125 ;
        RECT 55.885 109.385 56.215 110.075 ;
        RECT 56.445 109.935 57.655 110.105 ;
        RECT 57.825 110.055 58.345 110.365 ;
        RECT 58.515 110.955 58.935 111.295 ;
        RECT 59.225 110.955 59.635 111.285 ;
        RECT 58.515 110.185 58.705 110.955 ;
        RECT 59.805 110.825 59.975 111.555 ;
        RECT 61.120 111.385 61.290 111.715 ;
        RECT 61.460 111.555 61.790 111.935 ;
        RECT 60.145 111.005 60.495 111.375 ;
        RECT 59.805 110.785 60.225 110.825 ;
        RECT 58.875 110.615 60.225 110.785 ;
        RECT 58.875 110.455 59.125 110.615 ;
        RECT 59.635 110.185 59.885 110.445 ;
        RECT 58.515 109.935 59.885 110.185 ;
        RECT 56.445 109.645 56.685 109.935 ;
        RECT 57.485 109.855 57.655 109.935 ;
        RECT 56.885 109.385 57.305 109.765 ;
        RECT 57.485 109.605 58.115 109.855 ;
        RECT 58.585 109.385 58.915 109.765 ;
        RECT 59.085 109.645 59.255 109.935 ;
        RECT 60.055 109.770 60.225 110.615 ;
        RECT 60.675 110.445 60.895 111.315 ;
        RECT 61.120 111.195 61.815 111.385 ;
        RECT 60.395 110.065 60.895 110.445 ;
        RECT 61.065 110.395 61.475 111.015 ;
        RECT 61.645 110.225 61.815 111.195 ;
        RECT 61.120 110.055 61.815 110.225 ;
        RECT 59.435 109.385 59.815 109.765 ;
        RECT 60.055 109.600 60.885 109.770 ;
        RECT 61.120 109.555 61.290 110.055 ;
        RECT 61.460 109.385 61.790 109.885 ;
        RECT 62.005 109.555 62.230 111.675 ;
        RECT 62.400 111.555 62.730 111.935 ;
        RECT 62.900 111.385 63.070 111.675 ;
        RECT 62.405 111.215 63.070 111.385 ;
        RECT 62.405 110.225 62.635 111.215 ;
        RECT 63.370 111.115 63.600 111.935 ;
        RECT 63.770 111.135 64.100 111.765 ;
        RECT 62.805 110.395 63.155 111.045 ;
        RECT 63.350 110.695 63.680 110.945 ;
        RECT 63.850 110.535 64.100 111.135 ;
        RECT 64.270 111.115 64.480 111.935 ;
        RECT 65.170 111.165 67.760 111.935 ;
        RECT 62.405 110.055 63.070 110.225 ;
        RECT 62.400 109.385 62.730 109.885 ;
        RECT 62.900 109.555 63.070 110.055 ;
        RECT 63.370 109.385 63.600 110.525 ;
        RECT 63.770 109.555 64.100 110.535 ;
        RECT 64.270 109.385 64.480 110.525 ;
        RECT 65.170 110.475 66.380 110.995 ;
        RECT 66.550 110.645 67.760 111.165 ;
        RECT 67.990 111.115 68.200 111.935 ;
        RECT 68.370 111.135 68.700 111.765 ;
        RECT 68.370 110.535 68.620 111.135 ;
        RECT 68.870 111.115 69.100 111.935 ;
        RECT 69.585 111.125 69.830 111.730 ;
        RECT 70.050 111.400 70.560 111.935 ;
        RECT 69.310 110.955 70.540 111.125 ;
        RECT 68.790 110.695 69.120 110.945 ;
        RECT 65.170 109.385 67.760 110.475 ;
        RECT 67.990 109.385 68.200 110.525 ;
        RECT 68.370 109.555 68.700 110.535 ;
        RECT 68.870 109.385 69.100 110.525 ;
        RECT 69.310 110.145 69.650 110.955 ;
        RECT 69.820 110.390 70.570 110.580 ;
        RECT 69.310 109.735 69.825 110.145 ;
        RECT 70.060 109.385 70.230 110.145 ;
        RECT 70.400 109.725 70.570 110.390 ;
        RECT 70.740 110.405 70.930 111.765 ;
        RECT 71.100 111.595 71.375 111.765 ;
        RECT 71.100 111.425 71.380 111.595 ;
        RECT 71.100 110.605 71.375 111.425 ;
        RECT 71.565 111.400 72.095 111.765 ;
        RECT 72.520 111.535 72.850 111.935 ;
        RECT 71.920 111.365 72.095 111.400 ;
        RECT 71.580 110.405 71.750 111.205 ;
        RECT 70.740 110.235 71.750 110.405 ;
        RECT 71.920 111.195 72.850 111.365 ;
        RECT 73.020 111.195 73.275 111.765 ;
        RECT 73.450 111.210 73.740 111.935 ;
        RECT 71.920 110.065 72.090 111.195 ;
        RECT 72.680 111.025 72.850 111.195 ;
        RECT 70.965 109.895 72.090 110.065 ;
        RECT 72.260 110.695 72.455 111.025 ;
        RECT 72.680 110.695 72.935 111.025 ;
        RECT 72.260 109.725 72.430 110.695 ;
        RECT 73.105 110.525 73.275 111.195 ;
        RECT 74.185 111.125 74.430 111.730 ;
        RECT 74.650 111.400 75.160 111.935 ;
        RECT 73.910 110.955 75.140 111.125 ;
        RECT 70.400 109.555 72.430 109.725 ;
        RECT 72.600 109.385 72.770 110.525 ;
        RECT 72.940 109.555 73.275 110.525 ;
        RECT 73.450 109.385 73.740 110.550 ;
        RECT 73.910 110.145 74.250 110.955 ;
        RECT 74.420 110.390 75.170 110.580 ;
        RECT 73.910 109.735 74.425 110.145 ;
        RECT 74.660 109.385 74.830 110.145 ;
        RECT 75.000 109.725 75.170 110.390 ;
        RECT 75.340 110.405 75.530 111.765 ;
        RECT 75.700 110.915 75.975 111.765 ;
        RECT 76.165 111.400 76.695 111.765 ;
        RECT 77.120 111.535 77.450 111.935 ;
        RECT 76.520 111.365 76.695 111.400 ;
        RECT 75.700 110.745 75.980 110.915 ;
        RECT 75.700 110.605 75.975 110.745 ;
        RECT 76.180 110.405 76.350 111.205 ;
        RECT 75.340 110.235 76.350 110.405 ;
        RECT 76.520 111.195 77.450 111.365 ;
        RECT 77.620 111.195 77.875 111.765 ;
        RECT 76.520 110.065 76.690 111.195 ;
        RECT 77.280 111.025 77.450 111.195 ;
        RECT 75.565 109.895 76.690 110.065 ;
        RECT 76.860 110.695 77.055 111.025 ;
        RECT 77.280 110.695 77.535 111.025 ;
        RECT 76.860 109.725 77.030 110.695 ;
        RECT 77.705 110.525 77.875 111.195 ;
        RECT 78.710 111.305 79.040 111.665 ;
        RECT 79.660 111.475 79.910 111.935 ;
        RECT 80.080 111.475 80.640 111.765 ;
        RECT 81.185 111.595 81.440 111.755 ;
        RECT 78.710 111.115 80.100 111.305 ;
        RECT 79.930 111.025 80.100 111.115 ;
        RECT 75.000 109.555 77.030 109.725 ;
        RECT 77.200 109.385 77.370 110.525 ;
        RECT 77.540 109.555 77.875 110.525 ;
        RECT 78.525 110.695 79.200 110.945 ;
        RECT 79.420 110.695 79.760 110.945 ;
        RECT 79.930 110.695 80.220 111.025 ;
        RECT 78.525 110.335 78.790 110.695 ;
        RECT 79.930 110.445 80.100 110.695 ;
        RECT 79.160 110.275 80.100 110.445 ;
        RECT 78.710 109.385 78.990 110.055 ;
        RECT 79.160 109.725 79.460 110.275 ;
        RECT 80.390 110.105 80.640 111.475 ;
        RECT 81.100 111.425 81.440 111.595 ;
        RECT 81.620 111.475 81.905 111.935 ;
        RECT 79.660 109.385 79.990 110.105 ;
        RECT 80.180 109.555 80.640 110.105 ;
        RECT 81.185 111.225 81.440 111.425 ;
        RECT 81.185 110.365 81.365 111.225 ;
        RECT 82.085 111.025 82.335 111.675 ;
        RECT 81.535 110.695 82.335 111.025 ;
        RECT 81.185 109.695 81.440 110.365 ;
        RECT 81.620 109.385 81.905 110.185 ;
        RECT 82.085 110.105 82.335 110.695 ;
        RECT 82.535 111.340 82.855 111.670 ;
        RECT 83.035 111.455 83.695 111.935 ;
        RECT 83.895 111.545 84.745 111.715 ;
        RECT 82.535 110.445 82.725 111.340 ;
        RECT 83.045 111.015 83.705 111.285 ;
        RECT 83.375 110.955 83.705 111.015 ;
        RECT 82.895 110.785 83.225 110.845 ;
        RECT 83.895 110.785 84.065 111.545 ;
        RECT 85.305 111.475 85.625 111.935 ;
        RECT 85.825 111.295 86.075 111.725 ;
        RECT 86.365 111.495 86.775 111.935 ;
        RECT 86.945 111.555 87.960 111.755 ;
        RECT 84.235 111.125 85.485 111.295 ;
        RECT 84.235 111.005 84.565 111.125 ;
        RECT 82.895 110.615 84.795 110.785 ;
        RECT 82.535 110.275 84.455 110.445 ;
        RECT 82.535 110.255 82.855 110.275 ;
        RECT 82.085 109.595 82.415 110.105 ;
        RECT 82.685 109.645 82.855 110.255 ;
        RECT 84.625 110.105 84.795 110.615 ;
        RECT 84.965 110.545 85.145 110.955 ;
        RECT 85.315 110.365 85.485 111.125 ;
        RECT 83.025 109.385 83.355 110.075 ;
        RECT 83.585 109.935 84.795 110.105 ;
        RECT 84.965 110.055 85.485 110.365 ;
        RECT 85.655 110.955 86.075 111.295 ;
        RECT 86.365 110.955 86.775 111.285 ;
        RECT 85.655 110.185 85.845 110.955 ;
        RECT 86.945 110.825 87.115 111.555 ;
        RECT 88.260 111.385 88.430 111.715 ;
        RECT 88.600 111.555 88.930 111.935 ;
        RECT 87.285 111.005 87.635 111.375 ;
        RECT 86.945 110.785 87.365 110.825 ;
        RECT 86.015 110.615 87.365 110.785 ;
        RECT 86.015 110.455 86.265 110.615 ;
        RECT 86.775 110.185 87.025 110.445 ;
        RECT 85.655 109.935 87.025 110.185 ;
        RECT 83.585 109.645 83.825 109.935 ;
        RECT 84.625 109.855 84.795 109.935 ;
        RECT 84.025 109.385 84.445 109.765 ;
        RECT 84.625 109.605 85.255 109.855 ;
        RECT 85.725 109.385 86.055 109.765 ;
        RECT 86.225 109.645 86.395 109.935 ;
        RECT 87.195 109.770 87.365 110.615 ;
        RECT 87.815 110.445 88.035 111.315 ;
        RECT 88.260 111.195 88.955 111.385 ;
        RECT 87.535 110.065 88.035 110.445 ;
        RECT 88.205 110.395 88.615 111.015 ;
        RECT 88.785 110.225 88.955 111.195 ;
        RECT 88.260 110.055 88.955 110.225 ;
        RECT 86.575 109.385 86.955 109.765 ;
        RECT 87.195 109.600 88.025 109.770 ;
        RECT 88.260 109.555 88.430 110.055 ;
        RECT 88.600 109.385 88.930 109.885 ;
        RECT 89.145 109.555 89.370 111.675 ;
        RECT 89.540 111.555 89.870 111.935 ;
        RECT 90.040 111.385 90.210 111.675 ;
        RECT 89.545 111.215 90.210 111.385 ;
        RECT 89.545 110.225 89.775 111.215 ;
        RECT 90.475 111.195 90.730 111.765 ;
        RECT 90.900 111.535 91.230 111.935 ;
        RECT 91.655 111.400 92.185 111.765 ;
        RECT 92.375 111.595 92.650 111.765 ;
        RECT 92.370 111.425 92.650 111.595 ;
        RECT 91.655 111.365 91.830 111.400 ;
        RECT 90.900 111.195 91.830 111.365 ;
        RECT 89.945 110.395 90.295 111.045 ;
        RECT 90.475 110.525 90.645 111.195 ;
        RECT 90.900 111.025 91.070 111.195 ;
        RECT 90.815 110.695 91.070 111.025 ;
        RECT 91.295 110.695 91.490 111.025 ;
        RECT 89.545 110.055 90.210 110.225 ;
        RECT 89.540 109.385 89.870 109.885 ;
        RECT 90.040 109.555 90.210 110.055 ;
        RECT 90.475 109.555 90.810 110.525 ;
        RECT 90.980 109.385 91.150 110.525 ;
        RECT 91.320 109.725 91.490 110.695 ;
        RECT 91.660 110.065 91.830 111.195 ;
        RECT 92.000 110.405 92.170 111.205 ;
        RECT 92.375 110.605 92.650 111.425 ;
        RECT 92.820 110.405 93.010 111.765 ;
        RECT 93.190 111.400 93.700 111.935 ;
        RECT 93.920 111.125 94.165 111.730 ;
        RECT 94.885 111.125 95.130 111.730 ;
        RECT 95.350 111.400 95.860 111.935 ;
        RECT 93.210 110.955 94.440 111.125 ;
        RECT 92.000 110.235 93.010 110.405 ;
        RECT 93.180 110.390 93.930 110.580 ;
        RECT 91.660 109.895 92.785 110.065 ;
        RECT 93.180 109.725 93.350 110.390 ;
        RECT 94.100 110.145 94.440 110.955 ;
        RECT 91.320 109.555 93.350 109.725 ;
        RECT 93.520 109.385 93.690 110.145 ;
        RECT 93.925 109.735 94.440 110.145 ;
        RECT 94.610 110.955 95.840 111.125 ;
        RECT 94.610 110.145 94.950 110.955 ;
        RECT 95.120 110.390 95.870 110.580 ;
        RECT 94.610 109.735 95.125 110.145 ;
        RECT 95.360 109.385 95.530 110.145 ;
        RECT 95.700 109.725 95.870 110.390 ;
        RECT 96.040 110.405 96.230 111.765 ;
        RECT 96.400 111.255 96.675 111.765 ;
        RECT 96.865 111.400 97.395 111.765 ;
        RECT 97.820 111.535 98.150 111.935 ;
        RECT 97.220 111.365 97.395 111.400 ;
        RECT 96.400 111.085 96.680 111.255 ;
        RECT 96.400 110.605 96.675 111.085 ;
        RECT 96.880 110.405 97.050 111.205 ;
        RECT 96.040 110.235 97.050 110.405 ;
        RECT 97.220 111.195 98.150 111.365 ;
        RECT 98.320 111.195 98.575 111.765 ;
        RECT 99.210 111.210 99.500 111.935 ;
        RECT 100.135 111.390 105.480 111.935 ;
        RECT 105.655 111.390 111.000 111.935 ;
        RECT 97.220 110.065 97.390 111.195 ;
        RECT 97.980 111.025 98.150 111.195 ;
        RECT 96.265 109.895 97.390 110.065 ;
        RECT 97.560 110.695 97.755 111.025 ;
        RECT 97.980 110.695 98.235 111.025 ;
        RECT 97.560 109.725 97.730 110.695 ;
        RECT 98.405 110.525 98.575 111.195 ;
        RECT 95.700 109.555 97.730 109.725 ;
        RECT 97.900 109.385 98.070 110.525 ;
        RECT 98.240 109.555 98.575 110.525 ;
        RECT 99.210 109.385 99.500 110.550 ;
        RECT 101.725 109.820 102.075 111.070 ;
        RECT 103.555 110.560 103.895 111.390 ;
        RECT 107.245 109.820 107.595 111.070 ;
        RECT 109.075 110.560 109.415 111.390 ;
        RECT 111.170 111.185 112.380 111.935 ;
        RECT 111.170 110.475 111.690 111.015 ;
        RECT 111.860 110.645 112.380 111.185 ;
        RECT 100.135 109.385 105.480 109.820 ;
        RECT 105.655 109.385 111.000 109.820 ;
        RECT 111.170 109.385 112.380 110.475 ;
        RECT 18.165 109.215 112.465 109.385 ;
        RECT 18.250 108.125 19.460 109.215 ;
        RECT 20.095 108.780 25.440 109.215 ;
        RECT 25.615 108.780 30.960 109.215 ;
        RECT 18.250 107.415 18.770 107.955 ;
        RECT 18.940 107.585 19.460 108.125 ;
        RECT 21.685 107.530 22.035 108.780 ;
        RECT 18.250 106.665 19.460 107.415 ;
        RECT 23.515 107.210 23.855 108.040 ;
        RECT 27.205 107.530 27.555 108.780 ;
        RECT 31.170 108.075 31.400 109.215 ;
        RECT 31.570 108.065 31.900 109.045 ;
        RECT 32.070 108.075 32.280 109.215 ;
        RECT 32.510 108.495 32.970 109.045 ;
        RECT 33.160 108.495 33.490 109.215 ;
        RECT 29.035 107.210 29.375 108.040 ;
        RECT 31.150 107.655 31.480 107.905 ;
        RECT 20.095 106.665 25.440 107.210 ;
        RECT 25.615 106.665 30.960 107.210 ;
        RECT 31.170 106.665 31.400 107.485 ;
        RECT 31.650 107.465 31.900 108.065 ;
        RECT 31.570 106.835 31.900 107.465 ;
        RECT 32.070 106.665 32.280 107.485 ;
        RECT 32.510 107.125 32.760 108.495 ;
        RECT 33.690 108.325 33.990 108.875 ;
        RECT 34.160 108.545 34.440 109.215 ;
        RECT 33.050 108.155 33.990 108.325 ;
        RECT 33.050 107.905 33.220 108.155 ;
        RECT 34.360 107.905 34.625 108.265 ;
        RECT 34.810 108.050 35.100 109.215 ;
        RECT 36.190 108.455 36.705 108.865 ;
        RECT 36.940 108.455 37.110 109.215 ;
        RECT 37.280 108.875 39.310 109.045 ;
        RECT 32.930 107.575 33.220 107.905 ;
        RECT 33.390 107.655 33.730 107.905 ;
        RECT 33.950 107.655 34.625 107.905 ;
        RECT 33.050 107.485 33.220 107.575 ;
        RECT 36.190 107.645 36.530 108.455 ;
        RECT 37.280 108.210 37.450 108.875 ;
        RECT 37.845 108.535 38.970 108.705 ;
        RECT 36.700 108.020 37.450 108.210 ;
        RECT 37.620 108.195 38.630 108.365 ;
        RECT 33.050 107.295 34.440 107.485 ;
        RECT 36.190 107.475 37.420 107.645 ;
        RECT 32.510 106.835 33.070 107.125 ;
        RECT 33.240 106.665 33.490 107.125 ;
        RECT 34.110 106.935 34.440 107.295 ;
        RECT 34.810 106.665 35.100 107.390 ;
        RECT 36.465 106.870 36.710 107.475 ;
        RECT 36.930 106.665 37.440 107.200 ;
        RECT 37.620 106.835 37.810 108.195 ;
        RECT 37.980 107.855 38.255 107.995 ;
        RECT 37.980 107.685 38.260 107.855 ;
        RECT 37.980 106.835 38.255 107.685 ;
        RECT 38.460 107.395 38.630 108.195 ;
        RECT 38.800 107.405 38.970 108.535 ;
        RECT 39.140 107.905 39.310 108.875 ;
        RECT 39.480 108.075 39.650 109.215 ;
        RECT 39.820 108.075 40.155 109.045 ;
        RECT 39.140 107.575 39.335 107.905 ;
        RECT 39.560 107.575 39.815 107.905 ;
        RECT 39.560 107.405 39.730 107.575 ;
        RECT 39.985 107.405 40.155 108.075 ;
        RECT 40.330 108.455 40.845 108.865 ;
        RECT 41.080 108.455 41.250 109.215 ;
        RECT 41.420 108.875 43.450 109.045 ;
        RECT 40.330 107.645 40.670 108.455 ;
        RECT 41.420 108.210 41.590 108.875 ;
        RECT 41.985 108.535 43.110 108.705 ;
        RECT 40.840 108.020 41.590 108.210 ;
        RECT 41.760 108.195 42.770 108.365 ;
        RECT 40.330 107.475 41.560 107.645 ;
        RECT 38.800 107.235 39.730 107.405 ;
        RECT 38.800 107.200 38.975 107.235 ;
        RECT 38.445 106.835 38.975 107.200 ;
        RECT 39.400 106.665 39.730 107.065 ;
        RECT 39.900 106.835 40.155 107.405 ;
        RECT 40.605 106.870 40.850 107.475 ;
        RECT 41.070 106.665 41.580 107.200 ;
        RECT 41.760 106.835 41.950 108.195 ;
        RECT 42.120 107.855 42.395 107.995 ;
        RECT 42.120 107.685 42.400 107.855 ;
        RECT 42.120 106.835 42.395 107.685 ;
        RECT 42.600 107.395 42.770 108.195 ;
        RECT 42.940 107.405 43.110 108.535 ;
        RECT 43.280 107.905 43.450 108.875 ;
        RECT 43.620 108.075 43.790 109.215 ;
        RECT 43.960 108.075 44.295 109.045 ;
        RECT 43.280 107.575 43.475 107.905 ;
        RECT 43.700 107.575 43.955 107.905 ;
        RECT 43.700 107.405 43.870 107.575 ;
        RECT 44.125 107.405 44.295 108.075 ;
        RECT 44.845 108.235 45.100 108.905 ;
        RECT 45.280 108.415 45.565 109.215 ;
        RECT 45.745 108.495 46.075 109.005 ;
        RECT 44.845 107.855 45.025 108.235 ;
        RECT 45.745 107.905 45.995 108.495 ;
        RECT 46.345 108.345 46.515 108.955 ;
        RECT 46.685 108.525 47.015 109.215 ;
        RECT 47.245 108.665 47.485 108.955 ;
        RECT 47.685 108.835 48.105 109.215 ;
        RECT 48.285 108.745 48.915 108.995 ;
        RECT 49.385 108.835 49.715 109.215 ;
        RECT 48.285 108.665 48.455 108.745 ;
        RECT 49.885 108.665 50.055 108.955 ;
        RECT 50.235 108.835 50.615 109.215 ;
        RECT 50.855 108.830 51.685 109.000 ;
        RECT 47.245 108.495 48.455 108.665 ;
        RECT 44.760 107.685 45.025 107.855 ;
        RECT 42.940 107.235 43.870 107.405 ;
        RECT 42.940 107.200 43.115 107.235 ;
        RECT 42.585 106.835 43.115 107.200 ;
        RECT 43.540 106.665 43.870 107.065 ;
        RECT 44.040 106.835 44.295 107.405 ;
        RECT 44.845 107.375 45.025 107.685 ;
        RECT 45.195 107.575 45.995 107.905 ;
        RECT 44.845 106.845 45.100 107.375 ;
        RECT 45.280 106.665 45.565 107.125 ;
        RECT 45.745 106.925 45.995 107.575 ;
        RECT 46.195 108.325 46.515 108.345 ;
        RECT 46.195 108.155 48.115 108.325 ;
        RECT 46.195 107.260 46.385 108.155 ;
        RECT 48.285 107.985 48.455 108.495 ;
        RECT 48.625 108.235 49.145 108.545 ;
        RECT 46.555 107.815 48.455 107.985 ;
        RECT 46.555 107.755 46.885 107.815 ;
        RECT 47.035 107.585 47.365 107.645 ;
        RECT 46.705 107.315 47.365 107.585 ;
        RECT 46.195 106.930 46.515 107.260 ;
        RECT 46.695 106.665 47.355 107.145 ;
        RECT 47.555 107.055 47.725 107.815 ;
        RECT 48.625 107.645 48.805 108.055 ;
        RECT 47.895 107.475 48.225 107.595 ;
        RECT 48.975 107.475 49.145 108.235 ;
        RECT 47.895 107.305 49.145 107.475 ;
        RECT 49.315 108.415 50.685 108.665 ;
        RECT 49.315 107.645 49.505 108.415 ;
        RECT 50.435 108.155 50.685 108.415 ;
        RECT 49.675 107.985 49.925 108.145 ;
        RECT 50.855 107.985 51.025 108.830 ;
        RECT 51.920 108.545 52.090 109.045 ;
        RECT 52.260 108.715 52.590 109.215 ;
        RECT 51.195 108.155 51.695 108.535 ;
        RECT 51.920 108.375 52.615 108.545 ;
        RECT 49.675 107.815 51.025 107.985 ;
        RECT 50.605 107.775 51.025 107.815 ;
        RECT 49.315 107.305 49.735 107.645 ;
        RECT 50.025 107.315 50.435 107.645 ;
        RECT 47.555 106.885 48.405 107.055 ;
        RECT 48.965 106.665 49.285 107.125 ;
        RECT 49.485 106.875 49.735 107.305 ;
        RECT 50.025 106.665 50.435 107.105 ;
        RECT 50.605 107.045 50.775 107.775 ;
        RECT 50.945 107.225 51.295 107.595 ;
        RECT 51.475 107.285 51.695 108.155 ;
        RECT 51.865 107.585 52.275 108.205 ;
        RECT 52.445 107.405 52.615 108.375 ;
        RECT 51.920 107.215 52.615 107.405 ;
        RECT 50.605 106.845 51.620 107.045 ;
        RECT 51.920 106.885 52.090 107.215 ;
        RECT 52.260 106.665 52.590 107.045 ;
        RECT 52.805 106.925 53.030 109.045 ;
        RECT 53.200 108.715 53.530 109.215 ;
        RECT 53.700 108.545 53.870 109.045 ;
        RECT 53.205 108.375 53.870 108.545 ;
        RECT 53.205 107.385 53.435 108.375 ;
        RECT 53.605 107.555 53.955 108.205 ;
        RECT 54.590 108.125 56.260 109.215 ;
        RECT 56.430 108.455 56.945 108.865 ;
        RECT 57.180 108.455 57.350 109.215 ;
        RECT 57.520 108.875 59.550 109.045 ;
        RECT 54.590 107.605 55.340 108.125 ;
        RECT 55.510 107.435 56.260 107.955 ;
        RECT 56.430 107.645 56.770 108.455 ;
        RECT 57.520 108.210 57.690 108.875 ;
        RECT 58.085 108.535 59.210 108.705 ;
        RECT 56.940 108.020 57.690 108.210 ;
        RECT 57.860 108.195 58.870 108.365 ;
        RECT 56.430 107.475 57.660 107.645 ;
        RECT 53.205 107.215 53.870 107.385 ;
        RECT 53.200 106.665 53.530 107.045 ;
        RECT 53.700 106.925 53.870 107.215 ;
        RECT 54.590 106.665 56.260 107.435 ;
        RECT 56.705 106.870 56.950 107.475 ;
        RECT 57.170 106.665 57.680 107.200 ;
        RECT 57.860 106.835 58.050 108.195 ;
        RECT 58.220 107.855 58.495 107.995 ;
        RECT 58.220 107.685 58.500 107.855 ;
        RECT 58.220 106.835 58.495 107.685 ;
        RECT 58.700 107.395 58.870 108.195 ;
        RECT 59.040 107.405 59.210 108.535 ;
        RECT 59.380 107.905 59.550 108.875 ;
        RECT 59.720 108.075 59.890 109.215 ;
        RECT 60.060 108.075 60.395 109.045 ;
        RECT 59.380 107.575 59.575 107.905 ;
        RECT 59.800 107.575 60.055 107.905 ;
        RECT 59.800 107.405 59.970 107.575 ;
        RECT 60.225 107.405 60.395 108.075 ;
        RECT 60.570 108.050 60.860 109.215 ;
        RECT 61.120 108.285 61.290 109.045 ;
        RECT 61.505 108.455 61.835 109.215 ;
        RECT 61.120 108.115 61.835 108.285 ;
        RECT 62.005 108.140 62.260 109.045 ;
        RECT 61.030 107.565 61.385 107.935 ;
        RECT 61.665 107.905 61.835 108.115 ;
        RECT 61.665 107.575 61.920 107.905 ;
        RECT 59.040 107.235 59.970 107.405 ;
        RECT 59.040 107.200 59.215 107.235 ;
        RECT 58.685 106.835 59.215 107.200 ;
        RECT 59.640 106.665 59.970 107.065 ;
        RECT 60.140 106.835 60.395 107.405 ;
        RECT 60.570 106.665 60.860 107.390 ;
        RECT 61.665 107.385 61.835 107.575 ;
        RECT 62.090 107.410 62.260 108.140 ;
        RECT 62.435 108.065 62.695 109.215 ;
        RECT 62.870 108.125 65.460 109.215 ;
        RECT 66.005 108.875 66.260 108.905 ;
        RECT 65.920 108.705 66.260 108.875 ;
        RECT 66.005 108.235 66.260 108.705 ;
        RECT 66.440 108.415 66.725 109.215 ;
        RECT 66.905 108.495 67.235 109.005 ;
        RECT 62.870 107.605 64.080 108.125 ;
        RECT 61.120 107.215 61.835 107.385 ;
        RECT 61.120 106.835 61.290 107.215 ;
        RECT 61.505 106.665 61.835 107.045 ;
        RECT 62.005 106.835 62.260 107.410 ;
        RECT 62.435 106.665 62.695 107.505 ;
        RECT 64.250 107.435 65.460 107.955 ;
        RECT 62.870 106.665 65.460 107.435 ;
        RECT 66.005 107.375 66.185 108.235 ;
        RECT 66.905 107.905 67.155 108.495 ;
        RECT 67.505 108.345 67.675 108.955 ;
        RECT 67.845 108.525 68.175 109.215 ;
        RECT 68.405 108.665 68.645 108.955 ;
        RECT 68.845 108.835 69.265 109.215 ;
        RECT 69.445 108.745 70.075 108.995 ;
        RECT 70.545 108.835 70.875 109.215 ;
        RECT 69.445 108.665 69.615 108.745 ;
        RECT 71.045 108.665 71.215 108.955 ;
        RECT 71.395 108.835 71.775 109.215 ;
        RECT 72.015 108.830 72.845 109.000 ;
        RECT 68.405 108.495 69.615 108.665 ;
        RECT 66.355 107.575 67.155 107.905 ;
        RECT 66.005 106.845 66.260 107.375 ;
        RECT 66.440 106.665 66.725 107.125 ;
        RECT 66.905 106.925 67.155 107.575 ;
        RECT 67.355 108.325 67.675 108.345 ;
        RECT 67.355 108.155 69.275 108.325 ;
        RECT 67.355 107.260 67.545 108.155 ;
        RECT 69.445 107.985 69.615 108.495 ;
        RECT 69.785 108.235 70.305 108.545 ;
        RECT 67.715 107.815 69.615 107.985 ;
        RECT 67.715 107.755 68.045 107.815 ;
        RECT 68.195 107.585 68.525 107.645 ;
        RECT 67.865 107.315 68.525 107.585 ;
        RECT 67.355 106.930 67.675 107.260 ;
        RECT 67.855 106.665 68.515 107.145 ;
        RECT 68.715 107.055 68.885 107.815 ;
        RECT 69.785 107.645 69.965 108.055 ;
        RECT 69.055 107.475 69.385 107.595 ;
        RECT 70.135 107.475 70.305 108.235 ;
        RECT 69.055 107.305 70.305 107.475 ;
        RECT 70.475 108.415 71.845 108.665 ;
        RECT 70.475 107.645 70.665 108.415 ;
        RECT 71.595 108.155 71.845 108.415 ;
        RECT 70.835 107.985 71.085 108.145 ;
        RECT 72.015 107.985 72.185 108.830 ;
        RECT 73.080 108.545 73.250 109.045 ;
        RECT 73.420 108.715 73.750 109.215 ;
        RECT 72.355 108.155 72.855 108.535 ;
        RECT 73.080 108.375 73.775 108.545 ;
        RECT 70.835 107.815 72.185 107.985 ;
        RECT 71.765 107.775 72.185 107.815 ;
        RECT 70.475 107.305 70.895 107.645 ;
        RECT 71.185 107.315 71.595 107.645 ;
        RECT 68.715 106.885 69.565 107.055 ;
        RECT 70.125 106.665 70.445 107.125 ;
        RECT 70.645 106.875 70.895 107.305 ;
        RECT 71.185 106.665 71.595 107.105 ;
        RECT 71.765 107.045 71.935 107.775 ;
        RECT 72.105 107.225 72.455 107.595 ;
        RECT 72.635 107.285 72.855 108.155 ;
        RECT 73.025 107.585 73.435 108.205 ;
        RECT 73.605 107.405 73.775 108.375 ;
        RECT 73.080 107.215 73.775 107.405 ;
        RECT 71.765 106.845 72.780 107.045 ;
        RECT 73.080 106.885 73.250 107.215 ;
        RECT 73.420 106.665 73.750 107.045 ;
        RECT 73.965 106.925 74.190 109.045 ;
        RECT 74.360 108.715 74.690 109.215 ;
        RECT 74.860 108.545 75.030 109.045 ;
        RECT 74.365 108.375 75.030 108.545 ;
        RECT 75.380 108.545 75.550 109.045 ;
        RECT 75.720 108.715 76.050 109.215 ;
        RECT 75.380 108.375 76.045 108.545 ;
        RECT 74.365 107.385 74.595 108.375 ;
        RECT 74.765 107.555 75.115 108.205 ;
        RECT 75.295 107.555 75.645 108.205 ;
        RECT 75.815 107.385 76.045 108.375 ;
        RECT 74.365 107.215 75.030 107.385 ;
        RECT 74.360 106.665 74.690 107.045 ;
        RECT 74.860 106.925 75.030 107.215 ;
        RECT 75.380 107.215 76.045 107.385 ;
        RECT 75.380 106.925 75.550 107.215 ;
        RECT 75.720 106.665 76.050 107.045 ;
        RECT 76.220 106.925 76.445 109.045 ;
        RECT 76.660 108.715 76.990 109.215 ;
        RECT 77.160 108.545 77.330 109.045 ;
        RECT 77.565 108.830 78.395 109.000 ;
        RECT 78.635 108.835 79.015 109.215 ;
        RECT 76.635 108.375 77.330 108.545 ;
        RECT 76.635 107.405 76.805 108.375 ;
        RECT 76.975 107.585 77.385 108.205 ;
        RECT 77.555 108.155 78.055 108.535 ;
        RECT 76.635 107.215 77.330 107.405 ;
        RECT 77.555 107.285 77.775 108.155 ;
        RECT 78.225 107.985 78.395 108.830 ;
        RECT 79.195 108.665 79.365 108.955 ;
        RECT 79.535 108.835 79.865 109.215 ;
        RECT 80.335 108.745 80.965 108.995 ;
        RECT 81.145 108.835 81.565 109.215 ;
        RECT 80.795 108.665 80.965 108.745 ;
        RECT 81.765 108.665 82.005 108.955 ;
        RECT 78.565 108.415 79.935 108.665 ;
        RECT 78.565 108.155 78.815 108.415 ;
        RECT 79.325 107.985 79.575 108.145 ;
        RECT 78.225 107.815 79.575 107.985 ;
        RECT 78.225 107.775 78.645 107.815 ;
        RECT 77.955 107.225 78.305 107.595 ;
        RECT 76.660 106.665 76.990 107.045 ;
        RECT 77.160 106.885 77.330 107.215 ;
        RECT 78.475 107.045 78.645 107.775 ;
        RECT 79.745 107.645 79.935 108.415 ;
        RECT 78.815 107.315 79.225 107.645 ;
        RECT 79.515 107.305 79.935 107.645 ;
        RECT 80.105 108.235 80.625 108.545 ;
        RECT 80.795 108.495 82.005 108.665 ;
        RECT 82.235 108.525 82.565 109.215 ;
        RECT 80.105 107.475 80.275 108.235 ;
        RECT 80.445 107.645 80.625 108.055 ;
        RECT 80.795 107.985 80.965 108.495 ;
        RECT 82.735 108.345 82.905 108.955 ;
        RECT 83.175 108.495 83.505 109.005 ;
        RECT 82.735 108.325 83.055 108.345 ;
        RECT 81.135 108.155 83.055 108.325 ;
        RECT 80.795 107.815 82.695 107.985 ;
        RECT 81.025 107.475 81.355 107.595 ;
        RECT 80.105 107.305 81.355 107.475 ;
        RECT 77.630 106.845 78.645 107.045 ;
        RECT 78.815 106.665 79.225 107.105 ;
        RECT 79.515 106.875 79.765 107.305 ;
        RECT 79.965 106.665 80.285 107.125 ;
        RECT 81.525 107.055 81.695 107.815 ;
        RECT 82.365 107.755 82.695 107.815 ;
        RECT 81.885 107.585 82.215 107.645 ;
        RECT 81.885 107.315 82.545 107.585 ;
        RECT 82.865 107.260 83.055 108.155 ;
        RECT 80.845 106.885 81.695 107.055 ;
        RECT 81.895 106.665 82.555 107.145 ;
        RECT 82.735 106.930 83.055 107.260 ;
        RECT 83.255 107.905 83.505 108.495 ;
        RECT 83.685 108.415 83.970 109.215 ;
        RECT 84.150 108.875 84.405 108.905 ;
        RECT 84.150 108.705 84.490 108.875 ;
        RECT 84.150 108.235 84.405 108.705 ;
        RECT 83.255 107.575 84.055 107.905 ;
        RECT 83.255 106.925 83.505 107.575 ;
        RECT 84.225 107.375 84.405 108.235 ;
        RECT 85.010 108.075 85.220 109.215 ;
        RECT 85.390 108.065 85.720 109.045 ;
        RECT 85.890 108.075 86.120 109.215 ;
        RECT 83.685 106.665 83.970 107.125 ;
        RECT 84.150 106.845 84.405 107.375 ;
        RECT 85.010 106.665 85.220 107.485 ;
        RECT 85.390 107.465 85.640 108.065 ;
        RECT 86.330 108.050 86.620 109.215 ;
        RECT 86.790 108.245 87.100 109.045 ;
        RECT 87.270 108.415 87.580 109.215 ;
        RECT 87.750 108.585 88.010 109.045 ;
        RECT 88.180 108.755 88.435 109.215 ;
        RECT 88.610 108.585 88.870 109.045 ;
        RECT 87.750 108.415 88.870 108.585 ;
        RECT 88.230 108.365 88.400 108.415 ;
        RECT 86.790 108.075 87.820 108.245 ;
        RECT 85.810 107.655 86.140 107.905 ;
        RECT 85.390 106.835 85.720 107.465 ;
        RECT 85.890 106.665 86.120 107.485 ;
        RECT 86.330 106.665 86.620 107.390 ;
        RECT 86.790 107.165 86.960 108.075 ;
        RECT 87.130 107.335 87.480 107.905 ;
        RECT 87.650 107.825 87.820 108.075 ;
        RECT 88.610 108.165 88.870 108.415 ;
        RECT 89.040 108.345 89.325 109.215 ;
        RECT 88.610 107.995 89.365 108.165 ;
        RECT 89.590 108.075 89.820 109.215 ;
        RECT 89.990 108.065 90.320 109.045 ;
        RECT 90.490 108.075 90.700 109.215 ;
        RECT 91.020 108.545 91.190 109.045 ;
        RECT 91.360 108.715 91.690 109.215 ;
        RECT 91.020 108.375 91.685 108.545 ;
        RECT 87.650 107.655 88.790 107.825 ;
        RECT 88.960 107.485 89.365 107.995 ;
        RECT 89.570 107.655 89.900 107.905 ;
        RECT 87.715 107.315 89.365 107.485 ;
        RECT 86.790 106.835 87.090 107.165 ;
        RECT 87.260 106.665 87.535 107.145 ;
        RECT 87.715 106.925 88.010 107.315 ;
        RECT 88.180 106.665 88.435 107.145 ;
        RECT 88.610 106.925 88.870 107.315 ;
        RECT 89.040 106.665 89.320 107.145 ;
        RECT 89.590 106.665 89.820 107.485 ;
        RECT 90.070 107.465 90.320 108.065 ;
        RECT 90.935 107.555 91.285 108.205 ;
        RECT 89.990 106.835 90.320 107.465 ;
        RECT 90.490 106.665 90.700 107.485 ;
        RECT 91.455 107.385 91.685 108.375 ;
        RECT 91.020 107.215 91.685 107.385 ;
        RECT 91.020 106.925 91.190 107.215 ;
        RECT 91.360 106.665 91.690 107.045 ;
        RECT 91.860 106.925 92.085 109.045 ;
        RECT 92.300 108.715 92.630 109.215 ;
        RECT 92.800 108.545 92.970 109.045 ;
        RECT 93.205 108.830 94.035 109.000 ;
        RECT 94.275 108.835 94.655 109.215 ;
        RECT 92.275 108.375 92.970 108.545 ;
        RECT 92.275 107.405 92.445 108.375 ;
        RECT 92.615 107.585 93.025 108.205 ;
        RECT 93.195 108.155 93.695 108.535 ;
        RECT 92.275 107.215 92.970 107.405 ;
        RECT 93.195 107.285 93.415 108.155 ;
        RECT 93.865 107.985 94.035 108.830 ;
        RECT 94.835 108.665 95.005 108.955 ;
        RECT 95.175 108.835 95.505 109.215 ;
        RECT 95.975 108.745 96.605 108.995 ;
        RECT 96.785 108.835 97.205 109.215 ;
        RECT 96.435 108.665 96.605 108.745 ;
        RECT 97.405 108.665 97.645 108.955 ;
        RECT 94.205 108.415 95.575 108.665 ;
        RECT 94.205 108.155 94.455 108.415 ;
        RECT 94.965 107.985 95.215 108.145 ;
        RECT 93.865 107.815 95.215 107.985 ;
        RECT 93.865 107.775 94.285 107.815 ;
        RECT 93.595 107.225 93.945 107.595 ;
        RECT 92.300 106.665 92.630 107.045 ;
        RECT 92.800 106.885 92.970 107.215 ;
        RECT 94.115 107.045 94.285 107.775 ;
        RECT 95.385 107.645 95.575 108.415 ;
        RECT 94.455 107.315 94.865 107.645 ;
        RECT 95.155 107.305 95.575 107.645 ;
        RECT 95.745 108.235 96.265 108.545 ;
        RECT 96.435 108.495 97.645 108.665 ;
        RECT 97.875 108.525 98.205 109.215 ;
        RECT 95.745 107.475 95.915 108.235 ;
        RECT 96.085 107.645 96.265 108.055 ;
        RECT 96.435 107.985 96.605 108.495 ;
        RECT 98.375 108.345 98.545 108.955 ;
        RECT 98.815 108.495 99.145 109.005 ;
        RECT 98.375 108.325 98.695 108.345 ;
        RECT 96.775 108.155 98.695 108.325 ;
        RECT 96.435 107.815 98.335 107.985 ;
        RECT 96.665 107.475 96.995 107.595 ;
        RECT 95.745 107.305 96.995 107.475 ;
        RECT 93.270 106.845 94.285 107.045 ;
        RECT 94.455 106.665 94.865 107.105 ;
        RECT 95.155 106.875 95.405 107.305 ;
        RECT 95.605 106.665 95.925 107.125 ;
        RECT 97.165 107.055 97.335 107.815 ;
        RECT 98.005 107.755 98.335 107.815 ;
        RECT 97.525 107.585 97.855 107.645 ;
        RECT 97.525 107.315 98.185 107.585 ;
        RECT 98.505 107.260 98.695 108.155 ;
        RECT 96.485 106.885 97.335 107.055 ;
        RECT 97.535 106.665 98.195 107.145 ;
        RECT 98.375 106.930 98.695 107.260 ;
        RECT 98.895 107.905 99.145 108.495 ;
        RECT 99.325 108.415 99.610 109.215 ;
        RECT 99.790 108.875 100.045 108.905 ;
        RECT 99.790 108.705 100.130 108.875 ;
        RECT 99.790 108.235 100.045 108.705 ;
        RECT 98.895 107.575 99.695 107.905 ;
        RECT 98.895 106.925 99.145 107.575 ;
        RECT 99.865 107.375 100.045 108.235 ;
        RECT 100.650 108.075 100.860 109.215 ;
        RECT 101.030 108.065 101.360 109.045 ;
        RECT 101.530 108.075 101.760 109.215 ;
        RECT 101.970 108.125 105.480 109.215 ;
        RECT 105.655 108.780 111.000 109.215 ;
        RECT 99.325 106.665 99.610 107.125 ;
        RECT 99.790 106.845 100.045 107.375 ;
        RECT 100.650 106.665 100.860 107.485 ;
        RECT 101.030 107.465 101.280 108.065 ;
        RECT 101.450 107.655 101.780 107.905 ;
        RECT 101.970 107.605 103.660 108.125 ;
        RECT 101.030 106.835 101.360 107.465 ;
        RECT 101.530 106.665 101.760 107.485 ;
        RECT 103.830 107.435 105.480 107.955 ;
        RECT 107.245 107.530 107.595 108.780 ;
        RECT 111.170 108.125 112.380 109.215 ;
        RECT 101.970 106.665 105.480 107.435 ;
        RECT 109.075 107.210 109.415 108.040 ;
        RECT 111.170 107.585 111.690 108.125 ;
        RECT 111.860 107.415 112.380 107.955 ;
        RECT 105.655 106.665 111.000 107.210 ;
        RECT 111.170 106.665 112.380 107.415 ;
        RECT 18.165 106.495 112.465 106.665 ;
        RECT 18.250 105.745 19.460 106.495 ;
        RECT 18.250 105.205 18.770 105.745 ;
        RECT 20.090 105.725 21.760 106.495 ;
        RECT 21.930 105.770 22.220 106.495 ;
        RECT 23.310 105.725 26.820 106.495 ;
        RECT 26.995 105.950 32.340 106.495 ;
        RECT 32.515 105.950 37.860 106.495 ;
        RECT 38.405 106.155 38.660 106.315 ;
        RECT 38.320 105.985 38.660 106.155 ;
        RECT 38.840 106.035 39.125 106.495 ;
        RECT 18.940 105.035 19.460 105.575 ;
        RECT 18.250 103.945 19.460 105.035 ;
        RECT 20.090 105.035 20.840 105.555 ;
        RECT 21.010 105.205 21.760 105.725 ;
        RECT 20.090 103.945 21.760 105.035 ;
        RECT 21.930 103.945 22.220 105.110 ;
        RECT 23.310 105.035 25.000 105.555 ;
        RECT 25.170 105.205 26.820 105.725 ;
        RECT 23.310 103.945 26.820 105.035 ;
        RECT 28.585 104.380 28.935 105.630 ;
        RECT 30.415 105.120 30.755 105.950 ;
        RECT 34.105 104.380 34.455 105.630 ;
        RECT 35.935 105.120 36.275 105.950 ;
        RECT 38.405 105.785 38.660 105.985 ;
        RECT 38.405 104.925 38.585 105.785 ;
        RECT 39.305 105.585 39.555 106.235 ;
        RECT 38.755 105.255 39.555 105.585 ;
        RECT 26.995 103.945 32.340 104.380 ;
        RECT 32.515 103.945 37.860 104.380 ;
        RECT 38.405 104.255 38.660 104.925 ;
        RECT 38.840 103.945 39.125 104.745 ;
        RECT 39.305 104.665 39.555 105.255 ;
        RECT 39.755 105.900 40.075 106.230 ;
        RECT 40.255 106.015 40.915 106.495 ;
        RECT 41.115 106.105 41.965 106.275 ;
        RECT 39.755 105.005 39.945 105.900 ;
        RECT 40.265 105.575 40.925 105.845 ;
        RECT 40.595 105.515 40.925 105.575 ;
        RECT 40.115 105.345 40.445 105.405 ;
        RECT 41.115 105.345 41.285 106.105 ;
        RECT 42.525 106.035 42.845 106.495 ;
        RECT 43.045 105.855 43.295 106.285 ;
        RECT 43.585 106.055 43.995 106.495 ;
        RECT 44.165 106.115 45.180 106.315 ;
        RECT 41.455 105.685 42.705 105.855 ;
        RECT 41.455 105.565 41.785 105.685 ;
        RECT 40.115 105.175 42.015 105.345 ;
        RECT 39.755 104.835 41.675 105.005 ;
        RECT 39.755 104.815 40.075 104.835 ;
        RECT 39.305 104.155 39.635 104.665 ;
        RECT 39.905 104.205 40.075 104.815 ;
        RECT 41.845 104.665 42.015 105.175 ;
        RECT 42.185 105.105 42.365 105.515 ;
        RECT 42.535 104.925 42.705 105.685 ;
        RECT 40.245 103.945 40.575 104.635 ;
        RECT 40.805 104.495 42.015 104.665 ;
        RECT 42.185 104.615 42.705 104.925 ;
        RECT 42.875 105.515 43.295 105.855 ;
        RECT 43.585 105.515 43.995 105.845 ;
        RECT 42.875 104.745 43.065 105.515 ;
        RECT 44.165 105.385 44.335 106.115 ;
        RECT 45.480 105.945 45.650 106.275 ;
        RECT 45.820 106.115 46.150 106.495 ;
        RECT 44.505 105.565 44.855 105.935 ;
        RECT 44.165 105.345 44.585 105.385 ;
        RECT 43.235 105.175 44.585 105.345 ;
        RECT 43.235 105.015 43.485 105.175 ;
        RECT 43.995 104.745 44.245 105.005 ;
        RECT 42.875 104.495 44.245 104.745 ;
        RECT 40.805 104.205 41.045 104.495 ;
        RECT 41.845 104.415 42.015 104.495 ;
        RECT 41.245 103.945 41.665 104.325 ;
        RECT 41.845 104.165 42.475 104.415 ;
        RECT 42.945 103.945 43.275 104.325 ;
        RECT 43.445 104.205 43.615 104.495 ;
        RECT 44.415 104.330 44.585 105.175 ;
        RECT 45.035 105.005 45.255 105.875 ;
        RECT 45.480 105.755 46.175 105.945 ;
        RECT 44.755 104.625 45.255 105.005 ;
        RECT 45.425 104.955 45.835 105.575 ;
        RECT 46.005 104.785 46.175 105.755 ;
        RECT 45.480 104.615 46.175 104.785 ;
        RECT 43.795 103.945 44.175 104.325 ;
        RECT 44.415 104.160 45.245 104.330 ;
        RECT 45.480 104.115 45.650 104.615 ;
        RECT 45.820 103.945 46.150 104.445 ;
        RECT 46.365 104.115 46.590 106.235 ;
        RECT 46.760 106.115 47.090 106.495 ;
        RECT 47.260 105.945 47.430 106.235 ;
        RECT 46.765 105.775 47.430 105.945 ;
        RECT 46.765 104.785 46.995 105.775 ;
        RECT 47.690 105.770 47.980 106.495 ;
        RECT 48.150 105.745 49.360 106.495 ;
        RECT 49.840 106.025 50.010 106.495 ;
        RECT 50.180 105.845 50.510 106.325 ;
        RECT 50.680 106.025 50.850 106.495 ;
        RECT 51.020 105.845 51.350 106.325 ;
        RECT 47.165 104.955 47.515 105.605 ;
        RECT 46.765 104.615 47.430 104.785 ;
        RECT 46.760 103.945 47.090 104.445 ;
        RECT 47.260 104.115 47.430 104.615 ;
        RECT 47.690 103.945 47.980 105.110 ;
        RECT 48.150 105.035 48.670 105.575 ;
        RECT 48.840 105.205 49.360 105.745 ;
        RECT 49.585 105.675 51.350 105.845 ;
        RECT 51.520 105.685 51.690 106.495 ;
        RECT 51.890 106.115 52.960 106.285 ;
        RECT 51.890 105.760 52.210 106.115 ;
        RECT 49.585 105.125 49.995 105.675 ;
        RECT 51.885 105.505 52.210 105.760 ;
        RECT 50.180 105.295 52.210 105.505 ;
        RECT 51.865 105.285 52.210 105.295 ;
        RECT 52.380 105.545 52.620 105.945 ;
        RECT 52.790 105.885 52.960 106.115 ;
        RECT 53.130 106.055 53.320 106.495 ;
        RECT 53.490 106.045 54.440 106.325 ;
        RECT 54.660 106.135 55.010 106.305 ;
        RECT 52.790 105.715 53.320 105.885 ;
        RECT 48.150 103.945 49.360 105.035 ;
        RECT 49.585 104.955 51.310 105.125 ;
        RECT 49.840 103.945 50.010 104.785 ;
        RECT 50.220 104.115 50.470 104.955 ;
        RECT 50.680 103.945 50.850 104.785 ;
        RECT 51.020 104.115 51.310 104.955 ;
        RECT 51.520 103.945 51.690 105.005 ;
        RECT 51.865 104.665 52.035 105.285 ;
        RECT 52.380 105.175 52.920 105.545 ;
        RECT 53.100 105.435 53.320 105.715 ;
        RECT 53.490 105.265 53.660 106.045 ;
        RECT 53.255 105.095 53.660 105.265 ;
        RECT 53.830 105.255 54.180 105.875 ;
        RECT 53.255 105.005 53.425 105.095 ;
        RECT 54.350 105.085 54.560 105.875 ;
        RECT 52.205 104.835 53.425 105.005 ;
        RECT 53.885 104.925 54.560 105.085 ;
        RECT 51.865 104.495 52.665 104.665 ;
        RECT 51.985 103.945 52.315 104.325 ;
        RECT 52.495 104.205 52.665 104.495 ;
        RECT 53.255 104.455 53.425 104.835 ;
        RECT 53.595 104.915 54.560 104.925 ;
        RECT 54.750 105.745 55.010 106.135 ;
        RECT 55.220 106.035 55.550 106.495 ;
        RECT 56.425 106.105 57.280 106.275 ;
        RECT 57.485 106.105 57.980 106.275 ;
        RECT 58.150 106.135 58.480 106.495 ;
        RECT 54.750 105.055 54.920 105.745 ;
        RECT 55.090 105.395 55.260 105.575 ;
        RECT 55.430 105.565 56.220 105.815 ;
        RECT 56.425 105.395 56.595 106.105 ;
        RECT 56.765 105.595 57.120 105.815 ;
        RECT 55.090 105.225 56.780 105.395 ;
        RECT 53.595 104.625 54.055 104.915 ;
        RECT 54.750 104.885 56.250 105.055 ;
        RECT 54.750 104.745 54.920 104.885 ;
        RECT 54.360 104.575 54.920 104.745 ;
        RECT 52.835 103.945 53.085 104.405 ;
        RECT 53.255 104.115 54.125 104.455 ;
        RECT 54.360 104.115 54.530 104.575 ;
        RECT 55.365 104.545 56.440 104.715 ;
        RECT 54.700 103.945 55.070 104.405 ;
        RECT 55.365 104.205 55.535 104.545 ;
        RECT 55.705 103.945 56.035 104.375 ;
        RECT 56.270 104.205 56.440 104.545 ;
        RECT 56.610 104.445 56.780 105.225 ;
        RECT 56.950 105.005 57.120 105.595 ;
        RECT 57.290 105.195 57.640 105.815 ;
        RECT 56.950 104.615 57.415 105.005 ;
        RECT 57.810 104.745 57.980 106.105 ;
        RECT 58.150 104.915 58.610 105.965 ;
        RECT 57.585 104.575 57.980 104.745 ;
        RECT 57.585 104.445 57.755 104.575 ;
        RECT 56.610 104.115 57.290 104.445 ;
        RECT 57.505 104.115 57.755 104.445 ;
        RECT 57.925 103.945 58.175 104.405 ;
        RECT 58.345 104.130 58.670 104.915 ;
        RECT 58.840 104.115 59.010 106.235 ;
        RECT 59.180 106.115 59.510 106.495 ;
        RECT 59.680 105.945 59.935 106.235 ;
        RECT 60.420 106.025 60.590 106.495 ;
        RECT 59.185 105.775 59.935 105.945 ;
        RECT 60.760 105.845 61.090 106.325 ;
        RECT 61.260 106.025 61.430 106.495 ;
        RECT 61.600 105.845 61.930 106.325 ;
        RECT 59.185 104.785 59.415 105.775 ;
        RECT 60.165 105.675 61.930 105.845 ;
        RECT 62.100 105.685 62.270 106.495 ;
        RECT 62.470 106.115 63.540 106.285 ;
        RECT 62.470 105.760 62.790 106.115 ;
        RECT 59.585 104.955 59.935 105.605 ;
        RECT 60.165 105.125 60.575 105.675 ;
        RECT 62.465 105.505 62.790 105.760 ;
        RECT 60.760 105.295 62.790 105.505 ;
        RECT 62.445 105.285 62.790 105.295 ;
        RECT 62.960 105.545 63.200 105.945 ;
        RECT 63.370 105.885 63.540 106.115 ;
        RECT 63.710 106.055 63.900 106.495 ;
        RECT 64.070 106.045 65.020 106.325 ;
        RECT 65.240 106.135 65.590 106.305 ;
        RECT 63.370 105.715 63.900 105.885 ;
        RECT 60.165 104.955 61.890 105.125 ;
        RECT 59.185 104.615 59.935 104.785 ;
        RECT 59.180 103.945 59.510 104.445 ;
        RECT 59.680 104.115 59.935 104.615 ;
        RECT 60.420 103.945 60.590 104.785 ;
        RECT 60.800 104.115 61.050 104.955 ;
        RECT 61.260 103.945 61.430 104.785 ;
        RECT 61.600 104.115 61.890 104.955 ;
        RECT 62.100 103.945 62.270 105.005 ;
        RECT 62.445 104.665 62.615 105.285 ;
        RECT 62.960 105.175 63.500 105.545 ;
        RECT 63.680 105.435 63.900 105.715 ;
        RECT 64.070 105.265 64.240 106.045 ;
        RECT 63.835 105.095 64.240 105.265 ;
        RECT 64.410 105.255 64.760 105.875 ;
        RECT 63.835 105.005 64.005 105.095 ;
        RECT 64.930 105.085 65.140 105.875 ;
        RECT 62.785 104.835 64.005 105.005 ;
        RECT 64.465 104.925 65.140 105.085 ;
        RECT 62.445 104.495 63.245 104.665 ;
        RECT 62.565 103.945 62.895 104.325 ;
        RECT 63.075 104.205 63.245 104.495 ;
        RECT 63.835 104.455 64.005 104.835 ;
        RECT 64.175 104.915 65.140 104.925 ;
        RECT 65.330 105.745 65.590 106.135 ;
        RECT 65.800 106.035 66.130 106.495 ;
        RECT 67.005 106.105 67.860 106.275 ;
        RECT 68.065 106.105 68.560 106.275 ;
        RECT 68.730 106.135 69.060 106.495 ;
        RECT 65.330 105.055 65.500 105.745 ;
        RECT 65.670 105.395 65.840 105.575 ;
        RECT 66.010 105.565 66.800 105.815 ;
        RECT 67.005 105.395 67.175 106.105 ;
        RECT 67.345 105.595 67.700 105.815 ;
        RECT 65.670 105.225 67.360 105.395 ;
        RECT 64.175 104.625 64.635 104.915 ;
        RECT 65.330 104.885 66.830 105.055 ;
        RECT 65.330 104.745 65.500 104.885 ;
        RECT 64.940 104.575 65.500 104.745 ;
        RECT 63.415 103.945 63.665 104.405 ;
        RECT 63.835 104.115 64.705 104.455 ;
        RECT 64.940 104.115 65.110 104.575 ;
        RECT 65.945 104.545 67.020 104.715 ;
        RECT 65.280 103.945 65.650 104.405 ;
        RECT 65.945 104.205 66.115 104.545 ;
        RECT 66.285 103.945 66.615 104.375 ;
        RECT 66.850 104.205 67.020 104.545 ;
        RECT 67.190 104.445 67.360 105.225 ;
        RECT 67.530 105.005 67.700 105.595 ;
        RECT 67.870 105.195 68.220 105.815 ;
        RECT 67.530 104.615 67.995 105.005 ;
        RECT 68.390 104.745 68.560 106.105 ;
        RECT 68.730 104.915 69.190 105.965 ;
        RECT 68.165 104.575 68.560 104.745 ;
        RECT 68.165 104.445 68.335 104.575 ;
        RECT 67.190 104.115 67.870 104.445 ;
        RECT 68.085 104.115 68.335 104.445 ;
        RECT 68.505 103.945 68.755 104.405 ;
        RECT 68.925 104.130 69.250 104.915 ;
        RECT 69.420 104.115 69.590 106.235 ;
        RECT 69.760 106.115 70.090 106.495 ;
        RECT 70.260 105.945 70.515 106.235 ;
        RECT 69.765 105.775 70.515 105.945 ;
        RECT 69.765 104.785 69.995 105.775 ;
        RECT 70.690 105.725 73.280 106.495 ;
        RECT 73.450 105.770 73.740 106.495 ;
        RECT 70.165 104.955 70.515 105.605 ;
        RECT 70.690 105.035 71.900 105.555 ;
        RECT 72.070 105.205 73.280 105.725 ;
        RECT 74.410 105.675 74.640 106.495 ;
        RECT 74.810 105.695 75.140 106.325 ;
        RECT 74.390 105.255 74.720 105.505 ;
        RECT 69.765 104.615 70.515 104.785 ;
        RECT 69.760 103.945 70.090 104.445 ;
        RECT 70.260 104.115 70.515 104.615 ;
        RECT 70.690 103.945 73.280 105.035 ;
        RECT 73.450 103.945 73.740 105.110 ;
        RECT 74.890 105.095 75.140 105.695 ;
        RECT 75.310 105.675 75.520 106.495 ;
        RECT 76.060 106.025 76.230 106.495 ;
        RECT 76.400 105.845 76.730 106.325 ;
        RECT 76.900 106.025 77.070 106.495 ;
        RECT 77.240 105.845 77.570 106.325 ;
        RECT 75.805 105.675 77.570 105.845 ;
        RECT 77.740 105.685 77.910 106.495 ;
        RECT 78.110 106.115 79.180 106.285 ;
        RECT 78.110 105.760 78.430 106.115 ;
        RECT 74.410 103.945 74.640 105.085 ;
        RECT 74.810 104.115 75.140 105.095 ;
        RECT 75.805 105.125 76.215 105.675 ;
        RECT 78.105 105.505 78.430 105.760 ;
        RECT 76.400 105.295 78.430 105.505 ;
        RECT 78.085 105.285 78.430 105.295 ;
        RECT 78.600 105.545 78.840 105.945 ;
        RECT 79.010 105.885 79.180 106.115 ;
        RECT 79.350 106.055 79.540 106.495 ;
        RECT 79.710 106.045 80.660 106.325 ;
        RECT 80.880 106.135 81.230 106.305 ;
        RECT 79.010 105.715 79.540 105.885 ;
        RECT 75.310 103.945 75.520 105.085 ;
        RECT 75.805 104.955 77.530 105.125 ;
        RECT 76.060 103.945 76.230 104.785 ;
        RECT 76.440 104.115 76.690 104.955 ;
        RECT 76.900 103.945 77.070 104.785 ;
        RECT 77.240 104.115 77.530 104.955 ;
        RECT 77.740 103.945 77.910 105.005 ;
        RECT 78.085 104.665 78.255 105.285 ;
        RECT 78.600 105.175 79.140 105.545 ;
        RECT 79.320 105.435 79.540 105.715 ;
        RECT 79.710 105.265 79.880 106.045 ;
        RECT 79.475 105.095 79.880 105.265 ;
        RECT 80.050 105.255 80.400 105.875 ;
        RECT 79.475 105.005 79.645 105.095 ;
        RECT 80.570 105.085 80.780 105.875 ;
        RECT 78.425 104.835 79.645 105.005 ;
        RECT 80.105 104.925 80.780 105.085 ;
        RECT 78.085 104.495 78.885 104.665 ;
        RECT 78.205 103.945 78.535 104.325 ;
        RECT 78.715 104.205 78.885 104.495 ;
        RECT 79.475 104.455 79.645 104.835 ;
        RECT 79.815 104.915 80.780 104.925 ;
        RECT 80.970 105.745 81.230 106.135 ;
        RECT 81.440 106.035 81.770 106.495 ;
        RECT 82.645 106.105 83.500 106.275 ;
        RECT 83.705 106.105 84.200 106.275 ;
        RECT 84.370 106.135 84.700 106.495 ;
        RECT 80.970 105.055 81.140 105.745 ;
        RECT 81.310 105.395 81.480 105.575 ;
        RECT 81.650 105.565 82.440 105.815 ;
        RECT 82.645 105.395 82.815 106.105 ;
        RECT 82.985 105.595 83.340 105.815 ;
        RECT 81.310 105.225 83.000 105.395 ;
        RECT 79.815 104.625 80.275 104.915 ;
        RECT 80.970 104.885 82.470 105.055 ;
        RECT 80.970 104.745 81.140 104.885 ;
        RECT 80.580 104.575 81.140 104.745 ;
        RECT 79.055 103.945 79.305 104.405 ;
        RECT 79.475 104.115 80.345 104.455 ;
        RECT 80.580 104.115 80.750 104.575 ;
        RECT 81.585 104.545 82.660 104.715 ;
        RECT 80.920 103.945 81.290 104.405 ;
        RECT 81.585 104.205 81.755 104.545 ;
        RECT 81.925 103.945 82.255 104.375 ;
        RECT 82.490 104.205 82.660 104.545 ;
        RECT 82.830 104.445 83.000 105.225 ;
        RECT 83.170 105.005 83.340 105.595 ;
        RECT 83.510 105.195 83.860 105.815 ;
        RECT 83.170 104.615 83.635 105.005 ;
        RECT 84.030 104.745 84.200 106.105 ;
        RECT 84.370 104.915 84.830 105.965 ;
        RECT 83.805 104.575 84.200 104.745 ;
        RECT 83.805 104.445 83.975 104.575 ;
        RECT 82.830 104.115 83.510 104.445 ;
        RECT 83.725 104.115 83.975 104.445 ;
        RECT 84.145 103.945 84.395 104.405 ;
        RECT 84.565 104.130 84.890 104.915 ;
        RECT 85.060 104.115 85.230 106.235 ;
        RECT 85.400 106.115 85.730 106.495 ;
        RECT 85.900 105.945 86.155 106.235 ;
        RECT 86.640 106.025 86.810 106.495 ;
        RECT 85.405 105.775 86.155 105.945 ;
        RECT 86.980 105.845 87.310 106.325 ;
        RECT 87.480 106.025 87.650 106.495 ;
        RECT 87.820 105.845 88.150 106.325 ;
        RECT 85.405 104.785 85.635 105.775 ;
        RECT 86.385 105.675 88.150 105.845 ;
        RECT 88.320 105.685 88.490 106.495 ;
        RECT 88.690 106.115 89.760 106.285 ;
        RECT 88.690 105.760 89.010 106.115 ;
        RECT 85.805 104.955 86.155 105.605 ;
        RECT 86.385 105.125 86.795 105.675 ;
        RECT 88.685 105.505 89.010 105.760 ;
        RECT 86.980 105.295 89.010 105.505 ;
        RECT 88.665 105.285 89.010 105.295 ;
        RECT 89.180 105.545 89.420 105.945 ;
        RECT 89.590 105.885 89.760 106.115 ;
        RECT 89.930 106.055 90.120 106.495 ;
        RECT 90.290 106.045 91.240 106.325 ;
        RECT 91.460 106.135 91.810 106.305 ;
        RECT 89.590 105.715 90.120 105.885 ;
        RECT 86.385 104.955 88.110 105.125 ;
        RECT 85.405 104.615 86.155 104.785 ;
        RECT 85.400 103.945 85.730 104.445 ;
        RECT 85.900 104.115 86.155 104.615 ;
        RECT 86.640 103.945 86.810 104.785 ;
        RECT 87.020 104.115 87.270 104.955 ;
        RECT 87.480 103.945 87.650 104.785 ;
        RECT 87.820 104.115 88.110 104.955 ;
        RECT 88.320 103.945 88.490 105.005 ;
        RECT 88.665 104.665 88.835 105.285 ;
        RECT 89.180 105.175 89.720 105.545 ;
        RECT 89.900 105.435 90.120 105.715 ;
        RECT 90.290 105.265 90.460 106.045 ;
        RECT 90.055 105.095 90.460 105.265 ;
        RECT 90.630 105.255 90.980 105.875 ;
        RECT 90.055 105.005 90.225 105.095 ;
        RECT 91.150 105.085 91.360 105.875 ;
        RECT 89.005 104.835 90.225 105.005 ;
        RECT 90.685 104.925 91.360 105.085 ;
        RECT 88.665 104.495 89.465 104.665 ;
        RECT 88.785 103.945 89.115 104.325 ;
        RECT 89.295 104.205 89.465 104.495 ;
        RECT 90.055 104.455 90.225 104.835 ;
        RECT 90.395 104.915 91.360 104.925 ;
        RECT 91.550 105.745 91.810 106.135 ;
        RECT 92.020 106.035 92.350 106.495 ;
        RECT 93.225 106.105 94.080 106.275 ;
        RECT 94.285 106.105 94.780 106.275 ;
        RECT 94.950 106.135 95.280 106.495 ;
        RECT 91.550 105.055 91.720 105.745 ;
        RECT 91.890 105.395 92.060 105.575 ;
        RECT 92.230 105.565 93.020 105.815 ;
        RECT 93.225 105.395 93.395 106.105 ;
        RECT 93.565 105.595 93.920 105.815 ;
        RECT 91.890 105.225 93.580 105.395 ;
        RECT 90.395 104.625 90.855 104.915 ;
        RECT 91.550 104.885 93.050 105.055 ;
        RECT 91.550 104.745 91.720 104.885 ;
        RECT 91.160 104.575 91.720 104.745 ;
        RECT 89.635 103.945 89.885 104.405 ;
        RECT 90.055 104.115 90.925 104.455 ;
        RECT 91.160 104.115 91.330 104.575 ;
        RECT 92.165 104.545 93.240 104.715 ;
        RECT 91.500 103.945 91.870 104.405 ;
        RECT 92.165 104.205 92.335 104.545 ;
        RECT 92.505 103.945 92.835 104.375 ;
        RECT 93.070 104.205 93.240 104.545 ;
        RECT 93.410 104.445 93.580 105.225 ;
        RECT 93.750 105.005 93.920 105.595 ;
        RECT 94.090 105.195 94.440 105.815 ;
        RECT 93.750 104.615 94.215 105.005 ;
        RECT 94.610 104.745 94.780 106.105 ;
        RECT 94.950 104.915 95.410 105.965 ;
        RECT 94.385 104.575 94.780 104.745 ;
        RECT 94.385 104.445 94.555 104.575 ;
        RECT 93.410 104.115 94.090 104.445 ;
        RECT 94.305 104.115 94.555 104.445 ;
        RECT 94.725 103.945 94.975 104.405 ;
        RECT 95.145 104.130 95.470 104.915 ;
        RECT 95.640 104.115 95.810 106.235 ;
        RECT 95.980 106.115 96.310 106.495 ;
        RECT 96.480 105.945 96.735 106.235 ;
        RECT 95.985 105.775 96.735 105.945 ;
        RECT 95.985 104.785 96.215 105.775 ;
        RECT 97.370 105.725 99.040 106.495 ;
        RECT 99.210 105.770 99.500 106.495 ;
        RECT 100.135 105.950 105.480 106.495 ;
        RECT 105.655 105.950 111.000 106.495 ;
        RECT 96.385 104.955 96.735 105.605 ;
        RECT 97.370 105.035 98.120 105.555 ;
        RECT 98.290 105.205 99.040 105.725 ;
        RECT 95.985 104.615 96.735 104.785 ;
        RECT 95.980 103.945 96.310 104.445 ;
        RECT 96.480 104.115 96.735 104.615 ;
        RECT 97.370 103.945 99.040 105.035 ;
        RECT 99.210 103.945 99.500 105.110 ;
        RECT 101.725 104.380 102.075 105.630 ;
        RECT 103.555 105.120 103.895 105.950 ;
        RECT 107.245 104.380 107.595 105.630 ;
        RECT 109.075 105.120 109.415 105.950 ;
        RECT 111.170 105.745 112.380 106.495 ;
        RECT 111.170 105.035 111.690 105.575 ;
        RECT 111.860 105.205 112.380 105.745 ;
        RECT 100.135 103.945 105.480 104.380 ;
        RECT 105.655 103.945 111.000 104.380 ;
        RECT 111.170 103.945 112.380 105.035 ;
        RECT 18.165 103.775 112.465 103.945 ;
        RECT 18.250 102.685 19.460 103.775 ;
        RECT 18.250 101.975 18.770 102.515 ;
        RECT 18.940 102.145 19.460 102.685 ;
        RECT 20.090 102.685 21.760 103.775 ;
        RECT 20.090 102.165 20.840 102.685 ;
        RECT 21.930 102.610 22.220 103.775 ;
        RECT 22.390 102.685 23.600 103.775 ;
        RECT 23.775 103.340 29.120 103.775 ;
        RECT 29.295 103.340 34.640 103.775 ;
        RECT 21.010 101.995 21.760 102.515 ;
        RECT 22.390 102.145 22.910 102.685 ;
        RECT 18.250 101.225 19.460 101.975 ;
        RECT 20.090 101.225 21.760 101.995 ;
        RECT 23.080 101.975 23.600 102.515 ;
        RECT 25.365 102.090 25.715 103.340 ;
        RECT 21.930 101.225 22.220 101.950 ;
        RECT 22.390 101.225 23.600 101.975 ;
        RECT 27.195 101.770 27.535 102.600 ;
        RECT 30.885 102.090 31.235 103.340 ;
        RECT 34.810 102.610 35.100 103.775 ;
        RECT 35.270 102.685 36.480 103.775 ;
        RECT 36.655 103.340 42.000 103.775 ;
        RECT 42.175 103.340 47.520 103.775 ;
        RECT 32.715 101.770 33.055 102.600 ;
        RECT 35.270 102.145 35.790 102.685 ;
        RECT 35.960 101.975 36.480 102.515 ;
        RECT 38.245 102.090 38.595 103.340 ;
        RECT 23.775 101.225 29.120 101.770 ;
        RECT 29.295 101.225 34.640 101.770 ;
        RECT 34.810 101.225 35.100 101.950 ;
        RECT 35.270 101.225 36.480 101.975 ;
        RECT 40.075 101.770 40.415 102.600 ;
        RECT 43.765 102.090 44.115 103.340 ;
        RECT 47.690 102.610 47.980 103.775 ;
        RECT 48.155 103.340 53.500 103.775 ;
        RECT 45.595 101.770 45.935 102.600 ;
        RECT 49.745 102.090 50.095 103.340 ;
        RECT 53.730 102.635 53.940 103.775 ;
        RECT 54.110 102.625 54.440 103.605 ;
        RECT 54.610 102.635 54.840 103.775 ;
        RECT 55.055 103.340 60.400 103.775 ;
        RECT 36.655 101.225 42.000 101.770 ;
        RECT 42.175 101.225 47.520 101.770 ;
        RECT 47.690 101.225 47.980 101.950 ;
        RECT 51.575 101.770 51.915 102.600 ;
        RECT 48.155 101.225 53.500 101.770 ;
        RECT 53.730 101.225 53.940 102.045 ;
        RECT 54.110 102.025 54.360 102.625 ;
        RECT 54.530 102.215 54.860 102.465 ;
        RECT 56.645 102.090 56.995 103.340 ;
        RECT 60.570 102.610 60.860 103.775 ;
        RECT 61.030 102.685 62.240 103.775 ;
        RECT 54.110 101.395 54.440 102.025 ;
        RECT 54.610 101.225 54.840 102.045 ;
        RECT 58.475 101.770 58.815 102.600 ;
        RECT 61.030 102.145 61.550 102.685 ;
        RECT 62.450 102.635 62.680 103.775 ;
        RECT 62.850 102.625 63.180 103.605 ;
        RECT 63.350 102.635 63.560 103.775 ;
        RECT 64.250 102.685 67.760 103.775 ;
        RECT 67.935 103.340 73.280 103.775 ;
        RECT 61.720 101.975 62.240 102.515 ;
        RECT 62.430 102.215 62.760 102.465 ;
        RECT 55.055 101.225 60.400 101.770 ;
        RECT 60.570 101.225 60.860 101.950 ;
        RECT 61.030 101.225 62.240 101.975 ;
        RECT 62.450 101.225 62.680 102.045 ;
        RECT 62.930 102.025 63.180 102.625 ;
        RECT 64.250 102.165 65.940 102.685 ;
        RECT 62.850 101.395 63.180 102.025 ;
        RECT 63.350 101.225 63.560 102.045 ;
        RECT 66.110 101.995 67.760 102.515 ;
        RECT 69.525 102.090 69.875 103.340 ;
        RECT 73.450 102.610 73.740 103.775 ;
        RECT 74.375 103.340 79.720 103.775 ;
        RECT 64.250 101.225 67.760 101.995 ;
        RECT 71.355 101.770 71.695 102.600 ;
        RECT 75.965 102.090 76.315 103.340 ;
        RECT 79.950 102.635 80.160 103.775 ;
        RECT 80.330 102.625 80.660 103.605 ;
        RECT 80.830 102.635 81.060 103.775 ;
        RECT 81.270 102.685 82.480 103.775 ;
        RECT 82.650 102.685 86.160 103.775 ;
        RECT 67.935 101.225 73.280 101.770 ;
        RECT 73.450 101.225 73.740 101.950 ;
        RECT 77.795 101.770 78.135 102.600 ;
        RECT 74.375 101.225 79.720 101.770 ;
        RECT 79.950 101.225 80.160 102.045 ;
        RECT 80.330 102.025 80.580 102.625 ;
        RECT 80.750 102.215 81.080 102.465 ;
        RECT 81.270 102.145 81.790 102.685 ;
        RECT 80.330 101.395 80.660 102.025 ;
        RECT 80.830 101.225 81.060 102.045 ;
        RECT 81.960 101.975 82.480 102.515 ;
        RECT 82.650 102.165 84.340 102.685 ;
        RECT 86.330 102.610 86.620 103.775 ;
        RECT 86.790 102.685 88.000 103.775 ;
        RECT 88.175 103.340 93.520 103.775 ;
        RECT 93.695 103.340 99.040 103.775 ;
        RECT 84.510 101.995 86.160 102.515 ;
        RECT 86.790 102.145 87.310 102.685 ;
        RECT 81.270 101.225 82.480 101.975 ;
        RECT 82.650 101.225 86.160 101.995 ;
        RECT 87.480 101.975 88.000 102.515 ;
        RECT 89.765 102.090 90.115 103.340 ;
        RECT 86.330 101.225 86.620 101.950 ;
        RECT 86.790 101.225 88.000 101.975 ;
        RECT 91.595 101.770 91.935 102.600 ;
        RECT 95.285 102.090 95.635 103.340 ;
        RECT 99.210 102.610 99.500 103.775 ;
        RECT 100.135 103.340 105.480 103.775 ;
        RECT 105.655 103.340 111.000 103.775 ;
        RECT 97.115 101.770 97.455 102.600 ;
        RECT 101.725 102.090 102.075 103.340 ;
        RECT 88.175 101.225 93.520 101.770 ;
        RECT 93.695 101.225 99.040 101.770 ;
        RECT 99.210 101.225 99.500 101.950 ;
        RECT 103.555 101.770 103.895 102.600 ;
        RECT 107.245 102.090 107.595 103.340 ;
        RECT 111.170 102.685 112.380 103.775 ;
        RECT 109.075 101.770 109.415 102.600 ;
        RECT 111.170 102.145 111.690 102.685 ;
        RECT 111.860 101.975 112.380 102.515 ;
        RECT 100.135 101.225 105.480 101.770 ;
        RECT 105.655 101.225 111.000 101.770 ;
        RECT 111.170 101.225 112.380 101.975 ;
        RECT 18.165 101.055 112.465 101.225 ;
        RECT 19.165 66.070 30.165 66.940 ;
        RECT 19.165 54.930 20.835 66.070 ;
        RECT 21.465 65.555 26.465 65.725 ;
        RECT 21.235 55.300 21.405 65.340 ;
        RECT 26.525 55.300 26.695 65.340 ;
        RECT 27.095 54.930 27.265 66.070 ;
        RECT 27.895 65.555 28.895 65.725 ;
        RECT 27.665 55.300 27.835 65.340 ;
        RECT 28.955 55.300 29.125 65.340 ;
        RECT 29.525 54.930 30.165 66.070 ;
        RECT 19.165 52.860 30.165 54.930 ;
        RECT 19.165 49.370 21.005 52.860 ;
        RECT 22.765 52.780 30.165 52.860 ;
        RECT 21.635 52.350 22.135 52.520 ;
        RECT 21.405 50.095 21.575 52.135 ;
        RECT 22.195 50.095 22.365 52.135 ;
        RECT 21.635 49.710 22.135 49.880 ;
        RECT 22.765 49.370 25.085 52.780 ;
        RECT 25.715 52.270 26.215 52.440 ;
        RECT 19.165 48.650 25.085 49.370 ;
        RECT 19.135 48.040 23.045 48.260 ;
        RECT 19.135 45.640 20.855 48.040 ;
        RECT 21.485 47.530 21.985 47.700 ;
        RECT 21.255 46.320 21.425 47.360 ;
        RECT 22.045 46.320 22.215 47.360 ;
        RECT 21.485 45.980 21.985 46.150 ;
        RECT 22.615 45.640 23.045 48.040 ;
        RECT 24.025 46.290 25.085 48.650 ;
        RECT 25.485 47.015 25.655 52.055 ;
        RECT 26.275 47.015 26.445 52.055 ;
        RECT 25.715 46.630 26.215 46.800 ;
        RECT 26.845 46.290 27.015 52.780 ;
        RECT 27.645 52.270 28.145 52.440 ;
        RECT 27.415 47.015 27.585 52.055 ;
        RECT 28.205 47.015 28.375 52.055 ;
        RECT 27.645 46.630 28.145 46.800 ;
        RECT 28.775 46.290 30.165 52.780 ;
        RECT 30.365 66.080 41.365 66.950 ;
        RECT 30.365 54.940 32.035 66.080 ;
        RECT 32.665 65.565 37.665 65.735 ;
        RECT 32.435 55.310 32.605 65.350 ;
        RECT 37.725 55.310 37.895 65.350 ;
        RECT 38.295 54.940 38.465 66.080 ;
        RECT 39.095 65.565 40.095 65.735 ;
        RECT 38.865 55.310 39.035 65.350 ;
        RECT 40.155 55.310 40.325 65.350 ;
        RECT 40.725 54.940 41.365 66.080 ;
        RECT 30.365 52.870 41.365 54.940 ;
        RECT 30.365 49.380 32.205 52.870 ;
        RECT 33.965 52.790 41.365 52.870 ;
        RECT 32.835 52.360 33.335 52.530 ;
        RECT 32.605 50.105 32.775 52.145 ;
        RECT 33.395 50.105 33.565 52.145 ;
        RECT 32.835 49.720 33.335 49.890 ;
        RECT 33.965 49.380 36.285 52.790 ;
        RECT 36.915 52.280 37.415 52.450 ;
        RECT 30.365 48.660 36.285 49.380 ;
        RECT 24.025 45.800 30.165 46.290 ;
        RECT 30.335 48.050 34.245 48.270 ;
        RECT 19.135 45.370 23.045 45.640 ;
        RECT 30.335 45.650 32.055 48.050 ;
        RECT 32.685 47.540 33.185 47.710 ;
        RECT 32.455 46.330 32.625 47.370 ;
        RECT 33.245 46.330 33.415 47.370 ;
        RECT 32.685 45.990 33.185 46.160 ;
        RECT 33.815 45.650 34.245 48.050 ;
        RECT 35.225 46.300 36.285 48.660 ;
        RECT 36.685 47.025 36.855 52.065 ;
        RECT 37.475 47.025 37.645 52.065 ;
        RECT 36.915 46.640 37.415 46.810 ;
        RECT 38.045 46.300 38.215 52.790 ;
        RECT 38.845 52.280 39.345 52.450 ;
        RECT 38.615 47.025 38.785 52.065 ;
        RECT 39.405 47.025 39.575 52.065 ;
        RECT 38.845 46.640 39.345 46.810 ;
        RECT 39.975 46.300 41.365 52.790 ;
        RECT 41.585 66.050 52.585 66.920 ;
        RECT 41.585 54.910 43.255 66.050 ;
        RECT 43.885 65.535 48.885 65.705 ;
        RECT 43.655 55.280 43.825 65.320 ;
        RECT 48.945 55.280 49.115 65.320 ;
        RECT 49.515 54.910 49.685 66.050 ;
        RECT 50.315 65.535 51.315 65.705 ;
        RECT 50.085 55.280 50.255 65.320 ;
        RECT 51.375 55.280 51.545 65.320 ;
        RECT 51.945 54.910 52.585 66.050 ;
        RECT 41.585 52.840 52.585 54.910 ;
        RECT 41.585 49.350 43.425 52.840 ;
        RECT 45.185 52.760 52.585 52.840 ;
        RECT 44.055 52.330 44.555 52.500 ;
        RECT 43.825 50.075 43.995 52.115 ;
        RECT 44.615 50.075 44.785 52.115 ;
        RECT 44.055 49.690 44.555 49.860 ;
        RECT 45.185 49.350 47.505 52.760 ;
        RECT 48.135 52.250 48.635 52.420 ;
        RECT 41.585 48.630 47.505 49.350 ;
        RECT 35.225 45.810 41.365 46.300 ;
        RECT 41.555 48.020 45.465 48.240 ;
        RECT 30.335 45.380 34.245 45.650 ;
        RECT 41.555 45.620 43.275 48.020 ;
        RECT 43.905 47.510 44.405 47.680 ;
        RECT 43.675 46.300 43.845 47.340 ;
        RECT 44.465 46.300 44.635 47.340 ;
        RECT 43.905 45.960 44.405 46.130 ;
        RECT 45.035 45.620 45.465 48.020 ;
        RECT 46.445 46.270 47.505 48.630 ;
        RECT 47.905 46.995 48.075 52.035 ;
        RECT 48.695 46.995 48.865 52.035 ;
        RECT 48.135 46.610 48.635 46.780 ;
        RECT 49.265 46.270 49.435 52.760 ;
        RECT 50.065 52.250 50.565 52.420 ;
        RECT 49.835 46.995 50.005 52.035 ;
        RECT 50.625 46.995 50.795 52.035 ;
        RECT 50.065 46.610 50.565 46.780 ;
        RECT 51.195 46.270 52.585 52.760 ;
        RECT 52.835 66.030 63.835 66.900 ;
        RECT 52.835 54.890 54.505 66.030 ;
        RECT 55.135 65.515 60.135 65.685 ;
        RECT 54.905 55.260 55.075 65.300 ;
        RECT 60.195 55.260 60.365 65.300 ;
        RECT 60.765 54.890 60.935 66.030 ;
        RECT 61.565 65.515 62.565 65.685 ;
        RECT 61.335 55.260 61.505 65.300 ;
        RECT 62.625 55.260 62.795 65.300 ;
        RECT 63.195 54.890 63.835 66.030 ;
        RECT 52.835 52.820 63.835 54.890 ;
        RECT 52.835 49.330 54.675 52.820 ;
        RECT 56.435 52.740 63.835 52.820 ;
        RECT 55.305 52.310 55.805 52.480 ;
        RECT 55.075 50.055 55.245 52.095 ;
        RECT 55.865 50.055 56.035 52.095 ;
        RECT 55.305 49.670 55.805 49.840 ;
        RECT 56.435 49.330 58.755 52.740 ;
        RECT 59.385 52.230 59.885 52.400 ;
        RECT 52.835 48.610 58.755 49.330 ;
        RECT 46.445 45.780 52.585 46.270 ;
        RECT 52.805 48.000 56.715 48.220 ;
        RECT 41.555 45.350 45.465 45.620 ;
        RECT 52.805 45.600 54.525 48.000 ;
        RECT 55.155 47.490 55.655 47.660 ;
        RECT 54.925 46.280 55.095 47.320 ;
        RECT 55.715 46.280 55.885 47.320 ;
        RECT 55.155 45.940 55.655 46.110 ;
        RECT 56.285 45.600 56.715 48.000 ;
        RECT 57.695 46.250 58.755 48.610 ;
        RECT 59.155 46.975 59.325 52.015 ;
        RECT 59.945 46.975 60.115 52.015 ;
        RECT 59.385 46.590 59.885 46.760 ;
        RECT 60.515 46.250 60.685 52.740 ;
        RECT 61.315 52.230 61.815 52.400 ;
        RECT 61.085 46.975 61.255 52.015 ;
        RECT 61.875 46.975 62.045 52.015 ;
        RECT 61.315 46.590 61.815 46.760 ;
        RECT 62.445 46.250 63.835 52.740 ;
        RECT 64.055 66.020 75.055 66.890 ;
        RECT 64.055 54.880 65.725 66.020 ;
        RECT 66.355 65.505 71.355 65.675 ;
        RECT 66.125 55.250 66.295 65.290 ;
        RECT 71.415 55.250 71.585 65.290 ;
        RECT 71.985 54.880 72.155 66.020 ;
        RECT 72.785 65.505 73.785 65.675 ;
        RECT 72.555 55.250 72.725 65.290 ;
        RECT 73.845 55.250 74.015 65.290 ;
        RECT 74.415 54.880 75.055 66.020 ;
        RECT 64.055 52.810 75.055 54.880 ;
        RECT 64.055 49.320 65.895 52.810 ;
        RECT 67.655 52.730 75.055 52.810 ;
        RECT 66.525 52.300 67.025 52.470 ;
        RECT 66.295 50.045 66.465 52.085 ;
        RECT 67.085 50.045 67.255 52.085 ;
        RECT 66.525 49.660 67.025 49.830 ;
        RECT 67.655 49.320 69.975 52.730 ;
        RECT 70.605 52.220 71.105 52.390 ;
        RECT 64.055 48.600 69.975 49.320 ;
        RECT 57.695 45.760 63.835 46.250 ;
        RECT 64.025 47.990 67.935 48.210 ;
        RECT 52.805 45.330 56.715 45.600 ;
        RECT 64.025 45.590 65.745 47.990 ;
        RECT 66.375 47.480 66.875 47.650 ;
        RECT 66.145 46.270 66.315 47.310 ;
        RECT 66.935 46.270 67.105 47.310 ;
        RECT 66.375 45.930 66.875 46.100 ;
        RECT 67.505 45.590 67.935 47.990 ;
        RECT 68.915 46.240 69.975 48.600 ;
        RECT 70.375 46.965 70.545 52.005 ;
        RECT 71.165 46.965 71.335 52.005 ;
        RECT 70.605 46.580 71.105 46.750 ;
        RECT 71.735 46.240 71.905 52.730 ;
        RECT 72.535 52.220 73.035 52.390 ;
        RECT 72.305 46.965 72.475 52.005 ;
        RECT 73.095 46.965 73.265 52.005 ;
        RECT 72.535 46.580 73.035 46.750 ;
        RECT 73.665 46.240 75.055 52.730 ;
        RECT 75.295 66.010 86.295 66.880 ;
        RECT 75.295 54.870 76.965 66.010 ;
        RECT 77.595 65.495 82.595 65.665 ;
        RECT 77.365 55.240 77.535 65.280 ;
        RECT 82.655 55.240 82.825 65.280 ;
        RECT 83.225 54.870 83.395 66.010 ;
        RECT 84.025 65.495 85.025 65.665 ;
        RECT 83.795 55.240 83.965 65.280 ;
        RECT 85.085 55.240 85.255 65.280 ;
        RECT 85.655 54.870 86.295 66.010 ;
        RECT 75.295 52.800 86.295 54.870 ;
        RECT 75.295 49.310 77.135 52.800 ;
        RECT 78.895 52.720 86.295 52.800 ;
        RECT 77.765 52.290 78.265 52.460 ;
        RECT 77.535 50.035 77.705 52.075 ;
        RECT 78.325 50.035 78.495 52.075 ;
        RECT 77.765 49.650 78.265 49.820 ;
        RECT 78.895 49.310 81.215 52.720 ;
        RECT 81.845 52.210 82.345 52.380 ;
        RECT 75.295 48.590 81.215 49.310 ;
        RECT 68.915 45.750 75.055 46.240 ;
        RECT 75.265 47.980 79.175 48.200 ;
        RECT 64.025 45.320 67.935 45.590 ;
        RECT 75.265 45.580 76.985 47.980 ;
        RECT 77.615 47.470 78.115 47.640 ;
        RECT 77.385 46.260 77.555 47.300 ;
        RECT 78.175 46.260 78.345 47.300 ;
        RECT 77.615 45.920 78.115 46.090 ;
        RECT 78.745 45.580 79.175 47.980 ;
        RECT 80.155 46.230 81.215 48.590 ;
        RECT 81.615 46.955 81.785 51.995 ;
        RECT 82.405 46.955 82.575 51.995 ;
        RECT 81.845 46.570 82.345 46.740 ;
        RECT 82.975 46.230 83.145 52.720 ;
        RECT 83.775 52.210 84.275 52.380 ;
        RECT 83.545 46.955 83.715 51.995 ;
        RECT 84.335 46.955 84.505 51.995 ;
        RECT 83.775 46.570 84.275 46.740 ;
        RECT 84.905 46.230 86.295 52.720 ;
        RECT 86.545 66.020 97.545 66.890 ;
        RECT 131.125 66.880 140.025 66.890 ;
        RECT 86.545 54.880 88.215 66.020 ;
        RECT 88.845 65.505 93.845 65.675 ;
        RECT 88.615 55.250 88.785 65.290 ;
        RECT 93.905 55.250 94.075 65.290 ;
        RECT 94.475 54.880 94.645 66.020 ;
        RECT 95.275 65.505 96.275 65.675 ;
        RECT 95.045 55.250 95.215 65.290 ;
        RECT 96.335 55.250 96.505 65.290 ;
        RECT 96.905 54.880 97.545 66.020 ;
        RECT 86.545 52.810 97.545 54.880 ;
        RECT 86.545 49.320 88.385 52.810 ;
        RECT 90.145 52.730 97.545 52.810 ;
        RECT 89.015 52.300 89.515 52.470 ;
        RECT 88.785 50.045 88.955 52.085 ;
        RECT 89.575 50.045 89.745 52.085 ;
        RECT 89.015 49.660 89.515 49.830 ;
        RECT 90.145 49.320 92.465 52.730 ;
        RECT 93.095 52.220 93.595 52.390 ;
        RECT 86.545 48.600 92.465 49.320 ;
        RECT 80.155 45.740 86.295 46.230 ;
        RECT 86.515 47.990 90.425 48.210 ;
        RECT 75.265 45.310 79.175 45.580 ;
        RECT 86.515 45.590 88.235 47.990 ;
        RECT 88.865 47.480 89.365 47.650 ;
        RECT 88.635 46.270 88.805 47.310 ;
        RECT 89.425 46.270 89.595 47.310 ;
        RECT 88.865 45.930 89.365 46.100 ;
        RECT 89.995 45.590 90.425 47.990 ;
        RECT 91.405 46.240 92.465 48.600 ;
        RECT 92.865 46.965 93.035 52.005 ;
        RECT 93.655 46.965 93.825 52.005 ;
        RECT 93.095 46.580 93.595 46.750 ;
        RECT 94.225 46.240 94.395 52.730 ;
        RECT 95.025 52.220 95.525 52.390 ;
        RECT 94.795 46.965 94.965 52.005 ;
        RECT 95.585 46.965 95.755 52.005 ;
        RECT 95.025 46.580 95.525 46.750 ;
        RECT 96.155 46.240 97.545 52.730 ;
        RECT 97.825 66.010 108.825 66.880 ;
        RECT 97.825 54.870 99.495 66.010 ;
        RECT 100.125 65.495 105.125 65.665 ;
        RECT 99.895 55.240 100.065 65.280 ;
        RECT 105.185 55.240 105.355 65.280 ;
        RECT 105.755 54.870 105.925 66.010 ;
        RECT 106.555 65.495 107.555 65.665 ;
        RECT 106.325 55.240 106.495 65.280 ;
        RECT 107.615 55.240 107.785 65.280 ;
        RECT 108.185 54.870 108.825 66.010 ;
        RECT 97.825 52.800 108.825 54.870 ;
        RECT 97.825 49.310 99.665 52.800 ;
        RECT 101.425 52.720 108.825 52.800 ;
        RECT 100.295 52.290 100.795 52.460 ;
        RECT 100.065 50.035 100.235 52.075 ;
        RECT 100.855 50.035 101.025 52.075 ;
        RECT 100.295 49.650 100.795 49.820 ;
        RECT 101.425 49.310 103.745 52.720 ;
        RECT 104.375 52.210 104.875 52.380 ;
        RECT 97.825 48.590 103.745 49.310 ;
        RECT 91.405 45.750 97.545 46.240 ;
        RECT 97.795 47.980 101.705 48.200 ;
        RECT 86.515 45.320 90.425 45.590 ;
        RECT 97.795 45.580 99.515 47.980 ;
        RECT 100.145 47.470 100.645 47.640 ;
        RECT 99.915 46.260 100.085 47.300 ;
        RECT 100.705 46.260 100.875 47.300 ;
        RECT 100.145 45.920 100.645 46.090 ;
        RECT 101.275 45.580 101.705 47.980 ;
        RECT 102.685 46.230 103.745 48.590 ;
        RECT 104.145 46.955 104.315 51.995 ;
        RECT 104.935 46.955 105.105 51.995 ;
        RECT 104.375 46.570 104.875 46.740 ;
        RECT 105.505 46.230 105.675 52.720 ;
        RECT 106.305 52.210 106.805 52.380 ;
        RECT 106.075 46.955 106.245 51.995 ;
        RECT 106.865 46.955 107.035 51.995 ;
        RECT 106.305 46.570 106.805 46.740 ;
        RECT 107.435 46.230 108.825 52.720 ;
        RECT 109.095 66.010 120.095 66.880 ;
        RECT 109.095 54.870 110.765 66.010 ;
        RECT 111.395 65.495 116.395 65.665 ;
        RECT 111.165 55.240 111.335 65.280 ;
        RECT 116.455 55.240 116.625 65.280 ;
        RECT 117.025 54.870 117.195 66.010 ;
        RECT 117.825 65.495 118.825 65.665 ;
        RECT 117.595 55.240 117.765 65.280 ;
        RECT 118.885 55.240 119.055 65.280 ;
        RECT 119.455 54.870 120.095 66.010 ;
        RECT 109.095 52.800 120.095 54.870 ;
        RECT 109.095 49.310 110.935 52.800 ;
        RECT 112.695 52.720 120.095 52.800 ;
        RECT 111.565 52.290 112.065 52.460 ;
        RECT 111.335 50.035 111.505 52.075 ;
        RECT 112.125 50.035 112.295 52.075 ;
        RECT 111.565 49.650 112.065 49.820 ;
        RECT 112.695 49.310 115.015 52.720 ;
        RECT 115.645 52.210 116.145 52.380 ;
        RECT 109.095 48.590 115.015 49.310 ;
        RECT 102.685 45.740 108.825 46.230 ;
        RECT 109.065 47.980 112.975 48.200 ;
        RECT 97.795 45.310 101.705 45.580 ;
        RECT 109.065 45.580 110.785 47.980 ;
        RECT 111.415 47.470 111.915 47.640 ;
        RECT 111.185 46.260 111.355 47.300 ;
        RECT 111.975 46.260 112.145 47.300 ;
        RECT 111.415 45.920 111.915 46.090 ;
        RECT 112.545 45.580 112.975 47.980 ;
        RECT 113.955 46.230 115.015 48.590 ;
        RECT 115.415 46.955 115.585 51.995 ;
        RECT 116.205 46.955 116.375 51.995 ;
        RECT 115.645 46.570 116.145 46.740 ;
        RECT 116.775 46.230 116.945 52.720 ;
        RECT 117.575 52.210 118.075 52.380 ;
        RECT 117.345 46.955 117.515 51.995 ;
        RECT 118.135 46.955 118.305 51.995 ;
        RECT 117.575 46.570 118.075 46.740 ;
        RECT 118.705 46.230 120.095 52.720 ;
        RECT 120.345 66.010 140.025 66.880 ;
        RECT 120.345 54.870 122.015 66.010 ;
        RECT 122.645 65.495 127.645 65.665 ;
        RECT 122.415 55.240 122.585 65.280 ;
        RECT 127.705 55.240 127.875 65.280 ;
        RECT 128.275 54.870 128.445 66.010 ;
        RECT 130.705 65.980 140.025 66.010 ;
        RECT 129.075 65.495 130.075 65.665 ;
        RECT 128.845 55.240 129.015 65.280 ;
        RECT 130.135 55.240 130.305 65.280 ;
        RECT 130.705 54.870 132.765 65.980 ;
        RECT 133.395 65.465 138.395 65.635 ;
        RECT 133.165 55.210 133.335 65.250 ;
        RECT 138.455 55.210 138.625 65.250 ;
        RECT 120.345 54.840 132.765 54.870 ;
        RECT 139.025 54.840 140.025 65.980 ;
        RECT 120.345 54.720 140.025 54.840 ;
        RECT 120.345 53.550 140.035 54.720 ;
        RECT 120.345 52.800 131.345 53.550 ;
        RECT 120.345 49.310 122.185 52.800 ;
        RECT 123.945 52.720 131.345 52.800 ;
        RECT 122.815 52.290 123.315 52.460 ;
        RECT 122.585 50.035 122.755 52.075 ;
        RECT 123.375 50.035 123.545 52.075 ;
        RECT 122.815 49.650 123.315 49.820 ;
        RECT 123.945 49.310 126.265 52.720 ;
        RECT 126.895 52.210 127.395 52.380 ;
        RECT 120.345 48.590 126.265 49.310 ;
        RECT 113.955 45.740 120.095 46.230 ;
        RECT 120.315 47.980 124.225 48.200 ;
        RECT 109.065 45.310 112.975 45.580 ;
        RECT 120.315 45.580 122.035 47.980 ;
        RECT 122.665 47.470 123.165 47.640 ;
        RECT 122.435 46.260 122.605 47.300 ;
        RECT 123.225 46.260 123.395 47.300 ;
        RECT 122.665 45.920 123.165 46.090 ;
        RECT 123.795 45.580 124.225 47.980 ;
        RECT 125.205 46.230 126.265 48.590 ;
        RECT 126.665 46.955 126.835 51.995 ;
        RECT 127.455 46.955 127.625 51.995 ;
        RECT 126.895 46.570 127.395 46.740 ;
        RECT 128.025 46.230 128.195 52.720 ;
        RECT 128.825 52.210 129.325 52.380 ;
        RECT 128.595 46.955 128.765 51.995 ;
        RECT 129.385 46.955 129.555 51.995 ;
        RECT 128.825 46.570 129.325 46.740 ;
        RECT 129.955 46.230 131.345 52.720 ;
        RECT 125.205 45.740 131.345 46.230 ;
        RECT 120.315 45.310 124.225 45.580 ;
        RECT 25.695 39.770 29.605 40.040 ;
        RECT 18.575 39.120 24.715 39.610 ;
        RECT 18.575 32.630 19.965 39.120 ;
        RECT 20.595 38.610 21.095 38.780 ;
        RECT 20.365 33.355 20.535 38.395 ;
        RECT 21.155 33.355 21.325 38.395 ;
        RECT 20.595 32.970 21.095 33.140 ;
        RECT 21.725 32.630 21.895 39.120 ;
        RECT 22.525 38.610 23.025 38.780 ;
        RECT 22.295 33.355 22.465 38.395 ;
        RECT 23.085 33.355 23.255 38.395 ;
        RECT 23.655 36.760 24.715 39.120 ;
        RECT 25.695 37.370 26.125 39.770 ;
        RECT 26.755 39.260 27.255 39.430 ;
        RECT 26.525 38.050 26.695 39.090 ;
        RECT 27.315 38.050 27.485 39.090 ;
        RECT 26.755 37.710 27.255 37.880 ;
        RECT 27.885 37.370 29.605 39.770 ;
        RECT 36.975 39.770 40.885 40.040 ;
        RECT 25.695 37.150 29.605 37.370 ;
        RECT 29.855 39.120 35.995 39.610 ;
        RECT 23.655 36.040 29.575 36.760 ;
        RECT 22.525 32.970 23.025 33.140 ;
        RECT 23.655 32.630 25.975 36.040 ;
        RECT 26.605 35.530 27.105 35.700 ;
        RECT 26.375 33.275 26.545 35.315 ;
        RECT 27.165 33.275 27.335 35.315 ;
        RECT 26.605 32.890 27.105 33.060 ;
        RECT 18.575 32.550 25.975 32.630 ;
        RECT 27.735 32.550 29.575 36.040 ;
        RECT 18.575 30.480 29.575 32.550 ;
        RECT 18.575 19.340 19.215 30.480 ;
        RECT 19.615 20.070 19.785 30.110 ;
        RECT 20.905 20.070 21.075 30.110 ;
        RECT 19.845 19.685 20.845 19.855 ;
        RECT 21.475 19.340 21.645 30.480 ;
        RECT 22.045 20.070 22.215 30.110 ;
        RECT 27.335 20.070 27.505 30.110 ;
        RECT 22.275 19.685 27.275 19.855 ;
        RECT 27.905 19.340 29.575 30.480 ;
        RECT 18.575 18.470 29.575 19.340 ;
        RECT 29.855 32.630 31.245 39.120 ;
        RECT 31.875 38.610 32.375 38.780 ;
        RECT 31.645 33.355 31.815 38.395 ;
        RECT 32.435 33.355 32.605 38.395 ;
        RECT 31.875 32.970 32.375 33.140 ;
        RECT 33.005 32.630 33.175 39.120 ;
        RECT 33.805 38.610 34.305 38.780 ;
        RECT 33.575 33.355 33.745 38.395 ;
        RECT 34.365 33.355 34.535 38.395 ;
        RECT 34.935 36.760 35.995 39.120 ;
        RECT 36.975 37.370 37.405 39.770 ;
        RECT 38.035 39.260 38.535 39.430 ;
        RECT 37.805 38.050 37.975 39.090 ;
        RECT 38.595 38.050 38.765 39.090 ;
        RECT 38.035 37.710 38.535 37.880 ;
        RECT 39.165 37.370 40.885 39.770 ;
        RECT 48.265 39.750 52.175 40.020 ;
        RECT 36.975 37.150 40.885 37.370 ;
        RECT 41.145 39.100 47.285 39.590 ;
        RECT 34.935 36.040 40.855 36.760 ;
        RECT 33.805 32.970 34.305 33.140 ;
        RECT 34.935 32.630 37.255 36.040 ;
        RECT 37.885 35.530 38.385 35.700 ;
        RECT 37.655 33.275 37.825 35.315 ;
        RECT 38.445 33.275 38.615 35.315 ;
        RECT 37.885 32.890 38.385 33.060 ;
        RECT 29.855 32.550 37.255 32.630 ;
        RECT 39.015 32.550 40.855 36.040 ;
        RECT 29.855 30.480 40.855 32.550 ;
        RECT 29.855 19.340 30.495 30.480 ;
        RECT 30.895 20.070 31.065 30.110 ;
        RECT 32.185 20.070 32.355 30.110 ;
        RECT 31.125 19.685 32.125 19.855 ;
        RECT 32.755 19.340 32.925 30.480 ;
        RECT 33.325 20.070 33.495 30.110 ;
        RECT 38.615 20.070 38.785 30.110 ;
        RECT 33.555 19.685 38.555 19.855 ;
        RECT 39.185 19.340 40.855 30.480 ;
        RECT 29.855 18.470 40.855 19.340 ;
        RECT 41.145 32.610 42.535 39.100 ;
        RECT 43.165 38.590 43.665 38.760 ;
        RECT 42.935 33.335 43.105 38.375 ;
        RECT 43.725 33.335 43.895 38.375 ;
        RECT 43.165 32.950 43.665 33.120 ;
        RECT 44.295 32.610 44.465 39.100 ;
        RECT 45.095 38.590 45.595 38.760 ;
        RECT 44.865 33.335 45.035 38.375 ;
        RECT 45.655 33.335 45.825 38.375 ;
        RECT 46.225 36.740 47.285 39.100 ;
        RECT 48.265 37.350 48.695 39.750 ;
        RECT 49.325 39.240 49.825 39.410 ;
        RECT 49.095 38.030 49.265 39.070 ;
        RECT 49.885 38.030 50.055 39.070 ;
        RECT 49.325 37.690 49.825 37.860 ;
        RECT 50.455 37.350 52.175 39.750 ;
        RECT 59.485 39.750 63.395 40.020 ;
        RECT 48.265 37.130 52.175 37.350 ;
        RECT 52.365 39.100 58.505 39.590 ;
        RECT 46.225 36.020 52.145 36.740 ;
        RECT 45.095 32.950 45.595 33.120 ;
        RECT 46.225 32.610 48.545 36.020 ;
        RECT 49.175 35.510 49.675 35.680 ;
        RECT 48.945 33.255 49.115 35.295 ;
        RECT 49.735 33.255 49.905 35.295 ;
        RECT 49.175 32.870 49.675 33.040 ;
        RECT 41.145 32.530 48.545 32.610 ;
        RECT 50.305 32.530 52.145 36.020 ;
        RECT 41.145 30.460 52.145 32.530 ;
        RECT 41.145 19.320 41.785 30.460 ;
        RECT 42.185 20.050 42.355 30.090 ;
        RECT 43.475 20.050 43.645 30.090 ;
        RECT 42.415 19.665 43.415 19.835 ;
        RECT 44.045 19.320 44.215 30.460 ;
        RECT 44.615 20.050 44.785 30.090 ;
        RECT 49.905 20.050 50.075 30.090 ;
        RECT 44.845 19.665 49.845 19.835 ;
        RECT 50.475 19.320 52.145 30.460 ;
        RECT 41.145 18.450 52.145 19.320 ;
        RECT 52.365 32.610 53.755 39.100 ;
        RECT 54.385 38.590 54.885 38.760 ;
        RECT 54.155 33.335 54.325 38.375 ;
        RECT 54.945 33.335 55.115 38.375 ;
        RECT 54.385 32.950 54.885 33.120 ;
        RECT 55.515 32.610 55.685 39.100 ;
        RECT 56.315 38.590 56.815 38.760 ;
        RECT 56.085 33.335 56.255 38.375 ;
        RECT 56.875 33.335 57.045 38.375 ;
        RECT 57.445 36.740 58.505 39.100 ;
        RECT 59.485 37.350 59.915 39.750 ;
        RECT 60.545 39.240 61.045 39.410 ;
        RECT 60.315 38.030 60.485 39.070 ;
        RECT 61.105 38.030 61.275 39.070 ;
        RECT 60.545 37.690 61.045 37.860 ;
        RECT 61.675 37.350 63.395 39.750 ;
        RECT 70.685 39.750 74.595 40.020 ;
        RECT 59.485 37.130 63.395 37.350 ;
        RECT 63.565 39.100 69.705 39.590 ;
        RECT 57.445 36.020 63.365 36.740 ;
        RECT 56.315 32.950 56.815 33.120 ;
        RECT 57.445 32.610 59.765 36.020 ;
        RECT 60.395 35.510 60.895 35.680 ;
        RECT 60.165 33.255 60.335 35.295 ;
        RECT 60.955 33.255 61.125 35.295 ;
        RECT 60.395 32.870 60.895 33.040 ;
        RECT 52.365 32.530 59.765 32.610 ;
        RECT 61.525 32.530 63.365 36.020 ;
        RECT 52.365 30.460 63.365 32.530 ;
        RECT 52.365 19.320 53.005 30.460 ;
        RECT 53.405 20.050 53.575 30.090 ;
        RECT 54.695 20.050 54.865 30.090 ;
        RECT 53.635 19.665 54.635 19.835 ;
        RECT 55.265 19.320 55.435 30.460 ;
        RECT 55.835 20.050 56.005 30.090 ;
        RECT 61.125 20.050 61.295 30.090 ;
        RECT 56.065 19.665 61.065 19.835 ;
        RECT 61.695 19.320 63.365 30.460 ;
        RECT 52.365 18.450 63.365 19.320 ;
        RECT 63.565 32.610 64.955 39.100 ;
        RECT 65.585 38.590 66.085 38.760 ;
        RECT 65.355 33.335 65.525 38.375 ;
        RECT 66.145 33.335 66.315 38.375 ;
        RECT 65.585 32.950 66.085 33.120 ;
        RECT 66.715 32.610 66.885 39.100 ;
        RECT 67.515 38.590 68.015 38.760 ;
        RECT 67.285 33.335 67.455 38.375 ;
        RECT 68.075 33.335 68.245 38.375 ;
        RECT 68.645 36.740 69.705 39.100 ;
        RECT 70.685 37.350 71.115 39.750 ;
        RECT 71.745 39.240 72.245 39.410 ;
        RECT 71.515 38.030 71.685 39.070 ;
        RECT 72.305 38.030 72.475 39.070 ;
        RECT 71.745 37.690 72.245 37.860 ;
        RECT 72.875 37.350 74.595 39.750 ;
        RECT 81.975 39.740 85.885 40.010 ;
        RECT 70.685 37.130 74.595 37.350 ;
        RECT 74.855 39.090 80.995 39.580 ;
        RECT 68.645 36.020 74.565 36.740 ;
        RECT 67.515 32.950 68.015 33.120 ;
        RECT 68.645 32.610 70.965 36.020 ;
        RECT 71.595 35.510 72.095 35.680 ;
        RECT 71.365 33.255 71.535 35.295 ;
        RECT 72.155 33.255 72.325 35.295 ;
        RECT 71.595 32.870 72.095 33.040 ;
        RECT 63.565 32.530 70.965 32.610 ;
        RECT 72.725 32.530 74.565 36.020 ;
        RECT 63.565 30.460 74.565 32.530 ;
        RECT 63.565 19.320 64.205 30.460 ;
        RECT 64.605 20.050 64.775 30.090 ;
        RECT 65.895 20.050 66.065 30.090 ;
        RECT 64.835 19.665 65.835 19.835 ;
        RECT 66.465 19.320 66.635 30.460 ;
        RECT 67.035 20.050 67.205 30.090 ;
        RECT 72.325 20.050 72.495 30.090 ;
        RECT 67.265 19.665 72.265 19.835 ;
        RECT 72.895 19.320 74.565 30.460 ;
        RECT 63.565 18.450 74.565 19.320 ;
        RECT 74.855 32.600 76.245 39.090 ;
        RECT 76.875 38.580 77.375 38.750 ;
        RECT 76.645 33.325 76.815 38.365 ;
        RECT 77.435 33.325 77.605 38.365 ;
        RECT 76.875 32.940 77.375 33.110 ;
        RECT 78.005 32.600 78.175 39.090 ;
        RECT 78.805 38.580 79.305 38.750 ;
        RECT 78.575 33.325 78.745 38.365 ;
        RECT 79.365 33.325 79.535 38.365 ;
        RECT 79.935 36.730 80.995 39.090 ;
        RECT 81.975 37.340 82.405 39.740 ;
        RECT 83.035 39.230 83.535 39.400 ;
        RECT 82.805 38.020 82.975 39.060 ;
        RECT 83.595 38.020 83.765 39.060 ;
        RECT 83.035 37.680 83.535 37.850 ;
        RECT 84.165 37.340 85.885 39.740 ;
        RECT 93.215 39.760 97.125 40.030 ;
        RECT 81.975 37.120 85.885 37.340 ;
        RECT 86.095 39.110 92.235 39.600 ;
        RECT 79.935 36.010 85.855 36.730 ;
        RECT 78.805 32.940 79.305 33.110 ;
        RECT 79.935 32.600 82.255 36.010 ;
        RECT 82.885 35.500 83.385 35.670 ;
        RECT 82.655 33.245 82.825 35.285 ;
        RECT 83.445 33.245 83.615 35.285 ;
        RECT 82.885 32.860 83.385 33.030 ;
        RECT 74.855 32.520 82.255 32.600 ;
        RECT 84.015 32.520 85.855 36.010 ;
        RECT 74.855 30.450 85.855 32.520 ;
        RECT 74.855 19.310 75.495 30.450 ;
        RECT 75.895 20.040 76.065 30.080 ;
        RECT 77.185 20.040 77.355 30.080 ;
        RECT 76.125 19.655 77.125 19.825 ;
        RECT 77.755 19.310 77.925 30.450 ;
        RECT 78.325 20.040 78.495 30.080 ;
        RECT 83.615 20.040 83.785 30.080 ;
        RECT 78.555 19.655 83.555 19.825 ;
        RECT 84.185 19.310 85.855 30.450 ;
        RECT 74.855 18.440 85.855 19.310 ;
        RECT 86.095 32.620 87.485 39.110 ;
        RECT 88.115 38.600 88.615 38.770 ;
        RECT 87.885 33.345 88.055 38.385 ;
        RECT 88.675 33.345 88.845 38.385 ;
        RECT 88.115 32.960 88.615 33.130 ;
        RECT 89.245 32.620 89.415 39.110 ;
        RECT 90.045 38.600 90.545 38.770 ;
        RECT 89.815 33.345 89.985 38.385 ;
        RECT 90.605 33.345 90.775 38.385 ;
        RECT 91.175 36.750 92.235 39.110 ;
        RECT 93.215 37.360 93.645 39.760 ;
        RECT 94.275 39.250 94.775 39.420 ;
        RECT 94.045 38.040 94.215 39.080 ;
        RECT 94.835 38.040 95.005 39.080 ;
        RECT 94.275 37.700 94.775 37.870 ;
        RECT 95.405 37.360 97.125 39.760 ;
        RECT 104.425 39.780 108.335 40.050 ;
        RECT 93.215 37.140 97.125 37.360 ;
        RECT 97.305 39.130 103.445 39.620 ;
        RECT 91.175 36.030 97.095 36.750 ;
        RECT 90.045 32.960 90.545 33.130 ;
        RECT 91.175 32.620 93.495 36.030 ;
        RECT 94.125 35.520 94.625 35.690 ;
        RECT 93.895 33.265 94.065 35.305 ;
        RECT 94.685 33.265 94.855 35.305 ;
        RECT 94.125 32.880 94.625 33.050 ;
        RECT 86.095 32.540 93.495 32.620 ;
        RECT 95.255 32.540 97.095 36.030 ;
        RECT 86.095 30.470 97.095 32.540 ;
        RECT 86.095 19.330 86.735 30.470 ;
        RECT 87.135 20.060 87.305 30.100 ;
        RECT 88.425 20.060 88.595 30.100 ;
        RECT 87.365 19.675 88.365 19.845 ;
        RECT 88.995 19.330 89.165 30.470 ;
        RECT 89.565 20.060 89.735 30.100 ;
        RECT 94.855 20.060 95.025 30.100 ;
        RECT 89.795 19.675 94.795 19.845 ;
        RECT 95.425 19.330 97.095 30.470 ;
        RECT 86.095 18.460 97.095 19.330 ;
        RECT 97.305 32.640 98.695 39.130 ;
        RECT 99.325 38.620 99.825 38.790 ;
        RECT 99.095 33.365 99.265 38.405 ;
        RECT 99.885 33.365 100.055 38.405 ;
        RECT 99.325 32.980 99.825 33.150 ;
        RECT 100.455 32.640 100.625 39.130 ;
        RECT 101.255 38.620 101.755 38.790 ;
        RECT 101.025 33.365 101.195 38.405 ;
        RECT 101.815 33.365 101.985 38.405 ;
        RECT 102.385 36.770 103.445 39.130 ;
        RECT 104.425 37.380 104.855 39.780 ;
        RECT 105.485 39.270 105.985 39.440 ;
        RECT 105.255 38.060 105.425 39.100 ;
        RECT 106.045 38.060 106.215 39.100 ;
        RECT 105.485 37.720 105.985 37.890 ;
        RECT 106.615 37.380 108.335 39.780 ;
        RECT 115.625 39.820 119.535 40.090 ;
        RECT 104.425 37.160 108.335 37.380 ;
        RECT 108.505 39.170 114.645 39.660 ;
        RECT 102.385 36.050 108.305 36.770 ;
        RECT 101.255 32.980 101.755 33.150 ;
        RECT 102.385 32.640 104.705 36.050 ;
        RECT 105.335 35.540 105.835 35.710 ;
        RECT 105.105 33.285 105.275 35.325 ;
        RECT 105.895 33.285 106.065 35.325 ;
        RECT 105.335 32.900 105.835 33.070 ;
        RECT 97.305 32.560 104.705 32.640 ;
        RECT 106.465 32.560 108.305 36.050 ;
        RECT 97.305 30.490 108.305 32.560 ;
        RECT 97.305 19.350 97.945 30.490 ;
        RECT 98.345 20.080 98.515 30.120 ;
        RECT 99.635 20.080 99.805 30.120 ;
        RECT 98.575 19.695 99.575 19.865 ;
        RECT 100.205 19.350 100.375 30.490 ;
        RECT 100.775 20.080 100.945 30.120 ;
        RECT 106.065 20.080 106.235 30.120 ;
        RECT 101.005 19.695 106.005 19.865 ;
        RECT 106.635 19.350 108.305 30.490 ;
        RECT 97.305 18.480 108.305 19.350 ;
        RECT 108.505 32.680 109.895 39.170 ;
        RECT 110.525 38.660 111.025 38.830 ;
        RECT 110.295 33.405 110.465 38.445 ;
        RECT 111.085 33.405 111.255 38.445 ;
        RECT 110.525 33.020 111.025 33.190 ;
        RECT 111.655 32.680 111.825 39.170 ;
        RECT 112.455 38.660 112.955 38.830 ;
        RECT 112.225 33.405 112.395 38.445 ;
        RECT 113.015 33.405 113.185 38.445 ;
        RECT 113.585 36.810 114.645 39.170 ;
        RECT 115.625 37.420 116.055 39.820 ;
        RECT 116.685 39.310 117.185 39.480 ;
        RECT 116.455 38.100 116.625 39.140 ;
        RECT 117.245 38.100 117.415 39.140 ;
        RECT 116.685 37.760 117.185 37.930 ;
        RECT 117.815 37.420 119.535 39.820 ;
        RECT 126.835 39.840 130.745 40.110 ;
        RECT 115.625 37.200 119.535 37.420 ;
        RECT 119.715 39.190 125.855 39.680 ;
        RECT 113.585 36.090 119.505 36.810 ;
        RECT 112.455 33.020 112.955 33.190 ;
        RECT 113.585 32.680 115.905 36.090 ;
        RECT 116.535 35.580 117.035 35.750 ;
        RECT 116.305 33.325 116.475 35.365 ;
        RECT 117.095 33.325 117.265 35.365 ;
        RECT 116.535 32.940 117.035 33.110 ;
        RECT 108.505 32.600 115.905 32.680 ;
        RECT 117.665 32.600 119.505 36.090 ;
        RECT 108.505 30.530 119.505 32.600 ;
        RECT 108.505 19.390 109.145 30.530 ;
        RECT 109.545 20.120 109.715 30.160 ;
        RECT 110.835 20.120 111.005 30.160 ;
        RECT 109.775 19.735 110.775 19.905 ;
        RECT 111.405 19.390 111.575 30.530 ;
        RECT 111.975 20.120 112.145 30.160 ;
        RECT 117.265 20.120 117.435 30.160 ;
        RECT 112.205 19.735 117.205 19.905 ;
        RECT 117.835 19.390 119.505 30.530 ;
        RECT 108.505 18.520 119.505 19.390 ;
        RECT 119.715 32.700 121.105 39.190 ;
        RECT 121.735 38.680 122.235 38.850 ;
        RECT 121.505 33.425 121.675 38.465 ;
        RECT 122.295 33.425 122.465 38.465 ;
        RECT 121.735 33.040 122.235 33.210 ;
        RECT 122.865 32.700 123.035 39.190 ;
        RECT 123.665 38.680 124.165 38.850 ;
        RECT 123.435 33.425 123.605 38.465 ;
        RECT 124.225 33.425 124.395 38.465 ;
        RECT 124.795 36.830 125.855 39.190 ;
        RECT 126.835 37.440 127.265 39.840 ;
        RECT 127.895 39.330 128.395 39.500 ;
        RECT 127.665 38.120 127.835 39.160 ;
        RECT 128.455 38.120 128.625 39.160 ;
        RECT 127.895 37.780 128.395 37.950 ;
        RECT 129.025 37.440 130.745 39.840 ;
        RECT 126.835 37.220 130.745 37.440 ;
        RECT 124.795 36.110 130.715 36.830 ;
        RECT 123.665 33.040 124.165 33.210 ;
        RECT 124.795 32.700 127.115 36.110 ;
        RECT 127.745 35.600 128.245 35.770 ;
        RECT 127.515 33.345 127.685 35.385 ;
        RECT 128.305 33.345 128.475 35.385 ;
        RECT 127.745 32.960 128.245 33.130 ;
        RECT 119.715 32.620 127.115 32.700 ;
        RECT 128.875 32.620 130.715 36.110 ;
        RECT 119.715 31.140 130.715 32.620 ;
        RECT 119.715 30.550 139.465 31.140 ;
        RECT 119.715 19.410 120.355 30.550 ;
        RECT 120.755 20.140 120.925 30.180 ;
        RECT 122.045 20.140 122.215 30.180 ;
        RECT 120.985 19.755 121.985 19.925 ;
        RECT 122.615 19.410 122.785 30.550 ;
        RECT 129.045 30.520 139.465 30.550 ;
        RECT 123.185 20.140 123.355 30.180 ;
        RECT 128.475 20.140 128.645 30.180 ;
        RECT 123.415 19.755 128.415 19.925 ;
        RECT 129.045 19.410 132.075 30.520 ;
        RECT 132.475 20.110 132.645 30.150 ;
        RECT 137.765 20.110 137.935 30.150 ;
        RECT 132.705 19.725 137.705 19.895 ;
        RECT 119.715 19.380 132.075 19.410 ;
        RECT 138.335 19.380 139.465 30.520 ;
        RECT 119.715 18.540 139.465 19.380 ;
        RECT 131.925 18.520 139.465 18.540 ;
      LAYER met1 ;
        RECT 135.340 223.880 136.790 225.180 ;
        RECT 18.165 193.380 112.465 193.860 ;
        RECT 87.250 193.180 87.540 193.225 ;
        RECT 84.105 193.040 87.540 193.180 ;
        RECT 78.610 192.840 78.900 192.885 ;
        RECT 81.850 192.840 82.500 192.885 ;
        RECT 84.105 192.840 84.245 193.040 ;
        RECT 87.250 192.995 87.540 193.040 ;
        RECT 90.930 192.995 91.220 193.225 ;
        RECT 36.265 192.700 42.845 192.840 ;
        RECT 36.265 192.560 36.405 192.700 ;
        RECT 20.075 192.500 20.395 192.560 ;
        RECT 31.130 192.500 31.420 192.545 ;
        RECT 36.175 192.500 36.495 192.560 ;
        RECT 20.075 192.360 36.495 192.500 ;
        RECT 20.075 192.300 20.395 192.360 ;
        RECT 31.130 192.315 31.420 192.360 ;
        RECT 36.175 192.300 36.495 192.360 ;
        RECT 39.395 192.500 39.715 192.560 ;
        RECT 39.870 192.500 40.160 192.545 ;
        RECT 39.395 192.360 40.160 192.500 ;
        RECT 39.395 192.300 39.715 192.360 ;
        RECT 39.870 192.315 40.160 192.360 ;
        RECT 40.775 192.300 41.095 192.560 ;
        RECT 42.705 192.545 42.845 192.700 ;
        RECT 78.610 192.700 84.245 192.840 ;
        RECT 84.490 192.840 84.780 192.885 ;
        RECT 88.155 192.840 88.475 192.900 ;
        RECT 91.005 192.840 91.145 192.995 ;
        RECT 84.490 192.700 88.475 192.840 ;
        RECT 78.610 192.655 79.200 192.700 ;
        RECT 81.850 192.655 82.500 192.700 ;
        RECT 84.490 192.655 84.780 192.700 ;
        RECT 42.630 192.315 42.920 192.545 ;
        RECT 51.370 192.500 51.660 192.545 ;
        RECT 59.190 192.500 59.480 192.545 ;
        RECT 60.095 192.500 60.415 192.560 ;
        RECT 51.370 192.360 60.415 192.500 ;
        RECT 51.370 192.315 51.660 192.360 ;
        RECT 59.190 192.315 59.480 192.360 ;
        RECT 60.095 192.300 60.415 192.360 ;
        RECT 66.090 192.500 66.380 192.545 ;
        RECT 66.535 192.500 66.855 192.560 ;
        RECT 66.090 192.360 66.855 192.500 ;
        RECT 66.090 192.315 66.380 192.360 ;
        RECT 66.535 192.300 66.855 192.360 ;
        RECT 78.910 192.340 79.200 192.655 ;
        RECT 88.155 192.640 88.475 192.700 ;
        RECT 88.705 192.700 91.145 192.840 ;
        RECT 79.990 192.500 80.280 192.545 ;
        RECT 83.570 192.500 83.860 192.545 ;
        RECT 85.405 192.500 85.695 192.545 ;
        RECT 79.990 192.360 85.695 192.500 ;
        RECT 79.990 192.315 80.280 192.360 ;
        RECT 83.570 192.315 83.860 192.360 ;
        RECT 85.405 192.315 85.695 192.360 ;
        RECT 87.695 192.300 88.015 192.560 ;
        RECT 75.750 192.160 76.040 192.205 ;
        RECT 82.635 192.160 82.955 192.220 ;
        RECT 85.870 192.160 86.160 192.205 ;
        RECT 75.750 192.020 82.955 192.160 ;
        RECT 75.750 191.975 76.040 192.020 ;
        RECT 82.635 191.960 82.955 192.020 ;
        RECT 85.485 192.020 86.160 192.160 ;
        RECT 40.330 191.820 40.620 191.865 ;
        RECT 41.695 191.820 42.015 191.880 ;
        RECT 40.330 191.680 42.015 191.820 ;
        RECT 40.330 191.635 40.620 191.680 ;
        RECT 41.695 191.620 42.015 191.680 ;
        RECT 79.990 191.820 80.280 191.865 ;
        RECT 83.110 191.820 83.400 191.865 ;
        RECT 85.000 191.820 85.290 191.865 ;
        RECT 79.990 191.680 85.290 191.820 ;
        RECT 79.990 191.635 80.280 191.680 ;
        RECT 83.110 191.635 83.400 191.680 ;
        RECT 85.000 191.635 85.290 191.680 ;
        RECT 30.655 191.280 30.975 191.540 ;
        RECT 38.935 191.480 39.255 191.540 ;
        RECT 43.090 191.480 43.380 191.525 ;
        RECT 38.935 191.340 43.380 191.480 ;
        RECT 38.935 191.280 39.255 191.340 ;
        RECT 43.090 191.295 43.380 191.340 ;
        RECT 50.895 191.280 51.215 191.540 ;
        RECT 59.635 191.280 59.955 191.540 ;
        RECT 65.630 191.480 65.920 191.525 ;
        RECT 66.075 191.480 66.395 191.540 ;
        RECT 65.630 191.340 66.395 191.480 ;
        RECT 65.630 191.295 65.920 191.340 ;
        RECT 66.075 191.280 66.395 191.340 ;
        RECT 83.555 191.480 83.875 191.540 ;
        RECT 85.485 191.480 85.625 192.020 ;
        RECT 85.870 191.975 86.160 192.020 ;
        RECT 86.775 192.160 87.095 192.220 ;
        RECT 88.705 192.160 88.845 192.700 ;
        RECT 90.455 192.500 90.775 192.560 ;
        RECT 91.390 192.500 91.680 192.545 ;
        RECT 90.455 192.360 91.680 192.500 ;
        RECT 90.455 192.300 90.775 192.360 ;
        RECT 91.390 192.315 91.680 192.360 ;
        RECT 95.070 192.500 95.360 192.545 ;
        RECT 97.815 192.500 98.135 192.560 ;
        RECT 95.070 192.360 98.135 192.500 ;
        RECT 95.070 192.315 95.360 192.360 ;
        RECT 97.815 192.300 98.135 192.360 ;
        RECT 104.730 192.500 105.020 192.545 ;
        RECT 105.175 192.500 105.495 192.560 ;
        RECT 104.730 192.360 105.495 192.500 ;
        RECT 104.730 192.315 105.020 192.360 ;
        RECT 105.175 192.300 105.495 192.360 ;
        RECT 86.775 192.020 88.845 192.160 ;
        RECT 86.775 191.960 87.095 192.020 ;
        RECT 89.995 191.960 90.315 192.220 ;
        RECT 83.555 191.340 85.625 191.480 ;
        RECT 83.555 191.280 83.875 191.340 ;
        RECT 93.215 191.280 93.535 191.540 ;
        RECT 94.135 191.480 94.455 191.540 ;
        RECT 94.610 191.480 94.900 191.525 ;
        RECT 94.135 191.340 94.900 191.480 ;
        RECT 94.135 191.280 94.455 191.340 ;
        RECT 94.610 191.295 94.900 191.340 ;
        RECT 103.795 191.280 104.115 191.540 ;
        RECT 17.605 190.660 112.465 191.140 ;
        RECT 28.470 190.120 28.760 190.165 ;
        RECT 31.590 190.120 31.880 190.165 ;
        RECT 33.480 190.120 33.770 190.165 ;
        RECT 28.470 189.980 33.770 190.120 ;
        RECT 28.470 189.935 28.760 189.980 ;
        RECT 31.590 189.935 31.880 189.980 ;
        RECT 33.480 189.935 33.770 189.980 ;
        RECT 39.510 190.120 39.800 190.165 ;
        RECT 42.630 190.120 42.920 190.165 ;
        RECT 44.520 190.120 44.810 190.165 ;
        RECT 39.510 189.980 44.810 190.120 ;
        RECT 39.510 189.935 39.800 189.980 ;
        RECT 42.630 189.935 42.920 189.980 ;
        RECT 44.520 189.935 44.810 189.980 ;
        RECT 50.090 190.120 50.380 190.165 ;
        RECT 53.210 190.120 53.500 190.165 ;
        RECT 55.100 190.120 55.390 190.165 ;
        RECT 50.090 189.980 55.390 190.120 ;
        RECT 50.090 189.935 50.380 189.980 ;
        RECT 53.210 189.935 53.500 189.980 ;
        RECT 55.100 189.935 55.390 189.980 ;
        RECT 65.270 190.120 65.560 190.165 ;
        RECT 68.390 190.120 68.680 190.165 ;
        RECT 70.280 190.120 70.570 190.165 ;
        RECT 74.355 190.120 74.675 190.180 ;
        RECT 65.270 189.980 70.570 190.120 ;
        RECT 65.270 189.935 65.560 189.980 ;
        RECT 68.390 189.935 68.680 189.980 ;
        RECT 70.280 189.935 70.570 189.980 ;
        RECT 71.225 189.980 74.675 190.120 ;
        RECT 34.350 189.780 34.640 189.825 ;
        RECT 40.315 189.780 40.635 189.840 ;
        RECT 34.350 189.640 40.635 189.780 ;
        RECT 34.350 189.595 34.640 189.640 ;
        RECT 40.315 189.580 40.635 189.640 ;
        RECT 45.850 189.780 46.140 189.825 ;
        RECT 47.215 189.780 47.535 189.840 ;
        RECT 45.850 189.640 47.535 189.780 ;
        RECT 45.850 189.595 46.140 189.640 ;
        RECT 47.215 189.580 47.535 189.640 ;
        RECT 54.575 189.580 54.895 189.840 ;
        RECT 57.795 189.780 58.115 189.840 ;
        RECT 59.190 189.780 59.480 189.825 ;
        RECT 57.795 189.640 59.480 189.780 ;
        RECT 57.795 189.580 58.115 189.640 ;
        RECT 59.190 189.595 59.480 189.640 ;
        RECT 66.995 189.780 67.315 189.840 ;
        RECT 71.225 189.825 71.365 189.980 ;
        RECT 74.355 189.920 74.675 189.980 ;
        RECT 77.690 190.120 77.980 190.165 ;
        RECT 80.810 190.120 81.100 190.165 ;
        RECT 82.700 190.120 82.990 190.165 ;
        RECT 77.690 189.980 82.990 190.120 ;
        RECT 77.690 189.935 77.980 189.980 ;
        RECT 80.810 189.935 81.100 189.980 ;
        RECT 82.700 189.935 82.990 189.980 ;
        RECT 94.565 190.120 94.855 190.165 ;
        RECT 97.345 190.120 97.635 190.165 ;
        RECT 99.205 190.120 99.495 190.165 ;
        RECT 94.565 189.980 99.495 190.120 ;
        RECT 94.565 189.935 94.855 189.980 ;
        RECT 97.345 189.935 97.635 189.980 ;
        RECT 99.205 189.935 99.495 189.980 ;
        RECT 69.770 189.780 70.060 189.825 ;
        RECT 66.995 189.640 70.060 189.780 ;
        RECT 66.995 189.580 67.315 189.640 ;
        RECT 69.770 189.595 70.060 189.640 ;
        RECT 71.150 189.595 71.440 189.825 ;
        RECT 73.450 189.780 73.740 189.825 ;
        RECT 76.195 189.780 76.515 189.840 ;
        RECT 73.450 189.640 76.515 189.780 ;
        RECT 73.450 189.595 73.740 189.640 ;
        RECT 76.195 189.580 76.515 189.640 ;
        RECT 82.175 189.580 82.495 189.840 ;
        RECT 83.555 189.580 83.875 189.840 ;
        RECT 93.215 189.780 93.535 189.840 ;
        RECT 97.830 189.780 98.120 189.825 ;
        RECT 93.215 189.640 98.120 189.780 ;
        RECT 93.215 189.580 93.535 189.640 ;
        RECT 97.830 189.595 98.120 189.640 ;
        RECT 98.735 189.780 99.055 189.840 ;
        RECT 99.670 189.780 99.960 189.825 ;
        RECT 98.735 189.640 99.960 189.780 ;
        RECT 98.735 189.580 99.055 189.640 ;
        RECT 99.670 189.595 99.960 189.640 ;
        RECT 27.390 189.145 27.680 189.460 ;
        RECT 28.470 189.440 28.760 189.485 ;
        RECT 32.050 189.440 32.340 189.485 ;
        RECT 33.885 189.440 34.175 189.485 ;
        RECT 28.470 189.300 34.175 189.440 ;
        RECT 28.470 189.255 28.760 189.300 ;
        RECT 32.050 189.255 32.340 189.300 ;
        RECT 33.885 189.255 34.175 189.300 ;
        RECT 36.175 189.240 36.495 189.500 ;
        RECT 30.655 189.145 30.975 189.160 ;
        RECT 27.090 189.100 27.680 189.145 ;
        RECT 30.330 189.100 30.980 189.145 ;
        RECT 27.090 188.960 30.980 189.100 ;
        RECT 27.090 188.915 27.380 188.960 ;
        RECT 30.330 188.915 30.980 188.960 ;
        RECT 32.495 189.100 32.815 189.160 ;
        RECT 32.970 189.100 33.260 189.145 ;
        RECT 32.495 188.960 33.260 189.100 ;
        RECT 36.265 189.100 36.405 189.240 ;
        RECT 38.430 189.145 38.720 189.460 ;
        RECT 39.510 189.440 39.800 189.485 ;
        RECT 43.090 189.440 43.380 189.485 ;
        RECT 44.925 189.440 45.215 189.485 ;
        RECT 39.510 189.300 45.215 189.440 ;
        RECT 39.510 189.255 39.800 189.300 ;
        RECT 43.090 189.255 43.380 189.300 ;
        RECT 44.925 189.255 45.215 189.300 ;
        RECT 45.390 189.255 45.680 189.485 ;
        RECT 38.130 189.100 38.720 189.145 ;
        RECT 38.935 189.100 39.255 189.160 ;
        RECT 41.370 189.100 42.020 189.145 ;
        RECT 36.265 188.960 37.785 189.100 ;
        RECT 30.655 188.900 30.975 188.915 ;
        RECT 32.495 188.900 32.815 188.960 ;
        RECT 32.970 188.915 33.260 188.960 ;
        RECT 25.595 188.560 25.915 188.820 ;
        RECT 35.715 188.560 36.035 188.820 ;
        RECT 36.635 188.560 36.955 188.820 ;
        RECT 37.645 188.760 37.785 188.960 ;
        RECT 38.130 188.960 42.020 189.100 ;
        RECT 38.130 188.915 38.420 188.960 ;
        RECT 38.935 188.900 39.255 188.960 ;
        RECT 41.370 188.915 42.020 188.960 ;
        RECT 44.010 189.100 44.300 189.145 ;
        RECT 44.455 189.100 44.775 189.160 ;
        RECT 44.010 188.960 44.775 189.100 ;
        RECT 44.010 188.915 44.300 188.960 ;
        RECT 44.455 188.900 44.775 188.960 ;
        RECT 39.855 188.760 40.175 188.820 ;
        RECT 37.645 188.620 40.175 188.760 ;
        RECT 39.855 188.560 40.175 188.620 ;
        RECT 40.315 188.760 40.635 188.820 ;
        RECT 45.465 188.760 45.605 189.255 ;
        RECT 49.010 189.145 49.300 189.460 ;
        RECT 50.090 189.440 50.380 189.485 ;
        RECT 53.670 189.440 53.960 189.485 ;
        RECT 55.505 189.440 55.795 189.485 ;
        RECT 50.090 189.300 55.795 189.440 ;
        RECT 50.090 189.255 50.380 189.300 ;
        RECT 53.670 189.255 53.960 189.300 ;
        RECT 55.505 189.255 55.795 189.300 ;
        RECT 55.955 189.240 56.275 189.500 ;
        RECT 58.270 189.440 58.560 189.485 ;
        RECT 60.555 189.440 60.875 189.500 ;
        RECT 58.270 189.300 60.875 189.440 ;
        RECT 58.270 189.255 58.560 189.300 ;
        RECT 60.555 189.240 60.875 189.300 ;
        RECT 61.030 189.440 61.320 189.485 ;
        RECT 63.315 189.440 63.635 189.500 ;
        RECT 61.030 189.300 63.635 189.440 ;
        RECT 61.030 189.255 61.320 189.300 ;
        RECT 63.315 189.240 63.635 189.300 ;
        RECT 48.710 189.100 49.300 189.145 ;
        RECT 50.895 189.100 51.215 189.160 ;
        RECT 64.190 189.145 64.480 189.460 ;
        RECT 65.270 189.440 65.560 189.485 ;
        RECT 68.850 189.440 69.140 189.485 ;
        RECT 70.685 189.440 70.975 189.485 ;
        RECT 65.270 189.300 70.975 189.440 ;
        RECT 65.270 189.255 65.560 189.300 ;
        RECT 68.850 189.255 69.140 189.300 ;
        RECT 70.685 189.255 70.975 189.300 ;
        RECT 71.610 189.440 71.900 189.485 ;
        RECT 76.655 189.460 76.975 189.500 ;
        RECT 71.610 189.300 74.355 189.440 ;
        RECT 71.610 189.255 71.900 189.300 ;
        RECT 51.950 189.100 52.600 189.145 ;
        RECT 48.710 188.960 52.600 189.100 ;
        RECT 48.710 188.915 49.000 188.960 ;
        RECT 50.895 188.900 51.215 188.960 ;
        RECT 51.950 188.915 52.600 188.960 ;
        RECT 63.890 189.100 64.480 189.145 ;
        RECT 66.075 189.100 66.395 189.160 ;
        RECT 67.130 189.100 67.780 189.145 ;
        RECT 63.890 188.960 67.780 189.100 ;
        RECT 63.890 188.915 64.180 188.960 ;
        RECT 66.075 188.900 66.395 188.960 ;
        RECT 67.130 188.915 67.780 188.960 ;
        RECT 40.315 188.620 45.605 188.760 ;
        RECT 56.430 188.760 56.720 188.805 ;
        RECT 58.255 188.760 58.575 188.820 ;
        RECT 56.430 188.620 58.575 188.760 ;
        RECT 40.315 188.560 40.635 188.620 ;
        RECT 56.430 188.575 56.720 188.620 ;
        RECT 58.255 188.560 58.575 188.620 ;
        RECT 58.715 188.560 59.035 188.820 ;
        RECT 66.535 188.760 66.855 188.820 ;
        RECT 71.685 188.760 71.825 189.255 ;
        RECT 66.535 188.620 71.825 188.760 ;
        RECT 66.535 188.560 66.855 188.620 ;
        RECT 72.055 188.560 72.375 188.820 ;
        RECT 74.215 188.760 74.355 189.300 ;
        RECT 76.610 189.240 76.975 189.460 ;
        RECT 77.690 189.440 77.980 189.485 ;
        RECT 81.270 189.440 81.560 189.485 ;
        RECT 83.105 189.440 83.395 189.485 ;
        RECT 77.690 189.300 83.395 189.440 ;
        RECT 77.690 189.255 77.980 189.300 ;
        RECT 81.270 189.255 81.560 189.300 ;
        RECT 83.105 189.255 83.395 189.300 ;
        RECT 84.950 189.440 85.240 189.485 ;
        RECT 87.695 189.440 88.015 189.500 ;
        RECT 84.950 189.300 88.015 189.440 ;
        RECT 84.950 189.255 85.240 189.300 ;
        RECT 76.610 189.145 76.900 189.240 ;
        RECT 76.310 189.100 76.900 189.145 ;
        RECT 79.550 189.100 80.200 189.145 ;
        RECT 85.025 189.100 85.165 189.255 ;
        RECT 87.695 189.240 88.015 189.300 ;
        RECT 89.090 189.255 89.380 189.485 ;
        RECT 94.565 189.440 94.855 189.485 ;
        RECT 94.565 189.300 97.100 189.440 ;
        RECT 94.565 189.255 94.855 189.300 ;
        RECT 76.310 188.960 80.200 189.100 ;
        RECT 76.310 188.915 76.600 188.960 ;
        RECT 79.550 188.915 80.200 188.960 ;
        RECT 80.655 188.960 85.165 189.100 ;
        RECT 85.855 189.100 86.175 189.160 ;
        RECT 89.165 189.100 89.305 189.255 ;
        RECT 85.855 188.960 89.305 189.100 ;
        RECT 92.705 189.100 92.995 189.145 ;
        RECT 94.135 189.100 94.455 189.160 ;
        RECT 96.885 189.145 97.100 189.300 ;
        RECT 95.965 189.100 96.255 189.145 ;
        RECT 92.705 188.960 96.255 189.100 ;
        RECT 78.955 188.760 79.275 188.820 ;
        RECT 80.655 188.760 80.795 188.960 ;
        RECT 85.855 188.900 86.175 188.960 ;
        RECT 92.705 188.915 92.995 188.960 ;
        RECT 94.135 188.900 94.455 188.960 ;
        RECT 95.965 188.915 96.255 188.960 ;
        RECT 96.885 189.100 97.175 189.145 ;
        RECT 98.745 189.100 99.035 189.145 ;
        RECT 96.885 188.960 99.035 189.100 ;
        RECT 96.885 188.915 97.175 188.960 ;
        RECT 98.745 188.915 99.035 188.960 ;
        RECT 74.215 188.620 80.795 188.760 ;
        RECT 84.015 188.760 84.335 188.820 ;
        RECT 90.455 188.805 90.775 188.820 ;
        RECT 84.490 188.760 84.780 188.805 ;
        RECT 84.015 188.620 84.780 188.760 ;
        RECT 78.955 188.560 79.275 188.620 ;
        RECT 84.015 188.560 84.335 188.620 ;
        RECT 84.490 188.575 84.780 188.620 ;
        RECT 90.455 188.575 90.990 188.805 ;
        RECT 90.455 188.560 90.775 188.575 ;
        RECT 18.165 187.940 112.465 188.420 ;
        RECT 40.330 187.740 40.620 187.785 ;
        RECT 38.565 187.600 40.620 187.740 ;
        RECT 26.990 187.215 27.280 187.445 ;
        RECT 28.070 187.400 28.360 187.445 ;
        RECT 29.275 187.400 29.595 187.460 ;
        RECT 35.715 187.445 36.035 187.460 ;
        RECT 38.565 187.445 38.705 187.600 ;
        RECT 40.330 187.555 40.620 187.600 ;
        RECT 44.455 187.540 44.775 187.800 ;
        RECT 57.795 187.740 58.115 187.800 ;
        RECT 49.605 187.600 58.115 187.740 ;
        RECT 28.070 187.260 29.595 187.400 ;
        RECT 28.070 187.215 28.360 187.260 ;
        RECT 27.065 186.380 27.205 187.215 ;
        RECT 29.275 187.200 29.595 187.260 ;
        RECT 32.610 187.400 32.900 187.445 ;
        RECT 35.715 187.400 36.500 187.445 ;
        RECT 32.610 187.260 36.500 187.400 ;
        RECT 32.610 187.215 33.200 187.260 ;
        RECT 32.910 186.900 33.200 187.215 ;
        RECT 35.715 187.215 36.500 187.260 ;
        RECT 38.490 187.215 38.780 187.445 ;
        RECT 35.715 187.200 36.035 187.215 ;
        RECT 33.990 187.060 34.280 187.105 ;
        RECT 37.570 187.060 37.860 187.105 ;
        RECT 39.405 187.060 39.695 187.105 ;
        RECT 33.990 186.920 39.695 187.060 ;
        RECT 33.990 186.875 34.280 186.920 ;
        RECT 37.570 186.875 37.860 186.920 ;
        RECT 39.405 186.875 39.695 186.920 ;
        RECT 39.870 187.060 40.160 187.105 ;
        RECT 40.315 187.060 40.635 187.120 ;
        RECT 39.870 186.920 40.635 187.060 ;
        RECT 39.870 186.875 40.160 186.920 ;
        RECT 40.315 186.860 40.635 186.920 ;
        RECT 42.155 186.860 42.475 187.120 ;
        RECT 43.995 186.860 44.315 187.120 ;
        RECT 46.295 187.060 46.615 187.120 ;
        RECT 49.605 187.060 49.745 187.600 ;
        RECT 57.795 187.540 58.115 187.600 ;
        RECT 59.635 187.540 59.955 187.800 ;
        RECT 60.555 187.740 60.875 187.800 ;
        RECT 65.400 187.740 65.690 187.785 ;
        RECT 70.690 187.740 70.980 187.785 ;
        RECT 72.515 187.740 72.835 187.800 ;
        RECT 60.555 187.600 72.835 187.740 ;
        RECT 60.555 187.540 60.875 187.600 ;
        RECT 65.400 187.555 65.690 187.600 ;
        RECT 70.690 187.555 70.980 187.600 ;
        RECT 72.515 187.540 72.835 187.600 ;
        RECT 76.655 187.540 76.975 187.800 ;
        RECT 81.715 187.740 82.035 187.800 ;
        RECT 86.775 187.740 87.095 187.800 ;
        RECT 77.205 187.600 87.095 187.740 ;
        RECT 49.990 187.400 50.280 187.445 ;
        RECT 54.115 187.400 54.435 187.460 ;
        RECT 49.990 187.260 54.435 187.400 ;
        RECT 49.990 187.215 50.280 187.260 ;
        RECT 54.115 187.200 54.435 187.260 ;
        RECT 57.355 187.400 57.645 187.445 ;
        RECT 59.215 187.400 59.505 187.445 ;
        RECT 57.355 187.260 59.505 187.400 ;
        RECT 59.725 187.400 59.865 187.540 ;
        RECT 60.135 187.400 60.425 187.445 ;
        RECT 63.395 187.400 63.685 187.445 ;
        RECT 59.725 187.260 63.685 187.400 ;
        RECT 57.355 187.215 57.645 187.260 ;
        RECT 59.215 187.215 59.505 187.260 ;
        RECT 60.135 187.215 60.425 187.260 ;
        RECT 63.395 187.215 63.685 187.260 ;
        RECT 71.135 187.400 71.455 187.460 ;
        RECT 77.205 187.400 77.345 187.600 ;
        RECT 81.715 187.540 82.035 187.600 ;
        RECT 86.775 187.540 87.095 187.600 ;
        RECT 71.135 187.260 77.345 187.400 ;
        RECT 77.590 187.400 77.880 187.445 ;
        RECT 79.415 187.400 79.735 187.460 ;
        RECT 84.015 187.445 84.335 187.460 ;
        RECT 77.590 187.260 79.735 187.400 ;
        RECT 46.295 186.920 51.125 187.060 ;
        RECT 46.295 186.860 46.615 186.920 ;
        RECT 28.355 186.720 28.675 186.780 ;
        RECT 31.130 186.720 31.420 186.765 ;
        RECT 28.355 186.580 31.420 186.720 ;
        RECT 28.355 186.520 28.675 186.580 ;
        RECT 31.130 186.535 31.420 186.580 ;
        RECT 41.695 186.520 42.015 186.780 ;
        RECT 44.455 186.720 44.775 186.780 ;
        RECT 50.985 186.765 51.125 186.920 ;
        RECT 52.290 186.875 52.580 187.105 ;
        RECT 54.590 186.875 54.880 187.105 ;
        RECT 55.955 187.060 56.275 187.120 ;
        RECT 56.430 187.060 56.720 187.105 ;
        RECT 55.955 186.920 56.720 187.060 ;
        RECT 50.450 186.720 50.740 186.765 ;
        RECT 44.455 186.580 50.740 186.720 ;
        RECT 44.455 186.520 44.775 186.580 ;
        RECT 50.450 186.535 50.740 186.580 ;
        RECT 50.910 186.535 51.200 186.765 ;
        RECT 32.955 186.380 33.275 186.440 ;
        RECT 27.065 186.240 33.275 186.380 ;
        RECT 32.955 186.180 33.275 186.240 ;
        RECT 33.990 186.380 34.280 186.425 ;
        RECT 37.110 186.380 37.400 186.425 ;
        RECT 39.000 186.380 39.290 186.425 ;
        RECT 33.990 186.240 39.290 186.380 ;
        RECT 33.990 186.195 34.280 186.240 ;
        RECT 37.110 186.195 37.400 186.240 ;
        RECT 39.000 186.195 39.290 186.240 ;
        RECT 49.055 186.380 49.375 186.440 ;
        RECT 52.365 186.380 52.505 186.875 ;
        RECT 54.665 186.720 54.805 186.875 ;
        RECT 55.955 186.860 56.275 186.920 ;
        RECT 56.430 186.875 56.720 186.920 ;
        RECT 58.255 186.860 58.575 187.120 ;
        RECT 59.290 187.060 59.505 187.215 ;
        RECT 71.135 187.200 71.455 187.260 ;
        RECT 77.590 187.215 77.880 187.260 ;
        RECT 79.415 187.200 79.735 187.260 ;
        RECT 80.450 187.400 80.740 187.445 ;
        RECT 83.690 187.400 84.340 187.445 ;
        RECT 80.450 187.260 84.340 187.400 ;
        RECT 80.450 187.215 81.040 187.260 ;
        RECT 83.690 187.215 84.340 187.260 ;
        RECT 61.535 187.060 61.825 187.105 ;
        RECT 59.290 186.920 61.825 187.060 ;
        RECT 61.535 186.875 61.825 186.920 ;
        RECT 76.210 187.060 76.500 187.105 ;
        RECT 78.955 187.060 79.275 187.120 ;
        RECT 76.210 186.920 79.275 187.060 ;
        RECT 76.210 186.875 76.500 186.920 ;
        RECT 78.955 186.860 79.275 186.920 ;
        RECT 80.750 186.900 81.040 187.215 ;
        RECT 84.015 187.200 84.335 187.215 ;
        RECT 86.315 187.200 86.635 187.460 ;
        RECT 90.865 187.400 91.155 187.445 ;
        RECT 91.375 187.400 91.695 187.460 ;
        RECT 94.125 187.400 94.415 187.445 ;
        RECT 90.865 187.260 94.415 187.400 ;
        RECT 90.865 187.215 91.155 187.260 ;
        RECT 91.375 187.200 91.695 187.260 ;
        RECT 94.125 187.215 94.415 187.260 ;
        RECT 95.045 187.400 95.335 187.445 ;
        RECT 96.905 187.400 97.195 187.445 ;
        RECT 95.045 187.260 97.195 187.400 ;
        RECT 95.045 187.215 95.335 187.260 ;
        RECT 96.905 187.215 97.195 187.260 ;
        RECT 81.830 187.060 82.120 187.105 ;
        RECT 85.410 187.060 85.700 187.105 ;
        RECT 87.245 187.060 87.535 187.105 ;
        RECT 81.830 186.920 87.535 187.060 ;
        RECT 81.830 186.875 82.120 186.920 ;
        RECT 85.410 186.875 85.700 186.920 ;
        RECT 87.245 186.875 87.535 186.920 ;
        RECT 92.725 187.060 93.015 187.105 ;
        RECT 95.045 187.060 95.260 187.215 ;
        RECT 92.725 186.920 95.260 187.060 ;
        RECT 92.725 186.875 93.015 186.920 ;
        RECT 54.665 186.580 69.985 186.720 ;
        RECT 56.895 186.380 57.185 186.425 ;
        RECT 58.755 186.380 59.045 186.425 ;
        RECT 61.535 186.380 61.825 186.425 ;
        RECT 49.055 186.240 56.185 186.380 ;
        RECT 49.055 186.180 49.375 186.240 ;
        RECT 27.895 185.840 28.215 186.100 ;
        RECT 28.830 186.040 29.120 186.085 ;
        RECT 31.115 186.040 31.435 186.100 ;
        RECT 28.830 185.900 31.435 186.040 ;
        RECT 28.830 185.855 29.120 185.900 ;
        RECT 31.115 185.840 31.435 185.900 ;
        RECT 48.150 186.040 48.440 186.085 ;
        RECT 49.515 186.040 49.835 186.100 ;
        RECT 48.150 185.900 49.835 186.040 ;
        RECT 48.150 185.855 48.440 185.900 ;
        RECT 49.515 185.840 49.835 185.900 ;
        RECT 52.750 186.040 53.040 186.085 ;
        RECT 53.195 186.040 53.515 186.100 ;
        RECT 52.750 185.900 53.515 186.040 ;
        RECT 52.750 185.855 53.040 185.900 ;
        RECT 53.195 185.840 53.515 185.900 ;
        RECT 55.495 185.840 55.815 186.100 ;
        RECT 56.045 186.040 56.185 186.240 ;
        RECT 56.895 186.240 61.825 186.380 ;
        RECT 69.845 186.380 69.985 186.580 ;
        RECT 70.215 186.520 70.535 186.780 ;
        RECT 74.355 186.720 74.675 186.780 ;
        RECT 83.555 186.720 83.875 186.780 ;
        RECT 87.710 186.720 88.000 186.765 ;
        RECT 74.355 186.580 88.000 186.720 ;
        RECT 74.355 186.520 74.675 186.580 ;
        RECT 83.555 186.520 83.875 186.580 ;
        RECT 87.710 186.535 88.000 186.580 ;
        RECT 93.675 186.720 93.995 186.780 ;
        RECT 95.990 186.720 96.280 186.765 ;
        RECT 93.675 186.580 96.280 186.720 ;
        RECT 93.675 186.520 93.995 186.580 ;
        RECT 95.990 186.535 96.280 186.580 ;
        RECT 97.830 186.720 98.120 186.765 ;
        RECT 98.735 186.720 99.055 186.780 ;
        RECT 97.830 186.580 99.055 186.720 ;
        RECT 97.830 186.535 98.120 186.580 ;
        RECT 98.735 186.520 99.055 186.580 ;
        RECT 78.035 186.380 78.355 186.440 ;
        RECT 69.845 186.240 78.355 186.380 ;
        RECT 56.895 186.195 57.185 186.240 ;
        RECT 58.755 186.195 59.045 186.240 ;
        RECT 61.535 186.195 61.825 186.240 ;
        RECT 78.035 186.180 78.355 186.240 ;
        RECT 81.830 186.380 82.120 186.425 ;
        RECT 84.950 186.380 85.240 186.425 ;
        RECT 86.840 186.380 87.130 186.425 ;
        RECT 81.830 186.240 87.130 186.380 ;
        RECT 81.830 186.195 82.120 186.240 ;
        RECT 84.950 186.195 85.240 186.240 ;
        RECT 86.840 186.195 87.130 186.240 ;
        RECT 92.725 186.380 93.015 186.425 ;
        RECT 95.505 186.380 95.795 186.425 ;
        RECT 97.365 186.380 97.655 186.425 ;
        RECT 92.725 186.240 97.655 186.380 ;
        RECT 92.725 186.195 93.015 186.240 ;
        RECT 95.505 186.195 95.795 186.240 ;
        RECT 97.365 186.195 97.655 186.240 ;
        RECT 60.095 186.040 60.415 186.100 ;
        RECT 56.045 185.900 60.415 186.040 ;
        RECT 60.095 185.840 60.415 185.900 ;
        RECT 72.990 186.040 73.280 186.085 ;
        RECT 75.735 186.040 76.055 186.100 ;
        RECT 72.990 185.900 76.055 186.040 ;
        RECT 72.990 185.855 73.280 185.900 ;
        RECT 75.735 185.840 76.055 185.900 ;
        RECT 85.395 186.040 85.715 186.100 ;
        RECT 88.860 186.040 89.150 186.085 ;
        RECT 85.395 185.900 89.150 186.040 ;
        RECT 85.395 185.840 85.715 185.900 ;
        RECT 88.860 185.855 89.150 185.900 ;
        RECT 17.605 185.220 112.465 185.700 ;
        RECT 26.055 184.820 26.375 185.080 ;
        RECT 29.275 184.820 29.595 185.080 ;
        RECT 30.655 185.020 30.975 185.080 ;
        RECT 30.655 184.880 32.265 185.020 ;
        RECT 30.655 184.820 30.975 184.880 ;
        RECT 25.595 184.680 25.915 184.740 ;
        RECT 31.575 184.680 31.895 184.740 ;
        RECT 25.595 184.540 31.895 184.680 ;
        RECT 32.125 184.680 32.265 184.880 ;
        RECT 32.495 184.820 32.815 185.080 ;
        RECT 33.430 185.020 33.720 185.065 ;
        RECT 36.650 185.020 36.940 185.065 ;
        RECT 33.430 184.880 36.940 185.020 ;
        RECT 33.430 184.835 33.720 184.880 ;
        RECT 36.650 184.835 36.940 184.880 ;
        RECT 39.870 185.020 40.160 185.065 ;
        RECT 43.995 185.020 44.315 185.080 ;
        RECT 39.870 184.880 44.315 185.020 ;
        RECT 39.870 184.835 40.160 184.880 ;
        RECT 39.395 184.680 39.715 184.740 ;
        RECT 39.945 184.680 40.085 184.835 ;
        RECT 43.995 184.820 44.315 184.880 ;
        RECT 54.115 185.020 54.435 185.080 ;
        RECT 56.660 185.020 56.950 185.065 ;
        RECT 58.715 185.020 59.035 185.080 ;
        RECT 54.115 184.880 59.035 185.020 ;
        RECT 54.115 184.820 54.435 184.880 ;
        RECT 56.660 184.835 56.950 184.880 ;
        RECT 58.715 184.820 59.035 184.880 ;
        RECT 68.620 185.020 68.910 185.065 ;
        RECT 71.135 185.020 71.455 185.080 ;
        RECT 68.620 184.880 71.455 185.020 ;
        RECT 68.620 184.835 68.910 184.880 ;
        RECT 71.135 184.820 71.455 184.880 ;
        RECT 85.855 185.020 86.175 185.080 ;
        RECT 85.855 184.880 92.525 185.020 ;
        RECT 85.855 184.820 86.175 184.880 ;
        RECT 32.125 184.540 40.085 184.680 ;
        RECT 40.315 184.680 40.635 184.740 ;
        RECT 48.155 184.680 48.445 184.725 ;
        RECT 50.015 184.680 50.305 184.725 ;
        RECT 52.795 184.680 53.085 184.725 ;
        RECT 40.315 184.540 47.905 184.680 ;
        RECT 25.595 184.480 25.915 184.540 ;
        RECT 26.145 184.385 26.285 184.540 ;
        RECT 31.575 184.480 31.895 184.540 ;
        RECT 39.395 184.480 39.715 184.540 ;
        RECT 40.315 184.480 40.635 184.540 ;
        RECT 26.070 184.155 26.360 184.385 ;
        RECT 36.635 184.340 36.955 184.400 ;
        RECT 39.855 184.340 40.175 184.400 ;
        RECT 47.765 184.385 47.905 184.540 ;
        RECT 48.155 184.540 53.085 184.680 ;
        RECT 48.155 184.495 48.445 184.540 ;
        RECT 50.015 184.495 50.305 184.540 ;
        RECT 52.795 184.495 53.085 184.540 ;
        RECT 58.255 184.680 58.575 184.740 ;
        RECT 70.215 184.680 70.535 184.740 ;
        RECT 58.255 184.540 70.535 184.680 ;
        RECT 58.255 184.480 58.575 184.540 ;
        RECT 70.215 184.480 70.535 184.540 ;
        RECT 72.485 184.680 72.775 184.725 ;
        RECT 75.265 184.680 75.555 184.725 ;
        RECT 77.125 184.680 77.415 184.725 ;
        RECT 72.485 184.540 77.415 184.680 ;
        RECT 72.485 184.495 72.775 184.540 ;
        RECT 75.265 184.495 75.555 184.540 ;
        RECT 77.125 184.495 77.415 184.540 ;
        RECT 85.395 184.680 85.715 184.740 ;
        RECT 85.395 184.540 91.145 184.680 ;
        RECT 85.395 184.480 85.715 184.540 ;
        RECT 41.710 184.340 42.000 184.385 ;
        RECT 27.985 184.200 38.245 184.340 ;
        RECT 24.690 184.000 24.980 184.045 ;
        RECT 27.985 184.000 28.125 184.200 ;
        RECT 36.635 184.140 36.955 184.200 ;
        RECT 24.690 183.860 28.125 184.000 ;
        RECT 28.355 184.000 28.675 184.060 ;
        RECT 30.210 184.000 30.500 184.045 ;
        RECT 28.355 183.860 30.500 184.000 ;
        RECT 24.690 183.815 24.980 183.860 ;
        RECT 28.355 183.800 28.675 183.860 ;
        RECT 30.210 183.815 30.500 183.860 ;
        RECT 30.655 183.800 30.975 184.060 ;
        RECT 31.130 183.815 31.420 184.045 ;
        RECT 31.590 184.000 31.880 184.045 ;
        RECT 32.495 184.000 32.815 184.060 ;
        RECT 31.590 183.860 32.815 184.000 ;
        RECT 38.105 184.010 38.245 184.200 ;
        RECT 39.855 184.200 42.000 184.340 ;
        RECT 39.855 184.140 40.175 184.200 ;
        RECT 41.710 184.155 42.000 184.200 ;
        RECT 47.690 184.155 47.980 184.385 ;
        RECT 49.515 184.140 49.835 184.400 ;
        RECT 55.495 184.340 55.815 184.400 ;
        RECT 58.730 184.340 59.020 184.385 ;
        RECT 60.095 184.340 60.415 184.400 ;
        RECT 50.065 184.200 58.025 184.340 ;
        RECT 38.105 184.000 38.705 184.010 ;
        RECT 38.935 184.000 39.255 184.060 ;
        RECT 39.410 184.000 39.700 184.045 ;
        RECT 38.105 183.870 39.700 184.000 ;
        RECT 38.565 183.860 39.700 183.870 ;
        RECT 31.590 183.815 31.880 183.860 ;
        RECT 20.995 183.660 21.315 183.720 ;
        RECT 30.745 183.660 30.885 183.800 ;
        RECT 20.995 183.520 30.885 183.660 ;
        RECT 31.205 183.660 31.345 183.815 ;
        RECT 32.495 183.800 32.815 183.860 ;
        RECT 38.935 183.800 39.255 183.860 ;
        RECT 39.410 183.815 39.700 183.860 ;
        RECT 43.090 184.000 43.380 184.045 ;
        RECT 50.065 184.000 50.205 184.200 ;
        RECT 55.495 184.140 55.815 184.200 ;
        RECT 57.885 184.045 58.025 184.200 ;
        RECT 58.730 184.200 60.415 184.340 ;
        RECT 70.305 184.340 70.445 184.480 ;
        RECT 72.975 184.340 73.295 184.400 ;
        RECT 70.305 184.200 73.295 184.340 ;
        RECT 58.730 184.155 59.020 184.200 ;
        RECT 60.095 184.140 60.415 184.200 ;
        RECT 72.975 184.140 73.295 184.200 ;
        RECT 74.355 184.340 74.675 184.400 ;
        RECT 74.355 184.200 75.505 184.340 ;
        RECT 74.355 184.140 74.675 184.200 ;
        RECT 52.795 184.000 53.085 184.045 ;
        RECT 43.090 183.860 50.205 184.000 ;
        RECT 50.550 183.860 53.085 184.000 ;
        RECT 43.090 183.815 43.380 183.860 ;
        RECT 32.035 183.660 32.355 183.720 ;
        RECT 31.205 183.520 32.355 183.660 ;
        RECT 20.995 183.460 21.315 183.520 ;
        RECT 32.035 183.460 32.355 183.520 ;
        RECT 32.955 183.705 33.275 183.720 ;
        RECT 32.955 183.475 33.560 183.705 ;
        RECT 34.350 183.475 34.640 183.705 ;
        RECT 32.955 183.460 33.275 183.475 ;
        RECT 27.450 183.320 27.740 183.365 ;
        RECT 31.575 183.320 31.895 183.380 ;
        RECT 27.450 183.180 31.895 183.320 ;
        RECT 34.425 183.320 34.565 183.475 ;
        RECT 37.555 183.460 37.875 183.720 ;
        RECT 38.475 183.705 38.795 183.720 ;
        RECT 50.550 183.705 50.765 183.860 ;
        RECT 52.795 183.815 53.085 183.860 ;
        RECT 57.810 184.000 58.100 184.045 ;
        RECT 59.175 184.000 59.495 184.060 ;
        RECT 57.810 183.860 59.495 184.000 ;
        RECT 57.810 183.815 58.100 183.860 ;
        RECT 59.175 183.800 59.495 183.860 ;
        RECT 63.775 184.000 64.095 184.060 ;
        RECT 64.710 184.000 65.000 184.045 ;
        RECT 63.775 183.860 65.000 184.000 ;
        RECT 63.775 183.800 64.095 183.860 ;
        RECT 64.710 183.815 65.000 183.860 ;
        RECT 72.485 184.000 72.775 184.045 ;
        RECT 75.365 184.000 75.505 184.200 ;
        RECT 75.735 184.140 76.055 184.400 ;
        RECT 84.490 184.340 84.780 184.385 ;
        RECT 85.855 184.340 86.175 184.400 ;
        RECT 89.995 184.340 90.315 184.400 ;
        RECT 90.470 184.340 90.760 184.385 ;
        RECT 84.490 184.200 86.175 184.340 ;
        RECT 84.490 184.155 84.780 184.200 ;
        RECT 85.855 184.140 86.175 184.200 ;
        RECT 87.325 184.200 90.760 184.340 ;
        RECT 77.590 184.000 77.880 184.045 ;
        RECT 72.485 183.860 75.020 184.000 ;
        RECT 75.365 183.860 77.880 184.000 ;
        RECT 72.485 183.815 72.775 183.860 ;
        RECT 38.400 183.475 38.795 183.705 ;
        RECT 48.615 183.660 48.905 183.705 ;
        RECT 50.475 183.660 50.765 183.705 ;
        RECT 48.615 183.520 50.765 183.660 ;
        RECT 48.615 183.475 48.905 183.520 ;
        RECT 50.475 183.475 50.765 183.520 ;
        RECT 51.395 183.660 51.685 183.705 ;
        RECT 53.195 183.660 53.515 183.720 ;
        RECT 54.655 183.660 54.945 183.705 ;
        RECT 51.395 183.520 54.945 183.660 ;
        RECT 51.395 183.475 51.685 183.520 ;
        RECT 38.475 183.460 38.795 183.475 ;
        RECT 53.195 183.460 53.515 183.520 ;
        RECT 54.655 183.475 54.945 183.520 ;
        RECT 70.625 183.660 70.915 183.705 ;
        RECT 72.055 183.660 72.375 183.720 ;
        RECT 74.805 183.705 75.020 183.860 ;
        RECT 77.590 183.815 77.880 183.860 ;
        RECT 78.035 184.000 78.355 184.060 ;
        RECT 85.410 184.000 85.700 184.045 ;
        RECT 86.775 184.000 87.095 184.060 ;
        RECT 78.035 183.860 87.095 184.000 ;
        RECT 78.035 183.800 78.355 183.860 ;
        RECT 85.410 183.815 85.700 183.860 ;
        RECT 86.775 183.800 87.095 183.860 ;
        RECT 73.885 183.660 74.175 183.705 ;
        RECT 70.625 183.520 74.175 183.660 ;
        RECT 70.625 183.475 70.915 183.520 ;
        RECT 72.055 183.460 72.375 183.520 ;
        RECT 73.885 183.475 74.175 183.520 ;
        RECT 74.805 183.660 75.095 183.705 ;
        RECT 76.665 183.660 76.955 183.705 ;
        RECT 87.325 183.660 87.465 184.200 ;
        RECT 89.995 184.140 90.315 184.200 ;
        RECT 90.470 184.155 90.760 184.200 ;
        RECT 88.170 183.815 88.460 184.045 ;
        RECT 88.630 183.815 88.920 184.045 ;
        RECT 91.005 184.000 91.145 184.540 ;
        RECT 91.850 184.000 92.140 184.045 ;
        RECT 91.005 183.860 92.140 184.000 ;
        RECT 92.385 184.000 92.525 184.880 ;
        RECT 93.675 184.820 93.995 185.080 ;
        RECT 96.450 184.000 96.740 184.045 ;
        RECT 92.385 183.860 96.740 184.000 ;
        RECT 91.850 183.815 92.140 183.860 ;
        RECT 96.450 183.815 96.740 183.860 ;
        RECT 98.290 184.000 98.580 184.045 ;
        RECT 103.795 184.000 104.115 184.060 ;
        RECT 98.290 183.860 104.115 184.000 ;
        RECT 98.290 183.815 98.580 183.860 ;
        RECT 74.805 183.520 76.955 183.660 ;
        RECT 74.805 183.475 75.095 183.520 ;
        RECT 76.665 183.475 76.955 183.520 ;
        RECT 80.655 183.520 87.465 183.660 ;
        RECT 87.695 183.660 88.015 183.720 ;
        RECT 88.245 183.660 88.385 183.815 ;
        RECT 87.695 183.520 88.385 183.660 ;
        RECT 41.695 183.320 42.015 183.380 ;
        RECT 34.425 183.180 42.015 183.320 ;
        RECT 27.450 183.135 27.740 183.180 ;
        RECT 31.575 183.120 31.895 183.180 ;
        RECT 41.695 183.120 42.015 183.180 ;
        RECT 67.915 183.120 68.235 183.380 ;
        RECT 72.975 183.320 73.295 183.380 ;
        RECT 80.655 183.320 80.795 183.520 ;
        RECT 87.695 183.460 88.015 183.520 ;
        RECT 72.975 183.180 80.795 183.320 ;
        RECT 82.635 183.320 82.955 183.380 ;
        RECT 88.705 183.320 88.845 183.815 ;
        RECT 103.795 183.800 104.115 183.860 ;
        RECT 90.455 183.660 90.775 183.720 ;
        RECT 91.390 183.660 91.680 183.705 ;
        RECT 90.455 183.520 91.680 183.660 ;
        RECT 90.455 183.460 90.775 183.520 ;
        RECT 91.390 183.475 91.680 183.520 ;
        RECT 95.070 183.660 95.360 183.705 ;
        RECT 97.815 183.660 98.135 183.720 ;
        RECT 95.070 183.520 98.135 183.660 ;
        RECT 95.070 183.475 95.360 183.520 ;
        RECT 97.815 183.460 98.135 183.520 ;
        RECT 82.635 183.180 88.845 183.320 ;
        RECT 72.975 183.120 73.295 183.180 ;
        RECT 82.635 183.120 82.955 183.180 ;
        RECT 89.535 183.120 89.855 183.380 ;
        RECT 89.995 183.320 90.315 183.380 ;
        RECT 97.370 183.320 97.660 183.365 ;
        RECT 100.115 183.320 100.435 183.380 ;
        RECT 89.995 183.180 100.435 183.320 ;
        RECT 89.995 183.120 90.315 183.180 ;
        RECT 97.370 183.135 97.660 183.180 ;
        RECT 100.115 183.120 100.435 183.180 ;
        RECT 18.165 182.500 112.465 182.980 ;
        RECT 21.010 182.300 21.300 182.345 ;
        RECT 32.035 182.300 32.355 182.360 ;
        RECT 21.010 182.160 24.905 182.300 ;
        RECT 21.010 182.115 21.300 182.160 ;
        RECT 24.765 181.960 24.905 182.160 ;
        RECT 32.035 182.160 36.865 182.300 ;
        RECT 32.035 182.100 32.355 182.160 ;
        RECT 25.250 181.960 25.540 182.005 ;
        RECT 28.490 181.960 29.140 182.005 ;
        RECT 24.765 181.820 29.140 181.960 ;
        RECT 25.250 181.775 25.840 181.820 ;
        RECT 28.490 181.775 29.140 181.820 ;
        RECT 20.535 181.620 20.855 181.680 ;
        RECT 21.470 181.620 21.760 181.665 ;
        RECT 20.535 181.480 21.760 181.620 ;
        RECT 20.535 181.420 20.855 181.480 ;
        RECT 21.470 181.435 21.760 181.480 ;
        RECT 25.550 181.460 25.840 181.775 ;
        RECT 31.115 181.760 31.435 182.020 ;
        RECT 31.575 181.960 31.895 182.020 ;
        RECT 36.725 182.005 36.865 182.160 ;
        RECT 52.275 182.100 52.595 182.360 ;
        RECT 54.130 182.300 54.420 182.345 ;
        RECT 55.035 182.300 55.355 182.360 ;
        RECT 54.130 182.160 55.355 182.300 ;
        RECT 54.130 182.115 54.420 182.160 ;
        RECT 55.035 182.100 55.355 182.160 ;
        RECT 58.255 182.300 58.575 182.360 ;
        RECT 71.595 182.300 71.915 182.360 ;
        RECT 58.255 182.160 71.915 182.300 ;
        RECT 58.255 182.100 58.575 182.160 ;
        RECT 71.595 182.100 71.915 182.160 ;
        RECT 76.210 182.300 76.500 182.345 ;
        RECT 87.235 182.300 87.555 182.360 ;
        RECT 76.210 182.160 87.555 182.300 ;
        RECT 76.210 182.115 76.500 182.160 ;
        RECT 87.235 182.100 87.555 182.160 ;
        RECT 87.695 182.300 88.015 182.360 ;
        RECT 88.170 182.300 88.460 182.345 ;
        RECT 87.695 182.160 88.460 182.300 ;
        RECT 87.695 182.100 88.015 182.160 ;
        RECT 88.170 182.115 88.460 182.160 ;
        RECT 91.375 182.100 91.695 182.360 ;
        RECT 31.575 181.820 34.105 181.960 ;
        RECT 31.575 181.760 31.895 181.820 ;
        RECT 33.965 181.665 34.105 181.820 ;
        RECT 36.650 181.775 36.940 182.005 ;
        RECT 42.170 181.960 42.460 182.005 ;
        RECT 60.570 181.960 60.860 182.005 ;
        RECT 62.970 181.960 63.260 182.005 ;
        RECT 66.210 181.960 66.860 182.005 ;
        RECT 38.105 181.820 42.460 181.960 ;
        RECT 26.630 181.620 26.920 181.665 ;
        RECT 30.210 181.620 30.500 181.665 ;
        RECT 32.045 181.620 32.335 181.665 ;
        RECT 26.630 181.480 32.335 181.620 ;
        RECT 26.630 181.435 26.920 181.480 ;
        RECT 30.210 181.435 30.500 181.480 ;
        RECT 32.045 181.435 32.335 181.480 ;
        RECT 33.890 181.435 34.180 181.665 ;
        RECT 35.715 181.620 36.035 181.680 ;
        RECT 38.105 181.620 38.245 181.820 ;
        RECT 42.170 181.775 42.460 181.820 ;
        RECT 49.145 181.820 60.325 181.960 ;
        RECT 35.715 181.480 38.245 181.620 ;
        RECT 38.475 181.620 38.795 181.680 ;
        RECT 39.395 181.620 39.715 181.680 ;
        RECT 38.475 181.480 39.715 181.620 ;
        RECT 35.715 181.420 36.035 181.480 ;
        RECT 38.475 181.420 38.795 181.480 ;
        RECT 39.395 181.420 39.715 181.480 ;
        RECT 39.870 181.620 40.160 181.665 ;
        RECT 40.775 181.620 41.095 181.680 ;
        RECT 39.870 181.480 41.095 181.620 ;
        RECT 39.870 181.435 40.160 181.480 ;
        RECT 40.775 181.420 41.095 181.480 ;
        RECT 22.390 181.095 22.680 181.325 ;
        RECT 31.115 181.280 31.435 181.340 ;
        RECT 32.510 181.280 32.800 181.325 ;
        RECT 40.315 181.280 40.635 181.340 ;
        RECT 31.115 181.140 40.635 181.280 ;
        RECT 21.455 180.940 21.775 181.000 ;
        RECT 22.465 180.940 22.605 181.095 ;
        RECT 31.115 181.080 31.435 181.140 ;
        RECT 32.510 181.095 32.800 181.140 ;
        RECT 40.315 181.080 40.635 181.140 ;
        RECT 21.455 180.800 22.605 180.940 ;
        RECT 26.630 180.940 26.920 180.985 ;
        RECT 29.750 180.940 30.040 180.985 ;
        RECT 31.640 180.940 31.930 180.985 ;
        RECT 26.630 180.800 31.930 180.940 ;
        RECT 21.455 180.740 21.775 180.800 ;
        RECT 26.630 180.755 26.920 180.800 ;
        RECT 29.750 180.755 30.040 180.800 ;
        RECT 31.640 180.755 31.930 180.800 ;
        RECT 32.955 180.740 33.275 181.000 ;
        RECT 37.570 180.940 37.860 180.985 ;
        RECT 38.015 180.940 38.335 181.000 ;
        RECT 40.865 180.940 41.005 181.420 ;
        RECT 43.995 181.280 44.315 181.340 ;
        RECT 49.145 181.325 49.285 181.820 ;
        RECT 50.450 181.620 50.740 181.665 ;
        RECT 49.605 181.480 50.740 181.620 ;
        RECT 49.070 181.280 49.360 181.325 ;
        RECT 43.995 181.140 49.360 181.280 ;
        RECT 43.995 181.080 44.315 181.140 ;
        RECT 49.070 181.095 49.360 181.140 ;
        RECT 37.570 180.800 41.005 180.940 ;
        RECT 37.570 180.755 37.860 180.800 ;
        RECT 38.015 180.740 38.335 180.800 ;
        RECT 42.155 180.740 42.475 181.000 ;
        RECT 43.535 180.940 43.855 181.000 ;
        RECT 49.605 180.940 49.745 181.480 ;
        RECT 50.450 181.435 50.740 181.480 ;
        RECT 55.035 181.420 55.355 181.680 ;
        RECT 56.430 181.620 56.720 181.665 ;
        RECT 55.585 181.480 56.720 181.620 ;
        RECT 49.990 181.095 50.280 181.325 ;
        RECT 51.355 181.280 51.675 181.340 ;
        RECT 55.585 181.280 55.725 181.480 ;
        RECT 56.430 181.435 56.720 181.480 ;
        RECT 57.810 181.620 58.100 181.665 ;
        RECT 58.255 181.620 58.575 181.680 ;
        RECT 57.810 181.480 58.575 181.620 ;
        RECT 57.810 181.435 58.100 181.480 ;
        RECT 58.255 181.420 58.575 181.480 ;
        RECT 58.715 181.420 59.035 181.680 ;
        RECT 51.355 181.140 55.725 181.280 ;
        RECT 43.535 180.800 49.745 180.940 ;
        RECT 50.065 180.940 50.205 181.095 ;
        RECT 51.355 181.080 51.675 181.140 ;
        RECT 55.970 181.095 56.260 181.325 ;
        RECT 55.495 180.940 55.815 181.000 ;
        RECT 50.065 180.800 55.815 180.940 ;
        RECT 56.045 180.940 56.185 181.095 ;
        RECT 59.635 180.940 59.955 181.000 ;
        RECT 56.045 180.800 59.955 180.940 ;
        RECT 60.185 180.940 60.325 181.820 ;
        RECT 60.570 181.820 66.860 181.960 ;
        RECT 60.570 181.775 60.860 181.820 ;
        RECT 62.970 181.775 63.560 181.820 ;
        RECT 66.210 181.775 66.860 181.820 ;
        RECT 68.375 181.960 68.695 182.020 ;
        RECT 76.670 181.960 76.960 182.005 ;
        RECT 68.375 181.820 76.960 181.960 ;
        RECT 61.015 181.420 61.335 181.680 ;
        RECT 62.395 181.620 62.715 181.680 ;
        RECT 61.565 181.480 62.715 181.620 ;
        RECT 61.565 181.325 61.705 181.480 ;
        RECT 62.395 181.420 62.715 181.480 ;
        RECT 63.270 181.460 63.560 181.775 ;
        RECT 68.375 181.760 68.695 181.820 ;
        RECT 76.670 181.775 76.960 181.820 ;
        RECT 80.795 181.960 81.115 182.020 ;
        RECT 84.935 181.960 85.255 182.020 ;
        RECT 90.470 181.960 90.760 182.005 ;
        RECT 92.310 181.960 92.600 182.005 ;
        RECT 97.815 181.960 98.135 182.020 ;
        RECT 80.795 181.820 84.705 181.960 ;
        RECT 80.795 181.760 81.115 181.820 ;
        RECT 64.350 181.620 64.640 181.665 ;
        RECT 67.930 181.620 68.220 181.665 ;
        RECT 69.765 181.620 70.055 181.665 ;
        RECT 64.350 181.480 70.055 181.620 ;
        RECT 64.350 181.435 64.640 181.480 ;
        RECT 67.930 181.435 68.220 181.480 ;
        RECT 69.765 181.435 70.055 181.480 ;
        RECT 71.595 181.420 71.915 181.680 ;
        RECT 72.515 181.420 72.835 181.680 ;
        RECT 78.955 181.620 79.275 181.680 ;
        RECT 79.875 181.620 80.195 181.680 ;
        RECT 78.955 181.480 80.195 181.620 ;
        RECT 78.955 181.420 79.275 181.480 ;
        RECT 79.875 181.420 80.195 181.480 ;
        RECT 81.715 181.420 82.035 181.680 ;
        RECT 82.635 181.420 82.955 181.680 ;
        RECT 84.565 181.620 84.705 181.820 ;
        RECT 84.935 181.820 86.545 181.960 ;
        RECT 84.935 181.760 85.255 181.820 ;
        RECT 86.405 181.665 86.545 181.820 ;
        RECT 90.470 181.820 92.600 181.960 ;
        RECT 90.470 181.775 90.760 181.820 ;
        RECT 92.310 181.775 92.600 181.820 ;
        RECT 93.305 181.820 98.135 181.960 ;
        RECT 85.410 181.620 85.700 181.665 ;
        RECT 84.565 181.480 85.700 181.620 ;
        RECT 85.410 181.435 85.700 181.480 ;
        RECT 85.870 181.435 86.160 181.665 ;
        RECT 86.330 181.435 86.620 181.665 ;
        RECT 86.775 181.620 87.095 181.680 ;
        RECT 87.250 181.620 87.540 181.665 ;
        RECT 86.775 181.480 87.540 181.620 ;
        RECT 61.490 181.095 61.780 181.325 ;
        RECT 61.935 181.280 62.255 181.340 ;
        RECT 66.535 181.280 66.855 181.340 ;
        RECT 61.935 181.140 66.855 181.280 ;
        RECT 61.935 181.080 62.255 181.140 ;
        RECT 66.535 181.080 66.855 181.140 ;
        RECT 68.835 181.080 69.155 181.340 ;
        RECT 70.230 181.280 70.520 181.325 ;
        RECT 73.895 181.280 74.215 181.340 ;
        RECT 75.750 181.280 76.040 181.325 ;
        RECT 78.035 181.280 78.355 181.340 ;
        RECT 70.230 181.140 74.215 181.280 ;
        RECT 70.230 181.095 70.520 181.140 ;
        RECT 73.895 181.080 74.215 181.140 ;
        RECT 75.135 181.140 78.355 181.280 ;
        RECT 63.315 180.940 63.635 181.000 ;
        RECT 60.185 180.800 63.635 180.940 ;
        RECT 43.535 180.740 43.855 180.800 ;
        RECT 55.495 180.740 55.815 180.800 ;
        RECT 59.635 180.740 59.955 180.800 ;
        RECT 63.315 180.740 63.635 180.800 ;
        RECT 64.350 180.940 64.640 180.985 ;
        RECT 67.470 180.940 67.760 180.985 ;
        RECT 69.360 180.940 69.650 180.985 ;
        RECT 75.135 180.940 75.275 181.140 ;
        RECT 75.750 181.095 76.040 181.140 ;
        RECT 78.035 181.080 78.355 181.140 ;
        RECT 79.415 181.280 79.735 181.340 ;
        RECT 85.945 181.280 86.085 181.435 ;
        RECT 86.775 181.420 87.095 181.480 ;
        RECT 87.250 181.435 87.540 181.480 ;
        RECT 89.075 181.420 89.395 181.680 ;
        RECT 90.930 181.620 91.220 181.665 ;
        RECT 93.305 181.620 93.445 181.820 ;
        RECT 97.815 181.760 98.135 181.820 ;
        RECT 90.930 181.480 93.445 181.620 ;
        RECT 90.930 181.435 91.220 181.480 ;
        RECT 93.675 181.420 93.995 181.680 ;
        RECT 94.150 181.435 94.440 181.665 ;
        RECT 79.415 181.140 86.085 181.280 ;
        RECT 88.155 181.280 88.475 181.340 ;
        RECT 89.550 181.280 89.840 181.325 ;
        RECT 88.155 181.140 89.840 181.280 ;
        RECT 79.415 181.080 79.735 181.140 ;
        RECT 88.155 181.080 88.475 181.140 ;
        RECT 89.550 181.095 89.840 181.140 ;
        RECT 90.455 181.280 90.775 181.340 ;
        RECT 94.225 181.280 94.365 181.435 ;
        RECT 94.595 181.420 94.915 181.680 ;
        RECT 95.530 181.620 95.820 181.665 ;
        RECT 95.145 181.480 95.820 181.620 ;
        RECT 90.455 181.140 94.365 181.280 ;
        RECT 90.455 181.080 90.775 181.140 ;
        RECT 64.350 180.800 69.650 180.940 ;
        RECT 64.350 180.755 64.640 180.800 ;
        RECT 67.470 180.755 67.760 180.800 ;
        RECT 69.360 180.755 69.650 180.800 ;
        RECT 70.305 180.800 75.275 180.940 ;
        RECT 91.835 180.940 92.155 181.000 ;
        RECT 95.145 180.940 95.285 181.480 ;
        RECT 95.530 181.435 95.820 181.480 ;
        RECT 91.835 180.800 95.285 180.940 ;
        RECT 35.255 180.400 35.575 180.660 ;
        RECT 36.635 180.600 36.955 180.660 ;
        RECT 38.490 180.600 38.780 180.645 ;
        RECT 36.635 180.460 38.780 180.600 ;
        RECT 36.635 180.400 36.955 180.460 ;
        RECT 38.490 180.415 38.780 180.460 ;
        RECT 56.430 180.600 56.720 180.645 ;
        RECT 56.890 180.600 57.180 180.645 ;
        RECT 56.430 180.460 57.180 180.600 ;
        RECT 63.405 180.600 63.545 180.740 ;
        RECT 70.305 180.600 70.445 180.800 ;
        RECT 91.835 180.740 92.155 180.800 ;
        RECT 63.405 180.460 70.445 180.600 ;
        RECT 56.430 180.415 56.720 180.460 ;
        RECT 56.890 180.415 57.180 180.460 ;
        RECT 70.675 180.400 70.995 180.660 ;
        RECT 78.495 180.400 78.815 180.660 ;
        RECT 78.955 180.600 79.275 180.660 ;
        RECT 79.430 180.600 79.720 180.645 ;
        RECT 78.955 180.460 79.720 180.600 ;
        RECT 78.955 180.400 79.275 180.460 ;
        RECT 79.430 180.415 79.720 180.460 ;
        RECT 83.555 180.400 83.875 180.660 ;
        RECT 84.030 180.600 84.320 180.645 ;
        RECT 84.475 180.600 84.795 180.660 ;
        RECT 84.030 180.460 84.795 180.600 ;
        RECT 84.030 180.415 84.320 180.460 ;
        RECT 84.475 180.400 84.795 180.460 ;
        RECT 89.535 180.400 89.855 180.660 ;
        RECT 89.995 180.600 90.315 180.660 ;
        RECT 93.675 180.600 93.995 180.660 ;
        RECT 89.995 180.460 93.995 180.600 ;
        RECT 89.995 180.400 90.315 180.460 ;
        RECT 93.675 180.400 93.995 180.460 ;
        RECT 17.605 179.780 112.465 180.260 ;
        RECT 21.915 179.580 22.235 179.640 ;
        RECT 31.590 179.580 31.880 179.625 ;
        RECT 42.155 179.580 42.475 179.640 ;
        RECT 21.915 179.440 31.880 179.580 ;
        RECT 21.915 179.380 22.235 179.440 ;
        RECT 31.590 179.395 31.880 179.440 ;
        RECT 37.645 179.440 42.475 179.580 ;
        RECT 21.470 179.240 21.760 179.285 ;
        RECT 27.895 179.240 28.215 179.300 ;
        RECT 21.470 179.100 28.585 179.240 ;
        RECT 21.470 179.055 21.760 179.100 ;
        RECT 27.895 179.040 28.215 179.100 ;
        RECT 20.075 178.700 20.395 178.960 ;
        RECT 26.055 178.900 26.375 178.960 ;
        RECT 28.445 178.945 28.585 179.100 ;
        RECT 37.645 178.960 37.785 179.440 ;
        RECT 42.155 179.380 42.475 179.440 ;
        RECT 44.915 179.580 45.235 179.640 ;
        RECT 44.915 179.440 56.645 179.580 ;
        RECT 44.915 179.380 45.235 179.440 ;
        RECT 38.475 179.240 38.795 179.300 ;
        RECT 39.870 179.240 40.160 179.285 ;
        RECT 38.475 179.100 40.160 179.240 ;
        RECT 38.475 179.040 38.795 179.100 ;
        RECT 39.870 179.055 40.160 179.100 ;
        RECT 50.090 179.240 50.380 179.285 ;
        RECT 53.210 179.240 53.500 179.285 ;
        RECT 55.100 179.240 55.390 179.285 ;
        RECT 50.090 179.100 55.390 179.240 ;
        RECT 50.090 179.055 50.380 179.100 ;
        RECT 53.210 179.055 53.500 179.100 ;
        RECT 55.100 179.055 55.390 179.100 ;
        RECT 56.505 179.240 56.645 179.440 ;
        RECT 59.635 179.380 59.955 179.640 ;
        RECT 68.835 179.580 69.155 179.640 ;
        RECT 69.770 179.580 70.060 179.625 ;
        RECT 71.135 179.580 71.455 179.640 ;
        RECT 80.795 179.580 81.115 179.640 ;
        RECT 62.945 179.440 67.225 179.580 ;
        RECT 57.335 179.240 57.655 179.300 ;
        RECT 56.505 179.100 57.655 179.240 ;
        RECT 22.465 178.760 26.375 178.900 ;
        RECT 22.465 178.620 22.605 178.760 ;
        RECT 26.055 178.700 26.375 178.760 ;
        RECT 28.370 178.715 28.660 178.945 ;
        RECT 33.415 178.700 33.735 178.960 ;
        RECT 33.890 178.900 34.180 178.945 ;
        RECT 34.335 178.900 34.655 178.960 ;
        RECT 35.255 178.900 35.575 178.960 ;
        RECT 37.555 178.900 37.875 178.960 ;
        RECT 33.890 178.760 37.875 178.900 ;
        RECT 33.890 178.715 34.180 178.760 ;
        RECT 34.335 178.700 34.655 178.760 ;
        RECT 35.255 178.700 35.575 178.760 ;
        RECT 37.555 178.700 37.875 178.760 ;
        RECT 38.015 178.900 38.335 178.960 ;
        RECT 38.015 178.760 39.165 178.900 ;
        RECT 38.015 178.700 38.335 178.760 ;
        RECT 21.455 178.560 21.775 178.620 ;
        RECT 21.930 178.560 22.220 178.605 ;
        RECT 21.455 178.420 22.220 178.560 ;
        RECT 21.455 178.360 21.775 178.420 ;
        RECT 21.930 178.375 22.220 178.420 ;
        RECT 22.005 178.220 22.145 178.375 ;
        RECT 22.375 178.360 22.695 178.620 ;
        RECT 25.610 178.560 25.900 178.605 ;
        RECT 28.830 178.560 29.120 178.605 ;
        RECT 25.610 178.420 29.120 178.560 ;
        RECT 25.610 178.375 25.900 178.420 ;
        RECT 28.830 178.375 29.120 178.420 ;
        RECT 31.575 178.560 31.895 178.620 ;
        RECT 32.510 178.560 32.800 178.605 ;
        RECT 31.575 178.420 32.800 178.560 ;
        RECT 31.575 178.360 31.895 178.420 ;
        RECT 32.510 178.375 32.800 178.420 ;
        RECT 32.955 178.560 33.275 178.620 ;
        RECT 35.715 178.560 36.035 178.620 ;
        RECT 37.110 178.560 37.400 178.605 ;
        RECT 32.955 178.420 37.400 178.560 ;
        RECT 32.955 178.360 33.275 178.420 ;
        RECT 35.715 178.360 36.035 178.420 ;
        RECT 37.110 178.375 37.400 178.420 ;
        RECT 38.490 178.375 38.780 178.605 ;
        RECT 39.025 178.560 39.165 178.760 ;
        RECT 42.155 178.700 42.475 178.960 ;
        RECT 52.275 178.900 52.595 178.960 ;
        RECT 54.590 178.900 54.880 178.945 ;
        RECT 52.275 178.760 54.880 178.900 ;
        RECT 52.275 178.700 52.595 178.760 ;
        RECT 54.590 178.715 54.880 178.760 ;
        RECT 42.630 178.560 42.920 178.605 ;
        RECT 39.025 178.420 42.920 178.560 ;
        RECT 42.630 178.375 42.920 178.420 ;
        RECT 46.770 178.560 47.060 178.605 ;
        RECT 48.135 178.560 48.455 178.620 ;
        RECT 46.770 178.420 48.455 178.560 ;
        RECT 46.770 178.375 47.060 178.420 ;
        RECT 33.045 178.220 33.185 178.360 ;
        RECT 22.005 178.080 33.185 178.220 ;
        RECT 35.255 178.220 35.575 178.280 ;
        RECT 36.190 178.220 36.480 178.265 ;
        RECT 35.255 178.080 36.480 178.220 ;
        RECT 35.255 178.020 35.575 178.080 ;
        RECT 36.190 178.035 36.480 178.080 ;
        RECT 20.995 177.680 21.315 177.940 ;
        RECT 21.455 177.680 21.775 177.940 ;
        RECT 29.735 177.880 30.055 177.940 ;
        RECT 30.670 177.880 30.960 177.925 ;
        RECT 29.735 177.740 30.960 177.880 ;
        RECT 37.185 177.880 37.325 178.375 ;
        RECT 38.015 178.220 38.335 178.280 ;
        RECT 38.565 178.220 38.705 178.375 ;
        RECT 48.135 178.360 48.455 178.420 ;
        RECT 49.010 178.265 49.300 178.580 ;
        RECT 50.090 178.560 50.380 178.605 ;
        RECT 53.670 178.560 53.960 178.605 ;
        RECT 55.505 178.560 55.795 178.605 ;
        RECT 50.090 178.420 55.795 178.560 ;
        RECT 50.090 178.375 50.380 178.420 ;
        RECT 53.670 178.375 53.960 178.420 ;
        RECT 55.505 178.375 55.795 178.420 ;
        RECT 55.955 178.360 56.275 178.620 ;
        RECT 56.505 178.605 56.645 179.100 ;
        RECT 57.335 179.040 57.655 179.100 ;
        RECT 58.255 179.240 58.575 179.300 ;
        RECT 62.395 179.240 62.715 179.300 ;
        RECT 58.255 179.100 62.715 179.240 ;
        RECT 58.255 179.040 58.575 179.100 ;
        RECT 62.395 179.040 62.715 179.100 ;
        RECT 61.475 178.900 61.795 178.960 ;
        RECT 62.945 178.900 63.085 179.440 ;
        RECT 66.090 179.240 66.380 179.285 ;
        RECT 67.085 179.240 67.225 179.440 ;
        RECT 68.835 179.440 70.060 179.580 ;
        RECT 68.835 179.380 69.155 179.440 ;
        RECT 69.770 179.395 70.060 179.440 ;
        RECT 70.305 179.440 81.115 179.580 ;
        RECT 70.305 179.240 70.445 179.440 ;
        RECT 71.135 179.380 71.455 179.440 ;
        RECT 80.795 179.380 81.115 179.440 ;
        RECT 83.555 179.580 83.875 179.640 ;
        RECT 84.030 179.580 84.320 179.625 ;
        RECT 83.555 179.440 84.320 179.580 ;
        RECT 83.555 179.380 83.875 179.440 ;
        RECT 84.030 179.395 84.320 179.440 ;
        RECT 74.780 179.240 75.070 179.285 ;
        RECT 76.670 179.240 76.960 179.285 ;
        RECT 79.790 179.240 80.080 179.285 ;
        RECT 66.090 179.100 66.765 179.240 ;
        RECT 67.085 179.100 70.445 179.240 ;
        RECT 70.765 179.100 73.665 179.240 ;
        RECT 66.090 179.055 66.380 179.100 ;
        RECT 58.805 178.760 63.085 178.900 ;
        RECT 56.430 178.375 56.720 178.605 ;
        RECT 57.350 178.545 57.640 178.605 ;
        RECT 56.965 178.405 57.640 178.545 ;
        RECT 39.890 178.220 40.180 178.265 ;
        RECT 38.015 178.080 38.705 178.220 ;
        RECT 39.025 178.080 40.180 178.220 ;
        RECT 38.015 178.020 38.335 178.080 ;
        RECT 39.025 177.880 39.165 178.080 ;
        RECT 39.890 178.035 40.180 178.080 ;
        RECT 46.310 178.220 46.600 178.265 ;
        RECT 48.710 178.220 49.300 178.265 ;
        RECT 51.950 178.220 52.600 178.265 ;
        RECT 46.310 178.080 52.600 178.220 ;
        RECT 46.310 178.035 46.600 178.080 ;
        RECT 48.710 178.035 49.000 178.080 ;
        RECT 51.950 178.035 52.600 178.080 ;
        RECT 37.185 177.740 39.165 177.880 ;
        RECT 43.550 177.880 43.840 177.925 ;
        RECT 45.375 177.880 45.695 177.940 ;
        RECT 43.550 177.740 45.695 177.880 ;
        RECT 29.735 177.680 30.055 177.740 ;
        RECT 30.670 177.695 30.960 177.740 ;
        RECT 43.550 177.695 43.840 177.740 ;
        RECT 45.375 177.680 45.695 177.740 ;
        RECT 47.230 177.880 47.520 177.925 ;
        RECT 50.895 177.880 51.215 177.940 ;
        RECT 56.965 177.880 57.105 178.405 ;
        RECT 57.350 178.375 57.640 178.405 ;
        RECT 57.795 178.360 58.115 178.620 ;
        RECT 58.270 178.570 58.560 178.605 ;
        RECT 58.805 178.570 58.945 178.760 ;
        RECT 61.475 178.700 61.795 178.760 ;
        RECT 63.315 178.700 63.635 178.960 ;
        RECT 66.625 178.945 66.765 179.100 ;
        RECT 66.550 178.715 66.840 178.945 ;
        RECT 70.215 178.700 70.535 178.960 ;
        RECT 58.270 178.430 58.945 178.570 ;
        RECT 60.095 178.560 60.415 178.620 ;
        RECT 61.030 178.560 61.320 178.605 ;
        RECT 58.270 178.375 58.560 178.430 ;
        RECT 60.095 178.420 61.320 178.560 ;
        RECT 60.095 178.360 60.415 178.420 ;
        RECT 61.030 178.375 61.320 178.420 ;
        RECT 61.105 178.220 61.245 178.375 ;
        RECT 64.235 178.360 64.555 178.620 ;
        RECT 66.075 178.560 66.395 178.620 ;
        RECT 70.765 178.560 70.905 179.100 ;
        RECT 66.075 178.420 70.905 178.560 ;
        RECT 71.135 178.560 71.455 178.620 ;
        RECT 71.610 178.560 71.900 178.605 ;
        RECT 71.135 178.420 71.900 178.560 ;
        RECT 66.075 178.360 66.395 178.420 ;
        RECT 71.135 178.360 71.455 178.420 ;
        RECT 71.610 178.375 71.900 178.420 ;
        RECT 72.055 178.360 72.375 178.620 ;
        RECT 73.525 178.605 73.665 179.100 ;
        RECT 74.780 179.100 80.080 179.240 ;
        RECT 74.780 179.055 75.070 179.100 ;
        RECT 76.670 179.055 76.960 179.100 ;
        RECT 79.790 179.055 80.080 179.100 ;
        RECT 82.175 179.240 82.495 179.300 ;
        RECT 83.110 179.240 83.400 179.285 ;
        RECT 88.155 179.240 88.475 179.300 ;
        RECT 82.175 179.100 83.400 179.240 ;
        RECT 82.175 179.040 82.495 179.100 ;
        RECT 83.110 179.055 83.400 179.100 ;
        RECT 84.105 179.100 88.475 179.240 ;
        RECT 73.895 178.700 74.215 178.960 ;
        RECT 75.290 178.900 75.580 178.945 ;
        RECT 78.495 178.900 78.815 178.960 ;
        RECT 75.290 178.760 78.815 178.900 ;
        RECT 75.290 178.715 75.580 178.760 ;
        RECT 78.495 178.700 78.815 178.760 ;
        RECT 81.255 178.900 81.575 178.960 ;
        RECT 84.105 178.900 84.245 179.100 ;
        RECT 88.155 179.040 88.475 179.100 ;
        RECT 81.255 178.760 84.245 178.900 ;
        RECT 81.255 178.700 81.575 178.760 ;
        RECT 84.475 178.700 84.795 178.960 ;
        RECT 87.235 178.900 87.555 178.960 ;
        RECT 87.235 178.760 92.525 178.900 ;
        RECT 87.235 178.700 87.555 178.760 ;
        RECT 72.635 178.560 72.925 178.605 ;
        RECT 72.635 178.420 73.205 178.560 ;
        RECT 72.635 178.375 72.925 178.420 ;
        RECT 61.935 178.220 62.255 178.280 ;
        RECT 61.105 178.080 62.255 178.220 ;
        RECT 61.935 178.020 62.255 178.080 ;
        RECT 63.775 178.220 64.095 178.280 ;
        RECT 73.065 178.220 73.205 178.420 ;
        RECT 73.450 178.375 73.740 178.605 ;
        RECT 74.375 178.560 74.665 178.605 ;
        RECT 76.210 178.560 76.500 178.605 ;
        RECT 79.790 178.560 80.080 178.605 ;
        RECT 74.375 178.420 80.080 178.560 ;
        RECT 74.375 178.375 74.665 178.420 ;
        RECT 76.210 178.375 76.500 178.420 ;
        RECT 79.790 178.375 80.080 178.420 ;
        RECT 63.775 178.080 73.205 178.220 ;
        RECT 73.525 178.220 73.665 178.375 ;
        RECT 76.655 178.220 76.975 178.280 ;
        RECT 73.525 178.080 76.975 178.220 ;
        RECT 63.775 178.020 64.095 178.080 ;
        RECT 76.655 178.020 76.975 178.080 ;
        RECT 77.570 178.220 78.220 178.265 ;
        RECT 78.955 178.220 79.275 178.280 ;
        RECT 80.870 178.265 81.160 178.580 ;
        RECT 84.015 178.360 84.335 178.620 ;
        RECT 85.025 178.420 89.765 178.560 ;
        RECT 80.870 178.220 81.460 178.265 ;
        RECT 85.025 178.220 85.165 178.420 ;
        RECT 77.570 178.080 81.460 178.220 ;
        RECT 77.570 178.035 78.220 178.080 ;
        RECT 78.955 178.020 79.275 178.080 ;
        RECT 81.170 178.035 81.460 178.080 ;
        RECT 82.265 178.080 85.165 178.220 ;
        RECT 85.410 178.220 85.700 178.265 ;
        RECT 88.630 178.220 88.920 178.265 ;
        RECT 85.410 178.080 88.920 178.220 ;
        RECT 89.625 178.220 89.765 178.420 ;
        RECT 89.995 178.360 90.315 178.620 ;
        RECT 90.455 178.360 90.775 178.620 ;
        RECT 90.930 178.375 91.220 178.605 ;
        RECT 90.545 178.220 90.685 178.360 ;
        RECT 89.625 178.080 90.685 178.220 ;
        RECT 91.005 178.220 91.145 178.375 ;
        RECT 91.835 178.360 92.155 178.620 ;
        RECT 92.385 178.560 92.525 178.760 ;
        RECT 92.755 178.700 93.075 178.960 ;
        RECT 94.150 178.560 94.440 178.605 ;
        RECT 92.385 178.420 94.440 178.560 ;
        RECT 94.150 178.375 94.440 178.420 ;
        RECT 97.370 178.560 97.660 178.605 ;
        RECT 97.815 178.560 98.135 178.620 ;
        RECT 101.035 178.560 101.355 178.620 ;
        RECT 97.370 178.420 101.355 178.560 ;
        RECT 97.370 178.375 97.660 178.420 ;
        RECT 97.815 178.360 98.135 178.420 ;
        RECT 101.035 178.360 101.355 178.420 ;
        RECT 94.595 178.220 94.915 178.280 ;
        RECT 91.005 178.080 94.915 178.220 ;
        RECT 47.230 177.740 57.105 177.880 ;
        RECT 61.490 177.880 61.780 177.925 ;
        RECT 64.695 177.880 65.015 177.940 ;
        RECT 61.490 177.740 65.015 177.880 ;
        RECT 47.230 177.695 47.520 177.740 ;
        RECT 50.895 177.680 51.215 177.740 ;
        RECT 61.490 177.695 61.780 177.740 ;
        RECT 64.695 177.680 65.015 177.740 ;
        RECT 65.155 177.880 65.475 177.940 ;
        RECT 72.055 177.880 72.375 177.940 ;
        RECT 79.415 177.880 79.735 177.940 ;
        RECT 65.155 177.740 79.735 177.880 ;
        RECT 65.155 177.680 65.475 177.740 ;
        RECT 72.055 177.680 72.375 177.740 ;
        RECT 79.415 177.680 79.735 177.740 ;
        RECT 80.335 177.880 80.655 177.940 ;
        RECT 82.265 177.880 82.405 178.080 ;
        RECT 85.410 178.035 85.700 178.080 ;
        RECT 88.630 178.035 88.920 178.080 ;
        RECT 94.595 178.020 94.915 178.080 ;
        RECT 80.335 177.740 82.405 177.880 ;
        RECT 82.650 177.880 82.940 177.925 ;
        RECT 84.475 177.880 84.795 177.940 ;
        RECT 82.650 177.740 84.795 177.880 ;
        RECT 80.335 177.680 80.655 177.740 ;
        RECT 82.650 177.695 82.940 177.740 ;
        RECT 84.475 177.680 84.795 177.740 ;
        RECT 86.775 177.880 87.095 177.940 ;
        RECT 90.915 177.880 91.235 177.940 ;
        RECT 91.835 177.880 92.155 177.940 ;
        RECT 86.775 177.740 92.155 177.880 ;
        RECT 86.775 177.680 87.095 177.740 ;
        RECT 90.915 177.680 91.235 177.740 ;
        RECT 91.835 177.680 92.155 177.740 ;
        RECT 93.675 177.680 93.995 177.940 ;
        RECT 95.975 177.680 96.295 177.940 ;
        RECT 96.895 177.680 97.215 177.940 ;
        RECT 101.510 177.880 101.800 177.925 ;
        RECT 101.955 177.880 102.275 177.940 ;
        RECT 101.510 177.740 102.275 177.880 ;
        RECT 101.510 177.695 101.800 177.740 ;
        RECT 101.955 177.680 102.275 177.740 ;
        RECT 18.165 177.060 112.465 177.540 ;
        RECT 22.375 176.860 22.695 176.920 ;
        RECT 31.575 176.860 31.895 176.920 ;
        RECT 22.375 176.720 31.895 176.860 ;
        RECT 22.375 176.660 22.695 176.720 ;
        RECT 31.575 176.660 31.895 176.720 ;
        RECT 37.555 176.660 37.875 176.920 ;
        RECT 39.395 176.660 39.715 176.920 ;
        RECT 43.535 176.660 43.855 176.920 ;
        RECT 44.915 176.860 45.235 176.920 ;
        RECT 44.085 176.720 45.235 176.860 ;
        RECT 20.535 176.320 20.855 176.580 ;
        RECT 21.010 176.520 21.300 176.565 ;
        RECT 23.870 176.520 24.160 176.565 ;
        RECT 27.110 176.520 27.760 176.565 ;
        RECT 21.010 176.380 27.760 176.520 ;
        RECT 21.010 176.335 21.300 176.380 ;
        RECT 23.870 176.335 24.460 176.380 ;
        RECT 27.110 176.335 27.760 176.380 ;
        RECT 20.625 176.180 20.765 176.320 ;
        RECT 21.470 176.180 21.760 176.225 ;
        RECT 22.375 176.180 22.695 176.240 ;
        RECT 20.625 176.040 22.695 176.180 ;
        RECT 21.470 175.995 21.760 176.040 ;
        RECT 22.375 175.980 22.695 176.040 ;
        RECT 24.170 176.020 24.460 176.335 ;
        RECT 29.735 176.320 30.055 176.580 ;
        RECT 25.250 176.180 25.540 176.225 ;
        RECT 28.830 176.180 29.120 176.225 ;
        RECT 30.665 176.180 30.955 176.225 ;
        RECT 25.250 176.040 30.955 176.180 ;
        RECT 25.250 175.995 25.540 176.040 ;
        RECT 28.830 175.995 29.120 176.040 ;
        RECT 30.665 175.995 30.955 176.040 ;
        RECT 31.115 175.980 31.435 176.240 ;
        RECT 31.665 176.180 31.805 176.660 ;
        RECT 38.475 176.565 38.795 176.580 ;
        RECT 38.475 176.520 38.905 176.565 ;
        RECT 35.345 176.380 38.905 176.520 ;
        RECT 32.510 176.180 32.800 176.225 ;
        RECT 31.665 176.040 32.800 176.180 ;
        RECT 32.510 175.995 32.800 176.040 ;
        RECT 33.415 176.180 33.735 176.240 ;
        RECT 35.345 176.225 35.485 176.380 ;
        RECT 38.475 176.335 38.905 176.380 ;
        RECT 43.075 176.520 43.395 176.580 ;
        RECT 44.085 176.520 44.225 176.720 ;
        RECT 44.915 176.660 45.235 176.720 ;
        RECT 47.230 176.860 47.520 176.905 ;
        RECT 51.355 176.860 51.675 176.920 ;
        RECT 47.230 176.720 51.675 176.860 ;
        RECT 47.230 176.675 47.520 176.720 ;
        RECT 51.355 176.660 51.675 176.720 ;
        RECT 54.590 176.860 54.880 176.905 ;
        RECT 55.035 176.860 55.355 176.920 ;
        RECT 54.590 176.720 55.355 176.860 ;
        RECT 54.590 176.675 54.880 176.720 ;
        RECT 55.035 176.660 55.355 176.720 ;
        RECT 66.075 176.660 66.395 176.920 ;
        RECT 66.995 176.660 67.315 176.920 ;
        RECT 74.815 176.860 75.135 176.920 ;
        RECT 80.335 176.860 80.655 176.920 ;
        RECT 68.925 176.720 75.135 176.860 ;
        RECT 52.275 176.520 52.595 176.580 ;
        RECT 43.075 176.380 44.225 176.520 ;
        RECT 38.475 176.320 38.795 176.335 ;
        RECT 43.075 176.320 43.395 176.380 ;
        RECT 35.270 176.180 35.560 176.225 ;
        RECT 33.415 176.040 35.560 176.180 ;
        RECT 33.415 175.980 33.735 176.040 ;
        RECT 35.270 175.995 35.560 176.040 ;
        RECT 35.715 176.180 36.035 176.240 ;
        RECT 44.085 176.225 44.225 176.380 ;
        RECT 45.005 176.380 52.595 176.520 ;
        RECT 45.005 176.225 45.145 176.380 ;
        RECT 52.275 176.320 52.595 176.380 ;
        RECT 59.635 176.320 59.955 176.580 ;
        RECT 60.570 176.520 60.860 176.565 ;
        RECT 68.925 176.520 69.065 176.720 ;
        RECT 60.570 176.380 69.065 176.520 ;
        RECT 69.310 176.520 69.600 176.565 ;
        RECT 69.770 176.520 70.060 176.565 ;
        RECT 69.310 176.380 70.060 176.520 ;
        RECT 60.570 176.335 60.860 176.380 ;
        RECT 36.190 176.180 36.480 176.225 ;
        RECT 35.715 176.040 36.480 176.180 ;
        RECT 35.715 175.980 36.035 176.040 ;
        RECT 36.190 175.995 36.480 176.040 ;
        RECT 37.645 176.040 39.165 176.180 ;
        RECT 20.535 175.840 20.855 175.900 ;
        RECT 32.050 175.840 32.340 175.885 ;
        RECT 20.535 175.700 32.340 175.840 ;
        RECT 20.535 175.640 20.855 175.700 ;
        RECT 32.050 175.655 32.340 175.700 ;
        RECT 33.890 175.655 34.180 175.885 ;
        RECT 25.250 175.500 25.540 175.545 ;
        RECT 28.370 175.500 28.660 175.545 ;
        RECT 30.260 175.500 30.550 175.545 ;
        RECT 25.250 175.360 30.550 175.500 ;
        RECT 33.965 175.500 34.105 175.655 ;
        RECT 34.335 175.640 34.655 175.900 ;
        RECT 34.810 175.840 35.100 175.885 ;
        RECT 37.645 175.840 37.785 176.040 ;
        RECT 39.025 175.900 39.165 176.040 ;
        RECT 39.485 176.040 43.765 176.180 ;
        RECT 34.810 175.700 37.785 175.840 ;
        RECT 34.810 175.655 35.100 175.700 ;
        RECT 38.015 175.640 38.335 175.900 ;
        RECT 38.935 175.640 39.255 175.900 ;
        RECT 35.715 175.500 36.035 175.560 ;
        RECT 33.965 175.360 36.035 175.500 ;
        RECT 25.250 175.315 25.540 175.360 ;
        RECT 28.370 175.315 28.660 175.360 ;
        RECT 30.260 175.315 30.550 175.360 ;
        RECT 35.715 175.300 36.035 175.360 ;
        RECT 36.635 175.500 36.955 175.560 ;
        RECT 37.555 175.500 37.875 175.560 ;
        RECT 39.485 175.500 39.625 176.040 ;
        RECT 40.790 175.840 41.080 175.885 ;
        RECT 42.155 175.840 42.475 175.900 ;
        RECT 40.790 175.700 42.475 175.840 ;
        RECT 43.625 175.840 43.765 176.040 ;
        RECT 44.010 175.995 44.300 176.225 ;
        RECT 44.930 175.995 45.220 176.225 ;
        RECT 45.375 175.980 45.695 176.240 ;
        RECT 45.850 175.995 46.140 176.225 ;
        RECT 45.925 175.840 46.065 175.995 ;
        RECT 49.055 175.980 49.375 176.240 ;
        RECT 50.895 175.980 51.215 176.240 ;
        RECT 54.130 176.180 54.420 176.225 ;
        RECT 55.495 176.180 55.815 176.240 ;
        RECT 54.130 176.040 55.815 176.180 ;
        RECT 54.130 175.995 54.420 176.040 ;
        RECT 55.495 175.980 55.815 176.040 ;
        RECT 55.970 175.995 56.260 176.225 ;
        RECT 43.625 175.700 46.065 175.840 ;
        RECT 40.790 175.655 41.080 175.700 ;
        RECT 42.155 175.640 42.475 175.700 ;
        RECT 48.595 175.640 48.915 175.900 ;
        RECT 36.635 175.360 39.625 175.500 ;
        RECT 56.045 175.500 56.185 175.995 ;
        RECT 56.415 175.980 56.735 176.240 ;
        RECT 56.875 175.980 57.195 176.240 ;
        RECT 57.335 176.180 57.655 176.240 ;
        RECT 57.810 176.180 58.100 176.225 ;
        RECT 57.335 176.040 58.100 176.180 ;
        RECT 57.335 175.980 57.655 176.040 ;
        RECT 57.810 175.995 58.100 176.040 ;
        RECT 58.255 176.180 58.575 176.240 ;
        RECT 65.245 176.225 65.385 176.380 ;
        RECT 69.310 176.335 69.600 176.380 ;
        RECT 69.770 176.335 70.060 176.380 ;
        RECT 71.685 176.380 72.745 176.520 ;
        RECT 62.870 176.180 63.160 176.225 ;
        RECT 58.255 176.040 63.160 176.180 ;
        RECT 58.255 175.980 58.575 176.040 ;
        RECT 62.870 175.995 63.160 176.040 ;
        RECT 65.170 175.995 65.460 176.225 ;
        RECT 67.915 175.980 68.235 176.240 ;
        RECT 68.390 176.180 68.680 176.225 ;
        RECT 70.215 176.180 70.535 176.240 ;
        RECT 68.390 176.040 70.535 176.180 ;
        RECT 68.390 175.995 68.680 176.040 ;
        RECT 70.215 175.980 70.535 176.040 ;
        RECT 71.135 175.980 71.455 176.240 ;
        RECT 71.685 176.225 71.825 176.380 ;
        RECT 71.610 175.995 71.900 176.225 ;
        RECT 72.055 175.980 72.375 176.240 ;
        RECT 61.950 175.655 62.240 175.885 ;
        RECT 62.410 175.840 62.700 175.885 ;
        RECT 72.145 175.840 72.285 175.980 ;
        RECT 62.410 175.700 72.285 175.840 ;
        RECT 72.605 175.840 72.745 176.380 ;
        RECT 73.065 176.225 73.205 176.720 ;
        RECT 74.815 176.660 75.135 176.720 ;
        RECT 77.665 176.720 80.655 176.860 ;
        RECT 77.665 176.520 77.805 176.720 ;
        RECT 80.335 176.660 80.655 176.720 ;
        RECT 81.255 176.660 81.575 176.920 ;
        RECT 84.015 176.860 84.335 176.920 ;
        RECT 84.950 176.860 85.240 176.905 ;
        RECT 84.015 176.720 85.240 176.860 ;
        RECT 84.015 176.660 84.335 176.720 ;
        RECT 84.950 176.675 85.240 176.720 ;
        RECT 87.235 176.860 87.555 176.920 ;
        RECT 88.630 176.860 88.920 176.905 ;
        RECT 87.235 176.720 88.920 176.860 ;
        RECT 87.235 176.660 87.555 176.720 ;
        RECT 88.630 176.675 88.920 176.720 ;
        RECT 95.975 176.860 96.295 176.920 ;
        RECT 100.575 176.860 100.895 176.920 ;
        RECT 95.975 176.720 97.585 176.860 ;
        RECT 95.975 176.660 96.295 176.720 ;
        RECT 86.775 176.520 87.095 176.580 ;
        RECT 74.905 176.380 77.805 176.520 ;
        RECT 78.125 176.380 87.095 176.520 ;
        RECT 72.990 175.995 73.280 176.225 ;
        RECT 73.910 176.180 74.200 176.225 ;
        RECT 74.355 176.180 74.675 176.240 ;
        RECT 73.910 176.040 74.675 176.180 ;
        RECT 73.910 175.995 74.200 176.040 ;
        RECT 74.355 175.980 74.675 176.040 ;
        RECT 74.905 175.840 75.045 176.380 ;
        RECT 75.735 175.980 76.055 176.240 ;
        RECT 76.655 176.180 76.975 176.240 ;
        RECT 78.125 176.225 78.265 176.380 ;
        RECT 78.050 176.180 78.340 176.225 ;
        RECT 76.655 176.040 78.340 176.180 ;
        RECT 76.655 175.980 76.975 176.040 ;
        RECT 78.050 175.995 78.340 176.040 ;
        RECT 78.970 175.995 79.260 176.225 ;
        RECT 72.605 175.700 75.045 175.840 ;
        RECT 79.045 175.840 79.185 175.995 ;
        RECT 79.415 175.980 79.735 176.240 ;
        RECT 79.890 176.180 80.180 176.225 ;
        RECT 81.255 176.180 81.575 176.240 ;
        RECT 81.805 176.225 81.945 176.380 ;
        RECT 84.105 176.240 84.245 176.380 ;
        RECT 86.775 176.320 87.095 176.380 ;
        RECT 91.490 176.520 91.780 176.565 ;
        RECT 94.730 176.520 95.380 176.565 ;
        RECT 96.895 176.520 97.215 176.580 ;
        RECT 97.445 176.565 97.585 176.720 ;
        RECT 100.575 176.720 108.625 176.860 ;
        RECT 100.575 176.660 100.895 176.720 ;
        RECT 101.955 176.565 102.275 176.580 ;
        RECT 91.490 176.380 97.215 176.520 ;
        RECT 91.490 176.335 92.080 176.380 ;
        RECT 94.730 176.335 95.380 176.380 ;
        RECT 79.890 176.040 81.575 176.180 ;
        RECT 79.890 175.995 80.180 176.040 ;
        RECT 81.255 175.980 81.575 176.040 ;
        RECT 81.730 175.995 82.020 176.225 ;
        RECT 82.635 175.980 82.955 176.240 ;
        RECT 83.095 175.980 83.415 176.240 ;
        RECT 83.555 175.980 83.875 176.240 ;
        RECT 84.015 175.980 84.335 176.240 ;
        RECT 84.475 176.180 84.795 176.240 ;
        RECT 85.410 176.180 85.700 176.225 ;
        RECT 84.475 176.040 85.700 176.180 ;
        RECT 84.475 175.980 84.795 176.040 ;
        RECT 85.410 175.995 85.700 176.040 ;
        RECT 91.790 176.020 92.080 176.335 ;
        RECT 96.895 176.320 97.215 176.380 ;
        RECT 97.370 176.335 97.660 176.565 ;
        RECT 101.905 176.520 102.275 176.565 ;
        RECT 105.165 176.520 105.455 176.565 ;
        RECT 101.905 176.380 105.455 176.520 ;
        RECT 101.905 176.335 102.275 176.380 ;
        RECT 105.165 176.335 105.455 176.380 ;
        RECT 106.085 176.520 106.375 176.565 ;
        RECT 107.945 176.520 108.235 176.565 ;
        RECT 106.085 176.380 108.235 176.520 ;
        RECT 106.085 176.335 106.375 176.380 ;
        RECT 107.945 176.335 108.235 176.380 ;
        RECT 101.955 176.320 102.275 176.335 ;
        RECT 92.870 176.180 93.160 176.225 ;
        RECT 96.450 176.180 96.740 176.225 ;
        RECT 98.285 176.180 98.575 176.225 ;
        RECT 92.870 176.040 98.575 176.180 ;
        RECT 92.870 175.995 93.160 176.040 ;
        RECT 96.450 175.995 96.740 176.040 ;
        RECT 98.285 175.995 98.575 176.040 ;
        RECT 103.765 176.180 104.055 176.225 ;
        RECT 106.085 176.180 106.300 176.335 ;
        RECT 103.765 176.040 106.300 176.180 ;
        RECT 107.030 176.180 107.320 176.225 ;
        RECT 108.485 176.180 108.625 176.720 ;
        RECT 107.030 176.040 108.625 176.180 ;
        RECT 103.765 175.995 104.055 176.040 ;
        RECT 107.030 175.995 107.320 176.040 ;
        RECT 89.535 175.840 89.855 175.900 ;
        RECT 90.010 175.840 90.300 175.885 ;
        RECT 79.045 175.700 90.300 175.840 ;
        RECT 62.410 175.655 62.700 175.700 ;
        RECT 60.095 175.500 60.415 175.560 ;
        RECT 62.025 175.500 62.165 175.655 ;
        RECT 74.905 175.545 75.045 175.700 ;
        RECT 89.535 175.640 89.855 175.700 ;
        RECT 90.010 175.655 90.300 175.700 ;
        RECT 98.735 175.840 99.055 175.900 ;
        RECT 108.870 175.840 109.160 175.885 ;
        RECT 109.315 175.840 109.635 175.900 ;
        RECT 98.735 175.700 109.635 175.840 ;
        RECT 98.735 175.640 99.055 175.700 ;
        RECT 108.870 175.655 109.160 175.700 ;
        RECT 109.315 175.640 109.635 175.700 ;
        RECT 56.045 175.360 59.865 175.500 ;
        RECT 36.635 175.300 36.955 175.360 ;
        RECT 37.555 175.300 37.875 175.360 ;
        RECT 24.675 175.160 24.995 175.220 ;
        RECT 32.970 175.160 33.260 175.205 ;
        RECT 24.675 175.020 33.260 175.160 ;
        RECT 24.675 174.960 24.995 175.020 ;
        RECT 32.970 174.975 33.260 175.020 ;
        RECT 33.415 175.160 33.735 175.220 ;
        RECT 55.495 175.160 55.815 175.220 ;
        RECT 56.415 175.160 56.735 175.220 ;
        RECT 33.415 175.020 56.735 175.160 ;
        RECT 33.415 174.960 33.735 175.020 ;
        RECT 55.495 174.960 55.815 175.020 ;
        RECT 56.415 174.960 56.735 175.020 ;
        RECT 56.875 175.160 57.195 175.220 ;
        RECT 59.175 175.160 59.495 175.220 ;
        RECT 56.875 175.020 59.495 175.160 ;
        RECT 59.725 175.160 59.865 175.360 ;
        RECT 60.095 175.360 62.165 175.500 ;
        RECT 60.095 175.300 60.415 175.360 ;
        RECT 74.830 175.315 75.120 175.545 ;
        RECT 76.655 175.300 76.975 175.560 ;
        RECT 82.175 175.500 82.495 175.560 ;
        RECT 83.555 175.500 83.875 175.560 ;
        RECT 82.175 175.360 83.875 175.500 ;
        RECT 82.175 175.300 82.495 175.360 ;
        RECT 83.555 175.300 83.875 175.360 ;
        RECT 92.870 175.500 93.160 175.545 ;
        RECT 95.990 175.500 96.280 175.545 ;
        RECT 97.880 175.500 98.170 175.545 ;
        RECT 92.870 175.360 98.170 175.500 ;
        RECT 92.870 175.315 93.160 175.360 ;
        RECT 95.990 175.315 96.280 175.360 ;
        RECT 97.880 175.315 98.170 175.360 ;
        RECT 103.765 175.500 104.055 175.545 ;
        RECT 106.545 175.500 106.835 175.545 ;
        RECT 108.405 175.500 108.695 175.545 ;
        RECT 103.765 175.360 108.695 175.500 ;
        RECT 103.765 175.315 104.055 175.360 ;
        RECT 106.545 175.315 106.835 175.360 ;
        RECT 108.405 175.315 108.695 175.360 ;
        RECT 60.555 175.160 60.875 175.220 ;
        RECT 59.725 175.020 60.875 175.160 ;
        RECT 56.875 174.960 57.195 175.020 ;
        RECT 59.175 174.960 59.495 175.020 ;
        RECT 60.555 174.960 60.875 175.020 ;
        RECT 62.855 175.160 63.175 175.220 ;
        RECT 64.710 175.160 65.000 175.205 ;
        RECT 62.855 175.020 65.000 175.160 ;
        RECT 62.855 174.960 63.175 175.020 ;
        RECT 64.710 174.975 65.000 175.020 ;
        RECT 69.310 175.160 69.600 175.205 ;
        RECT 70.675 175.160 70.995 175.220 ;
        RECT 69.310 175.020 70.995 175.160 ;
        RECT 69.310 174.975 69.600 175.020 ;
        RECT 70.675 174.960 70.995 175.020 ;
        RECT 72.515 175.160 72.835 175.220 ;
        RECT 83.095 175.160 83.415 175.220 ;
        RECT 86.775 175.160 87.095 175.220 ;
        RECT 72.515 175.020 87.095 175.160 ;
        RECT 72.515 174.960 72.835 175.020 ;
        RECT 83.095 174.960 83.415 175.020 ;
        RECT 86.775 174.960 87.095 175.020 ;
        RECT 94.595 175.160 94.915 175.220 ;
        RECT 99.900 175.160 100.190 175.205 ;
        RECT 94.595 175.020 100.190 175.160 ;
        RECT 94.595 174.960 94.915 175.020 ;
        RECT 99.900 174.975 100.190 175.020 ;
        RECT 17.605 174.340 112.465 174.820 ;
        RECT 135.635 174.550 136.775 223.880 ;
        RECT 138.130 223.810 139.580 225.110 ;
        RECT 143.180 223.840 144.630 225.140 ;
        RECT 35.715 174.140 36.035 174.200 ;
        RECT 59.175 174.140 59.495 174.200 ;
        RECT 35.715 174.000 59.495 174.140 ;
        RECT 35.715 173.940 36.035 174.000 ;
        RECT 59.175 173.940 59.495 174.000 ;
        RECT 60.555 174.140 60.875 174.200 ;
        RECT 70.000 174.140 70.290 174.185 ;
        RECT 72.055 174.140 72.375 174.200 ;
        RECT 89.075 174.140 89.395 174.200 ;
        RECT 90.010 174.140 90.300 174.185 ;
        RECT 97.815 174.140 98.135 174.200 ;
        RECT 60.555 174.000 66.995 174.140 ;
        RECT 60.555 173.940 60.875 174.000 ;
        RECT 36.175 173.600 36.495 173.860 ;
        RECT 36.635 173.800 36.955 173.860 ;
        RECT 46.870 173.800 47.160 173.845 ;
        RECT 49.990 173.800 50.280 173.845 ;
        RECT 51.880 173.800 52.170 173.845 ;
        RECT 61.015 173.800 61.335 173.860 ;
        RECT 36.635 173.660 39.165 173.800 ;
        RECT 36.635 173.600 36.955 173.660 ;
        RECT 21.455 173.460 21.775 173.520 ;
        RECT 27.450 173.460 27.740 173.505 ;
        RECT 34.335 173.460 34.655 173.520 ;
        RECT 37.570 173.460 37.860 173.505 ;
        RECT 21.455 173.320 37.860 173.460 ;
        RECT 21.455 173.260 21.775 173.320 ;
        RECT 27.450 173.275 27.740 173.320 ;
        RECT 34.335 173.260 34.655 173.320 ;
        RECT 37.570 173.275 37.860 173.320 ;
        RECT 38.015 173.260 38.335 173.520 ;
        RECT 38.475 173.260 38.795 173.520 ;
        RECT 39.025 173.505 39.165 173.660 ;
        RECT 46.870 173.660 52.170 173.800 ;
        RECT 46.870 173.615 47.160 173.660 ;
        RECT 49.990 173.615 50.280 173.660 ;
        RECT 51.880 173.615 52.170 173.660 ;
        RECT 52.365 173.660 61.335 173.800 ;
        RECT 38.950 173.275 39.240 173.505 ;
        RECT 52.365 173.460 52.505 173.660 ;
        RECT 61.015 173.600 61.335 173.660 ;
        RECT 61.495 173.800 61.785 173.845 ;
        RECT 63.355 173.800 63.645 173.845 ;
        RECT 66.135 173.800 66.425 173.845 ;
        RECT 61.495 173.660 66.425 173.800 ;
        RECT 61.495 173.615 61.785 173.660 ;
        RECT 63.355 173.615 63.645 173.660 ;
        RECT 66.135 173.615 66.425 173.660 ;
        RECT 41.325 173.320 52.505 173.460 ;
        RECT 41.325 173.180 41.465 173.320 ;
        RECT 56.875 173.260 57.195 173.520 ;
        RECT 57.795 173.260 58.115 173.520 ;
        RECT 62.855 173.260 63.175 173.520 ;
        RECT 66.855 173.460 66.995 174.000 ;
        RECT 70.000 174.000 75.965 174.140 ;
        RECT 70.000 173.955 70.290 174.000 ;
        RECT 72.055 173.940 72.375 174.000 ;
        RECT 67.915 173.800 68.235 173.860 ;
        RECT 70.690 173.800 70.980 173.845 ;
        RECT 67.915 173.660 70.980 173.800 ;
        RECT 75.825 173.800 75.965 174.000 ;
        RECT 89.075 174.000 90.300 174.140 ;
        RECT 89.075 173.940 89.395 174.000 ;
        RECT 90.010 173.955 90.300 174.000 ;
        RECT 94.685 174.000 98.135 174.140 ;
        RECT 94.685 173.800 94.825 174.000 ;
        RECT 97.815 173.940 98.135 174.000 ;
        RECT 100.575 173.940 100.895 174.200 ;
        RECT 75.825 173.660 89.305 173.800 ;
        RECT 67.915 173.600 68.235 173.660 ;
        RECT 70.690 173.615 70.980 173.660 ;
        RECT 82.175 173.460 82.495 173.520 ;
        RECT 66.855 173.320 82.495 173.460 ;
        RECT 22.375 172.920 22.695 173.180 ;
        RECT 28.355 172.920 28.675 173.180 ;
        RECT 33.890 173.120 34.180 173.165 ;
        RECT 35.255 173.120 35.575 173.180 ;
        RECT 41.235 173.120 41.555 173.180 ;
        RECT 33.890 172.980 35.575 173.120 ;
        RECT 33.890 172.935 34.180 172.980 ;
        RECT 35.255 172.920 35.575 172.980 ;
        RECT 40.865 172.980 41.555 173.120 ;
        RECT 31.130 172.780 31.420 172.825 ;
        RECT 36.175 172.780 36.495 172.840 ;
        RECT 36.650 172.780 36.940 172.825 ;
        RECT 40.865 172.780 41.005 172.980 ;
        RECT 41.235 172.920 41.555 172.980 ;
        RECT 41.695 172.920 42.015 173.180 ;
        RECT 42.155 172.920 42.475 173.180 ;
        RECT 43.075 172.920 43.395 173.180 ;
        RECT 31.130 172.640 36.940 172.780 ;
        RECT 31.130 172.595 31.420 172.640 ;
        RECT 36.175 172.580 36.495 172.640 ;
        RECT 36.650 172.595 36.940 172.640 ;
        RECT 38.565 172.640 41.005 172.780 ;
        RECT 42.245 172.780 42.385 172.920 ;
        RECT 45.790 172.825 46.080 173.140 ;
        RECT 46.870 173.120 47.160 173.165 ;
        RECT 50.450 173.120 50.740 173.165 ;
        RECT 52.285 173.120 52.575 173.165 ;
        RECT 46.870 172.980 52.575 173.120 ;
        RECT 46.870 172.935 47.160 172.980 ;
        RECT 50.450 172.935 50.740 172.980 ;
        RECT 52.285 172.935 52.575 172.980 ;
        RECT 52.750 173.120 53.040 173.165 ;
        RECT 55.955 173.120 56.275 173.180 ;
        RECT 61.015 173.120 61.335 173.180 ;
        RECT 72.145 173.165 72.285 173.320 ;
        RECT 82.175 173.260 82.495 173.320 ;
        RECT 83.095 173.260 83.415 173.520 ;
        RECT 83.555 173.460 83.875 173.520 ;
        RECT 83.555 173.320 88.845 173.460 ;
        RECT 83.555 173.260 83.875 173.320 ;
        RECT 66.135 173.120 66.425 173.165 ;
        RECT 52.750 172.980 61.335 173.120 ;
        RECT 52.750 172.935 53.040 172.980 ;
        RECT 55.955 172.920 56.275 172.980 ;
        RECT 61.015 172.920 61.335 172.980 ;
        RECT 63.890 172.980 66.425 173.120 ;
        RECT 45.490 172.780 46.080 172.825 ;
        RECT 48.595 172.825 48.915 172.840 ;
        RECT 48.595 172.780 49.380 172.825 ;
        RECT 42.245 172.640 44.225 172.780 ;
        RECT 22.835 172.240 23.155 172.500 ;
        RECT 30.670 172.440 30.960 172.485 ;
        RECT 32.955 172.440 33.275 172.500 ;
        RECT 30.670 172.300 33.275 172.440 ;
        RECT 30.670 172.255 30.960 172.300 ;
        RECT 32.955 172.240 33.275 172.300 ;
        RECT 33.430 172.440 33.720 172.485 ;
        RECT 38.565 172.440 38.705 172.640 ;
        RECT 44.085 172.500 44.225 172.640 ;
        RECT 45.490 172.640 49.380 172.780 ;
        RECT 45.490 172.595 45.780 172.640 ;
        RECT 48.595 172.595 49.380 172.640 ;
        RECT 48.595 172.580 48.915 172.595 ;
        RECT 51.355 172.580 51.675 172.840 ;
        RECT 55.035 172.780 55.355 172.840 ;
        RECT 59.635 172.780 59.955 172.840 ;
        RECT 63.890 172.825 64.105 172.980 ;
        RECT 66.135 172.935 66.425 172.980 ;
        RECT 72.070 172.935 72.360 173.165 ;
        RECT 72.515 172.920 72.835 173.180 ;
        RECT 72.990 172.935 73.280 173.165 ;
        RECT 73.910 173.120 74.200 173.165 ;
        RECT 74.815 173.120 75.135 173.180 ;
        RECT 75.735 173.120 76.055 173.180 ;
        RECT 73.910 172.980 76.055 173.120 ;
        RECT 73.910 172.935 74.200 172.980 ;
        RECT 55.035 172.640 59.955 172.780 ;
        RECT 55.035 172.580 55.355 172.640 ;
        RECT 59.635 172.580 59.955 172.640 ;
        RECT 61.955 172.780 62.245 172.825 ;
        RECT 63.815 172.780 64.105 172.825 ;
        RECT 61.955 172.640 64.105 172.780 ;
        RECT 61.955 172.595 62.245 172.640 ;
        RECT 63.815 172.595 64.105 172.640 ;
        RECT 64.695 172.825 65.015 172.840 ;
        RECT 64.695 172.780 65.025 172.825 ;
        RECT 67.995 172.780 68.285 172.825 ;
        RECT 64.695 172.640 68.285 172.780 ;
        RECT 64.695 172.595 65.025 172.640 ;
        RECT 67.995 172.595 68.285 172.640 ;
        RECT 70.215 172.780 70.535 172.840 ;
        RECT 72.605 172.780 72.745 172.920 ;
        RECT 70.215 172.640 72.745 172.780 ;
        RECT 64.695 172.580 65.015 172.595 ;
        RECT 70.215 172.580 70.535 172.640 ;
        RECT 33.430 172.300 38.705 172.440 ;
        RECT 38.935 172.440 39.255 172.500 ;
        RECT 39.870 172.440 40.160 172.485 ;
        RECT 38.935 172.300 40.160 172.440 ;
        RECT 33.430 172.255 33.720 172.300 ;
        RECT 38.935 172.240 39.255 172.300 ;
        RECT 39.870 172.255 40.160 172.300 ;
        RECT 43.995 172.240 44.315 172.500 ;
        RECT 55.495 172.440 55.815 172.500 ;
        RECT 58.270 172.440 58.560 172.485 ;
        RECT 55.495 172.300 58.560 172.440 ;
        RECT 55.495 172.240 55.815 172.300 ;
        RECT 58.270 172.255 58.560 172.300 ;
        RECT 60.110 172.440 60.400 172.485 ;
        RECT 62.395 172.440 62.715 172.500 ;
        RECT 60.110 172.300 62.715 172.440 ;
        RECT 60.110 172.255 60.400 172.300 ;
        RECT 62.395 172.240 62.715 172.300 ;
        RECT 64.235 172.440 64.555 172.500 ;
        RECT 73.065 172.440 73.205 172.935 ;
        RECT 74.815 172.920 75.135 172.980 ;
        RECT 75.735 172.920 76.055 172.980 ;
        RECT 79.875 173.120 80.195 173.180 ;
        RECT 80.810 173.120 81.100 173.165 ;
        RECT 84.030 173.120 84.320 173.165 ;
        RECT 79.875 172.980 81.100 173.120 ;
        RECT 79.875 172.920 80.195 172.980 ;
        RECT 80.810 172.935 81.100 172.980 ;
        RECT 83.185 172.980 84.320 173.120 ;
        RECT 77.575 172.780 77.895 172.840 ;
        RECT 82.635 172.780 82.955 172.840 ;
        RECT 83.185 172.780 83.325 172.980 ;
        RECT 84.030 172.935 84.320 172.980 ;
        RECT 84.935 173.120 85.255 173.180 ;
        RECT 88.705 173.165 88.845 173.320 ;
        RECT 86.790 173.120 87.080 173.165 ;
        RECT 84.935 172.980 87.080 173.120 ;
        RECT 84.935 172.920 85.255 172.980 ;
        RECT 86.790 172.935 87.080 172.980 ;
        RECT 87.710 172.935 88.000 173.165 ;
        RECT 88.170 172.935 88.460 173.165 ;
        RECT 88.630 172.935 88.920 173.165 ;
        RECT 87.785 172.780 87.925 172.935 ;
        RECT 77.575 172.640 83.325 172.780 ;
        RECT 83.645 172.640 87.925 172.780 ;
        RECT 77.575 172.580 77.895 172.640 ;
        RECT 82.635 172.580 82.955 172.640 ;
        RECT 83.645 172.500 83.785 172.640 ;
        RECT 64.235 172.300 73.205 172.440 ;
        RECT 81.270 172.440 81.560 172.485 ;
        RECT 81.715 172.440 82.035 172.500 ;
        RECT 81.270 172.300 82.035 172.440 ;
        RECT 64.235 172.240 64.555 172.300 ;
        RECT 81.270 172.255 81.560 172.300 ;
        RECT 81.715 172.240 82.035 172.300 ;
        RECT 83.555 172.240 83.875 172.500 ;
        RECT 85.870 172.440 86.160 172.485 ;
        RECT 86.775 172.440 87.095 172.500 ;
        RECT 85.870 172.300 87.095 172.440 ;
        RECT 85.870 172.255 86.160 172.300 ;
        RECT 86.775 172.240 87.095 172.300 ;
        RECT 87.235 172.440 87.555 172.500 ;
        RECT 88.245 172.440 88.385 172.935 ;
        RECT 89.165 172.780 89.305 173.660 ;
        RECT 93.765 173.660 94.825 173.800 ;
        RECT 96.450 173.800 96.740 173.845 ;
        RECT 105.145 173.800 105.435 173.845 ;
        RECT 107.925 173.800 108.215 173.845 ;
        RECT 109.785 173.800 110.075 173.845 ;
        RECT 96.450 173.660 102.645 173.800 ;
        RECT 93.765 173.505 93.905 173.660 ;
        RECT 96.450 173.615 96.740 173.660 ;
        RECT 93.690 173.275 93.980 173.505 ;
        RECT 94.135 173.460 94.455 173.520 ;
        RECT 97.355 173.460 97.675 173.520 ;
        RECT 94.135 173.320 97.675 173.460 ;
        RECT 94.135 173.260 94.455 173.320 ;
        RECT 97.355 173.260 97.675 173.320 ;
        RECT 97.815 173.260 98.135 173.520 ;
        RECT 102.505 173.460 102.645 173.660 ;
        RECT 105.145 173.660 110.075 173.800 ;
        RECT 105.145 173.615 105.435 173.660 ;
        RECT 107.925 173.615 108.215 173.660 ;
        RECT 109.785 173.615 110.075 173.660 ;
        RECT 108.410 173.460 108.700 173.505 ;
        RECT 102.505 173.320 108.700 173.460 ;
        RECT 108.410 173.275 108.700 173.320 ;
        RECT 109.315 173.460 109.635 173.520 ;
        RECT 110.250 173.460 110.540 173.505 ;
        RECT 109.315 173.320 110.540 173.460 ;
        RECT 135.580 173.430 136.830 174.550 ;
        RECT 135.635 173.420 136.775 173.430 ;
        RECT 109.315 173.260 109.635 173.320 ;
        RECT 110.250 173.275 110.540 173.320 ;
        RECT 94.595 173.120 94.915 173.180 ;
        RECT 98.290 173.120 98.580 173.165 ;
        RECT 94.595 172.980 98.580 173.120 ;
        RECT 94.595 172.920 94.915 172.980 ;
        RECT 98.290 172.935 98.580 172.980 ;
        RECT 105.145 173.120 105.435 173.165 ;
        RECT 105.145 172.980 107.680 173.120 ;
        RECT 105.145 172.935 105.435 172.980 ;
        RECT 98.750 172.780 99.040 172.825 ;
        RECT 89.165 172.640 99.040 172.780 ;
        RECT 98.750 172.595 99.040 172.640 ;
        RECT 103.285 172.780 103.575 172.825 ;
        RECT 105.635 172.780 105.955 172.840 ;
        RECT 107.465 172.825 107.680 172.980 ;
        RECT 106.545 172.780 106.835 172.825 ;
        RECT 103.285 172.640 106.835 172.780 ;
        RECT 103.285 172.595 103.575 172.640 ;
        RECT 105.635 172.580 105.955 172.640 ;
        RECT 106.545 172.595 106.835 172.640 ;
        RECT 107.465 172.780 107.755 172.825 ;
        RECT 109.325 172.780 109.615 172.825 ;
        RECT 107.465 172.640 109.615 172.780 ;
        RECT 107.465 172.595 107.755 172.640 ;
        RECT 109.325 172.595 109.615 172.640 ;
        RECT 87.235 172.300 88.385 172.440 ;
        RECT 97.355 172.440 97.675 172.500 ;
        RECT 101.280 172.440 101.570 172.485 ;
        RECT 101.955 172.440 102.275 172.500 ;
        RECT 97.355 172.300 102.275 172.440 ;
        RECT 87.235 172.240 87.555 172.300 ;
        RECT 97.355 172.240 97.675 172.300 ;
        RECT 101.280 172.255 101.570 172.300 ;
        RECT 101.955 172.240 102.275 172.300 ;
        RECT 133.700 172.190 134.930 172.680 ;
        RECT 18.165 171.620 112.465 172.100 ;
        RECT 133.700 171.930 136.690 172.190 ;
        RECT 138.330 171.930 139.470 223.810 ;
        RECT 26.070 171.420 26.360 171.465 ;
        RECT 26.070 171.280 30.425 171.420 ;
        RECT 26.070 171.235 26.360 171.280 ;
        RECT 28.370 171.080 28.660 171.125 ;
        RECT 28.815 171.080 29.135 171.140 ;
        RECT 28.370 170.940 29.135 171.080 ;
        RECT 30.285 171.080 30.425 171.280 ;
        RECT 35.715 171.220 36.035 171.480 ;
        RECT 39.855 171.420 40.175 171.480 ;
        RECT 43.075 171.420 43.395 171.480 ;
        RECT 39.485 171.280 43.395 171.420 ;
        RECT 30.650 171.080 31.300 171.125 ;
        RECT 34.250 171.080 34.540 171.125 ;
        RECT 30.285 170.940 34.540 171.080 ;
        RECT 28.370 170.895 28.660 170.940 ;
        RECT 28.815 170.880 29.135 170.940 ;
        RECT 30.650 170.895 31.300 170.940 ;
        RECT 33.950 170.895 34.540 170.940 ;
        RECT 20.550 170.740 20.840 170.785 ;
        RECT 21.915 170.740 22.235 170.800 ;
        RECT 20.550 170.600 22.235 170.740 ;
        RECT 20.550 170.555 20.840 170.600 ;
        RECT 21.915 170.540 22.235 170.600 ;
        RECT 22.850 170.740 23.140 170.785 ;
        RECT 23.295 170.740 23.615 170.800 ;
        RECT 22.850 170.600 23.615 170.740 ;
        RECT 22.850 170.555 23.140 170.600 ;
        RECT 23.295 170.540 23.615 170.600 ;
        RECT 26.530 170.555 26.820 170.785 ;
        RECT 27.455 170.740 27.745 170.785 ;
        RECT 29.290 170.740 29.580 170.785 ;
        RECT 32.870 170.740 33.160 170.785 ;
        RECT 27.455 170.600 33.160 170.740 ;
        RECT 27.455 170.555 27.745 170.600 ;
        RECT 29.290 170.555 29.580 170.600 ;
        RECT 32.870 170.555 33.160 170.600 ;
        RECT 33.950 170.580 34.240 170.895 ;
        RECT 21.455 169.520 21.775 169.780 ;
        RECT 23.770 169.720 24.060 169.765 ;
        RECT 26.055 169.720 26.375 169.780 ;
        RECT 23.770 169.580 26.375 169.720 ;
        RECT 26.605 169.720 26.745 170.555 ;
        RECT 36.175 170.540 36.495 170.800 ;
        RECT 38.475 170.740 38.795 170.800 ;
        RECT 39.485 170.785 39.625 171.280 ;
        RECT 39.855 171.220 40.175 171.280 ;
        RECT 43.075 171.220 43.395 171.280 ;
        RECT 43.995 171.420 44.315 171.480 ;
        RECT 44.930 171.420 45.220 171.465 ;
        RECT 43.995 171.280 45.220 171.420 ;
        RECT 43.995 171.220 44.315 171.280 ;
        RECT 44.930 171.235 45.220 171.280 ;
        RECT 51.355 171.220 51.675 171.480 ;
        RECT 51.815 171.420 52.135 171.480 ;
        RECT 52.290 171.420 52.580 171.465 ;
        RECT 51.815 171.280 52.580 171.420 ;
        RECT 51.815 171.220 52.135 171.280 ;
        RECT 52.290 171.235 52.580 171.280 ;
        RECT 52.735 171.420 53.055 171.480 ;
        RECT 55.280 171.420 55.570 171.465 ;
        RECT 57.795 171.420 58.115 171.480 ;
        RECT 52.735 171.280 58.115 171.420 ;
        RECT 52.735 171.220 53.055 171.280 ;
        RECT 55.280 171.235 55.570 171.280 ;
        RECT 57.795 171.220 58.115 171.280 ;
        RECT 58.255 171.420 58.575 171.480 ;
        RECT 70.215 171.420 70.535 171.480 ;
        RECT 58.255 171.280 70.535 171.420 ;
        RECT 58.255 171.220 58.575 171.280 ;
        RECT 70.215 171.220 70.535 171.280 ;
        RECT 70.690 171.420 70.980 171.465 ;
        RECT 77.575 171.420 77.895 171.480 ;
        RECT 70.690 171.280 77.895 171.420 ;
        RECT 70.690 171.235 70.980 171.280 ;
        RECT 77.575 171.220 77.895 171.280 ;
        RECT 79.660 171.420 79.950 171.465 ;
        RECT 83.555 171.420 83.875 171.480 ;
        RECT 79.660 171.280 83.875 171.420 ;
        RECT 79.660 171.235 79.950 171.280 ;
        RECT 83.555 171.220 83.875 171.280 ;
        RECT 105.190 171.420 105.480 171.465 ;
        RECT 105.635 171.420 105.955 171.480 ;
        RECT 105.190 171.280 105.955 171.420 ;
        RECT 105.190 171.235 105.480 171.280 ;
        RECT 105.635 171.220 105.955 171.280 ;
        RECT 57.285 171.080 57.575 171.125 ;
        RECT 59.635 171.080 59.955 171.140 ;
        RECT 81.715 171.125 82.035 171.140 ;
        RECT 60.545 171.080 60.835 171.125 ;
        RECT 39.945 170.940 55.725 171.080 ;
        RECT 39.945 170.785 40.085 170.940 ;
        RECT 55.585 170.800 55.725 170.940 ;
        RECT 57.285 170.940 60.835 171.080 ;
        RECT 57.285 170.895 57.575 170.940 ;
        RECT 59.635 170.880 59.955 170.940 ;
        RECT 60.545 170.895 60.835 170.940 ;
        RECT 61.465 171.080 61.755 171.125 ;
        RECT 63.325 171.080 63.615 171.125 ;
        RECT 81.665 171.080 82.035 171.125 ;
        RECT 84.925 171.080 85.215 171.125 ;
        RECT 61.465 170.940 63.615 171.080 ;
        RECT 61.465 170.895 61.755 170.940 ;
        RECT 63.325 170.895 63.615 170.940 ;
        RECT 73.985 170.940 80.105 171.080 ;
        RECT 38.950 170.740 39.240 170.785 ;
        RECT 38.475 170.600 39.240 170.740 ;
        RECT 38.475 170.540 38.795 170.600 ;
        RECT 38.950 170.555 39.240 170.600 ;
        RECT 39.410 170.555 39.700 170.785 ;
        RECT 39.870 170.555 40.160 170.785 ;
        RECT 40.315 170.740 40.635 170.800 ;
        RECT 40.790 170.740 41.080 170.785 ;
        RECT 42.615 170.740 42.935 170.800 ;
        RECT 40.315 170.600 42.935 170.740 ;
        RECT 40.315 170.540 40.635 170.600 ;
        RECT 40.790 170.555 41.080 170.600 ;
        RECT 42.615 170.540 42.935 170.600 ;
        RECT 43.090 170.555 43.380 170.785 ;
        RECT 45.390 170.740 45.680 170.785 ;
        RECT 45.005 170.600 45.680 170.740 ;
        RECT 26.990 170.400 27.280 170.445 ;
        RECT 30.655 170.400 30.975 170.460 ;
        RECT 26.990 170.260 30.975 170.400 ;
        RECT 26.990 170.215 27.280 170.260 ;
        RECT 30.655 170.200 30.975 170.260 ;
        RECT 32.035 170.400 32.355 170.460 ;
        RECT 37.570 170.400 37.860 170.445 ;
        RECT 43.165 170.400 43.305 170.555 ;
        RECT 32.035 170.260 37.860 170.400 ;
        RECT 32.035 170.200 32.355 170.260 ;
        RECT 37.570 170.215 37.860 170.260 ;
        RECT 40.405 170.260 43.305 170.400 ;
        RECT 27.860 170.060 28.150 170.105 ;
        RECT 29.750 170.060 30.040 170.105 ;
        RECT 32.870 170.060 33.160 170.105 ;
        RECT 40.405 170.060 40.545 170.260 ;
        RECT 43.995 170.200 44.315 170.460 ;
        RECT 27.860 169.920 33.160 170.060 ;
        RECT 27.860 169.875 28.150 169.920 ;
        RECT 29.750 169.875 30.040 169.920 ;
        RECT 32.870 169.875 33.160 169.920 ;
        RECT 36.725 169.920 40.545 170.060 ;
        RECT 40.775 170.060 41.095 170.120 ;
        RECT 45.005 170.060 45.145 170.600 ;
        RECT 45.390 170.555 45.680 170.600 ;
        RECT 45.835 170.740 46.155 170.800 ;
        RECT 53.210 170.740 53.500 170.785 ;
        RECT 45.835 170.600 53.500 170.740 ;
        RECT 45.835 170.540 46.155 170.600 ;
        RECT 53.210 170.555 53.500 170.600 ;
        RECT 53.655 170.740 53.975 170.800 ;
        RECT 54.590 170.740 54.880 170.785 ;
        RECT 55.035 170.740 55.355 170.800 ;
        RECT 53.655 170.600 55.355 170.740 ;
        RECT 48.150 170.215 48.440 170.445 ;
        RECT 53.285 170.400 53.425 170.555 ;
        RECT 53.655 170.540 53.975 170.600 ;
        RECT 54.590 170.555 54.880 170.600 ;
        RECT 55.035 170.540 55.355 170.600 ;
        RECT 55.495 170.540 55.815 170.800 ;
        RECT 59.145 170.740 59.435 170.785 ;
        RECT 61.465 170.740 61.680 170.895 ;
        RECT 59.145 170.600 61.680 170.740 ;
        RECT 59.145 170.555 59.435 170.600 ;
        RECT 62.395 170.540 62.715 170.800 ;
        RECT 67.915 170.740 68.235 170.800 ;
        RECT 73.985 170.785 74.125 170.940 ;
        RECT 79.965 170.800 80.105 170.940 ;
        RECT 81.665 170.940 85.215 171.080 ;
        RECT 81.665 170.895 82.035 170.940 ;
        RECT 84.925 170.895 85.215 170.940 ;
        RECT 85.845 171.080 86.135 171.125 ;
        RECT 87.705 171.080 87.995 171.125 ;
        RECT 85.845 170.940 87.995 171.080 ;
        RECT 85.845 170.895 86.135 170.940 ;
        RECT 87.705 170.895 87.995 170.940 ;
        RECT 81.715 170.880 82.035 170.895 ;
        RECT 71.150 170.740 71.440 170.785 ;
        RECT 67.915 170.600 71.440 170.740 ;
        RECT 67.915 170.540 68.235 170.600 ;
        RECT 71.150 170.555 71.440 170.600 ;
        RECT 73.910 170.555 74.200 170.785 ;
        RECT 74.355 170.540 74.675 170.800 ;
        RECT 78.955 170.540 79.275 170.800 ;
        RECT 79.875 170.540 80.195 170.800 ;
        RECT 83.525 170.740 83.815 170.785 ;
        RECT 85.845 170.740 86.060 170.895 ;
        RECT 83.525 170.600 86.060 170.740 ;
        RECT 83.525 170.555 83.815 170.600 ;
        RECT 86.775 170.540 87.095 170.800 ;
        RECT 89.535 170.540 89.855 170.800 ;
        RECT 101.035 170.740 101.355 170.800 ;
        RECT 105.650 170.740 105.940 170.785 ;
        RECT 106.095 170.740 106.415 170.800 ;
        RECT 101.035 170.600 106.415 170.740 ;
        RECT 101.035 170.540 101.355 170.600 ;
        RECT 105.650 170.555 105.940 170.600 ;
        RECT 106.095 170.540 106.415 170.600 ;
        RECT 133.700 170.790 139.470 171.930 ;
        RECT 133.700 170.600 136.690 170.790 ;
        RECT 58.715 170.400 59.035 170.460 ;
        RECT 61.015 170.400 61.335 170.460 ;
        RECT 64.250 170.400 64.540 170.445 ;
        RECT 53.285 170.260 55.725 170.400 ;
        RECT 40.775 169.920 45.145 170.060 ;
        RECT 47.230 170.060 47.520 170.105 ;
        RECT 48.225 170.060 48.365 170.215 ;
        RECT 47.230 169.920 48.365 170.060 ;
        RECT 31.575 169.720 31.895 169.780 ;
        RECT 36.725 169.720 36.865 169.920 ;
        RECT 40.775 169.860 41.095 169.920 ;
        RECT 47.230 169.875 47.520 169.920 ;
        RECT 26.605 169.580 36.865 169.720 ;
        RECT 23.770 169.535 24.060 169.580 ;
        RECT 26.055 169.520 26.375 169.580 ;
        RECT 31.575 169.520 31.895 169.580 ;
        RECT 37.095 169.520 37.415 169.780 ;
        RECT 38.015 169.720 38.335 169.780 ;
        RECT 40.315 169.720 40.635 169.780 ;
        RECT 38.015 169.580 40.635 169.720 ;
        RECT 38.015 169.520 38.335 169.580 ;
        RECT 40.315 169.520 40.635 169.580 ;
        RECT 42.630 169.720 42.920 169.765 ;
        RECT 43.075 169.720 43.395 169.780 ;
        RECT 42.630 169.580 43.395 169.720 ;
        RECT 42.630 169.535 42.920 169.580 ;
        RECT 43.075 169.520 43.395 169.580 ;
        RECT 43.535 169.720 43.855 169.780 ;
        RECT 51.815 169.720 52.135 169.780 ;
        RECT 43.535 169.580 52.135 169.720 ;
        RECT 43.535 169.520 43.855 169.580 ;
        RECT 51.815 169.520 52.135 169.580 ;
        RECT 54.130 169.720 54.420 169.765 ;
        RECT 55.035 169.720 55.355 169.780 ;
        RECT 54.130 169.580 55.355 169.720 ;
        RECT 55.585 169.720 55.725 170.260 ;
        RECT 58.715 170.260 64.540 170.400 ;
        RECT 58.715 170.200 59.035 170.260 ;
        RECT 61.015 170.200 61.335 170.260 ;
        RECT 64.250 170.215 64.540 170.260 ;
        RECT 66.995 170.400 67.315 170.460 ;
        RECT 69.770 170.400 70.060 170.445 ;
        RECT 88.630 170.400 88.920 170.445 ;
        RECT 66.995 170.260 70.060 170.400 ;
        RECT 66.995 170.200 67.315 170.260 ;
        RECT 69.770 170.215 70.060 170.260 ;
        RECT 73.985 170.260 88.920 170.400 ;
        RECT 59.145 170.060 59.435 170.105 ;
        RECT 61.925 170.060 62.215 170.105 ;
        RECT 63.785 170.060 64.075 170.105 ;
        RECT 59.145 169.920 64.075 170.060 ;
        RECT 69.845 170.060 69.985 170.215 ;
        RECT 73.985 170.120 74.125 170.260 ;
        RECT 88.630 170.215 88.920 170.260 ;
        RECT 94.135 170.200 94.455 170.460 ;
        RECT 133.700 170.120 134.930 170.600 ;
        RECT 69.845 169.920 73.665 170.060 ;
        RECT 59.145 169.875 59.435 169.920 ;
        RECT 61.925 169.875 62.215 169.920 ;
        RECT 63.785 169.875 64.075 169.920 ;
        RECT 63.315 169.720 63.635 169.780 ;
        RECT 55.585 169.580 63.635 169.720 ;
        RECT 54.130 169.535 54.420 169.580 ;
        RECT 55.035 169.520 55.355 169.580 ;
        RECT 63.315 169.520 63.635 169.580 ;
        RECT 71.595 169.720 71.915 169.780 ;
        RECT 72.990 169.720 73.280 169.765 ;
        RECT 71.595 169.580 73.280 169.720 ;
        RECT 73.525 169.720 73.665 169.920 ;
        RECT 73.895 169.860 74.215 170.120 ;
        RECT 82.635 170.060 82.955 170.120 ;
        RECT 74.445 169.920 82.955 170.060 ;
        RECT 74.445 169.720 74.585 169.920 ;
        RECT 82.635 169.860 82.955 169.920 ;
        RECT 83.525 170.060 83.815 170.105 ;
        RECT 86.305 170.060 86.595 170.105 ;
        RECT 88.165 170.060 88.455 170.105 ;
        RECT 83.525 169.920 88.455 170.060 ;
        RECT 83.525 169.875 83.815 169.920 ;
        RECT 86.305 169.875 86.595 169.920 ;
        RECT 88.165 169.875 88.455 169.920 ;
        RECT 73.525 169.580 74.585 169.720 ;
        RECT 74.815 169.720 75.135 169.780 ;
        RECT 78.050 169.720 78.340 169.765 ;
        RECT 74.815 169.580 78.340 169.720 ;
        RECT 71.595 169.520 71.915 169.580 ;
        RECT 72.990 169.535 73.280 169.580 ;
        RECT 74.815 169.520 75.135 169.580 ;
        RECT 78.050 169.535 78.340 169.580 ;
        RECT 78.955 169.720 79.275 169.780 ;
        RECT 81.255 169.720 81.575 169.780 ;
        RECT 85.855 169.720 86.175 169.780 ;
        RECT 78.955 169.580 86.175 169.720 ;
        RECT 78.955 169.520 79.275 169.580 ;
        RECT 81.255 169.520 81.575 169.580 ;
        RECT 85.855 169.520 86.175 169.580 ;
        RECT 92.310 169.720 92.600 169.765 ;
        RECT 93.215 169.720 93.535 169.780 ;
        RECT 92.310 169.580 93.535 169.720 ;
        RECT 92.310 169.535 92.600 169.580 ;
        RECT 93.215 169.520 93.535 169.580 ;
        RECT 96.910 169.720 97.200 169.765 ;
        RECT 97.355 169.720 97.675 169.780 ;
        RECT 96.910 169.580 97.675 169.720 ;
        RECT 96.910 169.535 97.200 169.580 ;
        RECT 97.355 169.520 97.675 169.580 ;
        RECT 17.605 168.900 112.465 169.380 ;
        RECT 26.055 168.700 26.375 168.760 ;
        RECT 38.015 168.700 38.335 168.760 ;
        RECT 26.055 168.560 38.335 168.700 ;
        RECT 26.055 168.500 26.375 168.560 ;
        RECT 38.015 168.500 38.335 168.560 ;
        RECT 59.635 168.700 59.955 168.760 ;
        RECT 61.490 168.700 61.780 168.745 ;
        RECT 75.275 168.700 75.595 168.760 ;
        RECT 59.635 168.560 61.780 168.700 ;
        RECT 59.635 168.500 59.955 168.560 ;
        RECT 61.490 168.515 61.780 168.560 ;
        RECT 65.705 168.560 75.595 168.700 ;
        RECT 23.870 168.360 24.160 168.405 ;
        RECT 26.990 168.360 27.280 168.405 ;
        RECT 28.880 168.360 29.170 168.405 ;
        RECT 33.415 168.360 33.735 168.420 ;
        RECT 23.870 168.220 29.170 168.360 ;
        RECT 23.870 168.175 24.160 168.220 ;
        RECT 26.990 168.175 27.280 168.220 ;
        RECT 28.880 168.175 29.170 168.220 ;
        RECT 29.365 168.220 33.735 168.360 ;
        RECT 26.515 168.020 26.835 168.080 ;
        RECT 29.365 168.020 29.505 168.220 ;
        RECT 33.415 168.160 33.735 168.220 ;
        RECT 26.515 167.880 29.505 168.020 ;
        RECT 29.750 168.020 30.040 168.065 ;
        RECT 30.655 168.020 30.975 168.080 ;
        RECT 29.750 167.880 30.975 168.020 ;
        RECT 26.515 167.820 26.835 167.880 ;
        RECT 29.750 167.835 30.040 167.880 ;
        RECT 30.655 167.820 30.975 167.880 ;
        RECT 31.590 167.835 31.880 168.065 ;
        RECT 32.050 168.020 32.340 168.065 ;
        RECT 35.715 168.020 36.035 168.080 ;
        RECT 32.050 167.880 36.035 168.020 ;
        RECT 32.050 167.835 32.340 167.880 ;
        RECT 22.835 167.700 23.155 167.740 ;
        RECT 22.790 167.480 23.155 167.700 ;
        RECT 23.870 167.680 24.160 167.725 ;
        RECT 27.450 167.680 27.740 167.725 ;
        RECT 29.285 167.680 29.575 167.725 ;
        RECT 23.870 167.540 29.575 167.680 ;
        RECT 31.665 167.680 31.805 167.835 ;
        RECT 35.715 167.820 36.035 167.880 ;
        RECT 37.110 168.020 37.400 168.065 ;
        RECT 40.315 168.020 40.635 168.080 ;
        RECT 42.170 168.020 42.460 168.065 ;
        RECT 43.535 168.020 43.855 168.080 ;
        RECT 45.835 168.020 46.155 168.080 ;
        RECT 37.110 167.880 41.005 168.020 ;
        RECT 37.110 167.835 37.400 167.880 ;
        RECT 40.315 167.820 40.635 167.880 ;
        RECT 31.665 167.540 35.945 167.680 ;
        RECT 23.870 167.495 24.160 167.540 ;
        RECT 27.450 167.495 27.740 167.540 ;
        RECT 29.285 167.495 29.575 167.540 ;
        RECT 19.615 167.140 19.935 167.400 ;
        RECT 22.790 167.385 23.080 167.480 ;
        RECT 35.805 167.400 35.945 167.540 ;
        RECT 36.190 167.495 36.480 167.725 ;
        RECT 38.030 167.495 38.320 167.725 ;
        RECT 40.865 167.680 41.005 167.880 ;
        RECT 42.170 167.880 46.155 168.020 ;
        RECT 42.170 167.835 42.460 167.880 ;
        RECT 43.535 167.820 43.855 167.880 ;
        RECT 45.835 167.820 46.155 167.880 ;
        RECT 55.495 168.020 55.815 168.080 ;
        RECT 58.270 168.020 58.560 168.065 ;
        RECT 55.495 167.880 58.560 168.020 ;
        RECT 55.495 167.820 55.815 167.880 ;
        RECT 58.270 167.835 58.560 167.880 ;
        RECT 59.190 168.020 59.480 168.065 ;
        RECT 60.095 168.020 60.415 168.080 ;
        RECT 65.705 168.020 65.845 168.560 ;
        RECT 75.275 168.500 75.595 168.560 ;
        RECT 77.575 168.700 77.895 168.760 ;
        RECT 78.740 168.700 79.030 168.745 ;
        RECT 77.575 168.560 79.030 168.700 ;
        RECT 77.575 168.500 77.895 168.560 ;
        RECT 78.740 168.515 79.030 168.560 ;
        RECT 86.315 168.700 86.635 168.760 ;
        RECT 86.790 168.700 87.080 168.745 ;
        RECT 86.315 168.560 87.080 168.700 ;
        RECT 86.315 168.500 86.635 168.560 ;
        RECT 86.790 168.515 87.080 168.560 ;
        RECT 87.710 168.515 88.000 168.745 ;
        RECT 91.375 168.700 91.695 168.760 ;
        RECT 94.135 168.700 94.455 168.760 ;
        RECT 96.910 168.700 97.200 168.745 ;
        RECT 91.375 168.560 92.985 168.700 ;
        RECT 70.235 168.360 70.525 168.405 ;
        RECT 72.095 168.360 72.385 168.405 ;
        RECT 74.875 168.360 75.165 168.405 ;
        RECT 70.235 168.220 75.165 168.360 ;
        RECT 70.235 168.175 70.525 168.220 ;
        RECT 72.095 168.175 72.385 168.220 ;
        RECT 74.875 168.175 75.165 168.220 ;
        RECT 81.730 168.360 82.020 168.405 ;
        RECT 87.785 168.360 87.925 168.515 ;
        RECT 91.375 168.500 91.695 168.560 ;
        RECT 81.730 168.220 87.925 168.360 ;
        RECT 90.915 168.360 91.235 168.420 ;
        RECT 90.915 168.220 92.525 168.360 ;
        RECT 81.730 168.175 82.020 168.220 ;
        RECT 90.915 168.160 91.235 168.220 ;
        RECT 59.190 167.880 60.415 168.020 ;
        RECT 59.190 167.835 59.480 167.880 ;
        RECT 60.095 167.820 60.415 167.880 ;
        RECT 65.245 167.880 65.845 168.020 ;
        RECT 66.550 168.020 66.840 168.065 ;
        RECT 66.995 168.020 67.315 168.080 ;
        RECT 66.550 167.880 67.315 168.020 ;
        RECT 43.090 167.680 43.380 167.725 ;
        RECT 44.455 167.680 44.775 167.740 ;
        RECT 40.865 167.540 44.775 167.680 ;
        RECT 43.090 167.495 43.380 167.540 ;
        RECT 22.490 167.340 23.080 167.385 ;
        RECT 25.730 167.340 26.380 167.385 ;
        RECT 22.490 167.200 26.380 167.340 ;
        RECT 22.490 167.155 22.780 167.200 ;
        RECT 25.730 167.155 26.380 167.200 ;
        RECT 28.355 167.140 28.675 167.400 ;
        RECT 35.715 167.140 36.035 167.400 ;
        RECT 36.265 167.340 36.405 167.495 ;
        RECT 37.095 167.340 37.415 167.400 ;
        RECT 36.265 167.200 37.415 167.340 ;
        RECT 38.105 167.340 38.245 167.495 ;
        RECT 44.455 167.480 44.775 167.540 ;
        RECT 46.310 167.680 46.600 167.725 ;
        RECT 49.055 167.680 49.375 167.740 ;
        RECT 57.810 167.680 58.100 167.725 ;
        RECT 46.310 167.540 49.375 167.680 ;
        RECT 46.310 167.495 46.600 167.540 ;
        RECT 49.055 167.480 49.375 167.540 ;
        RECT 53.055 167.540 58.100 167.680 ;
        RECT 42.155 167.340 42.475 167.400 ;
        RECT 38.105 167.200 42.475 167.340 ;
        RECT 37.095 167.140 37.415 167.200 ;
        RECT 42.155 167.140 42.475 167.200 ;
        RECT 46.755 167.140 47.075 167.400 ;
        RECT 48.135 167.340 48.455 167.400 ;
        RECT 53.055 167.340 53.195 167.540 ;
        RECT 57.810 167.495 58.100 167.540 ;
        RECT 61.935 167.480 62.255 167.740 ;
        RECT 65.245 167.725 65.385 167.880 ;
        RECT 66.550 167.835 66.840 167.880 ;
        RECT 66.995 167.820 67.315 167.880 ;
        RECT 71.595 167.820 71.915 168.080 ;
        RECT 73.895 168.020 74.215 168.080 ;
        RECT 72.145 167.880 74.215 168.020 ;
        RECT 65.170 167.495 65.460 167.725 ;
        RECT 67.470 167.680 67.760 167.725 ;
        RECT 65.705 167.540 67.760 167.680 ;
        RECT 48.135 167.200 53.195 167.340 ;
        RECT 55.510 167.340 55.800 167.385 ;
        RECT 58.715 167.340 59.035 167.400 ;
        RECT 55.510 167.200 59.035 167.340 ;
        RECT 48.135 167.140 48.455 167.200 ;
        RECT 55.510 167.155 55.800 167.200 ;
        RECT 58.715 167.140 59.035 167.200 ;
        RECT 59.175 167.340 59.495 167.400 ;
        RECT 65.705 167.340 65.845 167.540 ;
        RECT 67.470 167.495 67.760 167.540 ;
        RECT 69.770 167.680 70.060 167.725 ;
        RECT 72.145 167.680 72.285 167.880 ;
        RECT 73.895 167.820 74.215 167.880 ;
        RECT 82.635 167.820 82.955 168.080 ;
        RECT 86.315 168.020 86.635 168.080 ;
        RECT 83.185 167.880 86.635 168.020 ;
        RECT 74.875 167.680 75.165 167.725 ;
        RECT 69.770 167.540 72.285 167.680 ;
        RECT 72.630 167.540 75.165 167.680 ;
        RECT 69.770 167.495 70.060 167.540 ;
        RECT 59.175 167.200 65.845 167.340 ;
        RECT 67.010 167.340 67.300 167.385 ;
        RECT 67.915 167.340 68.235 167.400 ;
        RECT 72.630 167.385 72.845 167.540 ;
        RECT 74.875 167.495 75.165 167.540 ;
        RECT 80.350 167.495 80.640 167.725 ;
        RECT 80.810 167.680 81.100 167.725 ;
        RECT 82.175 167.680 82.495 167.740 ;
        RECT 83.185 167.680 83.325 167.880 ;
        RECT 86.315 167.820 86.635 167.880 ;
        RECT 88.615 167.820 88.935 168.080 ;
        RECT 90.455 168.020 90.775 168.080 ;
        RECT 90.455 167.880 91.605 168.020 ;
        RECT 90.455 167.820 90.775 167.880 ;
        RECT 80.810 167.540 83.325 167.680 ;
        RECT 83.555 167.680 83.875 167.740 ;
        RECT 84.030 167.680 84.320 167.725 ;
        RECT 83.555 167.540 84.320 167.680 ;
        RECT 80.810 167.495 81.100 167.540 ;
        RECT 67.010 167.200 68.235 167.340 ;
        RECT 59.175 167.140 59.495 167.200 ;
        RECT 67.010 167.155 67.300 167.200 ;
        RECT 67.915 167.140 68.235 167.200 ;
        RECT 70.695 167.340 70.985 167.385 ;
        RECT 72.555 167.340 72.845 167.385 ;
        RECT 70.695 167.200 72.845 167.340 ;
        RECT 70.695 167.155 70.985 167.200 ;
        RECT 72.555 167.155 72.845 167.200 ;
        RECT 73.475 167.340 73.765 167.385 ;
        RECT 74.355 167.340 74.675 167.400 ;
        RECT 76.735 167.340 77.025 167.385 ;
        RECT 73.475 167.200 77.025 167.340 ;
        RECT 80.425 167.340 80.565 167.495 ;
        RECT 82.175 167.480 82.495 167.540 ;
        RECT 83.555 167.480 83.875 167.540 ;
        RECT 84.030 167.495 84.320 167.540 ;
        RECT 86.775 167.680 87.095 167.740 ;
        RECT 87.710 167.680 88.000 167.725 ;
        RECT 86.775 167.540 88.000 167.680 ;
        RECT 86.775 167.480 87.095 167.540 ;
        RECT 87.710 167.495 88.000 167.540 ;
        RECT 89.995 167.680 90.315 167.740 ;
        RECT 91.465 167.725 91.605 167.880 ;
        RECT 90.930 167.680 91.220 167.725 ;
        RECT 89.995 167.540 91.220 167.680 ;
        RECT 89.995 167.480 90.315 167.540 ;
        RECT 90.930 167.495 91.220 167.540 ;
        RECT 91.390 167.495 91.680 167.725 ;
        RECT 91.850 167.495 92.140 167.725 ;
        RECT 92.385 167.680 92.525 168.220 ;
        RECT 92.845 168.020 92.985 168.560 ;
        RECT 94.135 168.560 97.200 168.700 ;
        RECT 94.135 168.500 94.455 168.560 ;
        RECT 96.910 168.515 97.200 168.560 ;
        RECT 93.675 168.020 93.995 168.080 ;
        RECT 92.845 167.880 93.995 168.020 ;
        RECT 93.675 167.820 93.995 167.880 ;
        RECT 98.275 168.020 98.595 168.080 ;
        RECT 100.590 168.020 100.880 168.065 ;
        RECT 98.275 167.880 100.880 168.020 ;
        RECT 98.275 167.820 98.595 167.880 ;
        RECT 100.590 167.835 100.880 167.880 ;
        RECT 92.770 167.680 93.060 167.725 ;
        RECT 92.385 167.540 93.060 167.680 ;
        RECT 92.770 167.495 93.060 167.540 ;
        RECT 93.215 167.680 93.535 167.740 ;
        RECT 95.070 167.680 95.360 167.725 ;
        RECT 93.215 167.540 95.360 167.680 ;
        RECT 84.935 167.340 85.255 167.400 ;
        RECT 80.425 167.200 85.255 167.340 ;
        RECT 73.475 167.155 73.765 167.200 ;
        RECT 74.355 167.140 74.675 167.200 ;
        RECT 76.735 167.155 77.025 167.200 ;
        RECT 84.935 167.140 85.255 167.200 ;
        RECT 89.090 167.340 89.380 167.385 ;
        RECT 89.550 167.340 89.840 167.385 ;
        RECT 89.090 167.200 89.840 167.340 ;
        RECT 91.925 167.340 92.065 167.495 ;
        RECT 93.215 167.480 93.535 167.540 ;
        RECT 95.070 167.495 95.360 167.540 ;
        RECT 101.955 167.480 102.275 167.740 ;
        RECT 105.650 167.680 105.940 167.725 ;
        RECT 106.095 167.680 106.415 167.740 ;
        RECT 105.650 167.540 106.415 167.680 ;
        RECT 105.650 167.495 105.940 167.540 ;
        RECT 106.095 167.480 106.415 167.540 ;
        RECT 97.815 167.340 98.135 167.400 ;
        RECT 101.510 167.340 101.800 167.385 ;
        RECT 91.925 167.200 101.800 167.340 ;
        RECT 89.090 167.155 89.380 167.200 ;
        RECT 89.550 167.155 89.840 167.200 ;
        RECT 97.815 167.140 98.135 167.200 ;
        RECT 101.510 167.155 101.800 167.200 ;
        RECT 32.510 167.000 32.800 167.045 ;
        RECT 33.415 167.000 33.735 167.060 ;
        RECT 32.510 166.860 33.735 167.000 ;
        RECT 32.510 166.815 32.800 166.860 ;
        RECT 33.415 166.800 33.735 166.860 ;
        RECT 34.335 166.800 34.655 167.060 ;
        RECT 35.255 166.800 35.575 167.060 ;
        RECT 40.775 166.800 41.095 167.060 ;
        RECT 42.615 166.800 42.935 167.060 ;
        RECT 44.915 166.800 45.235 167.060 ;
        RECT 45.375 167.000 45.695 167.060 ;
        RECT 45.850 167.000 46.140 167.045 ;
        RECT 45.375 166.860 46.140 167.000 ;
        RECT 45.375 166.800 45.695 166.860 ;
        RECT 45.850 166.815 46.140 166.860 ;
        RECT 55.970 167.000 56.260 167.045 ;
        RECT 56.875 167.000 57.195 167.060 ;
        RECT 55.970 166.860 57.195 167.000 ;
        RECT 55.970 166.815 56.260 166.860 ;
        RECT 56.875 166.800 57.195 166.860 ;
        RECT 64.695 166.800 65.015 167.060 ;
        RECT 67.455 167.000 67.775 167.060 ;
        RECT 69.310 167.000 69.600 167.045 ;
        RECT 67.455 166.860 69.600 167.000 ;
        RECT 67.455 166.800 67.775 166.860 ;
        RECT 69.310 166.815 69.600 166.860 ;
        RECT 83.570 167.000 83.860 167.045 ;
        RECT 84.475 167.000 84.795 167.060 ;
        RECT 83.570 166.860 84.795 167.000 ;
        RECT 83.570 166.815 83.860 166.860 ;
        RECT 84.475 166.800 84.795 166.860 ;
        RECT 85.855 166.800 86.175 167.060 ;
        RECT 89.995 167.000 90.315 167.060 ;
        RECT 94.610 167.000 94.900 167.045 ;
        RECT 89.995 166.860 94.900 167.000 ;
        RECT 89.995 166.800 90.315 166.860 ;
        RECT 94.610 166.815 94.900 166.860 ;
        RECT 103.795 166.800 104.115 167.060 ;
        RECT 105.190 167.000 105.480 167.045 ;
        RECT 105.635 167.000 105.955 167.060 ;
        RECT 105.190 166.860 105.955 167.000 ;
        RECT 105.190 166.815 105.480 166.860 ;
        RECT 105.635 166.800 105.955 166.860 ;
        RECT 18.165 166.180 112.465 166.660 ;
        RECT 23.755 165.780 24.075 166.040 ;
        RECT 26.515 165.780 26.835 166.040 ;
        RECT 27.450 165.980 27.740 166.025 ;
        RECT 28.355 165.980 28.675 166.040 ;
        RECT 27.450 165.840 28.675 165.980 ;
        RECT 27.450 165.795 27.740 165.840 ;
        RECT 28.355 165.780 28.675 165.840 ;
        RECT 28.815 165.980 29.135 166.040 ;
        RECT 30.210 165.980 30.500 166.025 ;
        RECT 32.035 165.980 32.355 166.040 ;
        RECT 28.815 165.840 30.500 165.980 ;
        RECT 28.815 165.780 29.135 165.840 ;
        RECT 30.210 165.795 30.500 165.840 ;
        RECT 30.745 165.840 32.355 165.980 ;
        RECT 20.535 165.440 20.855 165.700 ;
        RECT 21.470 165.640 21.760 165.685 ;
        RECT 23.295 165.640 23.615 165.700 ;
        RECT 21.470 165.500 23.615 165.640 ;
        RECT 21.470 165.455 21.760 165.500 ;
        RECT 23.295 165.440 23.615 165.500 ;
        RECT 24.215 165.640 24.535 165.700 ;
        RECT 25.150 165.640 25.440 165.685 ;
        RECT 24.215 165.500 25.440 165.640 ;
        RECT 24.215 165.440 24.535 165.500 ;
        RECT 25.150 165.455 25.440 165.500 ;
        RECT 29.750 165.640 30.040 165.685 ;
        RECT 30.745 165.640 30.885 165.840 ;
        RECT 32.035 165.780 32.355 165.840 ;
        RECT 32.955 165.980 33.275 166.040 ;
        RECT 36.175 165.980 36.495 166.040 ;
        RECT 32.955 165.840 36.495 165.980 ;
        RECT 32.955 165.780 33.275 165.840 ;
        RECT 33.890 165.640 34.180 165.685 ;
        RECT 29.750 165.500 30.885 165.640 ;
        RECT 31.205 165.500 34.180 165.640 ;
        RECT 35.345 165.640 35.485 165.840 ;
        RECT 36.175 165.780 36.495 165.840 ;
        RECT 37.800 165.980 38.090 166.025 ;
        RECT 40.315 165.980 40.635 166.040 ;
        RECT 37.800 165.840 40.635 165.980 ;
        RECT 37.800 165.795 38.090 165.840 ;
        RECT 40.315 165.780 40.635 165.840 ;
        RECT 49.760 165.980 50.050 166.025 ;
        RECT 55.495 165.980 55.815 166.040 ;
        RECT 49.760 165.840 55.815 165.980 ;
        RECT 49.760 165.795 50.050 165.840 ;
        RECT 55.495 165.780 55.815 165.840 ;
        RECT 64.235 165.780 64.555 166.040 ;
        RECT 89.995 165.780 90.315 166.040 ;
        RECT 106.095 165.980 106.415 166.040 ;
        RECT 91.005 165.840 106.415 165.980 ;
        RECT 43.075 165.685 43.395 165.700 ;
        RECT 55.035 165.685 55.355 165.700 ;
        RECT 39.805 165.640 40.095 165.685 ;
        RECT 43.065 165.640 43.395 165.685 ;
        RECT 35.345 165.500 35.945 165.640 ;
        RECT 29.750 165.455 30.040 165.500 ;
        RECT 22.850 165.300 23.140 165.345 ;
        RECT 24.675 165.300 24.995 165.360 ;
        RECT 22.850 165.160 24.995 165.300 ;
        RECT 22.850 165.115 23.140 165.160 ;
        RECT 24.675 165.100 24.995 165.160 ;
        RECT 28.370 165.300 28.660 165.345 ;
        RECT 31.205 165.300 31.345 165.500 ;
        RECT 33.890 165.455 34.180 165.500 ;
        RECT 28.370 165.160 31.345 165.300 ;
        RECT 33.430 165.300 33.720 165.345 ;
        RECT 34.335 165.300 34.655 165.360 ;
        RECT 33.430 165.160 34.655 165.300 ;
        RECT 28.370 165.115 28.660 165.160 ;
        RECT 33.430 165.115 33.720 165.160 ;
        RECT 34.335 165.100 34.655 165.160 ;
        RECT 34.795 165.300 35.115 165.360 ;
        RECT 35.805 165.345 35.945 165.500 ;
        RECT 39.805 165.500 43.395 165.640 ;
        RECT 39.805 165.455 40.095 165.500 ;
        RECT 43.065 165.455 43.395 165.500 ;
        RECT 43.075 165.440 43.395 165.455 ;
        RECT 43.985 165.640 44.275 165.685 ;
        RECT 45.845 165.640 46.135 165.685 ;
        RECT 43.985 165.500 46.135 165.640 ;
        RECT 43.985 165.455 44.275 165.500 ;
        RECT 45.845 165.455 46.135 165.500 ;
        RECT 51.765 165.640 52.055 165.685 ;
        RECT 55.025 165.640 55.355 165.685 ;
        RECT 51.765 165.500 55.355 165.640 ;
        RECT 51.765 165.455 52.055 165.500 ;
        RECT 55.025 165.455 55.355 165.500 ;
        RECT 35.270 165.300 35.560 165.345 ;
        RECT 34.795 165.160 35.560 165.300 ;
        RECT 34.795 165.100 35.115 165.160 ;
        RECT 35.270 165.115 35.560 165.160 ;
        RECT 35.730 165.115 36.020 165.345 ;
        RECT 36.190 165.115 36.480 165.345 ;
        RECT 37.110 165.300 37.400 165.345 ;
        RECT 38.015 165.300 38.335 165.360 ;
        RECT 37.110 165.160 38.335 165.300 ;
        RECT 37.110 165.115 37.400 165.160 ;
        RECT 29.290 164.775 29.580 165.005 ;
        RECT 29.735 164.960 30.055 165.020 ;
        RECT 36.265 164.960 36.405 165.115 ;
        RECT 38.015 165.100 38.335 165.160 ;
        RECT 41.665 165.300 41.955 165.345 ;
        RECT 43.985 165.300 44.200 165.455 ;
        RECT 55.035 165.440 55.355 165.455 ;
        RECT 55.945 165.640 56.235 165.685 ;
        RECT 57.805 165.640 58.095 165.685 ;
        RECT 55.945 165.500 58.095 165.640 ;
        RECT 55.945 165.455 56.235 165.500 ;
        RECT 57.805 165.455 58.095 165.500 ;
        RECT 41.665 165.160 44.200 165.300 ;
        RECT 41.665 165.115 41.955 165.160 ;
        RECT 44.915 165.100 45.235 165.360 ;
        RECT 46.770 165.115 47.060 165.345 ;
        RECT 48.150 165.300 48.440 165.345 ;
        RECT 48.595 165.300 48.915 165.360 ;
        RECT 52.735 165.300 53.055 165.360 ;
        RECT 48.150 165.160 53.055 165.300 ;
        RECT 48.150 165.115 48.440 165.160 ;
        RECT 29.735 164.820 36.405 164.960 ;
        RECT 36.635 164.960 36.955 165.020 ;
        RECT 46.845 164.960 46.985 165.115 ;
        RECT 48.595 165.100 48.915 165.160 ;
        RECT 52.735 165.100 53.055 165.160 ;
        RECT 53.625 165.300 53.915 165.345 ;
        RECT 55.945 165.300 56.160 165.455 ;
        RECT 53.625 165.160 56.160 165.300 ;
        RECT 53.625 165.115 53.915 165.160 ;
        RECT 56.875 165.100 57.195 165.360 ;
        RECT 61.030 165.300 61.320 165.345 ;
        RECT 64.325 165.300 64.465 165.780 ;
        RECT 64.695 165.640 65.015 165.700 ;
        RECT 65.730 165.640 66.020 165.685 ;
        RECT 68.970 165.640 69.620 165.685 ;
        RECT 78.050 165.640 78.340 165.685 ;
        RECT 64.695 165.500 69.620 165.640 ;
        RECT 64.695 165.440 65.015 165.500 ;
        RECT 65.730 165.455 66.320 165.500 ;
        RECT 68.970 165.455 69.620 165.500 ;
        RECT 73.985 165.500 78.340 165.640 ;
        RECT 61.030 165.160 64.465 165.300 ;
        RECT 61.030 165.115 61.320 165.160 ;
        RECT 66.030 165.140 66.320 165.455 ;
        RECT 73.985 165.360 74.125 165.500 ;
        RECT 78.050 165.455 78.340 165.500 ;
        RECT 81.205 165.640 81.495 165.685 ;
        RECT 84.465 165.640 84.755 165.685 ;
        RECT 81.205 165.500 84.755 165.640 ;
        RECT 81.205 165.455 81.495 165.500 ;
        RECT 84.465 165.455 84.755 165.500 ;
        RECT 85.385 165.640 85.675 165.685 ;
        RECT 87.245 165.640 87.535 165.685 ;
        RECT 85.385 165.500 87.535 165.640 ;
        RECT 85.385 165.455 85.675 165.500 ;
        RECT 87.245 165.455 87.535 165.500 ;
        RECT 67.110 165.300 67.400 165.345 ;
        RECT 70.690 165.300 70.980 165.345 ;
        RECT 72.525 165.300 72.815 165.345 ;
        RECT 67.110 165.160 72.815 165.300 ;
        RECT 67.110 165.115 67.400 165.160 ;
        RECT 70.690 165.115 70.980 165.160 ;
        RECT 72.525 165.115 72.815 165.160 ;
        RECT 72.990 165.300 73.280 165.345 ;
        RECT 73.895 165.300 74.215 165.360 ;
        RECT 72.990 165.160 74.215 165.300 ;
        RECT 72.990 165.115 73.280 165.160 ;
        RECT 73.895 165.100 74.215 165.160 ;
        RECT 74.815 165.100 75.135 165.360 ;
        RECT 75.290 165.300 75.580 165.345 ;
        RECT 81.345 165.300 81.485 165.455 ;
        RECT 75.290 165.160 81.485 165.300 ;
        RECT 83.065 165.300 83.355 165.345 ;
        RECT 85.385 165.300 85.600 165.455 ;
        RECT 83.065 165.160 85.600 165.300 ;
        RECT 85.855 165.300 86.175 165.360 ;
        RECT 86.330 165.300 86.620 165.345 ;
        RECT 85.855 165.160 86.620 165.300 ;
        RECT 75.290 165.115 75.580 165.160 ;
        RECT 83.065 165.115 83.355 165.160 ;
        RECT 85.855 165.100 86.175 165.160 ;
        RECT 86.330 165.115 86.620 165.160 ;
        RECT 89.550 165.300 89.840 165.345 ;
        RECT 91.005 165.300 91.145 165.840 ;
        RECT 106.095 165.780 106.415 165.840 ;
        RECT 91.490 165.640 91.780 165.685 ;
        RECT 94.730 165.640 95.380 165.685 ;
        RECT 91.490 165.500 95.380 165.640 ;
        RECT 91.490 165.455 92.080 165.500 ;
        RECT 94.730 165.455 95.380 165.500 ;
        RECT 89.550 165.160 91.145 165.300 ;
        RECT 89.550 165.115 89.840 165.160 ;
        RECT 91.790 165.140 92.080 165.455 ;
        RECT 97.355 165.440 97.675 165.700 ;
        RECT 97.815 165.640 98.135 165.700 ;
        RECT 101.280 165.640 101.570 165.685 ;
        RECT 97.815 165.500 101.570 165.640 ;
        RECT 97.815 165.440 98.135 165.500 ;
        RECT 101.280 165.455 101.570 165.500 ;
        RECT 103.285 165.640 103.575 165.685 ;
        RECT 105.635 165.640 105.955 165.700 ;
        RECT 106.545 165.640 106.835 165.685 ;
        RECT 103.285 165.500 106.835 165.640 ;
        RECT 103.285 165.455 103.575 165.500 ;
        RECT 105.635 165.440 105.955 165.500 ;
        RECT 106.545 165.455 106.835 165.500 ;
        RECT 107.465 165.640 107.755 165.685 ;
        RECT 109.325 165.640 109.615 165.685 ;
        RECT 107.465 165.500 109.615 165.640 ;
        RECT 107.465 165.455 107.755 165.500 ;
        RECT 109.325 165.455 109.615 165.500 ;
        RECT 135.580 165.470 136.830 166.590 ;
        RECT 92.870 165.300 93.160 165.345 ;
        RECT 96.450 165.300 96.740 165.345 ;
        RECT 98.285 165.300 98.575 165.345 ;
        RECT 92.870 165.160 98.575 165.300 ;
        RECT 36.635 164.820 46.985 164.960 ;
        RECT 29.365 164.620 29.505 164.775 ;
        RECT 29.735 164.760 30.055 164.820 ;
        RECT 36.635 164.760 36.955 164.820 ;
        RECT 58.715 164.760 59.035 165.020 ;
        RECT 63.790 164.960 64.080 165.005 ;
        RECT 67.915 164.960 68.235 165.020 ;
        RECT 63.790 164.820 68.235 164.960 ;
        RECT 63.790 164.775 64.080 164.820 ;
        RECT 67.915 164.760 68.235 164.820 ;
        RECT 71.595 164.760 71.915 165.020 ;
        RECT 85.395 164.960 85.715 165.020 ;
        RECT 88.170 164.960 88.460 165.005 ;
        RECT 85.395 164.820 88.460 164.960 ;
        RECT 85.395 164.760 85.715 164.820 ;
        RECT 88.170 164.775 88.460 164.820 ;
        RECT 89.090 164.960 89.380 165.005 ;
        RECT 91.925 164.960 92.065 165.140 ;
        RECT 92.870 165.115 93.160 165.160 ;
        RECT 96.450 165.115 96.740 165.160 ;
        RECT 98.285 165.115 98.575 165.160 ;
        RECT 105.145 165.300 105.435 165.345 ;
        RECT 107.465 165.300 107.680 165.455 ;
        RECT 105.145 165.160 107.680 165.300 ;
        RECT 105.145 165.115 105.435 165.160 ;
        RECT 98.750 164.960 99.040 165.005 ;
        RECT 99.195 164.960 99.515 165.020 ;
        RECT 89.090 164.820 92.065 164.960 ;
        RECT 92.385 164.820 99.515 164.960 ;
        RECT 89.090 164.775 89.380 164.820 ;
        RECT 38.935 164.620 39.255 164.680 ;
        RECT 29.365 164.480 39.255 164.620 ;
        RECT 38.935 164.420 39.255 164.480 ;
        RECT 41.665 164.620 41.955 164.665 ;
        RECT 44.445 164.620 44.735 164.665 ;
        RECT 46.305 164.620 46.595 164.665 ;
        RECT 41.665 164.480 46.595 164.620 ;
        RECT 41.665 164.435 41.955 164.480 ;
        RECT 44.445 164.435 44.735 164.480 ;
        RECT 46.305 164.435 46.595 164.480 ;
        RECT 46.755 164.620 47.075 164.680 ;
        RECT 53.625 164.620 53.915 164.665 ;
        RECT 56.405 164.620 56.695 164.665 ;
        RECT 58.265 164.620 58.555 164.665 ;
        RECT 46.755 164.480 53.195 164.620 ;
        RECT 46.755 164.420 47.075 164.480 ;
        RECT 29.750 164.280 30.040 164.325 ;
        RECT 35.255 164.280 35.575 164.340 ;
        RECT 29.750 164.140 35.575 164.280 ;
        RECT 29.750 164.095 30.040 164.140 ;
        RECT 35.255 164.080 35.575 164.140 ;
        RECT 48.610 164.280 48.900 164.325 ;
        RECT 49.515 164.280 49.835 164.340 ;
        RECT 48.610 164.140 49.835 164.280 ;
        RECT 53.055 164.280 53.195 164.480 ;
        RECT 53.625 164.480 58.555 164.620 ;
        RECT 53.625 164.435 53.915 164.480 ;
        RECT 56.405 164.435 56.695 164.480 ;
        RECT 58.265 164.435 58.555 164.480 ;
        RECT 67.110 164.620 67.400 164.665 ;
        RECT 70.230 164.620 70.520 164.665 ;
        RECT 72.120 164.620 72.410 164.665 ;
        RECT 67.110 164.480 72.410 164.620 ;
        RECT 67.110 164.435 67.400 164.480 ;
        RECT 70.230 164.435 70.520 164.480 ;
        RECT 72.120 164.435 72.410 164.480 ;
        RECT 83.065 164.620 83.355 164.665 ;
        RECT 85.845 164.620 86.135 164.665 ;
        RECT 87.705 164.620 87.995 164.665 ;
        RECT 83.065 164.480 87.995 164.620 ;
        RECT 88.245 164.620 88.385 164.775 ;
        RECT 92.385 164.620 92.525 164.820 ;
        RECT 98.750 164.775 99.040 164.820 ;
        RECT 99.195 164.760 99.515 164.820 ;
        RECT 103.795 164.960 104.115 165.020 ;
        RECT 108.410 164.960 108.700 165.005 ;
        RECT 103.795 164.820 108.700 164.960 ;
        RECT 103.795 164.760 104.115 164.820 ;
        RECT 108.410 164.775 108.700 164.820 ;
        RECT 109.315 164.960 109.635 165.020 ;
        RECT 110.250 164.960 110.540 165.005 ;
        RECT 109.315 164.820 110.540 164.960 ;
        RECT 109.315 164.760 109.635 164.820 ;
        RECT 110.250 164.775 110.540 164.820 ;
        RECT 88.245 164.480 92.525 164.620 ;
        RECT 92.870 164.620 93.160 164.665 ;
        RECT 95.990 164.620 96.280 164.665 ;
        RECT 97.880 164.620 98.170 164.665 ;
        RECT 92.870 164.480 98.170 164.620 ;
        RECT 83.065 164.435 83.355 164.480 ;
        RECT 85.845 164.435 86.135 164.480 ;
        RECT 87.705 164.435 87.995 164.480 ;
        RECT 92.870 164.435 93.160 164.480 ;
        RECT 95.990 164.435 96.280 164.480 ;
        RECT 97.880 164.435 98.170 164.480 ;
        RECT 105.145 164.620 105.435 164.665 ;
        RECT 107.925 164.620 108.215 164.665 ;
        RECT 109.785 164.620 110.075 164.665 ;
        RECT 105.145 164.480 110.075 164.620 ;
        RECT 105.145 164.435 105.435 164.480 ;
        RECT 107.925 164.435 108.215 164.480 ;
        RECT 109.785 164.435 110.075 164.480 ;
        RECT 61.015 164.280 61.335 164.340 ;
        RECT 53.055 164.140 61.335 164.280 ;
        RECT 48.610 164.095 48.900 164.140 ;
        RECT 49.515 164.080 49.835 164.140 ;
        RECT 61.015 164.080 61.335 164.140 ;
        RECT 79.200 164.280 79.490 164.325 ;
        RECT 84.475 164.280 84.795 164.340 ;
        RECT 79.200 164.140 84.795 164.280 ;
        RECT 79.200 164.095 79.490 164.140 ;
        RECT 84.475 164.080 84.795 164.140 ;
        RECT 17.605 163.460 112.465 163.940 ;
        RECT 25.610 163.260 25.900 163.305 ;
        RECT 29.735 163.260 30.055 163.320 ;
        RECT 25.610 163.120 30.055 163.260 ;
        RECT 25.610 163.075 25.900 163.120 ;
        RECT 22.390 162.580 22.680 162.625 ;
        RECT 25.685 162.580 25.825 163.075 ;
        RECT 29.735 163.060 30.055 163.120 ;
        RECT 30.655 163.260 30.975 163.320 ;
        RECT 32.495 163.260 32.815 163.320 ;
        RECT 36.635 163.260 36.955 163.320 ;
        RECT 30.655 163.120 36.955 163.260 ;
        RECT 30.655 163.060 30.975 163.120 ;
        RECT 32.495 163.060 32.815 163.120 ;
        RECT 28.470 162.920 28.760 162.965 ;
        RECT 31.590 162.920 31.880 162.965 ;
        RECT 33.480 162.920 33.770 162.965 ;
        RECT 28.470 162.780 33.770 162.920 ;
        RECT 28.470 162.735 28.760 162.780 ;
        RECT 31.590 162.735 31.880 162.780 ;
        RECT 33.480 162.735 33.770 162.780 ;
        RECT 32.955 162.580 33.275 162.640 ;
        RECT 34.425 162.625 34.565 163.120 ;
        RECT 36.635 163.060 36.955 163.120 ;
        RECT 37.095 163.260 37.415 163.320 ;
        RECT 38.935 163.260 39.255 163.320 ;
        RECT 37.095 163.120 39.255 163.260 ;
        RECT 37.095 163.060 37.415 163.120 ;
        RECT 38.935 163.060 39.255 163.120 ;
        RECT 48.135 163.060 48.455 163.320 ;
        RECT 60.095 163.260 60.415 163.320 ;
        RECT 62.395 163.260 62.715 163.320 ;
        RECT 53.285 163.120 62.715 163.260 ;
        RECT 22.390 162.440 25.825 162.580 ;
        RECT 27.065 162.440 33.275 162.580 ;
        RECT 22.390 162.395 22.680 162.440 ;
        RECT 21.470 162.240 21.760 162.285 ;
        RECT 21.915 162.240 22.235 162.300 ;
        RECT 21.470 162.100 22.235 162.240 ;
        RECT 21.470 162.055 21.760 162.100 ;
        RECT 21.915 162.040 22.235 162.100 ;
        RECT 25.150 162.240 25.440 162.285 ;
        RECT 27.065 162.240 27.205 162.440 ;
        RECT 32.955 162.380 33.275 162.440 ;
        RECT 34.350 162.395 34.640 162.625 ;
        RECT 41.695 162.580 42.015 162.640 ;
        RECT 53.285 162.625 53.425 163.120 ;
        RECT 60.095 163.060 60.415 163.120 ;
        RECT 62.395 163.060 62.715 163.120 ;
        RECT 70.230 163.260 70.520 163.305 ;
        RECT 71.595 163.260 71.915 163.320 ;
        RECT 70.230 163.120 71.915 163.260 ;
        RECT 70.230 163.075 70.520 163.120 ;
        RECT 71.595 163.060 71.915 163.120 ;
        RECT 73.450 163.260 73.740 163.305 ;
        RECT 73.895 163.260 74.215 163.320 ;
        RECT 73.450 163.120 74.215 163.260 ;
        RECT 73.450 163.075 73.740 163.120 ;
        RECT 73.895 163.060 74.215 163.120 ;
        RECT 55.035 162.920 55.355 162.980 ;
        RECT 55.970 162.920 56.260 162.965 ;
        RECT 55.035 162.780 56.260 162.920 ;
        RECT 55.035 162.720 55.355 162.780 ;
        RECT 55.970 162.735 56.260 162.780 ;
        RECT 61.015 162.920 61.335 162.980 ;
        RECT 99.670 162.920 99.960 162.965 ;
        RECT 104.225 162.920 104.515 162.965 ;
        RECT 107.005 162.920 107.295 162.965 ;
        RECT 108.865 162.920 109.155 162.965 ;
        RECT 61.015 162.780 66.995 162.920 ;
        RECT 61.015 162.720 61.335 162.780 ;
        RECT 44.930 162.580 45.220 162.625 ;
        RECT 41.695 162.440 47.445 162.580 ;
        RECT 41.695 162.380 42.015 162.440 ;
        RECT 44.930 162.395 45.220 162.440 ;
        RECT 25.150 162.100 27.205 162.240 ;
        RECT 25.150 162.055 25.440 162.100 ;
        RECT 27.390 161.945 27.680 162.260 ;
        RECT 28.470 162.240 28.760 162.285 ;
        RECT 32.050 162.240 32.340 162.285 ;
        RECT 33.885 162.240 34.175 162.285 ;
        RECT 28.470 162.100 34.175 162.240 ;
        RECT 28.470 162.055 28.760 162.100 ;
        RECT 32.050 162.055 32.340 162.100 ;
        RECT 33.885 162.055 34.175 162.100 ;
        RECT 44.010 162.240 44.300 162.285 ;
        RECT 46.755 162.240 47.075 162.300 ;
        RECT 44.010 162.100 47.075 162.240 ;
        RECT 44.010 162.055 44.300 162.100 ;
        RECT 46.755 162.040 47.075 162.100 ;
        RECT 27.090 161.900 27.680 161.945 ;
        RECT 30.195 161.945 30.515 161.960 ;
        RECT 30.195 161.900 30.980 161.945 ;
        RECT 27.090 161.760 30.980 161.900 ;
        RECT 27.090 161.715 27.380 161.760 ;
        RECT 30.195 161.715 30.980 161.760 ;
        RECT 30.195 161.700 30.515 161.715 ;
        RECT 32.955 161.700 33.275 161.960 ;
        RECT 47.305 161.900 47.445 162.440 ;
        RECT 53.210 162.395 53.500 162.625 ;
        RECT 54.205 162.440 60.325 162.580 ;
        RECT 49.055 162.040 49.375 162.300 ;
        RECT 54.205 162.285 54.345 162.440 ;
        RECT 51.830 162.240 52.120 162.285 ;
        RECT 54.130 162.240 54.420 162.285 ;
        RECT 51.830 162.100 54.420 162.240 ;
        RECT 51.830 162.055 52.120 162.100 ;
        RECT 54.130 162.055 54.420 162.100 ;
        RECT 59.175 162.040 59.495 162.300 ;
        RECT 59.635 162.040 59.955 162.300 ;
        RECT 60.185 162.240 60.325 162.440 ;
        RECT 62.395 162.380 62.715 162.640 ;
        RECT 62.870 162.240 63.160 162.285 ;
        RECT 60.185 162.100 63.160 162.240 ;
        RECT 66.855 162.240 66.995 162.780 ;
        RECT 99.670 162.780 101.495 162.920 ;
        RECT 99.670 162.735 99.960 162.780 ;
        RECT 67.455 162.380 67.775 162.640 ;
        RECT 82.635 162.580 82.955 162.640 ;
        RECT 83.110 162.580 83.400 162.625 ;
        RECT 82.635 162.440 83.400 162.580 ;
        RECT 82.635 162.380 82.955 162.440 ;
        RECT 83.110 162.395 83.400 162.440 ;
        RECT 95.975 162.580 96.295 162.640 ;
        RECT 96.450 162.580 96.740 162.625 ;
        RECT 97.355 162.580 97.675 162.640 ;
        RECT 95.975 162.440 97.675 162.580 ;
        RECT 101.355 162.580 101.495 162.780 ;
        RECT 104.225 162.780 109.155 162.920 ;
        RECT 104.225 162.735 104.515 162.780 ;
        RECT 107.005 162.735 107.295 162.780 ;
        RECT 108.865 162.735 109.155 162.780 ;
        RECT 107.490 162.580 107.780 162.625 ;
        RECT 101.355 162.440 107.780 162.580 ;
        RECT 95.975 162.380 96.295 162.440 ;
        RECT 96.450 162.395 96.740 162.440 ;
        RECT 97.355 162.380 97.675 162.440 ;
        RECT 107.490 162.395 107.780 162.440 ;
        RECT 79.890 162.240 80.180 162.285 ;
        RECT 66.855 162.100 84.245 162.240 ;
        RECT 62.870 162.055 63.160 162.100 ;
        RECT 79.890 162.055 80.180 162.100 ;
        RECT 53.670 161.900 53.960 161.945 ;
        RECT 47.305 161.760 53.960 161.900 ;
        RECT 53.670 161.715 53.960 161.760 ;
        RECT 58.715 161.900 59.035 161.960 ;
        RECT 60.095 161.900 60.415 161.960 ;
        RECT 81.715 161.900 82.035 161.960 ;
        RECT 58.715 161.760 60.415 161.900 ;
        RECT 58.715 161.700 59.035 161.760 ;
        RECT 60.095 161.700 60.415 161.760 ;
        RECT 63.405 161.760 82.035 161.900 ;
        RECT 20.550 161.560 20.840 161.605 ;
        RECT 37.095 161.560 37.415 161.620 ;
        RECT 20.550 161.420 37.415 161.560 ;
        RECT 20.550 161.375 20.840 161.420 ;
        RECT 37.095 161.360 37.415 161.420 ;
        RECT 59.175 161.560 59.495 161.620 ;
        RECT 63.405 161.605 63.545 161.760 ;
        RECT 81.715 161.700 82.035 161.760 ;
        RECT 82.650 161.900 82.940 161.945 ;
        RECT 83.555 161.900 83.875 161.960 ;
        RECT 82.650 161.760 83.875 161.900 ;
        RECT 84.105 161.900 84.245 162.100 ;
        RECT 85.395 162.040 85.715 162.300 ;
        RECT 95.530 162.240 95.820 162.285 ;
        RECT 99.195 162.240 99.515 162.300 ;
        RECT 95.530 162.100 99.515 162.240 ;
        RECT 95.530 162.055 95.820 162.100 ;
        RECT 99.195 162.040 99.515 162.100 ;
        RECT 104.225 162.240 104.515 162.285 ;
        RECT 104.225 162.100 106.760 162.240 ;
        RECT 104.225 162.055 104.515 162.100 ;
        RECT 86.790 161.900 87.080 161.945 ;
        RECT 84.105 161.760 87.080 161.900 ;
        RECT 82.650 161.715 82.940 161.760 ;
        RECT 83.555 161.700 83.875 161.760 ;
        RECT 86.790 161.715 87.080 161.760 ;
        RECT 97.815 161.700 98.135 161.960 ;
        RECT 105.635 161.945 105.955 161.960 ;
        RECT 102.365 161.900 102.655 161.945 ;
        RECT 105.625 161.900 105.955 161.945 ;
        RECT 102.365 161.760 105.955 161.900 ;
        RECT 102.365 161.715 102.655 161.760 ;
        RECT 105.625 161.715 105.955 161.760 ;
        RECT 106.545 161.945 106.760 162.100 ;
        RECT 109.315 162.040 109.635 162.300 ;
        RECT 106.545 161.900 106.835 161.945 ;
        RECT 108.405 161.900 108.695 161.945 ;
        RECT 106.545 161.760 108.695 161.900 ;
        RECT 106.545 161.715 106.835 161.760 ;
        RECT 108.405 161.715 108.695 161.760 ;
        RECT 105.635 161.700 105.955 161.715 ;
        RECT 63.330 161.560 63.620 161.605 ;
        RECT 59.175 161.420 63.620 161.560 ;
        RECT 59.175 161.360 59.495 161.420 ;
        RECT 63.330 161.375 63.620 161.420 ;
        RECT 65.170 161.560 65.460 161.605 ;
        RECT 66.075 161.560 66.395 161.620 ;
        RECT 65.170 161.420 66.395 161.560 ;
        RECT 65.170 161.375 65.460 161.420 ;
        RECT 66.075 161.360 66.395 161.420 ;
        RECT 80.335 161.360 80.655 161.620 ;
        RECT 82.190 161.560 82.480 161.605 ;
        RECT 84.475 161.560 84.795 161.620 ;
        RECT 82.190 161.420 84.795 161.560 ;
        RECT 82.190 161.375 82.480 161.420 ;
        RECT 84.475 161.360 84.795 161.420 ;
        RECT 96.895 161.560 97.215 161.620 ;
        RECT 100.575 161.605 100.895 161.620 ;
        RECT 97.370 161.560 97.660 161.605 ;
        RECT 100.360 161.560 100.895 161.605 ;
        RECT 96.895 161.420 100.895 161.560 ;
        RECT 96.895 161.360 97.215 161.420 ;
        RECT 97.370 161.375 97.660 161.420 ;
        RECT 100.360 161.375 100.895 161.420 ;
        RECT 100.575 161.360 100.895 161.375 ;
        RECT 18.165 160.740 112.465 161.220 ;
        RECT 21.010 160.540 21.300 160.585 ;
        RECT 21.010 160.400 24.905 160.540 ;
        RECT 21.010 160.355 21.300 160.400 ;
        RECT 24.765 160.200 24.905 160.400 ;
        RECT 32.955 160.340 33.275 160.600 ;
        RECT 33.875 160.540 34.195 160.600 ;
        RECT 34.810 160.540 35.100 160.585 ;
        RECT 33.875 160.400 35.100 160.540 ;
        RECT 33.875 160.340 34.195 160.400 ;
        RECT 34.810 160.355 35.100 160.400 ;
        RECT 37.110 160.355 37.400 160.585 ;
        RECT 25.250 160.200 25.540 160.245 ;
        RECT 28.490 160.200 29.140 160.245 ;
        RECT 24.765 160.060 29.140 160.200 ;
        RECT 25.250 160.015 25.840 160.060 ;
        RECT 28.490 160.015 29.140 160.060 ;
        RECT 31.130 160.200 31.420 160.245 ;
        RECT 37.185 160.200 37.325 160.355 ;
        RECT 38.015 160.340 38.335 160.600 ;
        RECT 40.775 160.540 41.095 160.600 ;
        RECT 44.930 160.540 45.220 160.585 ;
        RECT 55.495 160.540 55.815 160.600 ;
        RECT 40.775 160.400 45.220 160.540 ;
        RECT 40.775 160.340 41.095 160.400 ;
        RECT 44.930 160.355 45.220 160.400 ;
        RECT 49.145 160.400 55.815 160.540 ;
        RECT 31.130 160.060 37.325 160.200 ;
        RECT 38.105 160.200 38.245 160.340 ;
        RECT 43.535 160.200 43.855 160.260 ;
        RECT 38.105 160.060 41.005 160.200 ;
        RECT 31.130 160.015 31.420 160.060 ;
        RECT 21.455 159.660 21.775 159.920 ;
        RECT 22.375 159.660 22.695 159.920 ;
        RECT 25.550 159.700 25.840 160.015 ;
        RECT 26.630 159.860 26.920 159.905 ;
        RECT 30.210 159.860 30.500 159.905 ;
        RECT 32.045 159.860 32.335 159.905 ;
        RECT 26.630 159.720 32.335 159.860 ;
        RECT 26.630 159.675 26.920 159.720 ;
        RECT 30.210 159.675 30.500 159.720 ;
        RECT 32.045 159.675 32.335 159.720 ;
        RECT 32.495 159.660 32.815 159.920 ;
        RECT 34.335 159.860 34.655 159.920 ;
        RECT 38.030 159.860 38.320 159.905 ;
        RECT 34.335 159.720 38.320 159.860 ;
        RECT 34.335 159.660 34.655 159.720 ;
        RECT 38.030 159.675 38.320 159.720 ;
        RECT 33.415 159.520 33.735 159.580 ;
        RECT 35.270 159.520 35.560 159.565 ;
        RECT 33.415 159.380 35.560 159.520 ;
        RECT 33.415 159.320 33.735 159.380 ;
        RECT 35.270 159.335 35.560 159.380 ;
        RECT 35.715 159.320 36.035 159.580 ;
        RECT 26.630 159.180 26.920 159.225 ;
        RECT 29.750 159.180 30.040 159.225 ;
        RECT 31.640 159.180 31.930 159.225 ;
        RECT 38.475 159.180 38.615 160.060 ;
        RECT 39.395 159.660 39.715 159.920 ;
        RECT 40.865 159.580 41.005 160.060 ;
        RECT 41.785 160.060 43.855 160.200 ;
        RECT 41.235 159.660 41.555 159.920 ;
        RECT 41.785 159.905 41.925 160.060 ;
        RECT 43.535 160.000 43.855 160.060 ;
        RECT 45.390 160.200 45.680 160.245 ;
        RECT 49.145 160.200 49.285 160.400 ;
        RECT 55.495 160.340 55.815 160.400 ;
        RECT 71.150 160.540 71.440 160.585 ;
        RECT 74.140 160.540 74.430 160.585 ;
        RECT 83.555 160.540 83.875 160.600 ;
        RECT 71.150 160.400 83.875 160.540 ;
        RECT 71.150 160.355 71.440 160.400 ;
        RECT 74.140 160.355 74.430 160.400 ;
        RECT 83.555 160.340 83.875 160.400 ;
        RECT 84.015 160.540 84.335 160.600 ;
        RECT 85.395 160.540 85.715 160.600 ;
        RECT 84.015 160.400 85.715 160.540 ;
        RECT 84.015 160.340 84.335 160.400 ;
        RECT 85.395 160.340 85.715 160.400 ;
        RECT 86.775 160.340 87.095 160.600 ;
        RECT 87.710 160.540 88.000 160.585 ;
        RECT 88.615 160.540 88.935 160.600 ;
        RECT 87.710 160.400 88.935 160.540 ;
        RECT 87.710 160.355 88.000 160.400 ;
        RECT 88.615 160.340 88.935 160.400 ;
        RECT 90.455 160.540 90.775 160.600 ;
        RECT 105.190 160.540 105.480 160.585 ;
        RECT 105.635 160.540 105.955 160.600 ;
        RECT 90.455 160.400 101.265 160.540 ;
        RECT 90.455 160.340 90.775 160.400 ;
        RECT 45.390 160.060 49.285 160.200 ;
        RECT 49.515 160.200 49.835 160.260 ;
        RECT 50.090 160.200 50.380 160.245 ;
        RECT 53.330 160.200 53.980 160.245 ;
        RECT 49.515 160.060 53.980 160.200 ;
        RECT 45.390 160.015 45.680 160.060 ;
        RECT 49.515 160.000 49.835 160.060 ;
        RECT 50.090 160.015 50.680 160.060 ;
        RECT 53.330 160.015 53.980 160.060 ;
        RECT 59.635 160.200 59.955 160.260 ;
        RECT 60.210 160.200 60.500 160.245 ;
        RECT 63.450 160.200 64.100 160.245 ;
        RECT 59.635 160.060 64.100 160.200 ;
        RECT 41.710 159.675 42.000 159.905 ;
        RECT 42.155 159.660 42.475 159.920 ;
        RECT 43.090 159.860 43.380 159.905 ;
        RECT 48.135 159.860 48.455 159.920 ;
        RECT 43.090 159.720 48.455 159.860 ;
        RECT 43.090 159.675 43.380 159.720 ;
        RECT 38.950 159.520 39.240 159.565 ;
        RECT 39.870 159.520 40.160 159.565 ;
        RECT 38.950 159.380 40.160 159.520 ;
        RECT 38.950 159.335 39.240 159.380 ;
        RECT 39.870 159.335 40.160 159.380 ;
        RECT 40.775 159.520 41.095 159.580 ;
        RECT 43.165 159.520 43.305 159.675 ;
        RECT 48.135 159.660 48.455 159.720 ;
        RECT 50.390 159.700 50.680 160.015 ;
        RECT 59.635 160.000 59.955 160.060 ;
        RECT 60.210 160.015 60.800 160.060 ;
        RECT 63.450 160.015 64.100 160.060 ;
        RECT 51.470 159.860 51.760 159.905 ;
        RECT 55.050 159.860 55.340 159.905 ;
        RECT 56.885 159.860 57.175 159.905 ;
        RECT 51.470 159.720 57.175 159.860 ;
        RECT 51.470 159.675 51.760 159.720 ;
        RECT 55.050 159.675 55.340 159.720 ;
        RECT 56.885 159.675 57.175 159.720 ;
        RECT 60.510 159.700 60.800 160.015 ;
        RECT 66.075 160.000 66.395 160.260 ;
        RECT 76.145 160.200 76.435 160.245 ;
        RECT 77.115 160.200 77.435 160.260 ;
        RECT 79.405 160.200 79.695 160.245 ;
        RECT 76.145 160.060 79.695 160.200 ;
        RECT 76.145 160.015 76.435 160.060 ;
        RECT 77.115 160.000 77.435 160.060 ;
        RECT 79.405 160.015 79.695 160.060 ;
        RECT 80.325 160.200 80.615 160.245 ;
        RECT 82.185 160.200 82.475 160.245 ;
        RECT 96.450 160.200 96.740 160.245 ;
        RECT 98.275 160.200 98.595 160.260 ;
        RECT 80.325 160.060 82.475 160.200 ;
        RECT 80.325 160.015 80.615 160.060 ;
        RECT 82.185 160.015 82.475 160.060 ;
        RECT 82.725 160.060 98.595 160.200 ;
        RECT 61.590 159.860 61.880 159.905 ;
        RECT 65.170 159.860 65.460 159.905 ;
        RECT 67.005 159.860 67.295 159.905 ;
        RECT 61.590 159.720 67.295 159.860 ;
        RECT 61.590 159.675 61.880 159.720 ;
        RECT 65.170 159.675 65.460 159.720 ;
        RECT 67.005 159.675 67.295 159.720 ;
        RECT 67.930 159.860 68.220 159.905 ;
        RECT 74.815 159.860 75.135 159.920 ;
        RECT 67.930 159.720 75.135 159.860 ;
        RECT 67.930 159.675 68.220 159.720 ;
        RECT 74.815 159.660 75.135 159.720 ;
        RECT 78.005 159.860 78.295 159.905 ;
        RECT 80.325 159.860 80.540 160.015 ;
        RECT 78.005 159.720 80.540 159.860 ;
        RECT 80.795 159.860 81.115 159.920 ;
        RECT 81.270 159.860 81.560 159.905 ;
        RECT 80.795 159.720 81.560 159.860 ;
        RECT 78.005 159.675 78.295 159.720 ;
        RECT 80.795 159.660 81.115 159.720 ;
        RECT 81.270 159.675 81.560 159.720 ;
        RECT 81.715 159.860 82.035 159.920 ;
        RECT 82.725 159.860 82.865 160.060 ;
        RECT 96.450 160.015 96.740 160.060 ;
        RECT 98.275 160.000 98.595 160.060 ;
        RECT 81.715 159.720 82.865 159.860 ;
        RECT 81.715 159.660 82.035 159.720 ;
        RECT 83.570 159.675 83.860 159.905 ;
        RECT 40.775 159.380 43.305 159.520 ;
        RECT 40.775 159.320 41.095 159.380 ;
        RECT 43.995 159.320 44.315 159.580 ;
        RECT 55.955 159.320 56.275 159.580 ;
        RECT 57.350 159.520 57.640 159.565 ;
        RECT 60.095 159.520 60.415 159.580 ;
        RECT 67.470 159.520 67.760 159.565 ;
        RECT 57.350 159.380 67.760 159.520 ;
        RECT 57.350 159.335 57.640 159.380 ;
        RECT 60.095 159.320 60.415 159.380 ;
        RECT 67.470 159.335 67.760 159.380 ;
        RECT 69.770 159.335 70.060 159.565 ;
        RECT 26.630 159.040 31.930 159.180 ;
        RECT 26.630 158.995 26.920 159.040 ;
        RECT 29.750 158.995 30.040 159.040 ;
        RECT 31.640 158.995 31.930 159.040 ;
        RECT 33.505 159.040 38.615 159.180 ;
        RECT 41.695 159.180 42.015 159.240 ;
        RECT 48.610 159.180 48.900 159.225 ;
        RECT 41.695 159.040 48.900 159.180 ;
        RECT 33.505 158.900 33.645 159.040 ;
        RECT 41.695 158.980 42.015 159.040 ;
        RECT 48.610 158.995 48.900 159.040 ;
        RECT 51.470 159.180 51.760 159.225 ;
        RECT 54.590 159.180 54.880 159.225 ;
        RECT 56.480 159.180 56.770 159.225 ;
        RECT 51.470 159.040 56.770 159.180 ;
        RECT 51.470 158.995 51.760 159.040 ;
        RECT 54.590 158.995 54.880 159.040 ;
        RECT 56.480 158.995 56.770 159.040 ;
        RECT 61.590 159.180 61.880 159.225 ;
        RECT 64.710 159.180 65.000 159.225 ;
        RECT 66.600 159.180 66.890 159.225 ;
        RECT 69.845 159.180 69.985 159.335 ;
        RECT 70.675 159.320 70.995 159.580 ;
        RECT 73.895 159.520 74.215 159.580 ;
        RECT 83.110 159.520 83.400 159.565 ;
        RECT 73.895 159.380 83.400 159.520 ;
        RECT 73.895 159.320 74.215 159.380 ;
        RECT 83.110 159.335 83.400 159.380 ;
        RECT 61.590 159.040 66.890 159.180 ;
        RECT 61.590 158.995 61.880 159.040 ;
        RECT 64.710 158.995 65.000 159.040 ;
        RECT 66.600 158.995 66.890 159.040 ;
        RECT 67.545 159.040 69.985 159.180 ;
        RECT 78.005 159.180 78.295 159.225 ;
        RECT 80.785 159.180 81.075 159.225 ;
        RECT 82.645 159.180 82.935 159.225 ;
        RECT 78.005 159.040 82.935 159.180 ;
        RECT 67.545 158.900 67.685 159.040 ;
        RECT 78.005 158.995 78.295 159.040 ;
        RECT 80.785 158.995 81.075 159.040 ;
        RECT 82.645 158.995 82.935 159.040 ;
        RECT 33.415 158.640 33.735 158.900 ;
        RECT 38.015 158.640 38.335 158.900 ;
        RECT 41.235 158.840 41.555 158.900 ;
        RECT 44.915 158.840 45.235 158.900 ;
        RECT 41.235 158.700 45.235 158.840 ;
        RECT 41.235 158.640 41.555 158.700 ;
        RECT 44.915 158.640 45.235 158.700 ;
        RECT 47.215 158.640 47.535 158.900 ;
        RECT 49.055 158.840 49.375 158.900 ;
        RECT 50.435 158.840 50.755 158.900 ;
        RECT 58.730 158.840 59.020 158.885 ;
        RECT 49.055 158.700 59.020 158.840 ;
        RECT 49.055 158.640 49.375 158.700 ;
        RECT 50.435 158.640 50.755 158.700 ;
        RECT 58.730 158.655 59.020 158.700 ;
        RECT 67.455 158.640 67.775 158.900 ;
        RECT 68.390 158.840 68.680 158.885 ;
        RECT 68.835 158.840 69.155 158.900 ;
        RECT 68.390 158.700 69.155 158.840 ;
        RECT 68.390 158.655 68.680 158.700 ;
        RECT 68.835 158.640 69.155 158.700 ;
        RECT 72.975 158.640 73.295 158.900 ;
        RECT 83.645 158.840 83.785 159.675 ;
        RECT 84.475 159.660 84.795 159.920 ;
        RECT 84.950 159.675 85.240 159.905 ;
        RECT 85.025 159.520 85.165 159.675 ;
        RECT 85.395 159.660 85.715 159.920 ;
        RECT 89.075 159.660 89.395 159.920 ;
        RECT 89.535 159.660 89.855 159.920 ;
        RECT 89.995 159.660 90.315 159.920 ;
        RECT 90.915 159.660 91.235 159.920 ;
        RECT 96.895 159.660 97.215 159.920 ;
        RECT 99.655 159.660 99.975 159.920 ;
        RECT 100.575 159.660 100.895 159.920 ;
        RECT 101.125 159.905 101.265 160.400 ;
        RECT 105.190 160.400 105.955 160.540 ;
        RECT 105.190 160.355 105.480 160.400 ;
        RECT 105.635 160.340 105.955 160.400 ;
        RECT 101.050 159.675 101.340 159.905 ;
        RECT 101.495 159.660 101.815 159.920 ;
        RECT 103.350 159.675 103.640 159.905 ;
        RECT 87.235 159.520 87.555 159.580 ;
        RECT 85.025 159.380 87.555 159.520 ;
        RECT 90.085 159.520 90.225 159.660 ;
        RECT 91.390 159.520 91.680 159.565 ;
        RECT 90.085 159.380 91.680 159.520 ;
        RECT 85.485 159.240 85.625 159.380 ;
        RECT 87.235 159.320 87.555 159.380 ;
        RECT 91.390 159.335 91.680 159.380 ;
        RECT 95.975 159.320 96.295 159.580 ;
        RECT 97.355 159.520 97.675 159.580 ;
        RECT 103.425 159.520 103.565 159.675 ;
        RECT 105.635 159.660 105.955 159.920 ;
        RECT 97.355 159.380 103.565 159.520 ;
        RECT 97.355 159.320 97.675 159.380 ;
        RECT 85.395 158.980 85.715 159.240 ;
        RECT 88.155 159.180 88.475 159.240 ;
        RECT 102.890 159.180 103.180 159.225 ;
        RECT 88.155 159.040 96.665 159.180 ;
        RECT 88.155 158.980 88.475 159.040 ;
        RECT 90.915 158.840 91.235 158.900 ;
        RECT 83.645 158.700 91.235 158.840 ;
        RECT 90.915 158.640 91.235 158.700 ;
        RECT 94.595 158.640 94.915 158.900 ;
        RECT 96.525 158.840 96.665 159.040 ;
        RECT 97.445 159.040 103.180 159.180 ;
        RECT 97.445 158.840 97.585 159.040 ;
        RECT 102.890 158.995 103.180 159.040 ;
        RECT 96.525 158.700 97.585 158.840 ;
        RECT 98.735 158.640 99.055 158.900 ;
        RECT 103.795 158.640 104.115 158.900 ;
        RECT 17.605 158.020 112.465 158.500 ;
        RECT 30.195 157.620 30.515 157.880 ;
        RECT 34.335 157.620 34.655 157.880 ;
        RECT 37.110 157.820 37.400 157.865 ;
        RECT 38.015 157.820 38.335 157.880 ;
        RECT 37.110 157.680 38.335 157.820 ;
        RECT 37.110 157.635 37.400 157.680 ;
        RECT 38.015 157.620 38.335 157.680 ;
        RECT 39.395 157.620 39.715 157.880 ;
        RECT 42.155 157.820 42.475 157.880 ;
        RECT 43.090 157.820 43.380 157.865 ;
        RECT 42.155 157.680 43.380 157.820 ;
        RECT 42.155 157.620 42.475 157.680 ;
        RECT 43.090 157.635 43.380 157.680 ;
        RECT 48.135 157.820 48.455 157.880 ;
        RECT 51.355 157.820 51.675 157.880 ;
        RECT 48.135 157.680 51.675 157.820 ;
        RECT 48.135 157.620 48.455 157.680 ;
        RECT 51.355 157.620 51.675 157.680 ;
        RECT 58.715 157.820 59.035 157.880 ;
        RECT 60.555 157.820 60.875 157.880 ;
        RECT 58.715 157.680 60.875 157.820 ;
        RECT 58.715 157.620 59.035 157.680 ;
        RECT 60.555 157.620 60.875 157.680 ;
        RECT 62.945 157.680 76.885 157.820 ;
        RECT 31.575 157.480 31.895 157.540 ;
        RECT 35.730 157.480 36.020 157.525 ;
        RECT 42.615 157.480 42.935 157.540 ;
        RECT 31.575 157.340 36.020 157.480 ;
        RECT 31.575 157.280 31.895 157.340 ;
        RECT 35.730 157.295 36.020 157.340 ;
        RECT 39.025 157.340 42.935 157.480 ;
        RECT 31.665 157.140 31.805 157.280 ;
        RECT 36.175 157.140 36.495 157.200 ;
        RECT 39.025 157.185 39.165 157.340 ;
        RECT 42.615 157.280 42.935 157.340 ;
        RECT 45.950 157.480 46.240 157.525 ;
        RECT 49.070 157.480 49.360 157.525 ;
        RECT 50.960 157.480 51.250 157.525 ;
        RECT 60.095 157.480 60.415 157.540 ;
        RECT 45.950 157.340 51.250 157.480 ;
        RECT 45.950 157.295 46.240 157.340 ;
        RECT 49.070 157.295 49.360 157.340 ;
        RECT 50.960 157.295 51.250 157.340 ;
        RECT 51.905 157.340 60.415 157.480 ;
        RECT 30.745 157.000 31.805 157.140 ;
        RECT 32.585 157.000 36.495 157.140 ;
        RECT 22.390 156.800 22.680 156.845 ;
        RECT 24.675 156.800 24.995 156.860 ;
        RECT 22.390 156.660 24.995 156.800 ;
        RECT 22.390 156.615 22.680 156.660 ;
        RECT 24.675 156.600 24.995 156.660 ;
        RECT 30.195 156.800 30.515 156.860 ;
        RECT 30.745 156.845 30.885 157.000 ;
        RECT 30.670 156.800 30.960 156.845 ;
        RECT 30.195 156.660 30.960 156.800 ;
        RECT 30.195 156.600 30.515 156.660 ;
        RECT 30.670 156.615 30.960 156.660 ;
        RECT 31.130 156.615 31.420 156.845 ;
        RECT 31.205 156.460 31.345 156.615 ;
        RECT 32.035 156.600 32.355 156.860 ;
        RECT 32.585 156.845 32.725 157.000 ;
        RECT 36.175 156.940 36.495 157.000 ;
        RECT 38.950 156.955 39.240 157.185 ;
        RECT 46.755 157.140 47.075 157.200 ;
        RECT 40.865 157.000 47.075 157.140 ;
        RECT 32.510 156.615 32.800 156.845 ;
        RECT 32.970 156.800 33.260 156.845 ;
        RECT 34.795 156.800 35.115 156.860 ;
        RECT 32.970 156.660 35.115 156.800 ;
        RECT 32.970 156.615 33.260 156.660 ;
        RECT 34.795 156.600 35.115 156.660 ;
        RECT 36.650 156.615 36.940 156.845 ;
        RECT 38.030 156.615 38.320 156.845 ;
        RECT 38.475 156.800 38.795 156.860 ;
        RECT 40.865 156.845 41.005 157.000 ;
        RECT 46.755 156.940 47.075 157.000 ;
        RECT 47.215 157.140 47.535 157.200 ;
        RECT 51.905 157.185 52.045 157.340 ;
        RECT 60.095 157.280 60.415 157.340 ;
        RECT 50.450 157.140 50.740 157.185 ;
        RECT 47.215 157.000 50.740 157.140 ;
        RECT 47.215 156.940 47.535 157.000 ;
        RECT 50.450 156.955 50.740 157.000 ;
        RECT 51.830 156.955 52.120 157.185 ;
        RECT 40.790 156.800 41.080 156.845 ;
        RECT 38.475 156.660 41.080 156.800 ;
        RECT 33.415 156.460 33.735 156.520 ;
        RECT 31.205 156.320 33.735 156.460 ;
        RECT 33.415 156.260 33.735 156.320 ;
        RECT 23.310 156.120 23.600 156.165 ;
        RECT 25.135 156.120 25.455 156.180 ;
        RECT 23.310 155.980 25.455 156.120 ;
        RECT 36.725 156.120 36.865 156.615 ;
        RECT 38.105 156.460 38.245 156.615 ;
        RECT 38.475 156.600 38.795 156.660 ;
        RECT 40.790 156.615 41.080 156.660 ;
        RECT 41.250 156.615 41.540 156.845 ;
        RECT 38.935 156.460 39.255 156.520 ;
        RECT 38.105 156.320 39.255 156.460 ;
        RECT 38.935 156.260 39.255 156.320 ;
        RECT 39.855 156.460 40.175 156.520 ;
        RECT 41.325 156.460 41.465 156.615 ;
        RECT 41.695 156.600 42.015 156.860 ;
        RECT 42.155 156.800 42.475 156.860 ;
        RECT 42.630 156.800 42.920 156.845 ;
        RECT 42.155 156.660 42.920 156.800 ;
        RECT 42.155 156.600 42.475 156.660 ;
        RECT 42.630 156.615 42.920 156.660 ;
        RECT 43.995 156.460 44.315 156.520 ;
        RECT 44.870 156.505 45.160 156.820 ;
        RECT 45.950 156.800 46.240 156.845 ;
        RECT 49.530 156.800 49.820 156.845 ;
        RECT 51.365 156.800 51.655 156.845 ;
        RECT 45.950 156.660 51.655 156.800 ;
        RECT 45.950 156.615 46.240 156.660 ;
        RECT 49.530 156.615 49.820 156.660 ;
        RECT 51.365 156.615 51.655 156.660 ;
        RECT 52.275 156.600 52.595 156.860 ;
        RECT 55.495 156.800 55.815 156.860 ;
        RECT 57.795 156.800 58.115 156.860 ;
        RECT 55.495 156.660 58.115 156.800 ;
        RECT 55.495 156.600 55.815 156.660 ;
        RECT 57.795 156.600 58.115 156.660 ;
        RECT 58.255 156.600 58.575 156.860 ;
        RECT 58.730 156.615 59.020 156.845 ;
        RECT 39.855 156.320 44.315 156.460 ;
        RECT 39.855 156.260 40.175 156.320 ;
        RECT 43.995 156.260 44.315 156.320 ;
        RECT 44.570 156.460 45.160 156.505 ;
        RECT 45.375 156.460 45.695 156.520 ;
        RECT 47.810 156.460 48.460 156.505 ;
        RECT 44.570 156.320 48.460 156.460 ;
        RECT 44.570 156.275 44.860 156.320 ;
        RECT 45.375 156.260 45.695 156.320 ;
        RECT 47.810 156.275 48.460 156.320 ;
        RECT 56.415 156.460 56.735 156.520 ;
        RECT 58.805 156.460 58.945 156.615 ;
        RECT 59.175 156.600 59.495 156.860 ;
        RECT 60.110 156.800 60.400 156.845 ;
        RECT 60.555 156.800 60.875 156.860 ;
        RECT 62.945 156.845 63.085 157.680 ;
        RECT 70.645 157.480 70.935 157.525 ;
        RECT 73.425 157.480 73.715 157.525 ;
        RECT 75.285 157.480 75.575 157.525 ;
        RECT 70.645 157.340 75.575 157.480 ;
        RECT 76.745 157.480 76.885 157.680 ;
        RECT 77.115 157.620 77.435 157.880 ;
        RECT 82.175 157.820 82.495 157.880 ;
        RECT 89.075 157.820 89.395 157.880 ;
        RECT 77.665 157.680 89.395 157.820 ;
        RECT 77.665 157.480 77.805 157.680 ;
        RECT 82.175 157.620 82.495 157.680 ;
        RECT 89.075 157.620 89.395 157.680 ;
        RECT 98.275 157.865 98.595 157.880 ;
        RECT 98.275 157.635 98.810 157.865 ;
        RECT 98.275 157.620 98.595 157.635 ;
        RECT 76.745 157.340 77.805 157.480 ;
        RECT 81.255 157.480 81.575 157.540 ;
        RECT 97.355 157.480 97.675 157.540 ;
        RECT 81.255 157.340 97.675 157.480 ;
        RECT 70.645 157.295 70.935 157.340 ;
        RECT 73.425 157.295 73.715 157.340 ;
        RECT 75.285 157.295 75.575 157.340 ;
        RECT 81.255 157.280 81.575 157.340 ;
        RECT 97.355 157.280 97.675 157.340 ;
        RECT 102.385 157.480 102.675 157.525 ;
        RECT 105.165 157.480 105.455 157.525 ;
        RECT 107.025 157.480 107.315 157.525 ;
        RECT 102.385 157.340 107.315 157.480 ;
        RECT 102.385 157.295 102.675 157.340 ;
        RECT 105.165 157.295 105.455 157.340 ;
        RECT 107.025 157.295 107.315 157.340 ;
        RECT 72.515 157.140 72.835 157.200 ;
        RECT 63.405 157.000 72.835 157.140 ;
        RECT 63.405 156.860 63.545 157.000 ;
        RECT 72.515 156.940 72.835 157.000 ;
        RECT 72.975 157.140 73.295 157.200 ;
        RECT 73.910 157.140 74.200 157.185 ;
        RECT 72.975 157.000 74.200 157.140 ;
        RECT 72.975 156.940 73.295 157.000 ;
        RECT 73.910 156.955 74.200 157.000 ;
        RECT 74.355 157.140 74.675 157.200 ;
        RECT 75.750 157.140 76.040 157.185 ;
        RECT 74.355 157.000 76.040 157.140 ;
        RECT 74.355 156.940 74.675 157.000 ;
        RECT 75.750 156.955 76.040 157.000 ;
        RECT 60.110 156.660 60.875 156.800 ;
        RECT 60.110 156.615 60.400 156.660 ;
        RECT 60.555 156.600 60.875 156.660 ;
        RECT 62.870 156.615 63.160 156.845 ;
        RECT 63.315 156.600 63.635 156.860 ;
        RECT 63.790 156.615 64.080 156.845 ;
        RECT 64.710 156.800 65.000 156.845 ;
        RECT 65.615 156.800 65.935 156.860 ;
        RECT 64.710 156.660 65.935 156.800 ;
        RECT 64.710 156.615 65.000 156.660 ;
        RECT 56.415 156.320 58.945 156.460 ;
        RECT 59.635 156.460 59.955 156.520 ;
        RECT 63.865 156.460 64.005 156.615 ;
        RECT 65.615 156.600 65.935 156.660 ;
        RECT 70.645 156.800 70.935 156.845 ;
        RECT 75.275 156.800 75.595 156.860 ;
        RECT 81.345 156.845 81.485 157.280 ;
        RECT 81.730 157.140 82.020 157.185 ;
        RECT 83.095 157.140 83.415 157.200 ;
        RECT 85.395 157.140 85.715 157.200 ;
        RECT 81.730 157.000 83.415 157.140 ;
        RECT 81.730 156.955 82.020 157.000 ;
        RECT 83.095 156.940 83.415 157.000 ;
        RECT 84.105 157.000 85.715 157.140 ;
        RECT 76.670 156.800 76.960 156.845 ;
        RECT 70.645 156.660 73.180 156.800 ;
        RECT 70.645 156.615 70.935 156.660 ;
        RECT 65.155 156.460 65.475 156.520 ;
        RECT 68.835 156.505 69.155 156.520 ;
        RECT 72.965 156.505 73.180 156.660 ;
        RECT 75.275 156.660 76.960 156.800 ;
        RECT 75.275 156.600 75.595 156.660 ;
        RECT 76.670 156.615 76.960 156.660 ;
        RECT 81.270 156.615 81.560 156.845 ;
        RECT 82.650 156.615 82.940 156.845 ;
        RECT 59.635 156.320 62.625 156.460 ;
        RECT 63.865 156.320 65.475 156.460 ;
        RECT 56.415 156.260 56.735 156.320 ;
        RECT 59.635 156.260 59.955 156.320 ;
        RECT 48.595 156.120 48.915 156.180 ;
        RECT 52.735 156.120 53.055 156.180 ;
        RECT 36.725 155.980 53.055 156.120 ;
        RECT 23.310 155.935 23.600 155.980 ;
        RECT 25.135 155.920 25.455 155.980 ;
        RECT 48.595 155.920 48.915 155.980 ;
        RECT 52.735 155.920 53.055 155.980 ;
        RECT 55.495 156.120 55.815 156.180 ;
        RECT 56.890 156.120 57.180 156.165 ;
        RECT 55.495 155.980 57.180 156.120 ;
        RECT 55.495 155.920 55.815 155.980 ;
        RECT 56.890 155.935 57.180 155.980 ;
        RECT 61.475 155.920 61.795 156.180 ;
        RECT 62.485 156.120 62.625 156.320 ;
        RECT 65.155 156.260 65.475 156.320 ;
        RECT 68.785 156.460 69.155 156.505 ;
        RECT 72.045 156.460 72.335 156.505 ;
        RECT 68.785 156.320 72.335 156.460 ;
        RECT 68.785 156.275 69.155 156.320 ;
        RECT 72.045 156.275 72.335 156.320 ;
        RECT 72.965 156.460 73.255 156.505 ;
        RECT 74.825 156.460 75.115 156.505 ;
        RECT 72.965 156.320 75.115 156.460 ;
        RECT 72.965 156.275 73.255 156.320 ;
        RECT 74.825 156.275 75.115 156.320 ;
        RECT 75.735 156.460 76.055 156.520 ;
        RECT 82.725 156.460 82.865 156.615 ;
        RECT 83.555 156.600 83.875 156.860 ;
        RECT 84.105 156.845 84.245 157.000 ;
        RECT 85.395 156.940 85.715 157.000 ;
        RECT 85.945 157.000 92.525 157.140 ;
        RECT 84.030 156.615 84.320 156.845 ;
        RECT 84.475 156.600 84.795 156.860 ;
        RECT 85.945 156.800 86.085 157.000 ;
        RECT 85.025 156.660 86.085 156.800 ;
        RECT 85.025 156.460 85.165 156.660 ;
        RECT 87.235 156.600 87.555 156.860 ;
        RECT 87.695 156.600 88.015 156.860 ;
        RECT 89.075 156.800 89.395 156.860 ;
        RECT 90.470 156.800 90.760 156.845 ;
        RECT 89.075 156.660 90.760 156.800 ;
        RECT 89.075 156.600 89.395 156.660 ;
        RECT 90.470 156.615 90.760 156.660 ;
        RECT 90.930 156.615 91.220 156.845 ;
        RECT 89.535 156.460 89.855 156.520 ;
        RECT 91.005 156.460 91.145 156.615 ;
        RECT 91.375 156.600 91.695 156.860 ;
        RECT 92.385 156.845 92.525 157.000 ;
        RECT 93.675 156.940 93.995 157.200 ;
        RECT 98.735 157.140 99.055 157.200 ;
        RECT 105.650 157.140 105.940 157.185 ;
        RECT 94.225 157.000 95.285 157.140 ;
        RECT 92.310 156.800 92.600 156.845 ;
        RECT 94.225 156.800 94.365 157.000 ;
        RECT 92.310 156.660 94.365 156.800 ;
        RECT 92.310 156.615 92.600 156.660 ;
        RECT 94.595 156.600 94.915 156.860 ;
        RECT 95.145 156.800 95.285 157.000 ;
        RECT 98.735 157.000 105.940 157.140 ;
        RECT 98.735 156.940 99.055 157.000 ;
        RECT 105.650 156.955 105.940 157.000 ;
        RECT 99.655 156.800 99.975 156.860 ;
        RECT 95.145 156.660 99.975 156.800 ;
        RECT 99.655 156.600 99.975 156.660 ;
        RECT 102.385 156.800 102.675 156.845 ;
        RECT 107.490 156.800 107.780 156.845 ;
        RECT 109.315 156.800 109.635 156.860 ;
        RECT 102.385 156.660 104.920 156.800 ;
        RECT 102.385 156.615 102.675 156.660 ;
        RECT 75.735 156.320 85.165 156.460 ;
        RECT 85.485 156.320 91.145 156.460 ;
        RECT 91.465 156.460 91.605 156.600 ;
        RECT 103.795 156.505 104.115 156.520 ;
        RECT 94.150 156.460 94.440 156.505 ;
        RECT 91.465 156.320 94.440 156.460 ;
        RECT 68.835 156.260 69.155 156.275 ;
        RECT 75.735 156.260 76.055 156.320 ;
        RECT 66.780 156.120 67.070 156.165 ;
        RECT 70.675 156.120 70.995 156.180 ;
        RECT 62.485 155.980 70.995 156.120 ;
        RECT 66.780 155.935 67.070 155.980 ;
        RECT 70.675 155.920 70.995 155.980 ;
        RECT 72.515 156.120 72.835 156.180 ;
        RECT 79.415 156.120 79.735 156.180 ;
        RECT 85.485 156.120 85.625 156.320 ;
        RECT 89.535 156.260 89.855 156.320 ;
        RECT 94.150 156.275 94.440 156.320 ;
        RECT 100.525 156.460 100.815 156.505 ;
        RECT 103.785 156.460 104.115 156.505 ;
        RECT 100.525 156.320 104.115 156.460 ;
        RECT 100.525 156.275 100.815 156.320 ;
        RECT 103.785 156.275 104.115 156.320 ;
        RECT 104.705 156.505 104.920 156.660 ;
        RECT 107.105 156.660 109.635 156.800 ;
        RECT 104.705 156.460 104.995 156.505 ;
        RECT 106.565 156.460 106.855 156.505 ;
        RECT 104.705 156.320 106.855 156.460 ;
        RECT 104.705 156.275 104.995 156.320 ;
        RECT 106.565 156.275 106.855 156.320 ;
        RECT 103.795 156.260 104.115 156.275 ;
        RECT 72.515 155.980 85.625 156.120 ;
        RECT 85.870 156.120 86.160 156.165 ;
        RECT 86.775 156.120 87.095 156.180 ;
        RECT 85.870 155.980 87.095 156.120 ;
        RECT 72.515 155.920 72.835 155.980 ;
        RECT 79.415 155.920 79.735 155.980 ;
        RECT 85.870 155.935 86.160 155.980 ;
        RECT 86.775 155.920 87.095 155.980 ;
        RECT 88.615 155.920 88.935 156.180 ;
        RECT 89.075 155.920 89.395 156.180 ;
        RECT 96.450 156.120 96.740 156.165 ;
        RECT 96.895 156.120 97.215 156.180 ;
        RECT 96.450 155.980 97.215 156.120 ;
        RECT 96.450 155.935 96.740 155.980 ;
        RECT 96.895 155.920 97.215 155.980 ;
        RECT 99.195 156.120 99.515 156.180 ;
        RECT 107.105 156.120 107.245 156.660 ;
        RECT 107.490 156.615 107.780 156.660 ;
        RECT 109.315 156.600 109.635 156.660 ;
        RECT 99.195 155.980 107.245 156.120 ;
        RECT 99.195 155.920 99.515 155.980 ;
        RECT 18.165 155.300 112.465 155.780 ;
        RECT 21.455 155.100 21.775 155.160 ;
        RECT 38.475 155.100 38.795 155.160 ;
        RECT 38.950 155.100 39.240 155.145 ;
        RECT 21.455 154.960 29.505 155.100 ;
        RECT 21.455 154.900 21.775 154.960 ;
        RECT 21.545 154.465 21.685 154.900 ;
        RECT 22.375 154.560 22.695 154.820 ;
        RECT 25.250 154.760 25.540 154.805 ;
        RECT 28.490 154.760 29.140 154.805 ;
        RECT 25.250 154.620 29.140 154.760 ;
        RECT 29.365 154.760 29.505 154.960 ;
        RECT 38.475 154.960 39.240 155.100 ;
        RECT 38.475 154.900 38.795 154.960 ;
        RECT 38.950 154.915 39.240 154.960 ;
        RECT 42.615 155.100 42.935 155.160 ;
        RECT 44.470 155.100 44.760 155.145 ;
        RECT 42.615 154.960 44.760 155.100 ;
        RECT 42.615 154.900 42.935 154.960 ;
        RECT 44.470 154.915 44.760 154.960 ;
        RECT 44.915 155.100 45.235 155.160 ;
        RECT 44.915 154.960 50.205 155.100 ;
        RECT 44.915 154.900 45.235 154.960 ;
        RECT 42.170 154.760 42.460 154.805 ;
        RECT 48.150 154.760 48.440 154.805 ;
        RECT 29.365 154.620 34.105 154.760 ;
        RECT 25.250 154.575 25.840 154.620 ;
        RECT 28.490 154.575 29.140 154.620 ;
        RECT 21.470 154.235 21.760 154.465 ;
        RECT 25.550 154.260 25.840 154.575 ;
        RECT 26.630 154.420 26.920 154.465 ;
        RECT 30.210 154.420 30.500 154.465 ;
        RECT 32.045 154.420 32.335 154.465 ;
        RECT 26.630 154.280 32.335 154.420 ;
        RECT 21.010 154.080 21.300 154.125 ;
        RECT 25.685 154.080 25.825 154.260 ;
        RECT 26.630 154.235 26.920 154.280 ;
        RECT 30.210 154.235 30.500 154.280 ;
        RECT 32.045 154.235 32.335 154.280 ;
        RECT 32.495 154.220 32.815 154.480 ;
        RECT 33.965 154.465 34.105 154.620 ;
        RECT 42.170 154.620 48.440 154.760 ;
        RECT 42.170 154.575 42.460 154.620 ;
        RECT 48.150 154.575 48.440 154.620 ;
        RECT 50.065 154.480 50.205 154.960 ;
        RECT 55.955 154.900 56.275 155.160 ;
        RECT 85.395 155.100 85.715 155.160 ;
        RECT 59.725 154.960 85.715 155.100 ;
        RECT 59.725 154.760 59.865 154.960 ;
        RECT 85.395 154.900 85.715 154.960 ;
        RECT 59.265 154.620 59.865 154.760 ;
        RECT 62.510 154.760 62.800 154.805 ;
        RECT 64.695 154.760 65.015 154.820 ;
        RECT 65.750 154.760 66.400 154.805 ;
        RECT 62.510 154.620 66.400 154.760 ;
        RECT 33.890 154.235 34.180 154.465 ;
        RECT 35.270 154.420 35.560 154.465 ;
        RECT 36.635 154.420 36.955 154.480 ;
        RECT 35.270 154.280 36.955 154.420 ;
        RECT 35.270 154.235 35.560 154.280 ;
        RECT 36.635 154.220 36.955 154.280 ;
        RECT 38.015 154.220 38.335 154.480 ;
        RECT 38.935 154.420 39.255 154.480 ;
        RECT 40.790 154.420 41.080 154.465 ;
        RECT 38.935 154.280 41.080 154.420 ;
        RECT 38.935 154.220 39.255 154.280 ;
        RECT 40.790 154.235 41.080 154.280 ;
        RECT 44.010 154.420 44.300 154.465 ;
        RECT 44.455 154.420 44.775 154.480 ;
        RECT 44.010 154.280 44.775 154.420 ;
        RECT 44.010 154.235 44.300 154.280 ;
        RECT 44.455 154.220 44.775 154.280 ;
        RECT 46.755 154.420 47.075 154.480 ;
        RECT 49.515 154.420 49.835 154.480 ;
        RECT 46.755 154.280 49.835 154.420 ;
        RECT 46.755 154.220 47.075 154.280 ;
        RECT 49.515 154.220 49.835 154.280 ;
        RECT 49.975 154.220 50.295 154.480 ;
        RECT 50.435 154.220 50.755 154.480 ;
        RECT 51.355 154.220 51.675 154.480 ;
        RECT 53.210 154.420 53.500 154.465 ;
        RECT 55.035 154.420 55.355 154.480 ;
        RECT 53.210 154.280 55.355 154.420 ;
        RECT 53.210 154.235 53.500 154.280 ;
        RECT 55.035 154.220 55.355 154.280 ;
        RECT 58.715 154.220 59.035 154.480 ;
        RECT 59.265 154.465 59.405 154.620 ;
        RECT 62.510 154.575 63.100 154.620 ;
        RECT 59.190 154.235 59.480 154.465 ;
        RECT 59.635 154.220 59.955 154.480 ;
        RECT 60.555 154.420 60.875 154.480 ;
        RECT 60.555 154.280 62.625 154.420 ;
        RECT 60.555 154.220 60.875 154.280 ;
        RECT 21.010 153.940 25.825 154.080 ;
        RECT 31.130 154.080 31.420 154.125 ;
        RECT 41.235 154.080 41.555 154.140 ;
        RECT 31.130 153.940 41.555 154.080 ;
        RECT 21.010 153.895 21.300 153.940 ;
        RECT 31.130 153.895 31.420 153.940 ;
        RECT 41.235 153.880 41.555 153.940 ;
        RECT 41.710 153.895 42.000 154.125 ;
        RECT 43.075 154.080 43.395 154.140 ;
        RECT 43.550 154.080 43.840 154.125 ;
        RECT 44.915 154.080 45.235 154.140 ;
        RECT 43.075 153.940 45.235 154.080 ;
        RECT 26.630 153.740 26.920 153.785 ;
        RECT 29.750 153.740 30.040 153.785 ;
        RECT 31.640 153.740 31.930 153.785 ;
        RECT 40.775 153.740 41.095 153.800 ;
        RECT 26.630 153.600 31.930 153.740 ;
        RECT 26.630 153.555 26.920 153.600 ;
        RECT 29.750 153.555 30.040 153.600 ;
        RECT 31.640 153.555 31.930 153.600 ;
        RECT 33.965 153.600 41.095 153.740 ;
        RECT 41.785 153.740 41.925 153.895 ;
        RECT 43.075 153.880 43.395 153.940 ;
        RECT 43.550 153.895 43.840 153.940 ;
        RECT 44.915 153.880 45.235 153.940 ;
        RECT 46.295 154.080 46.615 154.140 ;
        RECT 52.275 154.080 52.595 154.140 ;
        RECT 61.030 154.080 61.320 154.125 ;
        RECT 46.295 153.940 61.320 154.080 ;
        RECT 62.485 154.080 62.625 154.280 ;
        RECT 62.810 154.260 63.100 154.575 ;
        RECT 64.695 154.560 65.015 154.620 ;
        RECT 65.750 154.575 66.400 154.620 ;
        RECT 77.065 154.760 77.355 154.805 ;
        RECT 79.415 154.760 79.735 154.820 ;
        RECT 80.325 154.760 80.615 154.805 ;
        RECT 77.065 154.620 80.615 154.760 ;
        RECT 77.065 154.575 77.355 154.620 ;
        RECT 79.415 154.560 79.735 154.620 ;
        RECT 80.325 154.575 80.615 154.620 ;
        RECT 81.245 154.760 81.535 154.805 ;
        RECT 83.105 154.760 83.395 154.805 ;
        RECT 81.245 154.620 83.395 154.760 ;
        RECT 81.245 154.575 81.535 154.620 ;
        RECT 83.105 154.575 83.395 154.620 ;
        RECT 84.935 154.760 85.255 154.820 ;
        RECT 95.055 154.805 95.375 154.820 ;
        RECT 86.790 154.760 87.080 154.805 ;
        RECT 84.935 154.620 87.080 154.760 ;
        RECT 63.890 154.420 64.180 154.465 ;
        RECT 67.470 154.420 67.760 154.465 ;
        RECT 69.305 154.420 69.595 154.465 ;
        RECT 63.890 154.280 69.595 154.420 ;
        RECT 63.890 154.235 64.180 154.280 ;
        RECT 67.470 154.235 67.760 154.280 ;
        RECT 69.305 154.235 69.595 154.280 ;
        RECT 69.770 154.420 70.060 154.465 ;
        RECT 73.895 154.420 74.215 154.480 ;
        RECT 69.770 154.280 74.215 154.420 ;
        RECT 69.770 154.235 70.060 154.280 ;
        RECT 73.895 154.220 74.215 154.280 ;
        RECT 78.925 154.420 79.215 154.465 ;
        RECT 81.245 154.420 81.460 154.575 ;
        RECT 84.935 154.560 85.255 154.620 ;
        RECT 86.790 154.575 87.080 154.620 ;
        RECT 91.785 154.760 92.075 154.805 ;
        RECT 95.045 154.760 95.375 154.805 ;
        RECT 91.785 154.620 95.375 154.760 ;
        RECT 91.785 154.575 92.075 154.620 ;
        RECT 95.045 154.575 95.375 154.620 ;
        RECT 95.055 154.560 95.375 154.575 ;
        RECT 95.965 154.760 96.255 154.805 ;
        RECT 97.825 154.760 98.115 154.805 ;
        RECT 95.965 154.620 98.115 154.760 ;
        RECT 95.965 154.575 96.255 154.620 ;
        RECT 97.825 154.575 98.115 154.620 ;
        RECT 104.250 154.760 104.900 154.805 ;
        RECT 107.015 154.760 107.335 154.820 ;
        RECT 107.850 154.760 108.140 154.805 ;
        RECT 104.250 154.620 108.140 154.760 ;
        RECT 104.250 154.575 104.900 154.620 ;
        RECT 78.925 154.280 81.460 154.420 ;
        RECT 78.925 154.235 79.215 154.280 ;
        RECT 82.175 154.220 82.495 154.480 ;
        RECT 87.235 154.220 87.555 154.480 ;
        RECT 93.645 154.420 93.935 154.465 ;
        RECT 95.965 154.420 96.180 154.575 ;
        RECT 107.015 154.560 107.335 154.620 ;
        RECT 107.550 154.575 108.140 154.620 ;
        RECT 93.645 154.280 96.180 154.420 ;
        RECT 93.645 154.235 93.935 154.280 ;
        RECT 96.895 154.220 97.215 154.480 ;
        RECT 101.055 154.420 101.345 154.465 ;
        RECT 102.890 154.420 103.180 154.465 ;
        RECT 106.470 154.420 106.760 154.465 ;
        RECT 101.055 154.280 106.760 154.420 ;
        RECT 101.055 154.235 101.345 154.280 ;
        RECT 102.890 154.235 103.180 154.280 ;
        RECT 106.470 154.235 106.760 154.280 ;
        RECT 107.550 154.260 107.840 154.575 ;
        RECT 110.695 154.560 111.015 154.820 ;
        RECT 65.615 154.080 65.935 154.140 ;
        RECT 62.485 153.940 65.935 154.080 ;
        RECT 46.295 153.880 46.615 153.940 ;
        RECT 52.275 153.880 52.595 153.940 ;
        RECT 61.030 153.895 61.320 153.940 ;
        RECT 65.615 153.880 65.935 153.940 ;
        RECT 68.375 153.880 68.695 154.140 ;
        RECT 73.985 154.080 74.125 154.220 ;
        RECT 84.030 154.080 84.320 154.125 ;
        RECT 73.985 153.940 84.320 154.080 ;
        RECT 84.030 153.895 84.320 153.940 ;
        RECT 84.935 154.080 85.255 154.140 ;
        RECT 85.870 154.080 86.160 154.125 ;
        RECT 84.935 153.940 86.160 154.080 ;
        RECT 84.935 153.880 85.255 153.940 ;
        RECT 85.870 153.895 86.160 153.940 ;
        RECT 87.695 154.080 88.015 154.140 ;
        RECT 89.780 154.080 90.070 154.125 ;
        RECT 91.375 154.080 91.695 154.140 ;
        RECT 87.695 153.940 91.695 154.080 ;
        RECT 87.695 153.880 88.015 153.940 ;
        RECT 89.780 153.895 90.070 153.940 ;
        RECT 91.375 153.880 91.695 153.940 ;
        RECT 98.735 154.080 99.055 154.140 ;
        RECT 100.590 154.080 100.880 154.125 ;
        RECT 98.735 153.940 100.880 154.080 ;
        RECT 98.735 153.880 99.055 153.940 ;
        RECT 100.590 153.895 100.880 153.940 ;
        RECT 101.955 153.880 102.275 154.140 ;
        RECT 43.995 153.740 44.315 153.800 ;
        RECT 41.785 153.600 44.315 153.740 ;
        RECT 30.195 153.400 30.515 153.460 ;
        RECT 33.965 153.400 34.105 153.600 ;
        RECT 40.775 153.540 41.095 153.600 ;
        RECT 43.995 153.540 44.315 153.600 ;
        RECT 49.975 153.740 50.295 153.800 ;
        RECT 52.735 153.740 53.055 153.800 ;
        RECT 56.415 153.740 56.735 153.800 ;
        RECT 49.975 153.600 56.735 153.740 ;
        RECT 49.975 153.540 50.295 153.600 ;
        RECT 52.735 153.540 53.055 153.600 ;
        RECT 56.415 153.540 56.735 153.600 ;
        RECT 63.890 153.740 64.180 153.785 ;
        RECT 67.010 153.740 67.300 153.785 ;
        RECT 68.900 153.740 69.190 153.785 ;
        RECT 63.890 153.600 69.190 153.740 ;
        RECT 63.890 153.555 64.180 153.600 ;
        RECT 67.010 153.555 67.300 153.600 ;
        RECT 68.900 153.555 69.190 153.600 ;
        RECT 78.925 153.740 79.215 153.785 ;
        RECT 81.705 153.740 81.995 153.785 ;
        RECT 83.565 153.740 83.855 153.785 ;
        RECT 78.925 153.600 83.855 153.740 ;
        RECT 78.925 153.555 79.215 153.600 ;
        RECT 81.705 153.555 81.995 153.600 ;
        RECT 83.565 153.555 83.855 153.600 ;
        RECT 93.645 153.740 93.935 153.785 ;
        RECT 96.425 153.740 96.715 153.785 ;
        RECT 98.285 153.740 98.575 153.785 ;
        RECT 93.645 153.600 98.575 153.740 ;
        RECT 93.645 153.555 93.935 153.600 ;
        RECT 96.425 153.555 96.715 153.600 ;
        RECT 98.285 153.555 98.575 153.600 ;
        RECT 101.460 153.740 101.750 153.785 ;
        RECT 103.350 153.740 103.640 153.785 ;
        RECT 106.470 153.740 106.760 153.785 ;
        RECT 101.460 153.600 106.760 153.740 ;
        RECT 101.460 153.555 101.750 153.600 ;
        RECT 103.350 153.555 103.640 153.600 ;
        RECT 106.470 153.555 106.760 153.600 ;
        RECT 30.195 153.260 34.105 153.400 ;
        RECT 34.350 153.400 34.640 153.445 ;
        RECT 34.795 153.400 35.115 153.460 ;
        RECT 34.350 153.260 35.115 153.400 ;
        RECT 30.195 153.200 30.515 153.260 ;
        RECT 34.350 153.215 34.640 153.260 ;
        RECT 34.795 153.200 35.115 153.260 ;
        RECT 36.175 153.200 36.495 153.460 ;
        RECT 39.855 153.200 40.175 153.460 ;
        RECT 42.155 153.200 42.475 153.460 ;
        RECT 46.310 153.400 46.600 153.445 ;
        RECT 46.755 153.400 47.075 153.460 ;
        RECT 46.310 153.260 47.075 153.400 ;
        RECT 46.310 153.215 46.600 153.260 ;
        RECT 46.755 153.200 47.075 153.260 ;
        RECT 54.115 153.400 54.435 153.460 ;
        RECT 57.350 153.400 57.640 153.445 ;
        RECT 54.115 153.260 57.640 153.400 ;
        RECT 54.115 153.200 54.435 153.260 ;
        RECT 57.350 153.215 57.640 153.260 ;
        RECT 57.795 153.400 58.115 153.460 ;
        RECT 62.395 153.400 62.715 153.460 ;
        RECT 57.795 153.260 62.715 153.400 ;
        RECT 57.795 153.200 58.115 153.260 ;
        RECT 62.395 153.200 62.715 153.260 ;
        RECT 65.155 153.400 65.475 153.460 ;
        RECT 75.060 153.400 75.350 153.445 ;
        RECT 80.335 153.400 80.655 153.460 ;
        RECT 65.155 153.260 80.655 153.400 ;
        RECT 65.155 153.200 65.475 153.260 ;
        RECT 75.060 153.215 75.350 153.260 ;
        RECT 80.335 153.200 80.655 153.260 ;
        RECT 89.090 153.400 89.380 153.445 ;
        RECT 89.535 153.400 89.855 153.460 ;
        RECT 89.090 153.260 89.855 153.400 ;
        RECT 89.090 153.215 89.380 153.260 ;
        RECT 89.535 153.200 89.855 153.260 ;
        RECT 17.605 152.580 112.465 153.060 ;
        RECT 25.610 152.380 25.900 152.425 ;
        RECT 26.055 152.380 26.375 152.440 ;
        RECT 32.035 152.380 32.355 152.440 ;
        RECT 25.610 152.240 32.355 152.380 ;
        RECT 25.610 152.195 25.900 152.240 ;
        RECT 26.055 152.180 26.375 152.240 ;
        RECT 32.035 152.180 32.355 152.240 ;
        RECT 36.635 152.380 36.955 152.440 ;
        RECT 36.635 152.240 38.245 152.380 ;
        RECT 36.635 152.180 36.955 152.240 ;
        RECT 28.470 152.040 28.760 152.085 ;
        RECT 31.590 152.040 31.880 152.085 ;
        RECT 33.480 152.040 33.770 152.085 ;
        RECT 28.470 151.900 33.770 152.040 ;
        RECT 38.105 152.040 38.245 152.240 ;
        RECT 38.935 152.180 39.255 152.440 ;
        RECT 41.235 152.380 41.555 152.440 ;
        RECT 53.210 152.380 53.500 152.425 ;
        RECT 41.235 152.240 53.500 152.380 ;
        RECT 41.235 152.180 41.555 152.240 ;
        RECT 53.210 152.195 53.500 152.240 ;
        RECT 55.510 152.380 55.800 152.425 ;
        RECT 61.030 152.380 61.320 152.425 ;
        RECT 55.510 152.240 61.320 152.380 ;
        RECT 55.510 152.195 55.800 152.240 ;
        RECT 61.030 152.195 61.320 152.240 ;
        RECT 67.010 152.380 67.300 152.425 ;
        RECT 68.375 152.380 68.695 152.440 ;
        RECT 82.175 152.380 82.495 152.440 ;
        RECT 82.650 152.380 82.940 152.425 ;
        RECT 67.010 152.240 68.695 152.380 ;
        RECT 67.010 152.195 67.300 152.240 ;
        RECT 68.375 152.180 68.695 152.240 ;
        RECT 73.065 152.240 80.105 152.380 ;
        RECT 39.640 152.040 39.930 152.085 ;
        RECT 42.615 152.040 42.935 152.100 ;
        RECT 38.105 151.900 39.165 152.040 ;
        RECT 28.470 151.855 28.760 151.900 ;
        RECT 31.590 151.855 31.880 151.900 ;
        RECT 33.480 151.855 33.770 151.900 ;
        RECT 32.495 151.700 32.815 151.760 ;
        RECT 34.350 151.700 34.640 151.745 ;
        RECT 32.495 151.560 34.640 151.700 ;
        RECT 32.495 151.500 32.815 151.560 ;
        RECT 34.350 151.515 34.640 151.560 ;
        RECT 35.255 151.700 35.575 151.760 ;
        RECT 35.255 151.560 37.785 151.700 ;
        RECT 35.255 151.500 35.575 151.560 ;
        RECT 27.390 151.065 27.680 151.380 ;
        RECT 28.470 151.360 28.760 151.405 ;
        RECT 32.050 151.360 32.340 151.405 ;
        RECT 33.885 151.360 34.175 151.405 ;
        RECT 28.470 151.220 34.175 151.360 ;
        RECT 28.470 151.175 28.760 151.220 ;
        RECT 32.050 151.175 32.340 151.220 ;
        RECT 33.885 151.175 34.175 151.220 ;
        RECT 35.730 151.360 36.020 151.405 ;
        RECT 36.175 151.360 36.495 151.420 ;
        RECT 35.730 151.220 36.495 151.360 ;
        RECT 35.730 151.175 36.020 151.220 ;
        RECT 27.090 151.020 27.680 151.065 ;
        RECT 29.735 151.020 30.055 151.080 ;
        RECT 30.330 151.020 30.980 151.065 ;
        RECT 27.090 150.880 30.980 151.020 ;
        RECT 27.090 150.835 27.380 150.880 ;
        RECT 29.735 150.820 30.055 150.880 ;
        RECT 30.330 150.835 30.980 150.880 ;
        RECT 32.970 151.020 33.260 151.065 ;
        RECT 34.335 151.020 34.655 151.080 ;
        RECT 32.970 150.880 34.655 151.020 ;
        RECT 32.970 150.835 33.260 150.880 ;
        RECT 34.335 150.820 34.655 150.880 ;
        RECT 35.805 150.680 35.945 151.175 ;
        RECT 36.175 151.160 36.495 151.220 ;
        RECT 36.635 151.160 36.955 151.420 ;
        RECT 37.095 151.160 37.415 151.420 ;
        RECT 37.645 151.405 37.785 151.560 ;
        RECT 39.025 151.420 39.165 151.900 ;
        RECT 39.640 151.900 42.935 152.040 ;
        RECT 39.640 151.855 39.930 151.900 ;
        RECT 42.615 151.840 42.935 151.900 ;
        RECT 43.505 152.040 43.795 152.085 ;
        RECT 46.285 152.040 46.575 152.085 ;
        RECT 48.145 152.040 48.435 152.085 ;
        RECT 61.475 152.040 61.795 152.100 ;
        RECT 69.540 152.040 69.830 152.085 ;
        RECT 71.135 152.040 71.455 152.100 ;
        RECT 43.505 151.900 48.435 152.040 ;
        RECT 43.505 151.855 43.795 151.900 ;
        RECT 46.285 151.855 46.575 151.900 ;
        RECT 48.145 151.855 48.435 151.900 ;
        RECT 55.125 151.900 61.795 152.040 ;
        RECT 46.755 151.500 47.075 151.760 ;
        RECT 55.125 151.745 55.265 151.900 ;
        RECT 61.475 151.840 61.795 151.900 ;
        RECT 62.945 151.900 71.455 152.040 ;
        RECT 55.050 151.515 55.340 151.745 ;
        RECT 56.875 151.500 57.195 151.760 ;
        RECT 62.945 151.745 63.085 151.900 ;
        RECT 69.540 151.855 69.830 151.900 ;
        RECT 71.135 151.840 71.455 151.900 ;
        RECT 57.350 151.700 57.640 151.745 ;
        RECT 62.870 151.700 63.160 151.745 ;
        RECT 57.350 151.560 63.160 151.700 ;
        RECT 57.350 151.515 57.640 151.560 ;
        RECT 62.870 151.515 63.160 151.560 ;
        RECT 64.250 151.700 64.540 151.745 ;
        RECT 73.065 151.700 73.205 152.240 ;
        RECT 73.405 152.040 73.695 152.085 ;
        RECT 76.185 152.040 76.475 152.085 ;
        RECT 78.045 152.040 78.335 152.085 ;
        RECT 73.405 151.900 78.335 152.040 ;
        RECT 73.405 151.855 73.695 151.900 ;
        RECT 76.185 151.855 76.475 151.900 ;
        RECT 78.045 151.855 78.335 151.900 ;
        RECT 79.965 152.040 80.105 152.240 ;
        RECT 82.175 152.240 82.940 152.380 ;
        RECT 82.175 152.180 82.495 152.240 ;
        RECT 82.650 152.195 82.940 152.240 ;
        RECT 88.615 152.180 88.935 152.440 ;
        RECT 93.675 152.380 93.995 152.440 ;
        RECT 89.165 152.240 93.995 152.380 ;
        RECT 89.165 152.040 89.305 152.240 ;
        RECT 93.675 152.180 93.995 152.240 ;
        RECT 94.595 152.380 94.915 152.440 ;
        RECT 95.530 152.380 95.820 152.425 ;
        RECT 94.595 152.240 95.820 152.380 ;
        RECT 94.595 152.180 94.915 152.240 ;
        RECT 95.530 152.195 95.820 152.240 ;
        RECT 106.570 152.380 106.860 152.425 ;
        RECT 107.015 152.380 107.335 152.440 ;
        RECT 106.570 152.240 107.335 152.380 ;
        RECT 106.570 152.195 106.860 152.240 ;
        RECT 107.015 152.180 107.335 152.240 ;
        RECT 79.965 151.900 89.305 152.040 ;
        RECT 90.470 152.040 90.760 152.085 ;
        RECT 101.955 152.040 102.275 152.100 ;
        RECT 90.470 151.900 102.275 152.040 ;
        RECT 64.250 151.560 73.205 151.700 ;
        RECT 73.895 151.700 74.215 151.760 ;
        RECT 73.895 151.560 76.425 151.700 ;
        RECT 64.250 151.515 64.540 151.560 ;
        RECT 73.895 151.500 74.215 151.560 ;
        RECT 37.570 151.175 37.860 151.405 ;
        RECT 38.935 151.160 39.255 151.420 ;
        RECT 43.505 151.360 43.795 151.405 ;
        RECT 43.505 151.220 46.040 151.360 ;
        RECT 43.505 151.175 43.795 151.220 ;
        RECT 41.645 151.020 41.935 151.065 ;
        RECT 43.075 151.020 43.395 151.080 ;
        RECT 45.825 151.065 46.040 151.220 ;
        RECT 48.595 151.160 48.915 151.420 ;
        RECT 54.115 151.160 54.435 151.420 ;
        RECT 55.495 151.160 55.815 151.420 ;
        RECT 61.475 151.360 61.795 151.420 ;
        RECT 61.950 151.360 62.240 151.405 ;
        RECT 61.475 151.220 62.240 151.360 ;
        RECT 61.475 151.160 61.795 151.220 ;
        RECT 61.950 151.175 62.240 151.220 ;
        RECT 62.395 151.360 62.715 151.420 ;
        RECT 64.710 151.360 65.000 151.405 ;
        RECT 62.395 151.220 65.000 151.360 ;
        RECT 44.905 151.020 45.195 151.065 ;
        RECT 41.645 150.880 45.195 151.020 ;
        RECT 41.645 150.835 41.935 150.880 ;
        RECT 43.075 150.820 43.395 150.880 ;
        RECT 44.905 150.835 45.195 150.880 ;
        RECT 45.825 151.020 46.115 151.065 ;
        RECT 47.685 151.020 47.975 151.065 ;
        RECT 60.555 151.020 60.875 151.080 ;
        RECT 45.825 150.880 47.975 151.020 ;
        RECT 45.825 150.835 46.115 150.880 ;
        RECT 47.685 150.835 47.975 150.880 ;
        RECT 53.055 150.880 60.875 151.020 ;
        RECT 62.025 151.020 62.165 151.175 ;
        RECT 62.395 151.160 62.715 151.220 ;
        RECT 64.710 151.175 65.000 151.220 ;
        RECT 65.155 151.160 65.475 151.420 ;
        RECT 73.405 151.360 73.695 151.405 ;
        RECT 76.285 151.360 76.425 151.560 ;
        RECT 76.655 151.500 76.975 151.760 ;
        RECT 79.965 151.745 80.105 151.900 ;
        RECT 90.470 151.855 90.760 151.900 ;
        RECT 101.955 151.840 102.275 151.900 ;
        RECT 79.890 151.515 80.180 151.745 ;
        RECT 80.335 151.500 80.655 151.760 ;
        RECT 86.775 151.700 87.095 151.760 ;
        RECT 86.775 151.560 88.845 151.700 ;
        RECT 86.775 151.500 87.095 151.560 ;
        RECT 78.510 151.360 78.800 151.405 ;
        RECT 73.405 151.220 75.940 151.360 ;
        RECT 76.285 151.220 78.800 151.360 ;
        RECT 73.405 151.175 73.695 151.220 ;
        RECT 63.315 151.020 63.635 151.080 ;
        RECT 74.815 151.065 75.135 151.080 ;
        RECT 62.025 150.880 63.635 151.020 ;
        RECT 47.215 150.680 47.535 150.740 ;
        RECT 53.055 150.680 53.195 150.880 ;
        RECT 60.555 150.820 60.875 150.880 ;
        RECT 63.315 150.820 63.635 150.880 ;
        RECT 71.545 151.020 71.835 151.065 ;
        RECT 74.805 151.020 75.135 151.065 ;
        RECT 71.545 150.880 75.135 151.020 ;
        RECT 71.545 150.835 71.835 150.880 ;
        RECT 74.805 150.835 75.135 150.880 ;
        RECT 75.725 151.065 75.940 151.220 ;
        RECT 78.510 151.175 78.800 151.220 ;
        RECT 80.810 151.360 81.100 151.405 ;
        RECT 87.695 151.360 88.015 151.420 ;
        RECT 80.810 151.220 88.015 151.360 ;
        RECT 80.810 151.175 81.100 151.220 ;
        RECT 87.695 151.160 88.015 151.220 ;
        RECT 88.155 151.160 88.475 151.420 ;
        RECT 88.705 151.360 88.845 151.560 ;
        RECT 89.075 151.500 89.395 151.760 ;
        RECT 89.550 151.360 89.840 151.405 ;
        RECT 88.705 151.220 89.840 151.360 ;
        RECT 89.550 151.175 89.840 151.220 ;
        RECT 95.990 151.360 96.280 151.405 ;
        RECT 105.635 151.360 105.955 151.420 ;
        RECT 106.110 151.360 106.400 151.405 ;
        RECT 95.990 151.220 106.400 151.360 ;
        RECT 95.990 151.175 96.280 151.220 ;
        RECT 105.635 151.160 105.955 151.220 ;
        RECT 106.110 151.175 106.400 151.220 ;
        RECT 75.725 151.020 76.015 151.065 ;
        RECT 77.585 151.020 77.875 151.065 ;
        RECT 75.725 150.880 77.875 151.020 ;
        RECT 75.725 150.835 76.015 150.880 ;
        RECT 77.585 150.835 77.875 150.880 ;
        RECT 74.815 150.820 75.135 150.835 ;
        RECT 85.395 150.820 85.715 151.080 ;
        RECT 92.310 151.020 92.600 151.065 ;
        RECT 93.675 151.020 93.995 151.080 ;
        RECT 92.310 150.880 93.995 151.020 ;
        RECT 92.310 150.835 92.600 150.880 ;
        RECT 93.675 150.820 93.995 150.880 ;
        RECT 35.805 150.540 53.195 150.680 ;
        RECT 57.335 150.680 57.655 150.740 ;
        RECT 57.810 150.680 58.100 150.725 ;
        RECT 57.335 150.540 58.100 150.680 ;
        RECT 47.215 150.480 47.535 150.540 ;
        RECT 57.335 150.480 57.655 150.540 ;
        RECT 57.810 150.495 58.100 150.540 ;
        RECT 59.635 150.480 59.955 150.740 ;
        RECT 73.435 150.680 73.755 150.740 ;
        RECT 84.030 150.680 84.320 150.725 ;
        RECT 84.935 150.680 85.255 150.740 ;
        RECT 73.435 150.540 85.255 150.680 ;
        RECT 73.435 150.480 73.755 150.540 ;
        RECT 84.030 150.495 84.320 150.540 ;
        RECT 84.935 150.480 85.255 150.540 ;
        RECT 18.165 149.860 112.465 150.340 ;
        RECT 21.010 149.660 21.300 149.705 ;
        RECT 39.855 149.660 40.175 149.720 ;
        RECT 21.010 149.520 24.905 149.660 ;
        RECT 21.010 149.475 21.300 149.520 ;
        RECT 24.765 149.320 24.905 149.520 ;
        RECT 31.205 149.520 40.175 149.660 ;
        RECT 31.205 149.365 31.345 149.520 ;
        RECT 39.855 149.460 40.175 149.520 ;
        RECT 43.075 149.460 43.395 149.720 ;
        RECT 43.995 149.460 44.315 149.720 ;
        RECT 44.455 149.660 44.775 149.720 ;
        RECT 52.520 149.660 52.810 149.705 ;
        RECT 57.335 149.660 57.655 149.720 ;
        RECT 44.455 149.520 57.655 149.660 ;
        RECT 44.455 149.460 44.775 149.520 ;
        RECT 52.520 149.475 52.810 149.520 ;
        RECT 57.335 149.460 57.655 149.520 ;
        RECT 64.250 149.660 64.540 149.705 ;
        RECT 64.695 149.660 65.015 149.720 ;
        RECT 64.250 149.520 65.015 149.660 ;
        RECT 64.250 149.475 64.540 149.520 ;
        RECT 64.695 149.460 65.015 149.520 ;
        RECT 71.135 149.460 71.455 149.720 ;
        RECT 72.990 149.475 73.280 149.705 ;
        RECT 74.370 149.660 74.660 149.705 ;
        RECT 74.815 149.660 75.135 149.720 ;
        RECT 74.370 149.520 75.135 149.660 ;
        RECT 74.370 149.475 74.660 149.520 ;
        RECT 25.250 149.320 25.540 149.365 ;
        RECT 28.490 149.320 29.140 149.365 ;
        RECT 24.765 149.180 29.140 149.320 ;
        RECT 25.250 149.135 25.840 149.180 ;
        RECT 28.490 149.135 29.140 149.180 ;
        RECT 31.130 149.135 31.420 149.365 ;
        RECT 34.450 149.320 34.740 149.365 ;
        RECT 37.690 149.320 38.340 149.365 ;
        RECT 34.450 149.180 38.340 149.320 ;
        RECT 34.450 149.135 35.040 149.180 ;
        RECT 37.690 149.135 38.340 149.180 ;
        RECT 21.455 148.780 21.775 149.040 ;
        RECT 25.550 148.820 25.840 149.135 ;
        RECT 34.750 149.040 35.040 149.135 ;
        RECT 40.315 149.120 40.635 149.380 ;
        RECT 40.775 149.320 41.095 149.380 ;
        RECT 43.535 149.320 43.855 149.380 ;
        RECT 54.525 149.320 54.815 149.365 ;
        RECT 55.955 149.320 56.275 149.380 ;
        RECT 57.785 149.320 58.075 149.365 ;
        RECT 40.775 149.180 42.845 149.320 ;
        RECT 40.775 149.120 41.095 149.180 ;
        RECT 26.630 148.980 26.920 149.025 ;
        RECT 30.210 148.980 30.500 149.025 ;
        RECT 32.045 148.980 32.335 149.025 ;
        RECT 26.630 148.840 32.335 148.980 ;
        RECT 26.630 148.795 26.920 148.840 ;
        RECT 30.210 148.795 30.500 148.840 ;
        RECT 32.045 148.795 32.335 148.840 ;
        RECT 32.495 148.780 32.815 149.040 ;
        RECT 34.750 148.820 35.115 149.040 ;
        RECT 42.705 149.025 42.845 149.180 ;
        RECT 43.535 149.180 46.065 149.320 ;
        RECT 43.535 149.120 43.855 149.180 ;
        RECT 34.795 148.780 35.115 148.820 ;
        RECT 35.830 148.980 36.120 149.025 ;
        RECT 39.410 148.980 39.700 149.025 ;
        RECT 41.245 148.980 41.535 149.025 ;
        RECT 35.830 148.840 41.535 148.980 ;
        RECT 35.830 148.795 36.120 148.840 ;
        RECT 39.410 148.795 39.700 148.840 ;
        RECT 41.245 148.795 41.535 148.840 ;
        RECT 42.630 148.795 42.920 149.025 ;
        RECT 45.375 148.780 45.695 149.040 ;
        RECT 45.925 149.025 46.065 149.180 ;
        RECT 54.525 149.180 58.075 149.320 ;
        RECT 54.525 149.135 54.815 149.180 ;
        RECT 55.955 149.120 56.275 149.180 ;
        RECT 57.785 149.135 58.075 149.180 ;
        RECT 58.705 149.320 58.995 149.365 ;
        RECT 60.565 149.320 60.855 149.365 ;
        RECT 58.705 149.180 60.855 149.320 ;
        RECT 73.065 149.320 73.205 149.475 ;
        RECT 74.815 149.460 75.135 149.520 ;
        RECT 78.970 149.660 79.260 149.705 ;
        RECT 79.415 149.660 79.735 149.720 ;
        RECT 78.970 149.520 79.735 149.660 ;
        RECT 78.970 149.475 79.260 149.520 ;
        RECT 79.415 149.460 79.735 149.520 ;
        RECT 76.655 149.320 76.975 149.380 ;
        RECT 73.065 149.180 76.975 149.320 ;
        RECT 58.705 149.135 58.995 149.180 ;
        RECT 60.565 149.135 60.855 149.180 ;
        RECT 45.850 148.795 46.140 149.025 ;
        RECT 46.295 148.780 46.615 149.040 ;
        RECT 47.215 148.780 47.535 149.040 ;
        RECT 56.385 148.980 56.675 149.025 ;
        RECT 58.705 148.980 58.920 149.135 ;
        RECT 76.655 149.120 76.975 149.180 ;
        RECT 83.095 149.320 83.415 149.380 ;
        RECT 84.425 149.320 84.715 149.365 ;
        RECT 87.685 149.320 87.975 149.365 ;
        RECT 83.095 149.180 87.975 149.320 ;
        RECT 83.095 149.120 83.415 149.180 ;
        RECT 84.425 149.135 84.715 149.180 ;
        RECT 87.685 149.135 87.975 149.180 ;
        RECT 88.605 149.320 88.895 149.365 ;
        RECT 90.465 149.320 90.755 149.365 ;
        RECT 88.605 149.180 90.755 149.320 ;
        RECT 88.605 149.135 88.895 149.180 ;
        RECT 90.465 149.135 90.755 149.180 ;
        RECT 56.385 148.840 58.920 148.980 ;
        RECT 56.385 148.795 56.675 148.840 ;
        RECT 59.635 148.780 59.955 149.040 ;
        RECT 60.095 148.980 60.415 149.040 ;
        RECT 61.490 148.980 61.780 149.025 ;
        RECT 60.095 148.840 61.780 148.980 ;
        RECT 60.095 148.780 60.415 148.840 ;
        RECT 61.490 148.795 61.780 148.840 ;
        RECT 61.935 148.980 62.255 149.040 ;
        RECT 63.790 148.980 64.080 149.025 ;
        RECT 61.935 148.840 64.080 148.980 ;
        RECT 61.935 148.780 62.255 148.840 ;
        RECT 63.790 148.795 64.080 148.840 ;
        RECT 74.830 148.980 75.120 149.025 ;
        RECT 75.275 148.980 75.595 149.040 ;
        RECT 74.830 148.840 75.595 148.980 ;
        RECT 74.830 148.795 75.120 148.840 ;
        RECT 75.275 148.780 75.595 148.840 ;
        RECT 79.430 148.980 79.720 149.025 ;
        RECT 79.875 148.980 80.195 149.040 ;
        RECT 79.430 148.840 80.195 148.980 ;
        RECT 79.430 148.795 79.720 148.840 ;
        RECT 79.875 148.780 80.195 148.840 ;
        RECT 86.285 148.980 86.575 149.025 ;
        RECT 88.605 148.980 88.820 149.135 ;
        RECT 86.285 148.840 88.820 148.980 ;
        RECT 86.285 148.795 86.575 148.840 ;
        RECT 89.535 148.780 89.855 149.040 ;
        RECT 91.390 148.980 91.680 149.025 ;
        RECT 98.735 148.980 99.055 149.040 ;
        RECT 91.390 148.840 99.055 148.980 ;
        RECT 91.390 148.795 91.680 148.840 ;
        RECT 98.735 148.780 99.055 148.840 ;
        RECT 101.050 148.795 101.340 149.025 ;
        RECT 22.375 148.440 22.695 148.700 ;
        RECT 32.585 148.640 32.725 148.780 ;
        RECT 41.710 148.640 42.000 148.685 ;
        RECT 32.585 148.500 42.000 148.640 ;
        RECT 41.710 148.455 42.000 148.500 ;
        RECT 44.915 148.640 45.235 148.700 ;
        RECT 56.875 148.640 57.195 148.700 ;
        RECT 69.770 148.640 70.060 148.685 ;
        RECT 44.915 148.500 70.060 148.640 ;
        RECT 26.630 148.300 26.920 148.345 ;
        RECT 29.750 148.300 30.040 148.345 ;
        RECT 31.640 148.300 31.930 148.345 ;
        RECT 26.630 148.160 31.930 148.300 ;
        RECT 26.630 148.115 26.920 148.160 ;
        RECT 29.750 148.115 30.040 148.160 ;
        RECT 31.640 148.115 31.930 148.160 ;
        RECT 35.830 148.300 36.120 148.345 ;
        RECT 38.950 148.300 39.240 148.345 ;
        RECT 40.840 148.300 41.130 148.345 ;
        RECT 35.830 148.160 41.130 148.300 ;
        RECT 41.785 148.300 41.925 148.455 ;
        RECT 44.915 148.440 45.235 148.500 ;
        RECT 56.875 148.440 57.195 148.500 ;
        RECT 69.770 148.455 70.060 148.500 ;
        RECT 70.690 148.640 70.980 148.685 ;
        RECT 82.420 148.640 82.710 148.685 ;
        RECT 87.235 148.640 87.555 148.700 ;
        RECT 70.690 148.500 87.555 148.640 ;
        RECT 101.125 148.640 101.265 148.795 ;
        RECT 101.495 148.780 101.815 149.040 ;
        RECT 102.890 148.640 103.180 148.685 ;
        RECT 107.475 148.640 107.795 148.700 ;
        RECT 101.125 148.500 107.795 148.640 ;
        RECT 70.690 148.455 70.980 148.500 ;
        RECT 82.420 148.455 82.710 148.500 ;
        RECT 87.235 148.440 87.555 148.500 ;
        RECT 102.890 148.455 103.180 148.500 ;
        RECT 107.475 148.440 107.795 148.500 ;
        RECT 48.595 148.300 48.915 148.360 ;
        RECT 41.785 148.160 48.915 148.300 ;
        RECT 35.830 148.115 36.120 148.160 ;
        RECT 38.950 148.115 39.240 148.160 ;
        RECT 40.840 148.115 41.130 148.160 ;
        RECT 48.595 148.100 48.915 148.160 ;
        RECT 56.385 148.300 56.675 148.345 ;
        RECT 59.165 148.300 59.455 148.345 ;
        RECT 61.025 148.300 61.315 148.345 ;
        RECT 56.385 148.160 61.315 148.300 ;
        RECT 56.385 148.115 56.675 148.160 ;
        RECT 59.165 148.115 59.455 148.160 ;
        RECT 61.025 148.115 61.315 148.160 ;
        RECT 86.285 148.300 86.575 148.345 ;
        RECT 89.065 148.300 89.355 148.345 ;
        RECT 90.925 148.300 91.215 148.345 ;
        RECT 86.285 148.160 91.215 148.300 ;
        RECT 86.285 148.115 86.575 148.160 ;
        RECT 89.065 148.115 89.355 148.160 ;
        RECT 90.925 148.115 91.215 148.160 ;
        RECT 100.115 148.300 100.435 148.360 ;
        RECT 100.590 148.300 100.880 148.345 ;
        RECT 100.115 148.160 100.880 148.300 ;
        RECT 100.115 148.100 100.435 148.160 ;
        RECT 100.590 148.115 100.880 148.160 ;
        RECT 32.955 147.960 33.275 148.020 ;
        RECT 36.635 147.960 36.955 148.020 ;
        RECT 32.955 147.820 36.955 147.960 ;
        RECT 32.955 147.760 33.275 147.820 ;
        RECT 36.635 147.760 36.955 147.820 ;
        RECT 17.605 147.140 112.465 147.620 ;
        RECT 29.735 146.740 30.055 147.000 ;
        RECT 34.335 146.740 34.655 147.000 ;
        RECT 39.410 146.940 39.700 146.985 ;
        RECT 40.315 146.940 40.635 147.000 ;
        RECT 39.410 146.800 40.635 146.940 ;
        RECT 39.410 146.755 39.700 146.800 ;
        RECT 40.315 146.740 40.635 146.800 ;
        RECT 42.155 146.940 42.475 147.000 ;
        RECT 43.090 146.940 43.380 146.985 ;
        RECT 42.155 146.800 43.380 146.940 ;
        RECT 42.155 146.740 42.475 146.800 ;
        RECT 43.090 146.755 43.380 146.800 ;
        RECT 55.955 146.740 56.275 147.000 ;
        RECT 28.830 146.600 29.120 146.645 ;
        RECT 60.095 146.600 60.415 146.660 ;
        RECT 62.855 146.600 63.175 146.660 ;
        RECT 28.830 146.460 32.265 146.600 ;
        RECT 28.830 146.415 29.120 146.460 ;
        RECT 26.055 146.060 26.375 146.320 ;
        RECT 32.125 146.305 32.265 146.460 ;
        RECT 50.985 146.460 63.175 146.600 ;
        RECT 31.590 146.075 31.880 146.305 ;
        RECT 32.050 146.260 32.340 146.305 ;
        RECT 33.875 146.260 34.195 146.320 ;
        RECT 32.050 146.120 34.195 146.260 ;
        RECT 32.050 146.075 32.340 146.120 ;
        RECT 30.195 145.720 30.515 145.980 ;
        RECT 31.665 145.920 31.805 146.075 ;
        RECT 33.875 146.060 34.195 146.120 ;
        RECT 35.715 146.260 36.035 146.320 ;
        RECT 50.985 146.305 51.125 146.460 ;
        RECT 60.095 146.400 60.415 146.460 ;
        RECT 62.855 146.400 63.175 146.460 ;
        RECT 100.545 146.600 100.835 146.645 ;
        RECT 103.325 146.600 103.615 146.645 ;
        RECT 105.185 146.600 105.475 146.645 ;
        RECT 100.545 146.460 105.475 146.600 ;
        RECT 100.545 146.415 100.835 146.460 ;
        RECT 103.325 146.415 103.615 146.460 ;
        RECT 105.185 146.415 105.475 146.460 ;
        RECT 36.190 146.260 36.480 146.305 ;
        RECT 35.715 146.120 36.480 146.260 ;
        RECT 35.715 146.060 36.035 146.120 ;
        RECT 36.190 146.075 36.480 146.120 ;
        RECT 50.910 146.075 51.200 146.305 ;
        RECT 101.495 146.260 101.815 146.320 ;
        RECT 79.045 146.120 81.945 146.260 ;
        RECT 33.415 145.920 33.735 145.980 ;
        RECT 35.805 145.920 35.945 146.060 ;
        RECT 31.665 145.780 35.945 145.920 ;
        RECT 33.415 145.720 33.735 145.780 ;
        RECT 37.555 145.720 37.875 145.980 ;
        RECT 43.995 145.720 44.315 145.980 ;
        RECT 44.455 145.720 44.775 145.980 ;
        RECT 55.035 145.920 55.355 145.980 ;
        RECT 79.045 145.965 79.185 146.120 ;
        RECT 81.805 145.965 81.945 146.120 ;
        RECT 86.375 146.120 101.815 146.260 ;
        RECT 55.510 145.920 55.800 145.965 ;
        RECT 55.035 145.780 55.800 145.920 ;
        RECT 55.035 145.720 55.355 145.780 ;
        RECT 55.510 145.735 55.800 145.780 ;
        RECT 78.970 145.735 79.260 145.965 ;
        RECT 80.350 145.735 80.640 145.965 ;
        RECT 81.730 145.920 82.020 145.965 ;
        RECT 82.635 145.920 82.955 145.980 ;
        RECT 86.375 145.920 86.515 146.120 ;
        RECT 101.495 146.060 101.815 146.120 ;
        RECT 81.730 145.780 82.955 145.920 ;
        RECT 81.730 145.735 82.020 145.780 ;
        RECT 61.015 145.380 61.335 145.640 ;
        RECT 69.755 145.380 70.075 145.640 ;
        RECT 80.425 145.580 80.565 145.735 ;
        RECT 82.635 145.720 82.955 145.780 ;
        RECT 83.185 145.780 86.515 145.920 ;
        RECT 83.185 145.580 83.325 145.780 ;
        RECT 88.615 145.720 88.935 145.980 ;
        RECT 89.535 145.720 89.855 145.980 ;
        RECT 90.930 145.735 91.220 145.965 ;
        RECT 91.375 145.920 91.695 145.980 ;
        RECT 92.310 145.920 92.600 145.965 ;
        RECT 91.375 145.780 92.600 145.920 ;
        RECT 80.425 145.440 83.325 145.580 ;
        RECT 85.855 145.580 86.175 145.640 ;
        RECT 91.005 145.580 91.145 145.735 ;
        RECT 91.375 145.720 91.695 145.780 ;
        RECT 92.310 145.735 92.600 145.780 ;
        RECT 100.545 145.920 100.835 145.965 ;
        RECT 100.545 145.780 103.080 145.920 ;
        RECT 100.545 145.735 100.835 145.780 ;
        RECT 85.855 145.440 91.145 145.580 ;
        RECT 91.850 145.580 92.140 145.625 ;
        RECT 93.675 145.580 93.995 145.640 ;
        RECT 91.850 145.440 93.995 145.580 ;
        RECT 85.855 145.380 86.175 145.440 ;
        RECT 91.850 145.395 92.140 145.440 ;
        RECT 93.675 145.380 93.995 145.440 ;
        RECT 98.685 145.580 98.975 145.625 ;
        RECT 100.115 145.580 100.435 145.640 ;
        RECT 102.865 145.625 103.080 145.780 ;
        RECT 103.795 145.720 104.115 145.980 ;
        RECT 105.650 145.920 105.940 145.965 ;
        RECT 106.095 145.920 106.415 145.980 ;
        RECT 105.650 145.780 106.415 145.920 ;
        RECT 105.650 145.735 105.940 145.780 ;
        RECT 106.095 145.720 106.415 145.780 ;
        RECT 107.030 145.920 107.320 145.965 ;
        RECT 107.475 145.920 107.795 145.980 ;
        RECT 107.030 145.780 107.795 145.920 ;
        RECT 107.030 145.735 107.320 145.780 ;
        RECT 107.475 145.720 107.795 145.780 ;
        RECT 101.945 145.580 102.235 145.625 ;
        RECT 98.685 145.440 102.235 145.580 ;
        RECT 98.685 145.395 98.975 145.440 ;
        RECT 100.115 145.380 100.435 145.440 ;
        RECT 101.945 145.395 102.235 145.440 ;
        RECT 102.865 145.580 103.155 145.625 ;
        RECT 104.725 145.580 105.015 145.625 ;
        RECT 102.865 145.440 105.015 145.580 ;
        RECT 102.865 145.395 103.155 145.440 ;
        RECT 104.725 145.395 105.015 145.440 ;
        RECT 32.495 145.240 32.815 145.300 ;
        RECT 37.110 145.240 37.400 145.285 ;
        RECT 32.495 145.100 37.400 145.240 ;
        RECT 32.495 145.040 32.815 145.100 ;
        RECT 37.110 145.055 37.400 145.100 ;
        RECT 50.895 145.240 51.215 145.300 ;
        RECT 51.370 145.240 51.660 145.285 ;
        RECT 50.895 145.100 51.660 145.240 ;
        RECT 50.895 145.040 51.215 145.100 ;
        RECT 51.370 145.055 51.660 145.100 ;
        RECT 51.815 145.040 52.135 145.300 ;
        RECT 52.275 145.240 52.595 145.300 ;
        RECT 53.670 145.240 53.960 145.285 ;
        RECT 52.275 145.100 53.960 145.240 ;
        RECT 52.275 145.040 52.595 145.100 ;
        RECT 53.670 145.055 53.960 145.100 ;
        RECT 79.430 145.240 79.720 145.285 ;
        RECT 81.715 145.240 82.035 145.300 ;
        RECT 79.430 145.100 82.035 145.240 ;
        RECT 79.430 145.055 79.720 145.100 ;
        RECT 81.715 145.040 82.035 145.100 ;
        RECT 94.595 145.240 94.915 145.300 ;
        RECT 96.680 145.240 96.970 145.285 ;
        RECT 94.595 145.100 96.970 145.240 ;
        RECT 94.595 145.040 94.915 145.100 ;
        RECT 96.680 145.055 96.970 145.100 ;
        RECT 97.355 145.240 97.675 145.300 ;
        RECT 105.175 145.240 105.495 145.300 ;
        RECT 97.355 145.100 105.495 145.240 ;
        RECT 97.355 145.040 97.675 145.100 ;
        RECT 105.175 145.040 105.495 145.100 ;
        RECT 106.555 145.040 106.875 145.300 ;
        RECT 18.165 144.420 112.465 144.900 ;
        RECT 31.590 144.220 31.880 144.265 ;
        RECT 32.495 144.220 32.815 144.280 ;
        RECT 31.590 144.080 32.815 144.220 ;
        RECT 31.590 144.035 31.880 144.080 ;
        RECT 32.495 144.020 32.815 144.080 ;
        RECT 43.535 144.220 43.855 144.280 ;
        RECT 48.840 144.220 49.130 144.265 ;
        RECT 59.175 144.220 59.495 144.280 ;
        RECT 71.150 144.220 71.440 144.265 ;
        RECT 43.535 144.080 71.440 144.220 ;
        RECT 43.535 144.020 43.855 144.080 ;
        RECT 48.840 144.035 49.130 144.080 ;
        RECT 59.175 144.020 59.495 144.080 ;
        RECT 71.150 144.035 71.440 144.080 ;
        RECT 89.995 144.220 90.315 144.280 ;
        RECT 90.915 144.220 91.235 144.280 ;
        RECT 94.595 144.220 94.915 144.280 ;
        RECT 96.450 144.220 96.740 144.265 ;
        RECT 89.995 144.080 93.445 144.220 ;
        RECT 89.995 144.020 90.315 144.080 ;
        RECT 90.915 144.020 91.235 144.080 ;
        RECT 46.770 143.880 47.060 143.925 ;
        RECT 50.845 143.880 51.135 143.925 ;
        RECT 54.105 143.880 54.395 143.925 ;
        RECT 46.770 143.740 54.395 143.880 ;
        RECT 46.770 143.695 47.060 143.740 ;
        RECT 50.845 143.695 51.135 143.740 ;
        RECT 54.105 143.695 54.395 143.740 ;
        RECT 55.025 143.880 55.315 143.925 ;
        RECT 56.885 143.880 57.175 143.925 ;
        RECT 55.025 143.740 57.175 143.880 ;
        RECT 55.025 143.695 55.315 143.740 ;
        RECT 56.885 143.695 57.175 143.740 ;
        RECT 61.130 143.880 61.420 143.925 ;
        RECT 64.370 143.880 65.020 143.925 ;
        RECT 61.130 143.740 65.020 143.880 ;
        RECT 61.130 143.695 61.720 143.740 ;
        RECT 64.370 143.695 65.020 143.740 ;
        RECT 70.215 143.880 70.535 143.940 ;
        RECT 70.690 143.880 70.980 143.925 ;
        RECT 70.215 143.740 70.980 143.880 ;
        RECT 32.955 143.540 33.275 143.600 ;
        RECT 34.350 143.540 34.640 143.585 ;
        RECT 32.955 143.400 34.640 143.540 ;
        RECT 32.955 143.340 33.275 143.400 ;
        RECT 34.350 143.355 34.640 143.400 ;
        RECT 44.930 143.540 45.220 143.585 ;
        RECT 46.310 143.540 46.600 143.585 ;
        RECT 44.930 143.400 46.600 143.540 ;
        RECT 44.930 143.355 45.220 143.400 ;
        RECT 46.310 143.355 46.600 143.400 ;
        RECT 52.705 143.540 52.995 143.585 ;
        RECT 55.025 143.540 55.240 143.695 ;
        RECT 52.705 143.400 55.240 143.540 ;
        RECT 61.430 143.600 61.720 143.695 ;
        RECT 70.215 143.680 70.535 143.740 ;
        RECT 70.690 143.695 70.980 143.740 ;
        RECT 74.835 143.880 75.125 143.925 ;
        RECT 76.695 143.880 76.985 143.925 ;
        RECT 74.835 143.740 76.985 143.880 ;
        RECT 74.835 143.695 75.125 143.740 ;
        RECT 76.695 143.695 76.985 143.740 ;
        RECT 77.615 143.880 77.905 143.925 ;
        RECT 80.335 143.880 80.655 143.940 ;
        RECT 80.875 143.880 81.165 143.925 ;
        RECT 91.375 143.880 91.695 143.940 ;
        RECT 92.295 143.880 92.615 143.940 ;
        RECT 93.305 143.925 93.445 144.080 ;
        RECT 94.595 144.080 96.740 144.220 ;
        RECT 94.595 144.020 94.915 144.080 ;
        RECT 96.450 144.035 96.740 144.080 ;
        RECT 96.910 144.220 97.200 144.265 ;
        RECT 97.355 144.220 97.675 144.280 ;
        RECT 96.910 144.080 97.675 144.220 ;
        RECT 96.910 144.035 97.200 144.080 ;
        RECT 97.355 144.020 97.675 144.080 ;
        RECT 98.750 144.220 99.040 144.265 ;
        RECT 103.795 144.220 104.115 144.280 ;
        RECT 98.750 144.080 104.115 144.220 ;
        RECT 98.750 144.035 99.040 144.080 ;
        RECT 103.795 144.020 104.115 144.080 ;
        RECT 105.175 144.220 105.495 144.280 ;
        RECT 108.640 144.220 108.930 144.265 ;
        RECT 105.175 144.080 108.930 144.220 ;
        RECT 105.175 144.020 105.495 144.080 ;
        RECT 108.640 144.035 108.930 144.080 ;
        RECT 77.615 143.740 81.165 143.880 ;
        RECT 77.615 143.695 77.905 143.740 ;
        RECT 52.705 143.355 52.995 143.400 ;
        RECT 61.430 143.380 61.795 143.600 ;
        RECT 45.390 142.520 45.680 142.565 ;
        RECT 45.835 142.520 46.155 142.580 ;
        RECT 45.390 142.380 46.155 142.520 ;
        RECT 46.385 142.520 46.525 143.355 ;
        RECT 61.475 143.340 61.795 143.380 ;
        RECT 62.510 143.540 62.800 143.585 ;
        RECT 66.090 143.540 66.380 143.585 ;
        RECT 67.925 143.540 68.215 143.585 ;
        RECT 62.510 143.400 68.215 143.540 ;
        RECT 62.510 143.355 62.800 143.400 ;
        RECT 66.090 143.355 66.380 143.400 ;
        RECT 67.925 143.355 68.215 143.400 ;
        RECT 68.390 143.540 68.680 143.585 ;
        RECT 75.750 143.540 76.040 143.585 ;
        RECT 76.195 143.540 76.515 143.600 ;
        RECT 68.390 143.400 74.125 143.540 ;
        RECT 68.390 143.355 68.680 143.400 ;
        RECT 54.575 143.200 54.895 143.260 ;
        RECT 55.970 143.200 56.260 143.245 ;
        RECT 54.575 143.060 56.260 143.200 ;
        RECT 54.575 143.000 54.895 143.060 ;
        RECT 55.970 143.015 56.260 143.060 ;
        RECT 57.810 143.200 58.100 143.245 ;
        RECT 58.255 143.200 58.575 143.260 ;
        RECT 57.810 143.060 58.575 143.200 ;
        RECT 57.810 143.015 58.100 143.060 ;
        RECT 58.255 143.000 58.575 143.060 ;
        RECT 59.635 143.000 59.955 143.260 ;
        RECT 66.535 143.200 66.855 143.260 ;
        RECT 67.010 143.200 67.300 143.245 ;
        RECT 66.535 143.060 67.300 143.200 ;
        RECT 66.535 143.000 66.855 143.060 ;
        RECT 67.010 143.015 67.300 143.060 ;
        RECT 70.230 143.200 70.520 143.245 ;
        RECT 71.595 143.200 71.915 143.260 ;
        RECT 73.985 143.245 74.125 143.400 ;
        RECT 75.750 143.400 76.515 143.540 ;
        RECT 76.770 143.540 76.985 143.695 ;
        RECT 80.335 143.680 80.655 143.740 ;
        RECT 80.875 143.695 81.165 143.740 ;
        RECT 84.565 143.740 92.615 143.880 ;
        RECT 79.015 143.540 79.305 143.585 ;
        RECT 76.770 143.400 79.305 143.540 ;
        RECT 75.750 143.355 76.040 143.400 ;
        RECT 76.195 143.340 76.515 143.400 ;
        RECT 79.015 143.355 79.305 143.400 ;
        RECT 83.095 143.540 83.415 143.600 ;
        RECT 84.565 143.585 84.705 143.740 ;
        RECT 84.490 143.540 84.780 143.585 ;
        RECT 83.095 143.400 84.780 143.540 ;
        RECT 83.095 143.340 83.415 143.400 ;
        RECT 84.490 143.355 84.780 143.400 ;
        RECT 85.855 143.340 86.175 143.600 ;
        RECT 86.790 143.355 87.080 143.585 ;
        RECT 70.230 143.060 71.915 143.200 ;
        RECT 70.230 143.015 70.520 143.060 ;
        RECT 71.595 143.000 71.915 143.060 ;
        RECT 73.910 143.200 74.200 143.245 ;
        RECT 75.275 143.200 75.595 143.260 ;
        RECT 73.910 143.060 75.595 143.200 ;
        RECT 73.910 143.015 74.200 143.060 ;
        RECT 75.275 143.000 75.595 143.060 ;
        RECT 76.655 143.200 76.975 143.260 ;
        RECT 86.865 143.200 87.005 143.355 ;
        RECT 88.155 143.340 88.475 143.600 ;
        RECT 89.165 143.585 89.305 143.740 ;
        RECT 91.375 143.680 91.695 143.740 ;
        RECT 92.295 143.680 92.615 143.740 ;
        RECT 93.230 143.880 93.520 143.925 ;
        RECT 94.135 143.880 94.455 143.940 ;
        RECT 106.555 143.925 106.875 143.940 ;
        RECT 93.230 143.740 94.455 143.880 ;
        RECT 93.230 143.695 93.520 143.740 ;
        RECT 94.135 143.680 94.455 143.740 ;
        RECT 100.595 143.880 100.885 143.925 ;
        RECT 102.455 143.880 102.745 143.925 ;
        RECT 100.595 143.740 102.745 143.880 ;
        RECT 100.595 143.695 100.885 143.740 ;
        RECT 102.455 143.695 102.745 143.740 ;
        RECT 103.375 143.880 103.665 143.925 ;
        RECT 106.555 143.880 106.925 143.925 ;
        RECT 103.375 143.740 106.925 143.880 ;
        RECT 103.375 143.695 103.665 143.740 ;
        RECT 106.555 143.695 106.925 143.740 ;
        RECT 89.090 143.355 89.380 143.585 ;
        RECT 90.010 143.355 90.300 143.585 ;
        RECT 90.455 143.540 90.775 143.600 ;
        RECT 91.850 143.540 92.140 143.585 ;
        RECT 90.455 143.400 92.140 143.540 ;
        RECT 76.655 143.060 87.005 143.200 ;
        RECT 90.085 143.200 90.225 143.355 ;
        RECT 90.455 143.340 90.775 143.400 ;
        RECT 91.850 143.355 92.140 143.400 ;
        RECT 94.610 143.355 94.900 143.585 ;
        RECT 99.195 143.540 99.515 143.600 ;
        RECT 101.510 143.540 101.800 143.585 ;
        RECT 99.195 143.400 101.800 143.540 ;
        RECT 102.530 143.540 102.745 143.695 ;
        RECT 106.555 143.680 106.875 143.695 ;
        RECT 104.775 143.540 105.065 143.585 ;
        RECT 102.530 143.400 105.065 143.540 ;
        RECT 94.150 143.200 94.440 143.245 ;
        RECT 90.085 143.060 94.440 143.200 ;
        RECT 76.655 143.000 76.975 143.060 ;
        RECT 52.705 142.860 52.995 142.905 ;
        RECT 55.485 142.860 55.775 142.905 ;
        RECT 57.345 142.860 57.635 142.905 ;
        RECT 59.725 142.860 59.865 143.000 ;
        RECT 52.705 142.720 57.635 142.860 ;
        RECT 52.705 142.675 52.995 142.720 ;
        RECT 55.485 142.675 55.775 142.720 ;
        RECT 57.345 142.675 57.635 142.720 ;
        RECT 58.345 142.720 59.865 142.860 ;
        RECT 62.510 142.860 62.800 142.905 ;
        RECT 65.630 142.860 65.920 142.905 ;
        RECT 67.520 142.860 67.810 142.905 ;
        RECT 62.510 142.720 67.810 142.860 ;
        RECT 58.345 142.520 58.485 142.720 ;
        RECT 62.510 142.675 62.800 142.720 ;
        RECT 65.630 142.675 65.920 142.720 ;
        RECT 67.520 142.675 67.810 142.720 ;
        RECT 74.375 142.860 74.665 142.905 ;
        RECT 76.235 142.860 76.525 142.905 ;
        RECT 79.015 142.860 79.305 142.905 ;
        RECT 84.950 142.860 85.240 142.905 ;
        RECT 74.375 142.720 79.305 142.860 ;
        RECT 74.375 142.675 74.665 142.720 ;
        RECT 76.235 142.675 76.525 142.720 ;
        RECT 79.015 142.675 79.305 142.720 ;
        RECT 79.505 142.720 85.240 142.860 ;
        RECT 46.385 142.380 58.485 142.520 ;
        RECT 58.715 142.520 59.035 142.580 ;
        RECT 59.650 142.520 59.940 142.565 ;
        RECT 58.715 142.380 59.940 142.520 ;
        RECT 45.390 142.335 45.680 142.380 ;
        RECT 45.835 142.320 46.155 142.380 ;
        RECT 58.715 142.320 59.035 142.380 ;
        RECT 59.650 142.335 59.940 142.380 ;
        RECT 72.975 142.320 73.295 142.580 ;
        RECT 78.035 142.520 78.355 142.580 ;
        RECT 79.505 142.520 79.645 142.720 ;
        RECT 84.950 142.675 85.240 142.720 ;
        RECT 85.855 142.860 86.175 142.920 ;
        RECT 90.085 142.860 90.225 143.060 ;
        RECT 94.150 143.015 94.440 143.060 ;
        RECT 85.855 142.720 90.225 142.860 ;
        RECT 85.855 142.660 86.175 142.720 ;
        RECT 78.035 142.380 79.645 142.520 ;
        RECT 82.175 142.520 82.495 142.580 ;
        RECT 82.880 142.520 83.170 142.565 ;
        RECT 82.175 142.380 83.170 142.520 ;
        RECT 78.035 142.320 78.355 142.380 ;
        RECT 82.175 142.320 82.495 142.380 ;
        RECT 82.880 142.335 83.170 142.380 ;
        RECT 87.235 142.520 87.555 142.580 ;
        RECT 89.550 142.520 89.840 142.565 ;
        RECT 87.235 142.380 89.840 142.520 ;
        RECT 94.685 142.520 94.825 143.355 ;
        RECT 99.195 143.340 99.515 143.400 ;
        RECT 101.510 143.355 101.800 143.400 ;
        RECT 104.775 143.355 105.065 143.400 ;
        RECT 110.695 143.340 111.015 143.600 ;
        RECT 95.990 143.200 96.280 143.245 ;
        RECT 97.815 143.200 98.135 143.260 ;
        RECT 95.990 143.060 98.135 143.200 ;
        RECT 95.990 143.015 96.280 143.060 ;
        RECT 97.815 143.000 98.135 143.060 ;
        RECT 99.655 143.200 99.975 143.260 ;
        RECT 106.095 143.200 106.415 143.260 ;
        RECT 99.655 143.060 106.415 143.200 ;
        RECT 99.655 143.000 99.975 143.060 ;
        RECT 106.095 143.000 106.415 143.060 ;
        RECT 100.135 142.860 100.425 142.905 ;
        RECT 101.995 142.860 102.285 142.905 ;
        RECT 104.775 142.860 105.065 142.905 ;
        RECT 100.135 142.720 105.065 142.860 ;
        RECT 100.135 142.675 100.425 142.720 ;
        RECT 101.995 142.675 102.285 142.720 ;
        RECT 104.775 142.675 105.065 142.720 ;
        RECT 109.790 142.520 110.080 142.565 ;
        RECT 94.685 142.380 110.080 142.520 ;
        RECT 87.235 142.320 87.555 142.380 ;
        RECT 89.550 142.335 89.840 142.380 ;
        RECT 109.790 142.335 110.080 142.380 ;
        RECT 17.605 141.700 112.465 142.180 ;
        RECT 54.575 141.300 54.895 141.560 ;
        RECT 61.475 141.300 61.795 141.560 ;
        RECT 66.090 141.500 66.380 141.545 ;
        RECT 66.535 141.500 66.855 141.560 ;
        RECT 66.090 141.360 66.855 141.500 ;
        RECT 66.090 141.315 66.380 141.360 ;
        RECT 66.535 141.300 66.855 141.360 ;
        RECT 135.635 141.220 136.775 165.470 ;
        RECT 46.755 141.160 47.075 141.220 ;
        RECT 36.725 141.020 47.075 141.160 ;
        RECT 21.915 140.480 22.235 140.540 ;
        RECT 36.725 140.525 36.865 141.020 ;
        RECT 46.755 140.960 47.075 141.020 ;
        RECT 49.025 141.160 49.315 141.205 ;
        RECT 51.805 141.160 52.095 141.205 ;
        RECT 53.665 141.160 53.955 141.205 ;
        RECT 66.995 141.160 67.315 141.220 ;
        RECT 49.025 141.020 53.955 141.160 ;
        RECT 49.025 140.975 49.315 141.020 ;
        RECT 51.805 140.975 52.095 141.020 ;
        RECT 53.665 140.975 53.955 141.020 ;
        RECT 57.425 141.020 67.315 141.160 ;
        RECT 45.835 140.820 46.155 140.880 ;
        RECT 39.025 140.680 42.845 140.820 ;
        RECT 30.670 140.480 30.960 140.525 ;
        RECT 36.650 140.480 36.940 140.525 ;
        RECT 21.915 140.340 36.940 140.480 ;
        RECT 21.915 140.280 22.235 140.340 ;
        RECT 30.670 140.295 30.960 140.340 ;
        RECT 36.650 140.295 36.940 140.340 ;
        RECT 38.475 140.480 38.795 140.540 ;
        RECT 39.025 140.525 39.165 140.680 ;
        RECT 38.950 140.480 39.240 140.525 ;
        RECT 38.475 140.340 39.240 140.480 ;
        RECT 38.475 140.280 38.795 140.340 ;
        RECT 38.950 140.295 39.240 140.340 ;
        RECT 39.395 140.280 39.715 140.540 ;
        RECT 39.870 140.295 40.160 140.525 ;
        RECT 40.790 140.480 41.080 140.525 ;
        RECT 41.695 140.480 42.015 140.540 ;
        RECT 42.705 140.525 42.845 140.680 ;
        RECT 45.835 140.680 52.045 140.820 ;
        RECT 45.835 140.620 46.155 140.680 ;
        RECT 40.790 140.340 42.015 140.480 ;
        RECT 40.790 140.295 41.080 140.340 ;
        RECT 34.335 140.140 34.655 140.200 ;
        RECT 37.570 140.140 37.860 140.185 ;
        RECT 34.335 140.000 37.860 140.140 ;
        RECT 39.945 140.140 40.085 140.295 ;
        RECT 41.695 140.280 42.015 140.340 ;
        RECT 42.630 140.295 42.920 140.525 ;
        RECT 43.075 140.280 43.395 140.540 ;
        RECT 43.535 140.280 43.855 140.540 ;
        RECT 44.455 140.280 44.775 140.540 ;
        RECT 49.025 140.480 49.315 140.525 ;
        RECT 51.905 140.480 52.045 140.680 ;
        RECT 52.275 140.620 52.595 140.880 ;
        RECT 52.735 140.820 53.055 140.880 ;
        RECT 57.425 140.820 57.565 141.020 ;
        RECT 66.995 140.960 67.315 141.020 ;
        RECT 72.025 141.160 72.315 141.205 ;
        RECT 74.805 141.160 75.095 141.205 ;
        RECT 76.665 141.160 76.955 141.205 ;
        RECT 72.025 141.020 76.955 141.160 ;
        RECT 72.025 140.975 72.315 141.020 ;
        RECT 74.805 140.975 75.095 141.020 ;
        RECT 76.665 140.975 76.955 141.020 ;
        RECT 80.335 141.160 80.655 141.220 ;
        RECT 82.190 141.160 82.480 141.205 ;
        RECT 80.335 141.020 82.480 141.160 ;
        RECT 80.335 140.960 80.655 141.020 ;
        RECT 82.190 140.975 82.480 141.020 ;
        RECT 86.315 141.160 86.635 141.220 ;
        RECT 88.630 141.160 88.920 141.205 ;
        RECT 94.595 141.160 94.915 141.220 ;
        RECT 86.315 141.020 88.920 141.160 ;
        RECT 86.315 140.960 86.635 141.020 ;
        RECT 88.630 140.975 88.920 141.020 ;
        RECT 91.465 141.020 94.915 141.160 ;
        RECT 52.735 140.680 57.565 140.820 ;
        RECT 57.810 140.820 58.100 140.865 ;
        RECT 60.095 140.820 60.415 140.880 ;
        RECT 63.330 140.820 63.620 140.865 ;
        RECT 57.810 140.680 63.620 140.820 ;
        RECT 52.735 140.620 53.055 140.680 ;
        RECT 57.810 140.635 58.100 140.680 ;
        RECT 60.095 140.620 60.415 140.680 ;
        RECT 63.330 140.635 63.620 140.680 ;
        RECT 68.160 140.820 68.450 140.865 ;
        RECT 70.215 140.820 70.535 140.880 ;
        RECT 68.160 140.680 70.535 140.820 ;
        RECT 68.160 140.635 68.450 140.680 ;
        RECT 52.825 140.480 52.965 140.620 ;
        RECT 49.025 140.340 51.560 140.480 ;
        RECT 51.905 140.340 52.965 140.480 ;
        RECT 49.025 140.295 49.315 140.340 ;
        RECT 45.160 140.140 45.450 140.185 ;
        RECT 46.295 140.140 46.615 140.200 ;
        RECT 51.345 140.185 51.560 140.340 ;
        RECT 54.130 140.295 54.420 140.525 ;
        RECT 56.890 140.480 57.180 140.525 ;
        RECT 59.175 140.480 59.495 140.540 ;
        RECT 56.890 140.340 59.495 140.480 ;
        RECT 56.890 140.295 57.180 140.340 ;
        RECT 47.165 140.140 47.455 140.185 ;
        RECT 50.425 140.140 50.715 140.185 ;
        RECT 39.945 140.000 46.065 140.140 ;
        RECT 34.335 139.940 34.655 140.000 ;
        RECT 37.570 139.955 37.860 140.000 ;
        RECT 45.160 139.955 45.450 140.000 ;
        RECT 30.195 139.600 30.515 139.860 ;
        RECT 36.190 139.800 36.480 139.845 ;
        RECT 36.635 139.800 36.955 139.860 ;
        RECT 36.190 139.660 36.955 139.800 ;
        RECT 36.190 139.615 36.480 139.660 ;
        RECT 36.635 139.600 36.955 139.660 ;
        RECT 40.775 139.800 41.095 139.860 ;
        RECT 41.250 139.800 41.540 139.845 ;
        RECT 40.775 139.660 41.540 139.800 ;
        RECT 45.925 139.800 46.065 140.000 ;
        RECT 46.295 140.000 50.715 140.140 ;
        RECT 46.295 139.940 46.615 140.000 ;
        RECT 47.165 139.955 47.455 140.000 ;
        RECT 50.425 139.955 50.715 140.000 ;
        RECT 51.345 140.140 51.635 140.185 ;
        RECT 53.205 140.140 53.495 140.185 ;
        RECT 51.345 140.000 53.495 140.140 ;
        RECT 54.205 140.140 54.345 140.295 ;
        RECT 59.175 140.280 59.495 140.340 ;
        RECT 59.635 140.480 59.955 140.540 ;
        RECT 61.030 140.480 61.320 140.525 ;
        RECT 59.635 140.340 61.320 140.480 ;
        RECT 63.405 140.480 63.545 140.635 ;
        RECT 70.215 140.620 70.535 140.680 ;
        RECT 71.595 140.620 71.915 140.880 ;
        RECT 72.975 140.820 73.295 140.880 ;
        RECT 75.290 140.820 75.580 140.865 ;
        RECT 85.855 140.820 86.175 140.880 ;
        RECT 86.790 140.820 87.080 140.865 ;
        RECT 72.975 140.680 75.580 140.820 ;
        RECT 72.975 140.620 73.295 140.680 ;
        RECT 75.290 140.635 75.580 140.680 ;
        RECT 84.565 140.680 87.080 140.820 ;
        RECT 71.685 140.480 71.825 140.620 ;
        RECT 63.405 140.340 71.825 140.480 ;
        RECT 72.025 140.480 72.315 140.525 ;
        RECT 75.735 140.480 76.055 140.540 ;
        RECT 77.130 140.480 77.420 140.525 ;
        RECT 72.025 140.340 74.560 140.480 ;
        RECT 59.635 140.280 59.955 140.340 ;
        RECT 61.030 140.295 61.320 140.340 ;
        RECT 72.025 140.295 72.315 140.340 ;
        RECT 58.255 140.140 58.575 140.200 ;
        RECT 54.205 140.000 58.575 140.140 ;
        RECT 51.345 139.955 51.635 140.000 ;
        RECT 53.205 139.955 53.495 140.000 ;
        RECT 58.255 139.940 58.575 140.000 ;
        RECT 70.165 140.140 70.455 140.185 ;
        RECT 72.515 140.140 72.835 140.200 ;
        RECT 74.345 140.185 74.560 140.340 ;
        RECT 75.735 140.340 77.420 140.480 ;
        RECT 75.735 140.280 76.055 140.340 ;
        RECT 77.130 140.295 77.420 140.340 ;
        RECT 78.495 140.280 78.815 140.540 ;
        RECT 82.635 140.280 82.955 140.540 ;
        RECT 84.565 140.525 84.705 140.680 ;
        RECT 85.855 140.620 86.175 140.680 ;
        RECT 86.790 140.635 87.080 140.680 ;
        RECT 89.995 140.820 90.315 140.880 ;
        RECT 89.995 140.680 90.685 140.820 ;
        RECT 89.995 140.620 90.315 140.680 ;
        RECT 83.110 140.295 83.400 140.525 ;
        RECT 84.490 140.295 84.780 140.525 ;
        RECT 84.950 140.295 85.240 140.525 ;
        RECT 73.425 140.140 73.715 140.185 ;
        RECT 70.165 140.000 73.715 140.140 ;
        RECT 70.165 139.955 70.455 140.000 ;
        RECT 72.515 139.940 72.835 140.000 ;
        RECT 73.425 139.955 73.715 140.000 ;
        RECT 74.345 140.140 74.635 140.185 ;
        RECT 76.205 140.140 76.495 140.185 ;
        RECT 74.345 140.000 76.495 140.140 ;
        RECT 74.345 139.955 74.635 140.000 ;
        RECT 76.205 139.955 76.495 140.000 ;
        RECT 81.270 140.140 81.560 140.185 ;
        RECT 83.185 140.140 83.325 140.295 ;
        RECT 81.270 140.000 83.325 140.140 ;
        RECT 83.555 140.140 83.875 140.200 ;
        RECT 84.030 140.140 84.320 140.185 ;
        RECT 83.555 140.000 84.320 140.140 ;
        RECT 85.025 140.140 85.165 140.295 ;
        RECT 87.695 140.280 88.015 140.540 ;
        RECT 90.545 140.525 90.685 140.680 ;
        RECT 90.470 140.295 90.760 140.525 ;
        RECT 90.915 140.280 91.235 140.540 ;
        RECT 91.465 140.525 91.605 141.020 ;
        RECT 94.595 140.960 94.915 141.020 ;
        RECT 96.450 141.160 96.740 141.205 ;
        RECT 99.195 141.160 99.515 141.220 ;
        RECT 96.450 141.020 99.515 141.160 ;
        RECT 96.450 140.975 96.740 141.020 ;
        RECT 99.195 140.960 99.515 141.020 ;
        RECT 101.005 141.160 101.295 141.205 ;
        RECT 103.785 141.160 104.075 141.205 ;
        RECT 105.645 141.160 105.935 141.205 ;
        RECT 101.005 141.020 105.935 141.160 ;
        RECT 101.005 140.975 101.295 141.020 ;
        RECT 103.785 140.975 104.075 141.020 ;
        RECT 105.645 140.975 105.935 141.020 ;
        RECT 93.690 140.635 93.980 140.865 ;
        RECT 94.150 140.820 94.440 140.865 ;
        RECT 97.355 140.820 97.675 140.880 ;
        RECT 94.150 140.680 97.675 140.820 ;
        RECT 94.150 140.635 94.440 140.680 ;
        RECT 91.390 140.295 91.680 140.525 ;
        RECT 92.295 140.280 92.615 140.540 ;
        RECT 93.765 140.480 93.905 140.635 ;
        RECT 97.355 140.620 97.675 140.680 ;
        RECT 98.735 140.820 99.055 140.880 ;
        RECT 104.270 140.820 104.560 140.865 ;
        RECT 98.735 140.680 104.560 140.820 ;
        RECT 98.735 140.620 99.055 140.680 ;
        RECT 104.270 140.635 104.560 140.680 ;
        RECT 106.095 140.620 106.415 140.880 ;
        RECT 95.055 140.480 95.375 140.540 ;
        RECT 97.815 140.480 98.135 140.540 ;
        RECT 93.765 140.340 98.135 140.480 ;
        RECT 95.055 140.280 95.375 140.340 ;
        RECT 97.815 140.280 98.135 140.340 ;
        RECT 101.005 140.480 101.295 140.525 ;
        RECT 101.005 140.340 103.540 140.480 ;
        RECT 101.005 140.295 101.295 140.340 ;
        RECT 89.995 140.140 90.315 140.200 ;
        RECT 91.005 140.140 91.145 140.280 ;
        RECT 85.025 140.000 89.305 140.140 ;
        RECT 81.270 139.955 81.560 140.000 ;
        RECT 83.555 139.940 83.875 140.000 ;
        RECT 84.030 139.955 84.320 140.000 ;
        RECT 50.895 139.800 51.215 139.860 ;
        RECT 56.430 139.800 56.720 139.845 ;
        RECT 45.925 139.660 56.720 139.800 ;
        RECT 40.775 139.600 41.095 139.660 ;
        RECT 41.250 139.615 41.540 139.660 ;
        RECT 50.895 139.600 51.215 139.660 ;
        RECT 56.430 139.615 56.720 139.660 ;
        RECT 59.175 139.600 59.495 139.860 ;
        RECT 61.935 139.800 62.255 139.860 ;
        RECT 63.790 139.800 64.080 139.845 ;
        RECT 61.935 139.660 64.080 139.800 ;
        RECT 61.935 139.600 62.255 139.660 ;
        RECT 63.790 139.615 64.080 139.660 ;
        RECT 64.250 139.800 64.540 139.845 ;
        RECT 64.695 139.800 65.015 139.860 ;
        RECT 78.495 139.800 78.815 139.860 ;
        RECT 64.250 139.660 78.815 139.800 ;
        RECT 64.250 139.615 64.540 139.660 ;
        RECT 64.695 139.600 65.015 139.660 ;
        RECT 78.495 139.600 78.815 139.660 ;
        RECT 85.870 139.800 86.160 139.845 ;
        RECT 86.775 139.800 87.095 139.860 ;
        RECT 89.165 139.845 89.305 140.000 ;
        RECT 89.995 140.000 91.145 140.140 ;
        RECT 99.145 140.140 99.435 140.185 ;
        RECT 100.115 140.140 100.435 140.200 ;
        RECT 103.325 140.185 103.540 140.340 ;
        RECT 135.580 140.230 136.830 141.220 ;
        RECT 102.405 140.140 102.695 140.185 ;
        RECT 99.145 140.000 102.695 140.140 ;
        RECT 89.995 139.940 90.315 140.000 ;
        RECT 99.145 139.955 99.435 140.000 ;
        RECT 100.115 139.940 100.435 140.000 ;
        RECT 102.405 139.955 102.695 140.000 ;
        RECT 103.325 140.140 103.615 140.185 ;
        RECT 105.185 140.140 105.475 140.185 ;
        RECT 135.635 140.155 136.775 140.230 ;
        RECT 103.325 140.000 105.475 140.140 ;
        RECT 103.325 139.955 103.615 140.000 ;
        RECT 105.185 139.955 105.475 140.000 ;
        RECT 85.870 139.660 87.095 139.800 ;
        RECT 85.870 139.615 86.160 139.660 ;
        RECT 86.775 139.600 87.095 139.660 ;
        RECT 89.090 139.800 89.380 139.845 ;
        RECT 90.915 139.800 91.235 139.860 ;
        RECT 89.090 139.660 91.235 139.800 ;
        RECT 89.090 139.615 89.380 139.660 ;
        RECT 90.915 139.600 91.235 139.660 ;
        RECT 94.595 139.800 94.915 139.860 ;
        RECT 97.140 139.800 97.430 139.845 ;
        RECT 94.595 139.660 97.430 139.800 ;
        RECT 94.595 139.600 94.915 139.660 ;
        RECT 97.140 139.615 97.430 139.660 ;
        RECT 18.165 138.980 112.465 139.460 ;
        RECT 132.510 139.190 135.210 140.010 ;
        RECT 143.370 139.390 144.510 223.840 ;
        RECT 137.240 139.380 144.510 139.390 ;
        RECT 136.210 139.190 144.510 139.380 ;
        RECT 32.510 138.780 32.800 138.825 ;
        RECT 32.955 138.780 33.275 138.840 ;
        RECT 32.510 138.640 33.275 138.780 ;
        RECT 32.510 138.595 32.800 138.640 ;
        RECT 32.955 138.580 33.275 138.640 ;
        RECT 33.875 138.780 34.195 138.840 ;
        RECT 38.935 138.780 39.255 138.840 ;
        RECT 33.875 138.640 39.255 138.780 ;
        RECT 33.875 138.580 34.195 138.640 ;
        RECT 38.935 138.580 39.255 138.640 ;
        RECT 39.395 138.780 39.715 138.840 ;
        RECT 43.075 138.780 43.395 138.840 ;
        RECT 43.995 138.780 44.315 138.840 ;
        RECT 45.835 138.780 46.155 138.840 ;
        RECT 39.395 138.640 46.155 138.780 ;
        RECT 39.395 138.580 39.715 138.640 ;
        RECT 43.075 138.580 43.395 138.640 ;
        RECT 43.995 138.580 44.315 138.640 ;
        RECT 45.835 138.580 46.155 138.640 ;
        RECT 49.300 138.780 49.590 138.825 ;
        RECT 51.815 138.780 52.135 138.840 ;
        RECT 59.175 138.780 59.495 138.840 ;
        RECT 49.300 138.640 52.135 138.780 ;
        RECT 49.300 138.595 49.590 138.640 ;
        RECT 51.815 138.580 52.135 138.640 ;
        RECT 55.125 138.640 59.495 138.780 ;
        RECT 27.430 138.440 28.080 138.485 ;
        RECT 30.195 138.440 30.515 138.500 ;
        RECT 31.030 138.440 31.320 138.485 ;
        RECT 27.430 138.300 31.320 138.440 ;
        RECT 27.430 138.255 28.080 138.300 ;
        RECT 30.195 138.240 30.515 138.300 ;
        RECT 30.730 138.255 31.320 138.300 ;
        RECT 34.450 138.440 34.740 138.485 ;
        RECT 36.635 138.440 36.955 138.500 ;
        RECT 37.690 138.440 38.340 138.485 ;
        RECT 34.450 138.300 38.340 138.440 ;
        RECT 34.450 138.255 35.040 138.300 ;
        RECT 21.470 138.100 21.760 138.145 ;
        RECT 21.915 138.100 22.235 138.160 ;
        RECT 21.470 137.960 22.235 138.100 ;
        RECT 21.470 137.915 21.760 137.960 ;
        RECT 21.915 137.900 22.235 137.960 ;
        RECT 24.235 138.100 24.525 138.145 ;
        RECT 26.070 138.100 26.360 138.145 ;
        RECT 29.650 138.100 29.940 138.145 ;
        RECT 24.235 137.960 29.940 138.100 ;
        RECT 24.235 137.915 24.525 137.960 ;
        RECT 26.070 137.915 26.360 137.960 ;
        RECT 29.650 137.915 29.940 137.960 ;
        RECT 30.730 137.940 31.020 138.255 ;
        RECT 34.750 137.940 35.040 138.255 ;
        RECT 36.635 138.240 36.955 138.300 ;
        RECT 37.690 138.255 38.340 138.300 ;
        RECT 41.695 138.440 42.015 138.500 ;
        RECT 42.615 138.440 42.935 138.500 ;
        RECT 44.455 138.440 44.775 138.500 ;
        RECT 51.305 138.440 51.595 138.485 ;
        RECT 54.565 138.440 54.855 138.485 ;
        RECT 55.125 138.440 55.265 138.640 ;
        RECT 59.175 138.580 59.495 138.640 ;
        RECT 72.070 138.780 72.360 138.825 ;
        RECT 72.515 138.780 72.835 138.840 ;
        RECT 72.070 138.640 72.835 138.780 ;
        RECT 72.070 138.595 72.360 138.640 ;
        RECT 72.515 138.580 72.835 138.640 ;
        RECT 76.195 138.780 76.515 138.840 ;
        RECT 77.590 138.780 77.880 138.825 ;
        RECT 76.195 138.640 77.880 138.780 ;
        RECT 76.195 138.580 76.515 138.640 ;
        RECT 77.590 138.595 77.880 138.640 ;
        RECT 78.495 138.780 78.815 138.840 ;
        RECT 79.660 138.780 79.950 138.825 ;
        RECT 78.495 138.640 79.950 138.780 ;
        RECT 78.495 138.580 78.815 138.640 ;
        RECT 79.660 138.595 79.950 138.640 ;
        RECT 83.555 138.780 83.875 138.840 ;
        RECT 95.055 138.780 95.375 138.840 ;
        RECT 83.555 138.640 95.375 138.780 ;
        RECT 83.555 138.580 83.875 138.640 ;
        RECT 95.055 138.580 95.375 138.640 ;
        RECT 98.735 138.580 99.055 138.840 ;
        RECT 132.510 138.530 144.510 139.190 ;
        RECT 41.695 138.300 47.445 138.440 ;
        RECT 41.695 138.240 42.015 138.300 ;
        RECT 42.615 138.240 42.935 138.300 ;
        RECT 44.455 138.240 44.775 138.300 ;
        RECT 35.830 138.100 36.120 138.145 ;
        RECT 39.410 138.100 39.700 138.145 ;
        RECT 41.245 138.100 41.535 138.145 ;
        RECT 35.830 137.960 41.535 138.100 ;
        RECT 35.830 137.915 36.120 137.960 ;
        RECT 39.410 137.915 39.700 137.960 ;
        RECT 41.245 137.915 41.535 137.960 ;
        RECT 43.535 137.900 43.855 138.160 ;
        RECT 45.375 137.900 45.695 138.160 ;
        RECT 45.835 137.900 46.155 138.160 ;
        RECT 47.305 138.145 47.445 138.300 ;
        RECT 51.305 138.300 55.265 138.440 ;
        RECT 55.485 138.440 55.775 138.485 ;
        RECT 57.345 138.440 57.635 138.485 ;
        RECT 55.485 138.300 57.635 138.440 ;
        RECT 51.305 138.255 51.595 138.300 ;
        RECT 54.565 138.255 54.855 138.300 ;
        RECT 55.485 138.255 55.775 138.300 ;
        RECT 57.345 138.255 57.635 138.300 ;
        RECT 66.995 138.440 67.315 138.500 ;
        RECT 81.715 138.485 82.035 138.500 ;
        RECT 75.750 138.440 76.040 138.485 ;
        RECT 66.995 138.300 69.985 138.440 ;
        RECT 46.310 137.915 46.600 138.145 ;
        RECT 47.230 137.915 47.520 138.145 ;
        RECT 53.165 138.100 53.455 138.145 ;
        RECT 55.485 138.100 55.700 138.255 ;
        RECT 66.995 138.240 67.315 138.300 ;
        RECT 53.165 137.960 55.700 138.100 ;
        RECT 55.955 138.100 56.275 138.160 ;
        RECT 58.715 138.100 59.035 138.160 ;
        RECT 55.955 137.960 59.035 138.100 ;
        RECT 53.165 137.915 53.455 137.960 ;
        RECT 23.770 137.760 24.060 137.805 ;
        RECT 41.710 137.760 42.000 137.805 ;
        RECT 23.770 137.620 42.000 137.760 ;
        RECT 46.385 137.760 46.525 137.915 ;
        RECT 55.955 137.900 56.275 137.960 ;
        RECT 58.715 137.900 59.035 137.960 ;
        RECT 59.175 138.100 59.495 138.160 ;
        RECT 60.095 138.100 60.415 138.160 ;
        RECT 59.175 137.960 60.415 138.100 ;
        RECT 59.175 137.900 59.495 137.960 ;
        RECT 60.095 137.900 60.415 137.960 ;
        RECT 63.775 137.900 64.095 138.160 ;
        RECT 64.235 137.900 64.555 138.160 ;
        RECT 64.695 137.900 65.015 138.160 ;
        RECT 65.630 138.100 65.920 138.145 ;
        RECT 66.075 138.100 66.395 138.160 ;
        RECT 69.845 138.145 69.985 138.300 ;
        RECT 70.765 138.300 76.040 138.440 ;
        RECT 65.630 137.960 66.395 138.100 ;
        RECT 65.630 137.915 65.920 137.960 ;
        RECT 66.075 137.900 66.395 137.960 ;
        RECT 69.310 137.915 69.600 138.145 ;
        RECT 69.770 137.915 70.060 138.145 ;
        RECT 70.215 138.100 70.535 138.160 ;
        RECT 70.765 138.100 70.905 138.300 ;
        RECT 75.750 138.255 76.040 138.300 ;
        RECT 81.665 138.440 82.035 138.485 ;
        RECT 84.925 138.440 85.215 138.485 ;
        RECT 81.665 138.300 85.215 138.440 ;
        RECT 81.665 138.255 82.035 138.300 ;
        RECT 84.925 138.255 85.215 138.300 ;
        RECT 85.845 138.440 86.135 138.485 ;
        RECT 87.705 138.440 87.995 138.485 ;
        RECT 96.910 138.440 97.200 138.485 ;
        RECT 85.845 138.300 87.995 138.440 ;
        RECT 85.845 138.255 86.135 138.300 ;
        RECT 87.705 138.255 87.995 138.300 ;
        RECT 90.085 138.300 97.200 138.440 ;
        RECT 81.715 138.240 82.035 138.255 ;
        RECT 70.215 137.960 70.905 138.100 ;
        RECT 55.035 137.760 55.355 137.820 ;
        RECT 46.385 137.620 55.355 137.760 ;
        RECT 23.770 137.575 24.060 137.620 ;
        RECT 34.885 137.480 35.025 137.620 ;
        RECT 41.710 137.575 42.000 137.620 ;
        RECT 55.035 137.560 55.355 137.620 ;
        RECT 55.495 137.760 55.815 137.820 ;
        RECT 56.430 137.760 56.720 137.805 ;
        RECT 55.495 137.620 56.720 137.760 ;
        RECT 55.495 137.560 55.815 137.620 ;
        RECT 56.430 137.575 56.720 137.620 ;
        RECT 58.255 137.560 58.575 137.820 ;
        RECT 69.385 137.760 69.525 137.915 ;
        RECT 70.215 137.900 70.535 137.960 ;
        RECT 71.150 137.915 71.440 138.145 ;
        RECT 72.055 138.100 72.375 138.160 ;
        RECT 72.530 138.100 72.820 138.145 ;
        RECT 82.635 138.100 82.955 138.160 ;
        RECT 72.055 137.960 82.955 138.100 ;
        RECT 59.725 137.620 69.525 137.760 ;
        RECT 24.640 137.420 24.930 137.465 ;
        RECT 26.530 137.420 26.820 137.465 ;
        RECT 29.650 137.420 29.940 137.465 ;
        RECT 24.640 137.280 29.940 137.420 ;
        RECT 24.640 137.235 24.930 137.280 ;
        RECT 26.530 137.235 26.820 137.280 ;
        RECT 29.650 137.235 29.940 137.280 ;
        RECT 34.795 137.220 35.115 137.480 ;
        RECT 35.830 137.420 36.120 137.465 ;
        RECT 38.950 137.420 39.240 137.465 ;
        RECT 40.840 137.420 41.130 137.465 ;
        RECT 35.830 137.280 41.130 137.420 ;
        RECT 35.830 137.235 36.120 137.280 ;
        RECT 38.950 137.235 39.240 137.280 ;
        RECT 40.840 137.235 41.130 137.280 ;
        RECT 53.165 137.420 53.455 137.465 ;
        RECT 55.945 137.420 56.235 137.465 ;
        RECT 57.805 137.420 58.095 137.465 ;
        RECT 53.165 137.280 58.095 137.420 ;
        RECT 53.165 137.235 53.455 137.280 ;
        RECT 55.945 137.235 56.235 137.280 ;
        RECT 57.805 137.235 58.095 137.280 ;
        RECT 20.995 136.880 21.315 137.140 ;
        RECT 23.295 137.080 23.615 137.140 ;
        RECT 25.060 137.080 25.350 137.125 ;
        RECT 23.295 136.940 25.350 137.080 ;
        RECT 23.295 136.880 23.615 136.940 ;
        RECT 25.060 136.895 25.350 136.940 ;
        RECT 32.495 137.080 32.815 137.140 ;
        RECT 32.970 137.080 33.260 137.125 ;
        RECT 32.495 136.940 33.260 137.080 ;
        RECT 32.495 136.880 32.815 136.940 ;
        RECT 32.970 136.895 33.260 136.940 ;
        RECT 40.425 137.080 40.715 137.125 ;
        RECT 41.235 137.080 41.555 137.140 ;
        RECT 40.425 136.940 41.555 137.080 ;
        RECT 40.425 136.895 40.715 136.940 ;
        RECT 41.235 136.880 41.555 136.940 ;
        RECT 42.615 136.880 42.935 137.140 ;
        RECT 43.075 137.080 43.395 137.140 ;
        RECT 44.010 137.080 44.300 137.125 ;
        RECT 43.075 136.940 44.300 137.080 ;
        RECT 43.075 136.880 43.395 136.940 ;
        RECT 44.010 136.895 44.300 136.940 ;
        RECT 54.575 137.080 54.895 137.140 ;
        RECT 59.725 137.080 59.865 137.620 ;
        RECT 61.935 137.220 62.255 137.480 ;
        RECT 66.535 137.420 66.855 137.480 ;
        RECT 71.225 137.420 71.365 137.915 ;
        RECT 72.055 137.900 72.375 137.960 ;
        RECT 72.530 137.915 72.820 137.960 ;
        RECT 82.635 137.900 82.955 137.960 ;
        RECT 83.525 138.100 83.815 138.145 ;
        RECT 85.845 138.100 86.060 138.255 ;
        RECT 83.525 137.960 86.060 138.100 ;
        RECT 83.525 137.915 83.815 137.960 ;
        RECT 86.775 137.900 87.095 138.160 ;
        RECT 90.085 138.100 90.225 138.300 ;
        RECT 87.325 137.960 90.225 138.100 ;
        RECT 71.595 137.760 71.915 137.820 ;
        RECT 74.355 137.760 74.675 137.820 ;
        RECT 71.595 137.620 74.675 137.760 ;
        RECT 71.595 137.560 71.915 137.620 ;
        RECT 74.355 137.560 74.675 137.620 ;
        RECT 75.290 137.760 75.580 137.805 ;
        RECT 82.175 137.760 82.495 137.820 ;
        RECT 87.325 137.760 87.465 137.960 ;
        RECT 90.455 137.900 90.775 138.160 ;
        RECT 91.465 138.145 91.605 138.300 ;
        RECT 96.910 138.255 97.200 138.300 ;
        RECT 104.250 138.440 104.900 138.485 ;
        RECT 107.015 138.440 107.335 138.500 ;
        RECT 107.850 138.440 108.140 138.485 ;
        RECT 104.250 138.300 108.140 138.440 ;
        RECT 104.250 138.255 104.900 138.300 ;
        RECT 107.015 138.240 107.335 138.300 ;
        RECT 107.550 138.255 108.140 138.300 ;
        RECT 90.930 137.915 91.220 138.145 ;
        RECT 91.390 137.915 91.680 138.145 ;
        RECT 91.835 138.100 92.155 138.160 ;
        RECT 92.310 138.100 92.600 138.145 ;
        RECT 91.835 137.960 92.600 138.100 ;
        RECT 75.290 137.620 87.465 137.760 ;
        RECT 88.630 137.760 88.920 137.805 ;
        RECT 89.075 137.760 89.395 137.820 ;
        RECT 91.005 137.760 91.145 137.915 ;
        RECT 91.835 137.900 92.155 137.960 ;
        RECT 92.310 137.915 92.600 137.960 ;
        RECT 99.655 138.100 99.975 138.160 ;
        RECT 100.590 138.100 100.880 138.145 ;
        RECT 99.655 137.960 100.880 138.100 ;
        RECT 99.655 137.900 99.975 137.960 ;
        RECT 100.590 137.915 100.880 137.960 ;
        RECT 101.055 138.100 101.345 138.145 ;
        RECT 102.890 138.100 103.180 138.145 ;
        RECT 106.470 138.100 106.760 138.145 ;
        RECT 101.055 137.960 106.760 138.100 ;
        RECT 101.055 137.915 101.345 137.960 ;
        RECT 102.890 137.915 103.180 137.960 ;
        RECT 106.470 137.915 106.760 137.960 ;
        RECT 107.550 137.940 107.840 138.255 ;
        RECT 110.695 138.240 111.015 138.500 ;
        RECT 132.510 138.190 135.210 138.530 ;
        RECT 136.210 138.250 144.510 138.530 ;
        RECT 136.210 138.240 138.350 138.250 ;
        RECT 88.630 137.620 89.395 137.760 ;
        RECT 75.290 137.575 75.580 137.620 ;
        RECT 82.175 137.560 82.495 137.620 ;
        RECT 88.630 137.575 88.920 137.620 ;
        RECT 89.075 137.560 89.395 137.620 ;
        RECT 90.545 137.620 91.145 137.760 ;
        RECT 72.975 137.420 73.295 137.480 ;
        RECT 82.635 137.420 82.955 137.480 ;
        RECT 66.535 137.280 82.955 137.420 ;
        RECT 66.535 137.220 66.855 137.280 ;
        RECT 72.975 137.220 73.295 137.280 ;
        RECT 82.635 137.220 82.955 137.280 ;
        RECT 83.525 137.420 83.815 137.465 ;
        RECT 86.305 137.420 86.595 137.465 ;
        RECT 88.165 137.420 88.455 137.465 ;
        RECT 83.525 137.280 88.455 137.420 ;
        RECT 83.525 137.235 83.815 137.280 ;
        RECT 86.305 137.235 86.595 137.280 ;
        RECT 88.165 137.235 88.455 137.280 ;
        RECT 89.995 137.420 90.315 137.480 ;
        RECT 90.545 137.420 90.685 137.620 ;
        RECT 95.975 137.560 96.295 137.820 ;
        RECT 96.450 137.575 96.740 137.805 ;
        RECT 89.995 137.280 90.685 137.420 ;
        RECT 91.835 137.420 92.155 137.480 ;
        RECT 94.595 137.420 94.915 137.480 ;
        RECT 96.525 137.420 96.665 137.575 ;
        RECT 91.835 137.280 96.665 137.420 ;
        RECT 101.460 137.420 101.750 137.465 ;
        RECT 103.350 137.420 103.640 137.465 ;
        RECT 106.470 137.420 106.760 137.465 ;
        RECT 101.460 137.280 106.760 137.420 ;
        RECT 89.995 137.220 90.315 137.280 ;
        RECT 91.835 137.220 92.155 137.280 ;
        RECT 94.595 137.220 94.915 137.280 ;
        RECT 101.460 137.235 101.750 137.280 ;
        RECT 103.350 137.235 103.640 137.280 ;
        RECT 106.470 137.235 106.760 137.280 ;
        RECT 54.575 136.940 59.865 137.080 ;
        RECT 60.095 137.080 60.415 137.140 ;
        RECT 62.410 137.080 62.700 137.125 ;
        RECT 60.095 136.940 62.700 137.080 ;
        RECT 54.575 136.880 54.895 136.940 ;
        RECT 60.095 136.880 60.415 136.940 ;
        RECT 62.410 136.895 62.700 136.940 ;
        RECT 65.155 137.080 65.475 137.140 ;
        RECT 67.930 137.080 68.220 137.125 ;
        RECT 65.155 136.940 68.220 137.080 ;
        RECT 65.155 136.880 65.475 136.940 ;
        RECT 67.930 136.895 68.220 136.940 ;
        RECT 80.335 137.080 80.655 137.140 ;
        RECT 89.090 137.080 89.380 137.125 ;
        RECT 80.335 136.940 89.380 137.080 ;
        RECT 80.335 136.880 80.655 136.940 ;
        RECT 89.090 136.895 89.380 136.940 ;
        RECT 90.455 137.080 90.775 137.140 ;
        RECT 101.880 137.080 102.170 137.125 ;
        RECT 90.455 136.940 102.170 137.080 ;
        RECT 90.455 136.880 90.775 136.940 ;
        RECT 101.880 136.895 102.170 136.940 ;
        RECT 17.605 136.260 112.465 136.740 ;
        RECT 23.295 135.860 23.615 136.120 ;
        RECT 25.135 136.060 25.455 136.120 ;
        RECT 37.095 136.060 37.415 136.120 ;
        RECT 25.135 135.920 37.415 136.060 ;
        RECT 25.135 135.860 25.455 135.920 ;
        RECT 37.095 135.860 37.415 135.920 ;
        RECT 41.235 135.860 41.555 136.120 ;
        RECT 45.375 136.060 45.695 136.120 ;
        RECT 54.575 136.060 54.895 136.120 ;
        RECT 43.625 135.920 54.895 136.060 ;
        RECT 30.670 135.720 30.960 135.765 ;
        RECT 35.255 135.720 35.575 135.780 ;
        RECT 26.605 135.580 30.960 135.720 ;
        RECT 26.605 135.425 26.745 135.580 ;
        RECT 30.670 135.535 30.960 135.580 ;
        RECT 33.505 135.580 35.575 135.720 ;
        RECT 33.505 135.440 33.645 135.580 ;
        RECT 35.255 135.520 35.575 135.580 ;
        RECT 26.530 135.195 26.820 135.425 ;
        RECT 27.450 135.380 27.740 135.425 ;
        RECT 32.495 135.380 32.815 135.440 ;
        RECT 27.450 135.240 32.815 135.380 ;
        RECT 27.450 135.195 27.740 135.240 ;
        RECT 32.495 135.180 32.815 135.240 ;
        RECT 33.415 135.180 33.735 135.440 ;
        RECT 37.555 135.380 37.875 135.440 ;
        RECT 34.425 135.240 37.875 135.380 ;
        RECT 22.390 135.040 22.680 135.085 ;
        RECT 24.215 135.040 24.535 135.100 ;
        RECT 30.655 135.040 30.975 135.100 ;
        RECT 22.390 134.900 30.975 135.040 ;
        RECT 22.390 134.855 22.680 134.900 ;
        RECT 24.215 134.840 24.535 134.900 ;
        RECT 30.655 134.840 30.975 134.900 ;
        RECT 32.955 135.040 33.275 135.100 ;
        RECT 34.425 135.040 34.565 135.240 ;
        RECT 37.555 135.180 37.875 135.240 ;
        RECT 38.490 135.380 38.780 135.425 ;
        RECT 42.155 135.380 42.475 135.440 ;
        RECT 38.490 135.240 42.475 135.380 ;
        RECT 38.490 135.195 38.780 135.240 ;
        RECT 42.155 135.180 42.475 135.240 ;
        RECT 32.955 134.900 34.565 135.040 ;
        RECT 32.955 134.840 33.275 134.900 ;
        RECT 37.095 134.840 37.415 135.100 ;
        RECT 38.015 135.040 38.335 135.100 ;
        RECT 43.625 135.085 43.765 135.920 ;
        RECT 45.375 135.860 45.695 135.920 ;
        RECT 54.575 135.860 54.895 135.920 ;
        RECT 55.495 135.860 55.815 136.120 ;
        RECT 62.855 136.060 63.175 136.120 ;
        RECT 66.535 136.060 66.855 136.120 ;
        RECT 68.850 136.060 69.140 136.105 ;
        RECT 62.855 135.920 69.140 136.060 ;
        RECT 62.855 135.860 63.175 135.920 ;
        RECT 66.535 135.860 66.855 135.920 ;
        RECT 68.850 135.875 69.140 135.920 ;
        RECT 72.070 136.060 72.360 136.105 ;
        RECT 74.355 136.060 74.675 136.120 ;
        RECT 83.555 136.060 83.875 136.120 ;
        RECT 87.710 136.060 88.000 136.105 ;
        RECT 72.070 135.920 74.675 136.060 ;
        RECT 72.070 135.875 72.360 135.920 ;
        RECT 74.355 135.860 74.675 135.920 ;
        RECT 77.665 135.920 88.000 136.060 ;
        RECT 53.195 135.720 53.515 135.780 ;
        RECT 61.935 135.720 62.255 135.780 ;
        RECT 77.665 135.720 77.805 135.920 ;
        RECT 83.555 135.860 83.875 135.920 ;
        RECT 87.710 135.875 88.000 135.920 ;
        RECT 100.115 135.860 100.435 136.120 ;
        RECT 101.495 136.060 101.815 136.120 ;
        RECT 101.970 136.060 102.260 136.105 ;
        RECT 101.495 135.920 102.260 136.060 ;
        RECT 101.495 135.860 101.815 135.920 ;
        RECT 101.970 135.875 102.260 135.920 ;
        RECT 106.570 136.060 106.860 136.105 ;
        RECT 107.015 136.060 107.335 136.120 ;
        RECT 106.570 135.920 107.335 136.060 ;
        RECT 106.570 135.875 106.860 135.920 ;
        RECT 107.015 135.860 107.335 135.920 ;
        RECT 80.795 135.720 81.115 135.780 ;
        RECT 84.015 135.720 84.335 135.780 ;
        RECT 85.870 135.720 86.160 135.765 ;
        RECT 52.825 135.580 53.515 135.720 ;
        RECT 52.825 135.425 52.965 135.580 ;
        RECT 53.195 135.520 53.515 135.580 ;
        RECT 53.745 135.580 62.255 135.720 ;
        RECT 52.750 135.195 53.040 135.425 ;
        RECT 43.550 135.040 43.840 135.085 ;
        RECT 38.015 134.900 43.840 135.040 ;
        RECT 38.015 134.840 38.335 134.900 ;
        RECT 43.550 134.855 43.840 134.900 ;
        RECT 43.995 134.840 44.315 135.100 ;
        RECT 44.470 135.040 44.760 135.085 ;
        RECT 44.915 135.040 45.235 135.100 ;
        RECT 44.470 134.900 45.235 135.040 ;
        RECT 44.470 134.855 44.760 134.900 ;
        RECT 44.915 134.840 45.235 134.900 ;
        RECT 45.390 134.855 45.680 135.085 ;
        RECT 46.295 135.040 46.615 135.100 ;
        RECT 51.815 135.040 52.135 135.100 ;
        RECT 53.745 135.085 53.885 135.580 ;
        RECT 61.935 135.520 62.255 135.580 ;
        RECT 72.145 135.580 77.805 135.720 ;
        RECT 78.125 135.580 82.865 135.720 ;
        RECT 56.890 135.380 57.180 135.425 ;
        RECT 57.335 135.380 57.655 135.440 ;
        RECT 56.890 135.240 57.655 135.380 ;
        RECT 56.890 135.195 57.180 135.240 ;
        RECT 57.335 135.180 57.655 135.240 ;
        RECT 59.175 135.180 59.495 135.440 ;
        RECT 64.235 135.380 64.555 135.440 ;
        RECT 63.405 135.240 64.555 135.380 ;
        RECT 53.210 135.040 53.500 135.085 ;
        RECT 46.295 134.900 53.500 135.040 ;
        RECT 30.210 134.700 30.500 134.745 ;
        RECT 32.510 134.700 32.800 134.745 ;
        RECT 38.950 134.700 39.240 134.745 ;
        RECT 30.210 134.560 39.240 134.700 ;
        RECT 30.210 134.515 30.500 134.560 ;
        RECT 32.510 134.515 32.800 134.560 ;
        RECT 38.950 134.515 39.240 134.560 ;
        RECT 42.615 134.700 42.935 134.760 ;
        RECT 45.465 134.700 45.605 134.855 ;
        RECT 46.295 134.840 46.615 134.900 ;
        RECT 51.815 134.840 52.135 134.900 ;
        RECT 53.210 134.855 53.500 134.900 ;
        RECT 53.670 134.855 53.960 135.085 ;
        RECT 56.430 135.040 56.720 135.085 ;
        RECT 59.265 135.040 59.405 135.180 ;
        RECT 63.405 135.085 63.545 135.240 ;
        RECT 64.235 135.180 64.555 135.240 ;
        RECT 64.710 135.380 65.000 135.425 ;
        RECT 66.995 135.380 67.315 135.440 ;
        RECT 64.710 135.240 67.315 135.380 ;
        RECT 64.710 135.195 65.000 135.240 ;
        RECT 66.995 135.180 67.315 135.240 ;
        RECT 56.430 134.900 59.405 135.040 ;
        RECT 56.430 134.855 56.720 134.900 ;
        RECT 60.110 134.855 60.400 135.085 ;
        RECT 63.330 134.855 63.620 135.085 ;
        RECT 63.775 135.040 64.095 135.100 ;
        RECT 68.390 135.040 68.680 135.085 ;
        RECT 63.775 134.900 68.680 135.040 ;
        RECT 72.145 135.040 72.285 135.580 ;
        RECT 76.195 135.380 76.515 135.440 ;
        RECT 78.125 135.425 78.265 135.580 ;
        RECT 80.795 135.520 81.115 135.580 ;
        RECT 82.725 135.425 82.865 135.580 ;
        RECT 84.015 135.580 86.160 135.720 ;
        RECT 84.015 135.520 84.335 135.580 ;
        RECT 85.870 135.535 86.160 135.580 ;
        RECT 74.905 135.240 76.515 135.380 ;
        RECT 72.530 135.040 72.820 135.085 ;
        RECT 72.145 134.900 72.820 135.040 ;
        RECT 42.615 134.560 45.605 134.700 ;
        RECT 46.755 134.700 47.075 134.760 ;
        RECT 60.185 134.700 60.325 134.855 ;
        RECT 63.775 134.840 64.095 134.900 ;
        RECT 68.390 134.855 68.680 134.900 ;
        RECT 72.530 134.855 72.820 134.900 ;
        RECT 72.975 135.040 73.295 135.100 ;
        RECT 74.905 135.085 75.045 135.240 ;
        RECT 76.195 135.180 76.515 135.240 ;
        RECT 78.050 135.195 78.340 135.425 ;
        RECT 82.650 135.195 82.940 135.425 ;
        RECT 89.995 135.380 90.315 135.440 ;
        RECT 97.355 135.380 97.675 135.440 ;
        RECT 89.995 135.240 91.605 135.380 ;
        RECT 89.995 135.180 90.315 135.240 ;
        RECT 73.450 135.040 73.740 135.085 ;
        RECT 74.370 135.040 74.660 135.085 ;
        RECT 72.975 134.900 73.740 135.040 ;
        RECT 72.975 134.840 73.295 134.900 ;
        RECT 73.450 134.855 73.740 134.900 ;
        RECT 73.985 134.900 74.660 135.040 ;
        RECT 73.985 134.760 74.125 134.900 ;
        RECT 74.370 134.855 74.660 134.900 ;
        RECT 74.830 134.855 75.120 135.085 ;
        RECT 75.275 134.840 75.595 135.100 ;
        RECT 78.970 135.040 79.260 135.085 ;
        RECT 79.875 135.040 80.195 135.100 ;
        RECT 83.570 135.040 83.860 135.085 ;
        RECT 78.970 134.900 83.860 135.040 ;
        RECT 78.970 134.855 79.260 134.900 ;
        RECT 79.875 134.840 80.195 134.900 ;
        RECT 83.570 134.855 83.860 134.900 ;
        RECT 87.235 134.840 87.555 135.100 ;
        RECT 91.465 135.085 91.605 135.240 ;
        RECT 94.225 135.240 97.675 135.380 ;
        RECT 90.930 134.855 91.220 135.085 ;
        RECT 91.390 134.855 91.680 135.085 ;
        RECT 61.475 134.700 61.795 134.760 ;
        RECT 61.950 134.700 62.240 134.745 ;
        RECT 46.755 134.560 62.240 134.700 ;
        RECT 42.615 134.500 42.935 134.560 ;
        RECT 46.755 134.500 47.075 134.560 ;
        RECT 61.475 134.500 61.795 134.560 ;
        RECT 61.950 134.515 62.240 134.560 ;
        RECT 65.630 134.700 65.920 134.745 ;
        RECT 73.895 134.700 74.215 134.760 ;
        RECT 78.510 134.700 78.800 134.745 ;
        RECT 65.630 134.560 78.800 134.700 ;
        RECT 65.630 134.515 65.920 134.560 ;
        RECT 73.895 134.500 74.215 134.560 ;
        RECT 78.510 134.515 78.800 134.560 ;
        RECT 21.930 134.360 22.220 134.405 ;
        RECT 27.895 134.360 28.215 134.420 ;
        RECT 35.715 134.360 36.035 134.420 ;
        RECT 21.930 134.220 36.035 134.360 ;
        RECT 21.930 134.175 22.220 134.220 ;
        RECT 27.895 134.160 28.215 134.220 ;
        RECT 35.715 134.160 36.035 134.220 ;
        RECT 36.190 134.360 36.480 134.405 ;
        RECT 38.015 134.360 38.335 134.420 ;
        RECT 36.190 134.220 38.335 134.360 ;
        RECT 36.190 134.175 36.480 134.220 ;
        RECT 38.015 134.160 38.335 134.220 ;
        RECT 39.395 134.160 39.715 134.420 ;
        RECT 42.155 134.160 42.475 134.420 ;
        RECT 64.695 134.360 65.015 134.420 ;
        RECT 65.170 134.360 65.460 134.405 ;
        RECT 64.695 134.220 65.460 134.360 ;
        RECT 64.695 134.160 65.015 134.220 ;
        RECT 65.170 134.175 65.460 134.220 ;
        RECT 67.455 134.160 67.775 134.420 ;
        RECT 76.655 134.160 76.975 134.420 ;
        RECT 80.810 134.360 81.100 134.405 ;
        RECT 81.255 134.360 81.575 134.420 ;
        RECT 80.810 134.220 81.575 134.360 ;
        RECT 80.810 134.175 81.100 134.220 ;
        RECT 81.255 134.160 81.575 134.220 ;
        RECT 83.555 134.360 83.875 134.420 ;
        RECT 84.030 134.360 84.320 134.405 ;
        RECT 83.555 134.220 84.320 134.360 ;
        RECT 83.555 134.160 83.875 134.220 ;
        RECT 84.030 134.175 84.320 134.220 ;
        RECT 85.395 134.360 85.715 134.420 ;
        RECT 89.550 134.360 89.840 134.405 ;
        RECT 85.395 134.220 89.840 134.360 ;
        RECT 91.005 134.360 91.145 134.855 ;
        RECT 91.465 134.700 91.605 134.855 ;
        RECT 91.835 134.840 92.155 135.100 ;
        RECT 92.295 135.040 92.615 135.100 ;
        RECT 94.225 135.085 94.365 135.240 ;
        RECT 97.355 135.180 97.675 135.240 ;
        RECT 92.770 135.040 93.060 135.085 ;
        RECT 93.230 135.040 93.520 135.085 ;
        RECT 92.295 134.900 93.520 135.040 ;
        RECT 92.295 134.840 92.615 134.900 ;
        RECT 92.770 134.855 93.060 134.900 ;
        RECT 93.230 134.855 93.520 134.900 ;
        RECT 94.150 134.855 94.440 135.085 ;
        RECT 94.610 134.855 94.900 135.085 ;
        RECT 94.685 134.700 94.825 134.855 ;
        RECT 95.055 134.840 95.375 135.100 ;
        RECT 99.670 134.855 99.960 135.085 ;
        RECT 100.575 135.040 100.895 135.100 ;
        RECT 101.510 135.040 101.800 135.085 ;
        RECT 100.575 134.900 101.800 135.040 ;
        RECT 91.465 134.560 94.825 134.700 ;
        RECT 99.745 134.700 99.885 134.855 ;
        RECT 100.575 134.840 100.895 134.900 ;
        RECT 101.510 134.855 101.800 134.900 ;
        RECT 107.030 135.040 107.320 135.085 ;
        RECT 107.475 135.040 107.795 135.100 ;
        RECT 107.030 134.900 107.795 135.040 ;
        RECT 107.030 134.855 107.320 134.900 ;
        RECT 105.175 134.700 105.495 134.760 ;
        RECT 107.105 134.700 107.245 134.855 ;
        RECT 107.475 134.840 107.795 134.900 ;
        RECT 99.745 134.560 107.245 134.700 ;
        RECT 105.175 134.500 105.495 134.560 ;
        RECT 135.660 134.480 136.800 134.510 ;
        RECT 94.135 134.360 94.455 134.420 ;
        RECT 91.005 134.220 94.455 134.360 ;
        RECT 85.395 134.160 85.715 134.220 ;
        RECT 89.550 134.175 89.840 134.220 ;
        RECT 94.135 134.160 94.455 134.220 ;
        RECT 96.450 134.360 96.740 134.405 ;
        RECT 97.815 134.360 98.135 134.420 ;
        RECT 96.450 134.220 98.135 134.360 ;
        RECT 96.450 134.175 96.740 134.220 ;
        RECT 97.815 134.160 98.135 134.220 ;
        RECT 18.165 133.540 112.465 134.020 ;
        RECT 135.590 133.400 136.850 134.480 ;
        RECT 35.715 133.340 36.035 133.400 ;
        RECT 38.475 133.340 38.795 133.400 ;
        RECT 35.715 133.200 38.795 133.340 ;
        RECT 35.715 133.140 36.035 133.200 ;
        RECT 38.475 133.140 38.795 133.200 ;
        RECT 39.395 133.340 39.715 133.400 ;
        RECT 60.555 133.385 60.875 133.400 ;
        RECT 60.340 133.340 60.875 133.385 ;
        RECT 64.695 133.340 65.015 133.400 ;
        RECT 39.395 133.200 65.015 133.340 ;
        RECT 39.395 133.140 39.715 133.200 ;
        RECT 60.340 133.155 60.875 133.200 ;
        RECT 60.555 133.140 60.875 133.155 ;
        RECT 64.695 133.140 65.015 133.200 ;
        RECT 72.975 133.340 73.295 133.400 ;
        RECT 82.635 133.340 82.955 133.400 ;
        RECT 72.975 133.200 83.785 133.340 ;
        RECT 72.975 133.140 73.295 133.200 ;
        RECT 82.635 133.140 82.955 133.200 ;
        RECT 21.010 133.000 21.300 133.045 ;
        RECT 27.550 133.000 27.840 133.045 ;
        RECT 30.790 133.000 31.440 133.045 ;
        RECT 21.010 132.860 31.440 133.000 ;
        RECT 21.010 132.815 21.300 132.860 ;
        RECT 27.550 132.815 28.140 132.860 ;
        RECT 30.790 132.815 31.440 132.860 ;
        RECT 32.955 133.000 33.275 133.060 ;
        RECT 43.995 133.000 44.315 133.060 ;
        RECT 51.010 133.000 51.300 133.045 ;
        RECT 51.815 133.000 52.135 133.060 ;
        RECT 54.250 133.000 54.900 133.045 ;
        RECT 32.955 132.860 39.165 133.000 ;
        RECT 21.455 132.460 21.775 132.720 ;
        RECT 27.850 132.500 28.140 132.815 ;
        RECT 32.955 132.800 33.275 132.860 ;
        RECT 28.930 132.660 29.220 132.705 ;
        RECT 32.510 132.660 32.800 132.705 ;
        RECT 34.345 132.660 34.635 132.705 ;
        RECT 28.930 132.520 34.635 132.660 ;
        RECT 28.930 132.475 29.220 132.520 ;
        RECT 32.510 132.475 32.800 132.520 ;
        RECT 34.345 132.475 34.635 132.520 ;
        RECT 36.190 132.660 36.480 132.705 ;
        RECT 36.635 132.660 36.955 132.720 ;
        RECT 36.190 132.520 36.955 132.660 ;
        RECT 36.190 132.475 36.480 132.520 ;
        RECT 36.635 132.460 36.955 132.520 ;
        RECT 38.015 132.460 38.335 132.720 ;
        RECT 38.475 132.460 38.795 132.720 ;
        RECT 39.025 132.705 39.165 132.860 ;
        RECT 39.945 132.860 47.445 133.000 ;
        RECT 39.945 132.705 40.085 132.860 ;
        RECT 43.995 132.800 44.315 132.860 ;
        RECT 38.950 132.475 39.240 132.705 ;
        RECT 39.870 132.475 40.160 132.705 ;
        RECT 41.235 132.660 41.555 132.720 ;
        RECT 45.390 132.660 45.680 132.705 ;
        RECT 41.235 132.520 45.680 132.660 ;
        RECT 41.235 132.460 41.555 132.520 ;
        RECT 45.390 132.475 45.680 132.520 ;
        RECT 45.835 132.460 46.155 132.720 ;
        RECT 47.305 132.705 47.445 132.860 ;
        RECT 51.010 132.860 54.900 133.000 ;
        RECT 51.010 132.815 51.600 132.860 ;
        RECT 46.310 132.475 46.600 132.705 ;
        RECT 47.230 132.475 47.520 132.705 ;
        RECT 51.310 132.500 51.600 132.815 ;
        RECT 51.815 132.800 52.135 132.860 ;
        RECT 54.250 132.815 54.900 132.860 ;
        RECT 55.495 133.000 55.815 133.060 ;
        RECT 56.890 133.000 57.180 133.045 ;
        RECT 55.495 132.860 57.180 133.000 ;
        RECT 55.495 132.800 55.815 132.860 ;
        RECT 56.890 132.815 57.180 132.860 ;
        RECT 57.335 133.000 57.655 133.060 ;
        RECT 83.645 133.045 83.785 133.200 ;
        RECT 62.345 133.000 62.635 133.045 ;
        RECT 65.605 133.000 65.895 133.045 ;
        RECT 57.335 132.860 65.895 133.000 ;
        RECT 57.335 132.800 57.655 132.860 ;
        RECT 62.345 132.815 62.635 132.860 ;
        RECT 65.605 132.815 65.895 132.860 ;
        RECT 66.525 133.000 66.815 133.045 ;
        RECT 68.385 133.000 68.675 133.045 ;
        RECT 66.525 132.860 68.675 133.000 ;
        RECT 66.525 132.815 66.815 132.860 ;
        RECT 68.385 132.815 68.675 132.860 ;
        RECT 76.145 133.000 76.435 133.045 ;
        RECT 79.405 133.000 79.695 133.045 ;
        RECT 76.145 132.860 79.695 133.000 ;
        RECT 76.145 132.815 76.435 132.860 ;
        RECT 79.405 132.815 79.695 132.860 ;
        RECT 80.325 133.000 80.615 133.045 ;
        RECT 82.185 133.000 82.475 133.045 ;
        RECT 80.325 132.860 82.475 133.000 ;
        RECT 80.325 132.815 80.615 132.860 ;
        RECT 82.185 132.815 82.475 132.860 ;
        RECT 83.570 132.815 83.860 133.045 ;
        RECT 94.595 133.000 94.915 133.060 ;
        RECT 96.450 133.000 96.740 133.045 ;
        RECT 94.595 132.860 96.740 133.000 ;
        RECT 52.390 132.660 52.680 132.705 ;
        RECT 55.970 132.660 56.260 132.705 ;
        RECT 57.805 132.660 58.095 132.705 ;
        RECT 52.390 132.520 58.095 132.660 ;
        RECT 52.390 132.475 52.680 132.520 ;
        RECT 55.970 132.475 56.260 132.520 ;
        RECT 57.805 132.475 58.095 132.520 ;
        RECT 64.205 132.660 64.495 132.705 ;
        RECT 66.525 132.660 66.740 132.815 ;
        RECT 64.205 132.520 66.740 132.660 ;
        RECT 64.205 132.475 64.495 132.520 ;
        RECT 22.850 132.320 23.140 132.365 ;
        RECT 22.850 132.180 34.565 132.320 ;
        RECT 22.850 132.135 23.140 132.180 ;
        RECT 28.930 131.980 29.220 132.025 ;
        RECT 32.050 131.980 32.340 132.025 ;
        RECT 33.940 131.980 34.230 132.025 ;
        RECT 28.930 131.840 34.230 131.980 ;
        RECT 34.425 131.980 34.565 132.180 ;
        RECT 34.795 132.120 35.115 132.380 ;
        RECT 37.555 132.320 37.875 132.380 ;
        RECT 35.345 132.180 37.875 132.320 ;
        RECT 35.345 131.980 35.485 132.180 ;
        RECT 37.555 132.120 37.875 132.180 ;
        RECT 40.790 132.320 41.080 132.365 ;
        RECT 46.385 132.320 46.525 132.475 ;
        RECT 67.455 132.460 67.775 132.720 ;
        RECT 72.055 132.460 72.375 132.720 ;
        RECT 72.530 132.660 72.820 132.705 ;
        RECT 76.285 132.660 76.425 132.815 ;
        RECT 72.530 132.520 76.425 132.660 ;
        RECT 78.005 132.660 78.295 132.705 ;
        RECT 80.325 132.660 80.540 132.815 ;
        RECT 94.595 132.800 94.915 132.860 ;
        RECT 96.450 132.815 96.740 132.860 ;
        RECT 96.910 133.000 97.200 133.045 ;
        RECT 97.355 133.000 97.675 133.060 ;
        RECT 96.910 132.860 97.675 133.000 ;
        RECT 96.910 132.815 97.200 132.860 ;
        RECT 97.355 132.800 97.675 132.860 ;
        RECT 99.195 133.000 99.515 133.060 ;
        RECT 101.970 133.000 102.260 133.045 ;
        RECT 99.195 132.860 102.260 133.000 ;
        RECT 99.195 132.800 99.515 132.860 ;
        RECT 101.970 132.815 102.260 132.860 ;
        RECT 104.250 133.000 104.900 133.045 ;
        RECT 105.635 133.000 105.955 133.060 ;
        RECT 107.850 133.000 108.140 133.045 ;
        RECT 104.250 132.860 108.140 133.000 ;
        RECT 104.250 132.815 104.900 132.860 ;
        RECT 105.635 132.800 105.955 132.860 ;
        RECT 107.550 132.815 108.140 132.860 ;
        RECT 78.005 132.520 80.540 132.660 ;
        RECT 72.530 132.475 72.820 132.520 ;
        RECT 78.005 132.475 78.295 132.520 ;
        RECT 81.255 132.460 81.575 132.720 ;
        RECT 89.075 132.660 89.395 132.720 ;
        RECT 92.295 132.660 92.615 132.720 ;
        RECT 99.655 132.660 99.975 132.720 ;
        RECT 100.575 132.660 100.895 132.720 ;
        RECT 89.075 132.520 100.895 132.660 ;
        RECT 89.075 132.460 89.395 132.520 ;
        RECT 92.295 132.460 92.615 132.520 ;
        RECT 99.655 132.460 99.975 132.520 ;
        RECT 100.575 132.460 100.895 132.520 ;
        RECT 101.055 132.660 101.345 132.705 ;
        RECT 102.890 132.660 103.180 132.705 ;
        RECT 106.470 132.660 106.760 132.705 ;
        RECT 101.055 132.520 106.760 132.660 ;
        RECT 101.055 132.475 101.345 132.520 ;
        RECT 102.890 132.475 103.180 132.520 ;
        RECT 106.470 132.475 106.760 132.520 ;
        RECT 107.550 132.500 107.840 132.815 ;
        RECT 110.695 132.800 111.015 133.060 ;
        RECT 49.530 132.320 49.820 132.365 ;
        RECT 40.790 132.180 49.820 132.320 ;
        RECT 40.790 132.135 41.080 132.180 ;
        RECT 49.530 132.135 49.820 132.180 ;
        RECT 56.415 132.320 56.735 132.380 ;
        RECT 58.255 132.320 58.575 132.380 ;
        RECT 56.415 132.180 58.575 132.320 ;
        RECT 56.415 132.120 56.735 132.180 ;
        RECT 58.255 132.120 58.575 132.180 ;
        RECT 69.310 132.320 69.600 132.365 ;
        RECT 73.895 132.320 74.215 132.380 ;
        RECT 69.310 132.180 72.745 132.320 ;
        RECT 69.310 132.135 69.600 132.180 ;
        RECT 72.605 132.040 72.745 132.180 ;
        RECT 73.895 132.120 74.355 132.320 ;
        RECT 83.095 132.120 83.415 132.380 ;
        RECT 94.135 132.320 94.455 132.380 ;
        RECT 95.530 132.320 95.820 132.365 ;
        RECT 94.135 132.180 95.820 132.320 ;
        RECT 94.135 132.120 94.455 132.180 ;
        RECT 95.530 132.135 95.820 132.180 ;
        RECT 34.425 131.840 35.485 131.980 ;
        RECT 37.095 131.980 37.415 132.040 ;
        RECT 44.010 131.980 44.300 132.025 ;
        RECT 37.095 131.840 44.300 131.980 ;
        RECT 28.930 131.795 29.220 131.840 ;
        RECT 32.050 131.795 32.340 131.840 ;
        RECT 33.940 131.795 34.230 131.840 ;
        RECT 37.095 131.780 37.415 131.840 ;
        RECT 44.010 131.795 44.300 131.840 ;
        RECT 52.390 131.980 52.680 132.025 ;
        RECT 55.510 131.980 55.800 132.025 ;
        RECT 57.400 131.980 57.690 132.025 ;
        RECT 52.390 131.840 57.690 131.980 ;
        RECT 52.390 131.795 52.680 131.840 ;
        RECT 55.510 131.795 55.800 131.840 ;
        RECT 57.400 131.795 57.690 131.840 ;
        RECT 64.205 131.980 64.495 132.025 ;
        RECT 66.985 131.980 67.275 132.025 ;
        RECT 68.845 131.980 69.135 132.025 ;
        RECT 64.205 131.840 69.135 131.980 ;
        RECT 64.205 131.795 64.495 131.840 ;
        RECT 66.985 131.795 67.275 131.840 ;
        RECT 68.845 131.795 69.135 131.840 ;
        RECT 72.515 131.780 72.835 132.040 ;
        RECT 25.595 131.440 25.915 131.700 ;
        RECT 26.055 131.440 26.375 131.700 ;
        RECT 33.415 131.685 33.735 131.700 ;
        RECT 33.415 131.455 33.785 131.685 ;
        RECT 33.415 131.440 33.735 131.455 ;
        RECT 35.715 131.440 36.035 131.700 ;
        RECT 36.175 131.640 36.495 131.700 ;
        RECT 36.650 131.640 36.940 131.685 ;
        RECT 36.175 131.500 36.940 131.640 ;
        RECT 36.175 131.440 36.495 131.500 ;
        RECT 36.650 131.455 36.940 131.500 ;
        RECT 43.535 131.440 43.855 131.700 ;
        RECT 61.015 131.640 61.335 131.700 ;
        RECT 72.975 131.640 73.295 131.700 ;
        RECT 74.215 131.685 74.355 132.120 ;
        RECT 78.005 131.980 78.295 132.025 ;
        RECT 80.785 131.980 81.075 132.025 ;
        RECT 82.645 131.980 82.935 132.025 ;
        RECT 78.005 131.840 82.935 131.980 ;
        RECT 78.005 131.795 78.295 131.840 ;
        RECT 80.785 131.795 81.075 131.840 ;
        RECT 82.645 131.795 82.935 131.840 ;
        RECT 101.460 131.980 101.750 132.025 ;
        RECT 103.350 131.980 103.640 132.025 ;
        RECT 106.470 131.980 106.760 132.025 ;
        RECT 101.460 131.840 106.760 131.980 ;
        RECT 101.460 131.795 101.750 131.840 ;
        RECT 103.350 131.795 103.640 131.840 ;
        RECT 106.470 131.795 106.760 131.840 ;
        RECT 61.015 131.500 73.295 131.640 ;
        RECT 61.015 131.440 61.335 131.500 ;
        RECT 72.975 131.440 73.295 131.500 ;
        RECT 74.140 131.455 74.430 131.685 ;
        RECT 98.750 131.640 99.040 131.685 ;
        RECT 99.655 131.640 99.975 131.700 ;
        RECT 98.750 131.500 99.975 131.640 ;
        RECT 98.750 131.455 99.040 131.500 ;
        RECT 99.655 131.440 99.975 131.500 ;
        RECT 17.605 130.820 112.465 131.300 ;
        RECT 25.595 130.620 25.915 130.680 ;
        RECT 30.655 130.620 30.975 130.680 ;
        RECT 33.415 130.620 33.735 130.680 ;
        RECT 33.890 130.620 34.180 130.665 ;
        RECT 25.595 130.480 30.425 130.620 ;
        RECT 25.595 130.420 25.915 130.480 ;
        RECT 23.870 130.280 24.160 130.325 ;
        RECT 26.990 130.280 27.280 130.325 ;
        RECT 28.880 130.280 29.170 130.325 ;
        RECT 23.870 130.140 29.170 130.280 ;
        RECT 23.870 130.095 24.160 130.140 ;
        RECT 26.990 130.095 27.280 130.140 ;
        RECT 28.880 130.095 29.170 130.140 ;
        RECT 19.615 129.060 19.935 129.320 ;
        RECT 20.995 129.260 21.315 129.320 ;
        RECT 22.790 129.305 23.080 129.620 ;
        RECT 23.870 129.600 24.160 129.645 ;
        RECT 27.450 129.600 27.740 129.645 ;
        RECT 29.285 129.600 29.575 129.645 ;
        RECT 23.870 129.460 29.575 129.600 ;
        RECT 23.870 129.415 24.160 129.460 ;
        RECT 27.450 129.415 27.740 129.460 ;
        RECT 29.285 129.415 29.575 129.460 ;
        RECT 29.750 129.415 30.040 129.645 ;
        RECT 30.285 129.600 30.425 130.480 ;
        RECT 30.655 130.480 32.725 130.620 ;
        RECT 30.655 130.420 30.975 130.480 ;
        RECT 32.035 130.280 32.355 130.340 ;
        RECT 31.205 130.140 32.355 130.280 ;
        RECT 32.585 130.280 32.725 130.480 ;
        RECT 33.415 130.480 34.180 130.620 ;
        RECT 33.415 130.420 33.735 130.480 ;
        RECT 33.890 130.435 34.180 130.480 ;
        RECT 41.695 130.620 42.015 130.680 ;
        RECT 45.835 130.620 46.155 130.680 ;
        RECT 41.695 130.480 46.155 130.620 ;
        RECT 41.695 130.420 42.015 130.480 ;
        RECT 45.835 130.420 46.155 130.480 ;
        RECT 52.735 130.620 53.055 130.680 ;
        RECT 105.635 130.620 105.955 130.680 ;
        RECT 106.110 130.620 106.400 130.665 ;
        RECT 52.735 130.480 62.165 130.620 ;
        RECT 52.735 130.420 53.055 130.480 ;
        RECT 48.595 130.280 48.915 130.340 ;
        RECT 32.585 130.140 48.915 130.280 ;
        RECT 31.205 129.985 31.345 130.140 ;
        RECT 32.035 130.080 32.355 130.140 ;
        RECT 48.595 130.080 48.915 130.140 ;
        RECT 31.130 129.755 31.420 129.985 ;
        RECT 33.415 129.940 33.735 130.000 ;
        RECT 35.255 129.940 35.575 130.000 ;
        RECT 33.415 129.800 35.575 129.940 ;
        RECT 33.415 129.740 33.735 129.800 ;
        RECT 35.255 129.740 35.575 129.800 ;
        RECT 36.635 129.940 36.955 130.000 ;
        RECT 52.275 129.940 52.595 130.000 ;
        RECT 62.025 129.985 62.165 130.480 ;
        RECT 105.635 130.480 106.400 130.620 ;
        RECT 105.635 130.420 105.955 130.480 ;
        RECT 106.110 130.435 106.400 130.480 ;
        RECT 69.870 130.280 70.160 130.325 ;
        RECT 72.990 130.280 73.280 130.325 ;
        RECT 74.880 130.280 75.170 130.325 ;
        RECT 69.870 130.140 75.170 130.280 ;
        RECT 69.870 130.095 70.160 130.140 ;
        RECT 72.990 130.095 73.280 130.140 ;
        RECT 74.880 130.095 75.170 130.140 ;
        RECT 80.765 130.280 81.055 130.325 ;
        RECT 83.545 130.280 83.835 130.325 ;
        RECT 85.405 130.280 85.695 130.325 ;
        RECT 80.765 130.140 85.695 130.280 ;
        RECT 80.765 130.095 81.055 130.140 ;
        RECT 83.545 130.095 83.835 130.140 ;
        RECT 85.405 130.095 85.695 130.140 ;
        RECT 97.930 130.280 98.220 130.325 ;
        RECT 101.050 130.280 101.340 130.325 ;
        RECT 102.940 130.280 103.230 130.325 ;
        RECT 97.930 130.140 103.230 130.280 ;
        RECT 97.930 130.095 98.220 130.140 ;
        RECT 101.050 130.095 101.340 130.140 ;
        RECT 102.940 130.095 103.230 130.140 ;
        RECT 61.950 129.940 62.240 129.985 ;
        RECT 70.675 129.940 70.995 130.000 ;
        RECT 36.635 129.800 59.405 129.940 ;
        RECT 36.635 129.740 36.955 129.800 ;
        RECT 52.275 129.740 52.595 129.800 ;
        RECT 59.265 129.660 59.405 129.800 ;
        RECT 61.950 129.800 70.995 129.940 ;
        RECT 61.950 129.755 62.240 129.800 ;
        RECT 70.675 129.740 70.995 129.800 ;
        RECT 71.595 129.940 71.915 130.000 ;
        RECT 74.370 129.940 74.660 129.985 ;
        RECT 83.095 129.940 83.415 130.000 ;
        RECT 71.595 129.800 74.660 129.940 ;
        RECT 71.595 129.740 71.915 129.800 ;
        RECT 74.370 129.755 74.660 129.800 ;
        RECT 75.825 129.800 83.785 129.940 ;
        RECT 75.825 129.660 75.965 129.800 ;
        RECT 83.095 129.740 83.415 129.800 ;
        RECT 32.050 129.600 32.340 129.645 ;
        RECT 30.285 129.460 32.340 129.600 ;
        RECT 32.050 129.415 32.340 129.460 ;
        RECT 22.490 129.260 23.080 129.305 ;
        RECT 25.730 129.260 26.380 129.305 ;
        RECT 20.995 129.120 26.380 129.260 ;
        RECT 20.995 129.060 21.315 129.120 ;
        RECT 22.490 129.075 22.780 129.120 ;
        RECT 25.730 129.075 26.380 129.120 ;
        RECT 28.370 129.075 28.660 129.305 ;
        RECT 29.825 129.260 29.965 129.415 ;
        RECT 55.955 129.400 56.275 129.660 ;
        RECT 59.175 129.400 59.495 129.660 ;
        RECT 32.955 129.260 33.275 129.320 ;
        RECT 34.795 129.260 35.115 129.320 ;
        RECT 35.730 129.260 36.020 129.305 ;
        RECT 29.825 129.120 36.020 129.260 ;
        RECT 28.445 128.920 28.585 129.075 ;
        RECT 32.955 129.060 33.275 129.120 ;
        RECT 34.795 129.060 35.115 129.120 ;
        RECT 35.730 129.075 36.020 129.120 ;
        RECT 44.470 129.260 44.760 129.305 ;
        RECT 47.675 129.260 47.995 129.320 ;
        RECT 61.015 129.260 61.335 129.320 ;
        RECT 44.470 129.120 61.335 129.260 ;
        RECT 44.470 129.075 44.760 129.120 ;
        RECT 47.675 129.060 47.995 129.120 ;
        RECT 61.015 129.060 61.335 129.120 ;
        RECT 62.870 129.260 63.160 129.305 ;
        RECT 67.915 129.260 68.235 129.320 ;
        RECT 68.790 129.305 69.080 129.620 ;
        RECT 69.870 129.600 70.160 129.645 ;
        RECT 73.450 129.600 73.740 129.645 ;
        RECT 75.285 129.600 75.575 129.645 ;
        RECT 69.870 129.460 75.575 129.600 ;
        RECT 69.870 129.415 70.160 129.460 ;
        RECT 73.450 129.415 73.740 129.460 ;
        RECT 75.285 129.415 75.575 129.460 ;
        RECT 75.735 129.400 76.055 129.660 ;
        RECT 80.765 129.600 81.055 129.645 ;
        RECT 83.645 129.600 83.785 129.800 ;
        RECT 84.015 129.740 84.335 130.000 ;
        RECT 89.535 129.940 89.855 130.000 ;
        RECT 95.055 129.940 95.375 130.000 ;
        RECT 89.535 129.800 95.375 129.940 ;
        RECT 89.535 129.740 89.855 129.800 ;
        RECT 95.055 129.740 95.375 129.800 ;
        RECT 100.575 129.940 100.895 130.000 ;
        RECT 103.795 129.940 104.115 130.000 ;
        RECT 100.575 129.800 104.115 129.940 ;
        RECT 100.575 129.740 100.895 129.800 ;
        RECT 103.795 129.740 104.115 129.800 ;
        RECT 85.870 129.600 86.160 129.645 ;
        RECT 80.765 129.460 83.300 129.600 ;
        RECT 83.645 129.460 86.160 129.600 ;
        RECT 80.765 129.415 81.055 129.460 ;
        RECT 83.085 129.305 83.300 129.460 ;
        RECT 85.870 129.415 86.160 129.460 ;
        RECT 92.295 129.400 92.615 129.660 ;
        RECT 92.770 129.415 93.060 129.645 ;
        RECT 68.490 129.260 69.080 129.305 ;
        RECT 71.730 129.260 72.380 129.305 ;
        RECT 62.870 129.120 67.685 129.260 ;
        RECT 62.870 129.075 63.160 129.120 ;
        RECT 30.195 128.920 30.515 128.980 ;
        RECT 28.445 128.780 30.515 128.920 ;
        RECT 30.195 128.720 30.515 128.780 ;
        RECT 31.590 128.920 31.880 128.965 ;
        RECT 32.035 128.920 32.355 128.980 ;
        RECT 31.590 128.780 32.355 128.920 ;
        RECT 31.590 128.735 31.880 128.780 ;
        RECT 32.035 128.720 32.355 128.780 ;
        RECT 59.635 128.720 59.955 128.980 ;
        RECT 62.395 128.720 62.715 128.980 ;
        RECT 64.235 128.920 64.555 128.980 ;
        RECT 64.710 128.920 65.000 128.965 ;
        RECT 64.235 128.780 65.000 128.920 ;
        RECT 64.235 128.720 64.555 128.780 ;
        RECT 64.710 128.735 65.000 128.780 ;
        RECT 65.615 128.920 65.935 128.980 ;
        RECT 67.010 128.920 67.300 128.965 ;
        RECT 65.615 128.780 67.300 128.920 ;
        RECT 67.545 128.920 67.685 129.120 ;
        RECT 67.915 129.120 72.380 129.260 ;
        RECT 67.915 129.060 68.235 129.120 ;
        RECT 68.490 129.075 68.780 129.120 ;
        RECT 71.730 129.075 72.380 129.120 ;
        RECT 78.905 129.260 79.195 129.305 ;
        RECT 82.165 129.260 82.455 129.305 ;
        RECT 83.085 129.260 83.375 129.305 ;
        RECT 84.945 129.260 85.235 129.305 ;
        RECT 78.905 129.120 82.865 129.260 ;
        RECT 78.905 129.075 79.195 129.120 ;
        RECT 82.165 129.075 82.455 129.120 ;
        RECT 69.295 128.920 69.615 128.980 ;
        RECT 67.545 128.780 69.615 128.920 ;
        RECT 65.615 128.720 65.935 128.780 ;
        RECT 67.010 128.735 67.300 128.780 ;
        RECT 69.295 128.720 69.615 128.780 ;
        RECT 76.900 128.920 77.190 128.965 ;
        RECT 79.875 128.920 80.195 128.980 ;
        RECT 76.900 128.780 80.195 128.920 ;
        RECT 82.725 128.920 82.865 129.120 ;
        RECT 83.085 129.120 85.235 129.260 ;
        RECT 83.085 129.075 83.375 129.120 ;
        RECT 84.945 129.075 85.235 129.120 ;
        RECT 89.075 129.260 89.395 129.320 ;
        RECT 92.845 129.260 92.985 129.415 ;
        RECT 96.850 129.305 97.140 129.620 ;
        RECT 97.930 129.600 98.220 129.645 ;
        RECT 101.510 129.600 101.800 129.645 ;
        RECT 103.345 129.600 103.635 129.645 ;
        RECT 97.930 129.460 103.635 129.600 ;
        RECT 97.930 129.415 98.220 129.460 ;
        RECT 101.510 129.415 101.800 129.460 ;
        RECT 103.345 129.415 103.635 129.460 ;
        RECT 105.175 129.600 105.495 129.660 ;
        RECT 105.650 129.600 105.940 129.645 ;
        RECT 105.175 129.460 105.940 129.600 ;
        RECT 105.175 129.400 105.495 129.460 ;
        RECT 105.650 129.415 105.940 129.460 ;
        RECT 89.075 129.120 92.985 129.260 ;
        RECT 96.550 129.260 97.140 129.305 ;
        RECT 98.735 129.260 99.055 129.320 ;
        RECT 99.790 129.260 100.440 129.305 ;
        RECT 96.550 129.120 100.440 129.260 ;
        RECT 89.075 129.060 89.395 129.120 ;
        RECT 96.550 129.075 96.840 129.120 ;
        RECT 98.735 129.060 99.055 129.120 ;
        RECT 99.790 129.075 100.440 129.120 ;
        RECT 102.430 129.260 102.720 129.305 ;
        RECT 102.875 129.260 103.195 129.320 ;
        RECT 102.430 129.120 103.195 129.260 ;
        RECT 102.430 129.075 102.720 129.120 ;
        RECT 102.875 129.060 103.195 129.120 ;
        RECT 93.230 128.920 93.520 128.965 ;
        RECT 82.725 128.780 93.520 128.920 ;
        RECT 76.900 128.735 77.190 128.780 ;
        RECT 79.875 128.720 80.195 128.780 ;
        RECT 93.230 128.735 93.520 128.780 ;
        RECT 94.595 128.920 94.915 128.980 ;
        RECT 95.070 128.920 95.360 128.965 ;
        RECT 95.515 128.920 95.835 128.980 ;
        RECT 94.595 128.780 95.835 128.920 ;
        RECT 94.595 128.720 94.915 128.780 ;
        RECT 95.070 128.735 95.360 128.780 ;
        RECT 95.515 128.720 95.835 128.780 ;
        RECT 18.165 128.100 112.465 128.580 ;
        RECT 21.010 127.900 21.300 127.945 ;
        RECT 38.935 127.900 39.255 127.960 ;
        RECT 21.010 127.760 24.905 127.900 ;
        RECT 21.010 127.715 21.300 127.760 ;
        RECT 24.765 127.560 24.905 127.760 ;
        RECT 36.265 127.760 39.255 127.900 ;
        RECT 25.250 127.560 25.540 127.605 ;
        RECT 28.490 127.560 29.140 127.605 ;
        RECT 24.765 127.420 29.140 127.560 ;
        RECT 25.250 127.375 25.840 127.420 ;
        RECT 28.490 127.375 29.140 127.420 ;
        RECT 21.470 127.220 21.760 127.265 ;
        RECT 21.915 127.220 22.235 127.280 ;
        RECT 24.215 127.220 24.535 127.280 ;
        RECT 21.470 127.080 24.535 127.220 ;
        RECT 21.470 127.035 21.760 127.080 ;
        RECT 21.915 127.020 22.235 127.080 ;
        RECT 24.215 127.020 24.535 127.080 ;
        RECT 25.550 127.060 25.840 127.375 ;
        RECT 26.630 127.220 26.920 127.265 ;
        RECT 30.210 127.220 30.500 127.265 ;
        RECT 32.045 127.220 32.335 127.265 ;
        RECT 26.630 127.080 32.335 127.220 ;
        RECT 26.630 127.035 26.920 127.080 ;
        RECT 30.210 127.035 30.500 127.080 ;
        RECT 32.045 127.035 32.335 127.080 ;
        RECT 33.875 127.020 34.195 127.280 ;
        RECT 34.795 127.220 35.115 127.280 ;
        RECT 36.265 127.220 36.405 127.760 ;
        RECT 38.935 127.700 39.255 127.760 ;
        RECT 51.815 127.700 52.135 127.960 ;
        RECT 55.495 127.900 55.815 127.960 ;
        RECT 56.430 127.900 56.720 127.945 ;
        RECT 88.615 127.900 88.935 127.960 ;
        RECT 92.295 127.900 92.615 127.960 ;
        RECT 98.290 127.900 98.580 127.945 ;
        RECT 98.735 127.900 99.055 127.960 ;
        RECT 55.495 127.760 56.720 127.900 ;
        RECT 55.495 127.700 55.815 127.760 ;
        RECT 56.430 127.715 56.720 127.760 ;
        RECT 58.805 127.760 65.845 127.900 ;
        RECT 38.015 127.560 38.335 127.620 ;
        RECT 36.725 127.420 38.335 127.560 ;
        RECT 36.725 127.265 36.865 127.420 ;
        RECT 38.015 127.360 38.335 127.420 ;
        RECT 39.870 127.560 40.160 127.605 ;
        RECT 40.315 127.560 40.635 127.620 ;
        RECT 43.535 127.560 43.855 127.620 ;
        RECT 45.390 127.560 45.680 127.605 ;
        RECT 52.275 127.560 52.595 127.620 ;
        RECT 39.870 127.420 40.635 127.560 ;
        RECT 39.870 127.375 40.160 127.420 ;
        RECT 40.315 127.360 40.635 127.420 ;
        RECT 40.865 127.420 43.305 127.560 ;
        RECT 34.795 127.080 36.405 127.220 ;
        RECT 34.795 127.020 35.115 127.080 ;
        RECT 22.375 126.680 22.695 126.940 ;
        RECT 31.115 126.680 31.435 126.940 ;
        RECT 32.510 126.880 32.800 126.925 ;
        RECT 32.955 126.880 33.275 126.940 ;
        RECT 32.510 126.740 33.275 126.880 ;
        RECT 36.265 126.880 36.405 127.080 ;
        RECT 36.650 127.035 36.940 127.265 ;
        RECT 37.110 127.035 37.400 127.265 ;
        RECT 37.185 126.880 37.325 127.035 ;
        RECT 37.555 127.020 37.875 127.280 ;
        RECT 38.490 127.220 38.780 127.265 ;
        RECT 39.395 127.220 39.715 127.280 ;
        RECT 40.865 127.220 41.005 127.420 ;
        RECT 38.490 127.080 41.005 127.220 ;
        RECT 38.490 127.035 38.780 127.080 ;
        RECT 39.395 127.020 39.715 127.080 ;
        RECT 41.235 127.020 41.555 127.280 ;
        RECT 41.695 127.020 42.015 127.280 ;
        RECT 43.165 127.265 43.305 127.420 ;
        RECT 43.535 127.420 45.680 127.560 ;
        RECT 43.535 127.360 43.855 127.420 ;
        RECT 45.390 127.375 45.680 127.420 ;
        RECT 51.445 127.420 52.595 127.560 ;
        RECT 42.170 127.035 42.460 127.265 ;
        RECT 43.090 127.220 43.380 127.265 ;
        RECT 43.995 127.220 44.315 127.280 ;
        RECT 43.090 127.080 44.315 127.220 ;
        RECT 43.090 127.035 43.380 127.080 ;
        RECT 36.265 126.740 37.325 126.880 ;
        RECT 38.015 126.880 38.335 126.940 ;
        RECT 42.245 126.880 42.385 127.035 ;
        RECT 43.995 127.020 44.315 127.080 ;
        RECT 38.015 126.740 42.385 126.880 ;
        RECT 32.510 126.695 32.800 126.740 ;
        RECT 32.955 126.680 33.275 126.740 ;
        RECT 38.015 126.680 38.335 126.740 ;
        RECT 44.470 126.695 44.760 126.925 ;
        RECT 26.630 126.540 26.920 126.585 ;
        RECT 29.750 126.540 30.040 126.585 ;
        RECT 31.640 126.540 31.930 126.585 ;
        RECT 26.630 126.400 31.930 126.540 ;
        RECT 26.630 126.355 26.920 126.400 ;
        RECT 29.750 126.355 30.040 126.400 ;
        RECT 31.640 126.355 31.930 126.400 ;
        RECT 34.810 126.540 35.100 126.585 ;
        RECT 39.395 126.540 39.715 126.600 ;
        RECT 34.810 126.400 39.715 126.540 ;
        RECT 44.545 126.540 44.685 126.695 ;
        RECT 44.915 126.680 45.235 126.940 ;
        RECT 45.465 126.880 45.605 127.375 ;
        RECT 47.215 127.220 47.535 127.280 ;
        RECT 51.445 127.265 51.585 127.420 ;
        RECT 52.275 127.360 52.595 127.420 ;
        RECT 55.955 127.560 56.275 127.620 ;
        RECT 58.805 127.560 58.945 127.760 ;
        RECT 55.955 127.420 58.945 127.560 ;
        RECT 59.125 127.560 59.415 127.605 ;
        RECT 59.635 127.560 59.955 127.620 ;
        RECT 62.385 127.560 62.675 127.605 ;
        RECT 59.125 127.420 62.675 127.560 ;
        RECT 55.955 127.360 56.275 127.420 ;
        RECT 59.125 127.375 59.415 127.420 ;
        RECT 59.635 127.360 59.955 127.420 ;
        RECT 62.385 127.375 62.675 127.420 ;
        RECT 63.305 127.560 63.595 127.605 ;
        RECT 65.165 127.560 65.455 127.605 ;
        RECT 63.305 127.420 65.455 127.560 ;
        RECT 63.305 127.375 63.595 127.420 ;
        RECT 65.165 127.375 65.455 127.420 ;
        RECT 48.150 127.220 48.440 127.265 ;
        RECT 47.215 127.080 48.440 127.220 ;
        RECT 47.215 127.020 47.535 127.080 ;
        RECT 48.150 127.035 48.440 127.080 ;
        RECT 51.370 127.035 51.660 127.265 ;
        RECT 54.130 127.220 54.420 127.265 ;
        RECT 51.905 127.080 54.420 127.220 ;
        RECT 51.905 126.880 52.045 127.080 ;
        RECT 54.130 127.035 54.420 127.080 ;
        RECT 54.590 127.035 54.880 127.265 ;
        RECT 60.985 127.220 61.275 127.265 ;
        RECT 63.305 127.220 63.520 127.375 ;
        RECT 60.985 127.080 63.520 127.220 ;
        RECT 60.985 127.035 61.275 127.080 ;
        RECT 45.465 126.740 52.045 126.880 ;
        RECT 52.735 126.880 53.055 126.940 ;
        RECT 53.210 126.880 53.500 126.925 ;
        RECT 52.735 126.740 53.500 126.880 ;
        RECT 54.665 126.880 54.805 127.035 ;
        RECT 64.235 127.020 64.555 127.280 ;
        RECT 65.705 127.220 65.845 127.760 ;
        RECT 88.615 127.760 94.825 127.900 ;
        RECT 88.615 127.700 88.935 127.760 ;
        RECT 92.295 127.700 92.615 127.760 ;
        RECT 73.895 127.560 74.215 127.620 ;
        RECT 68.925 127.420 74.215 127.560 ;
        RECT 66.090 127.220 66.380 127.265 ;
        RECT 65.705 127.080 66.380 127.220 ;
        RECT 66.090 127.035 66.380 127.080 ;
        RECT 67.915 127.220 68.235 127.280 ;
        RECT 68.925 127.265 69.065 127.420 ;
        RECT 73.895 127.360 74.215 127.420 ;
        RECT 82.635 127.360 82.955 127.620 ;
        RECT 85.805 127.560 86.095 127.605 ;
        RECT 87.235 127.560 87.555 127.620 ;
        RECT 89.065 127.560 89.355 127.605 ;
        RECT 85.805 127.420 89.355 127.560 ;
        RECT 85.805 127.375 86.095 127.420 ;
        RECT 87.235 127.360 87.555 127.420 ;
        RECT 89.065 127.375 89.355 127.420 ;
        RECT 89.985 127.560 90.275 127.605 ;
        RECT 91.845 127.560 92.135 127.605 ;
        RECT 89.985 127.420 92.135 127.560 ;
        RECT 89.985 127.375 90.275 127.420 ;
        RECT 91.845 127.375 92.135 127.420 ;
        RECT 68.390 127.220 68.680 127.265 ;
        RECT 67.915 127.080 68.680 127.220 ;
        RECT 67.915 127.020 68.235 127.080 ;
        RECT 68.390 127.035 68.680 127.080 ;
        RECT 68.850 127.035 69.140 127.265 ;
        RECT 71.135 127.020 71.455 127.280 ;
        RECT 72.515 127.220 72.835 127.280 ;
        RECT 74.370 127.220 74.660 127.265 ;
        RECT 75.735 127.220 76.055 127.280 ;
        RECT 72.515 127.080 76.055 127.220 ;
        RECT 72.515 127.020 72.835 127.080 ;
        RECT 74.370 127.035 74.660 127.080 ;
        RECT 75.735 127.020 76.055 127.080 ;
        RECT 83.555 127.265 83.875 127.280 ;
        RECT 83.555 127.035 84.090 127.265 ;
        RECT 87.665 127.220 87.955 127.265 ;
        RECT 89.985 127.220 90.200 127.375 ;
        RECT 87.665 127.080 90.200 127.220 ;
        RECT 91.375 127.220 91.695 127.280 ;
        RECT 92.770 127.220 93.060 127.265 ;
        RECT 94.135 127.220 94.455 127.280 ;
        RECT 94.685 127.265 94.825 127.760 ;
        RECT 98.290 127.760 99.055 127.900 ;
        RECT 98.290 127.715 98.580 127.760 ;
        RECT 98.735 127.700 99.055 127.760 ;
        RECT 102.875 127.700 103.195 127.960 ;
        RECT 105.175 127.560 105.495 127.620 ;
        RECT 103.425 127.420 105.495 127.560 ;
        RECT 91.375 127.080 94.455 127.220 ;
        RECT 87.665 127.035 87.955 127.080 ;
        RECT 83.555 127.020 83.875 127.035 ;
        RECT 91.375 127.020 91.695 127.080 ;
        RECT 92.770 127.035 93.060 127.080 ;
        RECT 94.135 127.020 94.455 127.080 ;
        RECT 94.610 127.035 94.900 127.265 ;
        RECT 95.055 127.020 95.375 127.280 ;
        RECT 95.515 127.020 95.835 127.280 ;
        RECT 96.450 127.035 96.740 127.265 ;
        RECT 98.750 127.035 99.040 127.265 ;
        RECT 57.120 126.880 57.410 126.925 ;
        RECT 62.395 126.880 62.715 126.940 ;
        RECT 54.665 126.740 62.715 126.880 ;
        RECT 52.735 126.680 53.055 126.740 ;
        RECT 53.210 126.695 53.500 126.740 ;
        RECT 57.120 126.695 57.410 126.740 ;
        RECT 62.395 126.680 62.715 126.740 ;
        RECT 69.770 126.695 70.060 126.925 ;
        RECT 70.690 126.880 70.980 126.925 ;
        RECT 79.415 126.880 79.735 126.940 ;
        RECT 70.690 126.740 79.735 126.880 ;
        RECT 70.690 126.695 70.980 126.740 ;
        RECT 51.355 126.540 51.675 126.600 ;
        RECT 52.825 126.540 52.965 126.680 ;
        RECT 44.545 126.400 52.965 126.540 ;
        RECT 60.985 126.540 61.275 126.585 ;
        RECT 63.765 126.540 64.055 126.585 ;
        RECT 65.625 126.540 65.915 126.585 ;
        RECT 60.985 126.400 65.915 126.540 ;
        RECT 34.810 126.355 35.100 126.400 ;
        RECT 39.395 126.340 39.715 126.400 ;
        RECT 51.355 126.340 51.675 126.400 ;
        RECT 60.985 126.355 61.275 126.400 ;
        RECT 63.765 126.355 64.055 126.400 ;
        RECT 65.625 126.355 65.915 126.400 ;
        RECT 69.845 126.540 69.985 126.695 ;
        RECT 79.415 126.680 79.735 126.740 ;
        RECT 85.855 126.880 86.175 126.940 ;
        RECT 90.930 126.880 91.220 126.925 ;
        RECT 85.855 126.740 91.220 126.880 ;
        RECT 85.855 126.680 86.175 126.740 ;
        RECT 90.930 126.695 91.220 126.740 ;
        RECT 93.215 126.880 93.535 126.940 ;
        RECT 96.525 126.880 96.665 127.035 ;
        RECT 93.215 126.740 96.665 126.880 ;
        RECT 98.825 126.880 98.965 127.035 ;
        RECT 99.655 127.020 99.975 127.280 ;
        RECT 103.425 126.880 103.565 127.420 ;
        RECT 105.175 127.360 105.495 127.420 ;
        RECT 103.810 127.035 104.100 127.265 ;
        RECT 98.825 126.740 103.565 126.880 ;
        RECT 93.215 126.680 93.535 126.740 ;
        RECT 78.955 126.540 79.275 126.600 ;
        RECT 69.845 126.400 79.275 126.540 ;
        RECT 32.495 126.200 32.815 126.260 ;
        RECT 35.270 126.200 35.560 126.245 ;
        RECT 32.495 126.060 35.560 126.200 ;
        RECT 32.495 126.000 32.815 126.060 ;
        RECT 35.270 126.015 35.560 126.060 ;
        RECT 45.375 126.200 45.695 126.260 ;
        RECT 47.230 126.200 47.520 126.245 ;
        RECT 45.375 126.060 47.520 126.200 ;
        RECT 45.375 126.000 45.695 126.060 ;
        RECT 47.230 126.015 47.520 126.060 ;
        RECT 53.195 126.200 53.515 126.260 ;
        RECT 69.845 126.200 69.985 126.400 ;
        RECT 78.955 126.340 79.275 126.400 ;
        RECT 87.665 126.540 87.955 126.585 ;
        RECT 90.445 126.540 90.735 126.585 ;
        RECT 92.305 126.540 92.595 126.585 ;
        RECT 87.665 126.400 92.595 126.540 ;
        RECT 87.665 126.355 87.955 126.400 ;
        RECT 90.445 126.355 90.735 126.400 ;
        RECT 92.305 126.355 92.595 126.400 ;
        RECT 92.755 126.540 93.075 126.600 ;
        RECT 95.055 126.540 95.375 126.600 ;
        RECT 92.755 126.400 95.375 126.540 ;
        RECT 92.755 126.340 93.075 126.400 ;
        RECT 95.055 126.340 95.375 126.400 ;
        RECT 100.575 126.540 100.895 126.600 ;
        RECT 103.885 126.540 104.025 127.035 ;
        RECT 100.575 126.400 104.025 126.540 ;
        RECT 100.575 126.340 100.895 126.400 ;
        RECT 53.195 126.060 69.985 126.200 ;
        RECT 53.195 126.000 53.515 126.060 ;
        RECT 72.975 126.000 73.295 126.260 ;
        RECT 89.995 126.200 90.315 126.260 ;
        RECT 93.230 126.200 93.520 126.245 ;
        RECT 89.995 126.060 93.520 126.200 ;
        RECT 89.995 126.000 90.315 126.060 ;
        RECT 93.230 126.015 93.520 126.060 ;
        RECT 94.595 126.200 94.915 126.260 ;
        RECT 104.270 126.200 104.560 126.245 ;
        RECT 94.595 126.060 104.560 126.200 ;
        RECT 94.595 126.000 94.915 126.060 ;
        RECT 104.270 126.015 104.560 126.060 ;
        RECT 17.605 125.380 112.465 125.860 ;
        RECT 30.195 125.180 30.515 125.240 ;
        RECT 35.270 125.180 35.560 125.225 ;
        RECT 30.195 125.040 35.560 125.180 ;
        RECT 30.195 124.980 30.515 125.040 ;
        RECT 35.270 124.995 35.560 125.040 ;
        RECT 37.570 124.995 37.860 125.225 ;
        RECT 42.615 125.180 42.935 125.240 ;
        RECT 56.875 125.180 57.195 125.240 ;
        RECT 66.535 125.180 66.855 125.240 ;
        RECT 42.615 125.040 48.365 125.180 ;
        RECT 37.645 124.840 37.785 124.995 ;
        RECT 42.615 124.980 42.935 125.040 ;
        RECT 39.395 124.840 39.715 124.900 ;
        RECT 37.645 124.700 39.715 124.840 ;
        RECT 39.395 124.640 39.715 124.700 ;
        RECT 40.890 124.840 41.180 124.885 ;
        RECT 44.010 124.840 44.300 124.885 ;
        RECT 45.900 124.840 46.190 124.885 ;
        RECT 40.890 124.700 46.190 124.840 ;
        RECT 40.890 124.655 41.180 124.700 ;
        RECT 44.010 124.655 44.300 124.700 ;
        RECT 45.900 124.655 46.190 124.700 ;
        RECT 26.055 124.300 26.375 124.560 ;
        RECT 31.590 124.500 31.880 124.545 ;
        RECT 33.415 124.500 33.735 124.560 ;
        RECT 36.635 124.500 36.955 124.560 ;
        RECT 31.590 124.360 36.955 124.500 ;
        RECT 31.590 124.315 31.880 124.360 ;
        RECT 33.415 124.300 33.735 124.360 ;
        RECT 36.635 124.300 36.955 124.360 ;
        RECT 37.095 124.300 37.415 124.560 ;
        RECT 43.075 124.500 43.395 124.560 ;
        RECT 37.645 124.360 43.395 124.500 ;
        RECT 21.455 123.960 21.775 124.220 ;
        RECT 28.830 124.160 29.120 124.205 ;
        RECT 32.035 124.160 32.355 124.220 ;
        RECT 32.510 124.160 32.800 124.205 ;
        RECT 28.830 124.020 32.800 124.160 ;
        RECT 28.830 123.975 29.120 124.020 ;
        RECT 32.035 123.960 32.355 124.020 ;
        RECT 32.510 123.975 32.800 124.020 ;
        RECT 36.175 123.960 36.495 124.220 ;
        RECT 37.645 124.205 37.785 124.360 ;
        RECT 43.075 124.300 43.395 124.360 ;
        RECT 45.375 124.300 45.695 124.560 ;
        RECT 37.570 123.975 37.860 124.205 ;
        RECT 24.675 123.620 24.995 123.880 ;
        RECT 35.255 123.820 35.575 123.880 ;
        RECT 28.445 123.680 35.575 123.820 ;
        RECT 21.915 123.280 22.235 123.540 ;
        RECT 24.230 123.480 24.520 123.525 ;
        RECT 28.445 123.480 28.585 123.680 ;
        RECT 35.255 123.620 35.575 123.680 ;
        RECT 35.715 123.820 36.035 123.880 ;
        RECT 39.810 123.865 40.100 124.180 ;
        RECT 40.890 124.160 41.180 124.205 ;
        RECT 44.470 124.160 44.760 124.205 ;
        RECT 46.305 124.160 46.595 124.205 ;
        RECT 40.890 124.020 46.595 124.160 ;
        RECT 40.890 123.975 41.180 124.020 ;
        RECT 44.470 123.975 44.760 124.020 ;
        RECT 46.305 123.975 46.595 124.020 ;
        RECT 46.770 123.975 47.060 124.205 ;
        RECT 47.230 124.160 47.520 124.205 ;
        RECT 47.675 124.160 47.995 124.220 ;
        RECT 47.230 124.020 47.995 124.160 ;
        RECT 48.225 124.160 48.365 125.040 ;
        RECT 56.875 125.040 66.855 125.180 ;
        RECT 56.875 124.980 57.195 125.040 ;
        RECT 62.395 124.840 62.715 124.900 ;
        RECT 62.395 124.700 63.545 124.840 ;
        RECT 62.395 124.640 62.715 124.700 ;
        RECT 48.595 124.500 48.915 124.560 ;
        RECT 60.555 124.500 60.875 124.560 ;
        RECT 48.595 124.360 58.485 124.500 ;
        RECT 48.595 124.300 48.915 124.360 ;
        RECT 56.875 124.160 57.195 124.220 ;
        RECT 58.345 124.205 58.485 124.360 ;
        RECT 60.555 124.360 63.085 124.500 ;
        RECT 60.555 124.300 60.875 124.360 ;
        RECT 48.225 124.020 57.195 124.160 ;
        RECT 47.230 123.975 47.520 124.020 ;
        RECT 39.510 123.820 40.100 123.865 ;
        RECT 42.750 123.820 43.400 123.865 ;
        RECT 35.715 123.680 43.400 123.820 ;
        RECT 46.845 123.820 46.985 123.975 ;
        RECT 47.675 123.960 47.995 124.020 ;
        RECT 56.875 123.960 57.195 124.020 ;
        RECT 57.810 123.975 58.100 124.205 ;
        RECT 58.270 123.975 58.560 124.205 ;
        RECT 55.955 123.820 56.275 123.880 ;
        RECT 46.845 123.680 56.275 123.820 ;
        RECT 57.885 123.820 58.025 123.975 ;
        RECT 58.715 123.960 59.035 124.220 ;
        RECT 61.015 124.160 61.335 124.220 ;
        RECT 59.265 124.020 61.335 124.160 ;
        RECT 59.265 123.820 59.405 124.020 ;
        RECT 61.015 123.960 61.335 124.020 ;
        RECT 62.395 123.960 62.715 124.220 ;
        RECT 62.945 124.205 63.085 124.360 ;
        RECT 63.405 124.205 63.545 124.700 ;
        RECT 64.325 124.205 64.465 125.040 ;
        RECT 66.535 124.980 66.855 125.040 ;
        RECT 71.595 124.980 71.915 125.240 ;
        RECT 79.415 125.180 79.735 125.240 ;
        RECT 81.040 125.180 81.330 125.225 ;
        RECT 79.415 125.040 81.330 125.180 ;
        RECT 79.415 124.980 79.735 125.040 ;
        RECT 81.040 124.995 81.330 125.040 ;
        RECT 72.535 124.840 72.825 124.885 ;
        RECT 74.395 124.840 74.685 124.885 ;
        RECT 77.175 124.840 77.465 124.885 ;
        RECT 72.535 124.700 77.465 124.840 ;
        RECT 81.115 124.840 81.255 124.995 ;
        RECT 85.855 124.980 86.175 125.240 ;
        RECT 87.695 125.180 88.015 125.240 ;
        RECT 98.735 125.180 99.055 125.240 ;
        RECT 87.695 125.040 99.055 125.180 ;
        RECT 87.695 124.980 88.015 125.040 ;
        RECT 98.735 124.980 99.055 125.040 ;
        RECT 84.015 124.840 84.335 124.900 ;
        RECT 87.785 124.840 87.925 124.980 ;
        RECT 81.115 124.700 83.325 124.840 ;
        RECT 72.535 124.655 72.825 124.700 ;
        RECT 74.395 124.655 74.685 124.700 ;
        RECT 77.175 124.655 77.465 124.700 ;
        RECT 66.995 124.500 67.315 124.560 ;
        RECT 68.850 124.500 69.140 124.545 ;
        RECT 72.975 124.500 73.295 124.560 ;
        RECT 73.910 124.500 74.200 124.545 ;
        RECT 66.995 124.360 71.825 124.500 ;
        RECT 66.995 124.300 67.315 124.360 ;
        RECT 68.850 124.315 69.140 124.360 ;
        RECT 62.870 123.975 63.160 124.205 ;
        RECT 63.330 123.975 63.620 124.205 ;
        RECT 64.250 123.975 64.540 124.205 ;
        RECT 69.770 123.820 70.060 123.865 ;
        RECT 57.885 123.680 59.405 123.820 ;
        RECT 59.725 123.680 70.060 123.820 ;
        RECT 35.715 123.620 36.035 123.680 ;
        RECT 39.510 123.635 39.800 123.680 ;
        RECT 42.750 123.635 43.400 123.680 ;
        RECT 55.955 123.620 56.275 123.680 ;
        RECT 24.230 123.340 28.585 123.480 ;
        RECT 32.050 123.480 32.340 123.525 ;
        RECT 33.415 123.480 33.735 123.540 ;
        RECT 32.050 123.340 33.735 123.480 ;
        RECT 24.230 123.295 24.520 123.340 ;
        RECT 32.050 123.295 32.340 123.340 ;
        RECT 33.415 123.280 33.735 123.340 ;
        RECT 33.875 123.480 34.195 123.540 ;
        RECT 34.350 123.480 34.640 123.525 ;
        RECT 33.875 123.340 34.640 123.480 ;
        RECT 33.875 123.280 34.195 123.340 ;
        RECT 34.350 123.295 34.640 123.340 ;
        RECT 36.635 123.480 36.955 123.540 ;
        RECT 38.015 123.480 38.335 123.540 ;
        RECT 36.635 123.340 38.335 123.480 ;
        RECT 36.635 123.280 36.955 123.340 ;
        RECT 38.015 123.280 38.335 123.340 ;
        RECT 44.455 123.480 44.775 123.540 ;
        RECT 59.725 123.480 59.865 123.680 ;
        RECT 69.770 123.635 70.060 123.680 ;
        RECT 44.455 123.340 59.865 123.480 ;
        RECT 60.110 123.480 60.400 123.525 ;
        RECT 60.555 123.480 60.875 123.540 ;
        RECT 60.110 123.340 60.875 123.480 ;
        RECT 44.455 123.280 44.775 123.340 ;
        RECT 60.110 123.295 60.400 123.340 ;
        RECT 60.555 123.280 60.875 123.340 ;
        RECT 61.015 123.280 61.335 123.540 ;
        RECT 63.775 123.480 64.095 123.540 ;
        RECT 65.615 123.480 65.935 123.540 ;
        RECT 63.775 123.340 65.935 123.480 ;
        RECT 63.775 123.280 64.095 123.340 ;
        RECT 65.615 123.280 65.935 123.340 ;
        RECT 68.375 123.480 68.695 123.540 ;
        RECT 69.310 123.480 69.600 123.525 ;
        RECT 71.135 123.480 71.455 123.540 ;
        RECT 68.375 123.340 71.455 123.480 ;
        RECT 71.685 123.480 71.825 124.360 ;
        RECT 72.975 124.360 74.200 124.500 ;
        RECT 72.975 124.300 73.295 124.360 ;
        RECT 73.910 124.315 74.200 124.360 ;
        RECT 78.955 124.500 79.275 124.560 ;
        RECT 82.650 124.500 82.940 124.545 ;
        RECT 78.955 124.360 82.940 124.500 ;
        RECT 78.955 124.300 79.275 124.360 ;
        RECT 82.650 124.315 82.940 124.360 ;
        RECT 83.185 124.220 83.325 124.700 ;
        RECT 84.015 124.700 87.925 124.840 ;
        RECT 88.155 124.840 88.475 124.900 ;
        RECT 89.535 124.840 89.855 124.900 ;
        RECT 88.155 124.700 89.855 124.840 ;
        RECT 84.015 124.640 84.335 124.700 ;
        RECT 88.155 124.640 88.475 124.700 ;
        RECT 89.535 124.640 89.855 124.700 ;
        RECT 93.675 124.640 93.995 124.900 ;
        RECT 96.450 124.840 96.740 124.885 ;
        RECT 97.355 124.840 97.675 124.900 ;
        RECT 96.450 124.700 97.675 124.840 ;
        RECT 96.450 124.655 96.740 124.700 ;
        RECT 97.355 124.640 97.675 124.700 ;
        RECT 99.770 124.840 100.060 124.885 ;
        RECT 102.890 124.840 103.180 124.885 ;
        RECT 104.780 124.840 105.070 124.885 ;
        RECT 99.770 124.700 105.070 124.840 ;
        RECT 99.770 124.655 100.060 124.700 ;
        RECT 102.890 124.655 103.180 124.700 ;
        RECT 104.780 124.655 105.070 124.700 ;
        RECT 83.555 124.500 83.875 124.560 ;
        RECT 86.315 124.500 86.635 124.560 ;
        RECT 93.215 124.500 93.535 124.560 ;
        RECT 83.555 124.360 86.635 124.500 ;
        RECT 83.555 124.300 83.875 124.360 ;
        RECT 86.315 124.300 86.635 124.360 ;
        RECT 87.785 124.360 93.535 124.500 ;
        RECT 93.765 124.500 93.905 124.640 ;
        RECT 100.575 124.500 100.895 124.560 ;
        RECT 93.765 124.360 100.895 124.500 ;
        RECT 87.785 124.220 87.925 124.360 ;
        RECT 93.215 124.300 93.535 124.360 ;
        RECT 100.575 124.300 100.895 124.360 ;
        RECT 103.795 124.500 104.115 124.560 ;
        RECT 105.650 124.500 105.940 124.545 ;
        RECT 103.795 124.360 105.940 124.500 ;
        RECT 103.795 124.300 104.115 124.360 ;
        RECT 105.650 124.315 105.940 124.360 ;
        RECT 72.070 124.160 72.360 124.205 ;
        RECT 72.515 124.160 72.835 124.220 ;
        RECT 77.175 124.160 77.465 124.205 ;
        RECT 72.070 124.020 72.835 124.160 ;
        RECT 72.070 123.975 72.360 124.020 ;
        RECT 72.515 123.960 72.835 124.020 ;
        RECT 74.930 124.020 77.465 124.160 ;
        RECT 74.930 123.865 75.145 124.020 ;
        RECT 77.175 123.975 77.465 124.020 ;
        RECT 83.095 124.160 83.415 124.220 ;
        RECT 84.030 124.160 84.320 124.205 ;
        RECT 83.095 124.020 84.320 124.160 ;
        RECT 83.095 123.960 83.415 124.020 ;
        RECT 84.030 123.975 84.320 124.020 ;
        RECT 87.695 123.960 88.015 124.220 ;
        RECT 88.630 123.975 88.920 124.205 ;
        RECT 89.090 123.975 89.380 124.205 ;
        RECT 72.995 123.820 73.285 123.865 ;
        RECT 74.855 123.820 75.145 123.865 ;
        RECT 72.995 123.680 75.145 123.820 ;
        RECT 72.995 123.635 73.285 123.680 ;
        RECT 74.855 123.635 75.145 123.680 ;
        RECT 75.735 123.865 76.055 123.880 ;
        RECT 75.735 123.820 76.065 123.865 ;
        RECT 79.035 123.820 79.325 123.865 ;
        RECT 75.735 123.680 79.325 123.820 ;
        RECT 75.735 123.635 76.065 123.680 ;
        RECT 79.035 123.635 79.325 123.680 ;
        RECT 79.875 123.820 80.195 123.880 ;
        RECT 88.705 123.820 88.845 123.975 ;
        RECT 79.875 123.680 88.845 123.820 ;
        RECT 75.735 123.620 76.055 123.635 ;
        RECT 79.875 123.620 80.195 123.680 ;
        RECT 80.795 123.480 81.115 123.540 ;
        RECT 71.685 123.340 81.115 123.480 ;
        RECT 68.375 123.280 68.695 123.340 ;
        RECT 69.310 123.295 69.600 123.340 ;
        RECT 71.135 123.280 71.455 123.340 ;
        RECT 80.795 123.280 81.115 123.340 ;
        RECT 84.475 123.480 84.795 123.540 ;
        RECT 88.155 123.480 88.475 123.540 ;
        RECT 84.475 123.340 88.475 123.480 ;
        RECT 84.475 123.280 84.795 123.340 ;
        RECT 88.155 123.280 88.475 123.340 ;
        RECT 88.615 123.480 88.935 123.540 ;
        RECT 89.165 123.480 89.305 123.975 ;
        RECT 89.535 123.960 89.855 124.220 ;
        RECT 93.690 124.160 93.980 124.205 ;
        RECT 93.690 124.020 96.665 124.160 ;
        RECT 93.690 123.975 93.980 124.020 ;
        RECT 96.525 123.540 96.665 124.020 ;
        RECT 98.690 123.865 98.980 124.180 ;
        RECT 99.770 124.160 100.060 124.205 ;
        RECT 103.350 124.160 103.640 124.205 ;
        RECT 105.185 124.160 105.475 124.205 ;
        RECT 99.770 124.020 105.475 124.160 ;
        RECT 99.770 123.975 100.060 124.020 ;
        RECT 103.350 123.975 103.640 124.020 ;
        RECT 105.185 123.975 105.475 124.020 ;
        RECT 98.390 123.820 98.980 123.865 ;
        RECT 101.630 123.820 102.280 123.865 ;
        RECT 102.875 123.820 103.195 123.880 ;
        RECT 104.270 123.820 104.560 123.865 ;
        RECT 98.390 123.680 102.645 123.820 ;
        RECT 98.390 123.635 98.680 123.680 ;
        RECT 101.630 123.635 102.280 123.680 ;
        RECT 88.615 123.340 89.305 123.480 ;
        RECT 90.930 123.480 91.220 123.525 ;
        RECT 91.375 123.480 91.695 123.540 ;
        RECT 90.930 123.340 91.695 123.480 ;
        RECT 88.615 123.280 88.935 123.340 ;
        RECT 90.930 123.295 91.220 123.340 ;
        RECT 91.375 123.280 91.695 123.340 ;
        RECT 92.295 123.480 92.615 123.540 ;
        RECT 95.055 123.480 95.375 123.540 ;
        RECT 92.295 123.340 95.375 123.480 ;
        RECT 92.295 123.280 92.615 123.340 ;
        RECT 95.055 123.280 95.375 123.340 ;
        RECT 96.435 123.480 96.755 123.540 ;
        RECT 96.910 123.480 97.200 123.525 ;
        RECT 96.435 123.340 97.200 123.480 ;
        RECT 102.505 123.480 102.645 123.680 ;
        RECT 102.875 123.680 104.560 123.820 ;
        RECT 102.875 123.620 103.195 123.680 ;
        RECT 104.270 123.635 104.560 123.680 ;
        RECT 103.795 123.480 104.115 123.540 ;
        RECT 102.505 123.340 104.115 123.480 ;
        RECT 96.435 123.280 96.755 123.340 ;
        RECT 96.910 123.295 97.200 123.340 ;
        RECT 103.795 123.280 104.115 123.340 ;
        RECT 18.165 122.660 112.465 123.140 ;
        RECT 21.915 122.460 22.235 122.520 ;
        RECT 33.415 122.460 33.735 122.520 ;
        RECT 38.015 122.460 38.335 122.520 ;
        RECT 38.950 122.460 39.240 122.505 ;
        RECT 21.915 122.320 32.495 122.460 ;
        RECT 21.915 122.260 22.235 122.320 ;
        RECT 26.055 122.120 26.375 122.180 ;
        RECT 26.055 121.980 27.665 122.120 ;
        RECT 26.055 121.920 26.375 121.980 ;
        RECT 24.215 121.780 24.535 121.840 ;
        RECT 24.690 121.780 24.980 121.825 ;
        RECT 24.215 121.640 24.980 121.780 ;
        RECT 24.215 121.580 24.535 121.640 ;
        RECT 24.690 121.595 24.980 121.640 ;
        RECT 26.515 121.580 26.835 121.840 ;
        RECT 27.525 121.825 27.665 121.980 ;
        RECT 31.575 121.920 31.895 122.180 ;
        RECT 32.355 122.120 32.495 122.320 ;
        RECT 33.415 122.320 39.240 122.460 ;
        RECT 33.415 122.260 33.735 122.320 ;
        RECT 38.015 122.260 38.335 122.320 ;
        RECT 38.950 122.275 39.240 122.320 ;
        RECT 43.090 122.460 43.380 122.505 ;
        RECT 44.455 122.460 44.775 122.520 ;
        RECT 43.090 122.320 44.775 122.460 ;
        RECT 43.090 122.275 43.380 122.320 ;
        RECT 33.870 122.120 34.520 122.165 ;
        RECT 37.470 122.120 37.760 122.165 ;
        RECT 32.355 121.980 37.760 122.120 ;
        RECT 33.870 121.935 34.520 121.980 ;
        RECT 37.170 121.935 37.760 121.980 ;
        RECT 27.450 121.595 27.740 121.825 ;
        RECT 27.895 121.580 28.215 121.840 ;
        RECT 28.355 121.580 28.675 121.840 ;
        RECT 30.675 121.780 30.965 121.825 ;
        RECT 32.510 121.780 32.800 121.825 ;
        RECT 36.090 121.780 36.380 121.825 ;
        RECT 30.675 121.640 36.380 121.780 ;
        RECT 30.675 121.595 30.965 121.640 ;
        RECT 32.510 121.595 32.800 121.640 ;
        RECT 36.090 121.595 36.380 121.640 ;
        RECT 37.170 121.620 37.460 121.935 ;
        RECT 39.025 121.780 39.165 122.275 ;
        RECT 44.455 122.260 44.775 122.320 ;
        RECT 44.930 122.460 45.220 122.505 ;
        RECT 45.375 122.460 45.695 122.520 ;
        RECT 44.930 122.320 45.695 122.460 ;
        RECT 44.930 122.275 45.220 122.320 ;
        RECT 45.375 122.260 45.695 122.320 ;
        RECT 46.755 122.460 47.075 122.520 ;
        RECT 47.230 122.460 47.520 122.505 ;
        RECT 46.755 122.320 47.520 122.460 ;
        RECT 46.755 122.260 47.075 122.320 ;
        RECT 47.230 122.275 47.520 122.320 ;
        RECT 50.895 122.460 51.215 122.520 ;
        RECT 51.830 122.460 52.120 122.505 ;
        RECT 50.895 122.320 52.120 122.460 ;
        RECT 50.895 122.260 51.215 122.320 ;
        RECT 51.830 122.275 52.120 122.320 ;
        RECT 58.270 122.460 58.560 122.505 ;
        RECT 66.550 122.460 66.840 122.505 ;
        RECT 68.375 122.460 68.695 122.520 ;
        RECT 58.270 122.320 64.465 122.460 ;
        RECT 58.270 122.275 58.560 122.320 ;
        RECT 51.370 122.120 51.660 122.165 ;
        RECT 58.345 122.120 58.485 122.275 ;
        RECT 51.370 121.980 58.485 122.120 ;
        RECT 59.635 122.120 59.955 122.180 ;
        RECT 64.325 122.120 64.465 122.320 ;
        RECT 66.550 122.320 68.695 122.460 ;
        RECT 66.550 122.275 66.840 122.320 ;
        RECT 68.375 122.260 68.695 122.320 ;
        RECT 69.295 122.460 69.615 122.520 ;
        RECT 75.290 122.460 75.580 122.505 ;
        RECT 69.295 122.320 75.580 122.460 ;
        RECT 69.295 122.260 69.615 122.320 ;
        RECT 75.290 122.275 75.580 122.320 ;
        RECT 78.955 122.460 79.275 122.520 ;
        RECT 80.810 122.460 81.100 122.505 ;
        RECT 78.955 122.320 81.100 122.460 ;
        RECT 78.955 122.260 79.275 122.320 ;
        RECT 80.810 122.275 81.100 122.320 ;
        RECT 85.025 122.320 86.085 122.460 ;
        RECT 68.850 122.120 69.140 122.165 ;
        RECT 77.575 122.120 77.895 122.180 ;
        RECT 79.430 122.120 79.720 122.165 ;
        RECT 59.635 121.980 64.005 122.120 ;
        RECT 64.325 121.980 69.140 122.120 ;
        RECT 51.370 121.935 51.660 121.980 ;
        RECT 59.635 121.920 59.955 121.980 ;
        RECT 39.870 121.780 40.160 121.825 ;
        RECT 39.025 121.640 40.160 121.780 ;
        RECT 39.870 121.595 40.160 121.640 ;
        RECT 42.615 121.780 42.935 121.840 ;
        RECT 44.915 121.780 45.235 121.840 ;
        RECT 45.390 121.780 45.680 121.825 ;
        RECT 42.615 121.640 45.680 121.780 ;
        RECT 42.615 121.580 42.935 121.640 ;
        RECT 44.915 121.580 45.235 121.640 ;
        RECT 45.390 121.595 45.680 121.640 ;
        RECT 49.530 121.780 49.820 121.825 ;
        RECT 52.735 121.780 53.055 121.840 ;
        RECT 61.565 121.825 61.705 121.980 ;
        RECT 49.530 121.640 53.055 121.780 ;
        RECT 49.530 121.595 49.820 121.640 ;
        RECT 52.735 121.580 53.055 121.640 ;
        RECT 61.030 121.595 61.320 121.825 ;
        RECT 61.490 121.595 61.780 121.825 ;
        RECT 30.195 121.240 30.515 121.500 ;
        RECT 35.255 121.440 35.575 121.500 ;
        RECT 41.235 121.440 41.555 121.500 ;
        RECT 35.255 121.300 41.555 121.440 ;
        RECT 35.255 121.240 35.575 121.300 ;
        RECT 41.235 121.240 41.555 121.300 ;
        RECT 44.470 121.440 44.760 121.485 ;
        RECT 50.910 121.440 51.200 121.485 ;
        RECT 51.355 121.440 51.675 121.500 ;
        RECT 44.470 121.300 51.675 121.440 ;
        RECT 44.470 121.255 44.760 121.300 ;
        RECT 50.910 121.255 51.200 121.300 ;
        RECT 51.355 121.240 51.675 121.300 ;
        RECT 51.815 121.440 52.135 121.500 ;
        RECT 55.050 121.440 55.340 121.485 ;
        RECT 51.815 121.300 55.340 121.440 ;
        RECT 61.105 121.440 61.245 121.595 ;
        RECT 61.935 121.580 62.255 121.840 ;
        RECT 62.855 121.580 63.175 121.840 ;
        RECT 63.865 121.780 64.005 121.980 ;
        RECT 68.850 121.935 69.140 121.980 ;
        RECT 72.605 121.980 77.345 122.120 ;
        RECT 66.535 121.795 66.855 121.840 ;
        RECT 66.535 121.780 66.995 121.795 ;
        RECT 72.605 121.780 72.745 121.980 ;
        RECT 75.365 121.840 75.505 121.980 ;
        RECT 63.865 121.640 65.385 121.780 ;
        RECT 62.395 121.440 62.715 121.500 ;
        RECT 63.775 121.440 64.095 121.500 ;
        RECT 61.105 121.300 62.165 121.440 ;
        RECT 51.815 121.240 52.135 121.300 ;
        RECT 55.050 121.255 55.340 121.300 ;
        RECT 62.025 121.160 62.165 121.300 ;
        RECT 62.395 121.300 64.095 121.440 ;
        RECT 65.245 121.440 65.385 121.640 ;
        RECT 66.535 121.640 72.745 121.780 ;
        RECT 66.535 121.580 66.855 121.640 ;
        RECT 72.975 121.580 73.295 121.840 ;
        RECT 73.895 121.580 74.215 121.840 ;
        RECT 75.275 121.580 75.595 121.840 ;
        RECT 77.205 121.780 77.345 121.980 ;
        RECT 77.575 121.980 79.720 122.120 ;
        RECT 77.575 121.920 77.895 121.980 ;
        RECT 79.430 121.935 79.720 121.980 ;
        RECT 83.095 122.120 83.415 122.180 ;
        RECT 85.025 122.120 85.165 122.320 ;
        RECT 83.095 121.980 85.165 122.120 ;
        RECT 83.095 121.920 83.415 121.980 ;
        RECT 84.475 121.810 84.795 121.840 ;
        RECT 84.105 121.780 84.795 121.810 ;
        RECT 77.205 121.670 84.795 121.780 ;
        RECT 77.205 121.640 84.245 121.670 ;
        RECT 84.475 121.580 84.795 121.670 ;
        RECT 84.935 121.580 85.255 121.840 ;
        RECT 85.515 121.780 85.805 121.825 ;
        RECT 85.945 121.780 86.085 122.320 ;
        RECT 86.315 122.260 86.635 122.520 ;
        RECT 87.695 122.460 88.015 122.520 ;
        RECT 87.695 122.320 90.225 122.460 ;
        RECT 87.695 122.260 88.015 122.320 ;
        RECT 86.405 122.120 86.545 122.260 ;
        RECT 86.405 121.980 89.305 122.120 ;
        RECT 85.515 121.640 86.085 121.780 ;
        RECT 86.315 121.780 86.635 121.840 ;
        RECT 87.695 121.780 88.015 121.840 ;
        RECT 86.315 121.640 88.015 121.780 ;
        RECT 85.515 121.595 85.805 121.640 ;
        RECT 86.315 121.580 86.635 121.640 ;
        RECT 87.695 121.580 88.015 121.640 ;
        RECT 88.155 121.580 88.475 121.840 ;
        RECT 88.615 121.580 88.935 121.840 ;
        RECT 89.165 121.825 89.305 121.980 ;
        RECT 90.085 121.825 90.225 122.320 ;
        RECT 102.875 122.260 103.195 122.520 ;
        RECT 103.795 122.260 104.115 122.520 ;
        RECT 96.435 122.120 96.755 122.180 ;
        RECT 92.385 121.980 96.755 122.120 ;
        RECT 89.090 121.595 89.380 121.825 ;
        RECT 90.010 121.780 90.300 121.825 ;
        RECT 91.390 121.780 91.680 121.825 ;
        RECT 91.835 121.780 92.155 121.840 ;
        RECT 92.385 121.825 92.525 121.980 ;
        RECT 96.435 121.920 96.755 121.980 ;
        RECT 90.010 121.640 92.155 121.780 ;
        RECT 90.010 121.595 90.300 121.640 ;
        RECT 91.390 121.595 91.680 121.640 ;
        RECT 91.835 121.580 92.155 121.640 ;
        RECT 92.310 121.595 92.600 121.825 ;
        RECT 92.755 121.580 93.075 121.840 ;
        RECT 93.230 121.780 93.520 121.825 ;
        RECT 95.055 121.780 95.375 121.840 ;
        RECT 93.230 121.640 95.375 121.780 ;
        RECT 93.230 121.595 93.520 121.640 ;
        RECT 65.245 121.300 66.995 121.440 ;
        RECT 62.395 121.240 62.715 121.300 ;
        RECT 63.775 121.240 64.095 121.300 ;
        RECT 31.080 121.100 31.370 121.145 ;
        RECT 32.970 121.100 33.260 121.145 ;
        RECT 36.090 121.100 36.380 121.145 ;
        RECT 31.080 120.960 36.380 121.100 ;
        RECT 31.080 120.915 31.370 120.960 ;
        RECT 32.970 120.915 33.260 120.960 ;
        RECT 36.090 120.915 36.380 120.960 ;
        RECT 61.935 120.900 62.255 121.160 ;
        RECT 66.855 121.100 66.995 121.300 ;
        RECT 69.295 121.240 69.615 121.500 ;
        RECT 70.230 121.440 70.520 121.485 ;
        RECT 70.675 121.440 70.995 121.500 ;
        RECT 72.515 121.440 72.835 121.500 ;
        RECT 70.230 121.300 72.835 121.440 ;
        RECT 73.065 121.440 73.205 121.580 ;
        RECT 74.815 121.440 75.135 121.500 ;
        RECT 73.065 121.300 75.135 121.440 ;
        RECT 70.230 121.255 70.520 121.300 ;
        RECT 70.675 121.240 70.995 121.300 ;
        RECT 72.515 121.240 72.835 121.300 ;
        RECT 74.815 121.240 75.135 121.300 ;
        RECT 78.495 121.240 78.815 121.500 ;
        RECT 79.875 121.440 80.195 121.500 ;
        RECT 84.015 121.440 84.335 121.500 ;
        RECT 79.875 121.300 84.335 121.440 ;
        RECT 79.875 121.240 80.195 121.300 ;
        RECT 84.015 121.240 84.335 121.300 ;
        RECT 76.195 121.100 76.515 121.160 ;
        RECT 84.935 121.100 85.255 121.160 ;
        RECT 88.705 121.100 88.845 121.580 ;
        RECT 89.535 121.440 89.855 121.500 ;
        RECT 93.305 121.440 93.445 121.595 ;
        RECT 95.055 121.580 95.375 121.640 ;
        RECT 96.910 121.780 97.200 121.825 ;
        RECT 97.355 121.780 97.675 121.840 ;
        RECT 96.910 121.640 97.675 121.780 ;
        RECT 96.910 121.595 97.200 121.640 ;
        RECT 97.355 121.580 97.675 121.640 ;
        RECT 101.495 121.780 101.815 121.840 ;
        RECT 103.350 121.780 103.640 121.825 ;
        RECT 101.495 121.640 103.640 121.780 ;
        RECT 101.495 121.580 101.815 121.640 ;
        RECT 103.350 121.595 103.640 121.640 ;
        RECT 94.595 121.440 94.915 121.500 ;
        RECT 95.530 121.440 95.820 121.485 ;
        RECT 89.535 121.300 93.445 121.440 ;
        RECT 93.765 121.300 95.820 121.440 ;
        RECT 89.535 121.240 89.855 121.300 ;
        RECT 66.855 120.960 88.845 121.100 ;
        RECT 76.195 120.900 76.515 120.960 ;
        RECT 84.935 120.900 85.255 120.960 ;
        RECT 24.230 120.760 24.520 120.805 ;
        RECT 24.675 120.760 24.995 120.820 ;
        RECT 24.230 120.620 24.995 120.760 ;
        RECT 24.230 120.575 24.520 120.620 ;
        RECT 24.675 120.560 24.995 120.620 ;
        RECT 29.735 120.560 30.055 120.820 ;
        RECT 49.055 120.560 49.375 120.820 ;
        RECT 53.670 120.760 53.960 120.805 ;
        RECT 55.495 120.760 55.815 120.820 ;
        RECT 53.670 120.620 55.815 120.760 ;
        RECT 53.670 120.575 53.960 120.620 ;
        RECT 55.495 120.560 55.815 120.620 ;
        RECT 59.650 120.760 59.940 120.805 ;
        RECT 64.235 120.760 64.555 120.820 ;
        RECT 59.650 120.620 64.555 120.760 ;
        RECT 59.650 120.575 59.940 120.620 ;
        RECT 64.235 120.560 64.555 120.620 ;
        RECT 67.010 120.760 67.300 120.805 ;
        RECT 67.455 120.760 67.775 120.820 ;
        RECT 67.010 120.620 67.775 120.760 ;
        RECT 67.010 120.575 67.300 120.620 ;
        RECT 67.455 120.560 67.775 120.620 ;
        RECT 74.370 120.760 74.660 120.805 ;
        RECT 75.735 120.760 76.055 120.820 ;
        RECT 74.370 120.620 76.055 120.760 ;
        RECT 74.370 120.575 74.660 120.620 ;
        RECT 75.735 120.560 76.055 120.620 ;
        RECT 81.255 120.760 81.575 120.820 ;
        RECT 83.110 120.760 83.400 120.805 ;
        RECT 81.255 120.620 83.400 120.760 ;
        RECT 81.255 120.560 81.575 120.620 ;
        RECT 83.110 120.575 83.400 120.620 ;
        RECT 84.475 120.760 84.795 120.820 ;
        RECT 86.790 120.760 87.080 120.805 ;
        RECT 84.475 120.620 87.080 120.760 ;
        RECT 84.475 120.560 84.795 120.620 ;
        RECT 86.790 120.575 87.080 120.620 ;
        RECT 92.295 120.760 92.615 120.820 ;
        RECT 93.765 120.760 93.905 121.300 ;
        RECT 94.595 121.240 94.915 121.300 ;
        RECT 95.530 121.255 95.820 121.300 ;
        RECT 99.670 121.255 99.960 121.485 ;
        RECT 98.750 121.100 99.040 121.145 ;
        RECT 99.745 121.100 99.885 121.255 ;
        RECT 98.750 120.960 99.885 121.100 ;
        RECT 98.750 120.915 99.040 120.960 ;
        RECT 92.295 120.620 93.905 120.760 ;
        RECT 92.295 120.560 92.615 120.620 ;
        RECT 94.595 120.560 94.915 120.820 ;
        RECT 17.605 119.940 112.465 120.420 ;
        RECT 26.515 119.740 26.835 119.800 ;
        RECT 31.130 119.740 31.420 119.785 ;
        RECT 31.575 119.740 31.895 119.800 ;
        RECT 43.075 119.740 43.395 119.800 ;
        RECT 26.515 119.600 30.885 119.740 ;
        RECT 26.515 119.540 26.835 119.600 ;
        RECT 23.870 119.400 24.160 119.445 ;
        RECT 26.990 119.400 27.280 119.445 ;
        RECT 28.880 119.400 29.170 119.445 ;
        RECT 23.870 119.260 29.170 119.400 ;
        RECT 30.745 119.400 30.885 119.600 ;
        RECT 31.130 119.600 31.895 119.740 ;
        RECT 31.130 119.555 31.420 119.600 ;
        RECT 31.575 119.540 31.895 119.600 ;
        RECT 38.565 119.600 43.395 119.740 ;
        RECT 37.555 119.400 37.875 119.460 ;
        RECT 38.565 119.400 38.705 119.600 ;
        RECT 43.075 119.540 43.395 119.600 ;
        RECT 48.150 119.740 48.440 119.785 ;
        RECT 50.435 119.740 50.755 119.800 ;
        RECT 51.815 119.740 52.135 119.800 ;
        RECT 48.150 119.600 52.135 119.740 ;
        RECT 48.150 119.555 48.440 119.600 ;
        RECT 50.435 119.540 50.755 119.600 ;
        RECT 51.815 119.540 52.135 119.600 ;
        RECT 60.110 119.740 60.400 119.785 ;
        RECT 61.030 119.740 61.320 119.785 ;
        RECT 60.110 119.600 61.320 119.740 ;
        RECT 60.110 119.555 60.400 119.600 ;
        RECT 61.030 119.555 61.320 119.600 ;
        RECT 65.615 119.540 65.935 119.800 ;
        RECT 70.215 119.740 70.535 119.800 ;
        RECT 70.215 119.600 77.345 119.740 ;
        RECT 70.215 119.540 70.535 119.600 ;
        RECT 30.745 119.260 38.705 119.400 ;
        RECT 23.870 119.215 24.160 119.260 ;
        RECT 26.990 119.215 27.280 119.260 ;
        RECT 28.880 119.215 29.170 119.260 ;
        RECT 37.555 119.200 37.875 119.260 ;
        RECT 33.875 118.860 34.195 119.120 ;
        RECT 34.795 119.060 35.115 119.120 ;
        RECT 34.795 118.920 37.325 119.060 ;
        RECT 34.795 118.860 35.115 118.920 ;
        RECT 19.615 118.180 19.935 118.440 ;
        RECT 22.790 118.425 23.080 118.740 ;
        RECT 23.870 118.720 24.160 118.765 ;
        RECT 27.450 118.720 27.740 118.765 ;
        RECT 29.285 118.720 29.575 118.765 ;
        RECT 23.870 118.580 29.575 118.720 ;
        RECT 23.870 118.535 24.160 118.580 ;
        RECT 27.450 118.535 27.740 118.580 ;
        RECT 29.285 118.535 29.575 118.580 ;
        RECT 29.750 118.720 30.040 118.765 ;
        RECT 30.195 118.720 30.515 118.780 ;
        RECT 32.955 118.720 33.275 118.780 ;
        RECT 29.750 118.580 33.275 118.720 ;
        RECT 29.750 118.535 30.040 118.580 ;
        RECT 30.195 118.520 30.515 118.580 ;
        RECT 32.955 118.520 33.275 118.580 ;
        RECT 36.175 118.720 36.495 118.780 ;
        RECT 37.185 118.765 37.325 118.920 ;
        RECT 36.650 118.720 36.940 118.765 ;
        RECT 36.175 118.580 36.940 118.720 ;
        RECT 36.175 118.520 36.495 118.580 ;
        RECT 36.650 118.535 36.940 118.580 ;
        RECT 37.110 118.535 37.400 118.765 ;
        RECT 37.570 118.720 37.860 118.765 ;
        RECT 38.015 118.720 38.335 118.780 ;
        RECT 38.565 118.765 38.705 119.260 ;
        RECT 39.820 119.400 40.110 119.445 ;
        RECT 41.710 119.400 42.000 119.445 ;
        RECT 44.830 119.400 45.120 119.445 ;
        RECT 39.820 119.260 45.120 119.400 ;
        RECT 39.820 119.215 40.110 119.260 ;
        RECT 41.710 119.215 42.000 119.260 ;
        RECT 44.830 119.215 45.120 119.260 ;
        RECT 51.010 119.400 51.300 119.445 ;
        RECT 54.130 119.400 54.420 119.445 ;
        RECT 56.020 119.400 56.310 119.445 ;
        RECT 60.555 119.400 60.875 119.460 ;
        RECT 51.010 119.260 56.310 119.400 ;
        RECT 51.010 119.215 51.300 119.260 ;
        RECT 54.130 119.215 54.420 119.260 ;
        RECT 56.020 119.215 56.310 119.260 ;
        RECT 58.805 119.260 60.875 119.400 ;
        RECT 38.935 119.060 39.255 119.120 ;
        RECT 47.215 119.060 47.535 119.120 ;
        RECT 38.935 118.920 47.535 119.060 ;
        RECT 38.935 118.860 39.255 118.920 ;
        RECT 47.215 118.860 47.535 118.920 ;
        RECT 55.495 118.860 55.815 119.120 ;
        RECT 37.570 118.580 38.335 118.720 ;
        RECT 37.570 118.535 37.860 118.580 ;
        RECT 38.015 118.520 38.335 118.580 ;
        RECT 38.490 118.535 38.780 118.765 ;
        RECT 39.415 118.720 39.705 118.765 ;
        RECT 41.250 118.720 41.540 118.765 ;
        RECT 44.830 118.720 45.120 118.765 ;
        RECT 39.415 118.580 45.120 118.720 ;
        RECT 39.415 118.535 39.705 118.580 ;
        RECT 41.250 118.535 41.540 118.580 ;
        RECT 44.830 118.535 45.120 118.580 ;
        RECT 22.490 118.380 23.080 118.425 ;
        RECT 24.675 118.380 24.995 118.440 ;
        RECT 25.730 118.380 26.380 118.425 ;
        RECT 22.490 118.240 26.380 118.380 ;
        RECT 22.490 118.195 22.780 118.240 ;
        RECT 24.675 118.180 24.995 118.240 ;
        RECT 25.730 118.195 26.380 118.240 ;
        RECT 28.370 118.380 28.660 118.425 ;
        RECT 32.035 118.380 32.355 118.440 ;
        RECT 45.910 118.425 46.200 118.740 ;
        RECT 28.370 118.240 32.355 118.380 ;
        RECT 28.370 118.195 28.660 118.240 ;
        RECT 32.035 118.180 32.355 118.240 ;
        RECT 40.330 118.195 40.620 118.425 ;
        RECT 42.610 118.380 43.260 118.425 ;
        RECT 45.910 118.380 46.500 118.425 ;
        RECT 49.055 118.380 49.375 118.440 ;
        RECT 49.930 118.425 50.220 118.740 ;
        RECT 51.010 118.720 51.300 118.765 ;
        RECT 54.590 118.720 54.880 118.765 ;
        RECT 56.425 118.720 56.715 118.765 ;
        RECT 51.010 118.580 56.715 118.720 ;
        RECT 51.010 118.535 51.300 118.580 ;
        RECT 54.590 118.535 54.880 118.580 ;
        RECT 56.425 118.535 56.715 118.580 ;
        RECT 56.875 118.520 57.195 118.780 ;
        RECT 58.805 118.765 58.945 119.260 ;
        RECT 60.555 119.200 60.875 119.260 ;
        RECT 66.960 119.400 67.250 119.445 ;
        RECT 68.850 119.400 69.140 119.445 ;
        RECT 71.970 119.400 72.260 119.445 ;
        RECT 66.960 119.260 72.260 119.400 ;
        RECT 66.960 119.215 67.250 119.260 ;
        RECT 68.850 119.215 69.140 119.260 ;
        RECT 71.970 119.215 72.260 119.260 ;
        RECT 72.515 119.400 72.835 119.460 ;
        RECT 77.205 119.400 77.345 119.600 ;
        RECT 80.795 119.540 81.115 119.800 ;
        RECT 84.565 119.600 86.515 119.740 ;
        RECT 84.565 119.400 84.705 119.600 ;
        RECT 72.515 119.260 76.425 119.400 ;
        RECT 77.205 119.260 84.705 119.400 ;
        RECT 86.375 119.400 86.515 119.600 ;
        RECT 87.235 119.540 87.555 119.800 ;
        RECT 93.675 119.740 93.995 119.800 ;
        RECT 104.730 119.740 105.020 119.785 ;
        RECT 93.675 119.600 105.020 119.740 ;
        RECT 93.675 119.540 93.995 119.600 ;
        RECT 104.730 119.555 105.020 119.600 ;
        RECT 92.755 119.400 93.075 119.460 ;
        RECT 86.375 119.260 93.075 119.400 ;
        RECT 72.515 119.200 72.835 119.260 ;
        RECT 76.285 119.120 76.425 119.260 ;
        RECT 59.650 119.060 59.940 119.105 ;
        RECT 61.015 119.060 61.335 119.120 ;
        RECT 59.650 118.920 61.335 119.060 ;
        RECT 59.650 118.875 59.940 118.920 ;
        RECT 61.015 118.860 61.335 118.920 ;
        RECT 67.455 118.860 67.775 119.120 ;
        RECT 69.295 119.060 69.615 119.120 ;
        RECT 69.295 118.920 74.125 119.060 ;
        RECT 69.295 118.860 69.615 118.920 ;
        RECT 58.730 118.535 59.020 118.765 ;
        RECT 60.095 118.520 60.415 118.780 ;
        RECT 61.935 118.520 62.255 118.780 ;
        RECT 62.855 118.520 63.175 118.780 ;
        RECT 64.235 118.520 64.555 118.780 ;
        RECT 64.695 118.520 65.015 118.780 ;
        RECT 65.155 118.720 65.475 118.780 ;
        RECT 65.630 118.720 65.920 118.765 ;
        RECT 65.155 118.580 65.920 118.720 ;
        RECT 65.155 118.520 65.475 118.580 ;
        RECT 65.630 118.535 65.920 118.580 ;
        RECT 66.090 118.535 66.380 118.765 ;
        RECT 66.555 118.720 66.845 118.765 ;
        RECT 68.390 118.720 68.680 118.765 ;
        RECT 71.970 118.720 72.260 118.765 ;
        RECT 66.555 118.580 72.260 118.720 ;
        RECT 66.555 118.535 66.845 118.580 ;
        RECT 68.390 118.535 68.680 118.580 ;
        RECT 71.970 118.535 72.260 118.580 ;
        RECT 42.610 118.240 49.375 118.380 ;
        RECT 42.610 118.195 43.260 118.240 ;
        RECT 46.210 118.195 46.500 118.240 ;
        RECT 35.270 118.040 35.560 118.085 ;
        RECT 35.715 118.040 36.035 118.100 ;
        RECT 35.270 117.900 36.035 118.040 ;
        RECT 40.405 118.040 40.545 118.195 ;
        RECT 49.055 118.180 49.375 118.240 ;
        RECT 49.630 118.380 50.220 118.425 ;
        RECT 52.275 118.380 52.595 118.440 ;
        RECT 52.870 118.380 53.520 118.425 ;
        RECT 49.630 118.240 53.520 118.380 ;
        RECT 56.965 118.380 57.105 118.520 ;
        RECT 66.165 118.380 66.305 118.535 ;
        RECT 56.965 118.240 66.305 118.380 ;
        RECT 69.750 118.380 70.400 118.425 ;
        RECT 71.135 118.380 71.455 118.440 ;
        RECT 73.050 118.425 73.340 118.740 ;
        RECT 73.985 118.720 74.125 118.920 ;
        RECT 76.195 118.860 76.515 119.120 ;
        RECT 75.735 118.720 76.055 118.780 ;
        RECT 77.130 118.720 77.420 118.765 ;
        RECT 73.985 118.580 77.420 118.720 ;
        RECT 75.735 118.520 76.055 118.580 ;
        RECT 77.130 118.535 77.420 118.580 ;
        RECT 78.955 118.720 79.275 118.780 ;
        RECT 80.350 118.720 80.640 118.765 ;
        RECT 78.955 118.580 80.640 118.720 ;
        RECT 78.955 118.520 79.275 118.580 ;
        RECT 80.350 118.535 80.640 118.580 ;
        RECT 84.015 118.520 84.335 118.780 ;
        RECT 84.565 118.765 84.705 119.260 ;
        RECT 87.235 119.060 87.555 119.120 ;
        RECT 88.170 119.060 88.460 119.105 ;
        RECT 87.235 118.920 88.460 119.060 ;
        RECT 87.235 118.860 87.555 118.920 ;
        RECT 88.170 118.875 88.460 118.920 ;
        RECT 84.475 118.535 84.765 118.765 ;
        RECT 84.950 118.535 85.240 118.765 ;
        RECT 85.840 118.720 86.130 118.765 ;
        RECT 86.315 118.720 86.635 118.780 ;
        RECT 85.840 118.580 86.635 118.720 ;
        RECT 85.840 118.535 86.130 118.580 ;
        RECT 73.050 118.380 73.640 118.425 ;
        RECT 69.750 118.240 73.640 118.380 ;
        RECT 49.630 118.195 49.920 118.240 ;
        RECT 52.275 118.180 52.595 118.240 ;
        RECT 52.870 118.195 53.520 118.240 ;
        RECT 69.750 118.195 70.400 118.240 ;
        RECT 71.135 118.180 71.455 118.240 ;
        RECT 73.350 118.195 73.640 118.240 ;
        RECT 76.670 118.380 76.960 118.425 ;
        RECT 83.555 118.380 83.875 118.440 ;
        RECT 85.025 118.380 85.165 118.535 ;
        RECT 86.315 118.520 86.635 118.580 ;
        RECT 86.790 118.705 87.080 118.765 ;
        RECT 88.615 118.720 88.935 118.780 ;
        RECT 87.325 118.705 88.935 118.720 ;
        RECT 86.790 118.580 88.935 118.705 ;
        RECT 86.790 118.565 87.465 118.580 ;
        RECT 86.790 118.535 87.080 118.565 ;
        RECT 88.615 118.520 88.935 118.580 ;
        RECT 89.535 118.520 89.855 118.780 ;
        RECT 90.085 118.765 90.225 119.260 ;
        RECT 92.755 119.200 93.075 119.260 ;
        RECT 96.860 119.400 97.150 119.445 ;
        RECT 98.750 119.400 99.040 119.445 ;
        RECT 101.870 119.400 102.160 119.445 ;
        RECT 96.860 119.260 102.160 119.400 ;
        RECT 96.860 119.215 97.150 119.260 ;
        RECT 98.750 119.215 99.040 119.260 ;
        RECT 101.870 119.215 102.160 119.260 ;
        RECT 90.545 118.920 92.065 119.060 ;
        RECT 90.545 118.765 90.685 118.920 ;
        RECT 90.010 118.535 90.300 118.765 ;
        RECT 90.470 118.535 90.760 118.765 ;
        RECT 91.390 118.535 91.680 118.765 ;
        RECT 91.925 118.720 92.065 118.920 ;
        RECT 92.295 118.860 92.615 119.120 ;
        RECT 94.135 119.060 94.455 119.120 ;
        RECT 95.990 119.060 96.280 119.105 ;
        RECT 100.115 119.060 100.435 119.120 ;
        RECT 94.135 118.920 100.435 119.060 ;
        RECT 94.135 118.860 94.455 118.920 ;
        RECT 95.990 118.875 96.280 118.920 ;
        RECT 100.115 118.860 100.435 118.920 ;
        RECT 93.675 118.720 93.995 118.780 ;
        RECT 91.925 118.580 93.995 118.720 ;
        RECT 89.625 118.380 89.765 118.520 ;
        RECT 76.670 118.240 85.165 118.380 ;
        RECT 87.325 118.240 89.765 118.380 ;
        RECT 91.465 118.380 91.605 118.535 ;
        RECT 93.675 118.520 93.995 118.580 ;
        RECT 96.455 118.720 96.745 118.765 ;
        RECT 98.290 118.720 98.580 118.765 ;
        RECT 101.870 118.720 102.160 118.765 ;
        RECT 96.455 118.580 102.160 118.720 ;
        RECT 96.455 118.535 96.745 118.580 ;
        RECT 98.290 118.535 98.580 118.580 ;
        RECT 101.870 118.535 102.160 118.580 ;
        RECT 91.835 118.380 92.155 118.440 ;
        RECT 91.465 118.240 92.155 118.380 ;
        RECT 76.670 118.195 76.960 118.240 ;
        RECT 83.555 118.180 83.875 118.240 ;
        RECT 43.535 118.040 43.855 118.100 ;
        RECT 40.405 117.900 43.855 118.040 ;
        RECT 35.270 117.855 35.560 117.900 ;
        RECT 35.715 117.840 36.035 117.900 ;
        RECT 43.535 117.840 43.855 117.900 ;
        RECT 45.375 118.040 45.695 118.100 ;
        RECT 47.690 118.040 47.980 118.085 ;
        RECT 45.375 117.900 47.980 118.040 ;
        RECT 45.375 117.840 45.695 117.900 ;
        RECT 47.690 117.855 47.980 117.900 ;
        RECT 57.810 118.040 58.100 118.085 ;
        RECT 58.255 118.040 58.575 118.100 ;
        RECT 57.810 117.900 58.575 118.040 ;
        RECT 57.810 117.855 58.100 117.900 ;
        RECT 58.255 117.840 58.575 117.900 ;
        RECT 63.330 118.040 63.620 118.085 ;
        RECT 68.835 118.040 69.155 118.100 ;
        RECT 63.330 117.900 69.155 118.040 ;
        RECT 63.330 117.855 63.620 117.900 ;
        RECT 68.835 117.840 69.155 117.900 ;
        RECT 72.515 118.040 72.835 118.100 ;
        RECT 74.830 118.040 75.120 118.085 ;
        RECT 72.515 117.900 75.120 118.040 ;
        RECT 72.515 117.840 72.835 117.900 ;
        RECT 74.830 117.855 75.120 117.900 ;
        RECT 78.970 118.040 79.260 118.085 ;
        RECT 79.415 118.040 79.735 118.100 ;
        RECT 78.970 117.900 79.735 118.040 ;
        RECT 78.970 117.855 79.260 117.900 ;
        RECT 79.415 117.840 79.735 117.900 ;
        RECT 80.795 118.040 81.115 118.100 ;
        RECT 82.650 118.040 82.940 118.085 ;
        RECT 80.795 117.900 82.940 118.040 ;
        RECT 80.795 117.840 81.115 117.900 ;
        RECT 82.650 117.855 82.940 117.900 ;
        RECT 84.015 118.040 84.335 118.100 ;
        RECT 87.325 118.040 87.465 118.240 ;
        RECT 91.835 118.180 92.155 118.240 ;
        RECT 93.230 118.380 93.520 118.425 ;
        RECT 95.975 118.380 96.295 118.440 ;
        RECT 102.950 118.425 103.240 118.740 ;
        RECT 93.230 118.240 96.295 118.380 ;
        RECT 93.230 118.195 93.520 118.240 ;
        RECT 95.975 118.180 96.295 118.240 ;
        RECT 97.370 118.195 97.660 118.425 ;
        RECT 99.650 118.380 100.300 118.425 ;
        RECT 102.950 118.380 103.540 118.425 ;
        RECT 104.715 118.380 105.035 118.440 ;
        RECT 99.650 118.240 105.035 118.380 ;
        RECT 99.650 118.195 100.300 118.240 ;
        RECT 103.250 118.195 103.540 118.240 ;
        RECT 84.015 117.900 87.465 118.040 ;
        RECT 88.615 118.040 88.935 118.100 ;
        RECT 93.690 118.040 93.980 118.085 ;
        RECT 88.615 117.900 93.980 118.040 ;
        RECT 84.015 117.840 84.335 117.900 ;
        RECT 88.615 117.840 88.935 117.900 ;
        RECT 93.690 117.855 93.980 117.900 ;
        RECT 95.530 118.040 95.820 118.085 ;
        RECT 97.445 118.040 97.585 118.195 ;
        RECT 104.715 118.180 105.035 118.240 ;
        RECT 95.530 117.900 97.585 118.040 ;
        RECT 95.530 117.855 95.820 117.900 ;
        RECT 18.165 117.220 112.465 117.700 ;
        RECT 39.410 117.020 39.700 117.065 ;
        RECT 42.615 117.020 42.935 117.080 ;
        RECT 39.410 116.880 42.935 117.020 ;
        RECT 39.410 116.835 39.700 116.880 ;
        RECT 42.615 116.820 42.935 116.880 ;
        RECT 43.535 116.820 43.855 117.080 ;
        RECT 43.995 117.020 44.315 117.080 ;
        RECT 43.995 116.880 51.585 117.020 ;
        RECT 43.995 116.820 44.315 116.880 ;
        RECT 25.710 116.680 26.000 116.725 ;
        RECT 26.515 116.680 26.835 116.740 ;
        RECT 28.950 116.680 29.600 116.725 ;
        RECT 25.710 116.540 29.600 116.680 ;
        RECT 25.710 116.495 26.300 116.540 ;
        RECT 26.010 116.180 26.300 116.495 ;
        RECT 26.515 116.480 26.835 116.540 ;
        RECT 28.950 116.495 29.600 116.540 ;
        RECT 35.255 116.480 35.575 116.740 ;
        RECT 38.935 116.680 39.255 116.740 ;
        RECT 36.265 116.540 39.255 116.680 ;
        RECT 27.090 116.340 27.380 116.385 ;
        RECT 30.670 116.340 30.960 116.385 ;
        RECT 32.505 116.340 32.795 116.385 ;
        RECT 27.090 116.200 32.795 116.340 ;
        RECT 27.090 116.155 27.380 116.200 ;
        RECT 30.670 116.155 30.960 116.200 ;
        RECT 32.505 116.155 32.795 116.200 ;
        RECT 32.955 116.340 33.275 116.400 ;
        RECT 36.265 116.340 36.405 116.540 ;
        RECT 38.935 116.480 39.255 116.540 ;
        RECT 43.090 116.680 43.380 116.725 ;
        RECT 50.895 116.680 51.215 116.740 ;
        RECT 43.090 116.540 51.215 116.680 ;
        RECT 43.090 116.495 43.380 116.540 ;
        RECT 50.895 116.480 51.215 116.540 ;
        RECT 32.955 116.200 36.405 116.340 ;
        RECT 32.955 116.140 33.275 116.200 ;
        RECT 36.635 116.140 36.955 116.400 ;
        RECT 38.475 116.340 38.795 116.400 ;
        RECT 41.235 116.340 41.555 116.400 ;
        RECT 38.475 116.200 46.065 116.340 ;
        RECT 38.475 116.140 38.795 116.200 ;
        RECT 41.235 116.140 41.555 116.200 ;
        RECT 22.835 115.800 23.155 116.060 ;
        RECT 31.590 116.000 31.880 116.045 ;
        RECT 34.795 116.000 35.115 116.060 ;
        RECT 31.590 115.860 35.115 116.000 ;
        RECT 31.590 115.815 31.880 115.860 ;
        RECT 34.795 115.800 35.115 115.860 ;
        RECT 39.395 116.000 39.715 116.060 ;
        RECT 39.870 116.000 40.160 116.045 ;
        RECT 45.375 116.000 45.695 116.060 ;
        RECT 39.395 115.860 45.695 116.000 ;
        RECT 45.925 116.000 46.065 116.200 ;
        RECT 46.755 116.140 47.075 116.400 ;
        RECT 49.515 116.340 49.835 116.400 ;
        RECT 47.305 116.200 49.835 116.340 ;
        RECT 47.305 116.000 47.445 116.200 ;
        RECT 49.515 116.140 49.835 116.200 ;
        RECT 49.990 116.155 50.280 116.385 ;
        RECT 50.065 116.000 50.205 116.155 ;
        RECT 50.435 116.140 50.755 116.400 ;
        RECT 51.445 116.385 51.585 116.880 ;
        RECT 52.275 116.820 52.595 117.080 ;
        RECT 70.215 117.020 70.535 117.080 ;
        RECT 56.505 116.880 70.535 117.020 ;
        RECT 51.370 116.155 51.660 116.385 ;
        RECT 52.735 116.140 53.055 116.400 ;
        RECT 56.505 116.000 56.645 116.880 ;
        RECT 63.775 116.725 64.095 116.740 ;
        RECT 57.815 116.680 58.105 116.725 ;
        RECT 59.675 116.680 59.965 116.725 ;
        RECT 57.815 116.540 59.965 116.680 ;
        RECT 57.815 116.495 58.105 116.540 ;
        RECT 59.675 116.495 59.965 116.540 ;
        RECT 60.595 116.680 60.885 116.725 ;
        RECT 63.775 116.680 64.145 116.725 ;
        RECT 60.595 116.540 64.145 116.680 ;
        RECT 60.595 116.495 60.885 116.540 ;
        RECT 63.775 116.495 64.145 116.540 ;
        RECT 64.695 116.680 65.015 116.740 ;
        RECT 67.010 116.680 67.300 116.725 ;
        RECT 64.695 116.540 67.300 116.680 ;
        RECT 58.715 116.140 59.035 116.400 ;
        RECT 59.750 116.340 59.965 116.495 ;
        RECT 63.775 116.480 64.095 116.495 ;
        RECT 64.695 116.480 65.015 116.540 ;
        RECT 67.010 116.495 67.300 116.540 ;
        RECT 68.925 116.385 69.065 116.880 ;
        RECT 70.215 116.820 70.535 116.880 ;
        RECT 71.135 116.820 71.455 117.080 ;
        RECT 86.315 117.020 86.635 117.080 ;
        RECT 72.145 116.880 86.635 117.020 ;
        RECT 72.145 116.680 72.285 116.880 ;
        RECT 86.315 116.820 86.635 116.880 ;
        RECT 88.170 117.020 88.460 117.065 ;
        RECT 88.615 117.020 88.935 117.080 ;
        RECT 88.170 116.880 88.935 117.020 ;
        RECT 88.170 116.835 88.460 116.880 ;
        RECT 88.615 116.820 88.935 116.880 ;
        RECT 90.455 117.020 90.775 117.080 ;
        RECT 92.310 117.020 92.600 117.065 ;
        RECT 90.455 116.880 92.600 117.020 ;
        RECT 90.455 116.820 90.775 116.880 ;
        RECT 92.310 116.835 92.600 116.880 ;
        RECT 95.975 116.820 96.295 117.080 ;
        RECT 97.815 116.820 98.135 117.080 ;
        RECT 98.750 117.020 99.040 117.065 ;
        RECT 99.195 117.020 99.515 117.080 ;
        RECT 98.750 116.880 99.515 117.020 ;
        RECT 98.750 116.835 99.040 116.880 ;
        RECT 99.195 116.820 99.515 116.880 ;
        RECT 104.715 116.820 105.035 117.080 ;
        RECT 70.305 116.540 72.285 116.680 ;
        RECT 72.530 116.680 72.820 116.725 ;
        RECT 78.490 116.680 79.140 116.725 ;
        RECT 82.090 116.680 82.380 116.725 ;
        RECT 84.015 116.680 84.335 116.740 ;
        RECT 72.530 116.540 82.380 116.680 ;
        RECT 70.305 116.400 70.445 116.540 ;
        RECT 72.530 116.495 72.820 116.540 ;
        RECT 78.490 116.495 79.140 116.540 ;
        RECT 81.790 116.495 82.380 116.540 ;
        RECT 83.185 116.540 84.335 116.680 ;
        RECT 61.995 116.340 62.285 116.385 ;
        RECT 59.750 116.200 62.285 116.340 ;
        RECT 61.995 116.155 62.285 116.200 ;
        RECT 68.390 116.155 68.680 116.385 ;
        RECT 68.850 116.155 69.140 116.385 ;
        RECT 69.310 116.155 69.600 116.385 ;
        RECT 45.925 115.860 47.445 116.000 ;
        RECT 49.605 115.860 56.645 116.000 ;
        RECT 56.875 116.000 57.195 116.060 ;
        RECT 59.635 116.000 59.955 116.060 ;
        RECT 56.875 115.860 59.955 116.000 ;
        RECT 39.395 115.800 39.715 115.860 ;
        RECT 39.870 115.815 40.160 115.860 ;
        RECT 45.375 115.800 45.695 115.860 ;
        RECT 27.090 115.660 27.380 115.705 ;
        RECT 30.210 115.660 30.500 115.705 ;
        RECT 32.100 115.660 32.390 115.705 ;
        RECT 27.090 115.520 32.390 115.660 ;
        RECT 27.090 115.475 27.380 115.520 ;
        RECT 30.210 115.475 30.500 115.520 ;
        RECT 32.100 115.475 32.390 115.520 ;
        RECT 34.350 115.660 34.640 115.705 ;
        RECT 38.935 115.660 39.255 115.720 ;
        RECT 41.695 115.660 42.015 115.720 ;
        RECT 49.605 115.660 49.745 115.860 ;
        RECT 56.875 115.800 57.195 115.860 ;
        RECT 59.635 115.800 59.955 115.860 ;
        RECT 60.095 116.000 60.415 116.060 ;
        RECT 68.465 116.000 68.605 116.155 ;
        RECT 69.385 116.000 69.525 116.155 ;
        RECT 70.215 116.140 70.535 116.400 ;
        RECT 70.690 116.340 70.980 116.385 ;
        RECT 71.595 116.340 71.915 116.400 ;
        RECT 70.690 116.200 71.915 116.340 ;
        RECT 70.690 116.155 70.980 116.200 ;
        RECT 71.595 116.140 71.915 116.200 ;
        RECT 72.070 116.340 72.360 116.385 ;
        RECT 73.895 116.340 74.215 116.400 ;
        RECT 72.070 116.200 74.215 116.340 ;
        RECT 72.070 116.155 72.360 116.200 ;
        RECT 73.895 116.140 74.215 116.200 ;
        RECT 75.295 116.340 75.585 116.385 ;
        RECT 77.130 116.340 77.420 116.385 ;
        RECT 80.710 116.340 81.000 116.385 ;
        RECT 75.295 116.200 81.000 116.340 ;
        RECT 75.295 116.155 75.585 116.200 ;
        RECT 77.130 116.155 77.420 116.200 ;
        RECT 80.710 116.155 81.000 116.200 ;
        RECT 81.790 116.180 82.080 116.495 ;
        RECT 72.515 116.000 72.835 116.060 ;
        RECT 60.095 115.860 69.065 116.000 ;
        RECT 69.385 115.860 72.835 116.000 ;
        RECT 60.095 115.800 60.415 115.860 ;
        RECT 34.350 115.520 49.745 115.660 ;
        RECT 57.355 115.660 57.645 115.705 ;
        RECT 59.215 115.660 59.505 115.705 ;
        RECT 61.995 115.660 62.285 115.705 ;
        RECT 57.355 115.520 62.285 115.660 ;
        RECT 68.925 115.660 69.065 115.860 ;
        RECT 72.515 115.800 72.835 115.860 ;
        RECT 74.815 115.800 75.135 116.060 ;
        RECT 83.185 116.000 83.325 116.540 ;
        RECT 84.015 116.480 84.335 116.540 ;
        RECT 89.995 116.480 90.315 116.740 ;
        RECT 91.835 116.680 92.155 116.740 ;
        RECT 96.450 116.680 96.740 116.725 ;
        RECT 97.905 116.680 98.045 116.820 ;
        RECT 91.835 116.540 94.365 116.680 ;
        RECT 91.835 116.480 92.155 116.540 ;
        RECT 90.915 116.340 91.235 116.400 ;
        RECT 91.390 116.340 91.680 116.385 ;
        RECT 90.915 116.200 91.680 116.340 ;
        RECT 90.915 116.140 91.235 116.200 ;
        RECT 91.390 116.155 91.680 116.200 ;
        RECT 93.230 116.340 93.520 116.385 ;
        RECT 93.675 116.340 93.995 116.400 ;
        RECT 93.230 116.200 93.995 116.340 ;
        RECT 94.225 116.340 94.365 116.540 ;
        RECT 96.450 116.540 98.045 116.680 ;
        RECT 100.665 116.540 103.105 116.680 ;
        RECT 96.450 116.495 96.740 116.540 ;
        RECT 97.830 116.340 98.120 116.385 ;
        RECT 94.225 116.200 98.120 116.340 ;
        RECT 93.230 116.155 93.520 116.200 ;
        RECT 93.675 116.140 93.995 116.200 ;
        RECT 97.830 116.155 98.120 116.200 ;
        RECT 98.735 116.340 99.055 116.400 ;
        RECT 100.665 116.385 100.805 116.540 ;
        RECT 100.590 116.340 100.880 116.385 ;
        RECT 98.735 116.200 100.880 116.340 ;
        RECT 98.735 116.140 99.055 116.200 ;
        RECT 100.590 116.155 100.880 116.200 ;
        RECT 101.035 116.140 101.355 116.400 ;
        RECT 102.965 116.385 103.105 116.540 ;
        RECT 102.890 116.155 103.180 116.385 ;
        RECT 105.175 116.140 105.495 116.400 ;
        RECT 75.365 115.860 83.325 116.000 ;
        RECT 83.555 116.000 83.875 116.060 ;
        RECT 84.950 116.000 85.240 116.045 ;
        RECT 83.555 115.860 85.240 116.000 ;
        RECT 75.365 115.660 75.505 115.860 ;
        RECT 83.555 115.800 83.875 115.860 ;
        RECT 84.950 115.815 85.240 115.860 ;
        RECT 90.455 115.800 90.775 116.060 ;
        RECT 94.595 116.000 94.915 116.060 ;
        RECT 96.910 116.000 97.200 116.045 ;
        RECT 94.595 115.860 97.200 116.000 ;
        RECT 94.595 115.800 94.915 115.860 ;
        RECT 96.910 115.815 97.200 115.860 ;
        RECT 98.275 116.000 98.595 116.060 ;
        RECT 103.810 116.000 104.100 116.045 ;
        RECT 98.275 115.860 104.100 116.000 ;
        RECT 98.275 115.800 98.595 115.860 ;
        RECT 103.810 115.815 104.100 115.860 ;
        RECT 68.925 115.520 75.505 115.660 ;
        RECT 75.700 115.660 75.990 115.705 ;
        RECT 77.590 115.660 77.880 115.705 ;
        RECT 80.710 115.660 81.000 115.705 ;
        RECT 75.700 115.520 81.000 115.660 ;
        RECT 34.350 115.475 34.640 115.520 ;
        RECT 38.935 115.460 39.255 115.520 ;
        RECT 41.695 115.460 42.015 115.520 ;
        RECT 57.355 115.475 57.645 115.520 ;
        RECT 59.215 115.475 59.505 115.520 ;
        RECT 61.995 115.475 62.285 115.520 ;
        RECT 75.700 115.475 75.990 115.520 ;
        RECT 77.590 115.475 77.880 115.520 ;
        RECT 80.710 115.475 81.000 115.520 ;
        RECT 91.835 115.660 92.155 115.720 ;
        RECT 99.670 115.660 99.960 115.705 ;
        RECT 91.835 115.520 99.960 115.660 ;
        RECT 91.835 115.460 92.155 115.520 ;
        RECT 99.670 115.475 99.960 115.520 ;
        RECT 36.635 115.320 36.955 115.380 ;
        RECT 48.150 115.320 48.440 115.365 ;
        RECT 36.635 115.180 48.440 115.320 ;
        RECT 36.635 115.120 36.955 115.180 ;
        RECT 48.150 115.135 48.440 115.180 ;
        RECT 49.515 115.320 49.835 115.380 ;
        RECT 60.095 115.320 60.415 115.380 ;
        RECT 49.515 115.180 60.415 115.320 ;
        RECT 49.515 115.120 49.835 115.180 ;
        RECT 60.095 115.120 60.415 115.180 ;
        RECT 60.555 115.320 60.875 115.380 ;
        RECT 65.860 115.320 66.150 115.365 ;
        RECT 66.535 115.320 66.855 115.380 ;
        RECT 76.195 115.365 76.515 115.380 ;
        RECT 60.555 115.180 66.855 115.320 ;
        RECT 60.555 115.120 60.875 115.180 ;
        RECT 65.860 115.135 66.150 115.180 ;
        RECT 66.535 115.120 66.855 115.180 ;
        RECT 76.150 115.135 76.515 115.365 ;
        RECT 76.195 115.120 76.515 115.135 ;
        RECT 84.015 115.320 84.335 115.380 ;
        RECT 90.010 115.320 90.300 115.365 ;
        RECT 84.015 115.180 90.300 115.320 ;
        RECT 84.015 115.120 84.335 115.180 ;
        RECT 90.010 115.135 90.300 115.180 ;
        RECT 97.830 115.320 98.120 115.365 ;
        RECT 101.970 115.320 102.260 115.365 ;
        RECT 97.830 115.180 102.260 115.320 ;
        RECT 97.830 115.135 98.120 115.180 ;
        RECT 101.970 115.135 102.260 115.180 ;
        RECT 17.605 114.500 112.465 114.980 ;
        RECT 26.515 114.100 26.835 114.360 ;
        RECT 32.970 114.115 33.260 114.345 ;
        RECT 35.255 114.300 35.575 114.360 ;
        RECT 61.935 114.300 62.255 114.360 ;
        RECT 35.255 114.160 62.255 114.300 ;
        RECT 31.590 113.960 31.880 114.005 ;
        RECT 33.045 113.960 33.185 114.115 ;
        RECT 35.255 114.100 35.575 114.160 ;
        RECT 61.935 114.100 62.255 114.160 ;
        RECT 62.410 114.300 62.700 114.345 ;
        RECT 70.215 114.300 70.535 114.360 ;
        RECT 62.410 114.160 70.535 114.300 ;
        RECT 62.410 114.115 62.700 114.160 ;
        RECT 70.215 114.100 70.535 114.160 ;
        RECT 75.735 114.100 76.055 114.360 ;
        RECT 76.195 114.100 76.515 114.360 ;
        RECT 79.890 114.115 80.180 114.345 ;
        RECT 85.870 114.300 86.160 114.345 ;
        RECT 91.835 114.300 92.155 114.360 ;
        RECT 85.870 114.160 92.155 114.300 ;
        RECT 85.870 114.115 86.160 114.160 ;
        RECT 40.315 113.960 40.635 114.020 ;
        RECT 31.590 113.820 33.185 113.960 ;
        RECT 33.965 113.820 40.635 113.960 ;
        RECT 31.590 113.775 31.880 113.820 ;
        RECT 33.965 113.665 34.105 113.820 ;
        RECT 40.315 113.760 40.635 113.820 ;
        RECT 72.070 113.960 72.360 114.005 ;
        RECT 79.965 113.960 80.105 114.115 ;
        RECT 91.835 114.100 92.155 114.160 ;
        RECT 72.070 113.820 80.105 113.960 ;
        RECT 72.070 113.775 72.360 113.820 ;
        RECT 83.570 113.775 83.860 114.005 ;
        RECT 96.405 113.960 96.695 114.005 ;
        RECT 99.185 113.960 99.475 114.005 ;
        RECT 101.045 113.960 101.335 114.005 ;
        RECT 96.405 113.820 101.335 113.960 ;
        RECT 96.405 113.775 96.695 113.820 ;
        RECT 99.185 113.775 99.475 113.820 ;
        RECT 101.045 113.775 101.335 113.820 ;
        RECT 29.825 113.480 30.885 113.620 ;
        RECT 24.215 113.280 24.535 113.340 ;
        RECT 26.070 113.280 26.360 113.325 ;
        RECT 24.215 113.140 26.360 113.280 ;
        RECT 24.215 113.080 24.535 113.140 ;
        RECT 26.070 113.095 26.360 113.140 ;
        RECT 27.895 113.080 28.215 113.340 ;
        RECT 28.370 113.280 28.660 113.325 ;
        RECT 29.825 113.280 29.965 113.480 ;
        RECT 28.370 113.140 29.965 113.280 ;
        RECT 28.370 113.095 28.660 113.140 ;
        RECT 30.195 113.080 30.515 113.340 ;
        RECT 30.745 113.325 30.885 113.480 ;
        RECT 32.125 113.480 33.645 113.620 ;
        RECT 30.670 113.280 30.960 113.325 ;
        RECT 32.125 113.280 32.265 113.480 ;
        RECT 30.670 113.140 32.265 113.280 ;
        RECT 32.495 113.280 32.815 113.340 ;
        RECT 32.970 113.280 33.260 113.325 ;
        RECT 32.495 113.140 33.260 113.280 ;
        RECT 33.505 113.280 33.645 113.480 ;
        RECT 33.890 113.435 34.180 113.665 ;
        RECT 41.235 113.620 41.555 113.680 ;
        RECT 55.495 113.620 55.815 113.680 ;
        RECT 56.890 113.620 57.180 113.665 ;
        RECT 34.885 113.480 36.405 113.620 ;
        RECT 34.885 113.290 35.025 113.480 ;
        RECT 33.965 113.280 35.025 113.290 ;
        RECT 33.505 113.150 35.025 113.280 ;
        RECT 35.255 113.280 35.575 113.340 ;
        RECT 35.730 113.280 36.020 113.325 ;
        RECT 33.505 113.140 34.105 113.150 ;
        RECT 35.255 113.140 36.020 113.280 ;
        RECT 36.265 113.280 36.405 113.480 ;
        RECT 38.105 113.480 41.005 113.620 ;
        RECT 36.650 113.280 36.940 113.325 ;
        RECT 37.555 113.280 37.875 113.340 ;
        RECT 36.265 113.140 37.875 113.280 ;
        RECT 30.670 113.095 30.960 113.140 ;
        RECT 32.495 113.080 32.815 113.140 ;
        RECT 32.970 113.095 33.260 113.140 ;
        RECT 35.255 113.080 35.575 113.140 ;
        RECT 35.730 113.095 36.020 113.140 ;
        RECT 36.650 113.095 36.940 113.140 ;
        RECT 37.555 113.080 37.875 113.140 ;
        RECT 29.290 112.940 29.580 112.985 ;
        RECT 34.350 112.940 34.640 112.985 ;
        RECT 38.105 112.940 38.245 113.480 ;
        RECT 38.475 113.080 38.795 113.340 ;
        RECT 38.935 113.080 39.255 113.340 ;
        RECT 39.395 113.080 39.715 113.340 ;
        RECT 40.330 113.095 40.620 113.325 ;
        RECT 40.865 113.280 41.005 113.480 ;
        RECT 41.235 113.480 47.445 113.620 ;
        RECT 41.235 113.420 41.555 113.480 ;
        RECT 41.695 113.280 42.015 113.340 ;
        RECT 40.865 113.140 42.015 113.280 ;
        RECT 40.405 112.940 40.545 113.095 ;
        RECT 41.695 113.080 42.015 113.140 ;
        RECT 46.310 113.095 46.600 113.325 ;
        RECT 29.290 112.800 33.185 112.940 ;
        RECT 29.290 112.755 29.580 112.800 ;
        RECT 33.045 112.660 33.185 112.800 ;
        RECT 34.350 112.800 38.245 112.940 ;
        RECT 39.485 112.800 40.545 112.940 ;
        RECT 34.350 112.755 34.640 112.800 ;
        RECT 31.115 112.600 31.435 112.660 ;
        RECT 32.050 112.600 32.340 112.645 ;
        RECT 31.115 112.460 32.340 112.600 ;
        RECT 31.115 112.400 31.435 112.460 ;
        RECT 32.050 112.415 32.340 112.460 ;
        RECT 32.955 112.400 33.275 112.660 ;
        RECT 33.415 112.600 33.735 112.660 ;
        RECT 37.110 112.600 37.400 112.645 ;
        RECT 33.415 112.460 37.400 112.600 ;
        RECT 33.415 112.400 33.735 112.460 ;
        RECT 37.110 112.415 37.400 112.460 ;
        RECT 38.015 112.600 38.335 112.660 ;
        RECT 39.485 112.600 39.625 112.800 ;
        RECT 45.375 112.740 45.695 113.000 ;
        RECT 46.385 112.940 46.525 113.095 ;
        RECT 46.755 113.080 47.075 113.340 ;
        RECT 47.305 113.280 47.445 113.480 ;
        RECT 53.055 113.480 57.180 113.620 ;
        RECT 53.055 113.280 53.195 113.480 ;
        RECT 55.495 113.420 55.815 113.480 ;
        RECT 56.890 113.435 57.180 113.480 ;
        RECT 61.565 113.480 71.365 113.620 ;
        RECT 47.305 113.140 53.195 113.280 ;
        RECT 55.050 113.095 55.340 113.325 ;
        RECT 55.955 113.280 56.275 113.340 ;
        RECT 61.565 113.280 61.705 113.480 ;
        RECT 55.955 113.140 61.705 113.280 ;
        RECT 61.950 113.280 62.240 113.325 ;
        RECT 63.315 113.280 63.635 113.340 ;
        RECT 61.950 113.140 63.635 113.280 ;
        RECT 50.895 112.940 51.215 113.000 ;
        RECT 46.385 112.800 51.215 112.940 ;
        RECT 50.895 112.740 51.215 112.800 ;
        RECT 51.355 112.940 51.675 113.000 ;
        RECT 55.125 112.940 55.265 113.095 ;
        RECT 55.955 113.080 56.275 113.140 ;
        RECT 61.950 113.095 62.240 113.140 ;
        RECT 63.315 113.080 63.635 113.140 ;
        RECT 65.615 113.280 65.935 113.340 ;
        RECT 68.465 113.325 68.605 113.480 ;
        RECT 71.225 113.340 71.365 113.480 ;
        RECT 72.515 113.420 72.835 113.680 ;
        RECT 79.415 113.420 79.735 113.680 ;
        RECT 80.795 113.420 81.115 113.680 ;
        RECT 83.645 113.340 83.785 113.775 ;
        RECT 85.410 113.620 85.700 113.665 ;
        RECT 87.235 113.620 87.555 113.680 ;
        RECT 85.410 113.480 87.555 113.620 ;
        RECT 85.410 113.435 85.700 113.480 ;
        RECT 87.235 113.420 87.555 113.480 ;
        RECT 88.155 113.620 88.475 113.680 ;
        RECT 88.630 113.620 88.920 113.665 ;
        RECT 93.675 113.620 93.995 113.680 ;
        RECT 88.155 113.480 93.995 113.620 ;
        RECT 88.155 113.420 88.475 113.480 ;
        RECT 88.630 113.435 88.920 113.480 ;
        RECT 93.675 113.420 93.995 113.480 ;
        RECT 99.655 113.420 99.975 113.680 ;
        RECT 100.115 113.620 100.435 113.680 ;
        RECT 101.510 113.620 101.800 113.665 ;
        RECT 100.115 113.480 101.800 113.620 ;
        RECT 100.115 113.420 100.435 113.480 ;
        RECT 101.510 113.435 101.800 113.480 ;
        RECT 67.470 113.280 67.760 113.325 ;
        RECT 65.615 113.140 67.760 113.280 ;
        RECT 65.615 113.080 65.935 113.140 ;
        RECT 67.470 113.095 67.760 113.140 ;
        RECT 68.390 113.095 68.680 113.325 ;
        RECT 68.850 113.095 69.140 113.325 ;
        RECT 70.690 113.095 70.980 113.325 ;
        RECT 51.355 112.800 55.265 112.940 ;
        RECT 57.810 112.940 58.100 112.985 ;
        RECT 62.855 112.940 63.175 113.000 ;
        RECT 64.235 112.940 64.555 113.000 ;
        RECT 57.810 112.800 64.555 112.940 ;
        RECT 51.355 112.740 51.675 112.800 ;
        RECT 57.810 112.755 58.100 112.800 ;
        RECT 62.855 112.740 63.175 112.800 ;
        RECT 64.235 112.740 64.555 112.800 ;
        RECT 66.535 112.940 66.855 113.000 ;
        RECT 68.925 112.940 69.065 113.095 ;
        RECT 66.535 112.800 69.065 112.940 ;
        RECT 70.765 112.940 70.905 113.095 ;
        RECT 71.135 113.080 71.455 113.340 ;
        RECT 71.595 113.280 71.915 113.340 ;
        RECT 73.435 113.280 73.755 113.340 ;
        RECT 79.890 113.280 80.180 113.325 ;
        RECT 80.335 113.280 80.655 113.340 ;
        RECT 71.595 113.140 76.425 113.280 ;
        RECT 71.595 113.080 71.915 113.140 ;
        RECT 73.435 113.080 73.755 113.140 ;
        RECT 75.735 112.940 76.055 113.000 ;
        RECT 70.765 112.800 76.055 112.940 ;
        RECT 76.285 112.940 76.425 113.140 ;
        RECT 79.890 113.140 80.655 113.280 ;
        RECT 79.890 113.095 80.180 113.140 ;
        RECT 80.335 113.080 80.655 113.140 ;
        RECT 81.255 113.080 81.575 113.340 ;
        RECT 83.555 113.080 83.875 113.340 ;
        RECT 84.475 113.080 84.795 113.340 ;
        RECT 85.855 113.080 86.175 113.340 ;
        RECT 87.710 113.280 88.000 113.325 ;
        RECT 89.075 113.280 89.395 113.340 ;
        RECT 87.710 113.140 89.395 113.280 ;
        RECT 87.710 113.095 88.000 113.140 ;
        RECT 80.795 112.940 81.115 113.000 ;
        RECT 87.785 112.940 87.925 113.095 ;
        RECT 89.075 113.080 89.395 113.140 ;
        RECT 90.010 113.280 90.300 113.325 ;
        RECT 95.055 113.280 95.375 113.340 ;
        RECT 90.010 113.140 95.375 113.280 ;
        RECT 90.010 113.095 90.300 113.140 ;
        RECT 95.055 113.080 95.375 113.140 ;
        RECT 96.405 113.280 96.695 113.325 ;
        RECT 96.405 113.140 98.940 113.280 ;
        RECT 96.405 113.095 96.695 113.140 ;
        RECT 97.815 112.985 98.135 113.000 ;
        RECT 76.285 112.800 87.925 112.940 ;
        RECT 89.550 112.940 89.840 112.985 ;
        RECT 92.540 112.940 92.830 112.985 ;
        RECT 94.545 112.940 94.835 112.985 ;
        RECT 97.805 112.940 98.135 112.985 ;
        RECT 89.550 112.800 94.365 112.940 ;
        RECT 66.535 112.740 66.855 112.800 ;
        RECT 75.735 112.740 76.055 112.800 ;
        RECT 80.795 112.740 81.115 112.800 ;
        RECT 89.550 112.755 89.840 112.800 ;
        RECT 92.540 112.755 92.830 112.800 ;
        RECT 38.015 112.460 39.625 112.600 ;
        RECT 39.855 112.600 40.175 112.660 ;
        RECT 41.695 112.600 42.015 112.660 ;
        RECT 39.855 112.460 42.015 112.600 ;
        RECT 38.015 112.400 38.335 112.460 ;
        RECT 39.855 112.400 40.175 112.460 ;
        RECT 41.695 112.400 42.015 112.460 ;
        RECT 42.155 112.400 42.475 112.660 ;
        RECT 42.615 112.400 42.935 112.660 ;
        RECT 44.455 112.400 44.775 112.660 ;
        RECT 55.510 112.600 55.800 112.645 ;
        RECT 55.955 112.600 56.275 112.660 ;
        RECT 55.510 112.460 56.275 112.600 ;
        RECT 55.510 112.415 55.800 112.460 ;
        RECT 55.955 112.400 56.275 112.460 ;
        RECT 56.415 112.600 56.735 112.660 ;
        RECT 58.270 112.600 58.560 112.645 ;
        RECT 56.415 112.460 58.560 112.600 ;
        RECT 56.415 112.400 56.735 112.460 ;
        RECT 58.270 112.415 58.560 112.460 ;
        RECT 60.110 112.600 60.400 112.645 ;
        RECT 61.015 112.600 61.335 112.660 ;
        RECT 60.110 112.460 61.335 112.600 ;
        RECT 60.110 112.415 60.400 112.460 ;
        RECT 61.015 112.400 61.335 112.460 ;
        RECT 68.375 112.600 68.695 112.660 ;
        RECT 71.595 112.600 71.915 112.660 ;
        RECT 68.375 112.460 71.915 112.600 ;
        RECT 68.375 112.400 68.695 112.460 ;
        RECT 71.595 112.400 71.915 112.460 ;
        RECT 82.190 112.600 82.480 112.645 ;
        RECT 84.475 112.600 84.795 112.660 ;
        RECT 82.190 112.460 84.795 112.600 ;
        RECT 82.190 112.415 82.480 112.460 ;
        RECT 84.475 112.400 84.795 112.460 ;
        RECT 86.315 112.600 86.635 112.660 ;
        RECT 87.250 112.600 87.540 112.645 ;
        RECT 86.315 112.460 87.540 112.600 ;
        RECT 86.315 112.400 86.635 112.460 ;
        RECT 87.250 112.415 87.540 112.460 ;
        RECT 91.375 112.600 91.695 112.660 ;
        RECT 91.850 112.600 92.140 112.645 ;
        RECT 91.375 112.460 92.140 112.600 ;
        RECT 94.225 112.600 94.365 112.800 ;
        RECT 94.545 112.800 98.135 112.940 ;
        RECT 94.545 112.755 94.835 112.800 ;
        RECT 97.805 112.755 98.135 112.800 ;
        RECT 98.725 112.985 98.940 113.140 ;
        RECT 98.725 112.940 99.015 112.985 ;
        RECT 100.585 112.940 100.875 112.985 ;
        RECT 98.725 112.800 100.875 112.940 ;
        RECT 98.725 112.755 99.015 112.800 ;
        RECT 100.585 112.755 100.875 112.800 ;
        RECT 97.815 112.740 98.135 112.755 ;
        RECT 96.435 112.600 96.755 112.660 ;
        RECT 94.225 112.460 96.755 112.600 ;
        RECT 91.375 112.400 91.695 112.460 ;
        RECT 91.850 112.415 92.140 112.460 ;
        RECT 96.435 112.400 96.755 112.460 ;
        RECT 18.165 111.780 112.465 112.260 ;
        RECT 32.035 111.380 32.355 111.640 ;
        RECT 34.795 111.380 35.115 111.640 ;
        RECT 40.775 111.580 41.095 111.640 ;
        RECT 39.485 111.440 41.095 111.580 ;
        RECT 29.735 111.240 30.055 111.300 ;
        RECT 29.735 111.100 32.495 111.240 ;
        RECT 29.735 111.040 30.055 111.100 ;
        RECT 24.215 110.900 24.535 110.960 ;
        RECT 30.670 110.900 30.960 110.945 ;
        RECT 24.215 110.760 30.960 110.900 ;
        RECT 32.355 110.900 32.495 111.100 ;
        RECT 34.335 111.040 34.655 111.300 ;
        RECT 36.635 111.240 36.955 111.300 ;
        RECT 36.265 111.100 36.955 111.240 ;
        RECT 32.970 110.900 33.260 110.945 ;
        RECT 32.355 110.760 33.260 110.900 ;
        RECT 24.215 110.700 24.535 110.760 ;
        RECT 30.670 110.715 30.960 110.760 ;
        RECT 32.970 110.715 33.260 110.760 ;
        RECT 33.415 110.700 33.735 110.960 ;
        RECT 35.715 110.700 36.035 110.960 ;
        RECT 36.265 110.945 36.405 111.100 ;
        RECT 36.635 111.040 36.955 111.100 ;
        RECT 37.110 111.240 37.400 111.285 ;
        RECT 39.485 111.240 39.625 111.440 ;
        RECT 40.775 111.380 41.095 111.440 ;
        RECT 41.695 111.580 42.015 111.640 ;
        RECT 45.375 111.580 45.695 111.640 ;
        RECT 41.695 111.440 45.695 111.580 ;
        RECT 41.695 111.380 42.015 111.440 ;
        RECT 45.375 111.380 45.695 111.440 ;
        RECT 46.755 111.580 47.075 111.640 ;
        RECT 53.900 111.580 54.190 111.625 ;
        RECT 56.415 111.580 56.735 111.640 ;
        RECT 46.755 111.440 56.735 111.580 ;
        RECT 46.755 111.380 47.075 111.440 ;
        RECT 53.900 111.395 54.190 111.440 ;
        RECT 56.415 111.380 56.735 111.440 ;
        RECT 63.775 111.380 64.095 111.640 ;
        RECT 64.235 111.580 64.555 111.640 ;
        RECT 71.150 111.580 71.440 111.625 ;
        RECT 81.040 111.580 81.330 111.625 ;
        RECT 92.310 111.580 92.600 111.625 ;
        RECT 64.235 111.440 71.440 111.580 ;
        RECT 64.235 111.380 64.555 111.440 ;
        RECT 71.150 111.395 71.440 111.440 ;
        RECT 79.965 111.440 92.600 111.580 ;
        RECT 39.855 111.285 40.175 111.300 ;
        RECT 55.955 111.285 56.275 111.300 ;
        RECT 37.110 111.100 39.625 111.240 ;
        RECT 39.805 111.240 40.175 111.285 ;
        RECT 43.065 111.240 43.355 111.285 ;
        RECT 39.805 111.100 43.355 111.240 ;
        RECT 37.110 111.055 37.400 111.100 ;
        RECT 39.805 111.055 40.175 111.100 ;
        RECT 43.065 111.055 43.355 111.100 ;
        RECT 43.985 111.240 44.275 111.285 ;
        RECT 45.845 111.240 46.135 111.285 ;
        RECT 43.985 111.100 46.135 111.240 ;
        RECT 43.985 111.055 44.275 111.100 ;
        RECT 45.845 111.055 46.135 111.100 ;
        RECT 55.905 111.240 56.275 111.285 ;
        RECT 59.165 111.240 59.455 111.285 ;
        RECT 55.905 111.100 59.455 111.240 ;
        RECT 55.905 111.055 56.275 111.100 ;
        RECT 59.165 111.055 59.455 111.100 ;
        RECT 60.085 111.240 60.375 111.285 ;
        RECT 61.945 111.240 62.235 111.285 ;
        RECT 60.085 111.100 62.235 111.240 ;
        RECT 60.085 111.055 60.375 111.100 ;
        RECT 61.945 111.055 62.235 111.100 ;
        RECT 66.535 111.240 66.855 111.300 ;
        RECT 70.690 111.240 70.980 111.285 ;
        RECT 79.965 111.240 80.105 111.440 ;
        RECT 81.040 111.395 81.330 111.440 ;
        RECT 92.310 111.395 92.600 111.440 ;
        RECT 98.290 111.580 98.580 111.625 ;
        RECT 99.655 111.580 99.975 111.640 ;
        RECT 98.290 111.440 99.975 111.580 ;
        RECT 98.290 111.395 98.580 111.440 ;
        RECT 99.655 111.380 99.975 111.440 ;
        RECT 86.315 111.285 86.635 111.300 ;
        RECT 66.535 111.100 69.525 111.240 ;
        RECT 39.855 111.040 40.175 111.055 ;
        RECT 36.190 110.715 36.480 110.945 ;
        RECT 41.665 110.900 41.955 110.945 ;
        RECT 43.985 110.900 44.200 111.055 ;
        RECT 55.955 111.040 56.275 111.055 ;
        RECT 41.665 110.760 44.200 110.900 ;
        RECT 44.455 110.900 44.775 110.960 ;
        RECT 44.930 110.900 45.220 110.945 ;
        RECT 44.455 110.760 45.220 110.900 ;
        RECT 41.665 110.715 41.955 110.760 ;
        RECT 44.455 110.700 44.775 110.760 ;
        RECT 44.930 110.715 45.220 110.760 ;
        RECT 49.070 110.900 49.360 110.945 ;
        RECT 51.355 110.900 51.675 110.960 ;
        RECT 49.070 110.760 51.675 110.900 ;
        RECT 49.070 110.715 49.360 110.760 ;
        RECT 51.355 110.700 51.675 110.760 ;
        RECT 57.765 110.900 58.055 110.945 ;
        RECT 60.085 110.900 60.300 111.055 ;
        RECT 66.535 111.040 66.855 111.100 ;
        RECT 57.765 110.760 60.300 110.900 ;
        RECT 57.765 110.715 58.055 110.760 ;
        RECT 61.015 110.700 61.335 110.960 ;
        RECT 63.315 110.700 63.635 110.960 ;
        RECT 68.375 110.900 68.695 110.960 ;
        RECT 68.850 110.900 69.140 110.945 ;
        RECT 68.375 110.760 69.140 110.900 ;
        RECT 69.385 110.900 69.525 111.100 ;
        RECT 70.690 111.100 80.105 111.240 ;
        RECT 83.045 111.240 83.335 111.285 ;
        RECT 86.305 111.240 86.635 111.285 ;
        RECT 83.045 111.100 86.635 111.240 ;
        RECT 70.690 111.055 70.980 111.100 ;
        RECT 75.290 110.900 75.580 110.945 ;
        RECT 69.385 110.760 75.580 110.900 ;
        RECT 68.375 110.700 68.695 110.760 ;
        RECT 68.850 110.715 69.140 110.760 ;
        RECT 75.290 110.715 75.580 110.760 ;
        RECT 75.735 110.700 76.055 110.960 ;
        RECT 79.045 110.945 79.185 111.100 ;
        RECT 83.045 111.055 83.335 111.100 ;
        RECT 86.305 111.055 86.635 111.100 ;
        RECT 86.315 111.040 86.635 111.055 ;
        RECT 87.225 111.240 87.515 111.285 ;
        RECT 89.085 111.240 89.375 111.285 ;
        RECT 95.990 111.240 96.280 111.285 ;
        RECT 87.225 111.100 89.375 111.240 ;
        RECT 87.225 111.055 87.515 111.100 ;
        RECT 89.085 111.055 89.375 111.100 ;
        RECT 89.625 111.100 96.280 111.240 ;
        RECT 78.970 110.715 79.260 110.945 ;
        RECT 79.430 110.900 79.720 110.945 ;
        RECT 79.875 110.900 80.195 110.960 ;
        RECT 79.430 110.760 80.195 110.900 ;
        RECT 79.430 110.715 79.720 110.760 ;
        RECT 79.875 110.700 80.195 110.760 ;
        RECT 80.350 110.900 80.640 110.945 ;
        RECT 84.015 110.900 84.335 110.960 ;
        RECT 80.350 110.760 84.335 110.900 ;
        RECT 80.350 110.715 80.640 110.760 ;
        RECT 84.015 110.700 84.335 110.760 ;
        RECT 84.905 110.900 85.195 110.945 ;
        RECT 87.225 110.900 87.440 111.055 ;
        RECT 84.905 110.760 87.440 110.900 ;
        RECT 87.695 110.900 88.015 110.960 ;
        RECT 89.625 110.900 89.765 111.100 ;
        RECT 95.990 111.055 96.280 111.100 ;
        RECT 96.435 111.240 96.755 111.300 ;
        RECT 101.035 111.240 101.355 111.300 ;
        RECT 96.435 111.100 101.355 111.240 ;
        RECT 96.435 111.040 96.755 111.100 ;
        RECT 101.035 111.040 101.355 111.100 ;
        RECT 87.695 110.760 89.765 110.900 ;
        RECT 90.010 110.900 90.300 110.945 ;
        RECT 90.915 110.900 91.235 110.960 ;
        RECT 94.135 110.900 94.455 110.960 ;
        RECT 105.175 110.900 105.495 110.960 ;
        RECT 90.010 110.760 94.455 110.900 ;
        RECT 84.905 110.715 85.195 110.760 ;
        RECT 87.695 110.700 88.015 110.760 ;
        RECT 90.010 110.715 90.300 110.760 ;
        RECT 90.915 110.700 91.235 110.760 ;
        RECT 94.135 110.700 94.455 110.760 ;
        RECT 101.355 110.760 105.495 110.900 ;
        RECT 27.895 110.560 28.215 110.620 ;
        RECT 37.800 110.560 38.090 110.605 ;
        RECT 42.615 110.560 42.935 110.620 ;
        RECT 27.895 110.420 42.935 110.560 ;
        RECT 27.895 110.360 28.215 110.420 ;
        RECT 37.800 110.375 38.090 110.420 ;
        RECT 42.615 110.360 42.935 110.420 ;
        RECT 46.770 110.560 47.060 110.605 ;
        RECT 47.215 110.560 47.535 110.620 ;
        RECT 46.770 110.420 47.535 110.560 ;
        RECT 46.770 110.375 47.060 110.420 ;
        RECT 47.215 110.360 47.535 110.420 ;
        RECT 59.635 110.560 59.955 110.620 ;
        RECT 62.870 110.560 63.160 110.605 ;
        RECT 69.770 110.560 70.060 110.605 ;
        RECT 74.370 110.560 74.660 110.605 ;
        RECT 59.635 110.420 63.160 110.560 ;
        RECT 59.635 110.360 59.955 110.420 ;
        RECT 62.870 110.375 63.160 110.420 ;
        RECT 68.005 110.420 74.660 110.560 ;
        RECT 75.825 110.560 75.965 110.700 ;
        RECT 87.785 110.560 87.925 110.700 ;
        RECT 75.825 110.420 87.925 110.560 ;
        RECT 88.170 110.560 88.460 110.605 ;
        RECT 88.170 110.420 90.685 110.560 ;
        RECT 31.130 110.220 31.420 110.265 ;
        RECT 39.855 110.220 40.175 110.280 ;
        RECT 31.130 110.080 40.175 110.220 ;
        RECT 31.130 110.035 31.420 110.080 ;
        RECT 39.855 110.020 40.175 110.080 ;
        RECT 41.665 110.220 41.955 110.265 ;
        RECT 44.445 110.220 44.735 110.265 ;
        RECT 46.305 110.220 46.595 110.265 ;
        RECT 41.665 110.080 46.595 110.220 ;
        RECT 41.665 110.035 41.955 110.080 ;
        RECT 44.445 110.035 44.735 110.080 ;
        RECT 46.305 110.035 46.595 110.080 ;
        RECT 57.765 110.220 58.055 110.265 ;
        RECT 60.545 110.220 60.835 110.265 ;
        RECT 62.405 110.220 62.695 110.265 ;
        RECT 57.765 110.080 62.695 110.220 ;
        RECT 57.765 110.035 58.055 110.080 ;
        RECT 60.545 110.035 60.835 110.080 ;
        RECT 62.405 110.035 62.695 110.080 ;
        RECT 32.955 109.680 33.275 109.940 ;
        RECT 33.415 109.880 33.735 109.940 ;
        RECT 35.730 109.880 36.020 109.925 ;
        RECT 33.415 109.740 36.020 109.880 ;
        RECT 33.415 109.680 33.735 109.740 ;
        RECT 35.730 109.695 36.020 109.740 ;
        RECT 38.015 109.880 38.335 109.940 ;
        RECT 42.155 109.880 42.475 109.940 ;
        RECT 38.015 109.740 42.475 109.880 ;
        RECT 38.015 109.680 38.335 109.740 ;
        RECT 42.155 109.680 42.475 109.740 ;
        RECT 48.610 109.880 48.900 109.925 ;
        RECT 49.055 109.880 49.375 109.940 ;
        RECT 48.610 109.740 49.375 109.880 ;
        RECT 48.610 109.695 48.900 109.740 ;
        RECT 49.055 109.680 49.375 109.740 ;
        RECT 55.495 109.880 55.815 109.940 ;
        RECT 68.005 109.880 68.145 110.420 ;
        RECT 69.770 110.375 70.060 110.420 ;
        RECT 74.370 110.375 74.660 110.420 ;
        RECT 88.170 110.375 88.460 110.420 ;
        RECT 74.445 110.220 74.585 110.375 ;
        RECT 90.545 110.265 90.685 110.420 ;
        RECT 92.770 110.375 93.060 110.605 ;
        RECT 93.675 110.560 93.995 110.620 ;
        RECT 95.530 110.560 95.820 110.605 ;
        RECT 93.675 110.420 95.820 110.560 ;
        RECT 84.905 110.220 85.195 110.265 ;
        RECT 87.685 110.220 87.975 110.265 ;
        RECT 89.545 110.220 89.835 110.265 ;
        RECT 74.445 110.080 84.705 110.220 ;
        RECT 55.495 109.740 68.145 109.880 ;
        RECT 55.495 109.680 55.815 109.740 ;
        RECT 68.375 109.680 68.695 109.940 ;
        RECT 72.975 109.680 73.295 109.940 ;
        RECT 77.115 109.880 77.435 109.940 ;
        RECT 77.590 109.880 77.880 109.925 ;
        RECT 77.115 109.740 77.880 109.880 ;
        RECT 84.565 109.880 84.705 110.080 ;
        RECT 84.905 110.080 89.835 110.220 ;
        RECT 84.905 110.035 85.195 110.080 ;
        RECT 87.685 110.035 87.975 110.080 ;
        RECT 89.545 110.035 89.835 110.080 ;
        RECT 90.470 110.035 90.760 110.265 ;
        RECT 92.845 110.220 92.985 110.375 ;
        RECT 93.675 110.360 93.995 110.420 ;
        RECT 95.530 110.375 95.820 110.420 ;
        RECT 95.055 110.220 95.375 110.280 ;
        RECT 98.275 110.220 98.595 110.280 ;
        RECT 92.845 110.080 98.595 110.220 ;
        RECT 95.055 110.020 95.375 110.080 ;
        RECT 98.275 110.020 98.595 110.080 ;
        RECT 88.155 109.880 88.475 109.940 ;
        RECT 84.565 109.740 88.475 109.880 ;
        RECT 77.115 109.680 77.435 109.740 ;
        RECT 77.590 109.695 77.880 109.740 ;
        RECT 88.155 109.680 88.475 109.740 ;
        RECT 89.995 109.880 90.315 109.940 ;
        RECT 101.355 109.880 101.495 110.760 ;
        RECT 105.175 110.700 105.495 110.760 ;
        RECT 89.995 109.740 101.495 109.880 ;
        RECT 89.995 109.680 90.315 109.740 ;
        RECT 17.605 109.060 112.465 109.540 ;
        RECT 32.510 108.860 32.800 108.905 ;
        RECT 32.955 108.860 33.275 108.920 ;
        RECT 46.755 108.860 47.075 108.920 ;
        RECT 32.510 108.720 33.275 108.860 ;
        RECT 32.510 108.675 32.800 108.720 ;
        RECT 32.955 108.660 33.275 108.720 ;
        RECT 41.785 108.720 47.075 108.860 ;
        RECT 30.195 108.520 30.515 108.580 ;
        RECT 30.195 108.380 37.785 108.520 ;
        RECT 30.195 108.320 30.515 108.380 ;
        RECT 36.175 108.180 36.495 108.240 ;
        RECT 37.645 108.225 37.785 108.380 ;
        RECT 33.505 108.040 36.495 108.180 ;
        RECT 24.215 107.840 24.535 107.900 ;
        RECT 33.505 107.885 33.645 108.040 ;
        RECT 36.175 107.980 36.495 108.040 ;
        RECT 37.110 107.995 37.400 108.225 ;
        RECT 37.570 108.180 37.860 108.225 ;
        RECT 37.570 108.040 39.625 108.180 ;
        RECT 37.570 107.995 37.860 108.040 ;
        RECT 31.130 107.840 31.420 107.885 ;
        RECT 24.215 107.700 31.420 107.840 ;
        RECT 24.215 107.640 24.535 107.700 ;
        RECT 31.130 107.655 31.420 107.700 ;
        RECT 33.430 107.655 33.720 107.885 ;
        RECT 34.350 107.840 34.640 107.885 ;
        RECT 36.635 107.840 36.955 107.900 ;
        RECT 34.350 107.700 36.955 107.840 ;
        RECT 34.350 107.655 34.640 107.700 ;
        RECT 36.635 107.640 36.955 107.700 ;
        RECT 37.185 107.500 37.325 107.995 ;
        RECT 38.015 107.640 38.335 107.900 ;
        RECT 39.485 107.840 39.625 108.040 ;
        RECT 41.235 107.980 41.555 108.240 ;
        RECT 41.785 108.225 41.925 108.720 ;
        RECT 46.755 108.660 47.075 108.720 ;
        RECT 52.735 108.860 53.055 108.920 ;
        RECT 58.715 108.860 59.035 108.920 ;
        RECT 60.110 108.860 60.400 108.905 ;
        RECT 52.735 108.720 58.485 108.860 ;
        RECT 52.735 108.660 53.055 108.720 ;
        RECT 44.010 108.335 44.300 108.565 ;
        RECT 48.565 108.520 48.855 108.565 ;
        RECT 51.345 108.520 51.635 108.565 ;
        RECT 53.205 108.520 53.495 108.565 ;
        RECT 48.565 108.380 53.495 108.520 ;
        RECT 58.345 108.520 58.485 108.720 ;
        RECT 58.715 108.720 60.400 108.860 ;
        RECT 58.715 108.660 59.035 108.720 ;
        RECT 60.110 108.675 60.400 108.720 ;
        RECT 64.235 108.860 64.555 108.920 ;
        RECT 65.860 108.860 66.150 108.905 ;
        RECT 64.235 108.720 66.150 108.860 ;
        RECT 64.235 108.660 64.555 108.720 ;
        RECT 65.860 108.675 66.150 108.720 ;
        RECT 84.260 108.860 84.550 108.905 ;
        RECT 87.695 108.860 88.015 108.920 ;
        RECT 84.260 108.720 88.015 108.860 ;
        RECT 84.260 108.675 84.550 108.720 ;
        RECT 87.695 108.660 88.015 108.720 ;
        RECT 98.275 108.860 98.595 108.920 ;
        RECT 99.900 108.860 100.190 108.905 ;
        RECT 98.275 108.720 100.190 108.860 ;
        RECT 98.275 108.660 98.595 108.720 ;
        RECT 99.900 108.675 100.190 108.720 ;
        RECT 61.950 108.520 62.240 108.565 ;
        RECT 63.315 108.520 63.635 108.580 ;
        RECT 58.345 108.380 63.635 108.520 ;
        RECT 48.565 108.335 48.855 108.380 ;
        RECT 51.345 108.335 51.635 108.380 ;
        RECT 53.205 108.335 53.495 108.380 ;
        RECT 61.950 108.335 62.240 108.380 ;
        RECT 41.710 107.995 42.000 108.225 ;
        RECT 44.085 108.180 44.225 108.335 ;
        RECT 63.315 108.320 63.635 108.380 ;
        RECT 69.725 108.520 70.015 108.565 ;
        RECT 72.505 108.520 72.795 108.565 ;
        RECT 74.365 108.520 74.655 108.565 ;
        RECT 69.725 108.380 74.655 108.520 ;
        RECT 69.725 108.335 70.015 108.380 ;
        RECT 72.505 108.335 72.795 108.380 ;
        RECT 74.365 108.335 74.655 108.380 ;
        RECT 75.755 108.520 76.045 108.565 ;
        RECT 77.615 108.520 77.905 108.565 ;
        RECT 80.395 108.520 80.685 108.565 ;
        RECT 75.755 108.380 80.685 108.520 ;
        RECT 75.755 108.335 76.045 108.380 ;
        RECT 77.615 108.335 77.905 108.380 ;
        RECT 80.395 108.335 80.685 108.380 ;
        RECT 88.155 108.320 88.475 108.580 ;
        RECT 91.395 108.520 91.685 108.565 ;
        RECT 93.255 108.520 93.545 108.565 ;
        RECT 96.035 108.520 96.325 108.565 ;
        RECT 91.395 108.380 96.325 108.520 ;
        RECT 91.395 108.335 91.685 108.380 ;
        RECT 93.255 108.335 93.545 108.380 ;
        RECT 96.035 108.335 96.325 108.380 ;
        RECT 97.815 108.520 98.135 108.580 ;
        RECT 101.050 108.520 101.340 108.565 ;
        RECT 97.815 108.380 101.340 108.520 ;
        RECT 97.815 108.320 98.135 108.380 ;
        RECT 101.050 108.335 101.340 108.380 ;
        RECT 51.830 108.180 52.120 108.225 ;
        RECT 44.085 108.040 52.120 108.180 ;
        RECT 51.830 107.995 52.120 108.040 ;
        RECT 55.495 108.180 55.815 108.240 ;
        RECT 56.890 108.180 57.180 108.225 ;
        RECT 55.495 108.040 57.180 108.180 ;
        RECT 55.495 107.980 55.815 108.040 ;
        RECT 56.890 107.995 57.180 108.040 ;
        RECT 72.975 107.980 73.295 108.240 ;
        RECT 77.115 107.980 77.435 108.240 ;
        RECT 90.915 107.980 91.235 108.240 ;
        RECT 42.170 107.840 42.460 107.885 ;
        RECT 44.700 107.840 44.990 107.885 ;
        RECT 39.485 107.700 44.990 107.840 ;
        RECT 42.170 107.655 42.460 107.700 ;
        RECT 44.700 107.655 44.990 107.700 ;
        RECT 48.565 107.840 48.855 107.885 ;
        RECT 48.565 107.700 51.100 107.840 ;
        RECT 48.565 107.655 48.855 107.700 ;
        RECT 41.235 107.500 41.555 107.560 ;
        RECT 37.185 107.360 41.555 107.500 ;
        RECT 41.235 107.300 41.555 107.360 ;
        RECT 42.615 107.500 42.935 107.560 ;
        RECT 46.705 107.500 46.995 107.545 ;
        RECT 49.055 107.500 49.375 107.560 ;
        RECT 50.885 107.545 51.100 107.700 ;
        RECT 53.670 107.655 53.960 107.885 ;
        RECT 58.270 107.840 58.560 107.885 ;
        RECT 60.555 107.840 60.875 107.900 ;
        RECT 58.270 107.700 60.875 107.840 ;
        RECT 58.270 107.655 58.560 107.700 ;
        RECT 49.965 107.500 50.255 107.545 ;
        RECT 42.615 107.360 46.065 107.500 ;
        RECT 42.615 107.300 42.935 107.360 ;
        RECT 31.590 107.160 31.880 107.205 ;
        RECT 37.555 107.160 37.875 107.220 ;
        RECT 31.590 107.020 37.875 107.160 ;
        RECT 31.590 106.975 31.880 107.020 ;
        RECT 37.555 106.960 37.875 107.020 ;
        RECT 39.870 107.160 40.160 107.205 ;
        RECT 45.375 107.160 45.695 107.220 ;
        RECT 39.870 107.020 45.695 107.160 ;
        RECT 45.925 107.160 46.065 107.360 ;
        RECT 46.705 107.360 50.255 107.500 ;
        RECT 46.705 107.315 46.995 107.360 ;
        RECT 49.055 107.300 49.375 107.360 ;
        RECT 49.965 107.315 50.255 107.360 ;
        RECT 50.885 107.500 51.175 107.545 ;
        RECT 52.745 107.500 53.035 107.545 ;
        RECT 50.885 107.360 53.035 107.500 ;
        RECT 53.745 107.500 53.885 107.655 ;
        RECT 60.555 107.640 60.875 107.700 ;
        RECT 61.030 107.840 61.320 107.885 ;
        RECT 61.475 107.840 61.795 107.900 ;
        RECT 61.030 107.700 61.795 107.840 ;
        RECT 61.030 107.655 61.320 107.700 ;
        RECT 61.475 107.640 61.795 107.700 ;
        RECT 69.725 107.840 70.015 107.885 ;
        RECT 74.830 107.840 75.120 107.885 ;
        RECT 75.275 107.840 75.595 107.900 ;
        RECT 80.395 107.840 80.685 107.885 ;
        RECT 69.725 107.700 72.260 107.840 ;
        RECT 69.725 107.655 70.015 107.700 ;
        RECT 59.635 107.500 59.955 107.560 ;
        RECT 53.745 107.360 59.955 107.500 ;
        RECT 50.885 107.315 51.175 107.360 ;
        RECT 52.745 107.315 53.035 107.360 ;
        RECT 59.635 107.300 59.955 107.360 ;
        RECT 67.865 107.500 68.155 107.545 ;
        RECT 68.375 107.500 68.695 107.560 ;
        RECT 72.045 107.545 72.260 107.700 ;
        RECT 74.830 107.700 75.595 107.840 ;
        RECT 74.830 107.655 75.120 107.700 ;
        RECT 75.275 107.640 75.595 107.700 ;
        RECT 78.150 107.700 80.685 107.840 ;
        RECT 78.150 107.545 78.365 107.700 ;
        RECT 80.395 107.655 80.685 107.700 ;
        RECT 85.870 107.655 86.160 107.885 ;
        RECT 86.775 107.840 87.095 107.900 ;
        RECT 87.250 107.840 87.540 107.885 ;
        RECT 86.775 107.700 87.540 107.840 ;
        RECT 71.125 107.500 71.415 107.545 ;
        RECT 67.865 107.360 71.415 107.500 ;
        RECT 67.865 107.315 68.155 107.360 ;
        RECT 68.375 107.300 68.695 107.360 ;
        RECT 71.125 107.315 71.415 107.360 ;
        RECT 72.045 107.500 72.335 107.545 ;
        RECT 73.905 107.500 74.195 107.545 ;
        RECT 72.045 107.360 74.195 107.500 ;
        RECT 72.045 107.315 72.335 107.360 ;
        RECT 73.905 107.315 74.195 107.360 ;
        RECT 76.215 107.500 76.505 107.545 ;
        RECT 78.075 107.500 78.365 107.545 ;
        RECT 78.995 107.500 79.285 107.545 ;
        RECT 82.255 107.500 82.545 107.545 ;
        RECT 76.215 107.360 78.365 107.500 ;
        RECT 76.215 107.315 76.505 107.360 ;
        RECT 78.075 107.315 78.365 107.360 ;
        RECT 78.585 107.360 82.545 107.500 ;
        RECT 85.945 107.500 86.085 107.655 ;
        RECT 86.775 107.640 87.095 107.700 ;
        RECT 87.250 107.655 87.540 107.700 ;
        RECT 89.550 107.840 89.840 107.885 ;
        RECT 89.995 107.840 90.315 107.900 ;
        RECT 89.550 107.700 90.315 107.840 ;
        RECT 89.550 107.655 89.840 107.700 ;
        RECT 89.625 107.500 89.765 107.655 ;
        RECT 89.995 107.640 90.315 107.700 ;
        RECT 91.375 107.840 91.695 107.900 ;
        RECT 92.770 107.840 93.060 107.885 ;
        RECT 96.035 107.840 96.325 107.885 ;
        RECT 91.375 107.700 93.060 107.840 ;
        RECT 91.375 107.640 91.695 107.700 ;
        RECT 92.770 107.655 93.060 107.700 ;
        RECT 93.790 107.700 96.325 107.840 ;
        RECT 93.790 107.545 94.005 107.700 ;
        RECT 96.035 107.655 96.325 107.700 ;
        RECT 101.510 107.840 101.800 107.885 ;
        RECT 105.175 107.840 105.495 107.900 ;
        RECT 101.510 107.700 105.495 107.840 ;
        RECT 101.510 107.655 101.800 107.700 ;
        RECT 105.175 107.640 105.495 107.700 ;
        RECT 85.945 107.360 89.765 107.500 ;
        RECT 91.855 107.500 92.145 107.545 ;
        RECT 93.715 107.500 94.005 107.545 ;
        RECT 94.635 107.500 94.925 107.545 ;
        RECT 97.895 107.500 98.185 107.545 ;
        RECT 91.855 107.360 94.005 107.500 ;
        RECT 57.810 107.160 58.100 107.205 ;
        RECT 45.925 107.020 58.100 107.160 ;
        RECT 39.870 106.975 40.160 107.020 ;
        RECT 45.375 106.960 45.695 107.020 ;
        RECT 57.810 106.975 58.100 107.020 ;
        RECT 74.815 107.160 75.135 107.220 ;
        RECT 78.585 107.160 78.725 107.360 ;
        RECT 78.995 107.315 79.285 107.360 ;
        RECT 82.255 107.315 82.545 107.360 ;
        RECT 91.855 107.315 92.145 107.360 ;
        RECT 93.715 107.315 94.005 107.360 ;
        RECT 94.225 107.360 98.185 107.500 ;
        RECT 74.815 107.020 78.725 107.160 ;
        RECT 85.410 107.160 85.700 107.205 ;
        RECT 85.855 107.160 86.175 107.220 ;
        RECT 85.410 107.020 86.175 107.160 ;
        RECT 74.815 106.960 75.135 107.020 ;
        RECT 85.410 106.975 85.700 107.020 ;
        RECT 85.855 106.960 86.175 107.020 ;
        RECT 90.010 107.160 90.300 107.205 ;
        RECT 94.225 107.160 94.365 107.360 ;
        RECT 94.635 107.315 94.925 107.360 ;
        RECT 97.895 107.315 98.185 107.360 ;
        RECT 90.010 107.020 94.365 107.160 ;
        RECT 90.010 106.975 90.300 107.020 ;
        RECT 18.165 106.340 112.465 106.820 ;
        RECT 135.660 106.690 136.800 133.400 ;
        RECT 133.100 106.600 136.850 106.690 ;
        RECT 38.015 106.185 38.335 106.200 ;
        RECT 38.015 105.955 38.550 106.185 ;
        RECT 38.015 105.940 38.335 105.955 ;
        RECT 74.815 105.940 75.135 106.200 ;
        RECT 83.555 106.140 83.875 106.200 ;
        RECT 83.555 106.000 95.285 106.140 ;
        RECT 83.555 105.940 83.875 106.000 ;
        RECT 37.555 105.800 37.875 105.860 ;
        RECT 40.265 105.800 40.555 105.845 ;
        RECT 43.525 105.800 43.815 105.845 ;
        RECT 37.555 105.660 43.815 105.800 ;
        RECT 37.555 105.600 37.875 105.660 ;
        RECT 40.265 105.615 40.555 105.660 ;
        RECT 43.525 105.615 43.815 105.660 ;
        RECT 44.445 105.800 44.735 105.845 ;
        RECT 46.305 105.800 46.595 105.845 ;
        RECT 44.445 105.660 46.595 105.800 ;
        RECT 44.445 105.615 44.735 105.660 ;
        RECT 46.305 105.615 46.595 105.660 ;
        RECT 52.390 105.800 52.680 105.845 ;
        RECT 54.575 105.800 54.895 105.860 ;
        RECT 55.630 105.800 56.280 105.845 ;
        RECT 52.390 105.660 56.280 105.800 ;
        RECT 52.390 105.615 52.980 105.660 ;
        RECT 42.125 105.460 42.415 105.505 ;
        RECT 44.445 105.460 44.660 105.615 ;
        RECT 42.125 105.320 44.660 105.460 ;
        RECT 42.125 105.275 42.415 105.320 ;
        RECT 45.375 105.260 45.695 105.520 ;
        RECT 47.215 105.260 47.535 105.520 ;
        RECT 52.690 105.300 52.980 105.615 ;
        RECT 54.575 105.600 54.895 105.660 ;
        RECT 55.630 105.615 56.280 105.660 ;
        RECT 58.255 105.600 58.575 105.860 ;
        RECT 62.970 105.800 63.260 105.845 ;
        RECT 66.210 105.800 66.860 105.845 ;
        RECT 62.970 105.660 66.860 105.800 ;
        RECT 62.970 105.615 63.560 105.660 ;
        RECT 66.210 105.615 66.860 105.660 ;
        RECT 63.270 105.520 63.560 105.615 ;
        RECT 68.835 105.600 69.155 105.860 ;
        RECT 78.610 105.800 78.900 105.845 ;
        RECT 79.415 105.800 79.735 105.860 ;
        RECT 81.850 105.800 82.500 105.845 ;
        RECT 78.610 105.660 82.500 105.800 ;
        RECT 78.610 105.615 79.200 105.660 ;
        RECT 53.770 105.460 54.060 105.505 ;
        RECT 57.350 105.460 57.640 105.505 ;
        RECT 59.185 105.460 59.475 105.505 ;
        RECT 53.770 105.320 59.475 105.460 ;
        RECT 53.770 105.275 54.060 105.320 ;
        RECT 57.350 105.275 57.640 105.320 ;
        RECT 59.185 105.275 59.475 105.320 ;
        RECT 59.635 105.260 59.955 105.520 ;
        RECT 63.270 105.300 63.635 105.520 ;
        RECT 63.315 105.260 63.635 105.300 ;
        RECT 64.350 105.460 64.640 105.505 ;
        RECT 67.930 105.460 68.220 105.505 ;
        RECT 69.765 105.460 70.055 105.505 ;
        RECT 64.350 105.320 70.055 105.460 ;
        RECT 64.350 105.275 64.640 105.320 ;
        RECT 67.930 105.275 68.220 105.320 ;
        RECT 69.765 105.275 70.055 105.320 ;
        RECT 73.895 105.460 74.215 105.520 ;
        RECT 74.370 105.460 74.660 105.505 ;
        RECT 73.895 105.320 74.660 105.460 ;
        RECT 73.895 105.260 74.215 105.320 ;
        RECT 74.370 105.275 74.660 105.320 ;
        RECT 75.750 105.460 76.040 105.505 ;
        RECT 78.035 105.460 78.355 105.520 ;
        RECT 75.750 105.320 78.355 105.460 ;
        RECT 75.750 105.275 76.040 105.320 ;
        RECT 78.035 105.260 78.355 105.320 ;
        RECT 78.910 105.300 79.200 105.615 ;
        RECT 79.415 105.600 79.735 105.660 ;
        RECT 81.850 105.615 82.500 105.660 ;
        RECT 84.475 105.600 84.795 105.860 ;
        RECT 85.855 105.800 86.175 105.860 ;
        RECT 95.145 105.845 95.285 106.000 ;
        RECT 89.190 105.800 89.480 105.845 ;
        RECT 92.430 105.800 93.080 105.845 ;
        RECT 85.855 105.660 93.080 105.800 ;
        RECT 85.855 105.600 86.175 105.660 ;
        RECT 89.190 105.615 89.780 105.660 ;
        RECT 92.430 105.615 93.080 105.660 ;
        RECT 95.070 105.615 95.360 105.845 ;
        RECT 129.700 105.630 136.850 106.600 ;
        RECT 79.990 105.460 80.280 105.505 ;
        RECT 83.570 105.460 83.860 105.505 ;
        RECT 85.405 105.460 85.695 105.505 ;
        RECT 79.990 105.320 85.695 105.460 ;
        RECT 79.990 105.275 80.280 105.320 ;
        RECT 83.570 105.275 83.860 105.320 ;
        RECT 85.405 105.275 85.695 105.320 ;
        RECT 89.490 105.300 89.780 105.615 ;
        RECT 90.570 105.460 90.860 105.505 ;
        RECT 94.150 105.460 94.440 105.505 ;
        RECT 95.985 105.460 96.275 105.505 ;
        RECT 133.100 105.500 136.850 105.630 ;
        RECT 90.570 105.320 96.275 105.460 ;
        RECT 90.570 105.275 90.860 105.320 ;
        RECT 94.150 105.275 94.440 105.320 ;
        RECT 95.985 105.275 96.275 105.320 ;
        RECT 49.530 105.120 49.820 105.165 ;
        RECT 50.435 105.120 50.755 105.180 ;
        RECT 49.530 104.980 50.755 105.120 ;
        RECT 49.530 104.935 49.820 104.980 ;
        RECT 50.435 104.920 50.755 104.980 ;
        RECT 60.095 104.920 60.415 105.180 ;
        RECT 70.230 105.120 70.520 105.165 ;
        RECT 75.275 105.120 75.595 105.180 ;
        RECT 85.870 105.120 86.160 105.165 ;
        RECT 70.230 104.980 86.160 105.120 ;
        RECT 70.230 104.935 70.520 104.980 ;
        RECT 75.275 104.920 75.595 104.980 ;
        RECT 85.870 104.935 86.160 104.980 ;
        RECT 86.330 104.935 86.620 105.165 ;
        RECT 94.595 105.120 94.915 105.180 ;
        RECT 96.450 105.120 96.740 105.165 ;
        RECT 94.595 104.980 96.740 105.120 ;
        RECT 42.125 104.780 42.415 104.825 ;
        RECT 44.905 104.780 45.195 104.825 ;
        RECT 46.765 104.780 47.055 104.825 ;
        RECT 42.125 104.640 47.055 104.780 ;
        RECT 42.125 104.595 42.415 104.640 ;
        RECT 44.905 104.595 45.195 104.640 ;
        RECT 46.765 104.595 47.055 104.640 ;
        RECT 53.770 104.780 54.060 104.825 ;
        RECT 56.890 104.780 57.180 104.825 ;
        RECT 58.780 104.780 59.070 104.825 ;
        RECT 53.770 104.640 59.070 104.780 ;
        RECT 53.770 104.595 54.060 104.640 ;
        RECT 56.890 104.595 57.180 104.640 ;
        RECT 58.780 104.595 59.070 104.640 ;
        RECT 64.350 104.780 64.640 104.825 ;
        RECT 67.470 104.780 67.760 104.825 ;
        RECT 69.360 104.780 69.650 104.825 ;
        RECT 64.350 104.640 69.650 104.780 ;
        RECT 64.350 104.595 64.640 104.640 ;
        RECT 67.470 104.595 67.760 104.640 ;
        RECT 69.360 104.595 69.650 104.640 ;
        RECT 79.990 104.780 80.280 104.825 ;
        RECT 83.110 104.780 83.400 104.825 ;
        RECT 85.000 104.780 85.290 104.825 ;
        RECT 79.990 104.640 85.290 104.780 ;
        RECT 79.990 104.595 80.280 104.640 ;
        RECT 83.110 104.595 83.400 104.640 ;
        RECT 85.000 104.595 85.290 104.640 ;
        RECT 82.635 104.440 82.955 104.500 ;
        RECT 86.405 104.440 86.545 104.935 ;
        RECT 94.595 104.920 94.915 104.980 ;
        RECT 96.450 104.935 96.740 104.980 ;
        RECT 90.570 104.780 90.860 104.825 ;
        RECT 93.690 104.780 93.980 104.825 ;
        RECT 95.580 104.780 95.870 104.825 ;
        RECT 90.570 104.640 95.870 104.780 ;
        RECT 90.570 104.595 90.860 104.640 ;
        RECT 93.690 104.595 93.980 104.640 ;
        RECT 95.580 104.595 95.870 104.640 ;
        RECT 82.635 104.300 86.545 104.440 ;
        RECT 82.635 104.240 82.955 104.300 ;
        RECT 17.605 103.620 112.465 104.100 ;
        RECT 54.130 103.420 54.420 103.465 ;
        RECT 54.575 103.420 54.895 103.480 ;
        RECT 54.130 103.280 54.895 103.420 ;
        RECT 54.130 103.235 54.420 103.280 ;
        RECT 54.575 103.220 54.895 103.280 ;
        RECT 62.870 103.420 63.160 103.465 ;
        RECT 63.315 103.420 63.635 103.480 ;
        RECT 62.870 103.280 63.635 103.420 ;
        RECT 62.870 103.235 63.160 103.280 ;
        RECT 63.315 103.220 63.635 103.280 ;
        RECT 79.415 103.420 79.735 103.480 ;
        RECT 80.350 103.420 80.640 103.465 ;
        RECT 79.415 103.280 80.640 103.420 ;
        RECT 79.415 103.220 79.735 103.280 ;
        RECT 80.350 103.235 80.640 103.280 ;
        RECT 53.195 102.400 53.515 102.460 ;
        RECT 54.590 102.400 54.880 102.445 ;
        RECT 62.410 102.400 62.700 102.445 ;
        RECT 53.195 102.260 62.700 102.400 ;
        RECT 53.195 102.200 53.515 102.260 ;
        RECT 54.590 102.215 54.880 102.260 ;
        RECT 62.410 102.215 62.700 102.260 ;
        RECT 80.795 102.200 81.115 102.460 ;
        RECT 18.165 100.900 112.465 101.380 ;
        RECT 133.330 76.630 136.060 77.830 ;
        RECT 137.920 77.810 143.450 77.960 ;
        RECT 21.115 74.380 23.065 74.390 ;
        RECT 19.415 73.240 23.065 74.380 ;
        RECT 19.415 73.230 21.125 73.240 ;
        RECT 28.135 73.230 30.305 74.410 ;
        RECT 32.315 74.390 34.265 74.400 ;
        RECT 30.615 73.250 34.265 74.390 ;
        RECT 30.615 73.240 32.325 73.250 ;
        RECT 39.425 73.200 41.595 74.380 ;
        RECT 43.535 74.360 45.485 74.370 ;
        RECT 41.835 73.220 45.485 74.360 ;
        RECT 54.785 74.340 56.735 74.350 ;
        RECT 41.835 73.210 43.545 73.220 ;
        RECT 3.910 73.080 6.100 73.190 ;
        RECT 50.005 73.140 52.175 74.320 ;
        RECT 53.085 73.200 56.735 74.340 ;
        RECT 53.085 73.190 54.795 73.200 ;
        RECT 61.425 73.170 63.595 74.350 ;
        RECT 66.005 74.330 67.955 74.340 ;
        RECT 64.305 73.190 67.955 74.330 ;
        RECT 64.305 73.180 66.015 73.190 ;
        RECT 72.535 73.180 74.705 74.360 ;
        RECT 77.245 74.320 79.195 74.330 ;
        RECT 75.545 73.180 79.195 74.320 ;
        RECT 75.545 73.170 77.255 73.180 ;
        RECT 83.805 73.170 85.975 74.350 ;
        RECT 88.495 74.330 90.445 74.340 ;
        RECT 86.795 73.190 90.445 74.330 ;
        RECT 99.775 74.320 101.725 74.330 ;
        RECT 86.795 73.180 88.505 73.190 ;
        RECT 94.995 73.110 97.165 74.290 ;
        RECT 98.075 73.180 101.725 74.320 ;
        RECT 98.075 73.170 99.785 73.180 ;
        RECT 106.405 73.160 108.575 74.340 ;
        RECT 111.045 74.320 112.995 74.330 ;
        RECT 109.345 73.180 112.995 74.320 ;
        RECT 109.345 73.170 111.055 73.180 ;
        RECT 117.605 73.160 119.775 74.340 ;
        RECT 122.295 74.320 124.245 74.330 ;
        RECT 120.595 73.180 124.245 74.320 ;
        RECT 129.455 73.240 131.625 74.420 ;
        RECT 120.595 73.170 122.305 73.180 ;
        RECT 3.910 72.820 12.240 73.080 ;
        RECT 29.635 72.840 43.235 72.850 ;
        RECT 18.435 72.820 43.235 72.840 ;
        RECT 3.910 72.800 54.455 72.820 ;
        RECT 3.910 72.790 65.705 72.800 ;
        RECT 133.960 72.790 135.640 76.630 ;
        RECT 137.190 76.610 143.450 77.810 ;
        RECT 137.920 75.460 143.450 76.610 ;
        RECT 3.910 72.780 76.925 72.790 ;
        RECT 85.815 72.780 99.415 72.790 ;
        RECT 132.085 72.780 140.600 72.790 ;
        RECT 3.910 71.700 140.600 72.780 ;
        RECT 3.910 71.690 32.035 71.700 ;
        RECT 3.910 71.670 19.135 71.690 ;
        RECT 40.855 71.670 140.600 71.700 ;
        RECT 3.910 71.500 12.240 71.670 ;
        RECT 52.105 71.650 140.600 71.670 ;
        RECT 63.325 71.640 140.600 71.650 ;
        RECT 74.565 71.630 88.165 71.640 ;
        RECT 97.095 71.630 133.215 71.640 ;
        RECT 3.910 71.370 6.100 71.500 ;
        RECT 10.800 71.180 11.950 71.500 ;
        RECT 10.800 69.480 11.915 71.180 ;
        RECT 29.635 71.170 43.285 71.180 ;
        RECT 15.510 71.155 17.040 71.160 ;
        RECT 18.435 71.155 43.285 71.170 ;
        RECT 12.285 71.150 43.285 71.155 ;
        RECT 12.285 71.130 54.505 71.150 ;
        RECT 141.810 71.140 143.230 75.460 ;
        RECT 12.285 71.120 65.755 71.130 ;
        RECT 12.285 71.110 76.975 71.120 ;
        RECT 85.815 71.110 99.465 71.120 ;
        RECT 140.220 71.110 143.240 71.140 ;
        RECT 12.285 70.030 143.240 71.110 ;
        RECT 12.285 70.020 32.085 70.030 ;
        RECT 12.285 70.005 19.375 70.020 ;
        RECT 10.800 13.800 11.950 69.480 ;
        RECT 12.320 15.450 13.470 70.005 ;
        RECT 15.510 68.660 17.040 70.005 ;
        RECT 40.855 70.000 143.240 70.030 ;
        RECT 52.105 69.980 143.240 70.000 ;
        RECT 63.325 69.970 143.240 69.980 ;
        RECT 74.565 69.960 88.215 69.970 ;
        RECT 97.095 69.960 143.240 69.970 ;
        RECT 140.220 69.910 143.240 69.960 ;
        RECT 29.645 69.670 43.315 69.680 ;
        RECT 18.445 69.650 43.315 69.670 ;
        RECT 18.445 69.630 54.535 69.650 ;
        RECT 18.445 69.620 65.785 69.630 ;
        RECT 139.590 69.620 150.610 69.640 ;
        RECT 18.445 69.610 77.005 69.620 ;
        RECT 85.825 69.610 99.495 69.620 ;
        RECT 132.155 69.610 150.610 69.620 ;
        RECT 18.445 69.570 150.610 69.610 ;
        RECT 18.445 68.530 150.740 69.570 ;
        RECT 18.445 68.520 32.115 68.530 ;
        RECT 40.865 68.500 150.740 68.530 ;
        RECT 52.115 68.490 143.320 68.500 ;
        RECT 52.115 68.480 140.670 68.490 ;
        RECT 63.335 68.470 140.670 68.480 ;
        RECT 74.575 68.460 88.245 68.470 ;
        RECT 97.105 68.460 133.295 68.470 ;
        RECT 141.080 68.450 142.300 68.490 ;
        RECT 149.360 68.470 150.740 68.500 ;
        RECT 29.655 68.100 43.325 68.110 ;
        RECT 13.950 68.080 43.325 68.100 ;
        RECT 13.950 68.060 54.545 68.080 ;
        RECT 13.950 68.050 65.795 68.060 ;
        RECT 13.950 68.040 77.015 68.050 ;
        RECT 85.835 68.040 99.505 68.050 ;
        RECT 139.530 68.040 143.320 68.060 ;
        RECT 13.950 66.960 152.870 68.040 ;
        RECT 13.950 66.950 32.125 66.960 ;
        RECT 13.950 18.530 15.100 66.950 ;
        RECT 40.875 66.930 152.870 66.960 ;
        RECT 52.125 66.910 152.870 66.930 ;
        RECT 63.345 66.900 152.870 66.910 ;
        RECT 74.585 66.890 88.255 66.900 ;
        RECT 97.115 66.890 143.320 66.900 ;
        RECT 141.030 66.770 142.490 66.890 ;
        RECT 21.405 65.510 26.555 65.790 ;
        RECT 27.815 65.490 28.965 65.800 ;
        RECT 32.605 65.520 37.755 65.800 ;
        RECT 39.015 65.500 40.165 65.810 ;
        RECT 43.825 65.490 48.975 65.770 ;
        RECT 50.235 65.470 51.385 65.780 ;
        RECT 149.460 65.760 150.600 65.780 ;
        RECT 55.075 65.470 60.225 65.750 ;
        RECT 61.485 65.450 62.635 65.760 ;
        RECT 66.295 65.460 71.445 65.740 ;
        RECT 72.705 65.440 73.855 65.750 ;
        RECT 77.535 65.450 82.685 65.730 ;
        RECT 83.945 65.430 85.095 65.740 ;
        RECT 88.785 65.460 93.935 65.740 ;
        RECT 95.195 65.440 96.345 65.750 ;
        RECT 100.065 65.450 105.215 65.730 ;
        RECT 106.475 65.430 107.625 65.740 ;
        RECT 111.335 65.450 116.485 65.730 ;
        RECT 117.745 65.430 118.895 65.740 ;
        RECT 122.585 65.450 127.735 65.730 ;
        RECT 128.995 65.430 130.145 65.740 ;
        RECT 133.315 65.430 138.455 65.690 ;
        RECT 21.205 65.140 21.435 65.320 ;
        RECT 26.495 65.190 26.725 65.320 ;
        RECT 21.125 55.220 21.485 65.140 ;
        RECT 26.435 55.240 26.805 65.190 ;
        RECT 27.635 65.150 27.865 65.320 ;
        RECT 27.565 55.200 27.935 65.150 ;
        RECT 28.925 65.140 29.155 65.320 ;
        RECT 32.405 65.150 32.635 65.330 ;
        RECT 37.695 65.200 37.925 65.330 ;
        RECT 28.835 55.250 29.255 65.140 ;
        RECT 32.325 55.230 32.685 65.150 ;
        RECT 37.635 55.250 38.005 65.200 ;
        RECT 38.835 65.160 39.065 65.330 ;
        RECT 38.765 55.210 39.135 65.160 ;
        RECT 40.125 65.150 40.355 65.330 ;
        RECT 40.035 55.260 40.455 65.150 ;
        RECT 43.625 65.120 43.855 65.300 ;
        RECT 48.915 65.170 49.145 65.300 ;
        RECT 43.545 55.200 43.905 65.120 ;
        RECT 48.855 55.220 49.225 65.170 ;
        RECT 50.055 65.130 50.285 65.300 ;
        RECT 49.985 55.180 50.355 65.130 ;
        RECT 51.345 65.120 51.575 65.300 ;
        RECT 51.255 55.230 51.675 65.120 ;
        RECT 54.875 65.100 55.105 65.280 ;
        RECT 60.165 65.150 60.395 65.280 ;
        RECT 54.795 55.180 55.155 65.100 ;
        RECT 60.105 55.200 60.475 65.150 ;
        RECT 61.305 65.110 61.535 65.280 ;
        RECT 61.235 55.160 61.605 65.110 ;
        RECT 62.595 65.100 62.825 65.280 ;
        RECT 62.505 55.210 62.925 65.100 ;
        RECT 66.095 65.090 66.325 65.270 ;
        RECT 71.385 65.140 71.615 65.270 ;
        RECT 66.015 55.170 66.375 65.090 ;
        RECT 71.325 55.190 71.695 65.140 ;
        RECT 72.525 65.100 72.755 65.270 ;
        RECT 72.455 55.150 72.825 65.100 ;
        RECT 73.815 65.090 74.045 65.270 ;
        RECT 73.725 55.200 74.145 65.090 ;
        RECT 77.335 65.080 77.565 65.260 ;
        RECT 82.625 65.130 82.855 65.260 ;
        RECT 77.255 55.160 77.615 65.080 ;
        RECT 82.565 55.180 82.935 65.130 ;
        RECT 83.765 65.090 83.995 65.260 ;
        RECT 83.695 55.140 84.065 65.090 ;
        RECT 85.055 65.080 85.285 65.260 ;
        RECT 88.585 65.090 88.815 65.270 ;
        RECT 93.875 65.140 94.105 65.270 ;
        RECT 84.965 55.190 85.385 65.080 ;
        RECT 88.505 55.170 88.865 65.090 ;
        RECT 93.815 55.190 94.185 65.140 ;
        RECT 95.015 65.100 95.245 65.270 ;
        RECT 94.945 55.150 95.315 65.100 ;
        RECT 96.305 65.090 96.535 65.270 ;
        RECT 96.215 55.200 96.635 65.090 ;
        RECT 99.865 65.080 100.095 65.260 ;
        RECT 105.155 65.130 105.385 65.260 ;
        RECT 99.785 55.160 100.145 65.080 ;
        RECT 105.095 55.180 105.465 65.130 ;
        RECT 106.295 65.090 106.525 65.260 ;
        RECT 106.225 55.140 106.595 65.090 ;
        RECT 107.585 65.080 107.815 65.260 ;
        RECT 111.135 65.080 111.365 65.260 ;
        RECT 116.425 65.130 116.655 65.260 ;
        RECT 107.495 55.190 107.915 65.080 ;
        RECT 111.055 55.160 111.415 65.080 ;
        RECT 116.365 55.180 116.735 65.130 ;
        RECT 117.565 65.090 117.795 65.260 ;
        RECT 117.495 55.140 117.865 65.090 ;
        RECT 118.855 65.080 119.085 65.260 ;
        RECT 122.385 65.080 122.615 65.260 ;
        RECT 127.675 65.130 127.905 65.260 ;
        RECT 118.765 55.190 119.185 65.080 ;
        RECT 122.305 55.160 122.665 65.080 ;
        RECT 127.615 55.180 127.985 65.130 ;
        RECT 128.815 65.090 129.045 65.260 ;
        RECT 128.745 55.140 129.115 65.090 ;
        RECT 130.105 65.080 130.335 65.260 ;
        RECT 133.135 65.130 133.365 65.230 ;
        RECT 130.015 55.190 130.435 65.080 ;
        RECT 133.005 55.240 133.405 65.130 ;
        RECT 138.425 65.100 138.655 65.230 ;
        RECT 133.135 55.230 133.365 55.240 ;
        RECT 138.345 55.130 138.725 65.100 ;
        RECT 149.340 64.660 150.720 65.760 ;
        RECT 20.815 54.230 25.555 54.530 ;
        RECT 32.015 54.240 36.755 54.540 ;
        RECT 43.235 54.210 47.975 54.510 ;
        RECT 54.485 54.190 59.225 54.490 ;
        RECT 65.705 54.180 70.445 54.480 ;
        RECT 76.945 54.170 81.685 54.470 ;
        RECT 88.195 54.180 92.935 54.480 ;
        RECT 99.475 54.170 104.215 54.470 ;
        RECT 110.745 54.170 115.485 54.470 ;
        RECT 121.995 54.170 126.735 54.470 ;
        RECT 21.655 52.320 22.115 52.550 ;
        RECT 25.625 52.280 26.255 52.560 ;
        RECT 25.735 52.240 26.195 52.280 ;
        RECT 27.665 52.240 28.125 52.470 ;
        RECT 32.855 52.330 33.315 52.560 ;
        RECT 36.825 52.290 37.455 52.570 ;
        RECT 36.935 52.250 37.395 52.290 ;
        RECT 38.865 52.250 39.325 52.480 ;
        RECT 44.075 52.300 44.535 52.530 ;
        RECT 48.045 52.260 48.675 52.540 ;
        RECT 48.155 52.220 48.615 52.260 ;
        RECT 50.085 52.220 50.545 52.450 ;
        RECT 55.325 52.280 55.785 52.510 ;
        RECT 59.295 52.240 59.925 52.520 ;
        RECT 59.405 52.200 59.865 52.240 ;
        RECT 61.335 52.200 61.795 52.430 ;
        RECT 66.545 52.270 67.005 52.500 ;
        RECT 70.515 52.230 71.145 52.510 ;
        RECT 70.625 52.190 71.085 52.230 ;
        RECT 72.555 52.190 73.015 52.420 ;
        RECT 77.785 52.260 78.245 52.490 ;
        RECT 81.755 52.220 82.385 52.500 ;
        RECT 81.865 52.180 82.325 52.220 ;
        RECT 83.795 52.180 84.255 52.410 ;
        RECT 89.035 52.270 89.495 52.500 ;
        RECT 93.005 52.230 93.635 52.510 ;
        RECT 93.115 52.190 93.575 52.230 ;
        RECT 95.045 52.190 95.505 52.420 ;
        RECT 100.315 52.260 100.775 52.490 ;
        RECT 104.285 52.220 104.915 52.500 ;
        RECT 104.395 52.180 104.855 52.220 ;
        RECT 106.325 52.180 106.785 52.410 ;
        RECT 111.585 52.260 112.045 52.490 ;
        RECT 115.555 52.220 116.185 52.500 ;
        RECT 115.665 52.180 116.125 52.220 ;
        RECT 117.595 52.180 118.055 52.410 ;
        RECT 122.835 52.260 123.295 52.490 ;
        RECT 126.805 52.220 127.435 52.500 ;
        RECT 126.915 52.180 127.375 52.220 ;
        RECT 128.845 52.180 129.305 52.410 ;
        RECT 21.375 52.010 21.605 52.115 ;
        RECT 21.245 50.290 21.615 52.010 ;
        RECT 22.165 51.890 22.395 52.115 ;
        RECT 25.455 51.980 25.685 52.035 ;
        RECT 21.375 50.115 21.605 50.290 ;
        RECT 22.155 50.210 22.525 51.890 ;
        RECT 22.165 50.115 22.395 50.210 ;
        RECT 21.525 49.670 22.245 49.930 ;
        RECT 19.295 46.650 20.065 47.720 ;
        RECT 21.385 47.490 22.105 47.750 ;
        RECT 21.225 47.200 21.455 47.340 ;
        RECT 21.085 46.430 21.475 47.200 ;
        RECT 22.015 47.190 22.245 47.340 ;
        RECT 22.005 46.450 22.375 47.190 ;
        RECT 25.305 47.010 25.735 51.980 ;
        RECT 26.245 51.970 26.475 52.035 ;
        RECT 27.385 51.970 27.615 52.035 ;
        RECT 26.185 46.970 26.585 51.970 ;
        RECT 27.265 46.970 27.665 51.970 ;
        RECT 28.175 51.940 28.405 52.035 ;
        RECT 32.575 52.020 32.805 52.125 ;
        RECT 28.115 46.970 28.545 51.940 ;
        RECT 32.445 50.300 32.815 52.020 ;
        RECT 33.365 51.900 33.595 52.125 ;
        RECT 36.655 51.990 36.885 52.045 ;
        RECT 32.575 50.125 32.805 50.300 ;
        RECT 33.355 50.220 33.725 51.900 ;
        RECT 33.365 50.125 33.595 50.220 ;
        RECT 32.725 49.680 33.445 49.940 ;
        RECT 25.735 46.600 26.195 46.830 ;
        RECT 27.665 46.710 28.125 46.830 ;
        RECT 27.515 46.600 28.125 46.710 ;
        RECT 30.495 46.660 31.265 47.730 ;
        RECT 32.585 47.500 33.305 47.760 ;
        RECT 32.425 47.210 32.655 47.350 ;
        RECT 21.225 46.340 21.455 46.430 ;
        RECT 22.015 46.340 22.245 46.450 ;
        RECT 27.515 46.430 28.095 46.600 ;
        RECT 32.285 46.440 32.675 47.210 ;
        RECT 33.215 47.200 33.445 47.350 ;
        RECT 33.205 46.460 33.575 47.200 ;
        RECT 36.505 47.020 36.935 51.990 ;
        RECT 37.445 51.980 37.675 52.045 ;
        RECT 38.585 51.980 38.815 52.045 ;
        RECT 37.385 46.980 37.785 51.980 ;
        RECT 38.465 46.980 38.865 51.980 ;
        RECT 39.375 51.950 39.605 52.045 ;
        RECT 43.795 51.990 44.025 52.095 ;
        RECT 39.315 46.980 39.745 51.950 ;
        RECT 43.665 50.270 44.035 51.990 ;
        RECT 44.585 51.870 44.815 52.095 ;
        RECT 47.875 51.960 48.105 52.015 ;
        RECT 43.795 50.095 44.025 50.270 ;
        RECT 44.575 50.190 44.945 51.870 ;
        RECT 44.585 50.095 44.815 50.190 ;
        RECT 43.945 49.650 44.665 49.910 ;
        RECT 36.935 46.610 37.395 46.840 ;
        RECT 38.865 46.720 39.325 46.840 ;
        RECT 38.715 46.610 39.325 46.720 ;
        RECT 41.715 46.630 42.485 47.700 ;
        RECT 43.805 47.470 44.525 47.730 ;
        RECT 43.645 47.180 43.875 47.320 ;
        RECT 32.425 46.350 32.655 46.440 ;
        RECT 33.215 46.350 33.445 46.460 ;
        RECT 38.715 46.440 39.295 46.610 ;
        RECT 43.505 46.410 43.895 47.180 ;
        RECT 44.435 47.170 44.665 47.320 ;
        RECT 44.425 46.430 44.795 47.170 ;
        RECT 47.725 46.990 48.155 51.960 ;
        RECT 48.665 51.950 48.895 52.015 ;
        RECT 49.805 51.950 50.035 52.015 ;
        RECT 48.605 46.950 49.005 51.950 ;
        RECT 49.685 46.950 50.085 51.950 ;
        RECT 50.595 51.920 50.825 52.015 ;
        RECT 55.045 51.970 55.275 52.075 ;
        RECT 50.535 46.950 50.965 51.920 ;
        RECT 54.915 50.250 55.285 51.970 ;
        RECT 55.835 51.850 56.065 52.075 ;
        RECT 59.125 51.940 59.355 51.995 ;
        RECT 55.045 50.075 55.275 50.250 ;
        RECT 55.825 50.170 56.195 51.850 ;
        RECT 55.835 50.075 56.065 50.170 ;
        RECT 55.195 49.630 55.915 49.890 ;
        RECT 48.155 46.580 48.615 46.810 ;
        RECT 50.085 46.690 50.545 46.810 ;
        RECT 49.935 46.580 50.545 46.690 ;
        RECT 52.965 46.610 53.735 47.680 ;
        RECT 55.055 47.450 55.775 47.710 ;
        RECT 54.895 47.160 55.125 47.300 ;
        RECT 43.645 46.320 43.875 46.410 ;
        RECT 44.435 46.320 44.665 46.430 ;
        RECT 49.935 46.410 50.515 46.580 ;
        RECT 54.755 46.390 55.145 47.160 ;
        RECT 55.685 47.150 55.915 47.300 ;
        RECT 55.675 46.410 56.045 47.150 ;
        RECT 58.975 46.970 59.405 51.940 ;
        RECT 59.915 51.930 60.145 51.995 ;
        RECT 61.055 51.930 61.285 51.995 ;
        RECT 59.855 46.930 60.255 51.930 ;
        RECT 60.935 46.930 61.335 51.930 ;
        RECT 61.845 51.900 62.075 51.995 ;
        RECT 66.265 51.960 66.495 52.065 ;
        RECT 61.785 46.930 62.215 51.900 ;
        RECT 66.135 50.240 66.505 51.960 ;
        RECT 67.055 51.840 67.285 52.065 ;
        RECT 70.345 51.930 70.575 51.985 ;
        RECT 66.265 50.065 66.495 50.240 ;
        RECT 67.045 50.160 67.415 51.840 ;
        RECT 67.055 50.065 67.285 50.160 ;
        RECT 66.415 49.620 67.135 49.880 ;
        RECT 59.405 46.560 59.865 46.790 ;
        RECT 61.335 46.670 61.795 46.790 ;
        RECT 61.185 46.560 61.795 46.670 ;
        RECT 64.185 46.600 64.955 47.670 ;
        RECT 66.275 47.440 66.995 47.700 ;
        RECT 66.115 47.150 66.345 47.290 ;
        RECT 54.895 46.300 55.125 46.390 ;
        RECT 55.685 46.300 55.915 46.410 ;
        RECT 61.185 46.390 61.765 46.560 ;
        RECT 65.975 46.380 66.365 47.150 ;
        RECT 66.905 47.140 67.135 47.290 ;
        RECT 66.895 46.400 67.265 47.140 ;
        RECT 70.195 46.960 70.625 51.930 ;
        RECT 71.135 51.920 71.365 51.985 ;
        RECT 72.275 51.920 72.505 51.985 ;
        RECT 71.075 46.920 71.475 51.920 ;
        RECT 72.155 46.920 72.555 51.920 ;
        RECT 73.065 51.890 73.295 51.985 ;
        RECT 77.505 51.950 77.735 52.055 ;
        RECT 73.005 46.920 73.435 51.890 ;
        RECT 77.375 50.230 77.745 51.950 ;
        RECT 78.295 51.830 78.525 52.055 ;
        RECT 81.585 51.920 81.815 51.975 ;
        RECT 77.505 50.055 77.735 50.230 ;
        RECT 78.285 50.150 78.655 51.830 ;
        RECT 78.295 50.055 78.525 50.150 ;
        RECT 77.655 49.610 78.375 49.870 ;
        RECT 70.625 46.550 71.085 46.780 ;
        RECT 72.555 46.660 73.015 46.780 ;
        RECT 72.405 46.550 73.015 46.660 ;
        RECT 75.425 46.590 76.195 47.660 ;
        RECT 77.515 47.430 78.235 47.690 ;
        RECT 77.355 47.140 77.585 47.280 ;
        RECT 66.115 46.290 66.345 46.380 ;
        RECT 66.905 46.290 67.135 46.400 ;
        RECT 72.405 46.380 72.985 46.550 ;
        RECT 77.215 46.370 77.605 47.140 ;
        RECT 78.145 47.130 78.375 47.280 ;
        RECT 78.135 46.390 78.505 47.130 ;
        RECT 81.435 46.950 81.865 51.920 ;
        RECT 82.375 51.910 82.605 51.975 ;
        RECT 83.515 51.910 83.745 51.975 ;
        RECT 82.315 46.910 82.715 51.910 ;
        RECT 83.395 46.910 83.795 51.910 ;
        RECT 84.305 51.880 84.535 51.975 ;
        RECT 88.755 51.960 88.985 52.065 ;
        RECT 84.245 46.910 84.675 51.880 ;
        RECT 88.625 50.240 88.995 51.960 ;
        RECT 89.545 51.840 89.775 52.065 ;
        RECT 92.835 51.930 93.065 51.985 ;
        RECT 88.755 50.065 88.985 50.240 ;
        RECT 89.535 50.160 89.905 51.840 ;
        RECT 89.545 50.065 89.775 50.160 ;
        RECT 88.905 49.620 89.625 49.880 ;
        RECT 81.865 46.540 82.325 46.770 ;
        RECT 83.795 46.650 84.255 46.770 ;
        RECT 83.645 46.540 84.255 46.650 ;
        RECT 86.675 46.600 87.445 47.670 ;
        RECT 88.765 47.440 89.485 47.700 ;
        RECT 88.605 47.150 88.835 47.290 ;
        RECT 77.355 46.280 77.585 46.370 ;
        RECT 78.145 46.280 78.375 46.390 ;
        RECT 83.645 46.370 84.225 46.540 ;
        RECT 88.465 46.380 88.855 47.150 ;
        RECT 89.395 47.140 89.625 47.290 ;
        RECT 89.385 46.400 89.755 47.140 ;
        RECT 92.685 46.960 93.115 51.930 ;
        RECT 93.625 51.920 93.855 51.985 ;
        RECT 94.765 51.920 94.995 51.985 ;
        RECT 93.565 46.920 93.965 51.920 ;
        RECT 94.645 46.920 95.045 51.920 ;
        RECT 95.555 51.890 95.785 51.985 ;
        RECT 100.035 51.950 100.265 52.055 ;
        RECT 95.495 46.920 95.925 51.890 ;
        RECT 99.905 50.230 100.275 51.950 ;
        RECT 100.825 51.830 101.055 52.055 ;
        RECT 104.115 51.920 104.345 51.975 ;
        RECT 100.035 50.055 100.265 50.230 ;
        RECT 100.815 50.150 101.185 51.830 ;
        RECT 100.825 50.055 101.055 50.150 ;
        RECT 100.185 49.610 100.905 49.870 ;
        RECT 93.115 46.550 93.575 46.780 ;
        RECT 95.045 46.660 95.505 46.780 ;
        RECT 94.895 46.550 95.505 46.660 ;
        RECT 97.955 46.590 98.725 47.660 ;
        RECT 100.045 47.430 100.765 47.690 ;
        RECT 99.885 47.140 100.115 47.280 ;
        RECT 88.605 46.290 88.835 46.380 ;
        RECT 89.395 46.290 89.625 46.400 ;
        RECT 94.895 46.380 95.475 46.550 ;
        RECT 99.745 46.370 100.135 47.140 ;
        RECT 100.675 47.130 100.905 47.280 ;
        RECT 100.665 46.390 101.035 47.130 ;
        RECT 103.965 46.950 104.395 51.920 ;
        RECT 104.905 51.910 105.135 51.975 ;
        RECT 106.045 51.910 106.275 51.975 ;
        RECT 104.845 46.910 105.245 51.910 ;
        RECT 105.925 46.910 106.325 51.910 ;
        RECT 106.835 51.880 107.065 51.975 ;
        RECT 111.305 51.950 111.535 52.055 ;
        RECT 106.775 46.910 107.205 51.880 ;
        RECT 111.175 50.230 111.545 51.950 ;
        RECT 112.095 51.830 112.325 52.055 ;
        RECT 115.385 51.920 115.615 51.975 ;
        RECT 111.305 50.055 111.535 50.230 ;
        RECT 112.085 50.150 112.455 51.830 ;
        RECT 112.095 50.055 112.325 50.150 ;
        RECT 111.455 49.610 112.175 49.870 ;
        RECT 104.395 46.540 104.855 46.770 ;
        RECT 106.325 46.650 106.785 46.770 ;
        RECT 106.175 46.540 106.785 46.650 ;
        RECT 109.225 46.590 109.995 47.660 ;
        RECT 111.315 47.430 112.035 47.690 ;
        RECT 111.155 47.140 111.385 47.280 ;
        RECT 99.885 46.280 100.115 46.370 ;
        RECT 100.675 46.280 100.905 46.390 ;
        RECT 106.175 46.370 106.755 46.540 ;
        RECT 111.015 46.370 111.405 47.140 ;
        RECT 111.945 47.130 112.175 47.280 ;
        RECT 111.935 46.390 112.305 47.130 ;
        RECT 115.235 46.950 115.665 51.920 ;
        RECT 116.175 51.910 116.405 51.975 ;
        RECT 117.315 51.910 117.545 51.975 ;
        RECT 116.115 46.910 116.515 51.910 ;
        RECT 117.195 46.910 117.595 51.910 ;
        RECT 118.105 51.880 118.335 51.975 ;
        RECT 122.555 51.950 122.785 52.055 ;
        RECT 118.045 46.910 118.475 51.880 ;
        RECT 122.425 50.230 122.795 51.950 ;
        RECT 123.345 51.830 123.575 52.055 ;
        RECT 126.635 51.920 126.865 51.975 ;
        RECT 122.555 50.055 122.785 50.230 ;
        RECT 123.335 50.150 123.705 51.830 ;
        RECT 123.345 50.055 123.575 50.150 ;
        RECT 122.705 49.610 123.425 49.870 ;
        RECT 115.665 46.540 116.125 46.770 ;
        RECT 117.595 46.650 118.055 46.770 ;
        RECT 117.445 46.540 118.055 46.650 ;
        RECT 120.475 46.590 121.245 47.660 ;
        RECT 122.565 47.430 123.285 47.690 ;
        RECT 122.405 47.140 122.635 47.280 ;
        RECT 111.155 46.280 111.385 46.370 ;
        RECT 111.945 46.280 112.175 46.390 ;
        RECT 117.445 46.370 118.025 46.540 ;
        RECT 122.265 46.370 122.655 47.140 ;
        RECT 123.195 47.130 123.425 47.280 ;
        RECT 123.185 46.390 123.555 47.130 ;
        RECT 126.485 46.950 126.915 51.920 ;
        RECT 127.425 51.910 127.655 51.975 ;
        RECT 128.565 51.910 128.795 51.975 ;
        RECT 127.365 46.910 127.765 51.910 ;
        RECT 128.445 46.910 128.845 51.910 ;
        RECT 129.355 51.880 129.585 51.975 ;
        RECT 129.295 46.910 129.725 51.880 ;
        RECT 126.915 46.540 127.375 46.770 ;
        RECT 128.845 46.650 129.305 46.770 ;
        RECT 128.695 46.540 129.305 46.650 ;
        RECT 122.405 46.280 122.635 46.370 ;
        RECT 123.195 46.280 123.425 46.390 ;
        RECT 128.695 46.370 129.275 46.540 ;
        RECT 21.505 45.950 21.965 46.180 ;
        RECT 32.705 45.960 33.165 46.190 ;
        RECT 43.925 45.930 44.385 46.160 ;
        RECT 55.175 45.910 55.635 46.140 ;
        RECT 66.395 45.900 66.855 46.130 ;
        RECT 77.635 45.890 78.095 46.120 ;
        RECT 88.885 45.900 89.345 46.130 ;
        RECT 100.165 45.890 100.625 46.120 ;
        RECT 111.435 45.890 111.895 46.120 ;
        RECT 122.685 45.890 123.145 46.120 ;
        RECT 29.055 45.020 41.225 45.030 ;
        RECT 17.855 45.005 41.225 45.020 ;
        RECT 15.900 45.000 41.225 45.005 ;
        RECT 15.900 44.980 52.445 45.000 ;
        RECT 15.900 44.970 63.695 44.980 ;
        RECT 15.900 44.960 74.915 44.970 ;
        RECT 85.235 44.960 97.405 44.970 ;
        RECT 15.900 43.880 131.205 44.960 ;
        RECT 15.900 43.870 30.025 43.880 ;
        RECT 15.900 43.855 18.690 43.870 ;
        RECT 15.900 41.620 17.050 43.855 ;
        RECT 40.275 43.850 131.205 43.880 ;
        RECT 51.525 43.830 131.205 43.850 ;
        RECT 62.745 43.820 131.205 43.830 ;
        RECT 73.985 43.810 86.155 43.820 ;
        RECT 96.515 43.810 131.205 43.820 ;
        RECT 29.015 43.330 41.185 43.340 ;
        RECT 17.815 43.310 41.185 43.330 ;
        RECT 142.830 43.320 144.150 43.340 ;
        RECT 17.815 43.290 52.405 43.310 ;
        RECT 140.750 43.300 144.150 43.320 ;
        RECT 17.815 43.280 63.655 43.290 ;
        RECT 119.895 43.280 144.150 43.300 ;
        RECT 17.815 43.270 74.875 43.280 ;
        RECT 85.195 43.270 97.365 43.280 ;
        RECT 108.685 43.270 144.150 43.280 ;
        RECT 17.815 42.180 144.150 43.270 ;
        RECT 18.755 42.150 144.150 42.180 ;
        RECT 18.755 42.120 131.165 42.150 ;
        RECT 18.755 42.090 109.655 42.120 ;
        RECT 18.755 42.080 98.445 42.090 ;
        RECT 41.325 42.070 98.445 42.080 ;
        RECT 142.830 42.070 144.150 42.150 ;
        RECT 41.325 42.060 87.205 42.070 ;
        RECT 75.035 42.050 87.205 42.060 ;
        RECT 15.900 41.540 19.685 41.620 ;
        RECT 142.070 41.610 146.210 41.640 ;
        RECT 119.855 41.590 146.210 41.610 ;
        RECT 108.645 41.550 146.210 41.590 ;
        RECT 15.900 41.520 42.165 41.540 ;
        RECT 97.445 41.530 146.210 41.550 ;
        RECT 15.900 41.510 75.875 41.520 ;
        RECT 86.235 41.510 146.210 41.530 ;
        RECT 15.900 40.500 146.210 41.510 ;
        RECT 15.900 40.480 142.320 40.500 ;
        RECT 15.900 40.470 140.920 40.480 ;
        RECT 18.715 40.460 140.920 40.470 ;
        RECT 142.070 40.460 142.250 40.480 ;
        RECT 18.715 40.440 120.815 40.460 ;
        RECT 18.715 40.400 109.615 40.440 ;
        RECT 18.715 40.390 98.405 40.400 ;
        RECT 41.285 40.380 98.405 40.390 ;
        RECT 41.285 40.370 87.165 40.380 ;
        RECT 74.995 40.360 87.165 40.370 ;
        RECT 26.775 39.230 27.235 39.460 ;
        RECT 38.055 39.230 38.515 39.460 ;
        RECT 49.345 39.210 49.805 39.440 ;
        RECT 60.565 39.210 61.025 39.440 ;
        RECT 71.765 39.210 72.225 39.440 ;
        RECT 83.055 39.200 83.515 39.430 ;
        RECT 94.295 39.220 94.755 39.450 ;
        RECT 105.505 39.240 105.965 39.470 ;
        RECT 116.705 39.280 117.165 39.510 ;
        RECT 127.915 39.300 128.375 39.530 ;
        RECT 20.645 38.810 21.225 38.980 ;
        RECT 26.495 38.960 26.725 39.070 ;
        RECT 27.285 38.980 27.515 39.070 ;
        RECT 20.615 38.700 21.225 38.810 ;
        RECT 20.615 38.580 21.075 38.700 ;
        RECT 22.545 38.580 23.005 38.810 ;
        RECT 20.195 33.470 20.625 38.440 ;
        RECT 20.335 33.375 20.565 33.470 ;
        RECT 21.075 33.440 21.475 38.440 ;
        RECT 22.155 33.440 22.555 38.440 ;
        RECT 21.125 33.375 21.355 33.440 ;
        RECT 22.265 33.375 22.495 33.440 ;
        RECT 23.005 33.430 23.435 38.400 ;
        RECT 26.365 38.220 26.735 38.960 ;
        RECT 26.495 38.070 26.725 38.220 ;
        RECT 27.265 38.210 27.655 38.980 ;
        RECT 31.925 38.810 32.505 38.980 ;
        RECT 37.775 38.960 38.005 39.070 ;
        RECT 38.565 38.980 38.795 39.070 ;
        RECT 27.285 38.070 27.515 38.210 ;
        RECT 26.635 37.660 27.355 37.920 ;
        RECT 28.675 37.690 29.445 38.760 ;
        RECT 31.895 38.700 32.505 38.810 ;
        RECT 31.895 38.580 32.355 38.700 ;
        RECT 33.825 38.580 34.285 38.810 ;
        RECT 26.495 35.480 27.215 35.740 ;
        RECT 26.345 35.200 26.575 35.295 ;
        RECT 26.215 33.520 26.585 35.200 ;
        RECT 27.135 35.120 27.365 35.295 ;
        RECT 23.055 33.375 23.285 33.430 ;
        RECT 26.345 33.295 26.575 33.520 ;
        RECT 27.125 33.400 27.495 35.120 ;
        RECT 31.475 33.470 31.905 38.440 ;
        RECT 27.135 33.295 27.365 33.400 ;
        RECT 31.615 33.375 31.845 33.470 ;
        RECT 32.355 33.440 32.755 38.440 ;
        RECT 33.435 33.440 33.835 38.440 ;
        RECT 32.405 33.375 32.635 33.440 ;
        RECT 33.545 33.375 33.775 33.440 ;
        RECT 34.285 33.430 34.715 38.400 ;
        RECT 37.645 38.220 38.015 38.960 ;
        RECT 37.775 38.070 38.005 38.220 ;
        RECT 38.545 38.210 38.935 38.980 ;
        RECT 43.215 38.790 43.795 38.960 ;
        RECT 49.065 38.940 49.295 39.050 ;
        RECT 49.855 38.960 50.085 39.050 ;
        RECT 38.565 38.070 38.795 38.210 ;
        RECT 37.915 37.660 38.635 37.920 ;
        RECT 39.955 37.690 40.725 38.760 ;
        RECT 43.185 38.680 43.795 38.790 ;
        RECT 43.185 38.560 43.645 38.680 ;
        RECT 45.115 38.560 45.575 38.790 ;
        RECT 37.775 35.480 38.495 35.740 ;
        RECT 37.625 35.200 37.855 35.295 ;
        RECT 37.495 33.520 37.865 35.200 ;
        RECT 38.415 35.120 38.645 35.295 ;
        RECT 34.335 33.375 34.565 33.430 ;
        RECT 37.625 33.295 37.855 33.520 ;
        RECT 38.405 33.400 38.775 35.120 ;
        RECT 42.765 33.450 43.195 38.420 ;
        RECT 38.415 33.295 38.645 33.400 ;
        RECT 42.905 33.355 43.135 33.450 ;
        RECT 43.645 33.420 44.045 38.420 ;
        RECT 44.725 33.420 45.125 38.420 ;
        RECT 43.695 33.355 43.925 33.420 ;
        RECT 44.835 33.355 45.065 33.420 ;
        RECT 45.575 33.410 46.005 38.380 ;
        RECT 48.935 38.200 49.305 38.940 ;
        RECT 49.065 38.050 49.295 38.200 ;
        RECT 49.835 38.190 50.225 38.960 ;
        RECT 54.435 38.790 55.015 38.960 ;
        RECT 60.285 38.940 60.515 39.050 ;
        RECT 61.075 38.960 61.305 39.050 ;
        RECT 49.855 38.050 50.085 38.190 ;
        RECT 49.205 37.640 49.925 37.900 ;
        RECT 51.245 37.670 52.015 38.740 ;
        RECT 54.405 38.680 55.015 38.790 ;
        RECT 54.405 38.560 54.865 38.680 ;
        RECT 56.335 38.560 56.795 38.790 ;
        RECT 49.065 35.460 49.785 35.720 ;
        RECT 48.915 35.180 49.145 35.275 ;
        RECT 48.785 33.500 49.155 35.180 ;
        RECT 49.705 35.100 49.935 35.275 ;
        RECT 45.625 33.355 45.855 33.410 ;
        RECT 48.915 33.275 49.145 33.500 ;
        RECT 49.695 33.380 50.065 35.100 ;
        RECT 53.985 33.450 54.415 38.420 ;
        RECT 49.705 33.275 49.935 33.380 ;
        RECT 54.125 33.355 54.355 33.450 ;
        RECT 54.865 33.420 55.265 38.420 ;
        RECT 55.945 33.420 56.345 38.420 ;
        RECT 54.915 33.355 55.145 33.420 ;
        RECT 56.055 33.355 56.285 33.420 ;
        RECT 56.795 33.410 57.225 38.380 ;
        RECT 60.155 38.200 60.525 38.940 ;
        RECT 60.285 38.050 60.515 38.200 ;
        RECT 61.055 38.190 61.445 38.960 ;
        RECT 65.635 38.790 66.215 38.960 ;
        RECT 71.485 38.940 71.715 39.050 ;
        RECT 72.275 38.960 72.505 39.050 ;
        RECT 61.075 38.050 61.305 38.190 ;
        RECT 60.425 37.640 61.145 37.900 ;
        RECT 62.465 37.670 63.235 38.740 ;
        RECT 65.605 38.680 66.215 38.790 ;
        RECT 65.605 38.560 66.065 38.680 ;
        RECT 67.535 38.560 67.995 38.790 ;
        RECT 60.285 35.460 61.005 35.720 ;
        RECT 60.135 35.180 60.365 35.275 ;
        RECT 60.005 33.500 60.375 35.180 ;
        RECT 60.925 35.100 61.155 35.275 ;
        RECT 56.845 33.355 57.075 33.410 ;
        RECT 60.135 33.275 60.365 33.500 ;
        RECT 60.915 33.380 61.285 35.100 ;
        RECT 65.185 33.450 65.615 38.420 ;
        RECT 60.925 33.275 61.155 33.380 ;
        RECT 65.325 33.355 65.555 33.450 ;
        RECT 66.065 33.420 66.465 38.420 ;
        RECT 67.145 33.420 67.545 38.420 ;
        RECT 66.115 33.355 66.345 33.420 ;
        RECT 67.255 33.355 67.485 33.420 ;
        RECT 67.995 33.410 68.425 38.380 ;
        RECT 71.355 38.200 71.725 38.940 ;
        RECT 71.485 38.050 71.715 38.200 ;
        RECT 72.255 38.190 72.645 38.960 ;
        RECT 76.925 38.780 77.505 38.950 ;
        RECT 82.775 38.930 83.005 39.040 ;
        RECT 83.565 38.950 83.795 39.040 ;
        RECT 72.275 38.050 72.505 38.190 ;
        RECT 71.625 37.640 72.345 37.900 ;
        RECT 73.665 37.670 74.435 38.740 ;
        RECT 76.895 38.670 77.505 38.780 ;
        RECT 76.895 38.550 77.355 38.670 ;
        RECT 78.825 38.550 79.285 38.780 ;
        RECT 71.485 35.460 72.205 35.720 ;
        RECT 71.335 35.180 71.565 35.275 ;
        RECT 71.205 33.500 71.575 35.180 ;
        RECT 72.125 35.100 72.355 35.275 ;
        RECT 68.045 33.355 68.275 33.410 ;
        RECT 71.335 33.275 71.565 33.500 ;
        RECT 72.115 33.380 72.485 35.100 ;
        RECT 76.475 33.440 76.905 38.410 ;
        RECT 72.125 33.275 72.355 33.380 ;
        RECT 76.615 33.345 76.845 33.440 ;
        RECT 77.355 33.410 77.755 38.410 ;
        RECT 78.435 33.410 78.835 38.410 ;
        RECT 77.405 33.345 77.635 33.410 ;
        RECT 78.545 33.345 78.775 33.410 ;
        RECT 79.285 33.400 79.715 38.370 ;
        RECT 82.645 38.190 83.015 38.930 ;
        RECT 82.775 38.040 83.005 38.190 ;
        RECT 83.545 38.180 83.935 38.950 ;
        RECT 88.165 38.800 88.745 38.970 ;
        RECT 94.015 38.950 94.245 39.060 ;
        RECT 94.805 38.970 95.035 39.060 ;
        RECT 83.565 38.040 83.795 38.180 ;
        RECT 82.915 37.630 83.635 37.890 ;
        RECT 84.955 37.660 85.725 38.730 ;
        RECT 88.135 38.690 88.745 38.800 ;
        RECT 88.135 38.570 88.595 38.690 ;
        RECT 90.065 38.570 90.525 38.800 ;
        RECT 82.775 35.450 83.495 35.710 ;
        RECT 82.625 35.170 82.855 35.265 ;
        RECT 82.495 33.490 82.865 35.170 ;
        RECT 83.415 35.090 83.645 35.265 ;
        RECT 79.335 33.345 79.565 33.400 ;
        RECT 82.625 33.265 82.855 33.490 ;
        RECT 83.405 33.370 83.775 35.090 ;
        RECT 87.715 33.460 88.145 38.430 ;
        RECT 83.415 33.265 83.645 33.370 ;
        RECT 87.855 33.365 88.085 33.460 ;
        RECT 88.595 33.430 88.995 38.430 ;
        RECT 89.675 33.430 90.075 38.430 ;
        RECT 88.645 33.365 88.875 33.430 ;
        RECT 89.785 33.365 90.015 33.430 ;
        RECT 90.525 33.420 90.955 38.390 ;
        RECT 93.885 38.210 94.255 38.950 ;
        RECT 94.015 38.060 94.245 38.210 ;
        RECT 94.785 38.200 95.175 38.970 ;
        RECT 99.375 38.820 99.955 38.990 ;
        RECT 105.225 38.970 105.455 39.080 ;
        RECT 106.015 38.990 106.245 39.080 ;
        RECT 94.805 38.060 95.035 38.200 ;
        RECT 94.155 37.650 94.875 37.910 ;
        RECT 96.195 37.680 96.965 38.750 ;
        RECT 99.345 38.710 99.955 38.820 ;
        RECT 99.345 38.590 99.805 38.710 ;
        RECT 101.275 38.590 101.735 38.820 ;
        RECT 94.015 35.470 94.735 35.730 ;
        RECT 93.865 35.190 94.095 35.285 ;
        RECT 93.735 33.510 94.105 35.190 ;
        RECT 94.655 35.110 94.885 35.285 ;
        RECT 90.575 33.365 90.805 33.420 ;
        RECT 93.865 33.285 94.095 33.510 ;
        RECT 94.645 33.390 95.015 35.110 ;
        RECT 98.925 33.480 99.355 38.450 ;
        RECT 94.655 33.285 94.885 33.390 ;
        RECT 99.065 33.385 99.295 33.480 ;
        RECT 99.805 33.450 100.205 38.450 ;
        RECT 100.885 33.450 101.285 38.450 ;
        RECT 99.855 33.385 100.085 33.450 ;
        RECT 100.995 33.385 101.225 33.450 ;
        RECT 101.735 33.440 102.165 38.410 ;
        RECT 105.095 38.230 105.465 38.970 ;
        RECT 105.225 38.080 105.455 38.230 ;
        RECT 105.995 38.220 106.385 38.990 ;
        RECT 110.575 38.860 111.155 39.030 ;
        RECT 116.425 39.010 116.655 39.120 ;
        RECT 117.215 39.030 117.445 39.120 ;
        RECT 106.015 38.080 106.245 38.220 ;
        RECT 105.365 37.670 106.085 37.930 ;
        RECT 107.405 37.700 108.175 38.770 ;
        RECT 110.545 38.750 111.155 38.860 ;
        RECT 110.545 38.630 111.005 38.750 ;
        RECT 112.475 38.630 112.935 38.860 ;
        RECT 105.225 35.490 105.945 35.750 ;
        RECT 105.075 35.210 105.305 35.305 ;
        RECT 104.945 33.530 105.315 35.210 ;
        RECT 105.865 35.130 106.095 35.305 ;
        RECT 101.785 33.385 102.015 33.440 ;
        RECT 105.075 33.305 105.305 33.530 ;
        RECT 105.855 33.410 106.225 35.130 ;
        RECT 110.125 33.520 110.555 38.490 ;
        RECT 110.265 33.425 110.495 33.520 ;
        RECT 111.005 33.490 111.405 38.490 ;
        RECT 112.085 33.490 112.485 38.490 ;
        RECT 111.055 33.425 111.285 33.490 ;
        RECT 112.195 33.425 112.425 33.490 ;
        RECT 112.935 33.480 113.365 38.450 ;
        RECT 116.295 38.270 116.665 39.010 ;
        RECT 116.425 38.120 116.655 38.270 ;
        RECT 117.195 38.260 117.585 39.030 ;
        RECT 121.785 38.880 122.365 39.050 ;
        RECT 127.635 39.030 127.865 39.140 ;
        RECT 128.425 39.050 128.655 39.140 ;
        RECT 117.215 38.120 117.445 38.260 ;
        RECT 116.565 37.710 117.285 37.970 ;
        RECT 118.605 37.740 119.375 38.810 ;
        RECT 121.755 38.770 122.365 38.880 ;
        RECT 121.755 38.650 122.215 38.770 ;
        RECT 123.685 38.650 124.145 38.880 ;
        RECT 116.425 35.530 117.145 35.790 ;
        RECT 116.275 35.250 116.505 35.345 ;
        RECT 116.145 33.570 116.515 35.250 ;
        RECT 117.065 35.170 117.295 35.345 ;
        RECT 112.985 33.425 113.215 33.480 ;
        RECT 105.865 33.305 106.095 33.410 ;
        RECT 116.275 33.345 116.505 33.570 ;
        RECT 117.055 33.450 117.425 35.170 ;
        RECT 121.335 33.540 121.765 38.510 ;
        RECT 117.065 33.345 117.295 33.450 ;
        RECT 121.475 33.445 121.705 33.540 ;
        RECT 122.215 33.510 122.615 38.510 ;
        RECT 123.295 33.510 123.695 38.510 ;
        RECT 122.265 33.445 122.495 33.510 ;
        RECT 123.405 33.445 123.635 33.510 ;
        RECT 124.145 33.500 124.575 38.470 ;
        RECT 127.505 38.290 127.875 39.030 ;
        RECT 127.635 38.140 127.865 38.290 ;
        RECT 128.405 38.280 128.795 39.050 ;
        RECT 128.425 38.140 128.655 38.280 ;
        RECT 127.775 37.730 128.495 37.990 ;
        RECT 129.815 37.760 130.585 38.830 ;
        RECT 142.850 37.630 144.170 38.900 ;
        RECT 127.635 35.550 128.355 35.810 ;
        RECT 127.485 35.270 127.715 35.365 ;
        RECT 127.355 33.590 127.725 35.270 ;
        RECT 128.275 35.190 128.505 35.365 ;
        RECT 124.195 33.445 124.425 33.500 ;
        RECT 127.485 33.365 127.715 33.590 ;
        RECT 128.265 33.470 128.635 35.190 ;
        RECT 128.275 33.365 128.505 33.470 ;
        RECT 20.615 32.940 21.075 33.170 ;
        RECT 22.545 33.130 23.005 33.170 ;
        RECT 22.485 32.850 23.115 33.130 ;
        RECT 26.625 32.860 27.085 33.090 ;
        RECT 31.895 32.940 32.355 33.170 ;
        RECT 33.825 33.130 34.285 33.170 ;
        RECT 33.765 32.850 34.395 33.130 ;
        RECT 37.905 32.860 38.365 33.090 ;
        RECT 43.185 32.920 43.645 33.150 ;
        RECT 45.115 33.110 45.575 33.150 ;
        RECT 45.055 32.830 45.685 33.110 ;
        RECT 49.195 32.840 49.655 33.070 ;
        RECT 54.405 32.920 54.865 33.150 ;
        RECT 56.335 33.110 56.795 33.150 ;
        RECT 56.275 32.830 56.905 33.110 ;
        RECT 60.415 32.840 60.875 33.070 ;
        RECT 65.605 32.920 66.065 33.150 ;
        RECT 67.535 33.110 67.995 33.150 ;
        RECT 67.475 32.830 68.105 33.110 ;
        RECT 71.615 32.840 72.075 33.070 ;
        RECT 76.895 32.910 77.355 33.140 ;
        RECT 78.825 33.100 79.285 33.140 ;
        RECT 78.765 32.820 79.395 33.100 ;
        RECT 82.905 32.830 83.365 33.060 ;
        RECT 88.135 32.930 88.595 33.160 ;
        RECT 90.065 33.120 90.525 33.160 ;
        RECT 90.005 32.840 90.635 33.120 ;
        RECT 94.145 32.850 94.605 33.080 ;
        RECT 99.345 32.950 99.805 33.180 ;
        RECT 101.275 33.140 101.735 33.180 ;
        RECT 101.215 32.860 101.845 33.140 ;
        RECT 105.355 32.870 105.815 33.100 ;
        RECT 110.545 32.990 111.005 33.220 ;
        RECT 112.475 33.180 112.935 33.220 ;
        RECT 112.415 32.900 113.045 33.180 ;
        RECT 116.555 32.910 117.015 33.140 ;
        RECT 121.755 33.010 122.215 33.240 ;
        RECT 123.685 33.200 124.145 33.240 ;
        RECT 123.625 32.920 124.255 33.200 ;
        RECT 127.765 32.930 128.225 33.160 ;
        RECT 23.185 30.880 27.925 31.180 ;
        RECT 34.465 30.880 39.205 31.180 ;
        RECT 45.755 30.860 50.495 31.160 ;
        RECT 56.975 30.860 61.715 31.160 ;
        RECT 68.175 30.860 72.915 31.160 ;
        RECT 79.465 30.850 84.205 31.150 ;
        RECT 90.705 30.870 95.445 31.170 ;
        RECT 101.915 30.890 106.655 31.190 ;
        RECT 113.115 30.930 117.855 31.230 ;
        RECT 124.325 30.950 129.065 31.250 ;
        RECT 19.485 20.270 19.905 30.160 ;
        RECT 19.585 20.090 19.815 20.270 ;
        RECT 20.805 20.260 21.175 30.210 ;
        RECT 20.875 20.090 21.105 20.260 ;
        RECT 21.935 20.220 22.305 30.170 ;
        RECT 27.255 20.270 27.615 30.190 ;
        RECT 30.765 20.270 31.185 30.160 ;
        RECT 22.015 20.090 22.245 20.220 ;
        RECT 27.305 20.090 27.535 20.270 ;
        RECT 30.865 20.090 31.095 20.270 ;
        RECT 32.085 20.260 32.455 30.210 ;
        RECT 32.155 20.090 32.385 20.260 ;
        RECT 33.215 20.220 33.585 30.170 ;
        RECT 38.535 20.270 38.895 30.190 ;
        RECT 33.295 20.090 33.525 20.220 ;
        RECT 38.585 20.090 38.815 20.270 ;
        RECT 42.055 20.250 42.475 30.140 ;
        RECT 42.155 20.070 42.385 20.250 ;
        RECT 43.375 20.240 43.745 30.190 ;
        RECT 43.445 20.070 43.675 20.240 ;
        RECT 44.505 20.200 44.875 30.150 ;
        RECT 49.825 20.250 50.185 30.170 ;
        RECT 53.275 20.250 53.695 30.140 ;
        RECT 44.585 20.070 44.815 20.200 ;
        RECT 49.875 20.070 50.105 20.250 ;
        RECT 53.375 20.070 53.605 20.250 ;
        RECT 54.595 20.240 54.965 30.190 ;
        RECT 54.665 20.070 54.895 20.240 ;
        RECT 55.725 20.200 56.095 30.150 ;
        RECT 61.045 20.250 61.405 30.170 ;
        RECT 64.475 20.250 64.895 30.140 ;
        RECT 55.805 20.070 56.035 20.200 ;
        RECT 61.095 20.070 61.325 20.250 ;
        RECT 64.575 20.070 64.805 20.250 ;
        RECT 65.795 20.240 66.165 30.190 ;
        RECT 65.865 20.070 66.095 20.240 ;
        RECT 66.925 20.200 67.295 30.150 ;
        RECT 72.245 20.250 72.605 30.170 ;
        RECT 67.005 20.070 67.235 20.200 ;
        RECT 72.295 20.070 72.525 20.250 ;
        RECT 75.765 20.240 76.185 30.130 ;
        RECT 75.865 20.060 76.095 20.240 ;
        RECT 77.085 20.230 77.455 30.180 ;
        RECT 77.155 20.060 77.385 20.230 ;
        RECT 78.215 20.190 78.585 30.140 ;
        RECT 83.535 20.240 83.895 30.160 ;
        RECT 87.005 20.260 87.425 30.150 ;
        RECT 78.295 20.060 78.525 20.190 ;
        RECT 83.585 20.060 83.815 20.240 ;
        RECT 87.105 20.080 87.335 20.260 ;
        RECT 88.325 20.250 88.695 30.200 ;
        RECT 88.395 20.080 88.625 20.250 ;
        RECT 89.455 20.210 89.825 30.160 ;
        RECT 94.775 20.260 95.135 30.180 ;
        RECT 98.215 20.280 98.635 30.170 ;
        RECT 89.535 20.080 89.765 20.210 ;
        RECT 94.825 20.080 95.055 20.260 ;
        RECT 98.315 20.100 98.545 20.280 ;
        RECT 99.535 20.270 99.905 30.220 ;
        RECT 99.605 20.100 99.835 20.270 ;
        RECT 100.665 20.230 101.035 30.180 ;
        RECT 105.985 20.280 106.345 30.200 ;
        RECT 109.415 20.320 109.835 30.210 ;
        RECT 100.745 20.100 100.975 20.230 ;
        RECT 106.035 20.100 106.265 20.280 ;
        RECT 109.515 20.140 109.745 20.320 ;
        RECT 110.735 20.310 111.105 30.260 ;
        RECT 110.805 20.140 111.035 20.310 ;
        RECT 111.865 20.270 112.235 30.220 ;
        RECT 117.185 20.320 117.545 30.240 ;
        RECT 120.625 20.340 121.045 30.230 ;
        RECT 111.945 20.140 112.175 20.270 ;
        RECT 117.235 20.140 117.465 20.320 ;
        RECT 120.725 20.160 120.955 20.340 ;
        RECT 121.945 20.330 122.315 30.280 ;
        RECT 122.015 20.160 122.245 20.330 ;
        RECT 123.075 20.290 123.445 30.240 ;
        RECT 128.395 20.340 128.755 30.260 ;
        RECT 123.155 20.160 123.385 20.290 ;
        RECT 128.445 20.160 128.675 20.340 ;
        RECT 132.345 20.170 132.755 30.180 ;
        RECT 137.735 30.120 137.965 30.130 ;
        RECT 132.445 20.130 132.675 20.170 ;
        RECT 137.665 20.080 138.055 30.120 ;
        RECT 19.775 19.610 20.925 19.920 ;
        RECT 22.185 19.620 27.335 19.900 ;
        RECT 31.055 19.610 32.205 19.920 ;
        RECT 33.465 19.620 38.615 19.900 ;
        RECT 42.345 19.590 43.495 19.900 ;
        RECT 44.755 19.600 49.905 19.880 ;
        RECT 53.565 19.590 54.715 19.900 ;
        RECT 55.975 19.600 61.125 19.880 ;
        RECT 64.765 19.590 65.915 19.900 ;
        RECT 67.175 19.600 72.325 19.880 ;
        RECT 76.055 19.580 77.205 19.890 ;
        RECT 78.465 19.590 83.615 19.870 ;
        RECT 87.295 19.600 88.445 19.910 ;
        RECT 89.705 19.610 94.855 19.890 ;
        RECT 98.505 19.620 99.655 19.930 ;
        RECT 100.915 19.630 106.065 19.910 ;
        RECT 109.705 19.660 110.855 19.970 ;
        RECT 112.115 19.670 117.265 19.950 ;
        RECT 120.915 19.680 122.065 19.990 ;
        RECT 123.325 19.690 128.475 19.970 ;
        RECT 132.635 19.640 138.025 19.930 ;
        RECT 142.940 19.110 144.080 37.630 ;
        RECT 13.940 18.460 17.635 18.530 ;
        RECT 117.755 18.510 131.425 18.530 ;
        RECT 106.545 18.470 131.425 18.510 ;
        RECT 13.940 18.440 41.565 18.460 ;
        RECT 95.345 18.450 131.425 18.470 ;
        RECT 13.940 18.430 75.275 18.440 ;
        RECT 84.135 18.430 131.425 18.450 ;
        RECT 13.940 17.380 131.425 18.430 ;
        RECT 142.890 17.990 144.140 19.110 ;
        RECT 145.070 18.880 146.210 40.500 ;
        RECT 145.030 17.960 146.250 18.880 ;
        RECT 13.950 17.370 15.100 17.380 ;
        RECT 16.615 17.360 120.215 17.380 ;
        RECT 16.615 17.320 109.015 17.360 ;
        RECT 16.615 17.310 97.805 17.320 ;
        RECT 39.185 17.300 97.805 17.310 ;
        RECT 39.185 17.290 86.565 17.300 ;
        RECT 72.895 17.280 86.565 17.290 ;
        RECT 117.765 16.950 140.620 16.960 ;
        RECT 142.040 16.950 148.010 16.980 ;
        RECT 117.765 16.940 148.010 16.950 ;
        RECT 106.555 16.900 148.010 16.940 ;
        RECT 16.625 16.870 41.575 16.890 ;
        RECT 95.355 16.880 148.010 16.900 ;
        RECT 16.625 16.860 75.285 16.870 ;
        RECT 84.145 16.860 148.010 16.880 ;
        RECT 16.625 15.840 148.010 16.860 ;
        RECT 16.625 15.820 142.660 15.840 ;
        RECT 16.625 15.810 140.620 15.820 ;
        RECT 142.040 15.810 142.660 15.820 ;
        RECT 16.625 15.790 120.225 15.810 ;
        RECT 16.625 15.750 109.025 15.790 ;
        RECT 16.625 15.740 97.815 15.750 ;
        RECT 39.195 15.730 97.815 15.740 ;
        RECT 39.195 15.720 86.575 15.730 ;
        RECT 72.905 15.710 86.575 15.720 ;
        RECT 131.215 15.460 132.585 15.470 ;
        RECT 12.290 15.390 17.625 15.450 ;
        RECT 117.795 15.440 132.785 15.460 ;
        RECT 106.585 15.400 132.785 15.440 ;
        RECT 12.290 15.370 41.585 15.390 ;
        RECT 95.385 15.380 132.785 15.400 ;
        RECT 12.290 15.360 75.295 15.370 ;
        RECT 84.175 15.360 132.785 15.380 ;
        RECT 12.290 14.320 132.785 15.360 ;
        RECT 142.905 15.040 144.045 15.050 ;
        RECT 12.290 14.310 131.445 14.320 ;
        RECT 12.290 14.300 120.235 14.310 ;
        RECT 12.320 14.280 13.470 14.300 ;
        RECT 16.655 14.290 120.235 14.300 ;
        RECT 16.655 14.250 109.035 14.290 ;
        RECT 16.655 14.240 97.825 14.250 ;
        RECT 39.225 14.230 97.825 14.240 ;
        RECT 39.225 14.220 86.585 14.230 ;
        RECT 72.935 14.210 86.585 14.220 ;
        RECT 142.850 13.920 144.100 15.040 ;
        RECT 145.020 14.870 146.160 14.980 ;
        RECT 144.980 13.950 146.200 14.870 ;
        RECT 16.965 13.800 17.435 13.810 ;
        RECT 10.800 13.780 17.435 13.800 ;
        RECT 10.800 13.720 17.555 13.780 ;
        RECT 117.845 13.770 131.445 13.790 ;
        RECT 106.635 13.730 131.445 13.770 ;
        RECT 10.800 13.700 41.585 13.720 ;
        RECT 95.435 13.710 131.445 13.730 ;
        RECT 10.800 13.690 75.295 13.700 ;
        RECT 84.225 13.690 131.445 13.710 ;
        RECT 10.800 12.650 131.445 13.690 ;
        RECT 16.705 12.640 131.445 12.650 ;
        RECT 16.705 12.620 120.235 12.640 ;
        RECT 16.705 12.580 109.035 12.620 ;
        RECT 16.705 12.570 97.825 12.580 ;
        RECT 39.275 12.560 97.825 12.570 ;
        RECT 39.275 12.550 86.585 12.560 ;
        RECT 72.985 12.540 86.585 12.550 ;
        RECT 128.755 12.240 130.465 12.250 ;
        RECT 117.545 12.220 119.255 12.230 ;
        RECT 106.345 12.180 108.055 12.190 ;
        RECT 27.615 12.170 29.325 12.180 ;
        RECT 38.895 12.170 40.605 12.180 ;
        RECT 25.675 11.030 29.325 12.170 ;
        RECT 36.955 11.030 40.605 12.170 ;
        RECT 95.135 12.160 96.845 12.170 ;
        RECT 50.185 12.150 51.895 12.160 ;
        RECT 61.405 12.150 63.115 12.160 ;
        RECT 72.605 12.150 74.315 12.160 ;
        RECT 25.675 11.020 27.625 11.030 ;
        RECT 36.955 11.020 38.905 11.030 ;
        RECT 48.245 11.010 51.895 12.150 ;
        RECT 59.465 11.010 63.115 12.150 ;
        RECT 70.665 11.010 74.315 12.150 ;
        RECT 83.895 12.140 85.605 12.150 ;
        RECT 48.245 11.000 50.195 11.010 ;
        RECT 59.465 11.000 61.415 11.010 ;
        RECT 70.665 11.000 72.615 11.010 ;
        RECT 81.955 11.000 85.605 12.140 ;
        RECT 93.195 11.020 96.845 12.160 ;
        RECT 104.405 11.040 108.055 12.180 ;
        RECT 115.605 11.080 119.255 12.220 ;
        RECT 126.815 11.100 130.465 12.240 ;
        RECT 126.815 11.090 128.765 11.100 ;
        RECT 115.605 11.070 117.555 11.080 ;
        RECT 104.405 11.030 106.355 11.040 ;
        RECT 93.195 11.010 95.145 11.020 ;
        RECT 81.955 10.990 83.905 11.000 ;
        RECT 142.905 8.580 144.045 13.920 ;
        RECT 74.420 7.440 144.045 8.580 ;
        RECT 74.420 1.410 75.560 7.440 ;
        RECT 145.020 6.630 146.160 13.950 ;
        RECT 93.650 5.490 146.160 6.630 ;
        RECT 93.650 1.480 94.790 5.490 ;
        RECT 146.870 4.560 148.010 15.840 ;
        RECT 113.130 3.420 148.010 4.560 ;
        RECT 113.130 1.610 114.270 3.420 ;
        RECT 149.460 2.770 150.600 64.660 ;
        RECT 131.940 1.880 150.600 2.770 ;
        RECT 131.800 1.630 150.600 1.880 ;
        RECT 74.290 0.160 75.680 1.410 ;
        RECT 93.500 0.230 94.890 1.480 ;
        RECT 112.900 0.360 114.290 1.610 ;
        RECT 131.800 1.380 133.490 1.630 ;
        RECT 151.730 1.420 152.870 66.900 ;
        RECT 131.800 0.430 133.540 1.380 ;
        RECT 113.130 0.330 114.270 0.360 ;
        RECT 151.600 0.300 152.970 1.420 ;
        RECT 93.650 0.150 94.790 0.230 ;
      LAYER met2 ;
        RECT 135.390 223.830 136.740 225.230 ;
        RECT 138.180 223.760 139.530 225.160 ;
        RECT 143.230 223.790 144.580 225.190 ;
        RECT 47.235 194.340 47.515 196.340 ;
        RECT 63.335 194.340 63.615 196.340 ;
        RECT 76.215 194.340 76.495 196.340 ;
        RECT 79.435 194.340 79.715 196.340 ;
        RECT 82.655 194.340 82.935 196.340 ;
        RECT 105.195 194.340 105.475 196.340 ;
        RECT 20.105 192.270 20.365 192.590 ;
        RECT 36.205 192.270 36.465 192.590 ;
        RECT 39.425 192.270 39.685 192.590 ;
        RECT 40.805 192.270 41.065 192.590 ;
        RECT 17.635 190.715 19.175 191.085 ;
        RECT 17.635 185.275 19.175 185.645 ;
        RECT 20.165 182.610 20.305 192.270 ;
        RECT 30.685 191.250 30.945 191.570 ;
        RECT 30.745 189.190 30.885 191.250 ;
        RECT 36.265 189.530 36.405 192.270 ;
        RECT 38.965 191.250 39.225 191.570 ;
        RECT 36.205 189.210 36.465 189.530 ;
        RECT 39.025 189.190 39.165 191.250 ;
        RECT 30.685 188.870 30.945 189.190 ;
        RECT 32.525 188.870 32.785 189.190 ;
        RECT 38.965 188.870 39.225 189.190 ;
        RECT 25.625 188.530 25.885 188.850 ;
        RECT 25.685 184.770 25.825 188.530 ;
        RECT 29.305 187.170 29.565 187.490 ;
        RECT 28.385 186.490 28.645 186.810 ;
        RECT 27.925 185.810 28.185 186.130 ;
        RECT 26.085 184.790 26.345 185.110 ;
        RECT 25.625 184.450 25.885 184.770 ;
        RECT 21.025 183.430 21.285 183.750 ;
        RECT 20.165 182.470 20.765 182.610 ;
        RECT 20.625 181.710 20.765 182.470 ;
        RECT 20.565 181.390 20.825 181.710 ;
        RECT 17.635 179.835 19.175 180.205 ;
        RECT 20.095 178.815 20.375 179.185 ;
        RECT 20.105 178.670 20.365 178.815 ;
        RECT 20.625 176.610 20.765 181.390 ;
        RECT 21.085 177.970 21.225 183.430 ;
        RECT 21.485 180.710 21.745 181.030 ;
        RECT 21.545 178.650 21.685 180.710 ;
        RECT 21.945 179.350 22.205 179.670 ;
        RECT 21.485 178.330 21.745 178.650 ;
        RECT 21.025 177.650 21.285 177.970 ;
        RECT 21.485 177.650 21.745 177.970 ;
        RECT 20.565 176.290 20.825 176.610 ;
        RECT 20.565 175.610 20.825 175.930 ;
        RECT 17.635 174.395 19.175 174.765 ;
        RECT 17.635 168.955 19.175 169.325 ;
        RECT 19.645 167.110 19.905 167.430 ;
        RECT 19.705 165.585 19.845 167.110 ;
        RECT 20.625 165.730 20.765 175.610 ;
        RECT 21.545 173.550 21.685 177.650 ;
        RECT 21.485 173.230 21.745 173.550 ;
        RECT 22.005 170.830 22.145 179.350 ;
        RECT 26.145 178.990 26.285 184.790 ;
        RECT 27.985 179.330 28.125 185.810 ;
        RECT 28.445 184.090 28.585 186.490 ;
        RECT 29.365 185.110 29.505 187.170 ;
        RECT 31.145 185.810 31.405 186.130 ;
        RECT 29.305 184.790 29.565 185.110 ;
        RECT 30.685 184.790 30.945 185.110 ;
        RECT 30.745 184.090 30.885 184.790 ;
        RECT 28.385 183.770 28.645 184.090 ;
        RECT 30.685 183.770 30.945 184.090 ;
        RECT 27.925 179.010 28.185 179.330 ;
        RECT 26.085 178.670 26.345 178.990 ;
        RECT 22.405 178.330 22.665 178.650 ;
        RECT 22.465 176.950 22.605 178.330 ;
        RECT 23.315 178.135 23.595 178.505 ;
        RECT 22.405 176.630 22.665 176.950 ;
        RECT 22.405 175.950 22.665 176.270 ;
        RECT 22.465 173.210 22.605 175.950 ;
        RECT 22.405 172.890 22.665 173.210 ;
        RECT 21.945 170.510 22.205 170.830 ;
        RECT 21.485 169.665 21.745 169.810 ;
        RECT 21.475 169.295 21.755 169.665 ;
        RECT 19.635 165.215 19.915 165.585 ;
        RECT 20.565 165.410 20.825 165.730 ;
        RECT 17.635 163.515 19.175 163.885 ;
        RECT 22.005 162.330 22.145 170.510 ;
        RECT 21.945 162.010 22.205 162.330 ;
        RECT 22.465 161.390 22.605 172.890 ;
        RECT 22.865 172.210 23.125 172.530 ;
        RECT 22.925 167.770 23.065 172.210 ;
        RECT 23.385 170.830 23.525 178.135 ;
        RECT 24.235 176.095 24.515 176.465 ;
        RECT 23.325 170.510 23.585 170.830 ;
        RECT 22.865 167.450 23.125 167.770 ;
        RECT 23.385 165.730 23.525 170.510 ;
        RECT 23.785 165.750 24.045 166.070 ;
        RECT 23.325 165.410 23.585 165.730 ;
        RECT 23.845 165.585 23.985 165.750 ;
        RECT 24.305 165.730 24.445 176.095 ;
        RECT 24.705 174.930 24.965 175.250 ;
        RECT 23.775 165.215 24.055 165.585 ;
        RECT 24.245 165.410 24.505 165.730 ;
        RECT 21.545 161.250 22.605 161.390 ;
        RECT 21.545 159.950 21.685 161.250 ;
        RECT 21.485 159.630 21.745 159.950 ;
        RECT 22.395 159.775 22.675 160.145 ;
        RECT 22.405 159.630 22.665 159.775 ;
        RECT 17.635 158.075 19.175 158.445 ;
        RECT 21.545 155.190 21.685 159.630 ;
        RECT 21.485 154.870 21.745 155.190 ;
        RECT 22.395 155.015 22.675 155.385 ;
        RECT 17.635 152.635 19.175 153.005 ;
        RECT 21.545 149.070 21.685 154.870 ;
        RECT 22.465 154.850 22.605 155.015 ;
        RECT 22.405 154.530 22.665 154.850 ;
        RECT 21.485 148.750 21.745 149.070 ;
        RECT 22.405 148.585 22.665 148.730 ;
        RECT 22.395 148.215 22.675 148.585 ;
        RECT 17.635 147.195 19.175 147.565 ;
        RECT 17.635 141.755 19.175 142.125 ;
        RECT 21.945 140.250 22.205 140.570 ;
        RECT 22.005 138.190 22.145 140.250 ;
        RECT 21.945 137.870 22.205 138.190 ;
        RECT 21.025 136.850 21.285 137.170 ;
        RECT 17.635 136.315 19.175 136.685 ;
        RECT 17.635 130.875 19.175 131.245 ;
        RECT 21.085 129.350 21.225 136.850 ;
        RECT 21.485 132.430 21.745 132.750 ;
        RECT 21.545 132.265 21.685 132.430 ;
        RECT 21.475 131.895 21.755 132.265 ;
        RECT 19.645 129.030 19.905 129.350 ;
        RECT 21.025 129.030 21.285 129.350 ;
        RECT 17.635 125.435 19.175 125.805 ;
        RECT 19.705 124.785 19.845 129.030 ;
        RECT 19.635 124.415 19.915 124.785 ;
        RECT 21.545 124.250 21.685 131.895 ;
        RECT 22.005 127.310 22.145 137.870 ;
        RECT 23.325 136.850 23.585 137.170 ;
        RECT 23.385 136.150 23.525 136.850 ;
        RECT 23.325 135.830 23.585 136.150 ;
        RECT 24.305 135.130 24.445 165.410 ;
        RECT 24.765 165.390 24.905 174.930 ;
        RECT 28.445 173.210 28.585 183.770 ;
        RECT 31.205 182.050 31.345 185.810 ;
        RECT 32.585 185.110 32.725 188.870 ;
        RECT 35.745 188.530 36.005 188.850 ;
        RECT 36.665 188.530 36.925 188.850 ;
        RECT 35.805 187.490 35.945 188.530 ;
        RECT 35.745 187.170 36.005 187.490 ;
        RECT 32.985 186.150 33.245 186.470 ;
        RECT 32.525 184.790 32.785 185.110 ;
        RECT 31.605 184.680 31.865 184.770 ;
        RECT 31.605 184.540 32.265 184.680 ;
        RECT 31.605 184.450 31.865 184.540 ;
        RECT 32.125 183.750 32.265 184.540 ;
        RECT 32.525 183.770 32.785 184.090 ;
        RECT 32.065 183.430 32.325 183.750 ;
        RECT 31.605 183.090 31.865 183.410 ;
        RECT 31.665 182.050 31.805 183.090 ;
        RECT 32.125 182.390 32.265 183.430 ;
        RECT 32.065 182.070 32.325 182.390 ;
        RECT 31.145 181.730 31.405 182.050 ;
        RECT 31.605 181.730 31.865 182.050 ;
        RECT 31.145 181.050 31.405 181.370 ;
        RECT 29.765 177.650 30.025 177.970 ;
        RECT 29.825 176.610 29.965 177.650 ;
        RECT 29.765 176.290 30.025 176.610 ;
        RECT 31.205 176.270 31.345 181.050 ;
        RECT 31.605 178.330 31.865 178.650 ;
        RECT 32.585 178.560 32.725 183.770 ;
        RECT 33.045 183.750 33.185 186.150 ;
        RECT 36.725 184.430 36.865 188.530 ;
        RECT 39.485 184.770 39.625 192.270 ;
        RECT 40.345 189.550 40.605 189.870 ;
        RECT 40.405 188.850 40.545 189.550 ;
        RECT 39.885 188.530 40.145 188.850 ;
        RECT 40.345 188.530 40.605 188.850 ;
        RECT 39.425 184.510 39.685 184.770 ;
        RECT 38.565 184.450 39.685 184.510 ;
        RECT 36.665 184.110 36.925 184.430 ;
        RECT 38.565 184.370 39.625 184.450 ;
        RECT 39.945 184.430 40.085 188.530 ;
        RECT 40.405 187.150 40.545 188.530 ;
        RECT 40.345 186.830 40.605 187.150 ;
        RECT 40.405 184.770 40.545 186.830 ;
        RECT 40.345 184.450 40.605 184.770 ;
        RECT 38.565 183.750 38.705 184.370 ;
        RECT 38.965 183.770 39.225 184.090 ;
        RECT 32.985 183.430 33.245 183.750 ;
        RECT 37.585 183.430 37.845 183.750 ;
        RECT 38.505 183.430 38.765 183.750 ;
        RECT 33.045 181.030 33.185 183.430 ;
        RECT 35.745 181.390 36.005 181.710 ;
        RECT 32.985 180.710 33.245 181.030 ;
        RECT 35.285 180.370 35.545 180.690 ;
        RECT 33.435 178.815 33.715 179.185 ;
        RECT 35.345 178.990 35.485 180.370 ;
        RECT 33.445 178.670 33.705 178.815 ;
        RECT 34.365 178.670 34.625 178.990 ;
        RECT 35.285 178.670 35.545 178.990 ;
        RECT 32.985 178.560 33.245 178.650 ;
        RECT 32.585 178.420 33.245 178.560 ;
        RECT 32.985 178.330 33.245 178.420 ;
        RECT 31.665 176.950 31.805 178.330 ;
        RECT 31.605 176.630 31.865 176.950 ;
        RECT 33.505 176.270 33.645 178.670 ;
        RECT 31.145 176.180 31.405 176.270 ;
        RECT 30.745 176.040 31.405 176.180 ;
        RECT 28.385 172.890 28.645 173.210 ;
        RECT 28.845 170.850 29.105 171.170 ;
        RECT 26.085 169.490 26.345 169.810 ;
        RECT 26.145 168.790 26.285 169.490 ;
        RECT 26.085 168.470 26.345 168.790 ;
        RECT 26.545 167.790 26.805 168.110 ;
        RECT 26.605 166.070 26.745 167.790 ;
        RECT 28.385 167.110 28.645 167.430 ;
        RECT 28.445 166.070 28.585 167.110 ;
        RECT 28.905 166.070 29.045 170.850 ;
        RECT 30.745 170.490 30.885 176.040 ;
        RECT 31.145 175.950 31.405 176.040 ;
        RECT 33.445 175.950 33.705 176.270 ;
        RECT 34.425 175.930 34.565 178.670 ;
        RECT 35.805 178.650 35.945 181.390 ;
        RECT 37.645 180.940 37.785 183.430 ;
        RECT 38.505 181.390 38.765 181.710 ;
        RECT 38.045 180.940 38.305 181.030 ;
        RECT 37.645 180.800 38.305 180.940 ;
        RECT 38.045 180.710 38.305 180.800 ;
        RECT 36.665 180.370 36.925 180.690 ;
        RECT 35.745 178.330 36.005 178.650 ;
        RECT 35.285 177.990 35.545 178.310 ;
        RECT 34.365 175.610 34.625 175.930 ;
        RECT 33.445 174.930 33.705 175.250 ;
        RECT 32.975 172.695 33.255 173.065 ;
        RECT 33.045 172.530 33.185 172.695 ;
        RECT 32.985 172.210 33.245 172.530 ;
        RECT 30.685 170.170 30.945 170.490 ;
        RECT 32.065 170.170 32.325 170.490 ;
        RECT 30.745 168.110 30.885 170.170 ;
        RECT 31.605 169.490 31.865 169.810 ;
        RECT 30.685 167.790 30.945 168.110 ;
        RECT 26.545 165.750 26.805 166.070 ;
        RECT 28.385 165.750 28.645 166.070 ;
        RECT 28.845 165.750 29.105 166.070 ;
        RECT 24.705 165.070 24.965 165.390 ;
        RECT 24.765 156.890 24.905 165.070 ;
        RECT 29.765 164.730 30.025 165.050 ;
        RECT 29.825 163.350 29.965 164.730 ;
        RECT 30.745 163.350 30.885 167.790 ;
        RECT 29.765 163.030 30.025 163.350 ;
        RECT 30.685 163.030 30.945 163.350 ;
        RECT 30.225 161.670 30.485 161.990 ;
        RECT 30.285 157.910 30.425 161.670 ;
        RECT 30.225 157.590 30.485 157.910 ;
        RECT 31.665 157.570 31.805 169.490 ;
        RECT 32.125 166.070 32.265 170.170 ;
        RECT 33.505 168.450 33.645 174.930 ;
        RECT 34.425 173.550 34.565 175.610 ;
        RECT 34.365 173.230 34.625 173.550 ;
        RECT 35.345 173.210 35.485 177.990 ;
        RECT 35.805 176.270 35.945 178.330 ;
        RECT 35.745 175.950 36.005 176.270 ;
        RECT 35.805 175.590 35.945 175.950 ;
        RECT 36.725 175.590 36.865 180.370 ;
        RECT 38.105 179.185 38.245 180.710 ;
        RECT 38.565 179.330 38.705 181.390 ;
        RECT 37.585 178.670 37.845 178.990 ;
        RECT 38.035 178.815 38.315 179.185 ;
        RECT 38.505 179.010 38.765 179.330 ;
        RECT 38.045 178.670 38.305 178.815 ;
        RECT 37.645 176.950 37.785 178.670 ;
        RECT 38.565 178.390 38.705 179.010 ;
        RECT 38.105 178.310 38.705 178.390 ;
        RECT 38.045 178.250 38.705 178.310 ;
        RECT 38.045 177.990 38.305 178.250 ;
        RECT 37.585 176.630 37.845 176.950 ;
        RECT 38.105 175.930 38.245 177.990 ;
        RECT 38.505 176.290 38.765 176.610 ;
        RECT 38.045 175.610 38.305 175.930 ;
        RECT 35.745 175.270 36.005 175.590 ;
        RECT 36.665 175.270 36.925 175.590 ;
        RECT 37.585 175.270 37.845 175.590 ;
        RECT 35.805 174.990 35.945 175.270 ;
        RECT 35.805 174.850 36.865 174.990 ;
        RECT 35.745 173.910 36.005 174.230 ;
        RECT 35.285 172.890 35.545 173.210 ;
        RECT 35.805 171.510 35.945 173.910 ;
        RECT 36.725 173.890 36.865 174.850 ;
        RECT 36.205 173.745 36.465 173.890 ;
        RECT 36.195 173.375 36.475 173.745 ;
        RECT 36.665 173.570 36.925 173.890 ;
        RECT 36.205 172.550 36.465 172.870 ;
        RECT 35.745 171.190 36.005 171.510 ;
        RECT 33.445 168.130 33.705 168.450 ;
        RECT 33.505 167.510 33.645 168.130 ;
        RECT 35.805 168.110 35.945 171.190 ;
        RECT 36.265 170.830 36.405 172.550 ;
        RECT 36.205 170.510 36.465 170.830 ;
        RECT 37.125 169.665 37.385 169.810 ;
        RECT 37.115 169.295 37.395 169.665 ;
        RECT 35.745 167.790 36.005 168.110 ;
        RECT 33.045 167.370 33.645 167.510 ;
        RECT 33.045 166.070 33.185 167.370 ;
        RECT 35.745 167.110 36.005 167.430 ;
        RECT 37.125 167.110 37.385 167.430 ;
        RECT 33.445 166.770 33.705 167.090 ;
        RECT 34.365 166.770 34.625 167.090 ;
        RECT 35.285 166.770 35.545 167.090 ;
        RECT 32.065 165.750 32.325 166.070 ;
        RECT 32.985 165.750 33.245 166.070 ;
        RECT 32.525 163.030 32.785 163.350 ;
        RECT 32.585 159.950 32.725 163.030 ;
        RECT 33.505 162.750 33.645 166.770 ;
        RECT 34.425 165.390 34.565 166.770 ;
        RECT 34.365 165.070 34.625 165.390 ;
        RECT 34.815 165.215 35.095 165.585 ;
        RECT 34.825 165.070 35.085 165.215 ;
        RECT 33.045 162.670 33.645 162.750 ;
        RECT 32.985 162.610 33.645 162.670 ;
        RECT 32.985 162.350 33.245 162.610 ;
        RECT 32.985 161.670 33.245 161.990 ;
        RECT 33.045 160.630 33.185 161.670 ;
        RECT 32.985 160.310 33.245 160.630 ;
        RECT 32.525 159.630 32.785 159.950 ;
        RECT 31.605 157.250 31.865 157.570 ;
        RECT 24.705 156.570 24.965 156.890 ;
        RECT 30.225 156.570 30.485 156.890 ;
        RECT 32.065 156.570 32.325 156.890 ;
        RECT 25.165 155.890 25.425 156.210 ;
        RECT 25.225 136.150 25.365 155.890 ;
        RECT 30.285 153.490 30.425 156.570 ;
        RECT 30.225 153.170 30.485 153.490 ;
        RECT 26.085 152.150 26.345 152.470 ;
        RECT 26.145 146.350 26.285 152.150 ;
        RECT 29.765 150.790 30.025 151.110 ;
        RECT 29.825 147.030 29.965 150.790 ;
        RECT 29.765 146.710 30.025 147.030 ;
        RECT 26.085 146.030 26.345 146.350 ;
        RECT 30.285 146.010 30.425 153.170 ;
        RECT 32.125 152.470 32.265 156.570 ;
        RECT 32.585 154.510 32.725 159.630 ;
        RECT 33.505 159.610 33.645 162.610 ;
        RECT 33.905 160.310 34.165 160.630 ;
        RECT 33.445 159.290 33.705 159.610 ;
        RECT 33.445 158.610 33.705 158.930 ;
        RECT 33.505 156.550 33.645 158.610 ;
        RECT 33.445 156.230 33.705 156.550 ;
        RECT 32.525 154.190 32.785 154.510 ;
        RECT 32.065 152.150 32.325 152.470 ;
        RECT 32.585 151.790 32.725 154.190 ;
        RECT 32.525 151.470 32.785 151.790 ;
        RECT 32.585 149.070 32.725 151.470 ;
        RECT 32.525 148.750 32.785 149.070 ;
        RECT 32.985 147.730 33.245 148.050 ;
        RECT 30.225 145.690 30.485 146.010 ;
        RECT 32.525 145.010 32.785 145.330 ;
        RECT 32.585 144.310 32.725 145.010 ;
        RECT 32.525 143.990 32.785 144.310 ;
        RECT 33.045 143.630 33.185 147.730 ;
        RECT 33.965 146.350 34.105 160.310 ;
        RECT 34.365 159.630 34.625 159.950 ;
        RECT 34.425 157.910 34.565 159.630 ;
        RECT 34.365 157.590 34.625 157.910 ;
        RECT 34.885 156.890 35.025 165.070 ;
        RECT 35.345 164.370 35.485 166.770 ;
        RECT 35.285 164.050 35.545 164.370 ;
        RECT 35.805 159.610 35.945 167.110 ;
        RECT 36.205 165.750 36.465 166.070 ;
        RECT 35.745 159.290 36.005 159.610 ;
        RECT 34.825 156.800 35.085 156.890 ;
        RECT 34.825 156.660 35.485 156.800 ;
        RECT 34.825 156.570 35.085 156.660 ;
        RECT 34.825 153.170 35.085 153.490 ;
        RECT 34.365 150.790 34.625 151.110 ;
        RECT 34.425 147.030 34.565 150.790 ;
        RECT 34.885 149.070 35.025 153.170 ;
        RECT 35.345 151.790 35.485 156.660 ;
        RECT 35.285 151.470 35.545 151.790 ;
        RECT 34.825 148.750 35.085 149.070 ;
        RECT 34.365 146.710 34.625 147.030 ;
        RECT 35.805 146.350 35.945 159.290 ;
        RECT 36.265 157.230 36.405 165.750 ;
        RECT 36.665 164.730 36.925 165.050 ;
        RECT 36.725 163.350 36.865 164.730 ;
        RECT 37.185 163.350 37.325 167.110 ;
        RECT 36.665 163.030 36.925 163.350 ;
        RECT 37.125 163.030 37.385 163.350 ;
        RECT 37.185 161.650 37.325 163.030 ;
        RECT 37.125 161.330 37.385 161.650 ;
        RECT 36.205 157.140 36.465 157.230 ;
        RECT 36.205 157.000 37.325 157.140 ;
        RECT 36.205 156.910 36.465 157.000 ;
        RECT 36.665 154.190 36.925 154.510 ;
        RECT 36.205 153.170 36.465 153.490 ;
        RECT 36.265 151.450 36.405 153.170 ;
        RECT 36.725 152.470 36.865 154.190 ;
        RECT 36.665 152.150 36.925 152.470 ;
        RECT 37.185 151.450 37.325 157.000 ;
        RECT 37.645 154.420 37.785 175.270 ;
        RECT 38.105 173.550 38.245 175.610 ;
        RECT 38.565 173.550 38.705 176.290 ;
        RECT 39.025 175.930 39.165 183.770 ;
        RECT 39.485 181.710 39.625 184.370 ;
        RECT 39.885 184.110 40.145 184.430 ;
        RECT 39.425 181.390 39.685 181.710 ;
        RECT 40.405 181.370 40.545 184.450 ;
        RECT 40.865 181.710 41.005 192.270 ;
        RECT 41.725 191.590 41.985 191.910 ;
        RECT 41.785 186.810 41.925 191.590 ;
        RECT 47.305 189.870 47.445 194.340 ;
        RECT 53.205 193.435 54.745 193.805 ;
        RECT 60.125 192.270 60.385 192.590 ;
        RECT 50.925 191.250 51.185 191.570 ;
        RECT 59.665 191.250 59.925 191.570 ;
        RECT 47.245 189.550 47.505 189.870 ;
        RECT 50.985 189.190 51.125 191.250 ;
        RECT 56.505 190.715 58.045 191.085 ;
        RECT 54.605 189.780 54.865 189.870 ;
        RECT 54.605 189.640 55.265 189.780 ;
        RECT 54.605 189.550 54.865 189.640 ;
        RECT 44.485 188.870 44.745 189.190 ;
        RECT 50.925 188.870 51.185 189.190 ;
        RECT 44.545 187.830 44.685 188.870 ;
        RECT 53.205 187.995 54.745 188.365 ;
        RECT 44.485 187.510 44.745 187.830 ;
        RECT 54.145 187.170 54.405 187.490 ;
        RECT 42.185 186.830 42.445 187.150 ;
        RECT 44.025 186.830 44.285 187.150 ;
        RECT 46.325 186.830 46.585 187.150 ;
        RECT 41.725 186.490 41.985 186.810 ;
        RECT 41.785 183.410 41.925 186.490 ;
        RECT 41.725 183.090 41.985 183.410 ;
        RECT 40.805 181.390 41.065 181.710 ;
        RECT 40.345 181.050 40.605 181.370 ;
        RECT 42.245 181.030 42.385 186.830 ;
        RECT 44.085 185.110 44.225 186.830 ;
        RECT 44.485 186.490 44.745 186.810 ;
        RECT 44.025 184.790 44.285 185.110 ;
        RECT 44.025 181.050 44.285 181.370 ;
        RECT 42.185 180.710 42.445 181.030 ;
        RECT 43.565 180.710 43.825 181.030 ;
        RECT 42.245 179.670 42.385 180.710 ;
        RECT 42.185 179.350 42.445 179.670 ;
        RECT 42.245 178.990 42.385 179.350 ;
        RECT 42.185 178.670 42.445 178.990 ;
        RECT 43.625 176.950 43.765 180.710 ;
        RECT 39.425 176.630 39.685 176.950 ;
        RECT 43.565 176.630 43.825 176.950 ;
        RECT 39.485 176.465 39.625 176.630 ;
        RECT 39.415 176.095 39.695 176.465 ;
        RECT 41.715 176.095 41.995 176.465 ;
        RECT 43.105 176.290 43.365 176.610 ;
        RECT 38.965 175.610 39.225 175.930 ;
        RECT 38.045 173.230 38.305 173.550 ;
        RECT 38.505 173.230 38.765 173.550 ;
        RECT 41.785 173.210 41.925 176.095 ;
        RECT 42.185 175.610 42.445 175.930 ;
        RECT 42.245 173.210 42.385 175.610 ;
        RECT 43.165 173.210 43.305 176.290 ;
        RECT 44.085 175.670 44.225 181.050 ;
        RECT 43.625 175.530 44.225 175.670 ;
        RECT 41.265 172.890 41.525 173.210 ;
        RECT 41.725 173.065 41.985 173.210 ;
        RECT 38.965 172.210 39.225 172.530 ;
        RECT 38.505 170.510 38.765 170.830 ;
        RECT 38.045 169.490 38.305 169.810 ;
        RECT 38.105 168.790 38.245 169.490 ;
        RECT 38.045 168.470 38.305 168.790 ;
        RECT 38.105 165.390 38.245 168.470 ;
        RECT 38.045 165.070 38.305 165.390 ;
        RECT 38.105 160.630 38.245 165.070 ;
        RECT 38.045 160.310 38.305 160.630 ;
        RECT 38.045 158.610 38.305 158.930 ;
        RECT 38.105 157.910 38.245 158.610 ;
        RECT 38.045 157.590 38.305 157.910 ;
        RECT 38.565 156.890 38.705 170.510 ;
        RECT 39.025 164.710 39.165 172.210 ;
        RECT 39.885 171.190 40.145 171.510 ;
        RECT 38.965 164.390 39.225 164.710 ;
        RECT 38.965 163.030 39.225 163.350 ;
        RECT 38.505 156.570 38.765 156.890 ;
        RECT 38.565 155.190 38.705 156.570 ;
        RECT 39.025 156.550 39.165 163.030 ;
        RECT 39.425 159.630 39.685 159.950 ;
        RECT 39.485 157.910 39.625 159.630 ;
        RECT 39.425 157.590 39.685 157.910 ;
        RECT 39.945 156.550 40.085 171.190 ;
        RECT 40.345 170.510 40.605 170.830 ;
        RECT 40.405 169.810 40.545 170.510 ;
        RECT 40.805 169.830 41.065 170.150 ;
        RECT 40.345 169.490 40.605 169.810 ;
        RECT 40.345 167.790 40.605 168.110 ;
        RECT 40.405 166.070 40.545 167.790 ;
        RECT 40.865 167.090 41.005 169.830 ;
        RECT 40.805 166.770 41.065 167.090 ;
        RECT 40.345 165.750 40.605 166.070 ;
        RECT 40.865 160.630 41.005 166.770 ;
        RECT 40.805 160.310 41.065 160.630 ;
        RECT 41.325 159.950 41.465 172.890 ;
        RECT 41.715 172.695 41.995 173.065 ;
        RECT 42.185 172.890 42.445 173.210 ;
        RECT 43.105 173.120 43.365 173.210 ;
        RECT 42.705 172.980 43.365 173.120 ;
        RECT 42.705 170.830 42.845 172.980 ;
        RECT 43.105 172.890 43.365 172.980 ;
        RECT 43.105 171.190 43.365 171.510 ;
        RECT 42.645 170.510 42.905 170.830 ;
        RECT 43.165 170.230 43.305 171.190 ;
        RECT 43.625 170.910 43.765 175.530 ;
        RECT 44.025 172.210 44.285 172.530 ;
        RECT 44.085 171.510 44.225 172.210 ;
        RECT 44.025 171.190 44.285 171.510 ;
        RECT 43.625 170.770 44.225 170.910 ;
        RECT 44.085 170.490 44.225 170.770 ;
        RECT 43.165 170.090 43.765 170.230 ;
        RECT 44.025 170.170 44.285 170.490 ;
        RECT 43.625 169.810 43.765 170.090 ;
        RECT 43.105 169.490 43.365 169.810 ;
        RECT 43.565 169.490 43.825 169.810 ;
        RECT 42.185 167.110 42.445 167.430 ;
        RECT 41.725 162.350 41.985 162.670 ;
        RECT 41.265 159.630 41.525 159.950 ;
        RECT 40.805 159.290 41.065 159.610 ;
        RECT 38.965 156.230 39.225 156.550 ;
        RECT 39.885 156.230 40.145 156.550 ;
        RECT 39.025 155.270 39.165 156.230 ;
        RECT 40.865 155.950 41.005 159.290 ;
        RECT 41.325 158.930 41.465 159.630 ;
        RECT 41.785 159.270 41.925 162.350 ;
        RECT 42.245 159.950 42.385 167.110 ;
        RECT 42.645 166.770 42.905 167.090 ;
        RECT 42.185 159.630 42.445 159.950 ;
        RECT 41.725 158.950 41.985 159.270 ;
        RECT 41.265 158.610 41.525 158.930 ;
        RECT 41.785 156.890 41.925 158.950 ;
        RECT 42.245 157.910 42.385 159.630 ;
        RECT 42.185 157.590 42.445 157.910 ;
        RECT 42.705 157.570 42.845 166.770 ;
        RECT 43.165 165.730 43.305 169.490 ;
        RECT 43.565 167.790 43.825 168.110 ;
        RECT 43.105 165.410 43.365 165.730 ;
        RECT 43.625 164.790 43.765 167.790 ;
        RECT 43.165 164.650 43.765 164.790 ;
        RECT 42.645 157.250 42.905 157.570 ;
        RECT 41.725 156.570 41.985 156.890 ;
        RECT 42.185 156.570 42.445 156.890 ;
        RECT 42.245 155.950 42.385 156.570 ;
        RECT 40.865 155.810 42.385 155.950 ;
        RECT 38.505 154.870 38.765 155.190 ;
        RECT 39.025 155.130 39.625 155.270 ;
        RECT 42.705 155.190 42.845 157.250 ;
        RECT 38.045 154.420 38.305 154.510 ;
        RECT 37.645 154.280 38.305 154.420 ;
        RECT 38.045 154.190 38.305 154.280 ;
        RECT 37.575 153.655 37.855 154.025 ;
        RECT 36.205 151.130 36.465 151.450 ;
        RECT 36.665 151.130 36.925 151.450 ;
        RECT 37.125 151.130 37.385 151.450 ;
        RECT 36.725 148.050 36.865 151.130 ;
        RECT 36.665 147.730 36.925 148.050 ;
        RECT 33.905 146.030 34.165 146.350 ;
        RECT 35.745 146.030 36.005 146.350 ;
        RECT 37.645 146.010 37.785 153.655 ;
        RECT 38.105 149.265 38.245 154.190 ;
        RECT 38.035 148.895 38.315 149.265 ;
        RECT 33.445 145.690 33.705 146.010 ;
        RECT 37.585 145.690 37.845 146.010 ;
        RECT 32.985 143.310 33.245 143.630 ;
        RECT 30.225 139.570 30.485 139.890 ;
        RECT 30.285 138.530 30.425 139.570 ;
        RECT 32.985 138.550 33.245 138.870 ;
        RECT 30.225 138.210 30.485 138.530 ;
        RECT 32.525 136.850 32.785 137.170 ;
        RECT 25.165 135.830 25.425 136.150 ;
        RECT 32.585 135.470 32.725 136.850 ;
        RECT 32.525 135.150 32.785 135.470 ;
        RECT 24.245 134.810 24.505 135.130 ;
        RECT 30.685 134.810 30.945 135.130 ;
        RECT 27.925 134.130 28.185 134.450 ;
        RECT 25.625 131.410 25.885 131.730 ;
        RECT 26.085 131.410 26.345 131.730 ;
        RECT 25.685 130.710 25.825 131.410 ;
        RECT 25.625 130.390 25.885 130.710 ;
        RECT 21.945 126.990 22.205 127.310 ;
        RECT 24.245 126.990 24.505 127.310 ;
        RECT 22.405 126.650 22.665 126.970 ;
        RECT 21.485 123.930 21.745 124.250 ;
        RECT 21.945 123.250 22.205 123.570 ;
        RECT 22.005 122.550 22.145 123.250 ;
        RECT 21.945 122.230 22.205 122.550 ;
        RECT 22.465 121.385 22.605 126.650 ;
        RECT 24.305 121.870 24.445 126.990 ;
        RECT 26.145 124.590 26.285 131.410 ;
        RECT 26.085 124.270 26.345 124.590 ;
        RECT 24.695 123.735 24.975 124.105 ;
        RECT 24.705 123.590 24.965 123.735 ;
        RECT 26.145 122.210 26.285 124.270 ;
        RECT 26.085 121.890 26.345 122.210 ;
        RECT 27.985 121.870 28.125 134.130 ;
        RECT 30.745 130.710 30.885 134.810 ;
        RECT 32.585 134.310 32.725 135.150 ;
        RECT 33.045 135.130 33.185 138.550 ;
        RECT 33.505 135.470 33.645 145.690 ;
        RECT 38.565 140.570 38.705 154.870 ;
        RECT 38.965 154.190 39.225 154.510 ;
        RECT 39.025 152.470 39.165 154.190 ;
        RECT 38.965 152.150 39.225 152.470 ;
        RECT 38.965 151.130 39.225 151.450 ;
        RECT 38.505 140.250 38.765 140.570 ;
        RECT 34.365 139.910 34.625 140.230 ;
        RECT 33.905 138.550 34.165 138.870 ;
        RECT 33.445 135.150 33.705 135.470 ;
        RECT 32.985 134.810 33.245 135.130 ;
        RECT 32.585 134.170 33.185 134.310 ;
        RECT 33.045 133.090 33.185 134.170 ;
        RECT 32.985 132.770 33.245 133.090 ;
        RECT 33.445 131.410 33.705 131.730 ;
        RECT 33.505 130.710 33.645 131.410 ;
        RECT 30.685 130.390 30.945 130.710 ;
        RECT 33.445 130.390 33.705 130.710 ;
        RECT 32.065 130.110 32.325 130.370 ;
        RECT 32.065 130.050 33.645 130.110 ;
        RECT 32.125 130.030 33.645 130.050 ;
        RECT 32.125 129.970 33.705 130.030 ;
        RECT 33.445 129.710 33.705 129.970 ;
        RECT 32.985 129.030 33.245 129.350 ;
        RECT 30.225 128.690 30.485 129.010 ;
        RECT 32.065 128.690 32.325 129.010 ;
        RECT 30.285 125.270 30.425 128.690 ;
        RECT 31.145 126.650 31.405 126.970 ;
        RECT 30.225 124.950 30.485 125.270 ;
        RECT 24.245 121.550 24.505 121.870 ;
        RECT 26.545 121.550 26.805 121.870 ;
        RECT 27.925 121.550 28.185 121.870 ;
        RECT 28.385 121.550 28.645 121.870 ;
        RECT 22.395 121.015 22.675 121.385 ;
        RECT 17.635 119.995 19.175 120.365 ;
        RECT 19.645 118.150 19.905 118.470 ;
        RECT 19.705 117.985 19.845 118.150 ;
        RECT 19.635 117.615 19.915 117.985 ;
        RECT 22.865 115.945 23.125 116.090 ;
        RECT 22.855 115.575 23.135 115.945 ;
        RECT 17.635 114.555 19.175 114.925 ;
        RECT 24.305 113.370 24.445 121.550 ;
        RECT 24.705 120.530 24.965 120.850 ;
        RECT 24.765 118.470 24.905 120.530 ;
        RECT 26.605 119.830 26.745 121.550 ;
        RECT 26.545 119.510 26.805 119.830 ;
        RECT 28.445 119.345 28.585 121.550 ;
        RECT 30.225 121.210 30.485 121.530 ;
        RECT 29.765 120.530 30.025 120.850 ;
        RECT 28.375 118.975 28.655 119.345 ;
        RECT 24.705 118.150 24.965 118.470 ;
        RECT 26.545 116.450 26.805 116.770 ;
        RECT 26.605 114.390 26.745 116.450 ;
        RECT 26.545 114.070 26.805 114.390 ;
        RECT 24.245 113.050 24.505 113.370 ;
        RECT 27.925 113.050 28.185 113.370 ;
        RECT 24.305 110.990 24.445 113.050 ;
        RECT 24.245 110.670 24.505 110.990 ;
        RECT 17.635 109.115 19.175 109.485 ;
        RECT 24.305 107.930 24.445 110.670 ;
        RECT 27.985 110.650 28.125 113.050 ;
        RECT 29.825 111.330 29.965 120.530 ;
        RECT 30.285 118.810 30.425 121.210 ;
        RECT 30.225 118.490 30.485 118.810 ;
        RECT 30.225 113.050 30.485 113.370 ;
        RECT 29.765 111.010 30.025 111.330 ;
        RECT 27.925 110.330 28.185 110.650 ;
        RECT 30.285 108.610 30.425 113.050 ;
        RECT 31.205 112.690 31.345 126.650 ;
        RECT 32.125 124.250 32.265 128.690 ;
        RECT 33.045 126.970 33.185 129.030 ;
        RECT 32.985 126.650 33.245 126.970 ;
        RECT 32.525 125.970 32.785 126.290 ;
        RECT 32.065 123.930 32.325 124.250 ;
        RECT 31.605 121.890 31.865 122.210 ;
        RECT 31.665 119.830 31.805 121.890 ;
        RECT 31.605 119.510 31.865 119.830 ;
        RECT 32.065 118.150 32.325 118.470 ;
        RECT 31.145 112.370 31.405 112.690 ;
        RECT 32.125 111.670 32.265 118.150 ;
        RECT 32.585 113.370 32.725 125.970 ;
        RECT 33.045 118.810 33.185 126.650 ;
        RECT 33.505 124.590 33.645 129.710 ;
        RECT 33.965 127.310 34.105 138.550 ;
        RECT 33.905 126.990 34.165 127.310 ;
        RECT 33.445 124.270 33.705 124.590 ;
        RECT 33.445 123.250 33.705 123.570 ;
        RECT 33.905 123.250 34.165 123.570 ;
        RECT 33.505 122.550 33.645 123.250 ;
        RECT 33.445 122.230 33.705 122.550 ;
        RECT 33.965 119.150 34.105 123.250 ;
        RECT 33.905 118.830 34.165 119.150 ;
        RECT 32.985 118.490 33.245 118.810 ;
        RECT 33.045 116.430 33.185 118.490 ;
        RECT 32.985 116.110 33.245 116.430 ;
        RECT 32.525 113.050 32.785 113.370 ;
        RECT 32.985 112.370 33.245 112.690 ;
        RECT 33.445 112.370 33.705 112.690 ;
        RECT 32.065 111.350 32.325 111.670 ;
        RECT 33.045 110.390 33.185 112.370 ;
        RECT 33.505 110.990 33.645 112.370 ;
        RECT 34.425 111.330 34.565 139.910 ;
        RECT 36.665 139.570 36.925 139.890 ;
        RECT 36.725 138.530 36.865 139.570 ;
        RECT 36.665 138.210 36.925 138.530 ;
        RECT 34.825 137.190 35.085 137.510 ;
        RECT 34.885 132.410 35.025 137.190 ;
        RECT 37.125 135.830 37.385 136.150 ;
        RECT 35.285 135.490 35.545 135.810 ;
        RECT 34.825 132.090 35.085 132.410 ;
        RECT 34.885 129.350 35.025 132.090 ;
        RECT 35.345 130.030 35.485 135.490 ;
        RECT 37.185 135.130 37.325 135.830 ;
        RECT 37.585 135.150 37.845 135.470 ;
        RECT 37.125 134.810 37.385 135.130 ;
        RECT 35.745 134.130 36.005 134.450 ;
        RECT 35.805 133.430 35.945 134.130 ;
        RECT 35.745 133.110 36.005 133.430 ;
        RECT 37.185 132.945 37.325 134.810 ;
        RECT 36.665 132.430 36.925 132.750 ;
        RECT 37.115 132.575 37.395 132.945 ;
        RECT 35.745 131.410 36.005 131.730 ;
        RECT 36.205 131.410 36.465 131.730 ;
        RECT 35.285 129.710 35.545 130.030 ;
        RECT 34.825 129.030 35.085 129.350 ;
        RECT 34.825 126.990 35.085 127.310 ;
        RECT 34.885 122.065 35.025 126.990 ;
        RECT 35.805 123.910 35.945 131.410 ;
        RECT 36.265 124.250 36.405 131.410 ;
        RECT 36.725 130.030 36.865 132.430 ;
        RECT 37.645 132.410 37.785 135.150 ;
        RECT 38.045 135.040 38.305 135.130 ;
        RECT 38.565 135.040 38.705 140.250 ;
        RECT 39.025 138.870 39.165 151.130 ;
        RECT 39.485 148.585 39.625 155.130 ;
        RECT 42.645 154.870 42.905 155.190 ;
        RECT 41.265 153.850 41.525 154.170 ;
        RECT 40.805 153.510 41.065 153.830 ;
        RECT 39.885 153.170 40.145 153.490 ;
        RECT 39.945 149.750 40.085 153.170 ;
        RECT 39.885 149.430 40.145 149.750 ;
        RECT 40.865 149.410 41.005 153.510 ;
        RECT 41.325 152.470 41.465 153.850 ;
        RECT 42.185 153.170 42.445 153.490 ;
        RECT 41.265 152.150 41.525 152.470 ;
        RECT 40.345 149.090 40.605 149.410 ;
        RECT 40.805 149.090 41.065 149.410 ;
        RECT 39.415 148.215 39.695 148.585 ;
        RECT 40.405 147.030 40.545 149.090 ;
        RECT 42.245 147.030 42.385 153.170 ;
        RECT 42.705 152.130 42.845 154.870 ;
        RECT 43.165 154.170 43.305 164.650 ;
        RECT 43.565 159.970 43.825 160.290 ;
        RECT 43.625 156.745 43.765 159.970 ;
        RECT 44.085 159.610 44.225 170.170 ;
        RECT 44.545 167.770 44.685 186.490 ;
        RECT 44.945 179.350 45.205 179.670 ;
        RECT 45.005 176.950 45.145 179.350 ;
        RECT 45.405 177.650 45.665 177.970 ;
        RECT 44.945 176.630 45.205 176.950 ;
        RECT 45.465 176.270 45.605 177.650 ;
        RECT 45.405 176.180 45.665 176.270 ;
        RECT 45.405 176.040 46.065 176.180 ;
        RECT 45.405 175.950 45.665 176.040 ;
        RECT 45.925 170.830 46.065 176.040 ;
        RECT 45.865 170.510 46.125 170.830 ;
        RECT 46.385 168.700 46.525 186.830 ;
        RECT 49.085 186.150 49.345 186.470 ;
        RECT 48.165 178.560 48.425 178.650 ;
        RECT 49.145 178.560 49.285 186.150 ;
        RECT 49.545 185.810 49.805 186.130 ;
        RECT 53.225 185.810 53.485 186.130 ;
        RECT 49.605 184.430 49.745 185.810 ;
        RECT 49.545 184.110 49.805 184.430 ;
        RECT 53.285 183.750 53.425 185.810 ;
        RECT 54.205 185.110 54.345 187.170 ;
        RECT 54.145 184.790 54.405 185.110 ;
        RECT 53.225 183.430 53.485 183.750 ;
        RECT 53.205 182.555 54.745 182.925 ;
        RECT 55.125 182.390 55.265 189.640 ;
        RECT 57.825 189.550 58.085 189.870 ;
        RECT 55.985 189.210 56.245 189.530 ;
        RECT 56.045 187.150 56.185 189.210 ;
        RECT 57.885 187.830 58.025 189.550 ;
        RECT 58.285 188.530 58.545 188.850 ;
        RECT 58.745 188.530 59.005 188.850 ;
        RECT 57.825 187.510 58.085 187.830 ;
        RECT 55.985 186.830 56.245 187.150 ;
        RECT 55.525 185.810 55.785 186.130 ;
        RECT 55.585 184.430 55.725 185.810 ;
        RECT 55.525 184.110 55.785 184.430 ;
        RECT 52.305 182.070 52.565 182.390 ;
        RECT 55.065 182.070 55.325 182.390 ;
        RECT 51.385 181.050 51.645 181.370 ;
        RECT 48.165 178.420 49.285 178.560 ;
        RECT 48.165 178.330 48.425 178.420 ;
        RECT 49.145 176.270 49.285 178.420 ;
        RECT 50.925 177.650 51.185 177.970 ;
        RECT 50.985 176.270 51.125 177.650 ;
        RECT 51.445 176.950 51.585 181.050 ;
        RECT 51.835 178.815 52.115 179.185 ;
        RECT 52.365 178.990 52.505 182.070 ;
        RECT 55.065 181.390 55.325 181.710 ;
        RECT 51.385 176.630 51.645 176.950 ;
        RECT 49.085 175.950 49.345 176.270 ;
        RECT 50.925 175.950 51.185 176.270 ;
        RECT 48.625 175.610 48.885 175.930 ;
        RECT 48.685 172.870 48.825 175.610 ;
        RECT 48.625 172.550 48.885 172.870 ;
        RECT 45.925 168.560 46.525 168.700 ;
        RECT 45.925 168.110 46.065 168.560 ;
        RECT 45.865 167.790 46.125 168.110 ;
        RECT 49.145 167.770 49.285 175.950 ;
        RECT 51.385 172.550 51.645 172.870 ;
        RECT 51.445 171.510 51.585 172.550 ;
        RECT 51.905 171.510 52.045 178.815 ;
        RECT 52.305 178.670 52.565 178.990 ;
        RECT 53.205 177.115 54.745 177.485 ;
        RECT 55.125 176.950 55.265 181.390 ;
        RECT 55.525 180.710 55.785 181.030 ;
        RECT 55.585 177.145 55.725 180.710 ;
        RECT 56.045 178.650 56.185 186.830 ;
        RECT 57.885 186.040 58.025 187.510 ;
        RECT 58.345 187.150 58.485 188.530 ;
        RECT 58.285 186.830 58.545 187.150 ;
        RECT 57.885 185.900 58.485 186.040 ;
        RECT 56.505 185.275 58.045 185.645 ;
        RECT 58.345 184.770 58.485 185.900 ;
        RECT 58.805 185.110 58.945 188.530 ;
        RECT 59.725 187.830 59.865 191.250 ;
        RECT 59.665 187.510 59.925 187.830 ;
        RECT 60.185 186.130 60.325 192.270 ;
        RECT 63.405 189.530 63.545 194.340 ;
        RECT 66.565 192.270 66.825 192.590 ;
        RECT 66.105 191.250 66.365 191.570 ;
        RECT 60.585 189.210 60.845 189.530 ;
        RECT 63.345 189.210 63.605 189.530 ;
        RECT 60.645 187.830 60.785 189.210 ;
        RECT 66.165 189.190 66.305 191.250 ;
        RECT 66.105 188.870 66.365 189.190 ;
        RECT 66.625 188.850 66.765 192.270 ;
        RECT 74.385 189.890 74.645 190.210 ;
        RECT 67.025 189.550 67.285 189.870 ;
        RECT 66.565 188.530 66.825 188.850 ;
        RECT 60.585 187.510 60.845 187.830 ;
        RECT 60.125 185.810 60.385 186.130 ;
        RECT 58.745 184.790 59.005 185.110 ;
        RECT 58.285 184.450 58.545 184.770 ;
        RECT 58.285 182.070 58.545 182.390 ;
        RECT 58.345 181.710 58.485 182.070 ;
        RECT 58.805 181.710 58.945 184.790 ;
        RECT 60.185 184.430 60.325 185.810 ;
        RECT 60.125 184.110 60.385 184.430 ;
        RECT 59.205 183.770 59.465 184.090 ;
        RECT 58.285 181.390 58.545 181.710 ;
        RECT 58.745 181.390 59.005 181.710 ;
        RECT 56.505 179.835 58.045 180.205 ;
        RECT 58.345 179.330 58.485 181.390 ;
        RECT 57.365 179.010 57.625 179.330 ;
        RECT 58.285 179.010 58.545 179.330 ;
        RECT 55.985 178.330 56.245 178.650 ;
        RECT 55.065 176.630 55.325 176.950 ;
        RECT 55.515 176.775 55.795 177.145 ;
        RECT 52.305 176.290 52.565 176.610 ;
        RECT 51.385 171.190 51.645 171.510 ;
        RECT 51.845 171.190 52.105 171.510 ;
        RECT 52.365 171.420 52.505 176.290 ;
        RECT 55.585 176.270 55.725 176.775 ;
        RECT 55.525 175.950 55.785 176.270 ;
        RECT 55.525 174.930 55.785 175.250 ;
        RECT 55.585 173.065 55.725 174.930 ;
        RECT 56.045 173.210 56.185 178.330 ;
        RECT 57.425 176.270 57.565 179.010 ;
        RECT 57.825 178.330 58.085 178.650 ;
        RECT 57.885 177.825 58.025 178.330 ;
        RECT 57.815 177.455 58.095 177.825 ;
        RECT 57.885 176.465 58.025 177.455 ;
        RECT 56.445 175.950 56.705 176.270 ;
        RECT 56.905 175.950 57.165 176.270 ;
        RECT 57.365 175.950 57.625 176.270 ;
        RECT 57.815 176.095 58.095 176.465 ;
        RECT 58.285 175.950 58.545 176.270 ;
        RECT 58.735 176.095 59.015 176.465 ;
        RECT 56.505 175.250 56.645 175.950 ;
        RECT 56.965 175.250 57.105 175.950 ;
        RECT 56.445 174.930 56.705 175.250 ;
        RECT 56.905 174.930 57.165 175.250 ;
        RECT 56.505 174.395 58.045 174.765 ;
        RECT 56.895 173.375 57.175 173.745 ;
        RECT 57.825 173.460 58.085 173.550 ;
        RECT 58.345 173.460 58.485 175.950 ;
        RECT 56.905 173.230 57.165 173.375 ;
        RECT 57.825 173.320 58.485 173.460 ;
        RECT 57.825 173.230 58.085 173.320 ;
        RECT 55.065 172.550 55.325 172.870 ;
        RECT 55.515 172.695 55.795 173.065 ;
        RECT 55.985 172.890 56.245 173.210 ;
        RECT 53.205 171.675 54.745 172.045 ;
        RECT 52.765 171.420 53.025 171.510 ;
        RECT 52.365 171.280 53.025 171.420 ;
        RECT 52.765 171.190 53.025 171.280 ;
        RECT 51.905 169.810 52.045 171.190 ;
        RECT 55.125 170.830 55.265 172.550 ;
        RECT 55.525 172.210 55.785 172.530 ;
        RECT 55.585 170.830 55.725 172.210 ;
        RECT 57.885 171.510 58.025 173.230 ;
        RECT 58.275 172.695 58.555 173.065 ;
        RECT 58.345 171.510 58.485 172.695 ;
        RECT 57.825 171.190 58.085 171.510 ;
        RECT 58.285 171.190 58.545 171.510 ;
        RECT 58.805 170.910 58.945 176.095 ;
        RECT 59.265 175.670 59.405 183.770 ;
        RECT 59.665 180.710 59.925 181.030 ;
        RECT 59.725 179.670 59.865 180.710 ;
        RECT 59.665 179.350 59.925 179.670 ;
        RECT 60.185 178.650 60.325 184.110 ;
        RECT 63.805 183.770 64.065 184.090 ;
        RECT 63.865 181.790 64.005 183.770 ;
        RECT 62.485 181.710 64.005 181.790 ;
        RECT 61.045 181.390 61.305 181.710 ;
        RECT 62.425 181.650 64.005 181.710 ;
        RECT 62.425 181.390 62.685 181.650 ;
        RECT 61.105 181.110 61.245 181.390 ;
        RECT 61.965 181.110 62.225 181.370 ;
        RECT 61.105 181.050 62.225 181.110 ;
        RECT 61.105 180.970 62.165 181.050 ;
        RECT 63.345 180.710 63.605 181.030 ;
        RECT 62.425 179.010 62.685 179.330 ;
        RECT 61.505 178.900 61.765 178.990 ;
        RECT 61.105 178.760 61.765 178.900 ;
        RECT 59.655 178.135 59.935 178.505 ;
        RECT 60.125 178.330 60.385 178.650 ;
        RECT 59.725 176.610 59.865 178.135 ;
        RECT 59.665 176.290 59.925 176.610 ;
        RECT 59.265 175.530 59.865 175.670 ;
        RECT 59.205 174.930 59.465 175.250 ;
        RECT 59.265 174.230 59.405 174.930 ;
        RECT 59.205 173.910 59.465 174.230 ;
        RECT 53.685 170.510 53.945 170.830 ;
        RECT 55.065 170.510 55.325 170.830 ;
        RECT 55.525 170.510 55.785 170.830 ;
        RECT 58.345 170.770 58.945 170.910 ;
        RECT 51.845 169.490 52.105 169.810 ;
        RECT 44.485 167.450 44.745 167.770 ;
        RECT 49.085 167.450 49.345 167.770 ;
        RECT 46.785 167.110 47.045 167.430 ;
        RECT 48.165 167.110 48.425 167.430 ;
        RECT 53.745 167.340 53.885 170.510 ;
        RECT 55.065 169.490 55.325 169.810 ;
        RECT 52.825 167.200 53.885 167.340 ;
        RECT 44.945 166.770 45.205 167.090 ;
        RECT 45.405 166.770 45.665 167.090 ;
        RECT 45.005 165.390 45.145 166.770 ;
        RECT 44.945 165.070 45.205 165.390 ;
        RECT 44.025 159.290 44.285 159.610 ;
        RECT 44.945 158.610 45.205 158.930 ;
        RECT 43.555 156.375 43.835 156.745 ;
        RECT 43.105 153.850 43.365 154.170 ;
        RECT 42.645 151.810 42.905 152.130 ;
        RECT 43.105 150.790 43.365 151.110 ;
        RECT 43.165 149.750 43.305 150.790 ;
        RECT 43.105 149.430 43.365 149.750 ;
        RECT 43.625 149.410 43.765 156.375 ;
        RECT 44.025 156.230 44.285 156.550 ;
        RECT 44.085 155.270 44.225 156.230 ;
        RECT 45.005 155.950 45.145 158.610 ;
        RECT 45.465 156.550 45.605 166.770 ;
        RECT 46.845 164.710 46.985 167.110 ;
        RECT 46.785 164.390 47.045 164.710 ;
        RECT 46.845 162.330 46.985 164.390 ;
        RECT 48.225 163.350 48.365 167.110 ;
        RECT 52.825 165.390 52.965 167.200 ;
        RECT 53.205 166.235 54.745 166.605 ;
        RECT 55.125 165.730 55.265 169.490 ;
        RECT 55.585 168.110 55.725 170.510 ;
        RECT 56.505 168.955 58.045 169.325 ;
        RECT 55.525 167.790 55.785 168.110 ;
        RECT 55.585 166.070 55.725 167.790 ;
        RECT 56.905 166.770 57.165 167.090 ;
        RECT 55.525 165.750 55.785 166.070 ;
        RECT 55.065 165.410 55.325 165.730 ;
        RECT 56.965 165.390 57.105 166.770 ;
        RECT 48.625 165.070 48.885 165.390 ;
        RECT 52.765 165.070 53.025 165.390 ;
        RECT 56.905 165.070 57.165 165.390 ;
        RECT 48.165 163.030 48.425 163.350 ;
        RECT 46.785 162.010 47.045 162.330 ;
        RECT 48.165 159.630 48.425 159.950 ;
        RECT 47.245 158.610 47.505 158.930 ;
        RECT 47.305 157.230 47.445 158.610 ;
        RECT 48.225 157.910 48.365 159.630 ;
        RECT 48.165 157.590 48.425 157.910 ;
        RECT 46.785 156.910 47.045 157.230 ;
        RECT 47.245 156.910 47.505 157.230 ;
        RECT 45.405 156.230 45.665 156.550 ;
        RECT 45.005 155.810 45.605 155.950 ;
        RECT 44.085 155.190 45.145 155.270 ;
        RECT 44.085 155.130 45.205 155.190 ;
        RECT 44.945 154.870 45.205 155.130 ;
        RECT 44.485 154.190 44.745 154.510 ;
        RECT 44.025 153.510 44.285 153.830 ;
        RECT 44.085 149.750 44.225 153.510 ;
        RECT 44.545 149.750 44.685 154.190 ;
        RECT 44.945 153.850 45.205 154.170 ;
        RECT 44.025 149.430 44.285 149.750 ;
        RECT 44.485 149.430 44.745 149.750 ;
        RECT 43.565 149.090 43.825 149.410 ;
        RECT 44.015 148.215 44.295 148.585 ;
        RECT 40.345 146.710 40.605 147.030 ;
        RECT 42.185 146.710 42.445 147.030 ;
        RECT 44.085 146.010 44.225 148.215 ;
        RECT 44.545 146.010 44.685 149.430 ;
        RECT 45.005 148.730 45.145 153.850 ;
        RECT 45.465 149.070 45.605 155.810 ;
        RECT 46.845 154.510 46.985 156.910 ;
        RECT 48.685 156.210 48.825 165.070 ;
        RECT 49.545 164.050 49.805 164.370 ;
        RECT 49.085 162.010 49.345 162.330 ;
        RECT 49.145 158.930 49.285 162.010 ;
        RECT 49.605 160.290 49.745 164.050 ;
        RECT 56.505 163.515 58.045 163.885 ;
        RECT 55.065 162.690 55.325 163.010 ;
        RECT 53.205 160.795 54.745 161.165 ;
        RECT 49.545 159.970 49.805 160.290 ;
        RECT 49.085 158.610 49.345 158.930 ;
        RECT 50.465 158.610 50.725 158.930 ;
        RECT 48.625 155.890 48.885 156.210 ;
        RECT 46.785 154.190 47.045 154.510 ;
        RECT 49.535 154.335 49.815 154.705 ;
        RECT 50.525 154.510 50.665 158.610 ;
        RECT 51.385 157.590 51.645 157.910 ;
        RECT 51.445 154.510 51.585 157.590 ;
        RECT 52.305 156.570 52.565 156.890 ;
        RECT 49.545 154.190 49.805 154.335 ;
        RECT 50.005 154.190 50.265 154.510 ;
        RECT 50.465 154.190 50.725 154.510 ;
        RECT 51.385 154.190 51.645 154.510 ;
        RECT 46.325 153.850 46.585 154.170 ;
        RECT 46.385 149.070 46.525 153.850 ;
        RECT 50.065 153.830 50.205 154.190 ;
        RECT 52.365 154.170 52.505 156.570 ;
        RECT 52.765 155.890 53.025 156.210 ;
        RECT 52.825 154.590 52.965 155.890 ;
        RECT 53.205 155.355 54.745 155.725 ;
        RECT 52.825 154.450 53.885 154.590 ;
        RECT 55.125 154.510 55.265 162.690 ;
        RECT 55.525 160.310 55.785 160.630 ;
        RECT 55.585 156.890 55.725 160.310 ;
        RECT 55.985 159.290 56.245 159.610 ;
        RECT 55.525 156.570 55.785 156.890 ;
        RECT 55.525 155.890 55.785 156.210 ;
        RECT 52.305 153.850 52.565 154.170 ;
        RECT 53.745 153.910 53.885 154.450 ;
        RECT 55.065 154.190 55.325 154.510 ;
        RECT 50.005 153.510 50.265 153.830 ;
        RECT 52.765 153.510 53.025 153.830 ;
        RECT 53.745 153.770 55.265 153.910 ;
        RECT 46.785 153.170 47.045 153.490 ;
        RECT 46.845 151.790 46.985 153.170 ;
        RECT 46.785 151.470 47.045 151.790 ;
        RECT 48.625 151.130 48.885 151.450 ;
        RECT 47.245 150.450 47.505 150.770 ;
        RECT 47.305 149.070 47.445 150.450 ;
        RECT 45.405 148.750 45.665 149.070 ;
        RECT 46.325 148.750 46.585 149.070 ;
        RECT 47.245 148.750 47.505 149.070 ;
        RECT 44.945 148.410 45.205 148.730 ;
        RECT 48.685 148.390 48.825 151.130 ;
        RECT 48.625 148.070 48.885 148.390 ;
        RECT 44.025 145.690 44.285 146.010 ;
        RECT 44.485 145.690 44.745 146.010 ;
        RECT 50.925 145.010 51.185 145.330 ;
        RECT 51.845 145.010 52.105 145.330 ;
        RECT 52.305 145.010 52.565 145.330 ;
        RECT 43.565 143.990 43.825 144.310 ;
        RECT 42.175 140.735 42.455 141.105 ;
        RECT 39.425 140.250 39.685 140.570 ;
        RECT 41.725 140.250 41.985 140.570 ;
        RECT 39.485 138.870 39.625 140.250 ;
        RECT 40.805 139.570 41.065 139.890 ;
        RECT 38.965 138.550 39.225 138.870 ;
        RECT 39.425 138.550 39.685 138.870 ;
        RECT 39.025 138.385 39.165 138.550 ;
        RECT 38.955 138.015 39.235 138.385 ;
        RECT 38.045 134.900 38.705 135.040 ;
        RECT 38.045 134.810 38.305 134.900 ;
        RECT 38.045 134.130 38.305 134.450 ;
        RECT 39.425 134.130 39.685 134.450 ;
        RECT 38.105 132.750 38.245 134.130 ;
        RECT 39.485 133.430 39.625 134.130 ;
        RECT 38.505 133.110 38.765 133.430 ;
        RECT 39.425 133.110 39.685 133.430 ;
        RECT 38.565 132.750 38.705 133.110 ;
        RECT 38.045 132.430 38.305 132.750 ;
        RECT 38.505 132.660 38.765 132.750 ;
        RECT 38.505 132.520 39.165 132.660 ;
        RECT 38.505 132.430 38.765 132.520 ;
        RECT 37.585 132.090 37.845 132.410 ;
        RECT 37.125 131.750 37.385 132.070 ;
        RECT 36.665 129.710 36.925 130.030 ;
        RECT 36.655 126.455 36.935 126.825 ;
        RECT 36.725 124.590 36.865 126.455 ;
        RECT 37.185 124.590 37.325 131.750 ;
        RECT 37.645 127.310 37.785 132.090 ;
        RECT 38.105 127.650 38.245 132.430 ;
        RECT 39.025 127.990 39.165 132.520 ;
        RECT 38.965 127.670 39.225 127.990 ;
        RECT 38.045 127.560 38.305 127.650 ;
        RECT 38.045 127.420 38.705 127.560 ;
        RECT 38.045 127.330 38.305 127.420 ;
        RECT 37.585 126.990 37.845 127.310 ;
        RECT 38.045 126.650 38.305 126.970 ;
        RECT 36.665 124.270 36.925 124.590 ;
        RECT 37.125 124.270 37.385 124.590 ;
        RECT 36.205 123.930 36.465 124.250 ;
        RECT 35.285 123.590 35.545 123.910 ;
        RECT 35.745 123.590 36.005 123.910 ;
        RECT 34.815 121.695 35.095 122.065 ;
        RECT 34.885 119.150 35.025 121.695 ;
        RECT 35.345 121.530 35.485 123.590 ;
        RECT 38.105 123.570 38.245 126.650 ;
        RECT 36.665 123.250 36.925 123.570 ;
        RECT 38.045 123.250 38.305 123.570 ;
        RECT 35.285 121.210 35.545 121.530 ;
        RECT 34.825 118.830 35.085 119.150 ;
        RECT 36.195 118.975 36.475 119.345 ;
        RECT 36.265 118.810 36.405 118.975 ;
        RECT 36.205 118.490 36.465 118.810 ;
        RECT 35.745 117.810 36.005 118.130 ;
        RECT 35.275 116.935 35.555 117.305 ;
        RECT 35.345 116.770 35.485 116.935 ;
        RECT 35.285 116.450 35.545 116.770 ;
        RECT 34.825 115.770 35.085 116.090 ;
        RECT 34.885 111.670 35.025 115.770 ;
        RECT 35.275 115.575 35.555 115.945 ;
        RECT 35.345 114.390 35.485 115.575 ;
        RECT 35.285 114.070 35.545 114.390 ;
        RECT 35.345 113.370 35.485 114.070 ;
        RECT 35.285 113.050 35.545 113.370 ;
        RECT 34.825 111.350 35.085 111.670 ;
        RECT 34.365 111.010 34.625 111.330 ;
        RECT 35.805 110.990 35.945 117.810 ;
        RECT 36.725 116.430 36.865 123.250 ;
        RECT 38.045 122.230 38.305 122.550 ;
        RECT 37.585 119.170 37.845 119.490 ;
        RECT 36.665 116.110 36.925 116.430 ;
        RECT 36.665 115.090 36.925 115.410 ;
        RECT 36.725 111.330 36.865 115.090 ;
        RECT 37.645 113.790 37.785 119.170 ;
        RECT 38.105 118.810 38.245 122.230 ;
        RECT 38.565 119.345 38.705 127.420 ;
        RECT 40.345 127.330 40.605 127.650 ;
        RECT 39.425 126.990 39.685 127.310 ;
        RECT 39.485 126.630 39.625 126.990 ;
        RECT 39.425 126.310 39.685 126.630 ;
        RECT 39.425 124.610 39.685 124.930 ;
        RECT 38.495 118.975 38.775 119.345 ;
        RECT 39.485 119.230 39.625 124.610 ;
        RECT 38.965 118.830 39.225 119.150 ;
        RECT 39.485 119.090 40.085 119.230 ;
        RECT 38.045 118.490 38.305 118.810 ;
        RECT 39.025 116.770 39.165 118.830 ;
        RECT 38.965 116.450 39.225 116.770 ;
        RECT 38.505 116.110 38.765 116.430 ;
        RECT 37.645 113.650 38.245 113.790 ;
        RECT 37.585 113.225 37.845 113.370 ;
        RECT 37.575 112.855 37.855 113.225 ;
        RECT 36.665 111.010 36.925 111.330 ;
        RECT 33.445 110.670 33.705 110.990 ;
        RECT 35.745 110.670 36.005 110.990 ;
        RECT 33.045 110.250 33.645 110.390 ;
        RECT 33.505 109.970 33.645 110.250 ;
        RECT 32.985 109.650 33.245 109.970 ;
        RECT 33.445 109.650 33.705 109.970 ;
        RECT 37.645 109.710 37.785 112.855 ;
        RECT 38.105 112.690 38.245 113.650 ;
        RECT 38.565 113.370 38.705 116.110 ;
        RECT 39.425 115.770 39.685 116.090 ;
        RECT 38.965 115.430 39.225 115.750 ;
        RECT 39.025 113.370 39.165 115.430 ;
        RECT 39.485 113.370 39.625 115.770 ;
        RECT 38.505 113.050 38.765 113.370 ;
        RECT 38.965 113.050 39.225 113.370 ;
        RECT 39.425 113.050 39.685 113.370 ;
        RECT 39.945 112.690 40.085 119.090 ;
        RECT 40.405 114.050 40.545 127.330 ;
        RECT 40.345 113.730 40.605 114.050 ;
        RECT 38.045 112.370 38.305 112.690 ;
        RECT 39.885 112.370 40.145 112.690 ;
        RECT 40.865 111.670 41.005 139.570 ;
        RECT 41.785 138.530 41.925 140.250 ;
        RECT 41.725 138.210 41.985 138.530 ;
        RECT 41.265 136.850 41.525 137.170 ;
        RECT 41.325 136.150 41.465 136.850 ;
        RECT 41.265 135.830 41.525 136.150 ;
        RECT 42.245 135.470 42.385 140.735 ;
        RECT 43.625 140.570 43.765 143.990 ;
        RECT 45.865 142.350 46.125 142.610 ;
        RECT 45.865 142.290 46.525 142.350 ;
        RECT 45.925 142.210 46.525 142.290 ;
        RECT 45.865 140.590 46.125 140.910 ;
        RECT 43.105 140.250 43.365 140.570 ;
        RECT 43.565 140.250 43.825 140.570 ;
        RECT 44.485 140.250 44.745 140.570 ;
        RECT 43.165 138.870 43.305 140.250 ;
        RECT 43.105 138.550 43.365 138.870 ;
        RECT 44.025 138.550 44.285 138.870 ;
        RECT 42.645 138.210 42.905 138.530 ;
        RECT 42.705 137.170 42.845 138.210 ;
        RECT 43.555 138.015 43.835 138.385 ;
        RECT 43.565 137.870 43.825 138.015 ;
        RECT 42.645 136.850 42.905 137.170 ;
        RECT 43.105 136.850 43.365 137.170 ;
        RECT 42.185 135.150 42.445 135.470 ;
        RECT 42.705 134.790 42.845 136.850 ;
        RECT 42.645 134.470 42.905 134.790 ;
        RECT 42.185 134.130 42.445 134.450 ;
        RECT 41.265 132.430 41.525 132.750 ;
        RECT 41.325 127.310 41.465 132.430 ;
        RECT 41.725 130.390 41.985 130.710 ;
        RECT 41.785 127.310 41.925 130.390 ;
        RECT 41.265 126.990 41.525 127.310 ;
        RECT 41.725 126.990 41.985 127.310 ;
        RECT 41.325 121.530 41.465 126.990 ;
        RECT 41.265 121.210 41.525 121.530 ;
        RECT 41.325 116.430 41.465 121.210 ;
        RECT 41.265 116.110 41.525 116.430 ;
        RECT 41.785 115.750 41.925 126.990 ;
        RECT 41.725 115.430 41.985 115.750 ;
        RECT 41.265 113.390 41.525 113.710 ;
        RECT 40.805 111.350 41.065 111.670 ;
        RECT 39.885 111.010 40.145 111.330 ;
        RECT 39.945 110.310 40.085 111.010 ;
        RECT 39.885 109.990 40.145 110.310 ;
        RECT 33.045 108.950 33.185 109.650 ;
        RECT 36.265 109.570 37.785 109.710 ;
        RECT 38.045 109.650 38.305 109.970 ;
        RECT 32.985 108.630 33.245 108.950 ;
        RECT 30.225 108.290 30.485 108.610 ;
        RECT 36.265 108.270 36.405 109.570 ;
        RECT 36.205 107.950 36.465 108.270 ;
        RECT 38.105 107.930 38.245 109.650 ;
        RECT 41.325 108.270 41.465 113.390 ;
        RECT 41.725 113.280 41.985 113.370 ;
        RECT 42.245 113.280 42.385 134.130 ;
        RECT 42.705 125.270 42.845 134.470 ;
        RECT 42.645 124.950 42.905 125.270 ;
        RECT 42.705 123.990 42.845 124.950 ;
        RECT 43.165 124.590 43.305 136.850 ;
        RECT 44.085 135.130 44.225 138.550 ;
        RECT 44.545 138.530 44.685 140.250 ;
        RECT 45.925 138.870 46.065 140.590 ;
        RECT 46.385 140.230 46.525 142.210 ;
        RECT 46.785 140.930 47.045 141.250 ;
        RECT 46.325 139.910 46.585 140.230 ;
        RECT 45.865 138.550 46.125 138.870 ;
        RECT 44.485 138.210 44.745 138.530 ;
        RECT 45.925 138.190 46.065 138.550 ;
        RECT 45.405 137.870 45.665 138.190 ;
        RECT 45.865 137.870 46.125 138.190 ;
        RECT 45.465 136.150 45.605 137.870 ;
        RECT 45.405 135.830 45.665 136.150 ;
        RECT 44.025 134.810 44.285 135.130 ;
        RECT 44.945 135.040 45.205 135.130 ;
        RECT 46.325 135.040 46.585 135.130 ;
        RECT 44.945 134.900 46.585 135.040 ;
        RECT 44.945 134.810 45.205 134.900 ;
        RECT 46.325 134.810 46.585 134.900 ;
        RECT 46.845 134.790 46.985 140.930 ;
        RECT 50.985 139.890 51.125 145.010 ;
        RECT 50.925 139.570 51.185 139.890 ;
        RECT 51.905 138.870 52.045 145.010 ;
        RECT 52.365 140.910 52.505 145.010 ;
        RECT 52.825 140.910 52.965 153.510 ;
        RECT 54.145 153.170 54.405 153.490 ;
        RECT 54.205 151.450 54.345 153.170 ;
        RECT 54.145 151.130 54.405 151.450 ;
        RECT 53.205 149.915 54.745 150.285 ;
        RECT 55.125 146.010 55.265 153.770 ;
        RECT 55.585 151.450 55.725 155.890 ;
        RECT 56.045 155.190 56.185 159.290 ;
        RECT 56.505 158.075 58.045 158.445 ;
        RECT 58.345 156.890 58.485 170.770 ;
        RECT 58.745 170.170 59.005 170.490 ;
        RECT 58.805 167.430 58.945 170.170 ;
        RECT 59.265 167.430 59.405 173.910 ;
        RECT 59.725 172.870 59.865 175.530 ;
        RECT 60.125 175.270 60.385 175.590 ;
        RECT 60.185 173.745 60.325 175.270 ;
        RECT 60.585 174.930 60.845 175.250 ;
        RECT 60.645 174.230 60.785 174.930 ;
        RECT 60.585 173.910 60.845 174.230 ;
        RECT 60.115 173.375 60.395 173.745 ;
        RECT 59.665 172.550 59.925 172.870 ;
        RECT 59.665 170.850 59.925 171.170 ;
        RECT 59.725 168.790 59.865 170.850 ;
        RECT 59.665 168.470 59.925 168.790 ;
        RECT 60.185 168.110 60.325 173.375 ;
        RECT 60.125 167.790 60.385 168.110 ;
        RECT 58.745 167.110 59.005 167.430 ;
        RECT 59.205 167.110 59.465 167.430 ;
        RECT 58.805 165.050 58.945 167.110 ;
        RECT 58.745 164.730 59.005 165.050 ;
        RECT 58.805 161.990 58.945 164.730 ;
        RECT 60.185 163.350 60.325 167.790 ;
        RECT 60.645 165.585 60.785 173.910 ;
        RECT 61.105 173.890 61.245 178.760 ;
        RECT 61.505 178.670 61.765 178.760 ;
        RECT 61.965 177.990 62.225 178.310 ;
        RECT 61.045 173.570 61.305 173.890 ;
        RECT 61.045 172.890 61.305 173.210 ;
        RECT 61.105 170.490 61.245 172.890 ;
        RECT 61.045 170.170 61.305 170.490 ;
        RECT 62.025 167.770 62.165 177.990 ;
        RECT 62.485 172.950 62.625 179.010 ;
        RECT 63.405 178.990 63.545 180.710 ;
        RECT 63.345 178.670 63.605 178.990 ;
        RECT 63.865 178.310 64.005 181.650 ;
        RECT 66.625 181.370 66.765 188.530 ;
        RECT 66.565 181.050 66.825 181.370 ;
        RECT 64.265 178.330 64.525 178.650 ;
        RECT 66.105 178.330 66.365 178.650 ;
        RECT 63.805 177.990 64.065 178.310 ;
        RECT 64.325 177.145 64.465 178.330 ;
        RECT 64.725 177.650 64.985 177.970 ;
        RECT 65.185 177.825 65.445 177.970 ;
        RECT 64.255 176.775 64.535 177.145 ;
        RECT 62.885 174.930 63.145 175.250 ;
        RECT 62.945 173.550 63.085 174.930 ;
        RECT 62.885 173.230 63.145 173.550 ;
        RECT 62.485 172.810 63.085 172.950 ;
        RECT 64.785 172.870 64.925 177.650 ;
        RECT 65.175 177.455 65.455 177.825 ;
        RECT 66.165 176.950 66.305 178.330 ;
        RECT 67.085 176.950 67.225 189.550 ;
        RECT 72.085 188.530 72.345 188.850 ;
        RECT 71.165 187.170 71.425 187.490 ;
        RECT 70.245 186.490 70.505 186.810 ;
        RECT 70.305 184.770 70.445 186.490 ;
        RECT 71.225 185.110 71.365 187.170 ;
        RECT 71.165 184.790 71.425 185.110 ;
        RECT 70.245 184.450 70.505 184.770 ;
        RECT 72.145 183.750 72.285 188.530 ;
        RECT 72.545 187.510 72.805 187.830 ;
        RECT 72.085 183.430 72.345 183.750 ;
        RECT 67.945 183.090 68.205 183.410 ;
        RECT 68.005 182.610 68.145 183.090 ;
        RECT 68.005 182.470 68.605 182.610 ;
        RECT 68.465 182.050 68.605 182.470 ;
        RECT 71.625 182.070 71.885 182.390 ;
        RECT 68.405 181.730 68.665 182.050 ;
        RECT 71.685 181.710 71.825 182.070 ;
        RECT 72.605 181.710 72.745 187.510 ;
        RECT 74.445 186.810 74.585 189.890 ;
        RECT 76.285 189.870 76.425 194.340 ;
        RECT 76.225 189.550 76.485 189.870 ;
        RECT 76.685 189.210 76.945 189.530 ;
        RECT 76.745 187.830 76.885 189.210 ;
        RECT 78.985 188.530 79.245 188.850 ;
        RECT 76.685 187.510 76.945 187.830 ;
        RECT 79.045 187.150 79.185 188.530 ;
        RECT 79.505 187.490 79.645 194.340 ;
        RECT 82.725 192.250 82.865 194.340 ;
        RECT 92.075 193.435 93.615 193.805 ;
        RECT 88.185 192.610 88.445 192.930 ;
        RECT 87.725 192.270 87.985 192.590 ;
        RECT 82.665 191.930 82.925 192.250 ;
        RECT 86.805 191.930 87.065 192.250 ;
        RECT 83.585 191.250 83.845 191.570 ;
        RECT 83.645 189.870 83.785 191.250 ;
        RECT 82.205 189.550 82.465 189.870 ;
        RECT 83.585 189.550 83.845 189.870 ;
        RECT 81.745 187.510 82.005 187.830 ;
        RECT 79.445 187.170 79.705 187.490 ;
        RECT 78.985 186.830 79.245 187.150 ;
        RECT 74.385 186.490 74.645 186.810 ;
        RECT 74.445 184.430 74.585 186.490 ;
        RECT 78.065 186.150 78.325 186.470 ;
        RECT 75.765 185.810 76.025 186.130 ;
        RECT 75.825 184.430 75.965 185.810 ;
        RECT 73.005 184.110 73.265 184.430 ;
        RECT 74.385 184.110 74.645 184.430 ;
        RECT 75.765 184.110 76.025 184.430 ;
        RECT 73.065 183.410 73.205 184.110 ;
        RECT 73.005 183.090 73.265 183.410 ;
        RECT 73.065 182.610 73.205 183.090 ;
        RECT 74.445 182.610 74.585 184.110 ;
        RECT 78.125 184.090 78.265 186.150 ;
        RECT 78.065 183.770 78.325 184.090 ;
        RECT 73.065 182.470 73.665 182.610 ;
        RECT 71.625 181.390 71.885 181.710 ;
        RECT 72.545 181.390 72.805 181.710 ;
        RECT 68.865 181.050 69.125 181.370 ;
        RECT 68.925 179.670 69.065 181.050 ;
        RECT 70.705 180.370 70.965 180.690 ;
        RECT 68.865 179.350 69.125 179.670 ;
        RECT 70.245 178.670 70.505 178.990 ;
        RECT 66.105 176.630 66.365 176.950 ;
        RECT 67.025 176.630 67.285 176.950 ;
        RECT 70.305 176.270 70.445 178.670 ;
        RECT 67.945 175.950 68.205 176.270 ;
        RECT 70.245 175.950 70.505 176.270 ;
        RECT 68.005 173.890 68.145 175.950 ;
        RECT 70.765 175.250 70.905 180.370 ;
        RECT 71.165 179.350 71.425 179.670 ;
        RECT 71.225 178.650 71.365 179.350 ;
        RECT 71.165 178.330 71.425 178.650 ;
        RECT 71.685 177.145 71.825 181.390 ;
        RECT 72.085 178.330 72.345 178.650 ;
        RECT 72.145 177.970 72.285 178.330 ;
        RECT 72.085 177.650 72.345 177.970 ;
        RECT 71.615 176.775 71.895 177.145 ;
        RECT 71.165 175.950 71.425 176.270 ;
        RECT 72.085 175.950 72.345 176.270 ;
        RECT 71.225 175.785 71.365 175.950 ;
        RECT 71.155 175.415 71.435 175.785 ;
        RECT 70.705 174.930 70.965 175.250 ;
        RECT 72.145 174.230 72.285 175.950 ;
        RECT 72.545 174.930 72.805 175.250 ;
        RECT 72.085 173.910 72.345 174.230 ;
        RECT 67.945 173.570 68.205 173.890 ;
        RECT 72.605 173.210 72.745 174.930 ;
        RECT 72.545 172.890 72.805 173.210 ;
        RECT 62.425 172.210 62.685 172.530 ;
        RECT 62.485 170.830 62.625 172.210 ;
        RECT 62.425 170.510 62.685 170.830 ;
        RECT 61.965 167.450 62.225 167.770 ;
        RECT 60.575 165.215 60.855 165.585 ;
        RECT 60.125 163.030 60.385 163.350 ;
        RECT 59.205 162.185 59.465 162.330 ;
        RECT 58.745 161.670 59.005 161.990 ;
        RECT 59.195 161.815 59.475 162.185 ;
        RECT 59.665 162.010 59.925 162.330 ;
        RECT 59.205 161.330 59.465 161.650 ;
        RECT 58.745 157.590 59.005 157.910 ;
        RECT 57.825 156.570 58.085 156.890 ;
        RECT 58.285 156.570 58.545 156.890 ;
        RECT 56.445 156.230 56.705 156.550 ;
        RECT 55.985 154.870 56.245 155.190 ;
        RECT 56.505 153.830 56.645 156.230 ;
        RECT 56.445 153.510 56.705 153.830 ;
        RECT 57.885 153.490 58.025 156.570 ;
        RECT 58.345 154.705 58.485 156.570 ;
        RECT 58.275 154.335 58.555 154.705 ;
        RECT 58.805 154.510 58.945 157.590 ;
        RECT 59.265 156.890 59.405 161.330 ;
        RECT 59.725 160.290 59.865 162.010 ;
        RECT 60.125 161.670 60.385 161.990 ;
        RECT 59.665 159.970 59.925 160.290 ;
        RECT 60.185 159.610 60.325 161.670 ;
        RECT 60.125 159.290 60.385 159.610 ;
        RECT 60.185 157.570 60.325 159.290 ;
        RECT 60.645 157.910 60.785 165.215 ;
        RECT 61.045 164.050 61.305 164.370 ;
        RECT 61.105 163.010 61.245 164.050 ;
        RECT 61.045 162.690 61.305 163.010 ;
        RECT 60.585 157.590 60.845 157.910 ;
        RECT 60.125 157.250 60.385 157.570 ;
        RECT 59.205 156.570 59.465 156.890 ;
        RECT 59.665 156.230 59.925 156.550 ;
        RECT 59.725 154.510 59.865 156.230 ;
        RECT 58.745 154.190 59.005 154.510 ;
        RECT 59.665 154.190 59.925 154.510 ;
        RECT 59.725 154.025 59.865 154.190 ;
        RECT 59.655 153.655 59.935 154.025 ;
        RECT 57.825 153.170 58.085 153.490 ;
        RECT 56.505 152.635 58.045 153.005 ;
        RECT 56.905 151.470 57.165 151.790 ;
        RECT 55.525 151.130 55.785 151.450 ;
        RECT 55.985 149.090 56.245 149.410 ;
        RECT 56.045 147.030 56.185 149.090 ;
        RECT 56.965 148.730 57.105 151.470 ;
        RECT 57.365 150.450 57.625 150.770 ;
        RECT 59.665 150.450 59.925 150.770 ;
        RECT 57.425 149.750 57.565 150.450 ;
        RECT 57.365 149.430 57.625 149.750 ;
        RECT 59.725 149.070 59.865 150.450 ;
        RECT 60.185 149.070 60.325 157.250 ;
        RECT 60.585 156.570 60.845 156.890 ;
        RECT 60.645 154.510 60.785 156.570 ;
        RECT 60.585 154.190 60.845 154.510 ;
        RECT 60.645 151.110 60.785 154.190 ;
        RECT 60.585 150.790 60.845 151.110 ;
        RECT 59.665 148.750 59.925 149.070 ;
        RECT 60.125 148.750 60.385 149.070 ;
        RECT 56.905 148.410 57.165 148.730 ;
        RECT 56.505 147.195 58.045 147.565 ;
        RECT 55.985 146.710 56.245 147.030 ;
        RECT 60.125 146.370 60.385 146.690 ;
        RECT 55.065 145.690 55.325 146.010 ;
        RECT 53.205 144.475 54.745 144.845 ;
        RECT 59.205 143.990 59.465 144.310 ;
        RECT 54.605 142.970 54.865 143.290 ;
        RECT 58.285 142.970 58.545 143.290 ;
        RECT 54.665 141.590 54.805 142.970 ;
        RECT 56.505 141.755 58.045 142.125 ;
        RECT 54.605 141.270 54.865 141.590 ;
        RECT 52.305 140.590 52.565 140.910 ;
        RECT 52.765 140.590 53.025 140.910 ;
        RECT 58.345 140.230 58.485 142.970 ;
        RECT 58.745 142.290 59.005 142.610 ;
        RECT 58.285 139.910 58.545 140.230 ;
        RECT 53.205 139.035 54.745 139.405 ;
        RECT 51.845 138.550 52.105 138.870 ;
        RECT 51.905 135.130 52.045 138.550 ;
        RECT 55.125 138.190 56.185 138.270 ;
        RECT 55.125 138.130 56.245 138.190 ;
        RECT 55.125 137.850 55.265 138.130 ;
        RECT 55.985 137.870 56.245 138.130 ;
        RECT 58.345 137.850 58.485 139.910 ;
        RECT 58.805 138.190 58.945 142.290 ;
        RECT 59.265 140.570 59.405 143.990 ;
        RECT 59.665 142.970 59.925 143.290 ;
        RECT 59.725 140.570 59.865 142.970 ;
        RECT 60.185 140.910 60.325 146.370 ;
        RECT 61.105 145.670 61.245 162.690 ;
        RECT 62.025 162.185 62.165 167.450 ;
        RECT 62.425 163.030 62.685 163.350 ;
        RECT 62.485 162.670 62.625 163.030 ;
        RECT 62.425 162.350 62.685 162.670 ;
        RECT 61.955 161.815 62.235 162.185 ;
        RECT 61.505 155.890 61.765 156.210 ;
        RECT 61.565 152.130 61.705 155.890 ;
        RECT 61.505 151.810 61.765 152.130 ;
        RECT 61.505 151.130 61.765 151.450 ;
        RECT 61.565 148.585 61.705 151.130 ;
        RECT 62.025 149.070 62.165 161.815 ;
        RECT 62.485 153.910 62.625 162.350 ;
        RECT 62.945 154.760 63.085 172.810 ;
        RECT 64.725 172.550 64.985 172.870 ;
        RECT 70.245 172.550 70.505 172.870 ;
        RECT 64.265 172.210 64.525 172.530 ;
        RECT 63.345 169.490 63.605 169.810 ;
        RECT 63.405 165.470 63.545 169.490 ;
        RECT 64.325 166.070 64.465 172.210 ;
        RECT 70.305 171.510 70.445 172.550 ;
        RECT 70.245 171.190 70.505 171.510 ;
        RECT 67.945 170.510 68.205 170.830 ;
        RECT 67.025 170.170 67.285 170.490 ;
        RECT 67.085 168.110 67.225 170.170 ;
        RECT 67.025 167.790 67.285 168.110 ;
        RECT 64.725 166.770 64.985 167.090 ;
        RECT 64.265 165.750 64.525 166.070 ;
        RECT 64.785 165.730 64.925 166.770 ;
        RECT 63.405 165.330 64.465 165.470 ;
        RECT 64.725 165.410 64.985 165.730 ;
        RECT 63.345 156.745 63.605 156.890 ;
        RECT 63.335 156.375 63.615 156.745 ;
        RECT 62.945 154.620 63.545 154.760 ;
        RECT 62.485 153.770 63.085 153.910 ;
        RECT 62.425 153.170 62.685 153.490 ;
        RECT 62.485 151.450 62.625 153.170 ;
        RECT 62.425 151.130 62.685 151.450 ;
        RECT 61.965 148.750 62.225 149.070 ;
        RECT 61.495 148.215 61.775 148.585 ;
        RECT 62.945 146.690 63.085 153.770 ;
        RECT 63.405 151.110 63.545 154.620 ;
        RECT 63.345 150.790 63.605 151.110 ;
        RECT 63.795 148.895 64.075 149.265 ;
        RECT 62.885 146.370 63.145 146.690 ;
        RECT 61.045 145.350 61.305 145.670 ;
        RECT 60.125 140.590 60.385 140.910 ;
        RECT 59.205 140.250 59.465 140.570 ;
        RECT 59.665 140.250 59.925 140.570 ;
        RECT 59.205 139.570 59.465 139.890 ;
        RECT 59.265 138.870 59.405 139.570 ;
        RECT 59.725 138.950 59.865 140.250 ;
        RECT 59.205 138.550 59.465 138.870 ;
        RECT 59.725 138.810 60.325 138.950 ;
        RECT 60.185 138.190 60.325 138.810 ;
        RECT 58.745 137.870 59.005 138.190 ;
        RECT 59.205 137.870 59.465 138.190 ;
        RECT 60.125 137.870 60.385 138.190 ;
        RECT 55.065 137.530 55.325 137.850 ;
        RECT 55.525 137.530 55.785 137.850 ;
        RECT 58.285 137.530 58.545 137.850 ;
        RECT 54.605 136.850 54.865 137.170 ;
        RECT 54.665 136.150 54.805 136.850 ;
        RECT 55.585 136.150 55.725 137.530 ;
        RECT 56.505 136.315 58.045 136.685 ;
        RECT 54.605 135.830 54.865 136.150 ;
        RECT 55.525 135.830 55.785 136.150 ;
        RECT 53.225 135.490 53.485 135.810 ;
        RECT 51.845 134.810 52.105 135.130 ;
        RECT 53.285 134.870 53.425 135.490 ;
        RECT 57.365 135.150 57.625 135.470 ;
        RECT 54.595 134.870 54.875 134.985 ;
        RECT 46.785 134.470 47.045 134.790 ;
        RECT 53.285 134.730 54.875 134.870 ;
        RECT 54.595 134.615 54.875 134.730 ;
        RECT 53.205 133.595 54.745 133.965 ;
        RECT 57.425 133.090 57.565 135.150 ;
        RECT 44.025 132.770 44.285 133.090 ;
        RECT 51.845 132.770 52.105 133.090 ;
        RECT 55.525 132.770 55.785 133.090 ;
        RECT 57.365 132.770 57.625 133.090 ;
        RECT 43.565 131.410 43.825 131.730 ;
        RECT 43.625 127.650 43.765 131.410 ;
        RECT 43.565 127.330 43.825 127.650 ;
        RECT 44.085 127.310 44.225 132.770 ;
        RECT 45.865 132.430 46.125 132.750 ;
        RECT 45.925 130.710 46.065 132.430 ;
        RECT 45.865 130.390 46.125 130.710 ;
        RECT 48.625 130.050 48.885 130.370 ;
        RECT 47.705 129.030 47.965 129.350 ;
        RECT 44.025 126.990 44.285 127.310 ;
        RECT 47.245 126.990 47.505 127.310 ;
        RECT 43.105 124.270 43.365 124.590 ;
        RECT 42.705 123.850 43.305 123.990 ;
        RECT 42.645 121.550 42.905 121.870 ;
        RECT 42.705 117.110 42.845 121.550 ;
        RECT 43.165 119.830 43.305 123.850 ;
        RECT 43.105 119.510 43.365 119.830 ;
        RECT 43.565 117.810 43.825 118.130 ;
        RECT 43.625 117.110 43.765 117.810 ;
        RECT 44.085 117.110 44.225 126.990 ;
        RECT 44.945 126.650 45.205 126.970 ;
        RECT 44.485 123.250 44.745 123.570 ;
        RECT 44.545 122.550 44.685 123.250 ;
        RECT 44.485 122.230 44.745 122.550 ;
        RECT 45.005 121.870 45.145 126.650 ;
        RECT 45.405 125.970 45.665 126.290 ;
        RECT 45.465 124.590 45.605 125.970 ;
        RECT 45.405 124.270 45.665 124.590 ;
        RECT 45.405 122.230 45.665 122.550 ;
        RECT 46.785 122.230 47.045 122.550 ;
        RECT 44.945 121.550 45.205 121.870 ;
        RECT 45.465 118.130 45.605 122.230 ;
        RECT 45.405 117.810 45.665 118.130 ;
        RECT 42.645 116.790 42.905 117.110 ;
        RECT 43.565 116.790 43.825 117.110 ;
        RECT 44.025 116.790 44.285 117.110 ;
        RECT 45.465 116.090 45.605 117.810 ;
        RECT 46.845 116.430 46.985 122.230 ;
        RECT 47.305 119.150 47.445 126.990 ;
        RECT 47.765 124.250 47.905 129.030 ;
        RECT 48.685 124.590 48.825 130.050 ;
        RECT 51.905 127.990 52.045 132.770 ;
        RECT 52.765 130.390 53.025 130.710 ;
        RECT 52.305 129.710 52.565 130.030 ;
        RECT 51.845 127.670 52.105 127.990 ;
        RECT 52.365 127.650 52.505 129.710 ;
        RECT 52.305 127.330 52.565 127.650 ;
        RECT 51.385 126.310 51.645 126.630 ;
        RECT 48.625 124.270 48.885 124.590 ;
        RECT 47.705 123.930 47.965 124.250 ;
        RECT 50.925 122.230 51.185 122.550 ;
        RECT 49.085 120.530 49.345 120.850 ;
        RECT 47.245 118.830 47.505 119.150 ;
        RECT 46.785 116.110 47.045 116.430 ;
        RECT 45.405 115.770 45.665 116.090 ;
        RECT 41.725 113.140 42.385 113.280 ;
        RECT 41.725 113.050 41.985 113.140 ;
        RECT 46.785 113.050 47.045 113.370 ;
        RECT 45.405 112.710 45.665 113.030 ;
        RECT 41.725 112.370 41.985 112.690 ;
        RECT 42.185 112.370 42.445 112.690 ;
        RECT 42.645 112.370 42.905 112.690 ;
        RECT 44.485 112.370 44.745 112.690 ;
        RECT 41.785 111.670 41.925 112.370 ;
        RECT 41.725 111.350 41.985 111.670 ;
        RECT 42.245 109.970 42.385 112.370 ;
        RECT 42.705 110.650 42.845 112.370 ;
        RECT 44.545 110.990 44.685 112.370 ;
        RECT 45.465 111.670 45.605 112.710 ;
        RECT 46.845 111.670 46.985 113.050 ;
        RECT 45.405 111.350 45.665 111.670 ;
        RECT 46.785 111.350 47.045 111.670 ;
        RECT 44.485 110.670 44.745 110.990 ;
        RECT 42.645 110.330 42.905 110.650 ;
        RECT 42.185 109.650 42.445 109.970 ;
        RECT 41.265 107.950 41.525 108.270 ;
        RECT 24.245 107.610 24.505 107.930 ;
        RECT 36.665 107.670 36.925 107.930 ;
        RECT 38.045 107.670 38.305 107.930 ;
        RECT 36.665 107.610 38.305 107.670 ;
        RECT 36.725 107.530 38.245 107.610 ;
        RECT 41.325 107.590 41.465 107.950 ;
        RECT 42.705 107.590 42.845 110.330 ;
        RECT 46.845 108.950 46.985 111.350 ;
        RECT 47.305 110.650 47.445 118.830 ;
        RECT 49.145 118.470 49.285 120.530 ;
        RECT 50.465 119.510 50.725 119.830 ;
        RECT 49.085 118.150 49.345 118.470 ;
        RECT 50.525 116.430 50.665 119.510 ;
        RECT 50.985 116.770 51.125 122.230 ;
        RECT 51.445 121.530 51.585 126.310 ;
        RECT 51.385 121.210 51.645 121.530 ;
        RECT 51.845 121.210 52.105 121.530 ;
        RECT 51.905 119.830 52.045 121.210 ;
        RECT 51.845 119.510 52.105 119.830 ;
        RECT 52.365 119.230 52.505 127.330 ;
        RECT 52.825 126.970 52.965 130.390 ;
        RECT 53.205 128.155 54.745 128.525 ;
        RECT 55.585 127.990 55.725 132.770 ;
        RECT 58.345 132.410 58.485 137.530 ;
        RECT 59.265 135.470 59.405 137.870 ;
        RECT 60.125 136.850 60.385 137.170 ;
        RECT 59.205 135.150 59.465 135.470 ;
        RECT 58.735 132.575 59.015 132.945 ;
        RECT 56.445 132.320 56.705 132.410 ;
        RECT 56.045 132.180 56.705 132.320 ;
        RECT 56.045 129.690 56.185 132.180 ;
        RECT 56.445 132.090 56.705 132.180 ;
        RECT 58.285 132.090 58.545 132.410 ;
        RECT 56.505 130.875 58.045 131.245 ;
        RECT 55.985 129.370 56.245 129.690 ;
        RECT 55.525 127.670 55.785 127.990 ;
        RECT 56.045 127.650 56.185 129.370 ;
        RECT 55.985 127.330 56.245 127.650 ;
        RECT 52.765 126.650 53.025 126.970 ;
        RECT 53.215 126.455 53.495 126.825 ;
        RECT 53.285 126.290 53.425 126.455 ;
        RECT 53.225 125.970 53.485 126.290 ;
        RECT 56.045 123.910 56.185 127.330 ;
        RECT 56.505 125.435 58.045 125.805 ;
        RECT 56.905 124.950 57.165 125.270 ;
        RECT 56.965 124.250 57.105 124.950 ;
        RECT 58.805 124.250 58.945 132.575 ;
        RECT 59.265 129.690 59.405 135.150 ;
        RECT 59.205 129.370 59.465 129.690 ;
        RECT 59.665 128.690 59.925 129.010 ;
        RECT 59.725 127.650 59.865 128.690 ;
        RECT 59.665 127.330 59.925 127.650 ;
        RECT 56.905 123.930 57.165 124.250 ;
        RECT 58.745 123.930 59.005 124.250 ;
        RECT 55.985 123.590 56.245 123.910 ;
        RECT 53.205 122.715 54.745 123.085 ;
        RECT 52.765 121.550 53.025 121.870 ;
        RECT 51.445 119.090 52.505 119.230 ;
        RECT 50.925 116.450 51.185 116.770 ;
        RECT 49.545 116.110 49.805 116.430 ;
        RECT 50.465 116.110 50.725 116.430 ;
        RECT 49.605 115.410 49.745 116.110 ;
        RECT 49.545 115.090 49.805 115.410 ;
        RECT 50.915 112.855 51.195 113.225 ;
        RECT 51.445 113.030 51.585 119.090 ;
        RECT 52.305 118.150 52.565 118.470 ;
        RECT 52.365 117.110 52.505 118.150 ;
        RECT 52.305 116.790 52.565 117.110 ;
        RECT 52.825 116.430 52.965 121.550 ;
        RECT 55.525 120.530 55.785 120.850 ;
        RECT 55.585 119.150 55.725 120.530 ;
        RECT 55.525 118.830 55.785 119.150 ;
        RECT 56.045 118.720 56.185 123.590 ;
        RECT 59.665 122.065 59.925 122.210 ;
        RECT 59.655 121.695 59.935 122.065 ;
        RECT 56.505 119.995 58.045 120.365 ;
        RECT 60.185 118.810 60.325 136.850 ;
        RECT 60.585 133.110 60.845 133.430 ;
        RECT 60.645 125.180 60.785 133.110 ;
        RECT 61.105 131.730 61.245 145.350 ;
        RECT 61.505 143.310 61.765 143.630 ;
        RECT 61.565 141.590 61.705 143.310 ;
        RECT 61.505 141.270 61.765 141.590 ;
        RECT 61.965 139.570 62.225 139.890 ;
        RECT 62.025 137.510 62.165 139.570 ;
        RECT 63.335 138.015 63.615 138.385 ;
        RECT 63.865 138.190 64.005 148.895 ;
        RECT 64.325 138.190 64.465 165.330 ;
        RECT 67.085 162.070 67.225 167.790 ;
        RECT 68.005 167.430 68.145 170.510 ;
        RECT 71.625 169.490 71.885 169.810 ;
        RECT 71.685 168.110 71.825 169.490 ;
        RECT 71.625 167.790 71.885 168.110 ;
        RECT 67.945 167.110 68.205 167.430 ;
        RECT 67.485 166.770 67.745 167.090 ;
        RECT 67.545 162.670 67.685 166.770 ;
        RECT 68.005 165.050 68.145 167.110 ;
        RECT 67.945 164.730 68.205 165.050 ;
        RECT 71.625 164.730 71.885 165.050 ;
        RECT 71.685 163.350 71.825 164.730 ;
        RECT 71.625 163.030 71.885 163.350 ;
        RECT 67.485 162.350 67.745 162.670 ;
        RECT 67.085 161.930 67.685 162.070 ;
        RECT 66.105 161.330 66.365 161.650 ;
        RECT 66.165 160.290 66.305 161.330 ;
        RECT 66.105 159.970 66.365 160.290 ;
        RECT 67.545 158.930 67.685 161.930 ;
        RECT 70.705 159.290 70.965 159.610 ;
        RECT 67.485 158.610 67.745 158.930 ;
        RECT 68.865 158.610 69.125 158.930 ;
        RECT 65.645 156.570 65.905 156.890 ;
        RECT 65.185 156.230 65.445 156.550 ;
        RECT 64.725 154.530 64.985 154.850 ;
        RECT 64.785 149.750 64.925 154.530 ;
        RECT 65.245 153.490 65.385 156.230 ;
        RECT 65.705 154.170 65.845 156.570 ;
        RECT 65.645 153.850 65.905 154.170 ;
        RECT 65.185 153.170 65.445 153.490 ;
        RECT 65.245 151.450 65.385 153.170 ;
        RECT 65.185 151.130 65.445 151.450 ;
        RECT 64.725 149.430 64.985 149.750 ;
        RECT 66.565 142.970 66.825 143.290 ;
        RECT 66.625 141.590 66.765 142.970 ;
        RECT 66.565 141.270 66.825 141.590 ;
        RECT 67.025 140.930 67.285 141.250 ;
        RECT 64.725 139.570 64.985 139.890 ;
        RECT 64.785 138.190 64.925 139.570 ;
        RECT 67.085 138.530 67.225 140.930 ;
        RECT 67.025 138.210 67.285 138.530 ;
        RECT 61.965 137.190 62.225 137.510 ;
        RECT 62.025 135.810 62.165 137.190 ;
        RECT 62.885 135.830 63.145 136.150 ;
        RECT 61.965 135.490 62.225 135.810 ;
        RECT 61.505 134.470 61.765 134.790 ;
        RECT 61.045 131.410 61.305 131.730 ;
        RECT 61.105 129.350 61.245 131.410 ;
        RECT 61.045 129.030 61.305 129.350 ;
        RECT 60.645 125.040 61.245 125.180 ;
        RECT 60.575 124.415 60.855 124.785 ;
        RECT 60.585 124.270 60.845 124.415 ;
        RECT 61.105 124.250 61.245 125.040 ;
        RECT 61.045 123.930 61.305 124.250 ;
        RECT 60.585 123.250 60.845 123.570 ;
        RECT 61.045 123.250 61.305 123.570 ;
        RECT 60.645 119.490 60.785 123.250 ;
        RECT 60.585 119.170 60.845 119.490 ;
        RECT 61.105 119.150 61.245 123.250 ;
        RECT 61.045 118.830 61.305 119.150 ;
        RECT 56.905 118.720 57.165 118.810 ;
        RECT 56.045 118.580 57.165 118.720 ;
        RECT 56.905 118.490 57.165 118.580 ;
        RECT 60.125 118.490 60.385 118.810 ;
        RECT 53.205 117.275 54.745 117.645 ;
        RECT 52.765 116.110 53.025 116.430 ;
        RECT 50.925 112.710 51.185 112.855 ;
        RECT 51.385 112.710 51.645 113.030 ;
        RECT 51.445 110.990 51.585 112.710 ;
        RECT 51.385 110.670 51.645 110.990 ;
        RECT 47.245 110.330 47.505 110.650 ;
        RECT 46.785 108.630 47.045 108.950 ;
        RECT 37.585 106.930 37.845 107.250 ;
        RECT 37.645 105.890 37.785 106.930 ;
        RECT 38.105 106.230 38.245 107.530 ;
        RECT 41.265 107.270 41.525 107.590 ;
        RECT 42.645 107.270 42.905 107.590 ;
        RECT 45.405 106.930 45.665 107.250 ;
        RECT 38.045 105.910 38.305 106.230 ;
        RECT 37.585 105.570 37.845 105.890 ;
        RECT 45.465 105.550 45.605 106.930 ;
        RECT 47.305 105.550 47.445 110.330 ;
        RECT 49.085 109.650 49.345 109.970 ;
        RECT 49.145 107.590 49.285 109.650 ;
        RECT 52.825 108.950 52.965 116.110 ;
        RECT 56.965 116.090 57.105 118.490 ;
        RECT 58.285 117.810 58.545 118.130 ;
        RECT 56.905 115.770 57.165 116.090 ;
        RECT 56.505 114.555 58.045 114.925 ;
        RECT 55.525 113.390 55.785 113.710 ;
        RECT 53.205 111.835 54.745 112.205 ;
        RECT 55.585 109.970 55.725 113.390 ;
        RECT 55.985 113.225 56.245 113.370 ;
        RECT 55.975 112.855 56.255 113.225 ;
        RECT 55.985 112.370 56.245 112.690 ;
        RECT 56.445 112.370 56.705 112.690 ;
        RECT 56.045 111.330 56.185 112.370 ;
        RECT 56.505 111.670 56.645 112.370 ;
        RECT 56.445 111.350 56.705 111.670 ;
        RECT 55.985 111.010 56.245 111.330 ;
        RECT 55.525 109.650 55.785 109.970 ;
        RECT 52.765 108.630 53.025 108.950 ;
        RECT 49.085 107.270 49.345 107.590 ;
        RECT 45.405 105.230 45.665 105.550 ;
        RECT 47.245 105.230 47.505 105.550 ;
        RECT 50.465 104.890 50.725 105.210 ;
        RECT 17.635 103.675 19.175 104.045 ;
        RECT 50.525 98.340 50.665 104.890 ;
        RECT 52.825 102.400 52.965 108.630 ;
        RECT 55.585 108.270 55.725 109.650 ;
        RECT 56.505 109.115 58.045 109.485 ;
        RECT 55.525 107.950 55.785 108.270 ;
        RECT 53.205 106.395 54.745 106.765 ;
        RECT 58.345 105.890 58.485 117.810 ;
        RECT 58.745 116.110 59.005 116.430 ;
        RECT 58.805 108.950 58.945 116.110 ;
        RECT 59.665 115.770 59.925 116.090 ;
        RECT 60.125 115.770 60.385 116.090 ;
        RECT 59.725 110.650 59.865 115.770 ;
        RECT 60.185 115.410 60.325 115.770 ;
        RECT 60.125 115.090 60.385 115.410 ;
        RECT 60.585 115.090 60.845 115.410 ;
        RECT 59.665 110.330 59.925 110.650 ;
        RECT 58.745 108.630 59.005 108.950 ;
        RECT 59.725 107.590 59.865 110.330 ;
        RECT 60.645 107.930 60.785 115.090 ;
        RECT 61.045 112.370 61.305 112.690 ;
        RECT 61.105 110.990 61.245 112.370 ;
        RECT 61.045 110.670 61.305 110.990 ;
        RECT 61.565 107.930 61.705 134.470 ;
        RECT 62.425 128.690 62.685 129.010 ;
        RECT 62.485 126.970 62.625 128.690 ;
        RECT 62.425 126.650 62.685 126.970 ;
        RECT 62.485 124.930 62.625 126.650 ;
        RECT 62.425 124.610 62.685 124.930 ;
        RECT 62.425 124.105 62.685 124.250 ;
        RECT 62.415 123.735 62.695 124.105 ;
        RECT 62.025 121.870 62.625 121.950 ;
        RECT 62.945 121.870 63.085 135.830 ;
        RECT 63.405 135.040 63.545 138.015 ;
        RECT 63.805 137.870 64.065 138.190 ;
        RECT 64.265 137.870 64.525 138.190 ;
        RECT 64.725 137.870 64.985 138.190 ;
        RECT 66.105 137.870 66.365 138.190 ;
        RECT 65.185 136.850 65.445 137.170 ;
        RECT 64.255 135.295 64.535 135.665 ;
        RECT 64.265 135.150 64.525 135.295 ;
        RECT 63.805 135.040 64.065 135.130 ;
        RECT 63.405 134.900 64.065 135.040 ;
        RECT 61.965 121.810 62.625 121.870 ;
        RECT 61.965 121.550 62.225 121.810 ;
        RECT 62.485 121.530 62.625 121.810 ;
        RECT 62.885 121.550 63.145 121.870 ;
        RECT 62.425 121.210 62.685 121.530 ;
        RECT 61.965 120.870 62.225 121.190 ;
        RECT 62.025 119.345 62.165 120.870 ;
        RECT 61.955 118.975 62.235 119.345 ;
        RECT 61.965 118.490 62.225 118.810 ;
        RECT 62.885 118.490 63.145 118.810 ;
        RECT 62.025 114.390 62.165 118.490 ;
        RECT 61.965 114.070 62.225 114.390 ;
        RECT 62.945 113.030 63.085 118.490 ;
        RECT 63.405 113.370 63.545 134.900 ;
        RECT 63.805 134.810 64.065 134.900 ;
        RECT 64.325 132.265 64.465 135.150 ;
        RECT 64.725 134.130 64.985 134.450 ;
        RECT 64.785 133.430 64.925 134.130 ;
        RECT 64.725 133.110 64.985 133.430 ;
        RECT 64.255 131.895 64.535 132.265 ;
        RECT 64.265 128.690 64.525 129.010 ;
        RECT 64.325 127.310 64.465 128.690 ;
        RECT 64.265 126.990 64.525 127.310 ;
        RECT 63.805 123.250 64.065 123.570 ;
        RECT 63.865 121.530 64.005 123.250 ;
        RECT 63.805 121.210 64.065 121.530 ;
        RECT 64.265 120.530 64.525 120.850 ;
        RECT 64.325 118.810 64.465 120.530 ;
        RECT 65.245 118.810 65.385 136.850 ;
        RECT 66.165 135.550 66.305 137.870 ;
        RECT 67.545 137.590 67.685 158.610 ;
        RECT 68.925 156.550 69.065 158.610 ;
        RECT 68.865 156.230 69.125 156.550 ;
        RECT 70.765 156.210 70.905 159.290 ;
        RECT 73.005 158.610 73.265 158.930 ;
        RECT 73.065 157.230 73.205 158.610 ;
        RECT 72.545 156.910 72.805 157.230 ;
        RECT 73.005 156.910 73.265 157.230 ;
        RECT 72.605 156.210 72.745 156.910 ;
        RECT 70.705 155.890 70.965 156.210 ;
        RECT 72.545 155.890 72.805 156.210 ;
        RECT 68.405 153.850 68.665 154.170 ;
        RECT 68.465 152.470 68.605 153.850 ;
        RECT 68.405 152.150 68.665 152.470 ;
        RECT 71.165 151.810 71.425 152.130 ;
        RECT 71.225 149.750 71.365 151.810 ;
        RECT 73.525 150.770 73.665 182.470 ;
        RECT 73.985 182.470 74.585 182.610 ;
        RECT 73.985 181.370 74.125 182.470 ;
        RECT 79.045 181.710 79.185 186.830 ;
        RECT 80.825 181.730 81.085 182.050 ;
        RECT 78.985 181.390 79.245 181.710 ;
        RECT 79.905 181.390 80.165 181.710 ;
        RECT 73.925 181.050 74.185 181.370 ;
        RECT 78.065 181.050 78.325 181.370 ;
        RECT 79.445 181.050 79.705 181.370 ;
        RECT 73.985 178.990 74.125 181.050 ;
        RECT 78.125 179.185 78.265 181.050 ;
        RECT 78.525 180.370 78.785 180.690 ;
        RECT 78.985 180.370 79.245 180.690 ;
        RECT 73.925 178.670 74.185 178.990 ;
        RECT 74.375 178.815 74.655 179.185 ;
        RECT 78.055 178.815 78.335 179.185 ;
        RECT 78.585 178.990 78.725 180.370 ;
        RECT 73.985 170.150 74.125 178.670 ;
        RECT 74.445 176.270 74.585 178.815 ;
        RECT 78.525 178.670 78.785 178.990 ;
        RECT 79.045 178.310 79.185 180.370 ;
        RECT 76.685 177.990 76.945 178.310 ;
        RECT 78.985 177.990 79.245 178.310 ;
        RECT 74.845 176.630 75.105 176.950 ;
        RECT 74.385 175.950 74.645 176.270 ;
        RECT 74.905 173.210 75.045 176.630 ;
        RECT 75.755 176.095 76.035 176.465 ;
        RECT 76.745 176.270 76.885 177.990 ;
        RECT 79.505 177.970 79.645 181.050 ;
        RECT 79.445 177.650 79.705 177.970 ;
        RECT 79.505 176.270 79.645 177.650 ;
        RECT 75.765 175.950 76.025 176.095 ;
        RECT 76.685 175.950 76.945 176.270 ;
        RECT 79.445 175.950 79.705 176.270 ;
        RECT 76.675 175.415 76.955 175.785 ;
        RECT 76.685 175.270 76.945 175.415 ;
        RECT 74.845 172.890 75.105 173.210 ;
        RECT 75.765 172.890 76.025 173.210 ;
        RECT 74.385 170.510 74.645 170.830 ;
        RECT 73.925 169.830 74.185 170.150 ;
        RECT 73.985 168.110 74.125 169.830 ;
        RECT 73.925 167.790 74.185 168.110 ;
        RECT 73.985 165.390 74.125 167.790 ;
        RECT 74.445 167.430 74.585 170.510 ;
        RECT 74.845 169.490 75.105 169.810 ;
        RECT 74.905 168.870 75.045 169.490 ;
        RECT 74.905 168.790 75.505 168.870 ;
        RECT 74.905 168.730 75.565 168.790 ;
        RECT 74.385 167.110 74.645 167.430 ;
        RECT 74.905 165.390 75.045 168.730 ;
        RECT 75.305 168.470 75.565 168.730 ;
        RECT 73.925 165.070 74.185 165.390 ;
        RECT 74.845 165.070 75.105 165.390 ;
        RECT 73.985 163.350 74.125 165.070 ;
        RECT 73.925 163.030 74.185 163.350 ;
        RECT 73.985 159.610 74.125 163.030 ;
        RECT 74.905 159.950 75.045 165.070 ;
        RECT 74.845 159.630 75.105 159.950 ;
        RECT 73.925 159.290 74.185 159.610 ;
        RECT 73.985 157.310 74.125 159.290 ;
        RECT 73.985 157.230 74.585 157.310 ;
        RECT 73.985 157.170 74.645 157.230 ;
        RECT 73.985 154.510 74.125 157.170 ;
        RECT 74.385 156.910 74.645 157.170 ;
        RECT 74.905 156.800 75.045 159.630 ;
        RECT 75.305 156.800 75.565 156.890 ;
        RECT 74.905 156.660 75.565 156.800 ;
        RECT 75.305 156.570 75.565 156.660 ;
        RECT 73.925 154.190 74.185 154.510 ;
        RECT 73.985 151.790 74.125 154.190 ;
        RECT 73.925 151.470 74.185 151.790 ;
        RECT 74.845 150.790 75.105 151.110 ;
        RECT 73.465 150.450 73.725 150.770 ;
        RECT 74.905 149.750 75.045 150.790 ;
        RECT 71.165 149.430 71.425 149.750 ;
        RECT 74.845 149.430 75.105 149.750 ;
        RECT 75.365 149.070 75.505 156.570 ;
        RECT 75.825 156.550 75.965 172.890 ;
        RECT 77.605 172.550 77.865 172.870 ;
        RECT 77.665 171.510 77.805 172.550 ;
        RECT 77.605 171.190 77.865 171.510 ;
        RECT 77.665 168.790 77.805 171.190 ;
        RECT 78.985 170.510 79.245 170.830 ;
        RECT 79.045 169.810 79.185 170.510 ;
        RECT 78.985 169.490 79.245 169.810 ;
        RECT 77.605 168.470 77.865 168.790 ;
        RECT 77.145 159.970 77.405 160.290 ;
        RECT 77.205 157.910 77.345 159.970 ;
        RECT 77.145 157.590 77.405 157.910 ;
        RECT 75.765 156.230 76.025 156.550 ;
        RECT 79.505 156.210 79.645 175.950 ;
        RECT 79.965 173.210 80.105 181.390 ;
        RECT 80.885 179.670 81.025 181.730 ;
        RECT 81.805 181.710 81.945 187.510 ;
        RECT 81.745 181.390 82.005 181.710 ;
        RECT 80.825 179.350 81.085 179.670 ;
        RECT 80.365 177.650 80.625 177.970 ;
        RECT 80.425 176.950 80.565 177.650 ;
        RECT 80.365 176.630 80.625 176.950 ;
        RECT 80.885 176.180 81.025 179.350 ;
        RECT 82.265 179.330 82.405 189.550 ;
        RECT 83.645 186.810 83.785 189.550 ;
        RECT 85.885 188.870 86.145 189.190 ;
        RECT 84.045 188.530 84.305 188.850 ;
        RECT 84.105 187.490 84.245 188.530 ;
        RECT 84.045 187.170 84.305 187.490 ;
        RECT 83.585 186.490 83.845 186.810 ;
        RECT 85.425 185.810 85.685 186.130 ;
        RECT 85.485 184.770 85.625 185.810 ;
        RECT 85.945 185.110 86.085 188.870 ;
        RECT 86.865 187.830 87.005 191.930 ;
        RECT 87.785 189.530 87.925 192.270 ;
        RECT 87.725 189.210 87.985 189.530 ;
        RECT 86.805 187.510 87.065 187.830 ;
        RECT 86.345 187.170 86.605 187.490 ;
        RECT 85.885 184.790 86.145 185.110 ;
        RECT 85.425 184.450 85.685 184.770 ;
        RECT 82.665 183.090 82.925 183.410 ;
        RECT 82.725 181.710 82.865 183.090 ;
        RECT 84.965 181.730 85.225 182.050 ;
        RECT 82.665 181.390 82.925 181.710 ;
        RECT 82.205 179.010 82.465 179.330 ;
        RECT 81.285 178.670 81.545 178.990 ;
        RECT 81.345 176.950 81.485 178.670 ;
        RECT 81.735 177.030 82.015 177.145 ;
        RECT 82.725 177.030 82.865 181.390 ;
        RECT 83.585 180.370 83.845 180.690 ;
        RECT 84.505 180.370 84.765 180.690 ;
        RECT 83.645 179.670 83.785 180.370 ;
        RECT 83.585 179.350 83.845 179.670 ;
        RECT 84.565 178.990 84.705 180.370 ;
        RECT 84.505 178.670 84.765 178.990 ;
        RECT 84.045 178.330 84.305 178.650 ;
        RECT 85.025 178.390 85.165 181.730 ;
        RECT 81.285 176.630 81.545 176.950 ;
        RECT 81.735 176.890 82.865 177.030 ;
        RECT 84.105 176.950 84.245 178.330 ;
        RECT 84.565 178.250 85.165 178.390 ;
        RECT 84.565 177.970 84.705 178.250 ;
        RECT 84.505 177.650 84.765 177.970 ;
        RECT 81.735 176.775 82.015 176.890 ;
        RECT 81.285 176.180 81.545 176.270 ;
        RECT 80.885 176.040 81.545 176.180 ;
        RECT 81.285 175.950 81.545 176.040 ;
        RECT 79.905 172.890 80.165 173.210 ;
        RECT 79.965 170.830 80.105 172.890 ;
        RECT 79.905 170.510 80.165 170.830 ;
        RECT 79.445 155.890 79.705 156.210 ;
        RECT 79.445 154.530 79.705 154.850 ;
        RECT 76.685 151.470 76.945 151.790 ;
        RECT 76.745 149.410 76.885 151.470 ;
        RECT 79.505 149.750 79.645 154.530 ;
        RECT 79.445 149.430 79.705 149.750 ;
        RECT 76.685 149.090 76.945 149.410 ;
        RECT 79.965 149.070 80.105 170.510 ;
        RECT 81.345 170.400 81.485 175.950 ;
        RECT 81.805 172.950 81.945 176.775 ;
        RECT 84.045 176.630 84.305 176.950 ;
        RECT 84.565 176.270 84.705 177.650 ;
        RECT 82.665 175.950 82.925 176.270 ;
        RECT 83.125 175.950 83.385 176.270 ;
        RECT 83.585 175.950 83.845 176.270 ;
        RECT 84.045 175.950 84.305 176.270 ;
        RECT 84.505 175.950 84.765 176.270 ;
        RECT 82.205 175.270 82.465 175.590 ;
        RECT 82.265 173.550 82.405 175.270 ;
        RECT 82.205 173.230 82.465 173.550 ;
        RECT 81.805 172.810 82.405 172.950 ;
        RECT 82.725 172.870 82.865 175.950 ;
        RECT 83.185 175.250 83.325 175.950 ;
        RECT 83.645 175.590 83.785 175.950 ;
        RECT 83.585 175.270 83.845 175.590 ;
        RECT 83.125 174.930 83.385 175.250 ;
        RECT 83.645 173.550 83.785 175.270 ;
        RECT 83.125 173.230 83.385 173.550 ;
        RECT 83.585 173.230 83.845 173.550 ;
        RECT 84.105 173.460 84.245 175.950 ;
        RECT 84.105 173.320 84.705 173.460 ;
        RECT 81.745 172.210 82.005 172.530 ;
        RECT 81.805 171.170 81.945 172.210 ;
        RECT 81.745 170.850 82.005 171.170 ;
        RECT 81.345 170.260 81.945 170.400 ;
        RECT 81.285 169.490 81.545 169.810 ;
        RECT 80.365 161.330 80.625 161.650 ;
        RECT 80.425 159.860 80.565 161.330 ;
        RECT 80.825 159.860 81.085 159.950 ;
        RECT 80.425 159.720 81.085 159.860 ;
        RECT 80.825 159.630 81.085 159.720 ;
        RECT 81.345 157.570 81.485 169.490 ;
        RECT 81.805 167.000 81.945 170.260 ;
        RECT 82.265 167.770 82.405 172.810 ;
        RECT 82.665 172.550 82.925 172.870 ;
        RECT 83.185 170.230 83.325 173.230 ;
        RECT 83.645 172.950 83.785 173.230 ;
        RECT 84.565 173.120 84.705 173.320 ;
        RECT 84.965 173.120 85.225 173.210 ;
        RECT 84.565 172.980 85.225 173.120 ;
        RECT 83.645 172.810 84.245 172.950 ;
        RECT 84.965 172.890 85.225 172.980 ;
        RECT 83.585 172.210 83.845 172.530 ;
        RECT 83.645 171.510 83.785 172.210 ;
        RECT 83.585 171.190 83.845 171.510 ;
        RECT 82.725 170.150 83.325 170.230 ;
        RECT 82.665 170.090 83.325 170.150 ;
        RECT 82.665 169.830 82.925 170.090 ;
        RECT 82.725 168.110 82.865 169.830 ;
        RECT 82.665 167.790 82.925 168.110 ;
        RECT 82.205 167.450 82.465 167.770 ;
        RECT 81.805 166.860 82.405 167.000 ;
        RECT 81.745 161.670 82.005 161.990 ;
        RECT 81.805 159.950 81.945 161.670 ;
        RECT 81.745 159.630 82.005 159.950 ;
        RECT 82.265 157.910 82.405 166.860 ;
        RECT 82.725 162.670 82.865 167.790 ;
        RECT 83.645 167.770 83.785 171.190 ;
        RECT 83.585 167.450 83.845 167.770 ;
        RECT 82.665 162.350 82.925 162.670 ;
        RECT 83.585 161.670 83.845 161.990 ;
        RECT 83.645 160.630 83.785 161.670 ;
        RECT 84.105 160.630 84.245 172.810 ;
        RECT 84.965 167.340 85.225 167.430 ;
        RECT 85.485 167.340 85.625 184.450 ;
        RECT 85.945 184.430 86.085 184.790 ;
        RECT 85.885 184.110 86.145 184.430 ;
        RECT 85.945 169.810 86.085 184.110 ;
        RECT 85.885 169.490 86.145 169.810 ;
        RECT 86.405 168.790 86.545 187.170 ;
        RECT 88.245 184.510 88.385 192.610 ;
        RECT 105.265 192.590 105.405 194.340 ;
        RECT 90.485 192.270 90.745 192.590 ;
        RECT 97.845 192.270 98.105 192.590 ;
        RECT 105.205 192.270 105.465 192.590 ;
        RECT 90.025 191.930 90.285 192.250 ;
        RECT 87.325 184.370 88.385 184.510 ;
        RECT 90.085 184.430 90.225 191.930 ;
        RECT 90.545 188.850 90.685 192.270 ;
        RECT 93.245 191.250 93.505 191.570 ;
        RECT 94.165 191.250 94.425 191.570 ;
        RECT 93.305 189.870 93.445 191.250 ;
        RECT 93.245 189.550 93.505 189.870 ;
        RECT 94.225 189.190 94.365 191.250 ;
        RECT 95.375 190.715 96.915 191.085 ;
        RECT 94.165 188.870 94.425 189.190 ;
        RECT 90.485 188.530 90.745 188.850 ;
        RECT 86.805 183.770 87.065 184.090 ;
        RECT 86.865 183.265 87.005 183.770 ;
        RECT 86.795 182.895 87.075 183.265 ;
        RECT 87.325 183.150 87.465 184.370 ;
        RECT 90.025 184.110 90.285 184.430 ;
        RECT 90.545 183.830 90.685 188.530 ;
        RECT 92.075 187.995 93.615 188.365 ;
        RECT 91.405 187.170 91.665 187.490 ;
        RECT 87.785 183.750 90.685 183.830 ;
        RECT 87.725 183.690 90.745 183.750 ;
        RECT 87.725 183.430 87.985 183.690 ;
        RECT 90.485 183.430 90.745 183.690 ;
        RECT 87.325 183.010 87.925 183.150 ;
        RECT 89.565 183.090 89.825 183.410 ;
        RECT 90.025 183.265 90.285 183.410 ;
        RECT 87.785 182.390 87.925 183.010 ;
        RECT 87.265 182.070 87.525 182.390 ;
        RECT 87.725 182.070 87.985 182.390 ;
        RECT 86.805 181.390 87.065 181.710 ;
        RECT 86.865 177.970 87.005 181.390 ;
        RECT 87.325 178.990 87.465 182.070 ;
        RECT 89.105 181.390 89.365 181.710 ;
        RECT 88.185 181.050 88.445 181.370 ;
        RECT 88.245 179.330 88.385 181.050 ;
        RECT 88.185 179.010 88.445 179.330 ;
        RECT 87.265 178.670 87.525 178.990 ;
        RECT 86.805 177.650 87.065 177.970 ;
        RECT 86.865 176.610 87.005 177.650 ;
        RECT 87.325 176.950 87.465 178.670 ;
        RECT 87.265 176.630 87.525 176.950 ;
        RECT 86.805 176.290 87.065 176.610 ;
        RECT 86.805 174.930 87.065 175.250 ;
        RECT 86.865 172.950 87.005 174.930 ;
        RECT 89.165 174.230 89.305 181.390 ;
        RECT 89.625 180.690 89.765 183.090 ;
        RECT 90.015 182.895 90.295 183.265 ;
        RECT 91.465 182.390 91.605 187.170 ;
        RECT 93.705 186.490 93.965 186.810 ;
        RECT 93.765 185.110 93.905 186.490 ;
        RECT 95.375 185.275 96.915 185.645 ;
        RECT 93.705 184.790 93.965 185.110 ;
        RECT 97.905 183.750 98.045 192.270 ;
        RECT 103.825 191.250 104.085 191.570 ;
        RECT 98.765 189.550 99.025 189.870 ;
        RECT 98.825 186.810 98.965 189.550 ;
        RECT 98.765 186.490 99.025 186.810 ;
        RECT 97.845 183.430 98.105 183.750 ;
        RECT 92.075 182.555 93.615 182.925 ;
        RECT 91.405 182.070 91.665 182.390 ;
        RECT 97.905 182.050 98.045 183.430 ;
        RECT 97.845 181.730 98.105 182.050 ;
        RECT 93.705 181.390 93.965 181.710 ;
        RECT 94.625 181.390 94.885 181.710 ;
        RECT 90.485 181.050 90.745 181.370 ;
        RECT 89.565 180.370 89.825 180.690 ;
        RECT 90.025 180.370 90.285 180.690 ;
        RECT 90.085 178.650 90.225 180.370 ;
        RECT 90.545 178.650 90.685 181.050 ;
        RECT 91.865 180.710 92.125 181.030 ;
        RECT 91.395 178.815 91.675 179.185 ;
        RECT 90.025 178.330 90.285 178.650 ;
        RECT 90.485 178.330 90.745 178.650 ;
        RECT 89.565 175.610 89.825 175.930 ;
        RECT 90.085 175.785 90.225 178.330 ;
        RECT 89.105 173.910 89.365 174.230 ;
        RECT 86.865 172.810 87.465 172.950 ;
        RECT 87.325 172.530 87.465 172.810 ;
        RECT 86.805 172.210 87.065 172.530 ;
        RECT 87.265 172.210 87.525 172.530 ;
        RECT 86.865 170.830 87.005 172.210 ;
        RECT 86.805 170.510 87.065 170.830 ;
        RECT 86.345 168.470 86.605 168.790 ;
        RECT 86.345 167.790 86.605 168.110 ;
        RECT 84.965 167.200 85.625 167.340 ;
        RECT 84.965 167.110 85.225 167.200 ;
        RECT 84.505 166.770 84.765 167.090 ;
        RECT 84.565 164.370 84.705 166.770 ;
        RECT 84.505 164.050 84.765 164.370 ;
        RECT 84.565 161.650 84.705 164.050 ;
        RECT 84.505 161.330 84.765 161.650 ;
        RECT 83.585 160.310 83.845 160.630 ;
        RECT 84.045 160.310 84.305 160.630 ;
        RECT 82.205 157.590 82.465 157.910 ;
        RECT 81.285 157.250 81.545 157.570 ;
        RECT 83.125 156.910 83.385 157.230 ;
        RECT 82.205 154.190 82.465 154.510 ;
        RECT 80.365 153.170 80.625 153.490 ;
        RECT 80.425 151.790 80.565 153.170 ;
        RECT 82.265 152.470 82.405 154.190 ;
        RECT 82.205 152.150 82.465 152.470 ;
        RECT 80.365 151.470 80.625 151.790 ;
        RECT 83.185 149.410 83.325 156.910 ;
        RECT 83.645 156.890 83.785 160.310 ;
        RECT 83.585 156.570 83.845 156.890 ;
        RECT 84.105 156.800 84.245 160.310 ;
        RECT 84.565 159.950 84.705 161.330 ;
        RECT 84.505 159.630 84.765 159.950 ;
        RECT 84.505 156.800 84.765 156.890 ;
        RECT 84.105 156.660 84.765 156.800 ;
        RECT 84.505 156.570 84.765 156.660 ;
        RECT 85.025 154.850 85.165 167.110 ;
        RECT 85.885 166.770 86.145 167.090 ;
        RECT 85.945 165.390 86.085 166.770 ;
        RECT 85.885 165.070 86.145 165.390 ;
        RECT 85.425 164.730 85.685 165.050 ;
        RECT 85.485 162.330 85.625 164.730 ;
        RECT 85.425 162.010 85.685 162.330 ;
        RECT 85.425 160.310 85.685 160.630 ;
        RECT 85.485 159.950 85.625 160.310 ;
        RECT 85.425 159.630 85.685 159.950 ;
        RECT 85.425 158.950 85.685 159.270 ;
        RECT 85.485 157.230 85.625 158.950 ;
        RECT 86.405 157.310 86.545 167.790 ;
        RECT 86.805 167.450 87.065 167.770 ;
        RECT 86.865 160.630 87.005 167.450 ;
        RECT 86.805 160.310 87.065 160.630 ;
        RECT 87.325 159.610 87.465 172.210 ;
        RECT 89.625 170.830 89.765 175.610 ;
        RECT 90.015 175.415 90.295 175.785 ;
        RECT 89.565 170.510 89.825 170.830 ;
        RECT 88.645 167.790 88.905 168.110 ;
        RECT 88.705 160.630 88.845 167.790 ;
        RECT 90.085 167.770 90.225 175.415 ;
        RECT 90.545 168.110 90.685 178.330 ;
        RECT 90.945 177.650 91.205 177.970 ;
        RECT 91.005 168.450 91.145 177.650 ;
        RECT 91.465 168.790 91.605 178.815 ;
        RECT 91.925 178.650 92.065 180.710 ;
        RECT 93.765 180.690 93.905 181.390 ;
        RECT 93.705 180.370 93.965 180.690 ;
        RECT 92.775 178.815 93.055 179.185 ;
        RECT 94.685 178.900 94.825 181.390 ;
        RECT 95.375 179.835 96.915 180.205 ;
        RECT 92.785 178.670 93.045 178.815 ;
        RECT 94.225 178.760 94.825 178.900 ;
        RECT 91.865 178.330 92.125 178.650 ;
        RECT 91.925 177.970 92.065 178.330 ;
        RECT 91.865 177.650 92.125 177.970 ;
        RECT 93.705 177.650 93.965 177.970 ;
        RECT 92.075 177.115 93.615 177.485 ;
        RECT 92.075 171.675 93.615 172.045 ;
        RECT 93.245 169.720 93.505 169.810 ;
        RECT 93.765 169.720 93.905 177.650 ;
        RECT 94.225 173.550 94.365 178.760 ;
        RECT 97.905 178.650 98.045 181.730 ;
        RECT 97.845 178.330 98.105 178.650 ;
        RECT 94.625 177.990 94.885 178.310 ;
        RECT 94.685 175.250 94.825 177.990 ;
        RECT 96.005 177.650 96.265 177.970 ;
        RECT 96.925 177.650 97.185 177.970 ;
        RECT 96.065 176.950 96.205 177.650 ;
        RECT 96.005 176.630 96.265 176.950 ;
        RECT 96.985 176.610 97.125 177.650 ;
        RECT 96.925 176.290 97.185 176.610 ;
        RECT 98.825 175.930 98.965 186.490 ;
        RECT 103.885 184.090 104.025 191.250 ;
        RECT 103.825 183.770 104.085 184.090 ;
        RECT 100.145 183.090 100.405 183.410 ;
        RECT 98.765 175.610 99.025 175.930 ;
        RECT 94.625 174.930 94.885 175.250 ;
        RECT 94.165 173.230 94.425 173.550 ;
        RECT 94.685 173.210 94.825 174.930 ;
        RECT 95.375 174.395 96.915 174.765 ;
        RECT 97.845 173.910 98.105 174.230 ;
        RECT 97.905 173.550 98.045 173.910 ;
        RECT 97.385 173.230 97.645 173.550 ;
        RECT 97.845 173.230 98.105 173.550 ;
        RECT 94.625 172.890 94.885 173.210 ;
        RECT 97.445 172.530 97.585 173.230 ;
        RECT 97.385 172.210 97.645 172.530 ;
        RECT 94.165 170.170 94.425 170.490 ;
        RECT 93.245 169.580 93.905 169.720 ;
        RECT 93.245 169.490 93.505 169.580 ;
        RECT 91.405 168.470 91.665 168.790 ;
        RECT 90.945 168.130 91.205 168.450 ;
        RECT 90.485 167.790 90.745 168.110 ;
        RECT 90.025 167.625 90.285 167.770 ;
        RECT 90.015 167.255 90.295 167.625 ;
        RECT 90.025 166.770 90.285 167.090 ;
        RECT 90.085 166.070 90.225 166.770 ;
        RECT 90.025 165.750 90.285 166.070 ;
        RECT 88.645 160.310 88.905 160.630 ;
        RECT 90.085 159.950 90.225 165.750 ;
        RECT 90.545 160.630 90.685 167.790 ;
        RECT 90.485 160.310 90.745 160.630 ;
        RECT 89.105 159.630 89.365 159.950 ;
        RECT 89.565 159.630 89.825 159.950 ;
        RECT 90.025 159.630 90.285 159.950 ;
        RECT 87.265 159.290 87.525 159.610 ;
        RECT 88.185 158.950 88.445 159.270 ;
        RECT 85.425 156.910 85.685 157.230 ;
        RECT 86.405 157.170 87.925 157.310 ;
        RECT 85.485 155.190 85.625 156.910 ;
        RECT 87.785 156.890 87.925 157.170 ;
        RECT 87.265 156.570 87.525 156.890 ;
        RECT 87.725 156.570 87.985 156.890 ;
        RECT 86.805 155.890 87.065 156.210 ;
        RECT 85.425 154.870 85.685 155.190 ;
        RECT 84.965 154.530 85.225 154.850 ;
        RECT 84.965 153.850 85.225 154.170 ;
        RECT 85.025 150.770 85.165 153.850 ;
        RECT 86.865 151.790 87.005 155.890 ;
        RECT 87.325 154.510 87.465 156.570 ;
        RECT 87.265 154.190 87.525 154.510 ;
        RECT 86.805 151.470 87.065 151.790 ;
        RECT 85.425 150.790 85.685 151.110 ;
        RECT 84.965 150.450 85.225 150.770 ;
        RECT 83.125 149.090 83.385 149.410 ;
        RECT 75.305 148.750 75.565 149.070 ;
        RECT 79.905 148.750 80.165 149.070 ;
        RECT 85.485 148.110 85.625 150.790 ;
        RECT 87.325 148.730 87.465 154.190 ;
        RECT 87.725 153.850 87.985 154.170 ;
        RECT 87.785 151.450 87.925 153.850 ;
        RECT 88.245 151.450 88.385 158.950 ;
        RECT 89.165 157.910 89.305 159.630 ;
        RECT 89.105 157.590 89.365 157.910 ;
        RECT 89.165 156.890 89.305 157.590 ;
        RECT 89.105 156.570 89.365 156.890 ;
        RECT 89.625 156.550 89.765 159.630 ;
        RECT 89.565 156.230 89.825 156.550 ;
        RECT 88.645 155.890 88.905 156.210 ;
        RECT 89.105 155.890 89.365 156.210 ;
        RECT 88.705 152.470 88.845 155.890 ;
        RECT 88.645 152.150 88.905 152.470 ;
        RECT 89.165 151.790 89.305 155.890 ;
        RECT 89.565 153.170 89.825 153.490 ;
        RECT 89.105 151.470 89.365 151.790 ;
        RECT 87.725 151.130 87.985 151.450 ;
        RECT 88.185 151.130 88.445 151.450 ;
        RECT 89.625 149.070 89.765 153.170 ;
        RECT 89.565 148.750 89.825 149.070 ;
        RECT 87.265 148.410 87.525 148.730 ;
        RECT 85.485 147.970 86.545 148.110 ;
        RECT 82.665 145.690 82.925 146.010 ;
        RECT 69.785 145.350 70.045 145.670 ;
        RECT 66.565 137.190 66.825 137.510 ;
        RECT 67.085 137.450 67.685 137.590 ;
        RECT 66.625 136.150 66.765 137.190 ;
        RECT 66.565 135.830 66.825 136.150 ;
        RECT 66.165 135.410 66.765 135.550 ;
        RECT 67.085 135.470 67.225 137.450 ;
        RECT 65.645 128.690 65.905 129.010 ;
        RECT 65.705 123.570 65.845 128.690 ;
        RECT 66.625 125.270 66.765 135.410 ;
        RECT 67.025 135.150 67.285 135.470 ;
        RECT 66.565 124.950 66.825 125.270 ;
        RECT 67.085 124.590 67.225 135.150 ;
        RECT 67.485 134.130 67.745 134.450 ;
        RECT 67.545 132.750 67.685 134.130 ;
        RECT 67.485 132.430 67.745 132.750 ;
        RECT 67.945 129.030 68.205 129.350 ;
        RECT 68.005 127.310 68.145 129.030 ;
        RECT 69.325 128.690 69.585 129.010 ;
        RECT 67.945 126.990 68.205 127.310 ;
        RECT 67.025 124.270 67.285 124.590 ;
        RECT 65.645 123.250 65.905 123.570 ;
        RECT 68.405 123.250 68.665 123.570 ;
        RECT 68.465 122.550 68.605 123.250 ;
        RECT 69.385 122.550 69.525 128.690 ;
        RECT 68.405 122.230 68.665 122.550 ;
        RECT 69.325 122.230 69.585 122.550 ;
        RECT 66.565 121.550 66.825 121.870 ;
        RECT 65.645 119.510 65.905 119.830 ;
        RECT 64.265 118.490 64.525 118.810 ;
        RECT 64.725 118.490 64.985 118.810 ;
        RECT 65.185 118.490 65.445 118.810 ;
        RECT 64.785 116.770 64.925 118.490 ;
        RECT 63.805 116.450 64.065 116.770 ;
        RECT 64.725 116.450 64.985 116.770 ;
        RECT 63.345 113.050 63.605 113.370 ;
        RECT 62.885 112.710 63.145 113.030 ;
        RECT 63.865 111.670 64.005 116.450 ;
        RECT 65.705 113.370 65.845 119.510 ;
        RECT 66.625 119.345 66.765 121.550 ;
        RECT 69.325 121.210 69.585 121.530 ;
        RECT 67.485 120.530 67.745 120.850 ;
        RECT 66.555 118.975 66.835 119.345 ;
        RECT 67.545 119.150 67.685 120.530 ;
        RECT 69.385 119.150 69.525 121.210 ;
        RECT 67.485 118.830 67.745 119.150 ;
        RECT 69.325 118.830 69.585 119.150 ;
        RECT 68.865 117.810 69.125 118.130 ;
        RECT 66.565 115.090 66.825 115.410 ;
        RECT 65.645 113.050 65.905 113.370 ;
        RECT 66.625 113.030 66.765 115.090 ;
        RECT 64.265 112.710 64.525 113.030 ;
        RECT 66.565 112.710 66.825 113.030 ;
        RECT 64.325 111.670 64.465 112.710 ;
        RECT 63.805 111.350 64.065 111.670 ;
        RECT 64.265 111.350 64.525 111.670 ;
        RECT 63.345 110.670 63.605 110.990 ;
        RECT 63.405 108.610 63.545 110.670 ;
        RECT 64.325 108.950 64.465 111.350 ;
        RECT 66.625 111.330 66.765 112.710 ;
        RECT 68.405 112.370 68.665 112.690 ;
        RECT 66.565 111.010 66.825 111.330 ;
        RECT 68.465 110.990 68.605 112.370 ;
        RECT 68.405 110.670 68.665 110.990 ;
        RECT 68.405 109.650 68.665 109.970 ;
        RECT 64.265 108.630 64.525 108.950 ;
        RECT 63.345 108.290 63.605 108.610 ;
        RECT 60.585 107.610 60.845 107.930 ;
        RECT 61.505 107.610 61.765 107.930 ;
        RECT 68.465 107.590 68.605 109.650 ;
        RECT 59.665 107.270 59.925 107.590 ;
        RECT 68.405 107.270 68.665 107.590 ;
        RECT 54.605 105.570 54.865 105.890 ;
        RECT 58.285 105.570 58.545 105.890 ;
        RECT 54.665 103.510 54.805 105.570 ;
        RECT 59.725 105.550 59.865 107.270 ;
        RECT 68.925 105.890 69.065 117.810 ;
        RECT 69.845 107.785 69.985 145.350 ;
        RECT 81.745 145.010 82.005 145.330 ;
        RECT 70.245 143.650 70.505 143.970 ;
        RECT 80.365 143.650 80.625 143.970 ;
        RECT 70.305 140.910 70.445 143.650 ;
        RECT 76.225 143.310 76.485 143.630 ;
        RECT 71.625 142.970 71.885 143.290 ;
        RECT 75.305 143.200 75.565 143.290 ;
        RECT 75.305 143.060 75.965 143.200 ;
        RECT 75.305 142.970 75.565 143.060 ;
        RECT 71.685 140.910 71.825 142.970 ;
        RECT 73.005 142.290 73.265 142.610 ;
        RECT 73.065 140.910 73.205 142.290 ;
        RECT 70.245 140.590 70.505 140.910 ;
        RECT 71.625 140.590 71.885 140.910 ;
        RECT 73.005 140.590 73.265 140.910 ;
        RECT 70.305 138.190 70.445 140.590 ;
        RECT 70.245 137.870 70.505 138.190 ;
        RECT 71.685 137.850 71.825 140.590 ;
        RECT 75.825 140.570 75.965 143.060 ;
        RECT 75.765 140.250 76.025 140.570 ;
        RECT 72.545 139.910 72.805 140.230 ;
        RECT 72.605 138.870 72.745 139.910 ;
        RECT 72.545 138.550 72.805 138.870 ;
        RECT 72.085 137.870 72.345 138.190 ;
        RECT 71.625 137.530 71.885 137.850 ;
        RECT 72.145 132.750 72.285 137.870 ;
        RECT 74.385 137.530 74.645 137.850 ;
        RECT 73.005 137.190 73.265 137.510 ;
        RECT 73.065 135.130 73.205 137.190 ;
        RECT 74.445 136.150 74.585 137.530 ;
        RECT 74.385 135.830 74.645 136.150 ;
        RECT 73.005 134.810 73.265 135.130 ;
        RECT 75.305 134.810 75.565 135.130 ;
        RECT 73.925 134.470 74.185 134.790 ;
        RECT 73.005 133.110 73.265 133.430 ;
        RECT 72.085 132.430 72.345 132.750 ;
        RECT 70.705 129.710 70.965 130.030 ;
        RECT 71.625 129.710 71.885 130.030 ;
        RECT 70.765 121.530 70.905 129.710 ;
        RECT 71.165 126.990 71.425 127.310 ;
        RECT 71.225 123.570 71.365 126.990 ;
        RECT 71.685 125.270 71.825 129.710 ;
        RECT 71.625 124.950 71.885 125.270 ;
        RECT 71.165 123.250 71.425 123.570 ;
        RECT 70.705 121.210 70.965 121.530 ;
        RECT 70.245 119.510 70.505 119.830 ;
        RECT 70.305 117.110 70.445 119.510 ;
        RECT 71.165 118.150 71.425 118.470 ;
        RECT 71.225 117.110 71.365 118.150 ;
        RECT 70.245 116.790 70.505 117.110 ;
        RECT 71.165 116.790 71.425 117.110 ;
        RECT 70.245 116.110 70.505 116.430 ;
        RECT 71.625 116.340 71.885 116.430 ;
        RECT 72.145 116.340 72.285 132.430 ;
        RECT 72.545 131.750 72.805 132.070 ;
        RECT 72.605 127.310 72.745 131.750 ;
        RECT 73.065 131.730 73.205 133.110 ;
        RECT 73.985 132.410 74.125 134.470 ;
        RECT 73.925 132.090 74.185 132.410 ;
        RECT 73.005 131.410 73.265 131.730 ;
        RECT 73.925 127.330 74.185 127.650 ;
        RECT 72.545 126.990 72.805 127.310 ;
        RECT 72.605 124.250 72.745 126.990 ;
        RECT 73.005 125.970 73.265 126.290 ;
        RECT 73.065 124.590 73.205 125.970 ;
        RECT 73.005 124.270 73.265 124.590 ;
        RECT 72.545 123.990 72.805 124.250 ;
        RECT 72.545 123.930 73.205 123.990 ;
        RECT 72.605 123.850 73.205 123.930 ;
        RECT 73.065 121.870 73.205 123.850 ;
        RECT 73.985 121.870 74.125 127.330 ;
        RECT 75.365 121.870 75.505 134.810 ;
        RECT 75.825 129.690 75.965 140.250 ;
        RECT 76.285 138.870 76.425 143.310 ;
        RECT 76.685 142.970 76.945 143.290 ;
        RECT 76.225 138.550 76.485 138.870 ;
        RECT 76.225 135.380 76.485 135.470 ;
        RECT 76.745 135.380 76.885 142.970 ;
        RECT 78.065 142.290 78.325 142.610 ;
        RECT 78.125 141.105 78.265 142.290 ;
        RECT 80.425 141.250 80.565 143.650 ;
        RECT 78.055 140.735 78.335 141.105 ;
        RECT 80.365 140.930 80.625 141.250 ;
        RECT 76.225 135.240 76.885 135.380 ;
        RECT 76.225 135.150 76.485 135.240 ;
        RECT 75.765 129.370 76.025 129.690 ;
        RECT 75.825 127.310 75.965 129.370 ;
        RECT 75.765 126.990 76.025 127.310 ;
        RECT 75.765 123.590 76.025 123.910 ;
        RECT 73.005 121.550 73.265 121.870 ;
        RECT 73.925 121.550 74.185 121.870 ;
        RECT 75.305 121.550 75.565 121.870 ;
        RECT 72.545 121.210 72.805 121.530 ;
        RECT 72.605 119.490 72.745 121.210 ;
        RECT 72.545 119.170 72.805 119.490 ;
        RECT 73.985 119.345 74.125 121.550 ;
        RECT 74.845 121.210 75.105 121.530 ;
        RECT 73.915 118.975 74.195 119.345 ;
        RECT 72.545 117.810 72.805 118.130 ;
        RECT 71.625 116.200 72.285 116.340 ;
        RECT 71.625 116.110 71.885 116.200 ;
        RECT 70.305 114.390 70.445 116.110 ;
        RECT 70.245 114.070 70.505 114.390 ;
        RECT 71.685 113.370 71.825 116.110 ;
        RECT 72.605 116.090 72.745 117.810 ;
        RECT 73.985 116.430 74.125 118.975 ;
        RECT 73.925 116.110 74.185 116.430 ;
        RECT 74.905 116.090 75.045 121.210 ;
        RECT 75.825 120.850 75.965 123.590 ;
        RECT 76.285 121.190 76.425 135.150 ;
        RECT 76.685 134.130 76.945 134.450 ;
        RECT 78.125 134.310 78.265 140.735 ;
        RECT 78.525 140.250 78.785 140.570 ;
        RECT 78.585 139.890 78.725 140.250 ;
        RECT 78.525 139.570 78.785 139.890 ;
        RECT 78.585 138.870 78.725 139.570 ;
        RECT 78.525 138.550 78.785 138.870 ;
        RECT 81.805 138.530 81.945 145.010 ;
        RECT 82.205 142.290 82.465 142.610 ;
        RECT 81.745 138.210 82.005 138.530 ;
        RECT 82.265 137.850 82.405 142.290 ;
        RECT 82.725 140.570 82.865 145.690 ;
        RECT 85.885 145.350 86.145 145.670 ;
        RECT 85.945 143.630 86.085 145.350 ;
        RECT 83.125 143.310 83.385 143.630 ;
        RECT 85.885 143.310 86.145 143.630 ;
        RECT 82.665 140.250 82.925 140.570 ;
        RECT 82.725 138.190 82.865 140.250 ;
        RECT 82.665 137.870 82.925 138.190 ;
        RECT 82.205 137.530 82.465 137.850 ;
        RECT 83.185 137.590 83.325 143.310 ;
        RECT 85.945 142.950 86.085 143.310 ;
        RECT 85.885 142.630 86.145 142.950 ;
        RECT 85.945 140.910 86.085 142.630 ;
        RECT 86.405 141.250 86.545 147.970 ;
        RECT 88.645 145.690 88.905 146.010 ;
        RECT 89.565 145.690 89.825 146.010 ;
        RECT 88.185 143.310 88.445 143.630 ;
        RECT 87.265 142.290 87.525 142.610 ;
        RECT 86.345 140.930 86.605 141.250 ;
        RECT 85.885 140.590 86.145 140.910 ;
        RECT 83.585 139.910 83.845 140.230 ;
        RECT 83.645 138.870 83.785 139.910 ;
        RECT 83.585 138.550 83.845 138.870 ;
        RECT 82.725 137.510 83.325 137.590 ;
        RECT 82.665 137.450 83.325 137.510 ;
        RECT 82.665 137.190 82.925 137.450 ;
        RECT 80.365 136.850 80.625 137.170 ;
        RECT 79.905 134.810 80.165 135.130 ;
        RECT 77.665 134.170 78.265 134.310 ;
        RECT 76.225 120.870 76.485 121.190 ;
        RECT 75.765 120.530 76.025 120.850 ;
        RECT 76.225 118.830 76.485 119.150 ;
        RECT 75.765 118.490 76.025 118.810 ;
        RECT 72.545 115.770 72.805 116.090 ;
        RECT 74.845 116.000 75.105 116.090 ;
        RECT 74.845 115.860 75.505 116.000 ;
        RECT 74.845 115.770 75.105 115.860 ;
        RECT 72.605 113.710 72.745 115.770 ;
        RECT 72.545 113.390 72.805 113.710 ;
        RECT 71.165 113.225 71.425 113.370 ;
        RECT 71.155 112.855 71.435 113.225 ;
        RECT 71.625 113.050 71.885 113.370 ;
        RECT 73.465 113.050 73.725 113.370 ;
        RECT 71.685 112.690 71.825 113.050 ;
        RECT 71.625 112.370 71.885 112.690 ;
        RECT 73.005 109.650 73.265 109.970 ;
        RECT 73.065 108.270 73.205 109.650 ;
        RECT 73.005 107.950 73.265 108.270 ;
        RECT 69.775 107.415 70.055 107.785 ;
        RECT 68.865 105.570 69.125 105.890 ;
        RECT 73.525 105.630 73.665 113.050 ;
        RECT 75.365 107.930 75.505 115.860 ;
        RECT 75.825 114.390 75.965 118.490 ;
        RECT 76.285 117.305 76.425 118.830 ;
        RECT 76.215 116.935 76.495 117.305 ;
        RECT 76.745 116.625 76.885 134.130 ;
        RECT 77.665 122.210 77.805 134.170 ;
        RECT 79.965 129.010 80.105 134.810 ;
        RECT 79.905 128.690 80.165 129.010 ;
        RECT 78.515 126.455 78.795 126.825 ;
        RECT 79.445 126.650 79.705 126.970 ;
        RECT 77.605 121.890 77.865 122.210 ;
        RECT 78.585 121.530 78.725 126.455 ;
        RECT 78.985 126.310 79.245 126.630 ;
        RECT 79.045 124.590 79.185 126.310 ;
        RECT 79.505 125.270 79.645 126.650 ;
        RECT 79.445 124.950 79.705 125.270 ;
        RECT 78.985 124.270 79.245 124.590 ;
        RECT 79.045 122.550 79.185 124.270 ;
        RECT 79.965 123.910 80.105 128.690 ;
        RECT 79.905 123.590 80.165 123.910 ;
        RECT 78.985 122.230 79.245 122.550 ;
        RECT 78.525 121.210 78.785 121.530 ;
        RECT 79.045 118.810 79.185 122.230 ;
        RECT 79.905 121.210 80.165 121.530 ;
        RECT 78.985 118.490 79.245 118.810 ;
        RECT 79.445 117.810 79.705 118.130 ;
        RECT 76.675 116.255 76.955 116.625 ;
        RECT 76.225 115.090 76.485 115.410 ;
        RECT 76.285 114.390 76.425 115.090 ;
        RECT 75.765 114.070 76.025 114.390 ;
        RECT 76.225 114.070 76.485 114.390 ;
        RECT 79.505 113.710 79.645 117.810 ;
        RECT 79.445 113.390 79.705 113.710 ;
        RECT 79.965 113.225 80.105 121.210 ;
        RECT 80.425 113.370 80.565 136.850 ;
        RECT 83.645 136.150 83.785 138.550 ;
        RECT 83.585 135.830 83.845 136.150 ;
        RECT 80.825 135.490 81.085 135.810 ;
        RECT 84.045 135.490 84.305 135.810 ;
        RECT 80.885 123.570 81.025 135.490 ;
        RECT 81.285 134.130 81.545 134.450 ;
        RECT 83.585 134.130 83.845 134.450 ;
        RECT 81.345 132.750 81.485 134.130 ;
        RECT 82.665 133.110 82.925 133.430 ;
        RECT 81.285 132.430 81.545 132.750 ;
        RECT 82.725 127.650 82.865 133.110 ;
        RECT 83.125 132.090 83.385 132.410 ;
        RECT 83.185 130.030 83.325 132.090 ;
        RECT 83.125 129.710 83.385 130.030 ;
        RECT 82.665 127.330 82.925 127.650 ;
        RECT 83.645 127.310 83.785 134.130 ;
        RECT 84.105 130.030 84.245 135.490 ;
        RECT 85.425 134.130 85.685 134.450 ;
        RECT 84.045 129.710 84.305 130.030 ;
        RECT 83.585 126.990 83.845 127.310 ;
        RECT 83.645 124.590 83.785 126.990 ;
        RECT 84.045 124.610 84.305 124.930 ;
        RECT 85.485 124.670 85.625 134.130 ;
        RECT 85.885 126.650 86.145 126.970 ;
        RECT 85.945 125.270 86.085 126.650 ;
        RECT 86.405 125.465 86.545 140.930 ;
        RECT 86.805 139.570 87.065 139.890 ;
        RECT 86.865 138.190 87.005 139.570 ;
        RECT 86.805 137.870 87.065 138.190 ;
        RECT 87.325 135.130 87.465 142.290 ;
        RECT 87.725 140.250 87.985 140.570 ;
        RECT 87.265 134.985 87.525 135.130 ;
        RECT 87.255 134.615 87.535 134.985 ;
        RECT 87.265 127.330 87.525 127.650 ;
        RECT 85.885 124.950 86.145 125.270 ;
        RECT 86.335 125.095 86.615 125.465 ;
        RECT 83.585 124.270 83.845 124.590 ;
        RECT 83.125 123.930 83.385 124.250 ;
        RECT 80.825 123.250 81.085 123.570 ;
        RECT 80.885 119.830 81.025 123.250 ;
        RECT 83.185 122.210 83.325 123.930 ;
        RECT 83.125 121.890 83.385 122.210 ;
        RECT 84.105 121.530 84.245 124.610 ;
        RECT 85.485 124.530 86.085 124.670 ;
        RECT 84.505 123.250 84.765 123.570 ;
        RECT 84.565 121.870 84.705 123.250 ;
        RECT 84.505 121.550 84.765 121.870 ;
        RECT 84.965 121.550 85.225 121.870 ;
        RECT 84.045 121.210 84.305 121.530 ;
        RECT 85.025 121.190 85.165 121.550 ;
        RECT 84.965 120.870 85.225 121.190 ;
        RECT 81.285 120.530 81.545 120.850 ;
        RECT 84.505 120.530 84.765 120.850 ;
        RECT 80.825 119.510 81.085 119.830 ;
        RECT 80.825 117.810 81.085 118.130 ;
        RECT 80.885 113.710 81.025 117.810 ;
        RECT 80.825 113.390 81.085 113.710 ;
        RECT 81.345 113.370 81.485 120.530 ;
        RECT 84.045 118.490 84.305 118.810 ;
        RECT 83.585 118.150 83.845 118.470 ;
        RECT 83.645 116.090 83.785 118.150 ;
        RECT 84.105 118.130 84.245 118.490 ;
        RECT 84.045 117.810 84.305 118.130 ;
        RECT 84.105 116.770 84.245 117.810 ;
        RECT 84.045 116.450 84.305 116.770 ;
        RECT 83.585 115.770 83.845 116.090 ;
        RECT 84.045 115.090 84.305 115.410 ;
        RECT 75.765 112.710 76.025 113.030 ;
        RECT 79.895 112.855 80.175 113.225 ;
        RECT 80.365 113.050 80.625 113.370 ;
        RECT 81.285 113.050 81.545 113.370 ;
        RECT 83.585 113.050 83.845 113.370 ;
        RECT 75.825 110.990 75.965 112.710 ;
        RECT 79.965 110.990 80.105 112.855 ;
        RECT 80.825 112.710 81.085 113.030 ;
        RECT 75.765 110.670 76.025 110.990 ;
        RECT 79.905 110.670 80.165 110.990 ;
        RECT 77.145 109.650 77.405 109.970 ;
        RECT 77.205 108.270 77.345 109.650 ;
        RECT 77.145 107.950 77.405 108.270 ;
        RECT 75.305 107.610 75.565 107.930 ;
        RECT 74.845 106.930 75.105 107.250 ;
        RECT 74.905 106.230 75.045 106.930 ;
        RECT 74.845 105.910 75.105 106.230 ;
        RECT 73.525 105.550 74.125 105.630 ;
        RECT 59.665 105.230 59.925 105.550 ;
        RECT 63.345 105.230 63.605 105.550 ;
        RECT 73.525 105.490 74.185 105.550 ;
        RECT 73.925 105.230 74.185 105.490 ;
        RECT 60.125 104.890 60.385 105.210 ;
        RECT 56.505 103.675 58.045 104.045 ;
        RECT 54.605 103.190 54.865 103.510 ;
        RECT 53.225 102.400 53.485 102.490 ;
        RECT 52.825 102.260 53.485 102.400 ;
        RECT 53.225 102.170 53.485 102.260 ;
        RECT 53.205 100.955 54.745 101.325 ;
        RECT 60.185 98.340 60.325 104.890 ;
        RECT 63.405 103.510 63.545 105.230 ;
        RECT 75.365 105.210 75.505 107.610 ;
        RECT 79.445 105.570 79.705 105.890 ;
        RECT 78.065 105.230 78.325 105.550 ;
        RECT 75.305 104.890 75.565 105.210 ;
        RECT 63.345 103.190 63.605 103.510 ;
        RECT 50.455 96.340 50.735 98.340 ;
        RECT 60.115 96.340 60.395 98.340 ;
        RECT 78.125 98.150 78.265 105.230 ;
        RECT 79.505 103.510 79.645 105.570 ;
        RECT 79.445 103.190 79.705 103.510 ;
        RECT 80.885 102.490 81.025 112.710 ;
        RECT 83.645 106.230 83.785 113.050 ;
        RECT 84.105 110.990 84.245 115.090 ;
        RECT 84.565 113.370 84.705 120.530 ;
        RECT 85.945 113.370 86.085 124.530 ;
        RECT 86.345 124.270 86.605 124.590 ;
        RECT 86.405 122.550 86.545 124.270 ;
        RECT 86.795 123.735 87.075 124.105 ;
        RECT 86.345 122.230 86.605 122.550 ;
        RECT 86.345 121.550 86.605 121.870 ;
        RECT 86.405 118.810 86.545 121.550 ;
        RECT 86.345 118.490 86.605 118.810 ;
        RECT 86.405 117.110 86.545 118.490 ;
        RECT 86.345 116.790 86.605 117.110 ;
        RECT 84.505 113.050 84.765 113.370 ;
        RECT 85.885 113.050 86.145 113.370 ;
        RECT 84.505 112.370 84.765 112.690 ;
        RECT 86.345 112.370 86.605 112.690 ;
        RECT 84.045 110.670 84.305 110.990 ;
        RECT 83.585 105.910 83.845 106.230 ;
        RECT 84.565 105.890 84.705 112.370 ;
        RECT 86.405 111.330 86.545 112.370 ;
        RECT 86.345 111.010 86.605 111.330 ;
        RECT 86.865 107.930 87.005 123.735 ;
        RECT 87.325 119.830 87.465 127.330 ;
        RECT 87.785 125.270 87.925 140.250 ;
        RECT 87.725 124.950 87.985 125.270 ;
        RECT 88.245 124.930 88.385 143.310 ;
        RECT 88.705 127.990 88.845 145.690 ;
        RECT 89.105 137.530 89.365 137.850 ;
        RECT 89.165 132.750 89.305 137.530 ;
        RECT 89.105 132.430 89.365 132.750 ;
        RECT 89.625 130.030 89.765 145.690 ;
        RECT 90.025 143.990 90.285 144.310 ;
        RECT 90.085 140.910 90.225 143.990 ;
        RECT 90.545 143.630 90.685 160.310 ;
        RECT 91.005 159.950 91.145 168.130 ;
        RECT 93.305 167.770 93.445 169.490 ;
        RECT 94.225 168.790 94.365 170.170 ;
        RECT 97.385 169.490 97.645 169.810 ;
        RECT 97.905 169.720 98.045 173.230 ;
        RECT 97.905 169.580 98.505 169.720 ;
        RECT 95.375 168.955 96.915 169.325 ;
        RECT 94.165 168.470 94.425 168.790 ;
        RECT 93.705 167.790 93.965 168.110 ;
        RECT 91.395 167.255 91.675 167.625 ;
        RECT 93.245 167.450 93.505 167.770 ;
        RECT 91.465 160.145 91.605 167.255 ;
        RECT 92.075 166.235 93.615 166.605 ;
        RECT 92.075 160.795 93.615 161.165 ;
        RECT 90.945 159.630 91.205 159.950 ;
        RECT 91.395 159.775 91.675 160.145 ;
        RECT 91.005 158.930 91.145 159.630 ;
        RECT 90.945 158.610 91.205 158.930 ;
        RECT 91.465 157.990 91.605 159.775 ;
        RECT 91.005 157.850 91.605 157.990 ;
        RECT 91.005 144.310 91.145 157.850 ;
        RECT 93.765 157.230 93.905 167.790 ;
        RECT 97.445 165.730 97.585 169.490 ;
        RECT 98.365 168.110 98.505 169.580 ;
        RECT 98.305 167.790 98.565 168.110 ;
        RECT 97.845 167.110 98.105 167.430 ;
        RECT 97.905 165.730 98.045 167.110 ;
        RECT 97.385 165.410 97.645 165.730 ;
        RECT 97.845 165.410 98.105 165.730 ;
        RECT 95.375 163.515 96.915 163.885 ;
        RECT 96.005 162.350 96.265 162.670 ;
        RECT 97.385 162.350 97.645 162.670 ;
        RECT 96.065 159.610 96.205 162.350 ;
        RECT 96.925 161.330 97.185 161.650 ;
        RECT 97.445 161.390 97.585 162.350 ;
        RECT 97.905 161.990 98.045 165.410 ;
        RECT 97.845 161.670 98.105 161.990 ;
        RECT 98.365 161.390 98.505 167.790 ;
        RECT 99.225 164.730 99.485 165.050 ;
        RECT 99.285 162.330 99.425 164.730 ;
        RECT 99.225 162.010 99.485 162.330 ;
        RECT 96.985 159.950 97.125 161.330 ;
        RECT 97.445 161.250 98.505 161.390 ;
        RECT 96.925 159.630 97.185 159.950 ;
        RECT 96.005 159.290 96.265 159.610 ;
        RECT 97.385 159.290 97.645 159.610 ;
        RECT 94.625 158.610 94.885 158.930 ;
        RECT 93.705 156.910 93.965 157.230 ;
        RECT 91.405 156.570 91.665 156.890 ;
        RECT 91.465 154.170 91.605 156.570 ;
        RECT 92.075 155.355 93.615 155.725 ;
        RECT 91.405 153.850 91.665 154.170 ;
        RECT 93.765 152.470 93.905 156.910 ;
        RECT 94.685 156.890 94.825 158.610 ;
        RECT 95.375 158.075 96.915 158.445 ;
        RECT 97.445 157.570 97.585 159.290 ;
        RECT 97.385 157.250 97.645 157.570 ;
        RECT 94.625 156.570 94.885 156.890 ;
        RECT 96.925 155.890 97.185 156.210 ;
        RECT 95.085 154.530 95.345 154.850 ;
        RECT 95.145 153.740 95.285 154.530 ;
        RECT 96.985 154.510 97.125 155.890 ;
        RECT 96.925 154.190 97.185 154.510 ;
        RECT 94.685 153.600 95.285 153.740 ;
        RECT 94.685 152.470 94.825 153.600 ;
        RECT 95.375 152.635 96.915 153.005 ;
        RECT 93.705 152.150 93.965 152.470 ;
        RECT 94.625 152.150 94.885 152.470 ;
        RECT 93.705 150.790 93.965 151.110 ;
        RECT 92.075 149.915 93.615 150.285 ;
        RECT 91.405 145.690 91.665 146.010 ;
        RECT 90.945 143.990 91.205 144.310 ;
        RECT 91.465 143.970 91.605 145.690 ;
        RECT 93.765 145.670 93.905 150.790 ;
        RECT 95.375 147.195 96.915 147.565 ;
        RECT 93.705 145.350 93.965 145.670 ;
        RECT 92.075 144.475 93.615 144.845 ;
        RECT 91.405 143.650 91.665 143.970 ;
        RECT 92.325 143.650 92.585 143.970 ;
        RECT 90.485 143.540 90.745 143.630 ;
        RECT 90.485 143.400 91.145 143.540 ;
        RECT 90.485 143.310 90.745 143.400 ;
        RECT 90.025 140.820 90.285 140.910 ;
        RECT 90.025 140.680 90.685 140.820 ;
        RECT 90.025 140.590 90.285 140.680 ;
        RECT 90.025 139.910 90.285 140.230 ;
        RECT 90.085 137.510 90.225 139.910 ;
        RECT 90.545 138.190 90.685 140.680 ;
        RECT 91.005 140.570 91.145 143.400 ;
        RECT 92.385 140.570 92.525 143.650 ;
        RECT 90.945 140.250 91.205 140.570 ;
        RECT 92.325 140.250 92.585 140.570 ;
        RECT 90.945 139.570 91.205 139.890 ;
        RECT 92.385 139.800 92.525 140.250 ;
        RECT 91.465 139.660 92.525 139.800 ;
        RECT 90.485 137.870 90.745 138.190 ;
        RECT 90.025 137.190 90.285 137.510 ;
        RECT 90.085 135.470 90.225 137.190 ;
        RECT 90.485 136.850 90.745 137.170 ;
        RECT 90.025 135.150 90.285 135.470 ;
        RECT 89.565 129.710 89.825 130.030 ;
        RECT 89.105 129.030 89.365 129.350 ;
        RECT 88.645 127.670 88.905 127.990 ;
        RECT 88.185 124.610 88.445 124.930 ;
        RECT 87.725 123.930 87.985 124.250 ;
        RECT 87.785 122.550 87.925 123.930 ;
        RECT 88.245 123.570 88.385 124.610 ;
        RECT 88.185 123.250 88.445 123.570 ;
        RECT 88.645 123.250 88.905 123.570 ;
        RECT 87.725 122.230 87.985 122.550 ;
        RECT 87.785 121.870 87.925 122.230 ;
        RECT 88.245 121.870 88.385 123.250 ;
        RECT 88.705 121.870 88.845 123.250 ;
        RECT 87.725 121.550 87.985 121.870 ;
        RECT 88.185 121.550 88.445 121.870 ;
        RECT 88.645 121.550 88.905 121.870 ;
        RECT 87.265 119.510 87.525 119.830 ;
        RECT 87.265 118.830 87.525 119.150 ;
        RECT 88.635 118.975 88.915 119.345 ;
        RECT 87.325 113.710 87.465 118.830 ;
        RECT 88.705 118.810 88.845 118.975 ;
        RECT 88.645 118.490 88.905 118.810 ;
        RECT 88.645 117.810 88.905 118.130 ;
        RECT 88.705 117.110 88.845 117.810 ;
        RECT 88.645 116.790 88.905 117.110 ;
        RECT 87.265 113.390 87.525 113.710 ;
        RECT 88.185 113.390 88.445 113.710 ;
        RECT 87.725 110.670 87.985 110.990 ;
        RECT 87.785 108.950 87.925 110.670 ;
        RECT 88.245 109.970 88.385 113.390 ;
        RECT 89.165 113.370 89.305 129.030 ;
        RECT 90.025 125.970 90.285 126.290 ;
        RECT 89.565 124.610 89.825 124.930 ;
        RECT 89.625 124.250 89.765 124.610 ;
        RECT 89.565 123.930 89.825 124.250 ;
        RECT 89.565 121.210 89.825 121.530 ;
        RECT 89.625 118.810 89.765 121.210 ;
        RECT 89.565 118.490 89.825 118.810 ;
        RECT 90.085 116.770 90.225 125.970 ;
        RECT 90.545 117.110 90.685 136.850 ;
        RECT 90.485 116.790 90.745 117.110 ;
        RECT 90.025 116.450 90.285 116.770 ;
        RECT 90.475 116.255 90.755 116.625 ;
        RECT 91.005 116.430 91.145 139.570 ;
        RECT 91.465 138.270 91.605 139.660 ;
        RECT 92.075 139.035 93.615 139.405 ;
        RECT 91.465 138.130 92.525 138.270 ;
        RECT 91.865 137.870 92.125 138.130 ;
        RECT 91.865 137.190 92.125 137.510 ;
        RECT 91.925 135.130 92.065 137.190 ;
        RECT 92.385 135.130 92.525 138.130 ;
        RECT 91.865 134.810 92.125 135.130 ;
        RECT 92.325 134.810 92.585 135.130 ;
        RECT 92.075 133.595 93.615 133.965 ;
        RECT 92.325 132.430 92.585 132.750 ;
        RECT 92.385 129.690 92.525 132.430 ;
        RECT 92.325 129.600 92.585 129.690 ;
        RECT 91.465 129.460 92.585 129.600 ;
        RECT 91.465 127.310 91.605 129.460 ;
        RECT 92.325 129.370 92.585 129.460 ;
        RECT 92.075 128.155 93.615 128.525 ;
        RECT 92.325 127.670 92.585 127.990 ;
        RECT 91.405 126.990 91.665 127.310 ;
        RECT 92.385 123.570 92.525 127.670 ;
        RECT 93.245 126.650 93.505 126.970 ;
        RECT 92.785 126.310 93.045 126.630 ;
        RECT 91.405 123.250 91.665 123.570 ;
        RECT 92.325 123.250 92.585 123.570 ;
        RECT 92.845 123.480 92.985 126.310 ;
        RECT 93.305 124.590 93.445 126.650 ;
        RECT 93.765 124.930 93.905 145.350 ;
        RECT 94.625 145.010 94.885 145.330 ;
        RECT 97.385 145.010 97.645 145.330 ;
        RECT 94.685 144.310 94.825 145.010 ;
        RECT 97.445 144.310 97.585 145.010 ;
        RECT 94.625 143.990 94.885 144.310 ;
        RECT 97.385 143.990 97.645 144.310 ;
        RECT 94.165 143.650 94.425 143.970 ;
        RECT 94.225 135.040 94.365 143.650 ;
        RECT 94.685 141.250 94.825 143.990 ;
        RECT 95.375 141.755 96.915 142.125 ;
        RECT 94.625 140.930 94.885 141.250 ;
        RECT 97.445 140.910 97.585 143.990 ;
        RECT 97.905 143.290 98.045 161.250 ;
        RECT 98.305 159.970 98.565 160.290 ;
        RECT 98.365 157.910 98.505 159.970 ;
        RECT 98.765 158.610 99.025 158.930 ;
        RECT 98.305 157.590 98.565 157.910 ;
        RECT 98.825 157.230 98.965 158.610 ;
        RECT 98.765 156.910 99.025 157.230 ;
        RECT 99.285 156.210 99.425 162.010 ;
        RECT 99.685 159.630 99.945 159.950 ;
        RECT 99.745 156.890 99.885 159.630 ;
        RECT 99.685 156.570 99.945 156.890 ;
        RECT 99.225 155.890 99.485 156.210 ;
        RECT 98.765 154.080 99.025 154.170 ;
        RECT 99.285 154.080 99.425 155.890 ;
        RECT 98.765 153.940 99.425 154.080 ;
        RECT 98.765 153.850 99.025 153.940 ;
        RECT 98.825 149.070 98.965 153.850 ;
        RECT 98.765 148.750 99.025 149.070 ;
        RECT 100.205 148.980 100.345 183.090 ;
        RECT 101.065 178.330 101.325 178.650 ;
        RECT 100.605 176.630 100.865 176.950 ;
        RECT 100.665 174.230 100.805 176.630 ;
        RECT 100.605 173.910 100.865 174.230 ;
        RECT 101.125 170.830 101.265 178.330 ;
        RECT 101.985 177.650 102.245 177.970 ;
        RECT 102.045 176.610 102.185 177.650 ;
        RECT 101.985 176.290 102.245 176.610 ;
        RECT 109.345 175.610 109.605 175.930 ;
        RECT 109.405 173.550 109.545 175.610 ;
        RECT 109.345 173.230 109.605 173.550 ;
        RECT 135.630 173.380 136.780 174.600 ;
        RECT 105.665 172.550 105.925 172.870 ;
        RECT 101.985 172.210 102.245 172.530 ;
        RECT 101.065 170.510 101.325 170.830 ;
        RECT 102.045 167.770 102.185 172.210 ;
        RECT 105.725 171.510 105.865 172.550 ;
        RECT 105.665 171.190 105.925 171.510 ;
        RECT 106.125 170.510 106.385 170.830 ;
        RECT 106.185 167.770 106.325 170.510 ;
        RECT 101.985 167.450 102.245 167.770 ;
        RECT 106.125 167.450 106.385 167.770 ;
        RECT 103.825 166.770 104.085 167.090 ;
        RECT 105.665 166.770 105.925 167.090 ;
        RECT 103.885 165.050 104.025 166.770 ;
        RECT 105.725 165.730 105.865 166.770 ;
        RECT 106.185 166.070 106.325 167.450 ;
        RECT 106.125 165.750 106.385 166.070 ;
        RECT 105.665 165.410 105.925 165.730 ;
        RECT 103.825 164.730 104.085 165.050 ;
        RECT 105.665 161.670 105.925 161.990 ;
        RECT 100.605 161.330 100.865 161.650 ;
        RECT 100.665 159.950 100.805 161.330 ;
        RECT 105.725 160.630 105.865 161.670 ;
        RECT 105.665 160.310 105.925 160.630 ;
        RECT 100.605 159.630 100.865 159.950 ;
        RECT 101.515 159.775 101.795 160.145 ;
        RECT 106.185 160.030 106.325 165.750 ;
        RECT 109.405 165.050 109.545 173.230 ;
        RECT 133.750 170.070 134.880 172.730 ;
        RECT 135.630 166.640 136.740 173.380 ;
        RECT 135.630 165.420 136.780 166.640 ;
        RECT 109.345 164.730 109.605 165.050 ;
        RECT 109.405 162.330 109.545 164.730 ;
        RECT 109.345 162.010 109.605 162.330 ;
        RECT 105.725 159.950 106.325 160.030 ;
        RECT 105.665 159.890 106.325 159.950 ;
        RECT 101.525 159.630 101.785 159.775 ;
        RECT 105.665 159.630 105.925 159.890 ;
        RECT 103.825 158.610 104.085 158.930 ;
        RECT 103.885 156.550 104.025 158.610 ;
        RECT 103.825 156.230 104.085 156.550 ;
        RECT 101.985 153.850 102.245 154.170 ;
        RECT 102.045 152.130 102.185 153.850 ;
        RECT 101.985 151.810 102.245 152.130 ;
        RECT 105.725 151.450 105.865 159.630 ;
        RECT 109.405 156.890 109.545 162.010 ;
        RECT 109.345 156.570 109.605 156.890 ;
        RECT 110.715 155.015 110.995 155.385 ;
        RECT 110.785 154.850 110.925 155.015 ;
        RECT 107.045 154.530 107.305 154.850 ;
        RECT 110.725 154.530 110.985 154.850 ;
        RECT 107.105 152.470 107.245 154.530 ;
        RECT 107.045 152.150 107.305 152.470 ;
        RECT 105.665 151.130 105.925 151.450 ;
        RECT 100.205 148.840 100.805 148.980 ;
        RECT 100.145 148.070 100.405 148.390 ;
        RECT 100.205 145.670 100.345 148.070 ;
        RECT 100.145 145.350 100.405 145.670 ;
        RECT 99.225 143.310 99.485 143.630 ;
        RECT 97.845 142.970 98.105 143.290 ;
        RECT 97.385 140.590 97.645 140.910 ;
        RECT 95.085 140.250 95.345 140.570 ;
        RECT 94.625 139.570 94.885 139.890 ;
        RECT 94.685 137.510 94.825 139.570 ;
        RECT 95.145 138.870 95.285 140.250 ;
        RECT 95.085 138.780 95.345 138.870 ;
        RECT 95.085 138.640 96.205 138.780 ;
        RECT 95.085 138.550 95.345 138.640 ;
        RECT 96.065 137.850 96.205 138.640 ;
        RECT 96.005 137.530 96.265 137.850 ;
        RECT 94.625 137.190 94.885 137.510 ;
        RECT 95.375 136.315 96.915 136.685 ;
        RECT 97.445 135.470 97.585 140.590 ;
        RECT 97.905 140.570 98.045 142.970 ;
        RECT 99.285 141.250 99.425 143.310 ;
        RECT 99.685 142.970 99.945 143.290 ;
        RECT 99.225 140.930 99.485 141.250 ;
        RECT 98.765 140.590 99.025 140.910 ;
        RECT 97.845 140.250 98.105 140.570 ;
        RECT 98.825 138.870 98.965 140.590 ;
        RECT 98.765 138.550 99.025 138.870 ;
        RECT 99.745 138.190 99.885 142.970 ;
        RECT 100.145 139.910 100.405 140.230 ;
        RECT 99.685 137.870 99.945 138.190 ;
        RECT 97.385 135.150 97.645 135.470 ;
        RECT 95.085 135.040 95.345 135.130 ;
        RECT 94.225 134.900 95.345 135.040 ;
        RECT 94.225 134.450 94.365 134.900 ;
        RECT 95.085 134.810 95.345 134.900 ;
        RECT 94.165 134.130 94.425 134.450 ;
        RECT 97.845 134.130 98.105 134.450 ;
        RECT 94.625 132.770 94.885 133.090 ;
        RECT 97.385 132.770 97.645 133.090 ;
        RECT 94.165 132.090 94.425 132.410 ;
        RECT 94.225 128.070 94.365 132.090 ;
        RECT 94.685 129.010 94.825 132.770 ;
        RECT 95.375 130.875 96.915 131.245 ;
        RECT 95.085 129.710 95.345 130.030 ;
        RECT 94.625 128.690 94.885 129.010 ;
        RECT 94.225 127.930 94.825 128.070 ;
        RECT 94.165 126.990 94.425 127.310 ;
        RECT 93.705 124.610 93.965 124.930 ;
        RECT 93.245 124.270 93.505 124.590 ;
        RECT 92.845 123.340 93.905 123.480 ;
        RECT 91.465 116.680 91.605 123.250 ;
        RECT 92.075 122.715 93.615 123.085 ;
        RECT 91.865 121.550 92.125 121.870 ;
        RECT 92.785 121.780 93.045 121.870 ;
        RECT 93.765 121.780 93.905 123.340 ;
        RECT 92.785 121.640 93.905 121.780 ;
        RECT 92.785 121.550 93.045 121.640 ;
        RECT 91.925 118.470 92.065 121.550 ;
        RECT 92.325 120.530 92.585 120.850 ;
        RECT 92.385 119.150 92.525 120.530 ;
        RECT 92.845 119.490 92.985 121.550 ;
        RECT 93.705 119.510 93.965 119.830 ;
        RECT 92.785 119.170 93.045 119.490 ;
        RECT 92.325 118.830 92.585 119.150 ;
        RECT 92.385 118.665 92.525 118.830 ;
        RECT 93.765 118.810 93.905 119.510 ;
        RECT 94.225 119.150 94.365 126.990 ;
        RECT 94.685 126.290 94.825 127.930 ;
        RECT 95.145 127.310 95.285 129.710 ;
        RECT 95.545 128.690 95.805 129.010 ;
        RECT 95.605 127.310 95.745 128.690 ;
        RECT 95.085 126.990 95.345 127.310 ;
        RECT 95.545 126.990 95.805 127.310 ;
        RECT 95.145 126.630 95.285 126.990 ;
        RECT 95.605 126.825 95.745 126.990 ;
        RECT 95.085 126.310 95.345 126.630 ;
        RECT 95.535 126.455 95.815 126.825 ;
        RECT 94.625 125.970 94.885 126.290 ;
        RECT 94.685 121.530 94.825 125.970 ;
        RECT 95.375 125.435 96.915 125.805 ;
        RECT 97.445 124.930 97.585 132.770 ;
        RECT 97.385 124.610 97.645 124.930 ;
        RECT 95.085 123.250 95.345 123.570 ;
        RECT 96.465 123.250 96.725 123.570 ;
        RECT 95.145 121.870 95.285 123.250 ;
        RECT 96.525 122.210 96.665 123.250 ;
        RECT 96.465 121.890 96.725 122.210 ;
        RECT 95.085 121.550 95.345 121.870 ;
        RECT 97.385 121.550 97.645 121.870 ;
        RECT 94.625 121.210 94.885 121.530 ;
        RECT 94.625 120.530 94.885 120.850 ;
        RECT 94.165 118.830 94.425 119.150 ;
        RECT 91.865 118.150 92.125 118.470 ;
        RECT 92.315 118.295 92.595 118.665 ;
        RECT 93.705 118.490 93.965 118.810 ;
        RECT 92.075 117.275 93.615 117.645 ;
        RECT 91.865 116.680 92.125 116.770 ;
        RECT 91.465 116.540 92.125 116.680 ;
        RECT 91.865 116.450 92.125 116.540 ;
        RECT 93.765 116.430 93.905 118.490 ;
        RECT 90.545 116.090 90.685 116.255 ;
        RECT 90.945 116.110 91.205 116.430 ;
        RECT 93.705 116.110 93.965 116.430 ;
        RECT 90.485 115.770 90.745 116.090 ;
        RECT 91.865 115.430 92.125 115.750 ;
        RECT 91.925 114.390 92.065 115.430 ;
        RECT 91.865 114.070 92.125 114.390 ;
        RECT 93.705 113.390 93.965 113.710 ;
        RECT 89.105 113.050 89.365 113.370 ;
        RECT 91.405 112.370 91.665 112.690 ;
        RECT 90.945 110.670 91.205 110.990 ;
        RECT 88.185 109.650 88.445 109.970 ;
        RECT 90.025 109.650 90.285 109.970 ;
        RECT 87.725 108.630 87.985 108.950 ;
        RECT 88.245 108.610 88.385 109.650 ;
        RECT 88.185 108.290 88.445 108.610 ;
        RECT 90.085 107.930 90.225 109.650 ;
        RECT 91.005 108.270 91.145 110.670 ;
        RECT 90.945 107.950 91.205 108.270 ;
        RECT 91.465 107.930 91.605 112.370 ;
        RECT 92.075 111.835 93.615 112.205 ;
        RECT 93.765 110.650 93.905 113.390 ;
        RECT 94.225 110.990 94.365 118.830 ;
        RECT 94.685 116.090 94.825 120.530 ;
        RECT 95.375 119.995 96.915 120.365 ;
        RECT 96.005 118.380 96.265 118.470 ;
        RECT 97.445 118.380 97.585 121.550 ;
        RECT 96.005 118.240 97.585 118.380 ;
        RECT 96.005 118.150 96.265 118.240 ;
        RECT 96.065 117.110 96.205 118.150 ;
        RECT 97.905 117.110 98.045 134.130 ;
        RECT 99.225 132.770 99.485 133.090 ;
        RECT 98.765 129.030 99.025 129.350 ;
        RECT 98.825 127.990 98.965 129.030 ;
        RECT 98.765 127.670 99.025 127.990 ;
        RECT 98.765 124.950 99.025 125.270 ;
        RECT 96.005 116.790 96.265 117.110 ;
        RECT 97.845 116.790 98.105 117.110 ;
        RECT 98.825 116.430 98.965 124.950 ;
        RECT 99.285 117.110 99.425 132.770 ;
        RECT 99.745 132.750 99.885 137.870 ;
        RECT 100.205 136.150 100.345 139.910 ;
        RECT 100.145 135.830 100.405 136.150 ;
        RECT 100.665 135.665 100.805 148.840 ;
        RECT 101.525 148.750 101.785 149.070 ;
        RECT 101.585 146.350 101.725 148.750 ;
        RECT 107.505 148.410 107.765 148.730 ;
        RECT 101.525 146.030 101.785 146.350 ;
        RECT 101.585 136.150 101.725 146.030 ;
        RECT 107.565 146.010 107.705 148.410 ;
        RECT 103.825 145.690 104.085 146.010 ;
        RECT 106.125 145.690 106.385 146.010 ;
        RECT 107.505 145.690 107.765 146.010 ;
        RECT 103.885 144.310 104.025 145.690 ;
        RECT 105.205 145.010 105.465 145.330 ;
        RECT 105.265 144.310 105.405 145.010 ;
        RECT 103.825 143.990 104.085 144.310 ;
        RECT 105.205 143.990 105.465 144.310 ;
        RECT 106.185 143.290 106.325 145.690 ;
        RECT 106.585 145.010 106.845 145.330 ;
        RECT 106.645 143.970 106.785 145.010 ;
        RECT 106.585 143.650 106.845 143.970 ;
        RECT 106.125 142.970 106.385 143.290 ;
        RECT 106.185 140.910 106.325 142.970 ;
        RECT 106.125 140.590 106.385 140.910 ;
        RECT 107.045 138.210 107.305 138.530 ;
        RECT 107.105 136.150 107.245 138.210 ;
        RECT 101.525 135.830 101.785 136.150 ;
        RECT 107.045 135.830 107.305 136.150 ;
        RECT 100.595 135.295 100.875 135.665 ;
        RECT 100.665 135.130 100.805 135.295 ;
        RECT 100.605 134.810 100.865 135.130 ;
        RECT 99.685 132.430 99.945 132.750 ;
        RECT 100.605 132.430 100.865 132.750 ;
        RECT 99.685 131.410 99.945 131.730 ;
        RECT 99.745 127.310 99.885 131.410 ;
        RECT 100.665 130.030 100.805 132.430 ;
        RECT 100.605 129.710 100.865 130.030 ;
        RECT 99.685 126.990 99.945 127.310 ;
        RECT 100.605 126.310 100.865 126.630 ;
        RECT 100.665 124.590 100.805 126.310 ;
        RECT 100.605 124.270 100.865 124.590 ;
        RECT 101.585 121.870 101.725 135.830 ;
        RECT 107.565 135.130 107.705 145.690 ;
        RECT 110.715 144.815 110.995 145.185 ;
        RECT 110.785 143.630 110.925 144.815 ;
        RECT 110.725 143.310 110.985 143.630 ;
        RECT 110.715 141.415 110.995 141.785 ;
        RECT 110.785 138.530 110.925 141.415 ;
        RECT 135.630 141.200 136.780 141.270 ;
        RECT 135.630 140.180 136.800 141.200 ;
        RECT 110.725 138.210 110.985 138.530 ;
        RECT 132.560 138.140 135.160 140.060 ;
        RECT 107.505 134.810 107.765 135.130 ;
        RECT 105.205 134.470 105.465 134.790 ;
        RECT 110.715 134.615 110.995 134.985 ;
        RECT 103.825 129.710 104.085 130.030 ;
        RECT 102.905 129.030 103.165 129.350 ;
        RECT 102.965 127.990 103.105 129.030 ;
        RECT 102.905 127.670 103.165 127.990 ;
        RECT 103.885 124.590 104.025 129.710 ;
        RECT 105.265 129.690 105.405 134.470 ;
        RECT 110.785 133.090 110.925 134.615 ;
        RECT 135.640 133.320 136.800 140.180 ;
        RECT 105.665 132.770 105.925 133.090 ;
        RECT 110.725 132.770 110.985 133.090 ;
        RECT 105.725 130.710 105.865 132.770 ;
        RECT 105.665 130.390 105.925 130.710 ;
        RECT 105.205 129.370 105.465 129.690 ;
        RECT 105.265 127.650 105.405 129.370 ;
        RECT 105.205 127.330 105.465 127.650 ;
        RECT 103.825 124.270 104.085 124.590 ;
        RECT 102.905 123.590 103.165 123.910 ;
        RECT 102.965 122.550 103.105 123.590 ;
        RECT 103.825 123.250 104.085 123.570 ;
        RECT 103.885 122.550 104.025 123.250 ;
        RECT 102.905 122.230 103.165 122.550 ;
        RECT 103.825 122.230 104.085 122.550 ;
        RECT 101.525 121.550 101.785 121.870 ;
        RECT 101.585 119.345 101.725 121.550 ;
        RECT 100.145 118.830 100.405 119.150 ;
        RECT 101.515 118.975 101.795 119.345 ;
        RECT 99.225 116.790 99.485 117.110 ;
        RECT 98.765 116.110 99.025 116.430 ;
        RECT 94.625 115.770 94.885 116.090 ;
        RECT 98.305 115.770 98.565 116.090 ;
        RECT 95.375 114.555 96.915 114.925 ;
        RECT 95.085 113.050 95.345 113.370 ;
        RECT 94.165 110.670 94.425 110.990 ;
        RECT 93.705 110.330 93.965 110.650 ;
        RECT 86.805 107.610 87.065 107.930 ;
        RECT 90.025 107.610 90.285 107.930 ;
        RECT 91.405 107.610 91.665 107.930 ;
        RECT 85.885 106.930 86.145 107.250 ;
        RECT 85.945 105.890 86.085 106.930 ;
        RECT 92.075 106.395 93.615 106.765 ;
        RECT 84.505 105.570 84.765 105.890 ;
        RECT 85.885 105.570 86.145 105.890 ;
        RECT 94.225 105.120 94.365 110.670 ;
        RECT 95.145 110.310 95.285 113.050 ;
        RECT 97.845 112.710 98.105 113.030 ;
        RECT 96.465 112.370 96.725 112.690 ;
        RECT 96.525 111.330 96.665 112.370 ;
        RECT 96.465 111.010 96.725 111.330 ;
        RECT 95.085 109.990 95.345 110.310 ;
        RECT 95.375 109.115 96.915 109.485 ;
        RECT 97.905 108.610 98.045 112.710 ;
        RECT 98.365 110.310 98.505 115.770 ;
        RECT 100.205 113.710 100.345 118.830 ;
        RECT 104.745 118.150 105.005 118.470 ;
        RECT 104.805 117.110 104.945 118.150 ;
        RECT 104.745 116.790 105.005 117.110 ;
        RECT 105.265 116.430 105.405 127.330 ;
        RECT 101.065 116.110 101.325 116.430 ;
        RECT 105.205 116.110 105.465 116.430 ;
        RECT 99.685 113.390 99.945 113.710 ;
        RECT 100.145 113.390 100.405 113.710 ;
        RECT 99.745 111.670 99.885 113.390 ;
        RECT 99.685 111.350 99.945 111.670 ;
        RECT 101.125 111.330 101.265 116.110 ;
        RECT 101.065 111.010 101.325 111.330 ;
        RECT 105.265 110.990 105.405 116.110 ;
        RECT 105.205 110.670 105.465 110.990 ;
        RECT 98.305 109.990 98.565 110.310 ;
        RECT 98.365 108.950 98.505 109.990 ;
        RECT 98.305 108.630 98.565 108.950 ;
        RECT 97.845 108.290 98.105 108.610 ;
        RECT 105.265 107.930 105.405 110.670 ;
        RECT 105.205 107.610 105.465 107.930 ;
        RECT 129.750 105.580 133.160 106.650 ;
        RECT 94.625 105.120 94.885 105.210 ;
        RECT 94.225 104.980 94.885 105.120 ;
        RECT 94.625 104.890 94.885 104.980 ;
        RECT 82.665 104.210 82.925 104.530 ;
        RECT 80.825 102.170 81.085 102.490 ;
        RECT 79.045 98.690 79.645 98.830 ;
        RECT 79.045 98.150 79.185 98.690 ;
        RECT 79.505 98.340 79.645 98.690 ;
        RECT 82.725 98.340 82.865 104.210 ;
        RECT 95.375 103.675 96.915 104.045 ;
        RECT 92.075 100.955 93.615 101.325 ;
        RECT 78.125 98.010 79.185 98.150 ;
        RECT 79.435 96.340 79.715 98.340 ;
        RECT 82.655 96.340 82.935 98.340 ;
        RECT 13.920 85.550 15.140 89.420 ;
        RECT 19.910 85.980 21.130 89.850 ;
        RECT 67.730 89.640 68.670 89.840 ;
        RECT 25.730 85.120 26.950 88.990 ;
        RECT 31.780 85.510 33.000 89.380 ;
        RECT 37.750 88.780 38.970 89.290 ;
        RECT 37.680 88.620 38.970 88.780 ;
        RECT 43.810 88.630 45.030 89.530 ;
        RECT 49.740 88.640 50.960 89.040 ;
        RECT 37.680 86.810 39.070 88.620 ;
        RECT 37.750 85.420 38.970 86.810 ;
        RECT 43.810 86.720 45.140 88.630 ;
        RECT 49.740 86.920 51.010 88.640 ;
        RECT 43.810 85.660 45.030 86.720 ;
        RECT 49.740 85.170 50.960 86.920 ;
        RECT 55.530 85.320 56.750 89.190 ;
        RECT 61.720 88.640 62.940 88.870 ;
        RECT 61.720 86.600 63.130 88.640 ;
        RECT 61.720 85.000 62.940 86.600 ;
        RECT 67.580 85.770 68.800 89.640 ;
        RECT 73.850 84.290 75.070 88.160 ;
        RECT 79.730 84.310 80.950 88.180 ;
        RECT 74.090 80.440 74.370 84.290 ;
        RECT 20.140 80.160 74.370 80.440 ;
        RECT 20.140 75.650 20.420 80.160 ;
        RECT 80.070 79.800 80.350 84.310 ;
        RECT 85.470 84.100 86.690 87.970 ;
        RECT 91.460 84.500 92.680 88.320 ;
        RECT 97.600 84.630 98.820 88.240 ;
        RECT 103.650 84.740 104.870 88.610 ;
        RECT 109.620 85.420 110.840 89.290 ;
        RECT 115.740 85.700 116.960 89.570 ;
        RECT 121.520 85.700 122.740 89.570 ;
        RECT 31.380 79.520 80.350 79.800 ;
        RECT 31.380 75.850 31.660 79.520 ;
        RECT 86.050 79.170 86.330 84.100 ;
        RECT 42.510 78.890 86.330 79.170 ;
        RECT 3.960 71.320 6.050 73.240 ;
        RECT 19.330 73.120 21.890 75.650 ;
        RECT 28.185 73.180 30.255 74.460 ;
        RECT 30.670 73.320 33.230 75.850 ;
        RECT 42.510 75.750 42.790 78.890 ;
        RECT 92.030 78.570 92.310 84.500 ;
        RECT 53.830 78.290 92.310 78.570 ;
        RECT 53.830 75.820 54.110 78.290 ;
        RECT 98.010 77.990 98.290 84.630 ;
        RECT 64.900 77.710 98.290 77.990 ;
        RECT 19.005 71.800 19.865 72.640 ;
        RECT 15.560 68.610 16.990 71.210 ;
        RECT 19.305 68.570 19.845 71.800 ;
        RECT 20.145 70.600 20.555 73.120 ;
        RECT 30.205 71.810 31.065 72.650 ;
        RECT 19.325 47.770 19.825 68.570 ;
        RECT 20.165 49.090 20.555 70.600 ;
        RECT 20.955 70.010 21.845 70.740 ;
        RECT 21.055 65.190 21.315 70.010 ;
        RECT 22.695 68.620 25.405 69.470 ;
        RECT 22.895 65.840 24.825 68.620 ;
        RECT 30.505 68.580 31.045 71.810 ;
        RECT 31.345 70.610 31.755 73.320 ;
        RECT 39.475 73.150 41.545 74.430 ;
        RECT 41.910 73.220 44.470 75.750 ;
        RECT 41.425 71.780 42.285 72.620 ;
        RECT 27.795 67.130 28.915 67.810 ;
        RECT 28.075 65.850 28.745 67.130 ;
        RECT 21.455 65.460 26.505 65.840 ;
        RECT 27.865 65.440 28.915 65.850 ;
        RECT 21.055 63.640 21.435 65.190 ;
        RECT 21.175 55.800 21.435 63.640 ;
        RECT 26.485 63.200 26.755 65.240 ;
        RECT 27.615 63.200 27.885 65.200 ;
        RECT 26.485 56.510 27.885 63.200 ;
        RECT 21.085 55.290 21.445 55.800 ;
        RECT 21.065 54.860 21.445 55.290 ;
        RECT 26.485 55.190 26.755 56.510 ;
        RECT 27.615 55.150 27.885 56.510 ;
        RECT 28.885 55.260 29.205 65.190 ;
        RECT 28.885 55.200 29.215 55.260 ;
        RECT 21.065 54.580 21.315 54.860 ;
        RECT 20.865 54.180 25.505 54.580 ;
        RECT 26.405 54.290 27.535 54.300 ;
        RECT 28.895 54.290 29.215 55.200 ;
        RECT 21.065 52.060 21.315 54.180 ;
        RECT 25.765 53.490 26.125 54.110 ;
        RECT 25.845 52.610 26.105 53.490 ;
        RECT 26.385 53.240 29.215 54.290 ;
        RECT 25.675 52.230 26.205 52.610 ;
        RECT 21.065 51.970 21.565 52.060 ;
        RECT 21.055 51.240 21.565 51.970 ;
        RECT 21.295 50.240 21.565 51.240 ;
        RECT 22.205 50.990 22.475 51.940 ;
        RECT 22.205 50.840 22.675 50.990 ;
        RECT 22.205 50.160 22.765 50.840 ;
        RECT 22.285 50.150 22.765 50.160 ;
        RECT 21.575 49.620 22.195 49.980 ;
        RECT 21.615 49.090 22.045 49.620 ;
        RECT 20.165 48.670 22.045 49.090 ;
        RECT 22.535 48.960 22.765 50.150 ;
        RECT 21.615 47.800 22.045 48.670 ;
        RECT 22.455 48.360 22.835 48.960 ;
        RECT 19.325 47.060 20.015 47.770 ;
        RECT 21.435 47.440 22.055 47.800 ;
        RECT 21.135 47.060 21.425 47.250 ;
        RECT 19.325 46.620 21.425 47.060 ;
        RECT 19.325 46.600 20.015 46.620 ;
        RECT 21.135 46.380 21.425 46.620 ;
        RECT 22.055 46.990 22.325 47.240 ;
        RECT 22.535 46.990 22.765 48.360 ;
        RECT 25.355 47.010 25.685 52.030 ;
        RECT 26.405 52.020 27.535 53.240 ;
        RECT 28.895 53.220 29.215 53.240 ;
        RECT 22.055 46.880 22.765 46.990 ;
        RECT 25.345 46.960 25.685 47.010 ;
        RECT 26.235 47.780 27.615 52.020 ;
        RECT 22.055 46.570 22.715 46.880 ;
        RECT 22.055 46.400 22.325 46.570 ;
        RECT 25.345 45.000 25.625 46.960 ;
        RECT 26.235 46.920 26.535 47.780 ;
        RECT 27.315 46.920 27.615 47.780 ;
        RECT 28.165 46.920 28.495 51.990 ;
        RECT 27.565 46.380 28.045 46.760 ;
        RECT 27.665 45.760 27.915 46.380 ;
        RECT 27.565 45.160 27.945 45.760 ;
        RECT 24.825 44.230 25.925 45.000 ;
        RECT 28.215 44.930 28.495 46.920 ;
        RECT 30.525 47.780 31.025 68.580 ;
        RECT 31.365 49.100 31.755 70.610 ;
        RECT 32.155 70.020 33.045 70.750 ;
        RECT 32.255 65.200 32.515 70.020 ;
        RECT 33.895 68.630 36.605 69.480 ;
        RECT 34.095 65.850 36.025 68.630 ;
        RECT 41.725 68.550 42.265 71.780 ;
        RECT 42.565 70.580 42.975 73.220 ;
        RECT 50.055 73.090 52.125 74.370 ;
        RECT 53.150 73.290 55.710 75.820 ;
        RECT 64.900 75.810 65.180 77.710 ;
        RECT 103.990 77.230 104.270 84.740 ;
        RECT 76.140 76.950 104.270 77.230 ;
        RECT 52.675 71.760 53.535 72.600 ;
        RECT 38.995 67.140 40.115 67.820 ;
        RECT 39.275 65.860 39.945 67.140 ;
        RECT 32.655 65.470 37.705 65.850 ;
        RECT 39.065 65.450 40.115 65.860 ;
        RECT 32.255 63.650 32.635 65.200 ;
        RECT 32.375 55.810 32.635 63.650 ;
        RECT 37.685 63.210 37.955 65.250 ;
        RECT 38.815 63.210 39.085 65.210 ;
        RECT 37.685 56.520 39.085 63.210 ;
        RECT 32.285 55.300 32.645 55.810 ;
        RECT 32.265 54.870 32.645 55.300 ;
        RECT 37.685 55.200 37.955 56.520 ;
        RECT 38.815 55.160 39.085 56.520 ;
        RECT 40.085 55.270 40.405 65.200 ;
        RECT 40.085 55.210 40.415 55.270 ;
        RECT 32.265 54.590 32.515 54.870 ;
        RECT 32.065 54.190 36.705 54.590 ;
        RECT 37.605 54.300 38.735 54.310 ;
        RECT 40.095 54.300 40.415 55.210 ;
        RECT 32.265 52.070 32.515 54.190 ;
        RECT 36.965 53.500 37.325 54.120 ;
        RECT 37.045 52.620 37.305 53.500 ;
        RECT 37.585 53.250 40.415 54.300 ;
        RECT 36.875 52.240 37.405 52.620 ;
        RECT 32.265 51.980 32.765 52.070 ;
        RECT 32.255 51.250 32.765 51.980 ;
        RECT 32.495 50.250 32.765 51.250 ;
        RECT 33.405 51.000 33.675 51.950 ;
        RECT 33.405 50.850 33.875 51.000 ;
        RECT 33.405 50.170 33.965 50.850 ;
        RECT 33.485 50.160 33.965 50.170 ;
        RECT 32.775 49.630 33.395 49.990 ;
        RECT 32.815 49.100 33.245 49.630 ;
        RECT 31.365 48.680 33.245 49.100 ;
        RECT 33.735 48.970 33.965 50.160 ;
        RECT 32.815 47.810 33.245 48.680 ;
        RECT 33.655 48.370 34.035 48.970 ;
        RECT 30.525 47.070 31.215 47.780 ;
        RECT 32.635 47.450 33.255 47.810 ;
        RECT 32.335 47.070 32.625 47.260 ;
        RECT 30.525 46.630 32.625 47.070 ;
        RECT 30.525 46.610 31.215 46.630 ;
        RECT 32.335 46.390 32.625 46.630 ;
        RECT 33.255 47.000 33.525 47.250 ;
        RECT 33.735 47.000 33.965 48.370 ;
        RECT 36.555 47.020 36.885 52.040 ;
        RECT 37.605 52.030 38.735 53.250 ;
        RECT 40.095 53.230 40.415 53.250 ;
        RECT 33.255 46.890 33.965 47.000 ;
        RECT 36.545 46.970 36.885 47.020 ;
        RECT 37.435 47.790 38.815 52.030 ;
        RECT 33.255 46.580 33.915 46.890 ;
        RECT 33.255 46.410 33.525 46.580 ;
        RECT 36.545 45.010 36.825 46.970 ;
        RECT 37.435 46.930 37.735 47.790 ;
        RECT 38.515 46.930 38.815 47.790 ;
        RECT 39.365 46.930 39.695 52.000 ;
        RECT 38.765 46.390 39.245 46.770 ;
        RECT 38.865 45.770 39.115 46.390 ;
        RECT 38.765 45.170 39.145 45.770 ;
        RECT 28.215 43.200 28.515 44.930 ;
        RECT 36.025 44.240 37.125 45.010 ;
        RECT 39.415 44.940 39.695 46.930 ;
        RECT 41.745 47.750 42.245 68.550 ;
        RECT 42.585 49.070 42.975 70.580 ;
        RECT 43.375 69.990 44.265 70.720 ;
        RECT 43.475 65.170 43.735 69.990 ;
        RECT 45.115 68.600 47.825 69.450 ;
        RECT 45.315 65.820 47.245 68.600 ;
        RECT 52.975 68.530 53.515 71.760 ;
        RECT 53.815 70.560 54.225 73.290 ;
        RECT 61.475 73.120 63.545 74.400 ;
        RECT 64.400 73.280 66.960 75.810 ;
        RECT 76.140 75.740 76.420 76.950 ;
        RECT 109.970 76.610 110.250 85.420 ;
        RECT 87.580 76.330 110.250 76.610 ;
        RECT 87.580 75.760 87.860 76.330 ;
        RECT 115.950 76.030 116.230 85.700 ;
        RECT 98.850 75.840 116.230 76.030 ;
        RECT 63.895 71.750 64.755 72.590 ;
        RECT 50.215 67.110 51.335 67.790 ;
        RECT 50.495 65.830 51.165 67.110 ;
        RECT 43.875 65.440 48.925 65.820 ;
        RECT 50.285 65.420 51.335 65.830 ;
        RECT 43.475 63.620 43.855 65.170 ;
        RECT 43.595 55.780 43.855 63.620 ;
        RECT 48.905 63.180 49.175 65.220 ;
        RECT 50.035 63.180 50.305 65.180 ;
        RECT 48.905 56.490 50.305 63.180 ;
        RECT 43.505 55.270 43.865 55.780 ;
        RECT 43.485 54.840 43.865 55.270 ;
        RECT 48.905 55.170 49.175 56.490 ;
        RECT 50.035 55.130 50.305 56.490 ;
        RECT 51.305 55.240 51.625 65.170 ;
        RECT 51.305 55.180 51.635 55.240 ;
        RECT 43.485 54.560 43.735 54.840 ;
        RECT 43.285 54.160 47.925 54.560 ;
        RECT 48.825 54.270 49.955 54.280 ;
        RECT 51.315 54.270 51.635 55.180 ;
        RECT 43.485 52.040 43.735 54.160 ;
        RECT 48.185 53.470 48.545 54.090 ;
        RECT 48.265 52.590 48.525 53.470 ;
        RECT 48.805 53.220 51.635 54.270 ;
        RECT 48.095 52.210 48.625 52.590 ;
        RECT 43.485 51.950 43.985 52.040 ;
        RECT 43.475 51.220 43.985 51.950 ;
        RECT 43.715 50.220 43.985 51.220 ;
        RECT 44.625 50.970 44.895 51.920 ;
        RECT 44.625 50.820 45.095 50.970 ;
        RECT 44.625 50.140 45.185 50.820 ;
        RECT 44.705 50.130 45.185 50.140 ;
        RECT 43.995 49.600 44.615 49.960 ;
        RECT 44.035 49.070 44.465 49.600 ;
        RECT 42.585 48.650 44.465 49.070 ;
        RECT 44.955 48.940 45.185 50.130 ;
        RECT 44.035 47.780 44.465 48.650 ;
        RECT 44.875 48.340 45.255 48.940 ;
        RECT 41.745 47.040 42.435 47.750 ;
        RECT 43.855 47.420 44.475 47.780 ;
        RECT 43.555 47.040 43.845 47.230 ;
        RECT 41.745 46.600 43.845 47.040 ;
        RECT 41.745 46.580 42.435 46.600 ;
        RECT 43.555 46.360 43.845 46.600 ;
        RECT 44.475 46.970 44.745 47.220 ;
        RECT 44.955 46.970 45.185 48.340 ;
        RECT 47.775 46.990 48.105 52.010 ;
        RECT 48.825 52.000 49.955 53.220 ;
        RECT 51.315 53.200 51.635 53.220 ;
        RECT 44.475 46.860 45.185 46.970 ;
        RECT 47.765 46.940 48.105 46.990 ;
        RECT 48.655 47.760 50.035 52.000 ;
        RECT 44.475 46.550 45.135 46.860 ;
        RECT 44.475 46.380 44.745 46.550 ;
        RECT 47.765 44.980 48.045 46.940 ;
        RECT 48.655 46.900 48.955 47.760 ;
        RECT 49.735 46.900 50.035 47.760 ;
        RECT 50.585 46.900 50.915 51.970 ;
        RECT 49.985 46.360 50.465 46.740 ;
        RECT 50.085 45.740 50.335 46.360 ;
        RECT 49.985 45.140 50.365 45.740 ;
        RECT 39.415 43.210 39.715 44.940 ;
        RECT 47.245 44.210 48.345 44.980 ;
        RECT 50.635 44.910 50.915 46.900 ;
        RECT 52.995 47.730 53.495 68.530 ;
        RECT 53.835 49.050 54.225 70.560 ;
        RECT 54.625 69.970 55.515 70.700 ;
        RECT 54.725 65.150 54.985 69.970 ;
        RECT 56.365 68.580 59.075 69.430 ;
        RECT 56.565 65.800 58.495 68.580 ;
        RECT 64.195 68.520 64.735 71.750 ;
        RECT 65.035 70.550 65.445 73.280 ;
        RECT 72.585 73.130 74.655 74.410 ;
        RECT 75.550 73.210 78.110 75.740 ;
        RECT 75.135 71.740 75.995 72.580 ;
        RECT 61.465 67.090 62.585 67.770 ;
        RECT 61.745 65.810 62.415 67.090 ;
        RECT 55.125 65.420 60.175 65.800 ;
        RECT 61.535 65.400 62.585 65.810 ;
        RECT 54.725 63.600 55.105 65.150 ;
        RECT 54.845 55.760 55.105 63.600 ;
        RECT 60.155 63.160 60.425 65.200 ;
        RECT 61.285 63.160 61.555 65.160 ;
        RECT 60.155 56.470 61.555 63.160 ;
        RECT 54.755 55.250 55.115 55.760 ;
        RECT 54.735 54.820 55.115 55.250 ;
        RECT 60.155 55.150 60.425 56.470 ;
        RECT 61.285 55.110 61.555 56.470 ;
        RECT 62.555 55.220 62.875 65.150 ;
        RECT 62.555 55.160 62.885 55.220 ;
        RECT 54.735 54.540 54.985 54.820 ;
        RECT 54.535 54.140 59.175 54.540 ;
        RECT 60.075 54.250 61.205 54.260 ;
        RECT 62.565 54.250 62.885 55.160 ;
        RECT 54.735 52.020 54.985 54.140 ;
        RECT 59.435 53.450 59.795 54.070 ;
        RECT 59.515 52.570 59.775 53.450 ;
        RECT 60.055 53.200 62.885 54.250 ;
        RECT 59.345 52.190 59.875 52.570 ;
        RECT 54.735 51.930 55.235 52.020 ;
        RECT 54.725 51.200 55.235 51.930 ;
        RECT 54.965 50.200 55.235 51.200 ;
        RECT 55.875 50.950 56.145 51.900 ;
        RECT 55.875 50.800 56.345 50.950 ;
        RECT 55.875 50.120 56.435 50.800 ;
        RECT 55.955 50.110 56.435 50.120 ;
        RECT 55.245 49.580 55.865 49.940 ;
        RECT 55.285 49.050 55.715 49.580 ;
        RECT 53.835 48.630 55.715 49.050 ;
        RECT 56.205 48.920 56.435 50.110 ;
        RECT 55.285 47.760 55.715 48.630 ;
        RECT 56.125 48.320 56.505 48.920 ;
        RECT 52.995 47.020 53.685 47.730 ;
        RECT 55.105 47.400 55.725 47.760 ;
        RECT 54.805 47.020 55.095 47.210 ;
        RECT 52.995 46.580 55.095 47.020 ;
        RECT 52.995 46.560 53.685 46.580 ;
        RECT 54.805 46.340 55.095 46.580 ;
        RECT 55.725 46.950 55.995 47.200 ;
        RECT 56.205 46.950 56.435 48.320 ;
        RECT 59.025 46.970 59.355 51.990 ;
        RECT 60.075 51.980 61.205 53.200 ;
        RECT 62.565 53.180 62.885 53.200 ;
        RECT 55.725 46.840 56.435 46.950 ;
        RECT 59.015 46.920 59.355 46.970 ;
        RECT 59.905 47.740 61.285 51.980 ;
        RECT 55.725 46.530 56.385 46.840 ;
        RECT 55.725 46.360 55.995 46.530 ;
        RECT 59.015 44.960 59.295 46.920 ;
        RECT 59.905 46.880 60.205 47.740 ;
        RECT 60.985 46.880 61.285 47.740 ;
        RECT 61.835 46.880 62.165 51.950 ;
        RECT 61.235 46.340 61.715 46.720 ;
        RECT 61.335 45.720 61.585 46.340 ;
        RECT 61.235 45.120 61.615 45.720 ;
        RECT 19.865 42.210 21.245 42.780 ;
        RECT 27.495 42.630 28.875 43.200 ;
        RECT 31.145 42.210 32.525 42.780 ;
        RECT 38.695 42.640 40.075 43.210 ;
        RECT 50.635 43.180 50.935 44.910 ;
        RECT 58.495 44.190 59.595 44.960 ;
        RECT 61.885 44.890 62.165 46.880 ;
        RECT 64.215 47.720 64.715 68.520 ;
        RECT 65.055 49.040 65.445 70.550 ;
        RECT 65.845 69.960 66.735 70.690 ;
        RECT 65.945 65.140 66.205 69.960 ;
        RECT 67.585 68.570 70.295 69.420 ;
        RECT 67.785 65.790 69.715 68.570 ;
        RECT 75.435 68.510 75.975 71.740 ;
        RECT 76.275 70.540 76.685 73.210 ;
        RECT 83.855 73.120 85.925 74.400 ;
        RECT 86.850 73.230 89.410 75.760 ;
        RECT 98.150 75.750 116.230 75.840 ;
        RECT 86.385 71.750 87.245 72.590 ;
        RECT 72.685 67.080 73.805 67.760 ;
        RECT 72.965 65.800 73.635 67.080 ;
        RECT 66.345 65.410 71.395 65.790 ;
        RECT 72.755 65.390 73.805 65.800 ;
        RECT 65.945 63.590 66.325 65.140 ;
        RECT 66.065 55.750 66.325 63.590 ;
        RECT 71.375 63.150 71.645 65.190 ;
        RECT 72.505 63.150 72.775 65.150 ;
        RECT 71.375 56.460 72.775 63.150 ;
        RECT 65.975 55.240 66.335 55.750 ;
        RECT 65.955 54.810 66.335 55.240 ;
        RECT 71.375 55.140 71.645 56.460 ;
        RECT 72.505 55.100 72.775 56.460 ;
        RECT 73.775 55.210 74.095 65.140 ;
        RECT 73.775 55.150 74.105 55.210 ;
        RECT 65.955 54.530 66.205 54.810 ;
        RECT 65.755 54.130 70.395 54.530 ;
        RECT 71.295 54.240 72.425 54.250 ;
        RECT 73.785 54.240 74.105 55.150 ;
        RECT 65.955 52.010 66.205 54.130 ;
        RECT 70.655 53.440 71.015 54.060 ;
        RECT 70.735 52.560 70.995 53.440 ;
        RECT 71.275 53.190 74.105 54.240 ;
        RECT 70.565 52.180 71.095 52.560 ;
        RECT 65.955 51.920 66.455 52.010 ;
        RECT 65.945 51.190 66.455 51.920 ;
        RECT 66.185 50.190 66.455 51.190 ;
        RECT 67.095 50.940 67.365 51.890 ;
        RECT 67.095 50.790 67.565 50.940 ;
        RECT 67.095 50.110 67.655 50.790 ;
        RECT 67.175 50.100 67.655 50.110 ;
        RECT 66.465 49.570 67.085 49.930 ;
        RECT 66.505 49.040 66.935 49.570 ;
        RECT 65.055 48.620 66.935 49.040 ;
        RECT 67.425 48.910 67.655 50.100 ;
        RECT 66.505 47.750 66.935 48.620 ;
        RECT 67.345 48.310 67.725 48.910 ;
        RECT 64.215 47.010 64.905 47.720 ;
        RECT 66.325 47.390 66.945 47.750 ;
        RECT 66.025 47.010 66.315 47.200 ;
        RECT 64.215 46.570 66.315 47.010 ;
        RECT 64.215 46.550 64.905 46.570 ;
        RECT 66.025 46.330 66.315 46.570 ;
        RECT 66.945 46.940 67.215 47.190 ;
        RECT 67.425 46.940 67.655 48.310 ;
        RECT 70.245 46.960 70.575 51.980 ;
        RECT 71.295 51.970 72.425 53.190 ;
        RECT 73.785 53.170 74.105 53.190 ;
        RECT 66.945 46.830 67.655 46.940 ;
        RECT 70.235 46.910 70.575 46.960 ;
        RECT 71.125 47.730 72.505 51.970 ;
        RECT 66.945 46.520 67.605 46.830 ;
        RECT 66.945 46.350 67.215 46.520 ;
        RECT 70.235 44.950 70.515 46.910 ;
        RECT 71.125 46.870 71.425 47.730 ;
        RECT 72.205 46.870 72.505 47.730 ;
        RECT 73.055 46.870 73.385 51.940 ;
        RECT 72.455 46.330 72.935 46.710 ;
        RECT 72.555 45.710 72.805 46.330 ;
        RECT 72.455 45.110 72.835 45.710 ;
        RECT 20.225 40.480 20.525 42.210 ;
        RECT 20.245 38.490 20.525 40.480 ;
        RECT 22.815 40.410 23.915 41.180 ;
        RECT 31.505 40.480 31.805 42.210 ;
        RECT 42.435 42.190 43.815 42.760 ;
        RECT 49.915 42.610 51.295 43.180 ;
        RECT 61.885 43.160 62.185 44.890 ;
        RECT 69.715 44.180 70.815 44.950 ;
        RECT 73.105 44.880 73.385 46.870 ;
        RECT 75.455 47.710 75.955 68.510 ;
        RECT 76.295 49.030 76.685 70.540 ;
        RECT 77.085 69.950 77.975 70.680 ;
        RECT 77.185 65.130 77.445 69.950 ;
        RECT 78.825 68.560 81.535 69.410 ;
        RECT 79.025 65.780 80.955 68.560 ;
        RECT 86.685 68.520 87.225 71.750 ;
        RECT 87.525 70.550 87.935 73.230 ;
        RECT 95.045 73.060 97.115 74.340 ;
        RECT 98.150 73.310 100.710 75.750 ;
        RECT 109.390 75.480 111.950 75.560 ;
        RECT 121.930 75.480 122.210 85.700 ;
        RECT 127.550 85.510 128.770 89.380 ;
        RECT 127.910 76.040 128.190 85.510 ;
        RECT 133.380 76.580 136.010 77.880 ;
        RECT 137.240 76.560 139.870 77.860 ;
        RECT 109.390 75.200 122.210 75.480 ;
        RECT 97.665 71.740 98.525 72.580 ;
        RECT 83.925 67.070 85.045 67.750 ;
        RECT 84.205 65.790 84.875 67.070 ;
        RECT 77.585 65.400 82.635 65.780 ;
        RECT 83.995 65.380 85.045 65.790 ;
        RECT 77.185 63.580 77.565 65.130 ;
        RECT 77.305 55.740 77.565 63.580 ;
        RECT 82.615 63.140 82.885 65.180 ;
        RECT 83.745 63.140 84.015 65.140 ;
        RECT 82.615 56.450 84.015 63.140 ;
        RECT 77.215 55.230 77.575 55.740 ;
        RECT 77.195 54.800 77.575 55.230 ;
        RECT 82.615 55.130 82.885 56.450 ;
        RECT 83.745 55.090 84.015 56.450 ;
        RECT 85.015 55.200 85.335 65.130 ;
        RECT 85.015 55.140 85.345 55.200 ;
        RECT 77.195 54.520 77.445 54.800 ;
        RECT 76.995 54.120 81.635 54.520 ;
        RECT 82.535 54.230 83.665 54.240 ;
        RECT 85.025 54.230 85.345 55.140 ;
        RECT 77.195 52.000 77.445 54.120 ;
        RECT 81.895 53.430 82.255 54.050 ;
        RECT 81.975 52.550 82.235 53.430 ;
        RECT 82.515 53.180 85.345 54.230 ;
        RECT 81.805 52.170 82.335 52.550 ;
        RECT 77.195 51.910 77.695 52.000 ;
        RECT 77.185 51.180 77.695 51.910 ;
        RECT 77.425 50.180 77.695 51.180 ;
        RECT 78.335 50.930 78.605 51.880 ;
        RECT 78.335 50.780 78.805 50.930 ;
        RECT 78.335 50.100 78.895 50.780 ;
        RECT 78.415 50.090 78.895 50.100 ;
        RECT 77.705 49.560 78.325 49.920 ;
        RECT 77.745 49.030 78.175 49.560 ;
        RECT 76.295 48.610 78.175 49.030 ;
        RECT 78.665 48.900 78.895 50.090 ;
        RECT 77.745 47.740 78.175 48.610 ;
        RECT 78.585 48.300 78.965 48.900 ;
        RECT 75.455 47.000 76.145 47.710 ;
        RECT 77.565 47.380 78.185 47.740 ;
        RECT 77.265 47.000 77.555 47.190 ;
        RECT 75.455 46.560 77.555 47.000 ;
        RECT 75.455 46.540 76.145 46.560 ;
        RECT 77.265 46.320 77.555 46.560 ;
        RECT 78.185 46.930 78.455 47.180 ;
        RECT 78.665 46.930 78.895 48.300 ;
        RECT 81.485 46.950 81.815 51.970 ;
        RECT 82.535 51.960 83.665 53.180 ;
        RECT 85.025 53.160 85.345 53.180 ;
        RECT 78.185 46.820 78.895 46.930 ;
        RECT 81.475 46.900 81.815 46.950 ;
        RECT 82.365 47.720 83.745 51.960 ;
        RECT 78.185 46.510 78.845 46.820 ;
        RECT 78.185 46.340 78.455 46.510 ;
        RECT 81.475 44.940 81.755 46.900 ;
        RECT 82.365 46.860 82.665 47.720 ;
        RECT 83.445 46.860 83.745 47.720 ;
        RECT 84.295 46.860 84.625 51.930 ;
        RECT 83.695 46.320 84.175 46.700 ;
        RECT 83.795 45.700 84.045 46.320 ;
        RECT 83.695 45.100 84.075 45.700 ;
        RECT 53.655 42.190 55.035 42.760 ;
        RECT 61.165 42.590 62.545 43.160 ;
        RECT 73.105 43.150 73.405 44.880 ;
        RECT 80.955 44.170 82.055 44.940 ;
        RECT 84.345 44.870 84.625 46.860 ;
        RECT 86.705 47.720 87.205 68.520 ;
        RECT 87.545 49.040 87.935 70.550 ;
        RECT 88.335 69.960 89.225 70.690 ;
        RECT 88.435 65.140 88.695 69.960 ;
        RECT 90.075 68.570 92.785 69.420 ;
        RECT 90.275 65.790 92.205 68.570 ;
        RECT 97.965 68.510 98.505 71.740 ;
        RECT 98.805 70.540 99.215 73.310 ;
        RECT 106.455 73.110 108.525 74.390 ;
        RECT 109.390 73.030 111.950 75.200 ;
        RECT 125.760 74.810 128.190 76.040 ;
        RECT 121.290 74.790 128.190 74.810 ;
        RECT 120.600 74.530 128.190 74.790 ;
        RECT 117.655 73.110 119.725 74.390 ;
        RECT 120.600 73.180 128.160 74.530 ;
        RECT 129.505 73.190 131.575 74.470 ;
        RECT 120.600 73.110 126.160 73.180 ;
        RECT 108.935 71.740 109.795 72.580 ;
        RECT 95.175 67.080 96.295 67.760 ;
        RECT 95.455 65.800 96.125 67.080 ;
        RECT 88.835 65.410 93.885 65.790 ;
        RECT 95.245 65.390 96.295 65.800 ;
        RECT 88.435 63.590 88.815 65.140 ;
        RECT 88.555 55.750 88.815 63.590 ;
        RECT 93.865 63.150 94.135 65.190 ;
        RECT 94.995 63.150 95.265 65.150 ;
        RECT 93.865 56.460 95.265 63.150 ;
        RECT 88.465 55.240 88.825 55.750 ;
        RECT 88.445 54.810 88.825 55.240 ;
        RECT 93.865 55.140 94.135 56.460 ;
        RECT 94.995 55.100 95.265 56.460 ;
        RECT 96.265 55.210 96.585 65.140 ;
        RECT 96.265 55.150 96.595 55.210 ;
        RECT 88.445 54.530 88.695 54.810 ;
        RECT 88.245 54.130 92.885 54.530 ;
        RECT 93.785 54.240 94.915 54.250 ;
        RECT 96.275 54.240 96.595 55.150 ;
        RECT 88.445 52.010 88.695 54.130 ;
        RECT 93.145 53.440 93.505 54.060 ;
        RECT 93.225 52.560 93.485 53.440 ;
        RECT 93.765 53.190 96.595 54.240 ;
        RECT 93.055 52.180 93.585 52.560 ;
        RECT 88.445 51.920 88.945 52.010 ;
        RECT 88.435 51.190 88.945 51.920 ;
        RECT 88.675 50.190 88.945 51.190 ;
        RECT 89.585 50.940 89.855 51.890 ;
        RECT 89.585 50.790 90.055 50.940 ;
        RECT 89.585 50.110 90.145 50.790 ;
        RECT 89.665 50.100 90.145 50.110 ;
        RECT 88.955 49.570 89.575 49.930 ;
        RECT 88.995 49.040 89.425 49.570 ;
        RECT 87.545 48.620 89.425 49.040 ;
        RECT 89.915 48.910 90.145 50.100 ;
        RECT 88.995 47.750 89.425 48.620 ;
        RECT 89.835 48.310 90.215 48.910 ;
        RECT 86.705 47.010 87.395 47.720 ;
        RECT 88.815 47.390 89.435 47.750 ;
        RECT 88.515 47.010 88.805 47.200 ;
        RECT 86.705 46.570 88.805 47.010 ;
        RECT 86.705 46.550 87.395 46.570 ;
        RECT 88.515 46.330 88.805 46.570 ;
        RECT 89.435 46.940 89.705 47.190 ;
        RECT 89.915 46.940 90.145 48.310 ;
        RECT 92.735 46.960 93.065 51.980 ;
        RECT 93.785 51.970 94.915 53.190 ;
        RECT 96.275 53.170 96.595 53.190 ;
        RECT 89.435 46.830 90.145 46.940 ;
        RECT 92.725 46.910 93.065 46.960 ;
        RECT 93.615 47.730 94.995 51.970 ;
        RECT 89.435 46.520 90.095 46.830 ;
        RECT 89.435 46.350 89.705 46.520 ;
        RECT 92.725 44.950 93.005 46.910 ;
        RECT 93.615 46.870 93.915 47.730 ;
        RECT 94.695 46.870 94.995 47.730 ;
        RECT 95.545 46.870 95.875 51.940 ;
        RECT 94.945 46.330 95.425 46.710 ;
        RECT 95.045 45.710 95.295 46.330 ;
        RECT 94.945 45.110 95.325 45.710 ;
        RECT 64.855 42.190 66.235 42.760 ;
        RECT 72.385 42.580 73.765 43.150 ;
        RECT 84.345 43.140 84.645 44.870 ;
        RECT 92.205 44.180 93.305 44.950 ;
        RECT 95.595 44.880 95.875 46.870 ;
        RECT 97.985 47.710 98.485 68.510 ;
        RECT 98.825 49.030 99.215 70.540 ;
        RECT 99.615 69.950 100.505 70.680 ;
        RECT 99.715 65.130 99.975 69.950 ;
        RECT 101.355 68.560 104.065 69.410 ;
        RECT 101.555 65.780 103.485 68.560 ;
        RECT 109.235 68.510 109.775 71.740 ;
        RECT 110.075 70.540 110.485 73.030 ;
        RECT 120.185 71.740 121.045 72.580 ;
        RECT 106.455 67.070 107.575 67.750 ;
        RECT 106.735 65.790 107.405 67.070 ;
        RECT 100.115 65.400 105.165 65.780 ;
        RECT 106.525 65.380 107.575 65.790 ;
        RECT 99.715 63.580 100.095 65.130 ;
        RECT 99.835 55.740 100.095 63.580 ;
        RECT 105.145 63.140 105.415 65.180 ;
        RECT 106.275 63.140 106.545 65.140 ;
        RECT 105.145 56.450 106.545 63.140 ;
        RECT 99.745 55.230 100.105 55.740 ;
        RECT 99.725 54.800 100.105 55.230 ;
        RECT 105.145 55.130 105.415 56.450 ;
        RECT 106.275 55.090 106.545 56.450 ;
        RECT 107.545 55.200 107.865 65.130 ;
        RECT 107.545 55.140 107.875 55.200 ;
        RECT 99.725 54.520 99.975 54.800 ;
        RECT 99.525 54.120 104.165 54.520 ;
        RECT 105.065 54.230 106.195 54.240 ;
        RECT 107.555 54.230 107.875 55.140 ;
        RECT 99.725 52.000 99.975 54.120 ;
        RECT 104.425 53.430 104.785 54.050 ;
        RECT 104.505 52.550 104.765 53.430 ;
        RECT 105.045 53.180 107.875 54.230 ;
        RECT 104.335 52.170 104.865 52.550 ;
        RECT 99.725 51.910 100.225 52.000 ;
        RECT 99.715 51.180 100.225 51.910 ;
        RECT 99.955 50.180 100.225 51.180 ;
        RECT 100.865 50.930 101.135 51.880 ;
        RECT 100.865 50.780 101.335 50.930 ;
        RECT 100.865 50.100 101.425 50.780 ;
        RECT 100.945 50.090 101.425 50.100 ;
        RECT 100.235 49.560 100.855 49.920 ;
        RECT 100.275 49.030 100.705 49.560 ;
        RECT 98.825 48.610 100.705 49.030 ;
        RECT 101.195 48.900 101.425 50.090 ;
        RECT 100.275 47.740 100.705 48.610 ;
        RECT 101.115 48.300 101.495 48.900 ;
        RECT 97.985 47.000 98.675 47.710 ;
        RECT 100.095 47.380 100.715 47.740 ;
        RECT 99.795 47.000 100.085 47.190 ;
        RECT 97.985 46.560 100.085 47.000 ;
        RECT 97.985 46.540 98.675 46.560 ;
        RECT 99.795 46.320 100.085 46.560 ;
        RECT 100.715 46.930 100.985 47.180 ;
        RECT 101.195 46.930 101.425 48.300 ;
        RECT 104.015 46.950 104.345 51.970 ;
        RECT 105.065 51.960 106.195 53.180 ;
        RECT 107.555 53.160 107.875 53.180 ;
        RECT 100.715 46.820 101.425 46.930 ;
        RECT 104.005 46.900 104.345 46.950 ;
        RECT 104.895 47.720 106.275 51.960 ;
        RECT 100.715 46.510 101.375 46.820 ;
        RECT 100.715 46.340 100.985 46.510 ;
        RECT 104.005 44.940 104.285 46.900 ;
        RECT 104.895 46.860 105.195 47.720 ;
        RECT 105.975 46.860 106.275 47.720 ;
        RECT 106.825 46.860 107.155 51.930 ;
        RECT 106.225 46.320 106.705 46.700 ;
        RECT 106.325 45.700 106.575 46.320 ;
        RECT 106.225 45.100 106.605 45.700 ;
        RECT 95.595 43.150 95.895 44.880 ;
        RECT 103.485 44.170 104.585 44.940 ;
        RECT 106.875 44.870 107.155 46.860 ;
        RECT 109.255 47.710 109.755 68.510 ;
        RECT 110.095 49.030 110.485 70.540 ;
        RECT 110.885 69.950 111.775 70.680 ;
        RECT 110.985 65.130 111.245 69.950 ;
        RECT 112.625 68.560 115.335 69.410 ;
        RECT 112.825 65.780 114.755 68.560 ;
        RECT 120.485 68.510 121.025 71.740 ;
        RECT 121.325 70.540 121.735 73.110 ;
        RECT 132.925 70.810 133.225 70.900 ;
        RECT 117.725 67.070 118.845 67.750 ;
        RECT 118.005 65.790 118.675 67.070 ;
        RECT 111.385 65.400 116.435 65.780 ;
        RECT 117.795 65.380 118.845 65.790 ;
        RECT 110.985 63.580 111.365 65.130 ;
        RECT 111.105 55.740 111.365 63.580 ;
        RECT 116.415 63.140 116.685 65.180 ;
        RECT 117.545 63.140 117.815 65.140 ;
        RECT 116.415 56.450 117.815 63.140 ;
        RECT 111.015 55.230 111.375 55.740 ;
        RECT 110.995 54.800 111.375 55.230 ;
        RECT 116.415 55.130 116.685 56.450 ;
        RECT 117.545 55.090 117.815 56.450 ;
        RECT 118.815 55.200 119.135 65.130 ;
        RECT 118.815 55.140 119.145 55.200 ;
        RECT 110.995 54.520 111.245 54.800 ;
        RECT 110.795 54.120 115.435 54.520 ;
        RECT 116.335 54.230 117.465 54.240 ;
        RECT 118.825 54.230 119.145 55.140 ;
        RECT 110.995 52.000 111.245 54.120 ;
        RECT 115.695 53.430 116.055 54.050 ;
        RECT 115.775 52.550 116.035 53.430 ;
        RECT 116.315 53.180 119.145 54.230 ;
        RECT 115.605 52.170 116.135 52.550 ;
        RECT 110.995 51.910 111.495 52.000 ;
        RECT 110.985 51.180 111.495 51.910 ;
        RECT 111.225 50.180 111.495 51.180 ;
        RECT 112.135 50.930 112.405 51.880 ;
        RECT 112.135 50.780 112.605 50.930 ;
        RECT 112.135 50.100 112.695 50.780 ;
        RECT 112.215 50.090 112.695 50.100 ;
        RECT 111.505 49.560 112.125 49.920 ;
        RECT 111.545 49.030 111.975 49.560 ;
        RECT 110.095 48.610 111.975 49.030 ;
        RECT 112.465 48.900 112.695 50.090 ;
        RECT 111.545 47.740 111.975 48.610 ;
        RECT 112.385 48.300 112.765 48.900 ;
        RECT 109.255 47.000 109.945 47.710 ;
        RECT 111.365 47.380 111.985 47.740 ;
        RECT 111.065 47.000 111.355 47.190 ;
        RECT 109.255 46.560 111.355 47.000 ;
        RECT 109.255 46.540 109.945 46.560 ;
        RECT 111.065 46.320 111.355 46.560 ;
        RECT 111.985 46.930 112.255 47.180 ;
        RECT 112.465 46.930 112.695 48.300 ;
        RECT 115.285 46.950 115.615 51.970 ;
        RECT 116.335 51.960 117.465 53.180 ;
        RECT 118.825 53.160 119.145 53.180 ;
        RECT 111.985 46.820 112.695 46.930 ;
        RECT 115.275 46.900 115.615 46.950 ;
        RECT 116.165 47.720 117.545 51.960 ;
        RECT 111.985 46.510 112.645 46.820 ;
        RECT 111.985 46.340 112.255 46.510 ;
        RECT 115.275 44.940 115.555 46.900 ;
        RECT 116.165 46.860 116.465 47.720 ;
        RECT 117.245 46.860 117.545 47.720 ;
        RECT 118.095 46.860 118.425 51.930 ;
        RECT 117.495 46.320 117.975 46.700 ;
        RECT 117.595 45.700 117.845 46.320 ;
        RECT 117.495 45.100 117.875 45.700 ;
        RECT 20.795 39.650 21.175 40.250 ;
        RECT 20.825 39.030 21.075 39.650 ;
        RECT 20.695 38.650 21.175 39.030 ;
        RECT 20.245 33.420 20.575 38.490 ;
        RECT 21.125 37.630 21.425 38.490 ;
        RECT 22.205 37.630 22.505 38.490 ;
        RECT 23.115 38.450 23.395 40.410 ;
        RECT 26.415 38.840 26.685 39.010 ;
        RECT 26.025 38.530 26.685 38.840 ;
        RECT 21.125 33.390 22.505 37.630 ;
        RECT 23.055 38.400 23.395 38.450 ;
        RECT 25.975 38.420 26.685 38.530 ;
        RECT 19.525 32.170 19.845 32.190 ;
        RECT 21.205 32.170 22.335 33.390 ;
        RECT 23.055 33.380 23.385 38.400 ;
        RECT 25.975 37.050 26.205 38.420 ;
        RECT 26.415 38.170 26.685 38.420 ;
        RECT 27.315 38.790 27.605 39.030 ;
        RECT 28.725 38.790 29.415 38.810 ;
        RECT 27.315 38.350 29.415 38.790 ;
        RECT 27.315 38.160 27.605 38.350 ;
        RECT 26.685 37.610 27.305 37.970 ;
        RECT 28.725 37.640 29.415 38.350 ;
        RECT 25.905 36.450 26.285 37.050 ;
        RECT 26.695 36.740 27.125 37.610 ;
        RECT 25.975 35.260 26.205 36.450 ;
        RECT 26.695 36.320 28.575 36.740 ;
        RECT 26.695 35.790 27.125 36.320 ;
        RECT 26.545 35.430 27.165 35.790 ;
        RECT 25.975 35.250 26.455 35.260 ;
        RECT 25.975 34.570 26.535 35.250 ;
        RECT 26.065 34.420 26.535 34.570 ;
        RECT 26.265 33.470 26.535 34.420 ;
        RECT 27.175 34.170 27.445 35.170 ;
        RECT 27.175 33.440 27.685 34.170 ;
        RECT 27.175 33.350 27.675 33.440 ;
        RECT 22.535 32.800 23.065 33.180 ;
        RECT 19.525 31.120 22.355 32.170 ;
        RECT 22.635 31.920 22.895 32.800 ;
        RECT 22.615 31.300 22.975 31.920 ;
        RECT 27.425 31.230 27.675 33.350 ;
        RECT 19.525 30.210 19.845 31.120 ;
        RECT 21.205 31.110 22.335 31.120 ;
        RECT 23.235 30.830 27.875 31.230 ;
        RECT 27.425 30.550 27.675 30.830 ;
        RECT 19.525 30.150 19.855 30.210 ;
        RECT 19.535 20.220 19.855 30.150 ;
        RECT 20.855 28.900 21.125 30.260 ;
        RECT 21.985 28.900 22.255 30.220 ;
        RECT 27.295 30.120 27.675 30.550 ;
        RECT 27.295 29.610 27.655 30.120 ;
        RECT 20.855 22.210 22.255 28.900 ;
        RECT 20.855 20.210 21.125 22.210 ;
        RECT 21.985 20.170 22.255 22.210 ;
        RECT 27.305 21.770 27.565 29.610 ;
        RECT 27.305 20.220 27.685 21.770 ;
        RECT 19.825 19.560 20.875 19.970 ;
        RECT 22.235 19.570 27.285 19.950 ;
        RECT 19.995 18.280 20.665 19.560 ;
        RECT 19.825 17.600 20.945 18.280 ;
        RECT 23.915 16.790 25.845 19.570 ;
        RECT 23.335 15.940 26.045 16.790 ;
        RECT 27.425 15.400 27.685 20.220 ;
        RECT 26.895 14.670 27.785 15.400 ;
        RECT 28.185 14.810 28.575 36.320 ;
        RECT 28.915 16.840 29.415 37.640 ;
        RECT 31.525 38.490 31.805 40.480 ;
        RECT 34.095 40.410 35.195 41.180 ;
        RECT 42.795 40.460 43.095 42.190 ;
        RECT 32.075 39.650 32.455 40.250 ;
        RECT 32.105 39.030 32.355 39.650 ;
        RECT 31.975 38.650 32.455 39.030 ;
        RECT 31.525 33.420 31.855 38.490 ;
        RECT 32.405 37.630 32.705 38.490 ;
        RECT 33.485 37.630 33.785 38.490 ;
        RECT 34.395 38.450 34.675 40.410 ;
        RECT 37.695 38.840 37.965 39.010 ;
        RECT 37.305 38.530 37.965 38.840 ;
        RECT 32.405 33.390 33.785 37.630 ;
        RECT 34.335 38.400 34.675 38.450 ;
        RECT 37.255 38.420 37.965 38.530 ;
        RECT 30.805 32.170 31.125 32.190 ;
        RECT 32.485 32.170 33.615 33.390 ;
        RECT 34.335 33.380 34.665 38.400 ;
        RECT 37.255 37.050 37.485 38.420 ;
        RECT 37.695 38.170 37.965 38.420 ;
        RECT 38.595 38.790 38.885 39.030 ;
        RECT 40.005 38.790 40.695 38.810 ;
        RECT 38.595 38.350 40.695 38.790 ;
        RECT 38.595 38.160 38.885 38.350 ;
        RECT 37.965 37.610 38.585 37.970 ;
        RECT 40.005 37.640 40.695 38.350 ;
        RECT 37.185 36.450 37.565 37.050 ;
        RECT 37.975 36.740 38.405 37.610 ;
        RECT 37.255 35.260 37.485 36.450 ;
        RECT 37.975 36.320 39.855 36.740 ;
        RECT 37.975 35.790 38.405 36.320 ;
        RECT 37.825 35.430 38.445 35.790 ;
        RECT 37.255 35.250 37.735 35.260 ;
        RECT 37.255 34.570 37.815 35.250 ;
        RECT 37.345 34.420 37.815 34.570 ;
        RECT 37.545 33.470 37.815 34.420 ;
        RECT 38.455 34.170 38.725 35.170 ;
        RECT 38.455 33.440 38.965 34.170 ;
        RECT 38.455 33.350 38.955 33.440 ;
        RECT 33.815 32.800 34.345 33.180 ;
        RECT 30.805 31.120 33.635 32.170 ;
        RECT 33.915 31.920 34.175 32.800 ;
        RECT 33.895 31.300 34.255 31.920 ;
        RECT 38.705 31.230 38.955 33.350 ;
        RECT 30.805 30.210 31.125 31.120 ;
        RECT 32.485 31.110 33.615 31.120 ;
        RECT 34.515 30.830 39.155 31.230 ;
        RECT 38.705 30.550 38.955 30.830 ;
        RECT 30.805 30.150 31.135 30.210 ;
        RECT 30.815 20.220 31.135 30.150 ;
        RECT 32.135 28.900 32.405 30.260 ;
        RECT 33.265 28.900 33.535 30.220 ;
        RECT 38.575 30.120 38.955 30.550 ;
        RECT 38.575 29.610 38.935 30.120 ;
        RECT 32.135 22.210 33.535 28.900 ;
        RECT 32.135 20.210 32.405 22.210 ;
        RECT 33.265 20.170 33.535 22.210 ;
        RECT 38.585 21.770 38.845 29.610 ;
        RECT 38.585 20.220 38.965 21.770 ;
        RECT 31.105 19.560 32.155 19.970 ;
        RECT 33.515 19.570 38.565 19.950 ;
        RECT 31.275 18.280 31.945 19.560 ;
        RECT 31.105 17.600 32.225 18.280 ;
        RECT 28.185 12.290 28.595 14.810 ;
        RECT 28.895 13.610 29.435 16.840 ;
        RECT 35.195 16.790 37.125 19.570 ;
        RECT 34.615 15.940 37.325 16.790 ;
        RECT 38.705 15.400 38.965 20.220 ;
        RECT 38.175 14.670 39.065 15.400 ;
        RECT 39.465 14.810 39.855 36.320 ;
        RECT 40.195 16.840 40.695 37.640 ;
        RECT 42.815 38.470 43.095 40.460 ;
        RECT 45.385 40.390 46.485 41.160 ;
        RECT 54.015 40.460 54.315 42.190 ;
        RECT 43.365 39.630 43.745 40.230 ;
        RECT 43.395 39.010 43.645 39.630 ;
        RECT 43.265 38.630 43.745 39.010 ;
        RECT 42.815 33.400 43.145 38.470 ;
        RECT 43.695 37.610 43.995 38.470 ;
        RECT 44.775 37.610 45.075 38.470 ;
        RECT 45.685 38.430 45.965 40.390 ;
        RECT 48.985 38.820 49.255 38.990 ;
        RECT 48.595 38.510 49.255 38.820 ;
        RECT 43.695 33.370 45.075 37.610 ;
        RECT 45.625 38.380 45.965 38.430 ;
        RECT 48.545 38.400 49.255 38.510 ;
        RECT 42.095 32.150 42.415 32.170 ;
        RECT 43.775 32.150 44.905 33.370 ;
        RECT 45.625 33.360 45.955 38.380 ;
        RECT 48.545 37.030 48.775 38.400 ;
        RECT 48.985 38.150 49.255 38.400 ;
        RECT 49.885 38.770 50.175 39.010 ;
        RECT 51.295 38.770 51.985 38.790 ;
        RECT 49.885 38.330 51.985 38.770 ;
        RECT 49.885 38.140 50.175 38.330 ;
        RECT 49.255 37.590 49.875 37.950 ;
        RECT 51.295 37.620 51.985 38.330 ;
        RECT 48.475 36.430 48.855 37.030 ;
        RECT 49.265 36.720 49.695 37.590 ;
        RECT 48.545 35.240 48.775 36.430 ;
        RECT 49.265 36.300 51.145 36.720 ;
        RECT 49.265 35.770 49.695 36.300 ;
        RECT 49.115 35.410 49.735 35.770 ;
        RECT 48.545 35.230 49.025 35.240 ;
        RECT 48.545 34.550 49.105 35.230 ;
        RECT 48.635 34.400 49.105 34.550 ;
        RECT 48.835 33.450 49.105 34.400 ;
        RECT 49.745 34.150 50.015 35.150 ;
        RECT 49.745 33.420 50.255 34.150 ;
        RECT 49.745 33.330 50.245 33.420 ;
        RECT 45.105 32.780 45.635 33.160 ;
        RECT 42.095 31.100 44.925 32.150 ;
        RECT 45.205 31.900 45.465 32.780 ;
        RECT 45.185 31.280 45.545 31.900 ;
        RECT 49.995 31.210 50.245 33.330 ;
        RECT 42.095 30.190 42.415 31.100 ;
        RECT 43.775 31.090 44.905 31.100 ;
        RECT 45.805 30.810 50.445 31.210 ;
        RECT 49.995 30.530 50.245 30.810 ;
        RECT 42.095 30.130 42.425 30.190 ;
        RECT 42.105 20.200 42.425 30.130 ;
        RECT 43.425 28.880 43.695 30.240 ;
        RECT 44.555 28.880 44.825 30.200 ;
        RECT 49.865 30.100 50.245 30.530 ;
        RECT 49.865 29.590 50.225 30.100 ;
        RECT 43.425 22.190 44.825 28.880 ;
        RECT 43.425 20.190 43.695 22.190 ;
        RECT 44.555 20.150 44.825 22.190 ;
        RECT 49.875 21.750 50.135 29.590 ;
        RECT 49.875 20.200 50.255 21.750 ;
        RECT 42.395 19.540 43.445 19.950 ;
        RECT 44.805 19.550 49.855 19.930 ;
        RECT 42.565 18.260 43.235 19.540 ;
        RECT 42.395 17.580 43.515 18.260 ;
        RECT 28.875 12.770 29.735 13.610 ;
        RECT 28.185 11.950 30.415 12.290 ;
        RECT 39.465 11.990 39.875 14.810 ;
        RECT 40.175 13.610 40.715 16.840 ;
        RECT 46.485 16.770 48.415 19.550 ;
        RECT 45.905 15.920 48.615 16.770 ;
        RECT 49.995 15.380 50.255 20.200 ;
        RECT 49.465 14.650 50.355 15.380 ;
        RECT 50.755 14.790 51.145 36.300 ;
        RECT 51.485 16.820 51.985 37.620 ;
        RECT 54.035 38.470 54.315 40.460 ;
        RECT 56.605 40.390 57.705 41.160 ;
        RECT 65.215 40.460 65.515 42.190 ;
        RECT 76.145 42.180 77.525 42.750 ;
        RECT 83.625 42.570 85.005 43.140 ;
        RECT 87.385 42.200 88.765 42.770 ;
        RECT 94.875 42.580 96.255 43.150 ;
        RECT 106.875 43.140 107.175 44.870 ;
        RECT 114.755 44.170 115.855 44.940 ;
        RECT 118.145 44.870 118.425 46.860 ;
        RECT 120.505 47.710 121.005 68.510 ;
        RECT 121.345 49.030 121.735 70.540 ;
        RECT 122.135 69.950 123.025 70.680 ;
        RECT 132.615 70.040 134.265 70.810 ;
        RECT 122.235 65.130 122.495 69.950 ;
        RECT 123.875 68.560 126.585 69.410 ;
        RECT 124.075 65.780 126.005 68.560 ;
        RECT 128.975 67.070 130.095 67.750 ;
        RECT 129.255 65.790 129.925 67.070 ;
        RECT 122.635 65.400 127.685 65.780 ;
        RECT 129.045 65.380 130.095 65.790 ;
        RECT 132.925 65.180 133.225 70.040 ;
        RECT 137.675 68.690 139.075 69.460 ;
        RECT 138.385 65.740 138.645 68.690 ;
        RECT 149.410 68.420 150.690 69.620 ;
        RECT 149.480 65.810 150.640 68.420 ;
        RECT 133.365 65.380 138.645 65.740 ;
        RECT 122.235 63.580 122.615 65.130 ;
        RECT 122.355 55.740 122.615 63.580 ;
        RECT 127.665 63.140 127.935 65.180 ;
        RECT 128.795 63.140 129.065 65.140 ;
        RECT 127.665 56.450 129.065 63.140 ;
        RECT 122.265 55.230 122.625 55.740 ;
        RECT 122.245 54.800 122.625 55.230 ;
        RECT 127.665 55.130 127.935 56.450 ;
        RECT 128.795 55.090 129.065 56.450 ;
        RECT 130.065 55.200 130.385 65.130 ;
        RECT 132.925 61.010 133.355 65.180 ;
        RECT 138.385 65.150 138.645 65.380 ;
        RECT 138.385 64.770 138.675 65.150 ;
        RECT 130.065 55.140 130.395 55.200 ;
        RECT 133.055 55.190 133.355 61.010 ;
        RECT 122.245 54.520 122.495 54.800 ;
        RECT 122.045 54.120 126.685 54.520 ;
        RECT 127.585 54.230 128.715 54.240 ;
        RECT 130.075 54.230 130.395 55.140 ;
        RECT 138.395 55.080 138.675 64.770 ;
        RECT 149.390 64.610 150.670 65.810 ;
        RECT 122.245 52.000 122.495 54.120 ;
        RECT 126.945 53.430 127.305 54.050 ;
        RECT 127.025 52.550 127.285 53.430 ;
        RECT 127.565 53.180 130.395 54.230 ;
        RECT 126.855 52.170 127.385 52.550 ;
        RECT 122.245 51.910 122.745 52.000 ;
        RECT 122.235 51.180 122.745 51.910 ;
        RECT 122.475 50.180 122.745 51.180 ;
        RECT 123.385 50.930 123.655 51.880 ;
        RECT 123.385 50.780 123.855 50.930 ;
        RECT 123.385 50.100 123.945 50.780 ;
        RECT 123.465 50.090 123.945 50.100 ;
        RECT 122.755 49.560 123.375 49.920 ;
        RECT 122.795 49.030 123.225 49.560 ;
        RECT 121.345 48.610 123.225 49.030 ;
        RECT 123.715 48.900 123.945 50.090 ;
        RECT 122.795 47.740 123.225 48.610 ;
        RECT 123.635 48.300 124.015 48.900 ;
        RECT 120.505 47.000 121.195 47.710 ;
        RECT 122.615 47.380 123.235 47.740 ;
        RECT 122.315 47.000 122.605 47.190 ;
        RECT 120.505 46.560 122.605 47.000 ;
        RECT 120.505 46.540 121.195 46.560 ;
        RECT 122.315 46.320 122.605 46.560 ;
        RECT 123.235 46.930 123.505 47.180 ;
        RECT 123.715 46.930 123.945 48.300 ;
        RECT 126.535 46.950 126.865 51.970 ;
        RECT 127.585 51.960 128.715 53.180 ;
        RECT 130.075 53.160 130.395 53.180 ;
        RECT 123.235 46.820 123.945 46.930 ;
        RECT 126.525 46.900 126.865 46.950 ;
        RECT 127.415 47.720 128.795 51.960 ;
        RECT 123.235 46.510 123.895 46.820 ;
        RECT 123.235 46.340 123.505 46.510 ;
        RECT 126.525 44.940 126.805 46.900 ;
        RECT 127.415 46.860 127.715 47.720 ;
        RECT 128.495 46.860 128.795 47.720 ;
        RECT 129.345 46.860 129.675 51.930 ;
        RECT 128.745 46.320 129.225 46.700 ;
        RECT 128.845 45.700 129.095 46.320 ;
        RECT 128.745 45.100 129.125 45.700 ;
        RECT 118.145 43.140 118.445 44.870 ;
        RECT 126.005 44.170 127.105 44.940 ;
        RECT 129.395 44.870 129.675 46.860 ;
        RECT 129.395 43.140 129.695 44.870 ;
        RECT 98.595 42.220 99.975 42.790 ;
        RECT 106.155 42.570 107.535 43.140 ;
        RECT 109.795 42.260 111.175 42.830 ;
        RECT 117.425 42.570 118.805 43.140 ;
        RECT 121.005 42.280 122.385 42.850 ;
        RECT 128.675 42.570 130.055 43.140 ;
        RECT 54.585 39.630 54.965 40.230 ;
        RECT 54.615 39.010 54.865 39.630 ;
        RECT 54.485 38.630 54.965 39.010 ;
        RECT 54.035 33.400 54.365 38.470 ;
        RECT 54.915 37.610 55.215 38.470 ;
        RECT 55.995 37.610 56.295 38.470 ;
        RECT 56.905 38.430 57.185 40.390 ;
        RECT 60.205 38.820 60.475 38.990 ;
        RECT 59.815 38.510 60.475 38.820 ;
        RECT 54.915 33.370 56.295 37.610 ;
        RECT 56.845 38.380 57.185 38.430 ;
        RECT 59.765 38.400 60.475 38.510 ;
        RECT 53.315 32.150 53.635 32.170 ;
        RECT 54.995 32.150 56.125 33.370 ;
        RECT 56.845 33.360 57.175 38.380 ;
        RECT 59.765 37.030 59.995 38.400 ;
        RECT 60.205 38.150 60.475 38.400 ;
        RECT 61.105 38.770 61.395 39.010 ;
        RECT 62.515 38.770 63.205 38.790 ;
        RECT 61.105 38.330 63.205 38.770 ;
        RECT 61.105 38.140 61.395 38.330 ;
        RECT 60.475 37.590 61.095 37.950 ;
        RECT 62.515 37.620 63.205 38.330 ;
        RECT 59.695 36.430 60.075 37.030 ;
        RECT 60.485 36.720 60.915 37.590 ;
        RECT 59.765 35.240 59.995 36.430 ;
        RECT 60.485 36.300 62.365 36.720 ;
        RECT 60.485 35.770 60.915 36.300 ;
        RECT 60.335 35.410 60.955 35.770 ;
        RECT 59.765 35.230 60.245 35.240 ;
        RECT 59.765 34.550 60.325 35.230 ;
        RECT 59.855 34.400 60.325 34.550 ;
        RECT 60.055 33.450 60.325 34.400 ;
        RECT 60.965 34.150 61.235 35.150 ;
        RECT 60.965 33.420 61.475 34.150 ;
        RECT 60.965 33.330 61.465 33.420 ;
        RECT 56.325 32.780 56.855 33.160 ;
        RECT 53.315 31.100 56.145 32.150 ;
        RECT 56.425 31.900 56.685 32.780 ;
        RECT 56.405 31.280 56.765 31.900 ;
        RECT 61.215 31.210 61.465 33.330 ;
        RECT 53.315 30.190 53.635 31.100 ;
        RECT 54.995 31.090 56.125 31.100 ;
        RECT 57.025 30.810 61.665 31.210 ;
        RECT 61.215 30.530 61.465 30.810 ;
        RECT 53.315 30.130 53.645 30.190 ;
        RECT 53.325 20.200 53.645 30.130 ;
        RECT 54.645 28.880 54.915 30.240 ;
        RECT 55.775 28.880 56.045 30.200 ;
        RECT 61.085 30.100 61.465 30.530 ;
        RECT 61.085 29.590 61.445 30.100 ;
        RECT 54.645 22.190 56.045 28.880 ;
        RECT 54.645 20.190 54.915 22.190 ;
        RECT 55.775 20.150 56.045 22.190 ;
        RECT 61.095 21.750 61.355 29.590 ;
        RECT 61.095 20.200 61.475 21.750 ;
        RECT 53.615 19.540 54.665 19.950 ;
        RECT 56.025 19.550 61.075 19.930 ;
        RECT 53.785 18.260 54.455 19.540 ;
        RECT 53.615 17.580 54.735 18.260 ;
        RECT 40.155 12.770 41.015 13.610 ;
        RECT 50.755 12.170 51.165 14.790 ;
        RECT 51.465 13.590 52.005 16.820 ;
        RECT 57.705 16.770 59.635 19.550 ;
        RECT 57.125 15.920 59.835 16.770 ;
        RECT 61.215 15.380 61.475 20.200 ;
        RECT 60.685 14.650 61.575 15.380 ;
        RECT 61.975 14.790 62.365 36.300 ;
        RECT 62.705 16.820 63.205 37.620 ;
        RECT 65.235 38.470 65.515 40.460 ;
        RECT 67.805 40.390 68.905 41.160 ;
        RECT 76.505 40.450 76.805 42.180 ;
        RECT 65.785 39.630 66.165 40.230 ;
        RECT 65.815 39.010 66.065 39.630 ;
        RECT 65.685 38.630 66.165 39.010 ;
        RECT 65.235 33.400 65.565 38.470 ;
        RECT 66.115 37.610 66.415 38.470 ;
        RECT 67.195 37.610 67.495 38.470 ;
        RECT 68.105 38.430 68.385 40.390 ;
        RECT 71.405 38.820 71.675 38.990 ;
        RECT 71.015 38.510 71.675 38.820 ;
        RECT 66.115 33.370 67.495 37.610 ;
        RECT 68.045 38.380 68.385 38.430 ;
        RECT 70.965 38.400 71.675 38.510 ;
        RECT 64.515 32.150 64.835 32.170 ;
        RECT 66.195 32.150 67.325 33.370 ;
        RECT 68.045 33.360 68.375 38.380 ;
        RECT 70.965 37.030 71.195 38.400 ;
        RECT 71.405 38.150 71.675 38.400 ;
        RECT 72.305 38.770 72.595 39.010 ;
        RECT 73.715 38.770 74.405 38.790 ;
        RECT 72.305 38.330 74.405 38.770 ;
        RECT 72.305 38.140 72.595 38.330 ;
        RECT 71.675 37.590 72.295 37.950 ;
        RECT 73.715 37.620 74.405 38.330 ;
        RECT 70.895 36.430 71.275 37.030 ;
        RECT 71.685 36.720 72.115 37.590 ;
        RECT 70.965 35.240 71.195 36.430 ;
        RECT 71.685 36.300 73.565 36.720 ;
        RECT 71.685 35.770 72.115 36.300 ;
        RECT 71.535 35.410 72.155 35.770 ;
        RECT 70.965 35.230 71.445 35.240 ;
        RECT 70.965 34.550 71.525 35.230 ;
        RECT 71.055 34.400 71.525 34.550 ;
        RECT 71.255 33.450 71.525 34.400 ;
        RECT 72.165 34.150 72.435 35.150 ;
        RECT 72.165 33.420 72.675 34.150 ;
        RECT 72.165 33.330 72.665 33.420 ;
        RECT 67.525 32.780 68.055 33.160 ;
        RECT 64.515 31.100 67.345 32.150 ;
        RECT 67.625 31.900 67.885 32.780 ;
        RECT 67.605 31.280 67.965 31.900 ;
        RECT 72.415 31.210 72.665 33.330 ;
        RECT 64.515 30.190 64.835 31.100 ;
        RECT 66.195 31.090 67.325 31.100 ;
        RECT 68.225 30.810 72.865 31.210 ;
        RECT 72.415 30.530 72.665 30.810 ;
        RECT 64.515 30.130 64.845 30.190 ;
        RECT 64.525 20.200 64.845 30.130 ;
        RECT 65.845 28.880 66.115 30.240 ;
        RECT 66.975 28.880 67.245 30.200 ;
        RECT 72.285 30.100 72.665 30.530 ;
        RECT 72.285 29.590 72.645 30.100 ;
        RECT 65.845 22.190 67.245 28.880 ;
        RECT 65.845 20.190 66.115 22.190 ;
        RECT 66.975 20.150 67.245 22.190 ;
        RECT 72.295 21.750 72.555 29.590 ;
        RECT 72.295 20.200 72.675 21.750 ;
        RECT 64.815 19.540 65.865 19.950 ;
        RECT 67.225 19.550 72.275 19.930 ;
        RECT 64.985 18.260 65.655 19.540 ;
        RECT 64.815 17.580 65.935 18.260 ;
        RECT 51.445 12.750 52.305 13.590 ;
        RECT 27.865 11.130 30.415 11.950 ;
        RECT 28.395 11.090 30.415 11.130 ;
        RECT 39.115 10.980 41.565 11.990 ;
        RECT 50.335 10.970 52.355 12.170 ;
        RECT 61.975 12.160 62.385 14.790 ;
        RECT 62.685 13.590 63.225 16.820 ;
        RECT 68.905 16.770 70.835 19.550 ;
        RECT 68.325 15.920 71.035 16.770 ;
        RECT 72.415 15.380 72.675 20.200 ;
        RECT 71.885 14.650 72.775 15.380 ;
        RECT 73.175 14.790 73.565 36.300 ;
        RECT 73.905 16.820 74.405 37.620 ;
        RECT 76.525 38.460 76.805 40.450 ;
        RECT 79.095 40.380 80.195 41.150 ;
        RECT 87.745 40.470 88.045 42.200 ;
        RECT 77.075 39.620 77.455 40.220 ;
        RECT 77.105 39.000 77.355 39.620 ;
        RECT 76.975 38.620 77.455 39.000 ;
        RECT 76.525 33.390 76.855 38.460 ;
        RECT 77.405 37.600 77.705 38.460 ;
        RECT 78.485 37.600 78.785 38.460 ;
        RECT 79.395 38.420 79.675 40.380 ;
        RECT 82.695 38.810 82.965 38.980 ;
        RECT 82.305 38.500 82.965 38.810 ;
        RECT 77.405 33.360 78.785 37.600 ;
        RECT 79.335 38.370 79.675 38.420 ;
        RECT 82.255 38.390 82.965 38.500 ;
        RECT 75.805 32.140 76.125 32.160 ;
        RECT 77.485 32.140 78.615 33.360 ;
        RECT 79.335 33.350 79.665 38.370 ;
        RECT 82.255 37.020 82.485 38.390 ;
        RECT 82.695 38.140 82.965 38.390 ;
        RECT 83.595 38.760 83.885 39.000 ;
        RECT 85.005 38.760 85.695 38.780 ;
        RECT 83.595 38.320 85.695 38.760 ;
        RECT 83.595 38.130 83.885 38.320 ;
        RECT 82.965 37.580 83.585 37.940 ;
        RECT 85.005 37.610 85.695 38.320 ;
        RECT 82.185 36.420 82.565 37.020 ;
        RECT 82.975 36.710 83.405 37.580 ;
        RECT 82.255 35.230 82.485 36.420 ;
        RECT 82.975 36.290 84.855 36.710 ;
        RECT 82.975 35.760 83.405 36.290 ;
        RECT 82.825 35.400 83.445 35.760 ;
        RECT 82.255 35.220 82.735 35.230 ;
        RECT 82.255 34.540 82.815 35.220 ;
        RECT 82.345 34.390 82.815 34.540 ;
        RECT 82.545 33.440 82.815 34.390 ;
        RECT 83.455 34.140 83.725 35.140 ;
        RECT 83.455 33.410 83.965 34.140 ;
        RECT 83.455 33.320 83.955 33.410 ;
        RECT 78.815 32.770 79.345 33.150 ;
        RECT 75.805 31.090 78.635 32.140 ;
        RECT 78.915 31.890 79.175 32.770 ;
        RECT 78.895 31.270 79.255 31.890 ;
        RECT 83.705 31.200 83.955 33.320 ;
        RECT 75.805 30.180 76.125 31.090 ;
        RECT 77.485 31.080 78.615 31.090 ;
        RECT 79.515 30.800 84.155 31.200 ;
        RECT 83.705 30.520 83.955 30.800 ;
        RECT 75.805 30.120 76.135 30.180 ;
        RECT 75.815 20.190 76.135 30.120 ;
        RECT 77.135 28.870 77.405 30.230 ;
        RECT 78.265 28.870 78.535 30.190 ;
        RECT 83.575 30.090 83.955 30.520 ;
        RECT 83.575 29.580 83.935 30.090 ;
        RECT 77.135 22.180 78.535 28.870 ;
        RECT 77.135 20.180 77.405 22.180 ;
        RECT 78.265 20.140 78.535 22.180 ;
        RECT 83.585 21.740 83.845 29.580 ;
        RECT 83.585 20.190 83.965 21.740 ;
        RECT 76.105 19.530 77.155 19.940 ;
        RECT 78.515 19.540 83.565 19.920 ;
        RECT 76.275 18.250 76.945 19.530 ;
        RECT 76.105 17.570 77.225 18.250 ;
        RECT 62.665 12.750 63.525 13.590 ;
        RECT 73.175 12.190 73.585 14.790 ;
        RECT 73.885 13.590 74.425 16.820 ;
        RECT 80.195 16.760 82.125 19.540 ;
        RECT 79.615 15.910 82.325 16.760 ;
        RECT 83.705 15.370 83.965 20.190 ;
        RECT 83.175 14.640 84.065 15.370 ;
        RECT 84.465 14.780 84.855 36.290 ;
        RECT 85.195 16.810 85.695 37.610 ;
        RECT 87.765 38.480 88.045 40.470 ;
        RECT 90.335 40.400 91.435 41.170 ;
        RECT 98.955 40.490 99.255 42.220 ;
        RECT 88.315 39.640 88.695 40.240 ;
        RECT 88.345 39.020 88.595 39.640 ;
        RECT 88.215 38.640 88.695 39.020 ;
        RECT 87.765 33.410 88.095 38.480 ;
        RECT 88.645 37.620 88.945 38.480 ;
        RECT 89.725 37.620 90.025 38.480 ;
        RECT 90.635 38.440 90.915 40.400 ;
        RECT 93.935 38.830 94.205 39.000 ;
        RECT 93.545 38.520 94.205 38.830 ;
        RECT 88.645 33.380 90.025 37.620 ;
        RECT 90.575 38.390 90.915 38.440 ;
        RECT 93.495 38.410 94.205 38.520 ;
        RECT 87.045 32.160 87.365 32.180 ;
        RECT 88.725 32.160 89.855 33.380 ;
        RECT 90.575 33.370 90.905 38.390 ;
        RECT 93.495 37.040 93.725 38.410 ;
        RECT 93.935 38.160 94.205 38.410 ;
        RECT 94.835 38.780 95.125 39.020 ;
        RECT 96.245 38.780 96.935 38.800 ;
        RECT 94.835 38.340 96.935 38.780 ;
        RECT 94.835 38.150 95.125 38.340 ;
        RECT 94.205 37.600 94.825 37.960 ;
        RECT 96.245 37.630 96.935 38.340 ;
        RECT 93.425 36.440 93.805 37.040 ;
        RECT 94.215 36.730 94.645 37.600 ;
        RECT 93.495 35.250 93.725 36.440 ;
        RECT 94.215 36.310 96.095 36.730 ;
        RECT 94.215 35.780 94.645 36.310 ;
        RECT 94.065 35.420 94.685 35.780 ;
        RECT 93.495 35.240 93.975 35.250 ;
        RECT 93.495 34.560 94.055 35.240 ;
        RECT 93.585 34.410 94.055 34.560 ;
        RECT 93.785 33.460 94.055 34.410 ;
        RECT 94.695 34.160 94.965 35.160 ;
        RECT 94.695 33.430 95.205 34.160 ;
        RECT 94.695 33.340 95.195 33.430 ;
        RECT 90.055 32.790 90.585 33.170 ;
        RECT 87.045 31.110 89.875 32.160 ;
        RECT 90.155 31.910 90.415 32.790 ;
        RECT 90.135 31.290 90.495 31.910 ;
        RECT 94.945 31.220 95.195 33.340 ;
        RECT 87.045 30.200 87.365 31.110 ;
        RECT 88.725 31.100 89.855 31.110 ;
        RECT 90.755 30.820 95.395 31.220 ;
        RECT 94.945 30.540 95.195 30.820 ;
        RECT 87.045 30.140 87.375 30.200 ;
        RECT 87.055 20.210 87.375 30.140 ;
        RECT 88.375 28.890 88.645 30.250 ;
        RECT 89.505 28.890 89.775 30.210 ;
        RECT 94.815 30.110 95.195 30.540 ;
        RECT 94.815 29.600 95.175 30.110 ;
        RECT 88.375 22.200 89.775 28.890 ;
        RECT 88.375 20.200 88.645 22.200 ;
        RECT 89.505 20.160 89.775 22.200 ;
        RECT 94.825 21.760 95.085 29.600 ;
        RECT 94.825 20.210 95.205 21.760 ;
        RECT 87.345 19.550 88.395 19.960 ;
        RECT 89.755 19.560 94.805 19.940 ;
        RECT 87.515 18.270 88.185 19.550 ;
        RECT 87.345 17.590 88.465 18.270 ;
        RECT 73.865 12.750 74.725 13.590 ;
        RECT 61.415 10.960 63.435 12.160 ;
        RECT 72.725 10.990 74.745 12.190 ;
        RECT 84.465 12.180 84.875 14.780 ;
        RECT 85.175 13.580 85.715 16.810 ;
        RECT 91.435 16.780 93.365 19.560 ;
        RECT 90.855 15.930 93.565 16.780 ;
        RECT 94.945 15.390 95.205 20.210 ;
        RECT 94.415 14.660 95.305 15.390 ;
        RECT 95.705 14.800 96.095 36.310 ;
        RECT 96.435 16.830 96.935 37.630 ;
        RECT 98.975 38.500 99.255 40.490 ;
        RECT 101.545 40.420 102.645 41.190 ;
        RECT 110.155 40.530 110.455 42.260 ;
        RECT 99.525 39.660 99.905 40.260 ;
        RECT 99.555 39.040 99.805 39.660 ;
        RECT 99.425 38.660 99.905 39.040 ;
        RECT 98.975 33.430 99.305 38.500 ;
        RECT 99.855 37.640 100.155 38.500 ;
        RECT 100.935 37.640 101.235 38.500 ;
        RECT 101.845 38.460 102.125 40.420 ;
        RECT 105.145 38.850 105.415 39.020 ;
        RECT 104.755 38.540 105.415 38.850 ;
        RECT 99.855 33.400 101.235 37.640 ;
        RECT 101.785 38.410 102.125 38.460 ;
        RECT 104.705 38.430 105.415 38.540 ;
        RECT 98.255 32.180 98.575 32.200 ;
        RECT 99.935 32.180 101.065 33.400 ;
        RECT 101.785 33.390 102.115 38.410 ;
        RECT 104.705 37.060 104.935 38.430 ;
        RECT 105.145 38.180 105.415 38.430 ;
        RECT 106.045 38.800 106.335 39.040 ;
        RECT 107.455 38.800 108.145 38.820 ;
        RECT 106.045 38.360 108.145 38.800 ;
        RECT 106.045 38.170 106.335 38.360 ;
        RECT 105.415 37.620 106.035 37.980 ;
        RECT 107.455 37.650 108.145 38.360 ;
        RECT 104.635 36.460 105.015 37.060 ;
        RECT 105.425 36.750 105.855 37.620 ;
        RECT 104.705 35.270 104.935 36.460 ;
        RECT 105.425 36.330 107.305 36.750 ;
        RECT 105.425 35.800 105.855 36.330 ;
        RECT 105.275 35.440 105.895 35.800 ;
        RECT 104.705 35.260 105.185 35.270 ;
        RECT 104.705 34.580 105.265 35.260 ;
        RECT 104.795 34.430 105.265 34.580 ;
        RECT 104.995 33.480 105.265 34.430 ;
        RECT 105.905 34.180 106.175 35.180 ;
        RECT 105.905 33.450 106.415 34.180 ;
        RECT 105.905 33.360 106.405 33.450 ;
        RECT 101.265 32.810 101.795 33.190 ;
        RECT 98.255 31.130 101.085 32.180 ;
        RECT 101.365 31.930 101.625 32.810 ;
        RECT 101.345 31.310 101.705 31.930 ;
        RECT 106.155 31.240 106.405 33.360 ;
        RECT 98.255 30.220 98.575 31.130 ;
        RECT 99.935 31.120 101.065 31.130 ;
        RECT 101.965 30.840 106.605 31.240 ;
        RECT 106.155 30.560 106.405 30.840 ;
        RECT 98.255 30.160 98.585 30.220 ;
        RECT 98.265 20.230 98.585 30.160 ;
        RECT 99.585 28.910 99.855 30.270 ;
        RECT 100.715 28.910 100.985 30.230 ;
        RECT 106.025 30.130 106.405 30.560 ;
        RECT 106.025 29.620 106.385 30.130 ;
        RECT 99.585 22.220 100.985 28.910 ;
        RECT 99.585 20.220 99.855 22.220 ;
        RECT 100.715 20.180 100.985 22.220 ;
        RECT 106.035 21.780 106.295 29.620 ;
        RECT 106.035 20.230 106.415 21.780 ;
        RECT 98.555 19.570 99.605 19.980 ;
        RECT 100.965 19.580 106.015 19.960 ;
        RECT 98.725 18.290 99.395 19.570 ;
        RECT 98.555 17.610 99.675 18.290 ;
        RECT 85.155 12.740 86.015 13.580 ;
        RECT 95.705 12.180 96.115 14.800 ;
        RECT 96.415 13.600 96.955 16.830 ;
        RECT 102.645 16.800 104.575 19.580 ;
        RECT 102.065 15.950 104.775 16.800 ;
        RECT 106.155 15.410 106.415 20.230 ;
        RECT 105.625 14.680 106.515 15.410 ;
        RECT 106.915 14.820 107.305 36.330 ;
        RECT 107.645 16.850 108.145 37.650 ;
        RECT 110.175 38.540 110.455 40.530 ;
        RECT 112.745 40.460 113.845 41.230 ;
        RECT 121.365 40.550 121.665 42.280 ;
        RECT 142.880 42.020 144.100 43.390 ;
        RECT 110.725 39.700 111.105 40.300 ;
        RECT 110.755 39.080 111.005 39.700 ;
        RECT 110.625 38.700 111.105 39.080 ;
        RECT 110.175 33.470 110.505 38.540 ;
        RECT 111.055 37.680 111.355 38.540 ;
        RECT 112.135 37.680 112.435 38.540 ;
        RECT 113.045 38.500 113.325 40.460 ;
        RECT 116.345 38.890 116.615 39.060 ;
        RECT 115.955 38.580 116.615 38.890 ;
        RECT 111.055 33.440 112.435 37.680 ;
        RECT 112.985 38.450 113.325 38.500 ;
        RECT 115.905 38.470 116.615 38.580 ;
        RECT 109.455 32.220 109.775 32.240 ;
        RECT 111.135 32.220 112.265 33.440 ;
        RECT 112.985 33.430 113.315 38.450 ;
        RECT 115.905 37.100 116.135 38.470 ;
        RECT 116.345 38.220 116.615 38.470 ;
        RECT 117.245 38.840 117.535 39.080 ;
        RECT 118.655 38.840 119.345 38.860 ;
        RECT 117.245 38.400 119.345 38.840 ;
        RECT 117.245 38.210 117.535 38.400 ;
        RECT 116.615 37.660 117.235 38.020 ;
        RECT 118.655 37.690 119.345 38.400 ;
        RECT 115.835 36.500 116.215 37.100 ;
        RECT 116.625 36.790 117.055 37.660 ;
        RECT 115.905 35.310 116.135 36.500 ;
        RECT 116.625 36.370 118.505 36.790 ;
        RECT 116.625 35.840 117.055 36.370 ;
        RECT 116.475 35.480 117.095 35.840 ;
        RECT 115.905 35.300 116.385 35.310 ;
        RECT 115.905 34.620 116.465 35.300 ;
        RECT 115.995 34.470 116.465 34.620 ;
        RECT 116.195 33.520 116.465 34.470 ;
        RECT 117.105 34.220 117.375 35.220 ;
        RECT 117.105 33.490 117.615 34.220 ;
        RECT 117.105 33.400 117.605 33.490 ;
        RECT 112.465 32.850 112.995 33.230 ;
        RECT 109.455 31.170 112.285 32.220 ;
        RECT 112.565 31.970 112.825 32.850 ;
        RECT 112.545 31.350 112.905 31.970 ;
        RECT 117.355 31.280 117.605 33.400 ;
        RECT 109.455 30.260 109.775 31.170 ;
        RECT 111.135 31.160 112.265 31.170 ;
        RECT 113.165 30.880 117.805 31.280 ;
        RECT 117.355 30.600 117.605 30.880 ;
        RECT 109.455 30.200 109.785 30.260 ;
        RECT 109.465 20.270 109.785 30.200 ;
        RECT 110.785 28.950 111.055 30.310 ;
        RECT 111.915 28.950 112.185 30.270 ;
        RECT 117.225 30.170 117.605 30.600 ;
        RECT 117.225 29.660 117.585 30.170 ;
        RECT 110.785 22.260 112.185 28.950 ;
        RECT 110.785 20.260 111.055 22.260 ;
        RECT 111.915 20.220 112.185 22.260 ;
        RECT 117.235 21.820 117.495 29.660 ;
        RECT 117.235 20.270 117.615 21.820 ;
        RECT 109.755 19.610 110.805 20.020 ;
        RECT 112.165 19.620 117.215 20.000 ;
        RECT 109.925 18.330 110.595 19.610 ;
        RECT 109.755 17.650 110.875 18.330 ;
        RECT 96.395 12.760 97.255 13.600 ;
        RECT 106.915 12.230 107.325 14.820 ;
        RECT 107.625 13.620 108.165 16.850 ;
        RECT 113.845 16.840 115.775 19.620 ;
        RECT 113.265 15.990 115.975 16.840 ;
        RECT 117.355 15.450 117.615 20.270 ;
        RECT 116.825 14.720 117.715 15.450 ;
        RECT 118.115 14.860 118.505 36.370 ;
        RECT 118.845 16.890 119.345 37.690 ;
        RECT 121.385 38.560 121.665 40.550 ;
        RECT 123.955 40.480 125.055 41.250 ;
        RECT 121.935 39.720 122.315 40.320 ;
        RECT 121.965 39.100 122.215 39.720 ;
        RECT 121.835 38.720 122.315 39.100 ;
        RECT 121.385 33.490 121.715 38.560 ;
        RECT 122.265 37.700 122.565 38.560 ;
        RECT 123.345 37.700 123.645 38.560 ;
        RECT 124.255 38.520 124.535 40.480 ;
        RECT 127.555 38.910 127.825 39.080 ;
        RECT 127.165 38.600 127.825 38.910 ;
        RECT 122.265 33.460 123.645 37.700 ;
        RECT 124.195 38.470 124.535 38.520 ;
        RECT 127.115 38.490 127.825 38.600 ;
        RECT 120.665 32.240 120.985 32.260 ;
        RECT 122.345 32.240 123.475 33.460 ;
        RECT 124.195 33.450 124.525 38.470 ;
        RECT 127.115 37.120 127.345 38.490 ;
        RECT 127.555 38.240 127.825 38.490 ;
        RECT 128.455 38.860 128.745 39.100 ;
        RECT 142.940 38.950 144.100 42.020 ;
        RECT 129.865 38.860 130.555 38.880 ;
        RECT 128.455 38.420 130.555 38.860 ;
        RECT 128.455 38.230 128.745 38.420 ;
        RECT 127.825 37.680 128.445 38.040 ;
        RECT 129.865 37.710 130.555 38.420 ;
        RECT 127.045 36.520 127.425 37.120 ;
        RECT 127.835 36.810 128.265 37.680 ;
        RECT 127.115 35.330 127.345 36.520 ;
        RECT 127.835 36.390 129.715 36.810 ;
        RECT 127.835 35.860 128.265 36.390 ;
        RECT 127.685 35.500 128.305 35.860 ;
        RECT 127.115 35.320 127.595 35.330 ;
        RECT 127.115 34.640 127.675 35.320 ;
        RECT 127.205 34.490 127.675 34.640 ;
        RECT 127.405 33.540 127.675 34.490 ;
        RECT 128.315 34.240 128.585 35.240 ;
        RECT 128.315 33.510 128.825 34.240 ;
        RECT 128.315 33.420 128.815 33.510 ;
        RECT 123.675 32.870 124.205 33.250 ;
        RECT 120.665 31.190 123.495 32.240 ;
        RECT 123.775 31.990 124.035 32.870 ;
        RECT 123.755 31.370 124.115 31.990 ;
        RECT 128.565 31.300 128.815 33.420 ;
        RECT 120.665 30.280 120.985 31.190 ;
        RECT 122.345 31.180 123.475 31.190 ;
        RECT 124.375 30.900 129.015 31.300 ;
        RECT 128.565 30.620 128.815 30.900 ;
        RECT 120.665 30.220 120.995 30.280 ;
        RECT 120.675 20.290 120.995 30.220 ;
        RECT 121.995 28.970 122.265 30.330 ;
        RECT 123.125 28.970 123.395 30.290 ;
        RECT 128.435 30.190 128.815 30.620 ;
        RECT 128.435 29.680 128.795 30.190 ;
        RECT 121.995 22.280 123.395 28.970 ;
        RECT 121.995 20.280 122.265 22.280 ;
        RECT 123.125 20.240 123.395 22.280 ;
        RECT 128.445 21.840 128.705 29.680 ;
        RECT 128.445 20.290 128.825 21.840 ;
        RECT 120.965 19.630 122.015 20.040 ;
        RECT 123.375 19.640 128.425 20.020 ;
        RECT 121.135 18.350 121.805 19.630 ;
        RECT 120.965 17.670 122.085 18.350 ;
        RECT 107.605 12.780 108.465 13.620 ;
        RECT 118.115 12.230 118.525 14.860 ;
        RECT 118.825 13.660 119.365 16.890 ;
        RECT 125.055 16.860 126.985 19.640 ;
        RECT 124.475 16.010 127.185 16.860 ;
        RECT 128.565 15.470 128.825 20.290 ;
        RECT 128.035 14.740 128.925 15.470 ;
        RECT 129.325 14.880 129.715 36.390 ;
        RECT 130.055 16.910 130.555 37.710 ;
        RECT 142.900 37.580 144.120 38.950 ;
        RECT 132.395 24.340 132.705 30.230 ;
        RECT 132.195 20.120 132.705 24.340 ;
        RECT 118.805 12.820 119.665 13.660 ;
        RECT 129.325 12.260 129.735 14.880 ;
        RECT 130.035 13.680 130.575 16.910 ;
        RECT 132.195 15.510 132.505 20.120 ;
        RECT 137.715 19.980 138.005 30.170 ;
        RECT 132.685 19.590 138.005 19.980 ;
        RECT 137.715 16.940 138.005 19.590 ;
        RECT 142.940 17.940 144.090 19.160 ;
        RECT 145.080 18.760 146.200 18.930 ;
        RECT 137.395 15.890 138.295 16.940 ;
        RECT 137.715 15.720 138.005 15.890 ;
        RECT 131.975 14.270 132.735 15.510 ;
        RECT 142.940 15.090 144.050 17.940 ;
        RECT 142.900 13.870 144.050 15.090 ;
        RECT 145.070 14.920 146.200 18.760 ;
        RECT 145.030 13.970 146.200 14.920 ;
        RECT 145.030 13.900 146.150 13.970 ;
        RECT 130.015 12.840 130.875 13.680 ;
        RECT 83.845 10.980 85.865 12.180 ;
        RECT 95.145 10.980 97.165 12.180 ;
        RECT 106.335 11.030 108.355 12.230 ;
        RECT 117.565 11.030 119.585 12.230 ;
        RECT 128.865 11.060 130.885 12.260 ;
        RECT 74.340 0.110 75.630 1.460 ;
        RECT 93.550 0.180 94.840 1.530 ;
        RECT 112.950 0.310 114.240 1.660 ;
        RECT 131.850 0.380 133.490 1.930 ;
        RECT 151.650 0.250 152.920 1.470 ;
      LAYER met3 ;
        RECT 135.340 223.855 136.790 225.205 ;
        RECT 138.130 223.785 139.580 225.135 ;
        RECT 143.180 223.815 144.630 225.165 ;
        RECT 53.185 193.455 54.765 193.785 ;
        RECT 92.055 193.455 93.635 193.785 ;
        RECT 17.615 190.735 19.195 191.065 ;
        RECT 56.485 190.735 58.065 191.065 ;
        RECT 95.355 190.735 96.935 191.065 ;
        RECT 53.185 188.015 54.765 188.345 ;
        RECT 92.055 188.015 93.635 188.345 ;
        RECT 17.615 185.295 19.195 185.625 ;
        RECT 56.485 185.295 58.065 185.625 ;
        RECT 95.355 185.295 96.935 185.625 ;
        RECT 86.770 183.230 87.100 183.245 ;
        RECT 89.990 183.230 90.320 183.245 ;
        RECT 86.770 182.930 90.320 183.230 ;
        RECT 86.770 182.915 87.100 182.930 ;
        RECT 89.990 182.915 90.320 182.930 ;
        RECT 53.185 182.575 54.765 182.905 ;
        RECT 92.055 182.575 93.635 182.905 ;
        RECT 17.615 179.855 19.195 180.185 ;
        RECT 56.485 179.855 58.065 180.185 ;
        RECT 95.355 179.855 96.935 180.185 ;
        RECT 20.070 179.150 20.400 179.165 ;
        RECT 33.410 179.150 33.740 179.165 ;
        RECT 38.010 179.150 38.340 179.165 ;
        RECT 20.070 178.850 38.340 179.150 ;
        RECT 20.070 178.835 20.400 178.850 ;
        RECT 33.410 178.835 33.740 178.850 ;
        RECT 38.010 178.835 38.340 178.850 ;
        RECT 51.810 179.150 52.140 179.165 ;
        RECT 74.350 179.150 74.680 179.165 ;
        RECT 51.810 178.850 74.680 179.150 ;
        RECT 51.810 178.835 52.140 178.850 ;
        RECT 74.350 178.835 74.680 178.850 ;
        RECT 78.030 179.150 78.360 179.165 ;
        RECT 91.370 179.150 91.700 179.165 ;
        RECT 92.750 179.150 93.080 179.165 ;
        RECT 78.030 178.850 93.080 179.150 ;
        RECT 78.030 178.835 78.360 178.850 ;
        RECT 91.370 178.835 91.700 178.850 ;
        RECT 92.750 178.835 93.080 178.850 ;
        RECT 23.290 178.470 23.620 178.485 ;
        RECT 52.015 178.470 52.395 178.480 ;
        RECT 59.630 178.470 59.960 178.485 ;
        RECT 23.290 178.170 59.960 178.470 ;
        RECT 23.290 178.155 23.620 178.170 ;
        RECT 52.015 178.160 52.395 178.170 ;
        RECT 59.630 178.155 59.960 178.170 ;
        RECT 57.790 177.790 58.120 177.805 ;
        RECT 65.150 177.790 65.480 177.805 ;
        RECT 57.790 177.490 65.480 177.790 ;
        RECT 57.790 177.475 58.120 177.490 ;
        RECT 65.150 177.475 65.480 177.490 ;
        RECT 53.185 177.135 54.765 177.465 ;
        RECT 92.055 177.135 93.635 177.465 ;
        RECT 55.490 177.110 55.820 177.125 ;
        RECT 64.230 177.110 64.560 177.125 ;
        RECT 55.490 176.810 64.560 177.110 ;
        RECT 55.490 176.795 55.820 176.810 ;
        RECT 64.230 176.795 64.560 176.810 ;
        RECT 71.590 177.110 71.920 177.125 ;
        RECT 81.710 177.110 82.040 177.125 ;
        RECT 71.590 176.810 82.040 177.110 ;
        RECT 71.590 176.795 71.920 176.810 ;
        RECT 81.710 176.795 82.040 176.810 ;
        RECT 24.210 176.430 24.540 176.445 ;
        RECT 39.390 176.430 39.720 176.445 ;
        RECT 24.210 176.130 39.720 176.430 ;
        RECT 24.210 176.115 24.540 176.130 ;
        RECT 39.390 176.115 39.720 176.130 ;
        RECT 41.690 176.430 42.020 176.445 ;
        RECT 57.790 176.430 58.120 176.445 ;
        RECT 41.690 176.130 58.120 176.430 ;
        RECT 41.690 176.115 42.020 176.130 ;
        RECT 57.790 176.115 58.120 176.130 ;
        RECT 58.710 176.430 59.040 176.445 ;
        RECT 75.730 176.430 76.060 176.445 ;
        RECT 58.710 176.130 76.060 176.430 ;
        RECT 58.710 176.115 59.040 176.130 ;
        RECT 75.730 176.115 76.060 176.130 ;
        RECT 71.130 175.750 71.460 175.765 ;
        RECT 76.650 175.750 76.980 175.765 ;
        RECT 89.990 175.750 90.320 175.765 ;
        RECT 71.130 175.450 90.320 175.750 ;
        RECT 71.130 175.435 71.460 175.450 ;
        RECT 76.650 175.435 76.980 175.450 ;
        RECT 89.990 175.435 90.320 175.450 ;
        RECT 17.615 174.415 19.195 174.745 ;
        RECT 56.485 174.415 58.065 174.745 ;
        RECT 95.355 174.415 96.935 174.745 ;
        RECT 35.455 173.710 35.835 173.720 ;
        RECT 36.170 173.710 36.500 173.725 ;
        RECT 35.455 173.410 36.500 173.710 ;
        RECT 35.455 173.400 35.835 173.410 ;
        RECT 36.170 173.395 36.500 173.410 ;
        RECT 56.870 173.710 57.200 173.725 ;
        RECT 60.090 173.710 60.420 173.725 ;
        RECT 56.870 173.410 60.420 173.710 ;
        RECT 56.870 173.395 57.200 173.410 ;
        RECT 60.090 173.395 60.420 173.410 ;
        RECT 32.950 173.030 33.280 173.045 ;
        RECT 41.690 173.030 42.020 173.045 ;
        RECT 32.950 172.730 42.020 173.030 ;
        RECT 32.950 172.715 33.280 172.730 ;
        RECT 41.690 172.715 42.020 172.730 ;
        RECT 55.490 173.030 55.820 173.045 ;
        RECT 58.250 173.030 58.580 173.045 ;
        RECT 55.490 172.730 58.580 173.030 ;
        RECT 55.490 172.715 55.820 172.730 ;
        RECT 58.250 172.715 58.580 172.730 ;
        RECT 133.700 172.500 134.930 172.705 ;
        RECT 53.185 171.695 54.765 172.025 ;
        RECT 92.055 171.695 93.635 172.025 ;
        RECT 129.030 170.130 134.930 172.500 ;
        RECT 133.700 170.095 134.930 170.130 ;
        RECT 21.450 169.630 21.780 169.645 ;
        RECT 32.695 169.630 33.075 169.640 ;
        RECT 21.450 169.330 33.075 169.630 ;
        RECT 21.450 169.315 21.780 169.330 ;
        RECT 32.695 169.320 33.075 169.330 ;
        RECT 36.375 169.630 36.755 169.640 ;
        RECT 37.090 169.630 37.420 169.645 ;
        RECT 36.375 169.330 37.420 169.630 ;
        RECT 36.375 169.320 36.755 169.330 ;
        RECT 37.090 169.315 37.420 169.330 ;
        RECT 17.615 168.975 19.195 169.305 ;
        RECT 56.485 168.975 58.065 169.305 ;
        RECT 95.355 168.975 96.935 169.305 ;
        RECT 89.990 167.590 90.320 167.605 ;
        RECT 91.370 167.590 91.700 167.605 ;
        RECT 89.990 167.290 91.700 167.590 ;
        RECT 89.990 167.275 90.320 167.290 ;
        RECT 91.370 167.275 91.700 167.290 ;
        RECT 53.185 166.255 54.765 166.585 ;
        RECT 92.055 166.255 93.635 166.585 ;
        RECT 15.225 165.550 17.225 165.700 ;
        RECT 19.610 165.550 19.940 165.565 ;
        RECT 15.225 165.250 19.940 165.550 ;
        RECT 15.225 165.100 17.225 165.250 ;
        RECT 19.610 165.235 19.940 165.250 ;
        RECT 23.750 165.550 24.080 165.565 ;
        RECT 34.790 165.550 35.120 165.565 ;
        RECT 60.550 165.550 60.880 165.565 ;
        RECT 23.750 165.250 60.880 165.550 ;
        RECT 23.750 165.235 24.080 165.250 ;
        RECT 34.790 165.235 35.120 165.250 ;
        RECT 60.550 165.235 60.880 165.250 ;
        RECT 17.615 163.535 19.195 163.865 ;
        RECT 56.485 163.535 58.065 163.865 ;
        RECT 95.355 163.535 96.935 163.865 ;
        RECT 59.170 162.150 59.500 162.165 ;
        RECT 61.930 162.150 62.260 162.165 ;
        RECT 59.170 161.850 62.260 162.150 ;
        RECT 59.170 161.835 59.500 161.850 ;
        RECT 61.930 161.835 62.260 161.850 ;
        RECT 53.185 160.815 54.765 161.145 ;
        RECT 92.055 160.815 93.635 161.145 ;
        RECT 16.135 160.110 16.515 160.120 ;
        RECT 22.370 160.110 22.700 160.125 ;
        RECT 16.135 159.810 22.700 160.110 ;
        RECT 16.135 159.800 16.515 159.810 ;
        RECT 22.370 159.795 22.700 159.810 ;
        RECT 91.370 160.110 91.700 160.125 ;
        RECT 101.490 160.110 101.820 160.125 ;
        RECT 91.370 159.810 101.820 160.110 ;
        RECT 91.370 159.795 91.700 159.810 ;
        RECT 101.490 159.795 101.820 159.810 ;
        RECT 15.225 158.300 17.225 158.900 ;
        RECT 17.615 158.095 19.195 158.425 ;
        RECT 56.485 158.095 58.065 158.425 ;
        RECT 95.355 158.095 96.935 158.425 ;
        RECT 43.530 156.710 43.860 156.725 ;
        RECT 63.310 156.710 63.640 156.725 ;
        RECT 43.530 156.410 63.640 156.710 ;
        RECT 43.530 156.395 43.860 156.410 ;
        RECT 63.310 156.395 63.640 156.410 ;
        RECT 15.225 155.350 17.225 155.500 ;
        RECT 53.185 155.375 54.765 155.705 ;
        RECT 92.055 155.375 93.635 155.705 ;
        RECT 22.370 155.350 22.700 155.365 ;
        RECT 15.225 155.050 22.700 155.350 ;
        RECT 15.225 154.900 17.225 155.050 ;
        RECT 22.370 155.035 22.700 155.050 ;
        RECT 110.690 155.350 111.020 155.365 ;
        RECT 113.225 155.350 115.225 155.500 ;
        RECT 110.690 155.050 115.225 155.350 ;
        RECT 110.690 155.035 111.020 155.050 ;
        RECT 113.225 154.900 115.225 155.050 ;
        RECT 49.510 154.670 49.840 154.685 ;
        RECT 58.250 154.670 58.580 154.685 ;
        RECT 49.510 154.370 58.580 154.670 ;
        RECT 49.510 154.355 49.840 154.370 ;
        RECT 58.250 154.355 58.580 154.370 ;
        RECT 37.550 153.990 37.880 154.005 ;
        RECT 59.630 153.990 59.960 154.005 ;
        RECT 37.550 153.690 59.960 153.990 ;
        RECT 37.550 153.675 37.880 153.690 ;
        RECT 59.630 153.675 59.960 153.690 ;
        RECT 17.615 152.655 19.195 152.985 ;
        RECT 56.485 152.655 58.065 152.985 ;
        RECT 95.355 152.655 96.935 152.985 ;
        RECT 53.185 149.935 54.765 150.265 ;
        RECT 92.055 149.935 93.635 150.265 ;
        RECT 38.010 149.230 38.340 149.245 ;
        RECT 63.770 149.230 64.100 149.245 ;
        RECT 38.010 148.930 64.100 149.230 ;
        RECT 38.010 148.915 38.340 148.930 ;
        RECT 63.770 148.915 64.100 148.930 ;
        RECT 15.225 148.550 17.225 148.700 ;
        RECT 22.370 148.550 22.700 148.565 ;
        RECT 15.225 148.250 22.700 148.550 ;
        RECT 15.225 148.100 17.225 148.250 ;
        RECT 22.370 148.235 22.700 148.250 ;
        RECT 39.390 148.550 39.720 148.565 ;
        RECT 43.990 148.550 44.320 148.565 ;
        RECT 61.470 148.550 61.800 148.565 ;
        RECT 39.390 148.250 61.800 148.550 ;
        RECT 39.390 148.235 39.720 148.250 ;
        RECT 43.990 148.235 44.320 148.250 ;
        RECT 61.470 148.235 61.800 148.250 ;
        RECT 17.615 147.215 19.195 147.545 ;
        RECT 56.485 147.215 58.065 147.545 ;
        RECT 95.355 147.215 96.935 147.545 ;
        RECT 110.690 145.150 111.020 145.165 ;
        RECT 113.225 145.150 115.225 145.300 ;
        RECT 110.690 144.850 115.225 145.150 ;
        RECT 110.690 144.835 111.020 144.850 ;
        RECT 53.185 144.495 54.765 144.825 ;
        RECT 92.055 144.495 93.635 144.825 ;
        RECT 113.225 144.700 115.225 144.850 ;
        RECT 17.615 141.775 19.195 142.105 ;
        RECT 56.485 141.775 58.065 142.105 ;
        RECT 95.355 141.775 96.935 142.105 ;
        RECT 110.690 141.750 111.020 141.765 ;
        RECT 113.225 141.750 115.225 141.900 ;
        RECT 110.690 141.450 115.225 141.750 ;
        RECT 110.690 141.435 111.020 141.450 ;
        RECT 113.225 141.300 115.225 141.450 ;
        RECT 42.150 141.070 42.480 141.085 ;
        RECT 78.030 141.070 78.360 141.085 ;
        RECT 42.150 140.770 78.360 141.070 ;
        RECT 42.150 140.755 42.480 140.770 ;
        RECT 78.030 140.755 78.360 140.770 ;
        RECT 53.185 139.055 54.765 139.385 ;
        RECT 92.055 139.055 93.635 139.385 ;
        RECT 38.930 138.350 39.260 138.365 ;
        RECT 43.530 138.350 43.860 138.365 ;
        RECT 52.015 138.350 52.395 138.360 ;
        RECT 63.310 138.350 63.640 138.365 ;
        RECT 38.930 138.050 63.640 138.350 ;
        RECT 132.510 138.165 135.210 140.035 ;
        RECT 38.930 138.035 39.260 138.050 ;
        RECT 43.530 138.035 43.860 138.050 ;
        RECT 52.015 138.040 52.395 138.050 ;
        RECT 63.310 138.035 63.640 138.050 ;
        RECT 17.615 136.335 19.195 136.665 ;
        RECT 56.485 136.335 58.065 136.665 ;
        RECT 95.355 136.335 96.935 136.665 ;
        RECT 64.230 135.630 64.560 135.645 ;
        RECT 100.570 135.630 100.900 135.645 ;
        RECT 64.230 135.330 100.900 135.630 ;
        RECT 64.230 135.315 64.560 135.330 ;
        RECT 100.570 135.315 100.900 135.330 ;
        RECT 54.570 134.950 54.900 134.965 ;
        RECT 87.230 134.950 87.560 134.965 ;
        RECT 54.570 134.650 87.560 134.950 ;
        RECT 54.570 134.635 54.900 134.650 ;
        RECT 87.230 134.635 87.560 134.650 ;
        RECT 110.690 134.950 111.020 134.965 ;
        RECT 113.225 134.950 115.225 135.100 ;
        RECT 110.690 134.650 115.225 134.950 ;
        RECT 110.690 134.635 111.020 134.650 ;
        RECT 113.225 134.500 115.225 134.650 ;
        RECT 53.185 133.615 54.765 133.945 ;
        RECT 92.055 133.615 93.635 133.945 ;
        RECT 37.090 132.910 37.420 132.925 ;
        RECT 58.710 132.910 59.040 132.925 ;
        RECT 37.090 132.610 59.040 132.910 ;
        RECT 37.090 132.595 37.420 132.610 ;
        RECT 58.710 132.595 59.040 132.610 ;
        RECT 21.450 132.230 21.780 132.245 ;
        RECT 64.230 132.230 64.560 132.245 ;
        RECT 21.450 131.930 64.560 132.230 ;
        RECT 21.450 131.915 21.780 131.930 ;
        RECT 64.230 131.915 64.560 131.930 ;
        RECT 17.615 130.895 19.195 131.225 ;
        RECT 56.485 130.895 58.065 131.225 ;
        RECT 95.355 130.895 96.935 131.225 ;
        RECT 53.185 128.175 54.765 128.505 ;
        RECT 92.055 128.175 93.635 128.505 ;
        RECT 36.630 126.790 36.960 126.805 ;
        RECT 53.190 126.790 53.520 126.805 ;
        RECT 36.630 126.490 53.520 126.790 ;
        RECT 36.630 126.475 36.960 126.490 ;
        RECT 53.190 126.475 53.520 126.490 ;
        RECT 78.490 126.790 78.820 126.805 ;
        RECT 95.510 126.790 95.840 126.805 ;
        RECT 78.490 126.490 95.840 126.790 ;
        RECT 78.490 126.475 78.820 126.490 ;
        RECT 95.510 126.475 95.840 126.490 ;
        RECT 17.615 125.455 19.195 125.785 ;
        RECT 56.485 125.455 58.065 125.785 ;
        RECT 95.355 125.455 96.935 125.785 ;
        RECT 86.310 125.430 86.640 125.445 ;
        RECT 86.310 125.130 87.315 125.430 ;
        RECT 86.310 125.115 86.640 125.130 ;
        RECT 15.225 124.750 17.225 124.900 ;
        RECT 19.610 124.750 19.940 124.765 ;
        RECT 15.225 124.450 19.940 124.750 ;
        RECT 15.225 124.300 17.225 124.450 ;
        RECT 19.610 124.435 19.940 124.450 ;
        RECT 36.375 124.750 36.755 124.760 ;
        RECT 60.550 124.750 60.880 124.765 ;
        RECT 36.375 124.450 60.880 124.750 ;
        RECT 36.375 124.440 36.755 124.450 ;
        RECT 60.550 124.435 60.880 124.450 ;
        RECT 87.015 124.085 87.315 125.130 ;
        RECT 24.670 124.070 25.000 124.085 ;
        RECT 35.455 124.070 35.835 124.080 ;
        RECT 62.390 124.070 62.720 124.085 ;
        RECT 24.670 123.770 62.720 124.070 ;
        RECT 24.670 123.755 25.000 123.770 ;
        RECT 35.455 123.760 35.835 123.770 ;
        RECT 62.390 123.755 62.720 123.770 ;
        RECT 86.770 123.770 87.315 124.085 ;
        RECT 86.770 123.755 87.100 123.770 ;
        RECT 53.185 122.735 54.765 123.065 ;
        RECT 92.055 122.735 93.635 123.065 ;
        RECT 34.790 122.030 35.120 122.045 ;
        RECT 59.630 122.030 59.960 122.045 ;
        RECT 34.790 121.730 59.960 122.030 ;
        RECT 34.790 121.715 35.120 121.730 ;
        RECT 59.630 121.715 59.960 121.730 ;
        RECT 15.225 121.350 17.225 121.500 ;
        RECT 22.370 121.350 22.700 121.365 ;
        RECT 15.225 121.050 22.700 121.350 ;
        RECT 15.225 120.900 17.225 121.050 ;
        RECT 22.370 121.035 22.700 121.050 ;
        RECT 17.615 120.015 19.195 120.345 ;
        RECT 56.485 120.015 58.065 120.345 ;
        RECT 95.355 120.015 96.935 120.345 ;
        RECT 28.350 119.310 28.680 119.325 ;
        RECT 36.170 119.310 36.500 119.325 ;
        RECT 38.470 119.310 38.800 119.325 ;
        RECT 61.930 119.310 62.260 119.325 ;
        RECT 66.530 119.310 66.860 119.325 ;
        RECT 28.350 119.010 66.860 119.310 ;
        RECT 28.350 118.995 28.680 119.010 ;
        RECT 36.170 118.995 36.500 119.010 ;
        RECT 38.470 118.995 38.800 119.010 ;
        RECT 61.930 118.995 62.260 119.010 ;
        RECT 66.530 118.995 66.860 119.010 ;
        RECT 73.890 119.310 74.220 119.325 ;
        RECT 88.610 119.310 88.940 119.325 ;
        RECT 101.490 119.310 101.820 119.325 ;
        RECT 73.890 119.010 101.820 119.310 ;
        RECT 73.890 118.995 74.220 119.010 ;
        RECT 88.610 118.995 88.940 119.010 ;
        RECT 101.490 118.995 101.820 119.010 ;
        RECT 92.290 118.630 92.620 118.645 ;
        RECT 90.695 118.330 92.620 118.630 ;
        RECT 15.225 117.950 17.225 118.100 ;
        RECT 19.610 117.950 19.940 117.965 ;
        RECT 15.225 117.650 19.940 117.950 ;
        RECT 15.225 117.500 17.225 117.650 ;
        RECT 19.610 117.635 19.940 117.650 ;
        RECT 53.185 117.295 54.765 117.625 ;
        RECT 35.250 117.270 35.580 117.285 ;
        RECT 36.375 117.270 36.755 117.280 ;
        RECT 35.250 116.970 36.755 117.270 ;
        RECT 35.250 116.955 35.580 116.970 ;
        RECT 36.375 116.960 36.755 116.970 ;
        RECT 76.190 117.270 76.520 117.285 ;
        RECT 90.695 117.270 90.995 118.330 ;
        RECT 92.290 118.315 92.620 118.330 ;
        RECT 92.055 117.295 93.635 117.625 ;
        RECT 76.190 116.970 90.995 117.270 ;
        RECT 76.190 116.955 76.520 116.970 ;
        RECT 76.650 116.590 76.980 116.605 ;
        RECT 90.450 116.590 90.780 116.605 ;
        RECT 76.650 116.290 90.780 116.590 ;
        RECT 76.650 116.275 76.980 116.290 ;
        RECT 90.450 116.275 90.780 116.290 ;
        RECT 16.135 115.910 16.515 115.920 ;
        RECT 22.830 115.910 23.160 115.925 ;
        RECT 16.135 115.610 23.160 115.910 ;
        RECT 16.135 115.600 16.515 115.610 ;
        RECT 22.830 115.595 23.160 115.610 ;
        RECT 32.695 115.910 33.075 115.920 ;
        RECT 35.250 115.910 35.580 115.925 ;
        RECT 32.695 115.610 35.580 115.910 ;
        RECT 32.695 115.600 33.075 115.610 ;
        RECT 35.250 115.595 35.580 115.610 ;
        RECT 15.225 114.100 17.225 114.700 ;
        RECT 17.615 114.575 19.195 114.905 ;
        RECT 56.485 114.575 58.065 114.905 ;
        RECT 95.355 114.575 96.935 114.905 ;
        RECT 37.550 113.190 37.880 113.205 ;
        RECT 50.890 113.190 51.220 113.205 ;
        RECT 55.950 113.190 56.280 113.205 ;
        RECT 37.550 112.890 56.280 113.190 ;
        RECT 37.550 112.875 37.880 112.890 ;
        RECT 50.890 112.875 51.220 112.890 ;
        RECT 55.950 112.875 56.280 112.890 ;
        RECT 71.130 113.190 71.460 113.205 ;
        RECT 79.870 113.190 80.200 113.205 ;
        RECT 71.130 112.890 80.200 113.190 ;
        RECT 71.130 112.875 71.460 112.890 ;
        RECT 79.870 112.875 80.200 112.890 ;
        RECT 53.185 111.855 54.765 112.185 ;
        RECT 92.055 111.855 93.635 112.185 ;
        RECT 17.615 109.135 19.195 109.465 ;
        RECT 56.485 109.135 58.065 109.465 ;
        RECT 95.355 109.135 96.935 109.465 ;
        RECT 69.750 107.750 70.080 107.765 ;
        RECT 113.225 107.750 115.225 107.900 ;
        RECT 69.750 107.450 115.225 107.750 ;
        RECT 69.750 107.435 70.080 107.450 ;
        RECT 113.225 107.300 115.225 107.450 ;
        RECT 53.185 106.415 54.765 106.745 ;
        RECT 92.055 106.415 93.635 106.745 ;
        RECT 129.700 105.605 133.210 106.625 ;
        RECT 17.615 103.695 19.195 104.025 ;
        RECT 56.485 103.695 58.065 104.025 ;
        RECT 95.355 103.695 96.935 104.025 ;
        RECT 53.185 100.975 54.765 101.305 ;
        RECT 92.055 100.975 93.635 101.305 ;
        RECT 37.630 88.620 38.970 88.755 ;
        RECT 13.950 87.980 14.980 88.515 ;
        RECT 13.950 87.500 14.990 87.980 ;
        RECT 13.950 87.175 14.980 87.500 ;
        RECT 14.070 86.570 14.810 87.175 ;
        RECT 20.050 87.105 20.920 88.515 ;
        RECT 14.070 75.715 14.700 86.570 ;
        RECT 20.170 77.115 20.800 87.105 ;
        RECT 25.910 87.055 26.860 88.515 ;
        RECT 26.070 78.385 26.700 87.055 ;
        RECT 31.730 86.965 32.910 88.585 ;
        RECT 32.005 79.615 32.635 86.965 ;
        RECT 37.630 86.835 39.120 88.620 ;
        RECT 38.060 81.125 38.690 86.835 ;
        RECT 43.790 86.745 45.190 88.605 ;
        RECT 49.710 86.945 51.060 88.615 ;
        RECT 44.175 82.625 44.805 86.745 ;
        RECT 50.070 83.875 50.700 86.945 ;
        RECT 55.530 86.785 56.750 88.545 ;
        RECT 55.825 85.115 56.455 86.785 ;
        RECT 61.670 86.625 63.180 88.615 ;
        RECT 67.680 88.305 68.720 89.815 ;
        RECT 67.885 87.225 68.515 88.305 ;
        RECT 62.110 86.175 62.740 86.625 ;
        RECT 67.885 86.595 130.605 87.225 ;
        RECT 62.110 85.545 118.855 86.175 ;
        RECT 55.825 84.485 107.605 85.115 ;
        RECT 50.070 83.245 96.285 83.875 ;
        RECT 44.175 81.995 85.055 82.625 ;
        RECT 38.060 80.495 73.765 81.125 ;
        RECT 32.005 78.985 62.635 79.615 ;
        RECT 26.070 77.755 51.245 78.385 ;
        RECT 20.170 76.485 40.645 77.115 ;
        RECT 14.070 75.660 29.295 75.715 ;
        RECT 40.015 75.710 40.645 76.485 ;
        RECT 14.070 75.085 30.410 75.660 ;
        RECT 27.850 74.670 30.410 75.085 ;
        RECT 3.910 71.345 6.100 73.215 ;
        RECT 27.850 73.120 30.450 74.670 ;
        RECT 39.060 74.510 41.620 75.710 ;
        RECT 50.615 75.580 51.245 77.755 ;
        RECT 62.005 75.690 62.635 78.985 ;
        RECT 49.930 74.650 52.490 75.580 ;
        RECT 0.970 70.330 3.070 70.430 ;
        RECT 15.510 70.330 17.040 71.185 ;
        RECT 0.960 68.750 17.040 70.330 ;
        RECT 0.970 68.710 3.070 68.750 ;
        RECT 15.510 68.635 17.040 68.750 ;
        RECT 20.145 54.060 20.605 54.135 ;
        RECT 25.715 54.060 26.175 54.085 ;
        RECT 20.145 53.620 26.175 54.060 ;
        RECT 20.145 53.565 20.605 53.620 ;
        RECT 25.715 53.515 26.175 53.620 ;
        RECT 22.405 48.870 22.885 48.935 ;
        RECT 22.405 48.550 24.205 48.870 ;
        RECT 22.405 48.385 22.885 48.550 ;
        RECT 23.635 45.710 24.195 48.550 ;
        RECT 27.515 45.710 27.995 45.735 ;
        RECT 23.635 45.290 27.995 45.710 ;
        RECT 23.635 45.280 24.195 45.290 ;
        RECT 27.515 45.185 27.995 45.290 ;
        RECT 20.745 40.120 21.225 40.225 ;
        RECT 24.545 40.120 25.105 40.130 ;
        RECT 20.745 39.700 25.105 40.120 ;
        RECT 20.745 39.675 21.225 39.700 ;
        RECT 24.545 36.860 25.105 39.700 ;
        RECT 25.855 36.860 26.335 37.025 ;
        RECT 24.535 36.540 26.335 36.860 ;
        RECT 25.855 36.475 26.335 36.540 ;
        RECT 22.565 31.790 23.025 31.895 ;
        RECT 28.135 31.790 28.595 31.845 ;
        RECT 22.565 31.350 28.595 31.790 ;
        RECT 22.565 31.325 23.025 31.350 ;
        RECT 28.135 31.275 28.595 31.350 ;
        RECT 29.765 12.265 30.255 73.120 ;
        RECT 38.960 73.080 41.730 74.510 ;
        RECT 31.345 54.070 31.805 54.145 ;
        RECT 36.915 54.070 37.375 54.095 ;
        RECT 31.345 53.630 37.375 54.070 ;
        RECT 31.345 53.575 31.805 53.630 ;
        RECT 36.915 53.525 37.375 53.630 ;
        RECT 33.605 48.880 34.085 48.945 ;
        RECT 33.605 48.560 35.405 48.880 ;
        RECT 33.605 48.395 34.085 48.560 ;
        RECT 34.835 45.720 35.395 48.560 ;
        RECT 38.715 45.720 39.195 45.745 ;
        RECT 34.835 45.300 39.195 45.720 ;
        RECT 34.835 45.290 35.395 45.300 ;
        RECT 38.715 45.195 39.195 45.300 ;
        RECT 32.025 40.120 32.505 40.225 ;
        RECT 35.825 40.120 36.385 40.130 ;
        RECT 32.025 39.700 36.385 40.120 ;
        RECT 32.025 39.675 32.505 39.700 ;
        RECT 35.825 36.860 36.385 39.700 ;
        RECT 37.135 36.860 37.615 37.025 ;
        RECT 35.815 36.540 37.615 36.860 ;
        RECT 37.135 36.475 37.615 36.540 ;
        RECT 33.845 31.790 34.305 31.895 ;
        RECT 39.415 31.790 39.875 31.845 ;
        RECT 33.845 31.350 39.875 31.790 ;
        RECT 33.845 31.325 34.305 31.350 ;
        RECT 39.415 31.275 39.875 31.350 ;
        RECT 41.055 12.360 41.545 73.080 ;
        RECT 49.930 73.030 52.530 74.650 ;
        RECT 61.330 74.530 63.890 75.690 ;
        RECT 73.135 75.580 73.765 80.495 ;
        RECT 84.425 75.690 85.055 81.995 ;
        RECT 72.340 74.980 74.900 75.580 ;
        RECT 42.565 54.040 43.025 54.115 ;
        RECT 48.135 54.040 48.595 54.065 ;
        RECT 42.565 53.600 48.595 54.040 ;
        RECT 42.565 53.545 43.025 53.600 ;
        RECT 48.135 53.495 48.595 53.600 ;
        RECT 44.825 48.850 45.305 48.915 ;
        RECT 44.825 48.530 46.625 48.850 ;
        RECT 44.825 48.365 45.305 48.530 ;
        RECT 46.055 45.690 46.615 48.530 ;
        RECT 49.935 45.690 50.415 45.715 ;
        RECT 46.055 45.270 50.415 45.690 ;
        RECT 46.055 45.260 46.615 45.270 ;
        RECT 49.935 45.165 50.415 45.270 ;
        RECT 43.315 40.100 43.795 40.205 ;
        RECT 47.115 40.100 47.675 40.110 ;
        RECT 43.315 39.680 47.675 40.100 ;
        RECT 43.315 39.655 43.795 39.680 ;
        RECT 47.115 36.840 47.675 39.680 ;
        RECT 48.425 36.840 48.905 37.005 ;
        RECT 47.105 36.520 48.905 36.840 ;
        RECT 48.425 36.455 48.905 36.520 ;
        RECT 45.135 31.770 45.595 31.875 ;
        RECT 50.705 31.770 51.165 31.825 ;
        RECT 45.135 31.330 51.165 31.770 ;
        RECT 45.135 31.305 45.595 31.330 ;
        RECT 50.705 31.255 51.165 31.330 ;
        RECT 41.055 12.350 41.555 12.360 ;
        RECT 28.345 11.115 30.465 12.265 ;
        RECT 41.065 11.965 41.555 12.350 ;
        RECT 51.635 12.145 52.125 73.030 ;
        RECT 61.260 73.010 64.060 74.530 ;
        RECT 72.340 73.050 75.020 74.980 ;
        RECT 83.730 74.540 86.290 75.690 ;
        RECT 95.655 75.580 96.285 83.245 ;
        RECT 106.975 75.640 107.605 84.485 ;
        RECT 118.225 75.650 118.855 85.545 ;
        RECT 129.975 75.650 130.605 86.595 ;
        RECT 133.330 76.605 136.060 77.855 ;
        RECT 137.190 76.585 139.920 77.835 ;
        RECT 53.815 54.020 54.275 54.095 ;
        RECT 59.385 54.020 59.845 54.045 ;
        RECT 53.815 53.580 59.845 54.020 ;
        RECT 53.815 53.525 54.275 53.580 ;
        RECT 59.385 53.475 59.845 53.580 ;
        RECT 56.075 48.830 56.555 48.895 ;
        RECT 56.075 48.510 57.875 48.830 ;
        RECT 56.075 48.345 56.555 48.510 ;
        RECT 57.305 45.670 57.865 48.510 ;
        RECT 61.185 45.670 61.665 45.695 ;
        RECT 57.305 45.250 61.665 45.670 ;
        RECT 57.305 45.240 57.865 45.250 ;
        RECT 61.185 45.145 61.665 45.250 ;
        RECT 54.535 40.100 55.015 40.205 ;
        RECT 58.335 40.100 58.895 40.110 ;
        RECT 54.535 39.680 58.895 40.100 ;
        RECT 54.535 39.655 55.015 39.680 ;
        RECT 58.335 36.840 58.895 39.680 ;
        RECT 59.645 36.840 60.125 37.005 ;
        RECT 58.325 36.520 60.125 36.840 ;
        RECT 59.645 36.455 60.125 36.520 ;
        RECT 56.355 31.770 56.815 31.875 ;
        RECT 61.925 31.770 62.385 31.825 ;
        RECT 56.355 31.330 62.385 31.770 ;
        RECT 56.355 31.305 56.815 31.330 ;
        RECT 61.925 31.255 62.385 31.330 ;
        RECT 29.765 11.100 30.255 11.115 ;
        RECT 39.065 11.005 41.615 11.965 ;
        RECT 50.285 10.995 52.405 12.145 ;
        RECT 62.915 12.135 63.405 73.010 ;
        RECT 65.035 54.010 65.495 54.085 ;
        RECT 70.605 54.010 71.065 54.035 ;
        RECT 65.035 53.570 71.065 54.010 ;
        RECT 65.035 53.515 65.495 53.570 ;
        RECT 70.605 53.465 71.065 53.570 ;
        RECT 67.295 48.820 67.775 48.885 ;
        RECT 67.295 48.500 69.095 48.820 ;
        RECT 67.295 48.335 67.775 48.500 ;
        RECT 68.525 45.660 69.085 48.500 ;
        RECT 72.405 45.660 72.885 45.685 ;
        RECT 68.525 45.240 72.885 45.660 ;
        RECT 68.525 45.230 69.085 45.240 ;
        RECT 72.405 45.135 72.885 45.240 ;
        RECT 65.735 40.100 66.215 40.205 ;
        RECT 69.535 40.100 70.095 40.110 ;
        RECT 65.735 39.680 70.095 40.100 ;
        RECT 65.735 39.655 66.215 39.680 ;
        RECT 69.535 36.840 70.095 39.680 ;
        RECT 70.845 36.840 71.325 37.005 ;
        RECT 69.525 36.520 71.325 36.840 ;
        RECT 70.845 36.455 71.325 36.520 ;
        RECT 67.555 31.770 68.015 31.875 ;
        RECT 73.125 31.770 73.585 31.825 ;
        RECT 67.555 31.330 73.585 31.770 ;
        RECT 67.555 31.305 68.015 31.330 ;
        RECT 73.125 31.255 73.585 31.330 ;
        RECT 74.055 12.165 74.545 73.050 ;
        RECT 83.690 73.000 86.290 74.540 ;
        RECT 94.960 74.710 97.520 75.580 ;
        RECT 94.960 73.020 97.570 74.710 ;
        RECT 106.340 74.460 108.900 75.640 ;
        RECT 117.470 74.720 120.030 75.650 ;
        RECT 76.275 54.000 76.735 54.075 ;
        RECT 81.845 54.000 82.305 54.025 ;
        RECT 76.275 53.560 82.305 54.000 ;
        RECT 76.275 53.505 76.735 53.560 ;
        RECT 81.845 53.455 82.305 53.560 ;
        RECT 78.535 48.810 79.015 48.875 ;
        RECT 78.535 48.490 80.335 48.810 ;
        RECT 78.535 48.325 79.015 48.490 ;
        RECT 79.765 45.650 80.325 48.490 ;
        RECT 83.645 45.650 84.125 45.675 ;
        RECT 79.765 45.230 84.125 45.650 ;
        RECT 79.765 45.220 80.325 45.230 ;
        RECT 83.645 45.125 84.125 45.230 ;
        RECT 77.025 40.090 77.505 40.195 ;
        RECT 80.825 40.090 81.385 40.100 ;
        RECT 77.025 39.670 81.385 40.090 ;
        RECT 77.025 39.645 77.505 39.670 ;
        RECT 80.825 36.830 81.385 39.670 ;
        RECT 82.135 36.830 82.615 36.995 ;
        RECT 80.815 36.510 82.615 36.830 ;
        RECT 82.135 36.445 82.615 36.510 ;
        RECT 78.845 31.760 79.305 31.865 ;
        RECT 84.415 31.760 84.875 31.815 ;
        RECT 78.845 31.320 84.875 31.760 ;
        RECT 78.845 31.295 79.305 31.320 ;
        RECT 84.415 31.245 84.875 31.320 ;
        RECT 61.365 10.985 63.485 12.135 ;
        RECT 72.675 11.015 74.795 12.165 ;
        RECT 85.375 12.155 85.865 73.000 ;
        RECT 87.525 54.010 87.985 54.085 ;
        RECT 93.095 54.010 93.555 54.035 ;
        RECT 87.525 53.570 93.555 54.010 ;
        RECT 87.525 53.515 87.985 53.570 ;
        RECT 93.095 53.465 93.555 53.570 ;
        RECT 89.785 48.820 90.265 48.885 ;
        RECT 89.785 48.500 91.585 48.820 ;
        RECT 89.785 48.335 90.265 48.500 ;
        RECT 91.015 45.660 91.575 48.500 ;
        RECT 94.895 45.660 95.375 45.685 ;
        RECT 91.015 45.240 95.375 45.660 ;
        RECT 91.015 45.230 91.575 45.240 ;
        RECT 94.895 45.135 95.375 45.240 ;
        RECT 88.265 40.110 88.745 40.215 ;
        RECT 92.065 40.110 92.625 40.120 ;
        RECT 88.265 39.690 92.625 40.110 ;
        RECT 88.265 39.665 88.745 39.690 ;
        RECT 92.065 36.850 92.625 39.690 ;
        RECT 93.375 36.850 93.855 37.015 ;
        RECT 92.055 36.530 93.855 36.850 ;
        RECT 93.375 36.465 93.855 36.530 ;
        RECT 90.085 31.780 90.545 31.885 ;
        RECT 95.655 31.780 96.115 31.835 ;
        RECT 90.085 31.340 96.115 31.780 ;
        RECT 90.085 31.315 90.545 31.340 ;
        RECT 95.655 31.265 96.115 31.340 ;
        RECT 96.605 12.155 97.095 73.020 ;
        RECT 106.150 73.000 109.060 74.460 ;
        RECT 117.470 73.070 120.000 74.720 ;
        RECT 129.290 74.650 131.850 75.650 ;
        RECT 129.300 73.140 131.820 74.650 ;
        RECT 98.805 54.000 99.265 54.075 ;
        RECT 104.375 54.000 104.835 54.025 ;
        RECT 98.805 53.560 104.835 54.000 ;
        RECT 98.805 53.505 99.265 53.560 ;
        RECT 104.375 53.455 104.835 53.560 ;
        RECT 101.065 48.810 101.545 48.875 ;
        RECT 101.065 48.490 102.865 48.810 ;
        RECT 101.065 48.325 101.545 48.490 ;
        RECT 102.295 45.650 102.855 48.490 ;
        RECT 106.175 45.650 106.655 45.675 ;
        RECT 102.295 45.230 106.655 45.650 ;
        RECT 102.295 45.220 102.855 45.230 ;
        RECT 106.175 45.125 106.655 45.230 ;
        RECT 99.475 40.130 99.955 40.235 ;
        RECT 103.275 40.130 103.835 40.140 ;
        RECT 99.475 39.710 103.835 40.130 ;
        RECT 99.475 39.685 99.955 39.710 ;
        RECT 103.275 36.870 103.835 39.710 ;
        RECT 104.585 36.870 105.065 37.035 ;
        RECT 103.265 36.550 105.065 36.870 ;
        RECT 104.585 36.485 105.065 36.550 ;
        RECT 101.295 31.800 101.755 31.905 ;
        RECT 106.865 31.800 107.325 31.855 ;
        RECT 101.295 31.360 107.325 31.800 ;
        RECT 101.295 31.335 101.755 31.360 ;
        RECT 106.865 31.285 107.325 31.360 ;
        RECT 107.865 12.205 108.355 73.000 ;
        RECT 110.075 54.000 110.535 54.075 ;
        RECT 115.645 54.000 116.105 54.025 ;
        RECT 110.075 53.560 116.105 54.000 ;
        RECT 110.075 53.505 110.535 53.560 ;
        RECT 115.645 53.455 116.105 53.560 ;
        RECT 112.335 48.810 112.815 48.875 ;
        RECT 112.335 48.490 114.135 48.810 ;
        RECT 112.335 48.325 112.815 48.490 ;
        RECT 113.565 45.650 114.125 48.490 ;
        RECT 117.445 45.650 117.925 45.675 ;
        RECT 113.565 45.230 117.925 45.650 ;
        RECT 113.565 45.220 114.125 45.230 ;
        RECT 117.445 45.125 117.925 45.230 ;
        RECT 110.675 40.170 111.155 40.275 ;
        RECT 114.475 40.170 115.035 40.180 ;
        RECT 110.675 39.750 115.035 40.170 ;
        RECT 110.675 39.725 111.155 39.750 ;
        RECT 114.475 36.910 115.035 39.750 ;
        RECT 115.785 36.910 116.265 37.075 ;
        RECT 114.465 36.590 116.265 36.910 ;
        RECT 115.785 36.525 116.265 36.590 ;
        RECT 112.495 31.840 112.955 31.945 ;
        RECT 118.065 31.840 118.525 31.895 ;
        RECT 112.495 31.400 118.525 31.840 ;
        RECT 112.495 31.375 112.955 31.400 ;
        RECT 118.065 31.325 118.525 31.400 ;
        RECT 119.085 12.205 119.575 73.070 ;
        RECT 121.325 54.000 121.785 54.075 ;
        RECT 126.895 54.000 127.355 54.025 ;
        RECT 121.325 53.560 127.355 54.000 ;
        RECT 121.325 53.505 121.785 53.560 ;
        RECT 126.895 53.455 127.355 53.560 ;
        RECT 123.585 48.810 124.065 48.875 ;
        RECT 123.585 48.490 125.385 48.810 ;
        RECT 123.585 48.325 124.065 48.490 ;
        RECT 124.815 45.650 125.375 48.490 ;
        RECT 128.695 45.650 129.175 45.675 ;
        RECT 124.815 45.230 129.175 45.650 ;
        RECT 124.815 45.220 125.375 45.230 ;
        RECT 128.695 45.125 129.175 45.230 ;
        RECT 121.885 40.190 122.365 40.295 ;
        RECT 125.685 40.190 126.245 40.200 ;
        RECT 121.885 39.770 126.245 40.190 ;
        RECT 121.885 39.745 122.365 39.770 ;
        RECT 125.685 36.930 126.245 39.770 ;
        RECT 126.995 36.930 127.475 37.095 ;
        RECT 125.675 36.610 127.475 36.930 ;
        RECT 126.995 36.545 127.475 36.610 ;
        RECT 123.705 31.860 124.165 31.965 ;
        RECT 129.275 31.860 129.735 31.915 ;
        RECT 123.705 31.420 129.735 31.860 ;
        RECT 123.705 31.395 124.165 31.420 ;
        RECT 129.275 31.345 129.735 31.420 ;
        RECT 130.335 12.235 130.825 73.140 ;
        RECT 74.055 11.010 74.545 11.015 ;
        RECT 83.795 11.005 85.915 12.155 ;
        RECT 95.095 11.005 97.215 12.155 ;
        RECT 106.285 11.055 108.405 12.205 ;
        RECT 117.515 11.055 119.635 12.205 ;
        RECT 128.815 11.085 130.935 12.235 ;
        RECT 107.865 11.010 108.355 11.055 ;
        RECT 119.085 11.050 119.575 11.055 ;
        RECT 85.375 11.000 85.865 11.005 ;
        RECT 96.605 10.980 97.095 11.005 ;
        RECT 74.290 0.135 75.680 1.435 ;
        RECT 93.500 0.205 94.890 1.505 ;
        RECT 112.900 0.335 114.290 1.635 ;
        RECT 131.800 0.405 133.540 1.905 ;
        RECT 151.600 0.275 152.970 1.445 ;
      LAYER met4 ;
        RECT 30.420 225.130 30.670 225.140 ;
        RECT 30.300 224.760 30.670 225.130 ;
        RECT 30.970 224.760 33.430 225.140 ;
        RECT 33.730 224.760 36.190 225.140 ;
        RECT 36.490 224.760 38.950 225.140 ;
        RECT 39.250 224.760 41.710 225.140 ;
        RECT 42.010 224.760 44.470 225.140 ;
        RECT 44.770 224.760 47.230 225.140 ;
        RECT 47.530 224.760 49.990 225.140 ;
        RECT 50.290 224.760 52.750 225.140 ;
        RECT 53.050 224.760 55.510 225.140 ;
        RECT 55.810 224.760 58.270 225.140 ;
        RECT 58.570 224.760 61.030 225.140 ;
        RECT 61.330 224.760 63.790 225.140 ;
        RECT 64.090 224.760 66.550 225.140 ;
        RECT 66.850 224.760 69.310 225.140 ;
        RECT 69.610 224.760 72.070 225.140 ;
        RECT 72.370 224.760 74.830 225.140 ;
        RECT 75.130 224.760 77.590 225.140 ;
        RECT 77.890 224.760 80.350 225.140 ;
        RECT 80.650 224.760 83.110 225.140 ;
        RECT 83.410 224.760 85.870 225.140 ;
        RECT 86.170 224.760 88.630 225.140 ;
        RECT 88.930 224.760 91.390 225.140 ;
        RECT 91.690 224.760 94.150 225.140 ;
        RECT 94.450 224.760 96.910 225.140 ;
        RECT 97.210 224.760 99.670 225.140 ;
        RECT 99.970 224.760 102.430 225.140 ;
        RECT 102.730 224.760 105.190 225.140 ;
        RECT 105.490 224.760 107.950 225.140 ;
        RECT 108.250 224.760 110.710 225.140 ;
        RECT 111.010 224.760 113.470 225.140 ;
        RECT 113.770 224.760 116.230 225.140 ;
        RECT 116.530 224.760 118.990 225.140 ;
        RECT 119.290 224.760 121.750 225.140 ;
        RECT 122.050 224.760 124.510 225.140 ;
        RECT 124.810 224.760 127.270 225.140 ;
        RECT 127.570 224.760 130.030 225.140 ;
        RECT 130.330 224.760 132.790 225.140 ;
        RECT 133.090 224.760 133.520 225.140 ;
        RECT 30.300 224.240 133.520 224.760 ;
        RECT 135.385 224.760 135.550 225.185 ;
        RECT 135.850 224.760 136.745 225.185 ;
        RECT 30.300 219.100 31.660 224.240 ;
        RECT 135.385 223.875 136.745 224.760 ;
        RECT 138.175 224.760 138.310 225.115 ;
        RECT 138.610 224.760 139.535 225.115 ;
        RECT 138.175 223.805 139.535 224.760 ;
        RECT 143.225 224.760 143.830 225.145 ;
        RECT 144.130 224.760 144.585 225.145 ;
        RECT 143.225 223.835 144.585 224.760 ;
        RECT 6.000 218.040 31.660 219.100 ;
        RECT 30.300 217.960 31.660 218.040 ;
        RECT 16.160 159.795 16.490 160.125 ;
        RECT 16.175 158.765 16.475 159.795 ;
        RECT 16.160 158.435 16.490 158.765 ;
        RECT 16.160 115.595 16.490 115.925 ;
        RECT 16.175 114.565 16.475 115.595 ;
        RECT 16.160 114.235 16.490 114.565 ;
        RECT 17.605 100.900 19.205 193.860 ;
        RECT 52.040 178.155 52.370 178.485 ;
        RECT 35.480 173.395 35.810 173.725 ;
        RECT 32.720 169.315 33.050 169.645 ;
        RECT 32.735 115.925 33.035 169.315 ;
        RECT 35.495 124.085 35.795 173.395 ;
        RECT 36.400 169.315 36.730 169.645 ;
        RECT 36.415 124.765 36.715 169.315 ;
        RECT 52.055 138.365 52.355 178.155 ;
        RECT 52.040 138.035 52.370 138.365 ;
        RECT 36.400 124.435 36.730 124.765 ;
        RECT 35.480 123.755 35.810 124.085 ;
        RECT 36.415 117.285 36.715 124.435 ;
        RECT 36.400 116.955 36.730 117.285 ;
        RECT 32.720 115.595 33.050 115.925 ;
        RECT 53.175 100.900 54.775 193.860 ;
        RECT 56.475 100.900 58.075 193.860 ;
        RECT 92.045 100.900 93.645 193.860 ;
        RECT 95.345 100.900 96.945 193.860 ;
        RECT 118.110 97.700 120.130 99.670 ;
        RECT 121.810 97.750 123.830 99.720 ;
        RECT 118.130 93.980 120.130 97.700 ;
        RECT 121.820 96.830 123.820 97.750 ;
        RECT 121.820 94.830 139.410 96.830 ;
        RECT 118.130 91.980 135.580 93.980 ;
        RECT 133.580 77.835 135.580 91.980 ;
        RECT 133.375 76.625 136.015 77.835 ;
        RECT 137.410 77.815 139.410 94.830 ;
        RECT 137.235 76.605 139.875 77.815 ;
        RECT 3.955 71.365 4.000 73.195 ;
        RECT 6.000 71.365 6.055 73.195 ;
        RECT 3.000 68.705 3.025 70.435 ;
        RECT 15.555 68.655 16.995 71.165 ;
        RECT 74.335 1.000 75.635 1.415 ;
        RECT 74.335 0.155 74.530 1.000 ;
        RECT 75.430 0.155 75.635 1.000 ;
        RECT 93.545 1.000 94.845 1.485 ;
        RECT 93.545 0.225 93.850 1.000 ;
        RECT 94.750 0.225 94.845 1.000 ;
        RECT 112.945 1.000 114.245 1.615 ;
        RECT 112.945 0.355 113.170 1.000 ;
        RECT 114.070 0.355 114.245 1.000 ;
        RECT 131.845 1.000 133.495 1.885 ;
        RECT 131.845 0.425 132.490 1.000 ;
        RECT 133.390 0.425 133.495 1.000 ;
        RECT 151.645 1.000 152.925 1.425 ;
        RECT 151.645 0.295 151.810 1.000 ;
        RECT 152.710 0.295 152.925 1.000 ;
  END
END tt_um_08_sws
END LIBRARY

