VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_08_sws
  CLASS BLOCK ;
  FOREIGN tt_um_08_sws ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 200.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNADIFFAREA 394.109192 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 15.155 203.925 15.325 204.115 ;
        RECT 16.995 203.970 17.155 204.080 ;
        RECT 22.515 203.925 22.685 204.115 ;
        RECT 24.355 203.925 24.525 204.115 ;
        RECT 29.875 203.925 30.045 204.115 ;
        RECT 35.395 203.925 35.565 204.115 ;
        RECT 37.235 203.925 37.405 204.115 ;
        RECT 42.755 203.925 42.925 204.115 ;
        RECT 48.275 203.925 48.445 204.115 ;
        RECT 54.255 203.925 54.425 204.115 ;
        RECT 59.775 203.925 59.945 204.115 ;
        RECT 61.155 203.925 61.325 204.115 ;
        RECT 67.135 203.925 67.305 204.115 ;
        RECT 72.655 203.925 72.825 204.115 ;
        RECT 74.035 203.925 74.205 204.115 ;
        RECT 75.875 203.925 76.045 204.115 ;
        RECT 81.395 203.925 81.565 204.115 ;
        RECT 86.915 203.925 87.085 204.115 ;
        RECT 88.755 203.925 88.925 204.115 ;
        RECT 94.275 203.925 94.445 204.115 ;
        RECT 99.795 203.925 99.965 204.115 ;
        RECT 100.770 203.975 100.890 204.085 ;
        RECT 106.235 203.925 106.405 204.115 ;
        RECT 111.755 203.925 111.925 204.115 ;
        RECT 113.135 203.925 113.305 204.115 ;
        RECT 15.015 203.115 16.385 203.925 ;
        RECT 17.315 203.115 22.825 203.925 ;
        RECT 22.845 203.055 23.275 203.840 ;
        RECT 23.295 203.115 24.665 203.925 ;
        RECT 24.675 203.115 30.185 203.925 ;
        RECT 30.195 203.115 35.705 203.925 ;
        RECT 35.725 203.055 36.155 203.840 ;
        RECT 36.175 203.115 37.545 203.925 ;
        RECT 37.555 203.115 43.065 203.925 ;
        RECT 43.075 203.115 48.585 203.925 ;
        RECT 48.605 203.055 49.035 203.840 ;
        RECT 49.055 203.115 54.565 203.925 ;
        RECT 54.575 203.115 60.085 203.925 ;
        RECT 60.095 203.145 61.465 203.925 ;
        RECT 61.485 203.055 61.915 203.840 ;
        RECT 61.935 203.115 67.445 203.925 ;
        RECT 67.455 203.115 72.965 203.925 ;
        RECT 72.985 203.015 74.335 203.925 ;
        RECT 74.365 203.055 74.795 203.840 ;
        RECT 74.815 203.115 76.185 203.925 ;
        RECT 76.195 203.115 81.705 203.925 ;
        RECT 81.715 203.115 87.225 203.925 ;
        RECT 87.245 203.055 87.675 203.840 ;
        RECT 87.695 203.115 89.065 203.925 ;
        RECT 89.075 203.115 94.585 203.925 ;
        RECT 94.595 203.115 100.105 203.925 ;
        RECT 100.125 203.055 100.555 203.840 ;
        RECT 101.035 203.115 106.545 203.925 ;
        RECT 106.555 203.115 112.065 203.925 ;
        RECT 112.075 203.115 113.445 203.925 ;
      LAYER nwell ;
        RECT 14.820 199.895 113.640 202.725 ;
      LAYER pwell ;
        RECT 15.015 198.695 16.385 199.505 ;
        RECT 16.395 198.695 19.145 199.505 ;
        RECT 19.155 198.695 24.665 199.505 ;
        RECT 24.675 198.695 30.185 199.505 ;
        RECT 30.195 198.695 35.705 199.505 ;
        RECT 35.725 198.780 36.155 199.565 ;
        RECT 36.635 198.695 40.305 199.505 ;
        RECT 40.315 198.695 45.825 199.505 ;
        RECT 45.835 198.695 51.345 199.505 ;
        RECT 51.355 199.375 52.275 199.605 ;
        RECT 55.105 199.375 56.035 199.595 ;
        RECT 51.355 198.695 60.545 199.375 ;
        RECT 61.485 198.780 61.915 199.565 ;
        RECT 61.935 198.695 65.045 199.605 ;
        RECT 65.155 199.375 66.075 199.605 ;
        RECT 65.155 198.695 67.445 199.375 ;
        RECT 68.385 198.695 69.735 199.605 ;
        RECT 69.755 199.375 70.675 199.605 ;
        RECT 73.505 199.375 74.435 199.595 ;
        RECT 69.755 198.695 78.945 199.375 ;
        RECT 78.965 198.695 80.315 199.605 ;
        RECT 80.335 198.695 81.705 199.505 ;
        RECT 81.715 198.695 87.225 199.505 ;
        RECT 87.245 198.780 87.675 199.565 ;
        RECT 88.155 198.695 89.985 199.505 ;
        RECT 89.995 198.695 95.505 199.505 ;
        RECT 95.515 198.695 101.025 199.505 ;
        RECT 101.035 198.695 106.545 199.505 ;
        RECT 106.555 198.695 112.065 199.505 ;
        RECT 112.075 198.695 113.445 199.505 ;
        RECT 15.155 198.485 15.325 198.695 ;
        RECT 16.995 198.530 17.155 198.640 ;
        RECT 18.835 198.505 19.005 198.695 ;
        RECT 22.515 198.485 22.685 198.675 ;
        RECT 23.490 198.535 23.610 198.645 ;
        RECT 24.355 198.505 24.525 198.695 ;
        RECT 26.195 198.485 26.365 198.675 ;
        RECT 29.875 198.505 30.045 198.695 ;
        RECT 31.715 198.485 31.885 198.675 ;
        RECT 35.395 198.505 35.565 198.695 ;
        RECT 36.370 198.535 36.490 198.645 ;
        RECT 37.235 198.485 37.405 198.675 ;
        RECT 39.995 198.505 40.165 198.695 ;
        RECT 42.755 198.485 42.925 198.675 ;
        RECT 45.515 198.505 45.685 198.695 ;
        RECT 48.275 198.485 48.445 198.675 ;
        RECT 51.035 198.505 51.205 198.695 ;
        RECT 51.495 198.485 51.665 198.675 ;
        RECT 60.235 198.505 60.405 198.695 ;
        RECT 61.155 198.540 61.315 198.650 ;
        RECT 62.075 198.485 62.245 198.675 ;
        RECT 62.590 198.535 62.710 198.645 ;
        RECT 63.000 198.485 63.170 198.675 ;
        RECT 64.835 198.505 65.005 198.695 ;
        RECT 67.135 198.505 67.305 198.695 ;
        RECT 68.055 198.540 68.215 198.650 ;
        RECT 69.435 198.505 69.605 198.695 ;
        RECT 74.035 198.485 74.205 198.675 ;
        RECT 78.635 198.505 78.805 198.695 ;
        RECT 80.015 198.505 80.185 198.695 ;
        RECT 81.395 198.505 81.565 198.695 ;
        RECT 83.695 198.485 83.865 198.675 ;
        RECT 85.075 198.485 85.245 198.675 ;
        RECT 86.915 198.505 87.085 198.695 ;
        RECT 87.890 198.535 88.010 198.645 ;
        RECT 88.755 198.485 88.925 198.675 ;
        RECT 89.675 198.505 89.845 198.695 ;
        RECT 94.275 198.485 94.445 198.675 ;
        RECT 94.735 198.485 94.905 198.675 ;
        RECT 95.195 198.505 95.365 198.695 ;
        RECT 99.795 198.485 99.965 198.675 ;
        RECT 100.715 198.645 100.885 198.695 ;
        RECT 100.715 198.535 100.890 198.645 ;
        RECT 100.715 198.505 100.885 198.535 ;
        RECT 106.235 198.485 106.405 198.695 ;
        RECT 111.755 198.485 111.925 198.695 ;
        RECT 113.135 198.485 113.305 198.695 ;
        RECT 15.015 197.675 16.385 198.485 ;
        RECT 17.315 197.675 22.825 198.485 ;
        RECT 22.845 197.615 23.275 198.400 ;
        RECT 23.755 197.675 26.505 198.485 ;
        RECT 26.515 197.675 32.025 198.485 ;
        RECT 32.035 197.675 37.545 198.485 ;
        RECT 37.555 197.675 43.065 198.485 ;
        RECT 43.075 197.675 48.585 198.485 ;
        RECT 48.605 197.615 49.035 198.400 ;
        RECT 49.055 197.675 51.805 198.485 ;
        RECT 52.015 197.805 62.385 198.485 ;
        RECT 52.015 197.575 54.225 197.805 ;
        RECT 56.945 197.585 57.875 197.805 ;
        RECT 62.855 197.575 65.145 198.485 ;
        RECT 65.155 197.805 74.345 198.485 ;
        RECT 65.155 197.575 66.075 197.805 ;
        RECT 68.905 197.585 69.835 197.805 ;
        RECT 74.365 197.615 74.795 198.400 ;
        RECT 74.815 197.805 84.005 198.485 ;
        RECT 74.815 197.575 75.735 197.805 ;
        RECT 78.565 197.585 79.495 197.805 ;
        RECT 84.015 197.675 85.385 198.485 ;
        RECT 85.395 197.675 89.065 198.485 ;
        RECT 89.075 197.675 94.585 198.485 ;
        RECT 94.705 197.805 98.170 198.485 ;
        RECT 97.250 197.575 98.170 197.805 ;
        RECT 98.275 197.675 100.105 198.485 ;
        RECT 100.125 197.615 100.555 198.400 ;
        RECT 101.035 197.675 106.545 198.485 ;
        RECT 106.555 197.675 112.065 198.485 ;
        RECT 112.075 197.675 113.445 198.485 ;
      LAYER nwell ;
        RECT 14.820 194.455 113.640 197.285 ;
      LAYER pwell ;
        RECT 15.015 193.255 16.385 194.065 ;
        RECT 16.395 193.255 19.145 194.065 ;
        RECT 19.155 193.255 24.665 194.065 ;
        RECT 24.675 193.255 30.185 194.065 ;
        RECT 30.195 193.255 35.705 194.065 ;
        RECT 35.725 193.340 36.155 194.125 ;
        RECT 37.095 193.255 40.765 194.065 ;
        RECT 40.775 193.255 46.285 194.065 ;
        RECT 46.295 193.255 51.805 194.065 ;
        RECT 51.825 193.255 53.175 194.165 ;
        RECT 53.205 193.255 54.555 194.165 ;
        RECT 54.575 193.965 55.505 194.165 ;
        RECT 56.840 193.965 57.785 194.165 ;
        RECT 54.575 193.485 57.785 193.965 ;
        RECT 60.450 193.935 61.370 194.165 ;
        RECT 54.715 193.285 57.785 193.485 ;
        RECT 15.155 193.045 15.325 193.255 ;
        RECT 16.995 193.090 17.155 193.200 ;
        RECT 18.835 193.065 19.005 193.255 ;
        RECT 22.515 193.045 22.685 193.235 ;
        RECT 24.355 193.065 24.525 193.255 ;
        RECT 24.815 193.045 24.985 193.235 ;
        RECT 29.875 193.065 30.045 193.255 ;
        RECT 30.335 193.045 30.505 193.235 ;
        RECT 35.395 193.065 35.565 193.255 ;
        RECT 35.855 193.045 36.025 193.235 ;
        RECT 36.775 193.100 36.935 193.210 ;
        RECT 40.455 193.065 40.625 193.255 ;
        RECT 41.375 193.045 41.545 193.235 ;
        RECT 41.835 193.045 42.005 193.235 ;
        RECT 45.975 193.065 46.145 193.255 ;
        RECT 46.895 193.045 47.065 193.235 ;
        RECT 48.275 193.045 48.445 193.235 ;
        RECT 49.250 193.095 49.370 193.205 ;
        RECT 51.495 193.065 51.665 193.255 ;
        RECT 52.875 193.065 53.045 193.255 ;
        RECT 53.335 193.065 53.505 193.255 ;
        RECT 54.715 193.045 54.885 193.285 ;
        RECT 56.840 193.255 57.785 193.285 ;
        RECT 57.905 193.255 61.370 193.935 ;
        RECT 61.485 193.340 61.915 194.125 ;
        RECT 62.225 193.255 65.145 194.165 ;
        RECT 67.895 193.935 68.825 194.165 ;
        RECT 70.345 193.935 71.275 194.165 ;
        RECT 74.250 193.935 75.170 194.165 ;
        RECT 65.155 193.255 68.825 193.935 ;
        RECT 69.440 193.255 71.275 193.935 ;
        RECT 71.705 193.255 75.170 193.935 ;
        RECT 75.275 193.255 78.385 194.165 ;
        RECT 78.495 193.255 79.865 194.035 ;
        RECT 79.885 193.255 81.235 194.165 ;
        RECT 82.175 193.255 85.845 194.065 ;
        RECT 85.865 193.255 87.215 194.165 ;
        RECT 87.245 193.340 87.675 194.125 ;
        RECT 90.810 193.935 91.730 194.165 ;
        RECT 88.265 193.255 91.730 193.935 ;
        RECT 91.835 193.255 93.205 194.035 ;
        RECT 93.685 193.255 95.035 194.165 ;
        RECT 95.055 193.935 95.975 194.165 ;
        RECT 98.805 193.935 99.735 194.155 ;
        RECT 95.055 193.255 104.245 193.935 ;
        RECT 104.715 193.255 106.545 194.065 ;
        RECT 106.555 193.255 112.065 194.065 ;
        RECT 112.075 193.255 113.445 194.065 ;
        RECT 57.935 193.065 58.105 193.255 ;
        RECT 60.235 193.045 60.405 193.235 ;
        RECT 62.075 193.045 62.245 193.235 ;
        RECT 15.015 192.235 16.385 193.045 ;
        RECT 17.315 192.235 22.825 193.045 ;
        RECT 22.845 192.175 23.275 192.960 ;
        RECT 23.295 192.235 25.125 193.045 ;
        RECT 25.135 192.235 30.645 193.045 ;
        RECT 30.655 192.235 36.165 193.045 ;
        RECT 36.175 192.235 41.685 193.045 ;
        RECT 41.805 192.365 45.270 193.045 ;
        RECT 44.350 192.135 45.270 192.365 ;
        RECT 45.375 192.235 47.205 193.045 ;
        RECT 47.225 192.135 48.575 193.045 ;
        RECT 48.605 192.175 49.035 192.960 ;
        RECT 49.515 192.235 55.025 193.045 ;
        RECT 55.035 192.235 60.545 193.045 ;
        RECT 60.555 192.365 62.385 193.045 ;
        RECT 62.535 193.015 62.705 193.235 ;
        RECT 64.830 193.065 65.000 193.255 ;
        RECT 65.295 193.065 65.465 193.255 ;
        RECT 69.440 193.235 69.605 193.255 ;
        RECT 65.755 193.045 65.925 193.235 ;
        RECT 69.030 193.095 69.150 193.205 ;
        RECT 69.435 193.065 69.605 193.235 ;
        RECT 70.355 193.045 70.525 193.235 ;
        RECT 71.735 193.065 71.905 193.255 ;
        RECT 73.580 193.045 73.750 193.235 ;
        RECT 74.090 193.095 74.210 193.205 ;
        RECT 75.010 193.095 75.130 193.205 ;
        RECT 75.415 193.045 75.585 193.235 ;
        RECT 78.175 193.065 78.345 193.255 ;
        RECT 78.635 193.045 78.805 193.235 ;
        RECT 79.555 193.065 79.725 193.255 ;
        RECT 80.015 193.065 80.185 193.255 ;
        RECT 81.855 193.100 82.015 193.210 ;
        RECT 84.155 193.045 84.325 193.235 ;
        RECT 84.615 193.045 84.785 193.235 ;
        RECT 85.535 193.065 85.705 193.255 ;
        RECT 85.995 193.065 86.165 193.255 ;
        RECT 87.890 193.095 88.010 193.205 ;
        RECT 88.295 193.065 88.465 193.255 ;
        RECT 91.975 193.065 92.145 193.255 ;
        RECT 93.410 193.095 93.530 193.205 ;
        RECT 93.815 193.065 93.985 193.255 ;
        RECT 94.735 193.045 94.905 193.235 ;
        RECT 95.655 193.090 95.815 193.200 ;
        RECT 99.520 193.045 99.690 193.235 ;
        RECT 103.935 193.065 104.105 193.255 ;
        RECT 104.450 193.095 104.570 193.205 ;
        RECT 106.235 193.065 106.405 193.255 ;
        RECT 109.455 193.045 109.625 193.235 ;
        RECT 109.970 193.095 110.090 193.205 ;
        RECT 111.755 193.045 111.925 193.255 ;
        RECT 113.135 193.045 113.305 193.255 ;
        RECT 64.660 193.015 65.605 193.045 ;
        RECT 62.535 192.815 65.605 193.015 ;
        RECT 60.555 192.135 61.900 192.365 ;
        RECT 62.395 192.335 65.605 192.815 ;
        RECT 65.615 192.815 67.185 193.045 ;
        RECT 69.275 193.005 70.195 193.045 ;
        RECT 69.275 192.815 70.205 193.005 ;
        RECT 65.615 192.455 70.205 192.815 ;
        RECT 65.615 192.365 70.195 192.455 ;
        RECT 70.215 192.365 72.505 193.045 ;
        RECT 62.395 192.135 63.325 192.335 ;
        RECT 64.660 192.135 65.605 192.335 ;
        RECT 67.195 192.135 70.195 192.365 ;
        RECT 71.585 192.135 72.505 192.365 ;
        RECT 72.515 192.135 73.865 193.045 ;
        RECT 74.365 192.175 74.795 192.960 ;
        RECT 75.275 192.365 77.105 193.045 ;
        RECT 77.115 192.235 78.945 193.045 ;
        RECT 78.955 192.235 84.465 193.045 ;
        RECT 84.475 192.265 85.845 193.045 ;
        RECT 85.855 192.365 95.045 193.045 ;
        RECT 96.205 192.365 100.105 193.045 ;
        RECT 85.855 192.135 86.775 192.365 ;
        RECT 89.605 192.145 90.535 192.365 ;
        RECT 99.175 192.135 100.105 192.365 ;
        RECT 100.125 192.175 100.555 192.960 ;
        RECT 100.575 192.365 109.765 193.045 ;
        RECT 100.575 192.135 101.495 192.365 ;
        RECT 104.325 192.145 105.255 192.365 ;
        RECT 110.235 192.235 112.065 193.045 ;
        RECT 112.075 192.235 113.445 193.045 ;
      LAYER nwell ;
        RECT 14.820 189.015 113.640 191.845 ;
      LAYER pwell ;
        RECT 15.015 187.815 16.385 188.625 ;
        RECT 16.395 187.815 17.765 188.625 ;
        RECT 17.775 187.815 23.285 188.625 ;
        RECT 23.295 187.815 28.805 188.625 ;
        RECT 28.815 187.815 34.325 188.625 ;
        RECT 34.345 187.815 35.695 188.725 ;
        RECT 35.725 187.900 36.155 188.685 ;
        RECT 36.635 187.815 38.465 188.625 ;
        RECT 38.475 187.815 39.845 188.595 ;
        RECT 43.055 188.495 43.985 188.725 ;
        RECT 40.085 187.815 43.985 188.495 ;
        RECT 43.995 188.495 44.915 188.725 ;
        RECT 47.745 188.495 48.675 188.715 ;
        RECT 43.995 187.815 53.185 188.495 ;
        RECT 53.195 187.815 54.565 188.625 ;
        RECT 54.575 187.815 55.945 188.595 ;
        RECT 55.955 187.815 61.465 188.625 ;
        RECT 61.485 187.900 61.915 188.685 ;
        RECT 62.855 187.815 66.525 188.625 ;
        RECT 66.535 187.815 68.365 188.495 ;
        RECT 68.375 187.815 72.045 188.625 ;
        RECT 72.055 187.815 77.565 188.625 ;
        RECT 77.945 188.615 78.865 188.725 ;
        RECT 77.945 188.495 80.280 188.615 ;
        RECT 84.945 188.495 85.865 188.715 ;
        RECT 77.945 187.815 87.225 188.495 ;
        RECT 87.245 187.900 87.675 188.685 ;
        RECT 90.895 188.495 91.825 188.725 ;
        RECT 87.925 187.815 91.825 188.495 ;
        RECT 91.835 187.815 93.665 188.625 ;
        RECT 93.770 188.495 94.690 188.725 ;
        RECT 93.770 187.815 97.235 188.495 ;
        RECT 97.815 187.815 99.185 188.595 ;
        RECT 102.395 188.495 103.325 188.725 ;
        RECT 99.425 187.815 103.325 188.495 ;
        RECT 103.430 188.495 104.350 188.725 ;
        RECT 103.430 187.815 106.895 188.495 ;
        RECT 107.025 187.815 108.375 188.725 ;
        RECT 108.395 187.815 109.765 188.595 ;
        RECT 110.235 187.815 112.065 188.625 ;
        RECT 112.075 187.815 113.445 188.625 ;
        RECT 15.155 187.605 15.325 187.815 ;
        RECT 17.455 187.605 17.625 187.815 ;
        RECT 21.135 187.605 21.305 187.795 ;
        RECT 21.595 187.605 21.765 187.795 ;
        RECT 22.975 187.625 23.145 187.815 ;
        RECT 23.435 187.605 23.605 187.795 ;
        RECT 24.815 187.605 24.985 187.795 ;
        RECT 28.495 187.625 28.665 187.815 ;
        RECT 31.900 187.605 32.070 187.795 ;
        RECT 34.015 187.625 34.185 187.815 ;
        RECT 34.475 187.625 34.645 187.815 ;
        RECT 36.370 187.655 36.490 187.765 ;
        RECT 38.155 187.625 38.325 187.815 ;
        RECT 38.615 187.625 38.785 187.815 ;
        RECT 41.835 187.605 42.005 187.795 ;
        RECT 42.755 187.650 42.915 187.760 ;
        RECT 43.215 187.605 43.385 187.795 ;
        RECT 43.400 187.625 43.570 187.815 ;
        RECT 48.000 187.605 48.170 187.795 ;
        RECT 49.250 187.655 49.370 187.765 ;
        RECT 52.875 187.625 53.045 187.815 ;
        RECT 54.255 187.625 54.425 187.815 ;
        RECT 54.715 187.625 54.885 187.815 ;
        RECT 58.395 187.605 58.565 187.795 ;
        RECT 58.910 187.655 59.030 187.765 ;
        RECT 61.155 187.625 61.325 187.815 ;
        RECT 62.535 187.605 62.705 187.795 ;
        RECT 62.995 187.625 63.165 187.795 ;
        RECT 66.215 187.625 66.385 187.815 ;
        RECT 68.055 187.625 68.225 187.815 ;
        RECT 63.095 187.605 63.165 187.625 ;
        RECT 68.515 187.605 68.685 187.795 ;
        RECT 71.735 187.625 71.905 187.815 ;
        RECT 74.035 187.605 74.205 187.795 ;
        RECT 75.875 187.605 76.045 187.795 ;
        RECT 76.335 187.605 76.505 187.795 ;
        RECT 77.255 187.625 77.425 187.815 ;
        RECT 81.120 187.605 81.290 187.795 ;
        RECT 82.775 187.605 82.945 187.795 ;
        RECT 83.290 187.655 83.410 187.765 ;
        RECT 86.915 187.605 87.085 187.815 ;
        RECT 88.295 187.605 88.465 187.795 ;
        RECT 89.215 187.650 89.375 187.760 ;
        RECT 89.675 187.605 89.845 187.795 ;
        RECT 91.240 187.625 91.410 187.815 ;
        RECT 93.355 187.625 93.525 187.815 ;
        RECT 93.630 187.605 93.800 187.795 ;
        RECT 97.035 187.625 97.205 187.815 ;
        RECT 97.550 187.655 97.670 187.765 ;
        RECT 97.955 187.625 98.125 187.815 ;
        RECT 99.795 187.605 99.965 187.795 ;
        RECT 100.715 187.605 100.885 187.795 ;
        RECT 102.740 187.625 102.910 187.815 ;
        RECT 106.695 187.625 106.865 187.815 ;
        RECT 108.075 187.625 108.245 187.815 ;
        RECT 109.455 187.625 109.625 187.815 ;
        RECT 109.970 187.655 110.090 187.765 ;
        RECT 110.835 187.605 111.005 187.795 ;
        RECT 111.755 187.625 111.925 187.815 ;
        RECT 113.135 187.605 113.305 187.815 ;
        RECT 15.015 186.795 16.385 187.605 ;
        RECT 16.395 186.795 17.765 187.605 ;
        RECT 17.775 186.795 21.445 187.605 ;
        RECT 21.465 186.695 22.815 187.605 ;
        RECT 22.845 186.735 23.275 187.520 ;
        RECT 23.295 186.825 24.665 187.605 ;
        RECT 24.785 186.925 28.250 187.605 ;
        RECT 28.585 186.925 32.485 187.605 ;
        RECT 27.330 186.695 28.250 186.925 ;
        RECT 31.555 186.695 32.485 186.925 ;
        RECT 32.865 186.925 42.145 187.605 ;
        RECT 32.865 186.805 35.200 186.925 ;
        RECT 32.865 186.695 33.785 186.805 ;
        RECT 39.865 186.705 40.785 186.925 ;
        RECT 43.075 186.825 44.445 187.605 ;
        RECT 44.685 186.925 48.585 187.605 ;
        RECT 47.655 186.695 48.585 186.925 ;
        RECT 48.605 186.735 49.035 187.520 ;
        RECT 49.515 186.925 58.705 187.605 ;
        RECT 49.515 186.695 50.435 186.925 ;
        RECT 53.265 186.705 54.195 186.925 ;
        RECT 59.175 186.795 62.845 187.605 ;
        RECT 63.095 187.375 65.365 187.605 ;
        RECT 63.095 186.695 65.850 187.375 ;
        RECT 66.075 186.795 68.825 187.605 ;
        RECT 68.835 186.795 74.345 187.605 ;
        RECT 74.365 186.735 74.795 187.520 ;
        RECT 74.815 186.795 76.185 187.605 ;
        RECT 76.205 186.695 77.555 187.605 ;
        RECT 77.805 186.925 81.705 187.605 ;
        RECT 80.775 186.695 81.705 186.925 ;
        RECT 81.715 186.825 83.085 187.605 ;
        RECT 83.650 186.925 87.115 187.605 ;
        RECT 83.650 186.695 84.570 186.925 ;
        RECT 87.245 186.695 88.595 187.605 ;
        RECT 89.645 186.925 93.110 187.605 ;
        RECT 92.190 186.695 93.110 186.925 ;
        RECT 93.215 186.925 97.115 187.605 ;
        RECT 93.215 186.695 94.145 186.925 ;
        RECT 97.355 186.795 100.105 187.605 ;
        RECT 100.125 186.735 100.555 187.520 ;
        RECT 100.585 186.695 101.935 187.605 ;
        RECT 101.955 186.925 111.145 187.605 ;
        RECT 101.955 186.695 102.875 186.925 ;
        RECT 105.705 186.705 106.635 186.925 ;
        RECT 112.075 186.795 113.445 187.605 ;
      LAYER nwell ;
        RECT 14.820 183.575 113.640 186.405 ;
      LAYER pwell ;
        RECT 15.015 182.375 16.385 183.185 ;
        RECT 16.855 182.375 20.525 183.185 ;
        RECT 20.630 183.055 21.550 183.285 ;
        RECT 28.725 183.055 29.655 183.275 ;
        RECT 32.485 183.055 33.405 183.285 ;
        RECT 20.630 182.375 24.095 183.055 ;
        RECT 24.215 182.375 33.405 183.055 ;
        RECT 34.345 182.375 35.695 183.285 ;
        RECT 35.725 182.460 36.155 183.245 ;
        RECT 36.175 182.375 38.005 183.185 ;
        RECT 38.015 182.375 39.385 183.155 ;
        RECT 39.395 183.055 40.325 183.285 ;
        RECT 43.535 183.055 44.455 183.285 ;
        RECT 47.285 183.055 48.215 183.275 ;
        RECT 55.390 183.055 56.310 183.285 ;
        RECT 39.395 182.375 43.295 183.055 ;
        RECT 43.535 182.375 52.725 183.055 ;
        RECT 52.845 182.375 56.310 183.055 ;
        RECT 56.425 182.375 57.775 183.285 ;
        RECT 58.470 182.605 61.225 183.285 ;
        RECT 58.955 182.375 61.225 182.605 ;
        RECT 61.485 182.460 61.915 183.245 ;
        RECT 61.935 182.375 64.685 183.185 ;
        RECT 66.275 183.055 69.275 183.285 ;
        RECT 64.695 182.965 69.275 183.055 ;
        RECT 64.695 182.605 69.285 182.965 ;
        RECT 64.695 182.375 66.265 182.605 ;
        RECT 68.355 182.415 69.285 182.605 ;
        RECT 69.535 182.605 72.290 183.285 ;
        RECT 73.805 183.175 74.725 183.285 ;
        RECT 73.805 183.055 76.140 183.175 ;
        RECT 80.805 183.055 81.725 183.275 ;
        RECT 86.295 183.055 87.225 183.285 ;
        RECT 68.355 182.375 69.275 182.415 ;
        RECT 69.535 182.375 71.805 182.605 ;
        RECT 73.805 182.375 83.085 183.055 ;
        RECT 83.325 182.375 87.225 183.055 ;
        RECT 87.245 182.460 87.675 183.245 ;
        RECT 87.705 182.375 89.055 183.285 ;
        RECT 89.075 183.055 89.995 183.285 ;
        RECT 92.825 183.055 93.755 183.275 ;
        RECT 99.195 183.055 100.115 183.285 ;
        RECT 102.945 183.055 103.875 183.275 ;
        RECT 89.075 182.375 98.265 183.055 ;
        RECT 99.195 182.375 108.385 183.055 ;
        RECT 108.405 182.375 109.755 183.285 ;
        RECT 110.235 182.375 112.065 183.185 ;
        RECT 112.075 182.375 113.445 183.185 ;
        RECT 15.155 182.165 15.325 182.375 ;
        RECT 16.590 182.215 16.710 182.325 ;
        RECT 17.455 182.165 17.625 182.355 ;
        RECT 18.835 182.165 19.005 182.355 ;
        RECT 19.295 182.165 19.465 182.355 ;
        RECT 20.215 182.185 20.385 182.375 ;
        RECT 23.435 182.165 23.605 182.355 ;
        RECT 23.895 182.185 24.065 182.375 ;
        RECT 24.355 182.185 24.525 182.375 ;
        RECT 24.815 182.165 24.985 182.355 ;
        RECT 28.770 182.165 28.940 182.355 ;
        RECT 32.690 182.215 32.810 182.325 ;
        RECT 34.015 182.220 34.175 182.330 ;
        RECT 34.475 182.185 34.645 182.375 ;
        RECT 37.695 182.185 37.865 182.375 ;
        RECT 38.155 182.185 38.325 182.375 ;
        RECT 39.810 182.185 39.980 182.375 ;
        RECT 41.835 182.165 42.005 182.355 ;
        RECT 43.215 182.165 43.385 182.355 ;
        RECT 44.595 182.165 44.765 182.355 ;
        RECT 45.055 182.165 45.225 182.355 ;
        RECT 52.415 182.165 52.585 182.375 ;
        RECT 52.875 182.185 53.045 182.375 ;
        RECT 57.475 182.355 57.645 182.375 ;
        RECT 61.155 182.355 61.225 182.375 ;
        RECT 53.795 182.165 53.965 182.355 ;
        RECT 55.175 182.165 55.345 182.355 ;
        RECT 57.015 182.165 57.185 182.355 ;
        RECT 57.475 182.185 57.650 182.355 ;
        RECT 57.990 182.215 58.110 182.325 ;
        RECT 57.480 182.165 57.650 182.185 ;
        RECT 60.235 182.165 60.405 182.355 ;
        RECT 61.155 182.185 61.325 182.355 ;
        RECT 61.615 182.165 61.785 182.355 ;
        RECT 63.455 182.185 63.625 182.355 ;
        RECT 64.375 182.185 64.545 182.375 ;
        RECT 64.835 182.185 65.005 182.375 ;
        RECT 69.535 182.355 69.605 182.375 ;
        RECT 63.555 182.165 63.625 182.185 ;
        RECT 66.675 182.165 66.845 182.355 ;
        RECT 69.435 182.185 69.605 182.355 ;
        RECT 73.115 182.220 73.275 182.330 ;
        RECT 73.760 182.165 73.930 182.355 ;
        RECT 82.775 182.185 82.945 182.375 ;
        RECT 83.695 182.165 83.865 182.355 ;
        RECT 86.640 182.185 86.810 182.375 ;
        RECT 87.835 182.185 88.005 182.375 ;
        RECT 92.895 182.165 93.065 182.355 ;
        RECT 94.275 182.165 94.445 182.355 ;
        RECT 94.735 182.165 94.905 182.355 ;
        RECT 97.955 182.185 98.125 182.375 ;
        RECT 98.875 182.220 99.035 182.330 ;
        RECT 99.520 182.165 99.690 182.355 ;
        RECT 104.120 182.165 104.290 182.355 ;
        RECT 108.075 182.165 108.245 182.375 ;
        RECT 108.535 182.185 108.705 182.375 ;
        RECT 109.970 182.215 110.090 182.325 ;
        RECT 111.755 182.165 111.925 182.375 ;
        RECT 113.135 182.165 113.305 182.375 ;
        RECT 15.015 181.355 16.385 182.165 ;
        RECT 16.395 181.355 17.765 182.165 ;
        RECT 17.785 181.255 19.135 182.165 ;
        RECT 19.265 181.485 22.730 182.165 ;
        RECT 21.810 181.255 22.730 181.485 ;
        RECT 22.845 181.295 23.275 182.080 ;
        RECT 23.295 181.385 24.665 182.165 ;
        RECT 24.785 181.485 28.250 182.165 ;
        RECT 27.330 181.255 28.250 181.485 ;
        RECT 28.355 181.485 32.255 182.165 ;
        RECT 32.955 181.485 42.145 182.165 ;
        RECT 28.355 181.255 29.285 181.485 ;
        RECT 32.955 181.255 33.875 181.485 ;
        RECT 36.705 181.265 37.635 181.485 ;
        RECT 42.155 181.355 43.525 182.165 ;
        RECT 43.545 181.255 44.895 182.165 ;
        RECT 45.025 181.485 48.490 182.165 ;
        RECT 47.570 181.255 48.490 181.485 ;
        RECT 48.605 181.295 49.035 182.080 ;
        RECT 49.150 181.485 52.615 182.165 ;
        RECT 49.150 181.255 50.070 181.485 ;
        RECT 52.745 181.255 54.095 182.165 ;
        RECT 54.115 181.385 55.485 182.165 ;
        RECT 55.495 181.355 57.325 182.165 ;
        RECT 57.335 181.255 59.945 182.165 ;
        RECT 60.105 181.255 61.455 182.165 ;
        RECT 61.475 181.485 63.305 182.165 ;
        RECT 61.960 181.255 63.305 181.485 ;
        RECT 63.555 181.935 65.825 182.165 ;
        RECT 63.555 181.255 66.310 181.935 ;
        RECT 66.645 181.485 70.110 182.165 ;
        RECT 70.445 181.485 74.345 182.165 ;
        RECT 69.190 181.255 70.110 181.485 ;
        RECT 73.415 181.255 74.345 181.485 ;
        RECT 74.365 181.295 74.795 182.080 ;
        RECT 74.815 181.485 84.005 182.165 ;
        RECT 84.015 181.485 93.205 182.165 ;
        RECT 74.815 181.255 75.735 181.485 ;
        RECT 78.565 181.265 79.495 181.485 ;
        RECT 84.015 181.255 84.935 181.485 ;
        RECT 87.765 181.265 88.695 181.485 ;
        RECT 93.215 181.385 94.585 182.165 ;
        RECT 94.595 181.385 95.965 182.165 ;
        RECT 96.205 181.485 100.105 182.165 ;
        RECT 99.175 181.255 100.105 181.485 ;
        RECT 100.125 181.295 100.555 182.080 ;
        RECT 100.805 181.485 104.705 182.165 ;
        RECT 103.775 181.255 104.705 181.485 ;
        RECT 104.810 181.485 108.275 182.165 ;
        RECT 108.490 181.485 111.955 182.165 ;
        RECT 104.810 181.255 105.730 181.485 ;
        RECT 108.490 181.255 109.410 181.485 ;
        RECT 112.075 181.355 113.445 182.165 ;
      LAYER nwell ;
        RECT 14.820 178.135 113.640 180.965 ;
      LAYER pwell ;
        RECT 15.015 176.935 16.385 177.745 ;
        RECT 16.395 176.935 18.225 177.745 ;
        RECT 20.890 177.615 21.810 177.845 ;
        RECT 18.345 176.935 21.810 177.615 ;
        RECT 21.915 177.615 22.835 177.845 ;
        RECT 25.665 177.615 26.595 177.835 ;
        RECT 31.575 177.615 32.505 177.845 ;
        RECT 21.915 176.935 31.105 177.615 ;
        RECT 31.575 176.935 35.475 177.615 ;
        RECT 35.725 177.020 36.155 177.805 ;
        RECT 36.175 176.935 37.545 177.745 ;
        RECT 37.750 176.935 41.225 177.845 ;
        RECT 41.430 176.935 44.905 177.845 ;
        RECT 44.915 177.615 45.845 177.845 ;
        RECT 52.255 177.615 53.185 177.845 ;
        RECT 56.395 177.615 57.325 177.845 ;
        RECT 44.915 176.935 48.815 177.615 ;
        RECT 49.285 176.935 53.185 177.615 ;
        RECT 53.425 176.935 57.325 177.615 ;
        RECT 57.345 176.935 60.085 177.615 ;
        RECT 60.095 176.935 61.465 177.715 ;
        RECT 61.485 177.020 61.915 177.805 ;
        RECT 61.935 177.615 63.280 177.845 ;
        RECT 64.260 177.615 65.605 177.845 ;
        RECT 61.935 176.935 63.765 177.615 ;
        RECT 63.775 176.935 65.605 177.615 ;
        RECT 65.615 176.935 68.335 177.845 ;
        RECT 68.835 176.935 71.575 177.615 ;
        RECT 71.595 176.935 75.070 177.845 ;
        RECT 75.285 176.935 76.635 177.845 ;
        RECT 79.855 177.615 80.785 177.845 ;
        RECT 76.885 176.935 80.785 177.615 ;
        RECT 80.890 177.615 81.810 177.845 ;
        RECT 80.890 176.935 84.355 177.615 ;
        RECT 84.475 176.935 87.085 177.845 ;
        RECT 87.245 177.020 87.675 177.805 ;
        RECT 88.615 176.935 92.090 177.845 ;
        RECT 92.305 176.935 93.655 177.845 ;
        RECT 93.675 176.935 97.150 177.845 ;
        RECT 97.355 176.935 99.185 177.745 ;
        RECT 99.290 177.615 100.210 177.845 ;
        RECT 99.290 176.935 102.755 177.615 ;
        RECT 102.875 176.935 106.350 177.845 ;
        RECT 106.555 176.935 107.925 177.715 ;
        RECT 107.935 176.935 109.305 177.715 ;
        RECT 109.315 176.935 112.065 177.745 ;
        RECT 112.075 176.935 113.445 177.745 ;
        RECT 15.155 176.725 15.325 176.935 ;
        RECT 17.915 176.745 18.085 176.935 ;
        RECT 18.375 176.745 18.545 176.935 ;
        RECT 18.835 176.725 19.005 176.915 ;
        RECT 19.295 176.725 19.465 176.915 ;
        RECT 24.815 176.725 24.985 176.915 ;
        RECT 25.275 176.725 25.445 176.915 ;
        RECT 30.795 176.745 30.965 176.935 ;
        RECT 31.310 176.775 31.430 176.885 ;
        RECT 31.990 176.745 32.160 176.935 ;
        RECT 35.395 176.725 35.565 176.915 ;
        RECT 36.775 176.725 36.945 176.915 ;
        RECT 37.235 176.885 37.405 176.935 ;
        RECT 37.235 176.775 37.410 176.885 ;
        RECT 37.235 176.745 37.405 176.775 ;
        RECT 40.910 176.725 41.080 176.935 ;
        RECT 41.375 176.725 41.545 176.915 ;
        RECT 44.590 176.745 44.760 176.935 ;
        RECT 45.060 176.725 45.230 176.915 ;
        RECT 45.330 176.745 45.500 176.935 ;
        RECT 52.600 176.745 52.770 176.935 ;
        RECT 56.740 176.745 56.910 176.935 ;
        RECT 57.935 176.725 58.105 176.915 ;
        RECT 58.395 176.725 58.565 176.915 ;
        RECT 59.775 176.745 59.945 176.935 ;
        RECT 61.155 176.745 61.325 176.935 ;
        RECT 62.130 176.775 62.250 176.885 ;
        RECT 62.535 176.725 62.705 176.915 ;
        RECT 63.455 176.745 63.625 176.935 ;
        RECT 63.915 176.745 64.085 176.935 ;
        RECT 65.755 176.725 65.925 176.935 ;
        RECT 66.675 176.770 66.835 176.880 ;
        RECT 67.140 176.725 67.310 176.915 ;
        RECT 68.570 176.775 68.690 176.885 ;
        RECT 68.975 176.745 69.145 176.935 ;
        RECT 70.820 176.725 70.990 176.915 ;
        RECT 71.740 176.745 71.910 176.935 ;
        RECT 74.960 176.725 75.130 176.915 ;
        RECT 76.335 176.745 76.505 176.935 ;
        RECT 78.635 176.725 78.805 176.915 ;
        RECT 80.200 176.745 80.370 176.935 ;
        RECT 82.315 176.725 82.485 176.915 ;
        RECT 84.155 176.745 84.325 176.935 ;
        RECT 84.620 176.745 84.790 176.935 ;
        RECT 88.295 176.780 88.455 176.890 ;
        RECT 88.760 176.745 88.930 176.935 ;
        RECT 92.435 176.725 92.605 176.915 ;
        RECT 93.355 176.745 93.525 176.935 ;
        RECT 93.820 176.725 93.990 176.935 ;
        RECT 98.875 176.745 99.045 176.935 ;
        RECT 99.795 176.725 99.965 176.915 ;
        RECT 102.095 176.725 102.265 176.915 ;
        RECT 102.555 176.745 102.725 176.935 ;
        RECT 103.020 176.745 103.190 176.935 ;
        RECT 107.615 176.745 107.785 176.935 ;
        RECT 108.075 176.745 108.245 176.935 ;
        RECT 111.295 176.725 111.465 176.915 ;
        RECT 111.755 176.885 111.925 176.935 ;
        RECT 111.755 176.775 111.930 176.885 ;
        RECT 111.755 176.745 111.925 176.775 ;
        RECT 113.135 176.725 113.305 176.935 ;
        RECT 15.015 175.915 16.385 176.725 ;
        RECT 16.395 175.915 19.145 176.725 ;
        RECT 19.265 176.045 22.730 176.725 ;
        RECT 21.810 175.815 22.730 176.045 ;
        RECT 22.845 175.855 23.275 176.640 ;
        RECT 23.295 175.915 25.125 176.725 ;
        RECT 25.145 175.815 26.495 176.725 ;
        RECT 26.515 176.045 35.705 176.725 ;
        RECT 26.515 175.815 27.435 176.045 ;
        RECT 30.265 175.825 31.195 176.045 ;
        RECT 35.715 175.945 37.085 176.725 ;
        RECT 37.750 175.815 41.225 176.725 ;
        RECT 41.345 176.045 44.810 176.725 ;
        RECT 43.890 175.815 44.810 176.045 ;
        RECT 44.915 175.815 48.390 176.725 ;
        RECT 48.605 175.855 49.035 176.640 ;
        RECT 49.055 176.045 58.245 176.725 ;
        RECT 58.365 176.045 61.830 176.725 ;
        RECT 62.395 176.045 64.225 176.725 ;
        RECT 49.055 175.815 49.975 176.045 ;
        RECT 52.805 175.825 53.735 176.045 ;
        RECT 60.910 175.815 61.830 176.045 ;
        RECT 62.880 175.815 64.225 176.045 ;
        RECT 64.235 176.045 66.065 176.725 ;
        RECT 64.235 175.815 65.580 176.045 ;
        RECT 66.995 175.815 70.470 176.725 ;
        RECT 70.675 175.815 74.150 176.725 ;
        RECT 74.365 175.855 74.795 176.640 ;
        RECT 74.815 175.815 78.290 176.725 ;
        RECT 78.605 176.045 82.070 176.725 ;
        RECT 82.175 176.045 91.365 176.725 ;
        RECT 81.150 175.815 82.070 176.045 ;
        RECT 86.685 175.825 87.615 176.045 ;
        RECT 90.445 175.815 91.365 176.045 ;
        RECT 91.375 175.945 92.745 176.725 ;
        RECT 93.675 175.815 97.150 176.725 ;
        RECT 97.355 175.915 100.105 176.725 ;
        RECT 100.125 175.855 100.555 176.640 ;
        RECT 100.575 175.915 102.405 176.725 ;
        RECT 102.415 176.045 111.605 176.725 ;
        RECT 102.415 175.815 103.335 176.045 ;
        RECT 106.165 175.825 107.095 176.045 ;
        RECT 112.075 175.915 113.445 176.725 ;
      LAYER nwell ;
        RECT 14.820 172.695 113.640 175.525 ;
      LAYER pwell ;
        RECT 15.015 171.495 16.385 172.305 ;
        RECT 19.050 172.175 19.970 172.405 ;
        RECT 16.505 171.495 19.970 172.175 ;
        RECT 20.075 172.175 20.995 172.405 ;
        RECT 23.825 172.175 24.755 172.395 ;
        RECT 29.275 172.175 30.205 172.405 ;
        RECT 20.075 171.495 29.265 172.175 ;
        RECT 29.275 171.495 33.175 172.175 ;
        RECT 33.875 171.495 35.705 172.305 ;
        RECT 35.725 171.580 36.155 172.365 ;
        RECT 36.185 171.495 37.535 172.405 ;
        RECT 37.555 171.495 41.030 172.405 ;
        RECT 41.235 171.495 44.710 172.405 ;
        RECT 45.110 171.495 48.585 172.405 ;
        RECT 51.250 172.175 52.170 172.405 ;
        RECT 48.705 171.495 52.170 172.175 ;
        RECT 52.275 172.175 53.195 172.405 ;
        RECT 56.025 172.175 56.955 172.395 ;
        RECT 52.275 171.495 61.465 172.175 ;
        RECT 61.485 171.580 61.915 172.365 ;
        RECT 61.935 171.495 63.305 172.275 ;
        RECT 64.235 172.175 65.580 172.405 ;
        RECT 64.235 171.495 66.065 172.175 ;
        RECT 66.535 171.495 72.045 172.305 ;
        RECT 73.415 172.175 74.335 172.395 ;
        RECT 80.415 172.295 81.335 172.405 ;
        RECT 79.000 172.175 81.335 172.295 ;
        RECT 72.055 171.495 81.335 172.175 ;
        RECT 81.725 171.495 83.075 172.405 ;
        RECT 86.295 172.175 87.225 172.405 ;
        RECT 83.325 171.495 87.225 172.175 ;
        RECT 87.245 171.580 87.675 172.365 ;
        RECT 87.790 172.175 88.710 172.405 ;
        RECT 87.790 171.495 91.255 172.175 ;
        RECT 91.570 171.495 95.045 172.405 ;
        RECT 95.055 171.495 98.530 172.405 ;
        RECT 99.205 171.495 100.555 172.405 ;
        RECT 100.585 171.495 101.935 172.405 ;
        RECT 101.955 172.175 102.875 172.405 ;
        RECT 105.705 172.175 106.635 172.395 ;
        RECT 101.955 171.495 111.145 172.175 ;
        RECT 112.075 171.495 113.445 172.305 ;
        RECT 15.155 171.285 15.325 171.495 ;
        RECT 16.535 171.305 16.705 171.495 ;
        RECT 17.455 171.285 17.625 171.475 ;
        RECT 18.835 171.285 19.005 171.475 ;
        RECT 19.295 171.285 19.465 171.475 ;
        RECT 23.490 171.335 23.610 171.445 ;
        RECT 25.275 171.285 25.445 171.475 ;
        RECT 25.735 171.285 25.905 171.475 ;
        RECT 28.955 171.305 29.125 171.495 ;
        RECT 29.690 171.305 29.860 171.495 ;
        RECT 29.875 171.330 30.035 171.440 ;
        RECT 30.340 171.285 30.510 171.475 ;
        RECT 33.610 171.335 33.730 171.445 ;
        RECT 34.020 171.285 34.190 171.475 ;
        RECT 35.395 171.305 35.565 171.495 ;
        RECT 37.235 171.305 37.405 171.495 ;
        RECT 37.700 171.285 37.870 171.495 ;
        RECT 41.380 171.305 41.550 171.495 ;
        RECT 42.295 171.285 42.465 171.475 ;
        RECT 44.135 171.285 44.305 171.475 ;
        RECT 44.870 171.285 45.040 171.475 ;
        RECT 48.270 171.305 48.440 171.495 ;
        RECT 48.735 171.305 48.905 171.495 ;
        RECT 49.250 171.335 49.370 171.445 ;
        RECT 53.335 171.305 53.505 171.475 ;
        RECT 53.335 171.285 53.480 171.305 ;
        RECT 57.015 171.285 57.185 171.475 ;
        RECT 58.395 171.285 58.565 171.475 ;
        RECT 58.910 171.335 59.030 171.445 ;
        RECT 61.155 171.305 61.325 171.495 ;
        RECT 62.535 171.285 62.705 171.475 ;
        RECT 62.995 171.305 63.165 171.495 ;
        RECT 63.915 171.340 64.075 171.450 ;
        RECT 64.375 171.285 64.545 171.475 ;
        RECT 64.835 171.285 65.005 171.475 ;
        RECT 65.755 171.305 65.925 171.495 ;
        RECT 66.270 171.335 66.390 171.445 ;
        RECT 68.515 171.285 68.685 171.475 ;
        RECT 68.975 171.285 69.145 171.475 ;
        RECT 70.630 171.285 70.800 171.475 ;
        RECT 71.735 171.305 71.905 171.495 ;
        RECT 72.195 171.305 72.365 171.495 ;
        RECT 81.855 171.305 82.025 171.495 ;
        RECT 85.530 171.285 85.700 171.475 ;
        RECT 86.640 171.305 86.810 171.495 ;
        RECT 87.375 171.285 87.545 171.475 ;
        RECT 88.755 171.285 88.925 171.475 ;
        RECT 91.055 171.305 91.225 171.495 ;
        RECT 94.730 171.475 94.900 171.495 ;
        RECT 94.275 171.285 94.445 171.475 ;
        RECT 94.730 171.305 94.905 171.475 ;
        RECT 95.200 171.305 95.370 171.495 ;
        RECT 98.930 171.335 99.050 171.445 ;
        RECT 99.335 171.305 99.505 171.495 ;
        RECT 94.735 171.285 94.905 171.305 ;
        RECT 99.520 171.285 99.690 171.475 ;
        RECT 100.715 171.305 100.885 171.495 ;
        RECT 101.175 171.330 101.335 171.440 ;
        RECT 105.040 171.285 105.210 171.475 ;
        RECT 105.775 171.285 105.945 171.475 ;
        RECT 107.155 171.285 107.325 171.475 ;
        RECT 110.835 171.305 111.005 171.495 ;
        RECT 111.755 171.285 111.925 171.475 ;
        RECT 113.135 171.285 113.305 171.495 ;
        RECT 15.015 170.475 16.385 171.285 ;
        RECT 16.395 170.475 17.765 171.285 ;
        RECT 17.785 170.375 19.135 171.285 ;
        RECT 19.265 170.605 22.730 171.285 ;
        RECT 21.810 170.375 22.730 170.605 ;
        RECT 22.845 170.415 23.275 171.200 ;
        RECT 23.755 170.475 25.585 171.285 ;
        RECT 25.705 170.605 29.170 171.285 ;
        RECT 28.250 170.375 29.170 170.605 ;
        RECT 30.195 170.375 33.670 171.285 ;
        RECT 33.875 170.375 37.350 171.285 ;
        RECT 37.555 170.375 41.030 171.285 ;
        RECT 41.235 170.505 42.605 171.285 ;
        RECT 42.615 170.475 44.445 171.285 ;
        RECT 44.455 170.605 48.355 171.285 ;
        RECT 44.455 170.375 45.385 170.605 ;
        RECT 48.605 170.415 49.035 171.200 ;
        RECT 49.610 170.375 53.480 171.285 ;
        RECT 53.655 170.475 57.325 171.285 ;
        RECT 57.345 170.375 58.695 171.285 ;
        RECT 59.175 170.475 62.845 171.285 ;
        RECT 62.855 170.605 64.685 171.285 ;
        RECT 64.695 170.605 67.435 171.285 ;
        RECT 62.855 170.375 64.200 170.605 ;
        RECT 67.465 170.375 68.815 171.285 ;
        RECT 68.835 170.505 70.205 171.285 ;
        RECT 70.215 170.605 74.115 171.285 ;
        RECT 70.215 170.375 71.145 170.605 ;
        RECT 74.365 170.415 74.795 171.200 ;
        RECT 74.835 170.375 85.845 171.285 ;
        RECT 85.855 170.475 87.685 171.285 ;
        RECT 87.695 170.505 89.065 171.285 ;
        RECT 89.075 170.475 94.585 171.285 ;
        RECT 94.605 170.375 95.955 171.285 ;
        RECT 96.205 170.605 100.105 171.285 ;
        RECT 99.175 170.375 100.105 170.605 ;
        RECT 100.125 170.415 100.555 171.200 ;
        RECT 101.725 170.605 105.625 171.285 ;
        RECT 104.695 170.375 105.625 170.605 ;
        RECT 105.635 170.505 107.005 171.285 ;
        RECT 107.015 170.505 108.385 171.285 ;
        RECT 108.395 170.475 112.065 171.285 ;
        RECT 112.075 170.475 113.445 171.285 ;
      LAYER nwell ;
        RECT 14.820 167.255 113.640 170.085 ;
      LAYER pwell ;
        RECT 15.015 166.055 16.385 166.865 ;
        RECT 17.315 166.735 18.235 166.965 ;
        RECT 21.065 166.735 21.995 166.955 ;
        RECT 26.515 166.735 27.435 166.965 ;
        RECT 30.265 166.735 31.195 166.955 ;
        RECT 17.315 166.055 26.505 166.735 ;
        RECT 26.515 166.055 35.705 166.735 ;
        RECT 35.725 166.140 36.155 166.925 ;
        RECT 42.050 166.735 42.970 166.965 ;
        RECT 36.555 166.055 38.980 166.735 ;
        RECT 39.505 166.055 42.970 166.735 ;
        RECT 43.085 166.055 44.435 166.965 ;
        RECT 44.455 166.055 53.560 166.735 ;
        RECT 53.795 166.055 56.405 166.965 ;
        RECT 56.425 166.055 57.775 166.965 ;
        RECT 58.725 166.055 61.465 166.735 ;
        RECT 61.485 166.140 61.915 166.925 ;
        RECT 61.935 166.055 63.765 166.865 ;
        RECT 63.805 166.055 66.525 166.965 ;
        RECT 66.535 166.055 68.365 166.865 ;
        RECT 68.745 166.855 69.665 166.965 ;
        RECT 68.745 166.735 71.080 166.855 ;
        RECT 75.745 166.735 76.665 166.955 ;
        RECT 68.745 166.055 78.025 166.735 ;
        RECT 78.035 166.055 87.140 166.735 ;
        RECT 87.245 166.140 87.675 166.925 ;
        RECT 87.695 166.055 89.065 166.835 ;
        RECT 89.085 166.055 90.435 166.965 ;
        RECT 90.915 166.055 92.285 166.835 ;
        RECT 92.295 166.735 93.215 166.965 ;
        RECT 96.045 166.735 96.975 166.955 ;
        RECT 104.150 166.735 105.070 166.965 ;
        RECT 92.295 166.055 101.485 166.735 ;
        RECT 101.605 166.055 105.070 166.735 ;
        RECT 105.175 166.055 106.545 166.865 ;
        RECT 106.555 166.055 107.925 166.835 ;
        RECT 107.935 166.055 109.765 166.735 ;
        RECT 110.235 166.055 112.065 166.865 ;
        RECT 112.075 166.055 113.445 166.865 ;
        RECT 15.155 165.845 15.325 166.055 ;
        RECT 16.995 165.890 17.155 166.010 ;
        RECT 18.375 165.845 18.545 166.035 ;
        RECT 22.240 165.845 22.410 166.035 ;
        RECT 23.490 165.895 23.610 166.005 ;
        RECT 23.895 165.845 24.065 166.035 ;
        RECT 26.195 165.845 26.365 166.055 ;
        RECT 26.655 165.845 26.825 166.035 ;
        RECT 35.395 165.865 35.565 166.055 ;
        RECT 39.075 165.845 39.245 166.035 ;
        RECT 39.535 165.865 39.705 166.055 ;
        RECT 44.135 165.865 44.305 166.055 ;
        RECT 44.595 165.865 44.765 166.055 ;
        RECT 48.275 165.845 48.445 166.035 ;
        RECT 49.655 165.890 49.815 166.000 ;
        RECT 56.090 165.865 56.260 166.055 ;
        RECT 56.555 165.865 56.725 166.055 ;
        RECT 58.395 165.900 58.555 166.010 ;
        RECT 58.855 165.845 59.025 166.035 ;
        RECT 61.155 165.865 61.325 166.055 ;
        RECT 61.610 165.845 61.780 166.035 ;
        RECT 63.455 165.865 63.625 166.055 ;
        RECT 64.375 165.845 64.545 166.035 ;
        RECT 66.215 165.865 66.385 166.055 ;
        RECT 68.055 165.865 68.225 166.055 ;
        RECT 69.895 165.845 70.065 166.035 ;
        RECT 73.760 165.845 73.930 166.035 ;
        RECT 74.955 165.845 75.125 166.035 ;
        RECT 76.390 165.895 76.510 166.005 ;
        RECT 77.715 165.845 77.885 166.055 ;
        RECT 78.175 165.865 78.345 166.055 ;
        RECT 79.095 165.845 79.265 166.035 ;
        RECT 88.755 165.845 88.925 166.055 ;
        RECT 89.215 165.865 89.385 166.055 ;
        RECT 90.650 165.895 90.770 166.005 ;
        RECT 91.055 165.865 91.225 166.055 ;
        RECT 98.415 165.845 98.585 166.035 ;
        RECT 98.875 165.845 99.045 166.035 ;
        RECT 100.715 165.845 100.885 166.035 ;
        RECT 101.175 165.865 101.345 166.055 ;
        RECT 101.635 165.865 101.805 166.055 ;
        RECT 106.235 165.865 106.405 166.055 ;
        RECT 106.695 165.865 106.865 166.055 ;
        RECT 109.455 165.865 109.625 166.055 ;
        RECT 109.970 165.895 110.090 166.005 ;
        RECT 110.835 165.845 111.005 166.035 ;
        RECT 111.755 165.865 111.925 166.055 ;
        RECT 113.135 165.845 113.305 166.055 ;
        RECT 15.015 165.035 16.385 165.845 ;
        RECT 17.325 164.935 18.675 165.845 ;
        RECT 18.925 165.165 22.825 165.845 ;
        RECT 21.895 164.935 22.825 165.165 ;
        RECT 22.845 164.975 23.275 165.760 ;
        RECT 23.755 165.065 25.125 165.845 ;
        RECT 25.135 165.065 26.505 165.845 ;
        RECT 26.625 165.165 30.090 165.845 ;
        RECT 30.280 165.165 39.385 165.845 ;
        RECT 39.395 165.165 48.585 165.845 ;
        RECT 29.170 164.935 30.090 165.165 ;
        RECT 39.395 164.935 40.315 165.165 ;
        RECT 43.145 164.945 44.075 165.165 ;
        RECT 48.605 164.975 49.035 165.760 ;
        RECT 49.975 165.165 59.165 165.845 ;
        RECT 49.975 164.935 50.895 165.165 ;
        RECT 53.725 164.945 54.655 165.165 ;
        RECT 59.315 164.935 61.925 165.845 ;
        RECT 61.945 165.165 64.685 165.845 ;
        RECT 64.695 165.035 70.205 165.845 ;
        RECT 70.445 165.165 74.345 165.845 ;
        RECT 73.415 164.935 74.345 165.165 ;
        RECT 74.365 164.975 74.795 165.760 ;
        RECT 74.815 165.065 76.185 165.845 ;
        RECT 76.665 164.935 78.015 165.845 ;
        RECT 78.045 164.935 79.395 165.845 ;
        RECT 79.785 165.165 89.065 165.845 ;
        RECT 89.445 165.165 98.725 165.845 ;
        RECT 79.785 165.045 82.120 165.165 ;
        RECT 79.785 164.935 80.705 165.045 ;
        RECT 86.785 164.945 87.705 165.165 ;
        RECT 89.445 165.045 91.780 165.165 ;
        RECT 89.445 164.935 90.365 165.045 ;
        RECT 96.445 164.945 97.365 165.165 ;
        RECT 98.735 165.065 100.105 165.845 ;
        RECT 100.125 164.975 100.555 165.760 ;
        RECT 100.585 164.935 101.935 165.845 ;
        RECT 101.955 165.165 111.145 165.845 ;
        RECT 101.955 164.935 102.875 165.165 ;
        RECT 105.705 164.945 106.635 165.165 ;
        RECT 112.075 165.035 113.445 165.845 ;
      LAYER nwell ;
        RECT 14.820 161.815 113.640 164.645 ;
      LAYER pwell ;
        RECT 15.015 160.615 16.385 161.425 ;
        RECT 16.765 161.415 17.685 161.525 ;
        RECT 16.765 161.295 19.100 161.415 ;
        RECT 23.765 161.295 24.685 161.515 ;
        RECT 26.055 161.295 26.985 161.525 ;
        RECT 16.765 160.615 26.045 161.295 ;
        RECT 26.055 160.615 29.955 161.295 ;
        RECT 30.205 160.615 31.555 161.525 ;
        RECT 34.775 161.295 35.705 161.525 ;
        RECT 31.805 160.615 35.705 161.295 ;
        RECT 35.725 160.700 36.155 161.485 ;
        RECT 36.635 160.615 39.385 161.425 ;
        RECT 42.595 161.295 43.525 161.525 ;
        RECT 39.625 160.615 43.525 161.295 ;
        RECT 44.455 160.615 45.825 161.395 ;
        RECT 48.490 161.295 49.410 161.525 ;
        RECT 52.715 161.295 53.645 161.525 ;
        RECT 45.945 160.615 49.410 161.295 ;
        RECT 49.745 160.615 53.645 161.295 ;
        RECT 54.575 160.615 55.945 161.395 ;
        RECT 55.955 160.615 57.785 161.425 ;
        RECT 57.795 161.295 59.140 161.525 ;
        RECT 60.120 161.295 61.465 161.525 ;
        RECT 57.795 160.615 59.625 161.295 ;
        RECT 59.635 160.615 61.465 161.295 ;
        RECT 61.485 160.700 61.915 161.485 ;
        RECT 61.935 160.615 63.305 161.425 ;
        RECT 63.800 161.295 65.145 161.525 ;
        RECT 65.640 161.295 66.985 161.525 ;
        RECT 67.480 161.295 68.825 161.525 ;
        RECT 72.035 161.295 72.965 161.525 ;
        RECT 63.315 160.615 65.145 161.295 ;
        RECT 65.155 160.615 66.985 161.295 ;
        RECT 66.995 160.615 68.825 161.295 ;
        RECT 69.065 160.615 72.965 161.295 ;
        RECT 73.345 161.415 74.265 161.525 ;
        RECT 73.345 161.295 75.680 161.415 ;
        RECT 80.345 161.295 81.265 161.515 ;
        RECT 86.295 161.295 87.225 161.525 ;
        RECT 73.345 160.615 82.625 161.295 ;
        RECT 83.325 160.615 87.225 161.295 ;
        RECT 87.245 160.700 87.675 161.485 ;
        RECT 87.790 160.615 91.660 161.525 ;
        RECT 91.835 161.295 92.765 161.525 ;
        RECT 99.175 161.295 100.105 161.525 ;
        RECT 104.235 161.295 105.165 161.525 ;
        RECT 91.835 160.615 95.735 161.295 ;
        RECT 96.205 160.615 100.105 161.295 ;
        RECT 101.265 160.615 105.165 161.295 ;
        RECT 105.270 161.295 106.190 161.525 ;
        RECT 105.270 160.615 108.735 161.295 ;
        RECT 108.855 160.615 111.465 161.525 ;
        RECT 112.075 160.615 113.445 161.425 ;
        RECT 15.155 160.405 15.325 160.615 ;
        RECT 16.995 160.450 17.155 160.560 ;
        RECT 18.375 160.405 18.545 160.595 ;
        RECT 22.240 160.405 22.410 160.595 ;
        RECT 23.435 160.405 23.605 160.595 ;
        RECT 24.870 160.455 24.990 160.565 ;
        RECT 25.735 160.425 25.905 160.615 ;
        RECT 26.470 160.425 26.640 160.615 ;
        RECT 28.495 160.405 28.665 160.595 ;
        RECT 30.335 160.425 30.505 160.615 ;
        RECT 35.120 160.425 35.290 160.615 ;
        RECT 36.370 160.455 36.490 160.565 ;
        RECT 38.155 160.405 38.325 160.595 ;
        RECT 39.075 160.425 39.245 160.615 ;
        RECT 39.535 160.405 39.705 160.595 ;
        RECT 40.915 160.405 41.085 160.595 ;
        RECT 41.380 160.405 41.550 160.595 ;
        RECT 42.940 160.425 43.110 160.615 ;
        RECT 44.135 160.460 44.295 160.570 ;
        RECT 44.595 160.425 44.765 160.615 ;
        RECT 45.975 160.425 46.145 160.615 ;
        RECT 48.270 160.405 48.440 160.595 ;
        RECT 50.115 160.405 50.285 160.595 ;
        RECT 50.575 160.405 50.745 160.595 ;
        RECT 53.060 160.425 53.230 160.615 ;
        RECT 54.255 160.460 54.415 160.570 ;
        RECT 54.715 160.425 54.885 160.615 ;
        RECT 56.550 160.405 56.720 160.595 ;
        RECT 57.475 160.425 57.645 160.615 ;
        RECT 57.935 160.405 58.105 160.595 ;
        RECT 59.315 160.425 59.485 160.615 ;
        RECT 59.775 160.405 59.945 160.615 ;
        RECT 61.615 160.405 61.785 160.595 ;
        RECT 62.130 160.455 62.250 160.565 ;
        RECT 62.995 160.425 63.165 160.615 ;
        RECT 63.455 160.425 63.625 160.615 ;
        RECT 63.915 160.405 64.085 160.595 ;
        RECT 64.835 160.450 64.995 160.560 ;
        RECT 65.295 160.425 65.465 160.615 ;
        RECT 67.135 160.425 67.305 160.615 ;
        RECT 68.510 160.405 68.680 160.595 ;
        RECT 68.980 160.405 69.150 160.595 ;
        RECT 72.380 160.425 72.550 160.615 ;
        RECT 74.035 160.405 74.205 160.595 ;
        RECT 78.175 160.405 78.345 160.595 ;
        RECT 78.635 160.405 78.805 160.595 ;
        RECT 80.070 160.455 80.190 160.565 ;
        RECT 80.475 160.405 80.645 160.595 ;
        RECT 81.855 160.405 82.025 160.595 ;
        RECT 82.315 160.425 82.485 160.615 ;
        RECT 82.830 160.455 82.950 160.565 ;
        RECT 86.640 160.425 86.810 160.615 ;
        RECT 91.515 160.595 91.660 160.615 ;
        RECT 91.055 160.405 91.225 160.595 ;
        RECT 91.515 160.425 91.685 160.595 ;
        RECT 92.250 160.425 92.420 160.615 ;
        RECT 96.115 160.405 96.285 160.595 ;
        RECT 96.580 160.405 96.750 160.595 ;
        RECT 99.520 160.425 99.690 160.615 ;
        RECT 100.720 160.570 100.890 160.595 ;
        RECT 100.715 160.460 100.890 160.570 ;
        RECT 100.720 160.405 100.890 160.460 ;
        RECT 104.580 160.425 104.750 160.615 ;
        RECT 107.615 160.405 107.785 160.595 ;
        RECT 108.535 160.425 108.705 160.615 ;
        RECT 109.000 160.425 109.170 160.615 ;
        RECT 110.370 160.405 110.540 160.595 ;
        RECT 110.835 160.405 111.005 160.595 ;
        RECT 111.810 160.455 111.930 160.565 ;
        RECT 113.135 160.405 113.305 160.615 ;
        RECT 15.015 159.595 16.385 160.405 ;
        RECT 17.325 159.495 18.675 160.405 ;
        RECT 18.925 159.725 22.825 160.405 ;
        RECT 21.895 159.495 22.825 159.725 ;
        RECT 22.845 159.535 23.275 160.320 ;
        RECT 23.295 159.625 24.665 160.405 ;
        RECT 25.135 159.595 28.805 160.405 ;
        RECT 29.185 159.725 38.465 160.405 ;
        RECT 29.185 159.605 31.520 159.725 ;
        RECT 29.185 159.495 30.105 159.605 ;
        RECT 36.185 159.505 37.105 159.725 ;
        RECT 38.475 159.625 39.845 160.405 ;
        RECT 39.855 159.595 41.225 160.405 ;
        RECT 41.235 159.495 44.710 160.405 ;
        RECT 45.110 159.495 48.585 160.405 ;
        RECT 48.605 159.535 49.035 160.320 ;
        RECT 49.055 159.595 50.425 160.405 ;
        RECT 50.545 159.725 54.010 160.405 ;
        RECT 53.090 159.495 54.010 159.725 ;
        RECT 54.255 159.495 56.865 160.405 ;
        RECT 56.885 159.495 58.235 160.405 ;
        RECT 58.255 159.725 60.085 160.405 ;
        RECT 60.095 159.725 61.925 160.405 ;
        RECT 62.395 159.725 64.225 160.405 ;
        RECT 58.255 159.495 59.600 159.725 ;
        RECT 60.095 159.495 61.440 159.725 ;
        RECT 62.395 159.495 63.740 159.725 ;
        RECT 65.350 159.495 68.825 160.405 ;
        RECT 68.835 159.495 72.310 160.405 ;
        RECT 72.515 159.595 74.345 160.405 ;
        RECT 74.365 159.535 74.795 160.320 ;
        RECT 74.815 159.595 78.485 160.405 ;
        RECT 78.495 159.625 79.865 160.405 ;
        RECT 80.345 159.495 81.695 160.405 ;
        RECT 81.715 159.725 90.820 160.405 ;
        RECT 91.025 159.725 94.490 160.405 ;
        RECT 93.570 159.495 94.490 159.725 ;
        RECT 94.595 159.595 96.425 160.405 ;
        RECT 96.435 159.495 99.910 160.405 ;
        RECT 100.125 159.535 100.555 160.320 ;
        RECT 100.575 159.495 104.050 160.405 ;
        RECT 104.350 159.725 107.815 160.405 ;
        RECT 104.350 159.495 105.270 159.725 ;
        RECT 108.075 159.495 110.685 160.405 ;
        RECT 110.705 159.495 112.055 160.405 ;
        RECT 112.075 159.595 113.445 160.405 ;
      LAYER nwell ;
        RECT 14.820 156.375 113.640 159.205 ;
      LAYER pwell ;
        RECT 15.015 155.175 16.385 155.985 ;
        RECT 16.765 155.975 17.685 156.085 ;
        RECT 16.765 155.855 19.100 155.975 ;
        RECT 23.765 155.855 24.685 156.075 ;
        RECT 16.765 155.175 26.045 155.855 ;
        RECT 26.515 155.175 28.345 155.985 ;
        RECT 28.355 155.175 31.830 156.085 ;
        RECT 32.230 155.175 35.705 156.085 ;
        RECT 35.725 155.260 36.155 156.045 ;
        RECT 37.290 155.175 40.765 156.085 ;
        RECT 40.970 155.175 44.445 156.085 ;
        RECT 44.455 155.175 46.285 155.985 ;
        RECT 46.295 155.175 51.805 155.985 ;
        RECT 52.185 155.975 53.105 156.085 ;
        RECT 52.185 155.855 54.520 155.975 ;
        RECT 59.185 155.855 60.105 156.075 ;
        RECT 52.185 155.175 61.465 155.855 ;
        RECT 61.485 155.260 61.915 156.045 ;
        RECT 61.935 155.175 65.145 156.085 ;
        RECT 65.810 155.175 69.285 156.085 ;
        RECT 69.295 155.175 72.770 156.085 ;
        RECT 72.975 155.175 74.345 155.985 ;
        RECT 74.355 155.175 78.025 155.985 ;
        RECT 78.035 155.175 83.545 155.985 ;
        RECT 83.750 155.175 87.225 156.085 ;
        RECT 87.245 155.260 87.675 156.045 ;
        RECT 88.155 155.175 89.985 155.985 ;
        RECT 90.190 155.175 93.665 156.085 ;
        RECT 93.675 155.175 97.150 156.085 ;
        RECT 97.355 155.175 99.185 155.985 ;
        RECT 101.850 155.855 102.770 156.085 ;
        RECT 99.305 155.175 102.770 155.855 ;
        RECT 102.875 155.855 103.795 156.085 ;
        RECT 106.625 155.855 107.555 156.075 ;
        RECT 102.875 155.175 112.065 155.855 ;
        RECT 112.075 155.175 113.445 155.985 ;
        RECT 15.155 154.965 15.325 155.175 ;
        RECT 16.590 155.015 16.710 155.125 ;
        RECT 18.375 154.965 18.545 155.155 ;
        RECT 19.110 154.965 19.280 155.155 ;
        RECT 23.490 155.015 23.610 155.125 ;
        RECT 24.170 154.965 24.340 155.155 ;
        RECT 25.735 154.985 25.905 155.175 ;
        RECT 28.035 155.125 28.205 155.175 ;
        RECT 26.250 155.015 26.370 155.125 ;
        RECT 28.035 155.015 28.210 155.125 ;
        RECT 28.035 154.985 28.205 155.015 ;
        RECT 28.500 154.985 28.670 155.175 ;
        RECT 30.795 154.965 30.965 155.155 ;
        RECT 31.260 154.965 31.430 155.155 ;
        RECT 35.390 154.985 35.560 155.175 ;
        RECT 36.775 155.020 36.935 155.130 ;
        RECT 38.150 154.965 38.320 155.155 ;
        RECT 40.450 154.985 40.620 155.175 ;
        RECT 41.830 154.965 42.000 155.155 ;
        RECT 43.215 154.965 43.385 155.155 ;
        RECT 44.130 154.985 44.300 155.175 ;
        RECT 45.975 154.985 46.145 155.175 ;
        RECT 46.895 154.965 47.065 155.155 ;
        RECT 47.355 154.965 47.525 155.155 ;
        RECT 51.495 154.985 51.665 155.175 ;
        RECT 57.935 154.965 58.105 155.155 ;
        RECT 58.395 154.965 58.565 155.155 ;
        RECT 61.155 154.985 61.325 155.175 ;
        RECT 62.080 154.965 62.250 155.155 ;
        RECT 64.835 154.985 65.005 155.175 ;
        RECT 65.350 155.015 65.470 155.125 ;
        RECT 68.055 154.965 68.225 155.155 ;
        RECT 68.970 154.985 69.140 155.175 ;
        RECT 69.440 154.985 69.610 155.175 ;
        RECT 70.815 154.965 70.985 155.155 ;
        RECT 71.275 154.965 71.445 155.155 ;
        RECT 74.035 154.965 74.205 155.175 ;
        RECT 75.010 155.015 75.130 155.125 ;
        RECT 76.795 154.965 76.965 155.155 ;
        RECT 77.715 154.985 77.885 155.175 ;
        RECT 78.175 154.965 78.345 155.155 ;
        RECT 79.555 154.965 79.725 155.155 ;
        RECT 80.475 155.010 80.635 155.120 ;
        RECT 80.935 154.965 81.105 155.155 ;
        RECT 82.775 155.010 82.935 155.120 ;
        RECT 83.235 154.965 83.405 155.175 ;
        RECT 86.910 154.985 87.080 155.175 ;
        RECT 87.890 155.015 88.010 155.125 ;
        RECT 89.675 154.985 89.845 155.175 ;
        RECT 93.350 154.985 93.520 155.175 ;
        RECT 93.820 154.985 93.990 155.175 ;
        RECT 95.655 154.965 95.825 155.155 ;
        RECT 96.120 154.965 96.290 155.155 ;
        RECT 98.875 154.985 99.045 155.175 ;
        RECT 99.335 154.985 99.505 155.175 ;
        RECT 99.850 155.015 99.970 155.125 ;
        RECT 102.095 154.965 102.265 155.155 ;
        RECT 105.960 154.965 106.130 155.155 ;
        RECT 107.615 154.965 107.785 155.155 ;
        RECT 108.075 154.965 108.245 155.155 ;
        RECT 111.755 154.965 111.925 155.175 ;
        RECT 113.135 154.965 113.305 155.175 ;
        RECT 15.015 154.155 16.385 154.965 ;
        RECT 16.855 154.155 18.685 154.965 ;
        RECT 18.695 154.285 22.595 154.965 ;
        RECT 18.695 154.055 19.625 154.285 ;
        RECT 22.845 154.095 23.275 154.880 ;
        RECT 23.755 154.285 27.655 154.965 ;
        RECT 23.755 154.055 24.685 154.285 ;
        RECT 28.355 154.155 31.105 154.965 ;
        RECT 31.115 154.055 34.590 154.965 ;
        RECT 34.990 154.055 38.465 154.965 ;
        RECT 38.670 154.055 42.145 154.965 ;
        RECT 42.155 154.155 43.525 154.965 ;
        RECT 43.535 154.155 47.205 154.965 ;
        RECT 47.225 154.055 48.575 154.965 ;
        RECT 48.605 154.095 49.035 154.880 ;
        RECT 49.055 154.285 58.245 154.965 ;
        RECT 58.365 154.285 61.830 154.965 ;
        RECT 49.055 154.055 49.975 154.285 ;
        RECT 52.805 154.065 53.735 154.285 ;
        RECT 60.910 154.055 61.830 154.285 ;
        RECT 61.935 154.055 65.410 154.965 ;
        RECT 65.625 154.285 68.365 154.965 ;
        RECT 68.405 154.055 71.125 154.965 ;
        RECT 71.135 154.285 72.965 154.965 ;
        RECT 71.620 154.055 72.965 154.285 ;
        RECT 72.975 154.155 74.345 154.965 ;
        RECT 74.365 154.095 74.795 154.880 ;
        RECT 75.275 154.155 77.105 154.965 ;
        RECT 77.125 154.055 78.475 154.965 ;
        RECT 78.505 154.055 79.855 154.965 ;
        RECT 80.795 154.185 82.165 154.965 ;
        RECT 83.095 154.285 92.285 154.965 ;
        RECT 87.605 154.065 88.535 154.285 ;
        RECT 91.365 154.055 92.285 154.285 ;
        RECT 92.390 154.285 95.855 154.965 ;
        RECT 92.390 154.055 93.310 154.285 ;
        RECT 95.975 154.055 99.450 154.965 ;
        RECT 100.125 154.095 100.555 154.880 ;
        RECT 100.575 154.155 102.405 154.965 ;
        RECT 102.645 154.285 106.545 154.965 ;
        RECT 105.615 154.055 106.545 154.285 ;
        RECT 106.555 154.155 107.925 154.965 ;
        RECT 107.935 154.185 109.305 154.965 ;
        RECT 109.315 154.155 112.065 154.965 ;
        RECT 112.075 154.155 113.445 154.965 ;
      LAYER nwell ;
        RECT 14.820 150.935 113.640 153.765 ;
      LAYER pwell ;
        RECT 15.015 149.735 16.385 150.545 ;
        RECT 17.685 150.535 18.605 150.645 ;
        RECT 17.685 150.415 20.020 150.535 ;
        RECT 24.685 150.415 25.605 150.635 ;
        RECT 27.435 150.445 28.380 150.645 ;
        RECT 17.685 149.735 26.965 150.415 ;
        RECT 27.435 149.765 30.185 150.445 ;
        RECT 33.395 150.415 34.325 150.645 ;
        RECT 27.435 149.735 28.380 149.765 ;
        RECT 15.155 149.525 15.325 149.735 ;
        RECT 16.995 149.580 17.155 149.690 ;
        RECT 17.915 149.525 18.085 149.715 ;
        RECT 18.375 149.525 18.545 149.715 ;
        RECT 19.755 149.525 19.925 149.715 ;
        RECT 22.055 149.525 22.225 149.715 ;
        RECT 22.570 149.575 22.690 149.685 ;
        RECT 23.490 149.575 23.610 149.685 ;
        RECT 23.895 149.525 24.065 149.715 ;
        RECT 26.655 149.545 26.825 149.735 ;
        RECT 27.170 149.575 27.290 149.685 ;
        RECT 29.870 149.545 30.040 149.765 ;
        RECT 30.425 149.735 34.325 150.415 ;
        RECT 34.335 149.735 35.705 150.515 ;
        RECT 35.725 149.820 36.155 150.605 ;
        RECT 36.175 149.735 39.650 150.645 ;
        RECT 40.775 149.735 44.250 150.645 ;
        RECT 47.110 150.415 48.030 150.645 ;
        RECT 51.335 150.415 52.265 150.645 ;
        RECT 44.565 149.735 48.030 150.415 ;
        RECT 48.365 149.735 52.265 150.415 ;
        RECT 52.360 149.735 61.465 150.415 ;
        RECT 61.485 149.820 61.915 150.605 ;
        RECT 61.935 149.735 65.410 150.645 ;
        RECT 68.835 150.445 69.780 150.645 ;
        RECT 66.085 149.735 68.825 150.415 ;
        RECT 68.835 149.765 71.585 150.445 ;
        RECT 68.835 149.735 69.780 149.765 ;
        RECT 33.740 149.545 33.910 149.735 ;
        RECT 34.475 149.525 34.645 149.715 ;
        RECT 35.395 149.545 35.565 149.735 ;
        RECT 35.855 149.525 36.025 149.715 ;
        RECT 36.320 149.545 36.490 149.735 ;
        RECT 15.015 148.715 16.385 149.525 ;
        RECT 16.395 148.715 18.225 149.525 ;
        RECT 18.245 148.615 19.595 149.525 ;
        RECT 19.615 148.745 20.985 149.525 ;
        RECT 21.005 148.615 22.355 149.525 ;
        RECT 22.845 148.655 23.275 149.440 ;
        RECT 23.755 148.745 25.125 149.525 ;
        RECT 25.505 148.845 34.785 149.525 ;
        RECT 25.505 148.725 27.840 148.845 ;
        RECT 25.505 148.615 26.425 148.725 ;
        RECT 32.505 148.625 33.425 148.845 ;
        RECT 34.795 148.715 36.165 149.525 ;
        RECT 36.175 149.495 37.120 149.525 ;
        RECT 38.610 149.495 38.780 149.715 ;
        RECT 40.455 149.580 40.615 149.690 ;
        RECT 40.920 149.545 41.090 149.735 ;
        RECT 38.935 149.495 39.880 149.525 ;
        RECT 41.370 149.495 41.540 149.715 ;
        RECT 41.840 149.495 42.010 149.715 ;
        RECT 44.595 149.545 44.765 149.735 ;
        RECT 48.000 149.525 48.170 149.715 ;
        RECT 50.115 149.525 50.285 149.715 ;
        RECT 51.680 149.545 51.850 149.735 ;
        RECT 55.635 149.525 55.805 149.715 ;
        RECT 56.095 149.525 56.265 149.715 ;
        RECT 58.395 149.525 58.565 149.715 ;
        RECT 61.155 149.545 61.325 149.735 ;
        RECT 62.080 149.545 62.250 149.735 ;
        RECT 65.810 149.575 65.930 149.685 ;
        RECT 68.055 149.525 68.225 149.715 ;
        RECT 68.515 149.525 68.685 149.735 ;
        RECT 70.410 149.575 70.530 149.685 ;
        RECT 70.820 149.525 70.990 149.715 ;
        RECT 71.270 149.545 71.440 149.765 ;
        RECT 71.595 149.735 75.070 150.645 ;
        RECT 75.645 150.535 76.565 150.645 ;
        RECT 75.645 150.415 77.980 150.535 ;
        RECT 82.645 150.415 83.565 150.635 ;
        RECT 75.645 149.735 84.925 150.415 ;
        RECT 85.865 149.735 87.215 150.645 ;
        RECT 87.245 149.820 87.675 150.605 ;
        RECT 88.155 149.735 89.525 150.515 ;
        RECT 89.535 150.445 90.480 150.645 ;
        RECT 92.295 150.445 93.240 150.645 ;
        RECT 89.535 149.765 92.285 150.445 ;
        RECT 92.295 149.765 95.045 150.445 ;
        RECT 89.535 149.735 90.480 149.765 ;
        RECT 71.740 149.545 71.910 149.735 ;
        RECT 75.010 149.575 75.130 149.685 ;
        RECT 78.820 149.525 78.990 149.715 ;
        RECT 79.830 149.525 80.000 149.715 ;
        RECT 84.615 149.545 84.785 149.735 ;
        RECT 85.535 149.580 85.695 149.690 ;
        RECT 85.995 149.545 86.165 149.735 ;
        RECT 87.100 149.525 87.270 149.715 ;
        RECT 87.890 149.575 88.010 149.685 ;
        RECT 89.215 149.545 89.385 149.735 ;
        RECT 91.970 149.545 92.140 149.765 ;
        RECT 92.295 149.735 93.240 149.765 ;
        RECT 93.355 149.525 93.525 149.715 ;
        RECT 94.730 149.545 94.900 149.765 ;
        RECT 95.055 149.735 98.530 150.645 ;
        RECT 98.735 149.735 102.210 150.645 ;
        RECT 106.535 150.415 107.465 150.645 ;
        RECT 103.565 149.735 107.465 150.415 ;
        RECT 108.395 149.735 109.765 150.515 ;
        RECT 110.235 149.735 112.065 150.545 ;
        RECT 112.075 149.735 113.445 150.545 ;
        RECT 95.200 149.545 95.370 149.735 ;
        RECT 43.500 149.495 44.445 149.525 ;
        RECT 36.175 148.815 38.925 149.495 ;
        RECT 38.935 148.815 41.685 149.495 ;
        RECT 41.695 148.815 44.445 149.495 ;
        RECT 44.685 148.845 48.585 149.525 ;
        RECT 36.175 148.615 37.120 148.815 ;
        RECT 38.935 148.615 39.880 148.815 ;
        RECT 43.500 148.615 44.445 148.815 ;
        RECT 47.655 148.615 48.585 148.845 ;
        RECT 48.605 148.655 49.035 149.440 ;
        RECT 49.055 148.715 50.425 149.525 ;
        RECT 50.435 148.715 55.945 149.525 ;
        RECT 55.955 148.745 57.325 149.525 ;
        RECT 57.335 148.715 58.705 149.525 ;
        RECT 59.085 148.845 68.365 149.525 ;
        RECT 68.375 148.845 70.205 149.525 ;
        RECT 59.085 148.725 61.420 148.845 ;
        RECT 59.085 148.615 60.005 148.725 ;
        RECT 66.085 148.625 67.005 148.845 ;
        RECT 68.860 148.615 70.205 148.845 ;
        RECT 70.675 148.615 74.150 149.525 ;
        RECT 74.365 148.655 74.795 149.440 ;
        RECT 75.505 148.845 79.405 149.525 ;
        RECT 78.475 148.615 79.405 148.845 ;
        RECT 79.415 148.845 83.315 149.525 ;
        RECT 83.785 148.845 87.685 149.525 ;
        RECT 79.415 148.615 80.345 148.845 ;
        RECT 86.755 148.615 87.685 148.845 ;
        RECT 88.155 148.715 93.665 149.525 ;
        RECT 93.675 149.495 94.620 149.525 ;
        RECT 96.110 149.495 96.280 149.715 ;
        RECT 96.580 149.525 96.750 149.715 ;
        RECT 98.880 149.545 99.050 149.735 ;
        RECT 100.770 149.575 100.890 149.685 ;
        RECT 101.175 149.525 101.345 149.715 ;
        RECT 103.015 149.580 103.175 149.690 ;
        RECT 106.880 149.545 107.050 149.735 ;
        RECT 108.075 149.580 108.235 149.690 ;
        RECT 108.535 149.545 108.705 149.735 ;
        RECT 109.970 149.575 110.090 149.685 ;
        RECT 111.755 149.525 111.925 149.735 ;
        RECT 113.135 149.525 113.305 149.735 ;
        RECT 93.675 148.815 96.425 149.495 ;
        RECT 93.675 148.615 94.620 148.815 ;
        RECT 96.435 148.615 99.910 149.525 ;
        RECT 100.125 148.655 100.555 149.440 ;
        RECT 101.045 148.615 102.395 149.525 ;
        RECT 102.785 148.845 112.065 149.525 ;
        RECT 102.785 148.725 105.120 148.845 ;
        RECT 102.785 148.615 103.705 148.725 ;
        RECT 109.785 148.625 110.705 148.845 ;
        RECT 112.075 148.715 113.445 149.525 ;
      LAYER nwell ;
        RECT 14.820 145.495 113.640 148.325 ;
      LAYER pwell ;
        RECT 15.015 144.295 16.385 145.105 ;
        RECT 17.315 144.295 22.825 145.105 ;
        RECT 22.835 144.295 28.345 145.105 ;
        RECT 28.365 144.295 29.715 145.205 ;
        RECT 30.195 144.295 35.705 145.105 ;
        RECT 35.725 144.380 36.155 145.165 ;
        RECT 36.175 144.295 38.005 145.105 ;
        RECT 38.015 144.295 41.490 145.205 ;
        RECT 42.065 145.095 42.985 145.205 ;
        RECT 42.065 144.975 44.400 145.095 ;
        RECT 49.065 144.975 49.985 145.195 ;
        RECT 42.065 144.295 51.345 144.975 ;
        RECT 51.355 144.295 52.725 145.075 ;
        RECT 53.655 144.295 57.325 145.105 ;
        RECT 60.535 144.975 61.465 145.205 ;
        RECT 57.565 144.295 61.465 144.975 ;
        RECT 61.485 144.380 61.915 145.165 ;
        RECT 61.945 144.295 63.295 145.205 ;
        RECT 64.720 144.975 66.065 145.205 ;
        RECT 64.235 144.295 66.065 144.975 ;
        RECT 66.075 144.295 67.445 145.075 ;
        RECT 67.455 144.295 69.285 145.105 ;
        RECT 69.295 145.005 70.240 145.205 ;
        RECT 69.295 144.325 72.045 145.005 ;
        RECT 69.295 144.295 70.240 144.325 ;
        RECT 15.155 144.085 15.325 144.295 ;
        RECT 16.995 144.130 17.155 144.250 ;
        RECT 22.515 144.085 22.685 144.295 ;
        RECT 23.435 144.085 23.605 144.275 ;
        RECT 28.035 144.105 28.205 144.295 ;
        RECT 28.495 144.105 28.665 144.295 ;
        RECT 35.395 144.275 35.565 144.295 ;
        RECT 29.875 144.245 30.045 144.275 ;
        RECT 29.875 144.135 30.050 144.245 ;
        RECT 29.875 144.085 30.045 144.135 ;
        RECT 15.015 143.275 16.385 144.085 ;
        RECT 17.315 143.275 22.825 144.085 ;
        RECT 22.845 143.215 23.275 144.000 ;
        RECT 23.305 143.175 24.655 144.085 ;
        RECT 24.675 143.275 30.185 144.085 ;
        RECT 30.195 144.055 31.140 144.085 ;
        RECT 32.630 144.055 32.800 144.275 ;
        RECT 35.390 144.105 35.565 144.275 ;
        RECT 35.910 144.135 36.030 144.245 ;
        RECT 37.695 144.105 37.865 144.295 ;
        RECT 38.160 144.105 38.330 144.295 ;
        RECT 32.955 144.055 33.900 144.085 ;
        RECT 35.390 144.055 35.560 144.105 ;
        RECT 38.615 144.085 38.785 144.275 ;
        RECT 39.075 144.085 39.245 144.275 ;
        RECT 41.835 144.085 42.005 144.275 ;
        RECT 42.295 144.085 42.465 144.275 ;
        RECT 47.080 144.085 47.250 144.275 ;
        RECT 48.275 144.130 48.435 144.240 ;
        RECT 30.195 143.375 32.945 144.055 ;
        RECT 32.955 143.375 35.705 144.055 ;
        RECT 30.195 143.175 31.140 143.375 ;
        RECT 32.955 143.175 33.900 143.375 ;
        RECT 36.175 143.275 38.925 144.085 ;
        RECT 38.945 143.175 40.295 144.085 ;
        RECT 40.315 143.275 42.145 144.085 ;
        RECT 42.165 143.175 43.515 144.085 ;
        RECT 43.765 143.405 47.665 144.085 ;
        RECT 49.200 144.055 49.370 144.275 ;
        RECT 51.035 144.105 51.205 144.295 ;
        RECT 51.960 144.085 52.130 144.275 ;
        RECT 52.415 144.105 52.585 144.295 ;
        RECT 53.335 144.140 53.495 144.250 ;
        RECT 55.640 144.085 55.810 144.275 ;
        RECT 57.015 144.105 57.185 144.295 ;
        RECT 60.880 144.105 61.050 144.295 ;
        RECT 62.075 144.105 62.245 144.295 ;
        RECT 63.915 144.140 64.075 144.250 ;
        RECT 64.375 144.105 64.545 144.295 ;
        RECT 66.215 144.105 66.385 144.295 ;
        RECT 68.515 144.085 68.685 144.275 ;
        RECT 68.975 144.105 69.145 144.295 ;
        RECT 71.730 144.105 71.900 144.325 ;
        RECT 72.055 144.295 73.885 145.105 ;
        RECT 74.265 145.095 75.185 145.205 ;
        RECT 74.265 144.975 76.600 145.095 ;
        RECT 81.265 144.975 82.185 145.195 ;
        RECT 74.265 144.295 83.545 144.975 ;
        RECT 83.555 144.295 87.225 145.105 ;
        RECT 87.245 144.380 87.675 145.165 ;
        RECT 87.695 145.005 88.640 145.205 ;
        RECT 87.695 144.325 90.445 145.005 ;
        RECT 87.695 144.295 88.640 144.325 ;
        RECT 73.575 144.105 73.745 144.295 ;
        RECT 74.035 144.085 74.205 144.275 ;
        RECT 75.415 144.130 75.575 144.240 ;
        RECT 79.095 144.085 79.265 144.275 ;
        RECT 79.555 144.085 79.725 144.275 ;
        RECT 83.235 144.085 83.405 144.295 ;
        RECT 86.915 144.105 87.085 144.295 ;
        RECT 87.100 144.085 87.270 144.275 ;
        RECT 87.890 144.135 88.010 144.245 ;
        RECT 90.130 144.105 90.300 144.325 ;
        RECT 90.455 144.295 91.825 145.105 ;
        RECT 91.835 144.295 97.345 145.105 ;
        RECT 97.355 144.295 100.830 145.205 ;
        RECT 101.035 144.295 102.865 145.105 ;
        RECT 106.075 144.975 107.005 145.205 ;
        RECT 103.105 144.295 107.005 144.975 ;
        RECT 107.025 144.295 108.375 145.205 ;
        RECT 108.395 144.295 112.065 145.105 ;
        RECT 112.075 144.295 113.445 145.105 ;
        RECT 91.515 144.275 91.685 144.295 ;
        RECT 91.510 144.105 91.685 144.275 ;
        RECT 91.510 144.085 91.680 144.105 ;
        RECT 95.380 144.085 95.550 144.275 ;
        RECT 96.120 144.085 96.290 144.275 ;
        RECT 97.035 144.105 97.205 144.295 ;
        RECT 97.500 144.105 97.670 144.295 ;
        RECT 99.850 144.135 99.970 144.245 ;
        RECT 100.770 144.135 100.890 144.245 ;
        RECT 101.175 144.085 101.345 144.275 ;
        RECT 102.555 144.105 102.725 144.295 ;
        RECT 106.420 144.105 106.590 144.295 ;
        RECT 108.075 144.105 108.245 144.295 ;
        RECT 111.755 144.085 111.925 144.295 ;
        RECT 113.135 144.085 113.305 144.295 ;
        RECT 50.860 144.055 51.805 144.085 ;
        RECT 46.735 143.175 47.665 143.405 ;
        RECT 48.605 143.215 49.035 144.000 ;
        RECT 49.055 143.375 51.805 144.055 ;
        RECT 50.860 143.175 51.805 143.375 ;
        RECT 51.815 143.175 55.290 144.085 ;
        RECT 55.495 143.175 58.970 144.085 ;
        RECT 59.545 143.405 68.825 144.085 ;
        RECT 59.545 143.285 61.880 143.405 ;
        RECT 59.545 143.175 60.465 143.285 ;
        RECT 66.545 143.185 67.465 143.405 ;
        RECT 68.835 143.275 74.345 144.085 ;
        RECT 74.365 143.215 74.795 144.000 ;
        RECT 75.735 143.275 79.405 144.085 ;
        RECT 79.415 143.305 80.785 144.085 ;
        RECT 80.795 143.275 83.545 144.085 ;
        RECT 83.785 143.405 87.685 144.085 ;
        RECT 86.755 143.175 87.685 143.405 ;
        RECT 88.350 143.175 91.825 144.085 ;
        RECT 92.065 143.405 95.965 144.085 ;
        RECT 95.035 143.175 95.965 143.405 ;
        RECT 95.975 143.175 99.450 144.085 ;
        RECT 100.125 143.215 100.555 144.000 ;
        RECT 101.045 143.175 102.395 144.085 ;
        RECT 102.785 143.405 112.065 144.085 ;
        RECT 102.785 143.285 105.120 143.405 ;
        RECT 102.785 143.175 103.705 143.285 ;
        RECT 109.785 143.185 110.705 143.405 ;
        RECT 112.075 143.275 113.445 144.085 ;
      LAYER nwell ;
        RECT 14.820 140.055 113.640 142.885 ;
      LAYER pwell ;
        RECT 15.015 138.855 16.385 139.665 ;
        RECT 17.315 138.855 18.685 139.635 ;
        RECT 18.705 138.855 20.055 139.765 ;
        RECT 21.435 139.535 22.355 139.755 ;
        RECT 28.435 139.655 29.355 139.765 ;
        RECT 31.795 139.675 32.745 139.765 ;
        RECT 34.555 139.675 35.505 139.765 ;
        RECT 27.020 139.535 29.355 139.655 ;
        RECT 20.075 138.855 29.355 139.535 ;
        RECT 30.815 138.855 32.745 139.675 ;
        RECT 33.575 138.855 35.505 139.675 ;
        RECT 35.725 138.940 36.155 139.725 ;
        RECT 37.535 139.535 38.455 139.755 ;
        RECT 44.535 139.655 45.455 139.765 ;
        RECT 43.120 139.535 45.455 139.655 ;
        RECT 36.175 138.855 45.455 139.535 ;
        RECT 45.835 138.855 47.205 139.635 ;
        RECT 47.410 138.855 50.885 139.765 ;
        RECT 54.095 139.535 55.025 139.765 ;
        RECT 51.125 138.855 55.025 139.535 ;
        RECT 55.495 138.855 56.865 139.635 ;
        RECT 60.535 139.535 61.465 139.765 ;
        RECT 57.565 138.855 61.465 139.535 ;
        RECT 61.485 138.940 61.915 139.725 ;
        RECT 62.865 138.855 64.215 139.765 ;
        RECT 64.695 138.855 66.065 139.635 ;
        RECT 66.995 138.855 70.665 139.665 ;
        RECT 72.480 139.565 73.425 139.765 ;
        RECT 70.675 138.885 73.425 139.565 ;
        RECT 76.635 139.535 77.565 139.765 ;
        RECT 15.155 138.645 15.325 138.855 ;
        RECT 16.995 138.690 17.155 138.810 ;
        RECT 17.455 138.645 17.625 138.855 ;
        RECT 19.110 138.645 19.280 138.835 ;
        RECT 19.755 138.665 19.925 138.855 ;
        RECT 20.215 138.665 20.385 138.855 ;
        RECT 30.815 138.835 30.965 138.855 ;
        RECT 33.575 138.835 33.725 138.855 ;
        RECT 23.435 138.645 23.605 138.835 ;
        RECT 24.815 138.665 24.985 138.835 ;
        RECT 24.835 138.645 24.985 138.665 ;
        RECT 27.390 138.645 27.560 138.835 ;
        RECT 30.335 138.700 30.495 138.810 ;
        RECT 30.795 138.665 30.965 138.835 ;
        RECT 33.150 138.695 33.270 138.805 ;
        RECT 33.555 138.665 33.725 138.835 ;
        RECT 36.315 138.665 36.485 138.855 ;
        RECT 41.830 138.645 42.000 138.835 ;
        RECT 15.015 137.835 16.385 138.645 ;
        RECT 17.315 137.865 18.685 138.645 ;
        RECT 18.695 137.965 22.595 138.645 ;
        RECT 18.695 137.735 19.625 137.965 ;
        RECT 22.845 137.775 23.275 138.560 ;
        RECT 23.305 137.735 24.655 138.645 ;
        RECT 24.835 137.825 26.765 138.645 ;
        RECT 25.815 137.735 26.765 137.825 ;
        RECT 26.975 137.965 30.875 138.645 ;
        RECT 26.975 137.735 27.905 137.965 ;
        RECT 31.135 137.735 42.145 138.645 ;
        RECT 42.155 138.615 43.100 138.645 ;
        RECT 44.590 138.615 44.760 138.835 ;
        RECT 45.060 138.645 45.230 138.835 ;
        RECT 46.895 138.665 47.065 138.855 ;
        RECT 49.655 138.690 49.815 138.800 ;
        RECT 50.570 138.665 50.740 138.855 ;
        RECT 54.440 138.665 54.610 138.855 ;
        RECT 55.230 138.695 55.350 138.805 ;
        RECT 55.635 138.665 55.805 138.855 ;
        RECT 57.070 138.695 57.190 138.805 ;
        RECT 59.315 138.645 59.485 138.835 ;
        RECT 60.880 138.665 61.050 138.855 ;
        RECT 62.075 138.645 62.245 138.835 ;
        RECT 62.535 138.700 62.695 138.810 ;
        RECT 63.915 138.665 64.085 138.855 ;
        RECT 64.430 138.695 64.550 138.805 ;
        RECT 64.835 138.665 65.005 138.855 ;
        RECT 66.675 138.700 66.835 138.810 ;
        RECT 67.595 138.645 67.765 138.835 ;
        RECT 42.155 137.935 44.905 138.615 ;
        RECT 42.155 137.735 43.100 137.935 ;
        RECT 44.915 137.735 48.390 138.645 ;
        RECT 48.605 137.775 49.035 138.560 ;
        RECT 50.345 137.965 59.625 138.645 ;
        RECT 50.345 137.845 52.680 137.965 ;
        RECT 50.345 137.735 51.265 137.845 ;
        RECT 57.345 137.745 58.265 137.965 ;
        RECT 59.635 137.835 62.385 138.645 ;
        RECT 62.395 137.835 67.905 138.645 ;
        RECT 68.060 138.615 68.230 138.835 ;
        RECT 70.355 138.665 70.525 138.855 ;
        RECT 70.820 138.645 70.990 138.885 ;
        RECT 72.480 138.855 73.425 138.885 ;
        RECT 73.665 138.855 77.565 139.535 ;
        RECT 77.945 139.655 78.865 139.765 ;
        RECT 77.945 139.535 80.280 139.655 ;
        RECT 84.945 139.535 85.865 139.755 ;
        RECT 77.945 138.855 87.225 139.535 ;
        RECT 87.245 138.940 87.675 139.725 ;
        RECT 88.065 139.655 88.985 139.765 ;
        RECT 88.065 139.535 90.400 139.655 ;
        RECT 95.065 139.535 95.985 139.755 ;
        RECT 99.565 139.655 100.485 139.765 ;
        RECT 88.065 138.855 97.345 139.535 ;
        RECT 97.355 138.855 98.725 139.635 ;
        RECT 99.565 139.535 101.900 139.655 ;
        RECT 106.565 139.535 107.485 139.755 ;
        RECT 99.565 138.855 108.845 139.535 ;
        RECT 108.855 138.855 110.225 139.635 ;
        RECT 110.235 138.855 112.065 139.665 ;
        RECT 112.075 138.855 113.445 139.665 ;
        RECT 76.980 138.665 77.150 138.855 ;
        RECT 84.155 138.645 84.325 138.835 ;
        RECT 85.535 138.645 85.705 138.835 ;
        RECT 86.050 138.695 86.170 138.805 ;
        RECT 86.915 138.665 87.085 138.855 ;
        RECT 87.375 138.645 87.545 138.835 ;
        RECT 90.135 138.645 90.305 138.835 ;
        RECT 90.595 138.645 90.765 138.835 ;
        RECT 92.435 138.690 92.595 138.800 ;
        RECT 69.720 138.615 70.665 138.645 ;
        RECT 67.915 137.935 70.665 138.615 ;
        RECT 69.720 137.735 70.665 137.935 ;
        RECT 70.675 137.735 74.150 138.645 ;
        RECT 74.365 137.775 74.795 138.560 ;
        RECT 75.185 137.965 84.465 138.645 ;
        RECT 75.185 137.845 77.520 137.965 ;
        RECT 75.185 137.735 76.105 137.845 ;
        RECT 82.185 137.745 83.105 137.965 ;
        RECT 84.485 137.735 85.835 138.645 ;
        RECT 86.315 137.865 87.685 138.645 ;
        RECT 87.695 137.835 90.445 138.645 ;
        RECT 90.465 137.735 91.815 138.645 ;
        RECT 92.755 138.615 93.700 138.645 ;
        RECT 95.190 138.615 95.360 138.835 ;
        RECT 95.660 138.615 95.830 138.835 ;
        RECT 97.035 138.665 97.205 138.855 ;
        RECT 98.415 138.665 98.585 138.855 ;
        RECT 98.930 138.695 99.050 138.805 ;
        RECT 99.795 138.645 99.965 138.835 ;
        RECT 104.120 138.645 104.290 138.835 ;
        RECT 104.910 138.695 105.030 138.805 ;
        RECT 105.315 138.645 105.485 138.835 ;
        RECT 108.535 138.665 108.705 138.855 ;
        RECT 108.995 138.665 109.165 138.855 ;
        RECT 111.755 138.645 111.925 138.855 ;
        RECT 113.135 138.645 113.305 138.855 ;
        RECT 97.320 138.615 98.265 138.645 ;
        RECT 92.755 137.935 95.505 138.615 ;
        RECT 95.515 137.935 98.265 138.615 ;
        RECT 92.755 137.735 93.700 137.935 ;
        RECT 97.320 137.735 98.265 137.935 ;
        RECT 98.275 137.835 100.105 138.645 ;
        RECT 100.125 137.775 100.555 138.560 ;
        RECT 100.805 137.965 104.705 138.645 ;
        RECT 103.775 137.735 104.705 137.965 ;
        RECT 105.175 137.865 106.545 138.645 ;
        RECT 106.555 137.835 112.065 138.645 ;
        RECT 112.075 137.835 113.445 138.645 ;
      LAYER nwell ;
        RECT 14.820 134.615 113.640 137.445 ;
      LAYER pwell ;
        RECT 15.015 133.415 16.385 134.225 ;
        RECT 16.765 134.215 17.685 134.325 ;
        RECT 16.765 134.095 19.100 134.215 ;
        RECT 23.765 134.095 24.685 134.315 ;
        RECT 26.425 134.215 27.345 134.325 ;
        RECT 26.425 134.095 28.760 134.215 ;
        RECT 33.425 134.095 34.345 134.315 ;
        RECT 16.765 133.415 26.045 134.095 ;
        RECT 26.425 133.415 35.705 134.095 ;
        RECT 35.725 133.500 36.155 134.285 ;
        RECT 36.635 134.125 37.580 134.325 ;
        RECT 39.395 134.125 40.340 134.325 ;
        RECT 36.635 133.445 39.385 134.125 ;
        RECT 39.395 133.445 42.145 134.125 ;
        RECT 36.635 133.415 37.580 133.445 ;
        RECT 15.155 133.205 15.325 133.415 ;
        RECT 16.590 133.255 16.710 133.365 ;
        RECT 18.375 133.205 18.545 133.395 ;
        RECT 22.240 133.205 22.410 133.395 ;
        RECT 23.435 133.205 23.605 133.395 ;
        RECT 25.735 133.225 25.905 133.415 ;
        RECT 35.395 133.225 35.565 133.415 ;
        RECT 36.370 133.255 36.490 133.365 ;
        RECT 39.070 133.225 39.240 133.445 ;
        RECT 39.395 133.415 40.340 133.445 ;
        RECT 41.830 133.395 42.000 133.445 ;
        RECT 42.155 133.415 43.985 134.225 ;
        RECT 43.995 133.415 47.470 134.325 ;
        RECT 47.675 133.415 51.150 134.325 ;
        RECT 51.815 134.095 52.745 134.325 ;
        RECT 51.815 133.415 55.715 134.095 ;
        RECT 55.965 133.415 57.315 134.325 ;
        RECT 57.345 133.415 58.695 134.325 ;
        RECT 58.715 133.415 61.465 134.225 ;
        RECT 61.485 133.500 61.915 134.285 ;
        RECT 69.055 134.235 70.005 134.325 ;
        RECT 61.935 133.415 63.305 134.225 ;
        RECT 63.315 133.415 65.145 134.095 ;
        RECT 65.155 133.415 67.905 134.225 ;
        RECT 68.075 133.415 70.005 134.235 ;
        RECT 70.300 133.415 79.405 134.095 ;
        RECT 79.425 133.415 80.775 134.325 ;
        RECT 80.795 133.415 82.165 134.195 ;
        RECT 82.175 133.415 83.545 134.225 ;
        RECT 83.555 133.415 87.225 134.225 ;
        RECT 87.245 133.500 87.675 134.285 ;
        RECT 98.015 134.235 98.965 134.325 ;
        RECT 87.695 133.415 96.800 134.095 ;
        RECT 98.015 133.415 99.945 134.235 ;
        RECT 101.035 133.415 106.545 134.225 ;
        RECT 106.555 133.415 112.065 134.225 ;
        RECT 112.075 133.415 113.445 134.225 ;
        RECT 41.830 133.225 42.005 133.395 ;
        RECT 42.295 133.225 42.465 133.395 ;
        RECT 43.675 133.225 43.845 133.415 ;
        RECT 44.140 133.225 44.310 133.415 ;
        RECT 46.435 133.225 46.605 133.395 ;
        RECT 47.820 133.225 47.990 133.415 ;
        RECT 41.835 133.205 42.005 133.225 ;
        RECT 42.315 133.205 42.465 133.225 ;
        RECT 46.435 133.205 46.585 133.225 ;
        RECT 48.275 133.205 48.445 133.395 ;
        RECT 49.195 133.205 49.365 133.395 ;
        RECT 50.575 133.205 50.745 133.395 ;
        RECT 51.550 133.255 51.670 133.365 ;
        RECT 52.230 133.225 52.400 133.415 ;
        RECT 57.015 133.225 57.185 133.415 ;
        RECT 57.475 133.225 57.645 133.415 ;
        RECT 61.155 133.225 61.325 133.415 ;
        RECT 62.535 133.205 62.705 133.395 ;
        RECT 62.995 133.225 63.165 133.415 ;
        RECT 63.915 133.205 64.085 133.395 ;
        RECT 64.835 133.225 65.005 133.415 ;
        RECT 66.215 133.225 66.385 133.395 ;
        RECT 67.135 133.250 67.295 133.360 ;
        RECT 67.595 133.225 67.765 133.415 ;
        RECT 68.075 133.395 68.225 133.415 ;
        RECT 68.055 133.225 68.225 133.395 ;
        RECT 69.435 133.225 69.605 133.395 ;
        RECT 70.355 133.250 70.515 133.360 ;
        RECT 66.215 133.205 66.365 133.225 ;
        RECT 69.435 133.205 69.585 133.225 ;
        RECT 70.820 133.205 70.990 133.395 ;
        RECT 75.875 133.205 76.045 133.395 ;
        RECT 79.095 133.205 79.265 133.415 ;
        RECT 80.475 133.225 80.645 133.415 ;
        RECT 80.935 133.225 81.105 133.415 ;
        RECT 81.395 133.225 81.565 133.395 ;
        RECT 81.395 133.205 81.545 133.225 ;
        RECT 83.235 133.205 83.405 133.415 ;
        RECT 86.915 133.225 87.085 133.415 ;
        RECT 87.835 133.225 88.005 133.415 ;
        RECT 99.795 133.395 99.945 133.415 ;
        RECT 92.895 133.205 93.065 133.395 ;
        RECT 94.735 133.205 94.905 133.395 ;
        RECT 97.035 133.225 97.205 133.395 ;
        RECT 97.495 133.365 97.655 133.370 ;
        RECT 97.495 133.260 97.670 133.365 ;
        RECT 97.550 133.255 97.670 133.260 ;
        RECT 99.795 133.225 99.965 133.395 ;
        RECT 97.035 133.205 97.185 133.225 ;
        RECT 99.795 133.205 99.945 133.225 ;
        RECT 100.715 133.205 100.885 133.395 ;
        RECT 106.235 133.225 106.405 133.415 ;
        RECT 111.295 133.205 111.465 133.395 ;
        RECT 111.755 133.365 111.925 133.415 ;
        RECT 111.755 133.255 111.930 133.365 ;
        RECT 111.755 133.225 111.925 133.255 ;
        RECT 113.135 133.205 113.305 133.415 ;
        RECT 15.015 132.395 16.385 133.205 ;
        RECT 16.855 132.395 18.685 133.205 ;
        RECT 18.925 132.525 22.825 133.205 ;
        RECT 21.895 132.295 22.825 132.525 ;
        RECT 22.845 132.335 23.275 133.120 ;
        RECT 23.295 132.525 32.575 133.205 ;
        RECT 33.040 132.525 42.145 133.205 ;
        RECT 24.655 132.305 25.575 132.525 ;
        RECT 30.240 132.405 32.575 132.525 ;
        RECT 31.655 132.295 32.575 132.405 ;
        RECT 42.315 132.385 44.245 133.205 ;
        RECT 43.295 132.295 44.245 132.385 ;
        RECT 44.655 132.385 46.585 133.205 ;
        RECT 46.755 132.395 48.585 133.205 ;
        RECT 44.655 132.295 45.605 132.385 ;
        RECT 48.605 132.335 49.035 133.120 ;
        RECT 49.055 132.425 50.425 133.205 ;
        RECT 50.435 132.525 59.715 133.205 ;
        RECT 60.105 132.525 62.845 133.205 ;
        RECT 51.795 132.305 52.715 132.525 ;
        RECT 57.380 132.405 59.715 132.525 ;
        RECT 58.795 132.295 59.715 132.405 ;
        RECT 62.855 132.395 64.225 133.205 ;
        RECT 64.435 132.385 66.365 133.205 ;
        RECT 67.655 132.385 69.585 133.205 ;
        RECT 64.435 132.295 65.385 132.385 ;
        RECT 67.655 132.295 68.605 132.385 ;
        RECT 70.675 132.295 74.150 133.205 ;
        RECT 74.365 132.335 74.795 133.120 ;
        RECT 74.815 132.425 76.185 133.205 ;
        RECT 76.195 132.295 79.355 133.205 ;
        RECT 79.615 132.385 81.545 133.205 ;
        RECT 81.715 132.395 83.545 133.205 ;
        RECT 83.925 132.525 93.205 133.205 ;
        RECT 83.925 132.405 86.260 132.525 ;
        RECT 79.615 132.295 80.565 132.385 ;
        RECT 83.925 132.295 84.845 132.405 ;
        RECT 90.925 132.305 91.845 132.525 ;
        RECT 93.215 132.395 95.045 133.205 ;
        RECT 95.255 132.385 97.185 133.205 ;
        RECT 98.015 132.385 99.945 133.205 ;
        RECT 95.255 132.295 96.205 132.385 ;
        RECT 98.015 132.295 98.965 132.385 ;
        RECT 100.125 132.335 100.555 133.120 ;
        RECT 100.585 132.295 101.935 133.205 ;
        RECT 102.325 132.525 111.605 133.205 ;
        RECT 102.325 132.405 104.660 132.525 ;
        RECT 102.325 132.295 103.245 132.405 ;
        RECT 109.325 132.305 110.245 132.525 ;
        RECT 112.075 132.395 113.445 133.205 ;
      LAYER nwell ;
        RECT 14.820 129.175 113.640 132.005 ;
      LAYER pwell ;
        RECT 15.015 127.975 16.385 128.785 ;
        RECT 16.765 128.775 17.685 128.885 ;
        RECT 16.765 128.655 19.100 128.775 ;
        RECT 23.765 128.655 24.685 128.875 ;
        RECT 16.765 127.975 26.045 128.655 ;
        RECT 26.055 127.975 27.425 128.755 ;
        RECT 27.905 127.975 29.255 128.885 ;
        RECT 29.475 128.795 30.425 128.885 ;
        RECT 29.475 127.975 31.405 128.795 ;
        RECT 34.775 128.655 35.705 128.885 ;
        RECT 31.805 127.975 35.705 128.655 ;
        RECT 35.725 128.060 36.155 128.845 ;
        RECT 36.175 127.975 37.545 128.755 ;
        RECT 37.555 128.655 38.485 128.885 ;
        RECT 37.555 127.975 41.455 128.655 ;
        RECT 41.695 127.975 43.525 128.785 ;
        RECT 56.395 128.655 57.325 128.885 ;
        RECT 60.535 128.655 61.465 128.885 ;
        RECT 43.535 127.975 52.640 128.655 ;
        RECT 53.425 127.975 57.325 128.655 ;
        RECT 57.565 127.975 61.465 128.655 ;
        RECT 61.485 128.060 61.915 128.845 ;
        RECT 62.855 127.975 64.685 128.655 ;
        RECT 64.695 127.975 67.435 128.655 ;
        RECT 67.455 127.975 68.825 128.785 ;
        RECT 72.035 128.655 72.965 128.885 ;
        RECT 74.335 128.655 75.255 128.875 ;
        RECT 81.335 128.775 82.255 128.885 ;
        RECT 79.920 128.655 82.255 128.775 ;
        RECT 86.295 128.655 87.225 128.885 ;
        RECT 69.065 127.975 72.965 128.655 ;
        RECT 72.975 127.975 82.255 128.655 ;
        RECT 83.325 127.975 87.225 128.655 ;
        RECT 87.245 128.060 87.675 128.845 ;
        RECT 89.295 128.795 90.245 128.885 ;
        RECT 94.355 128.795 95.305 128.885 ;
        RECT 88.315 127.975 90.245 128.795 ;
        RECT 90.455 127.975 91.825 128.755 ;
        RECT 91.835 127.975 93.205 128.785 ;
        RECT 93.375 127.975 95.305 128.795 ;
        RECT 96.635 128.795 97.585 128.885 ;
        RECT 96.635 127.975 98.565 128.795 ;
        RECT 102.855 128.655 103.785 128.885 ;
        RECT 106.995 128.655 107.925 128.885 ;
        RECT 99.885 127.975 103.785 128.655 ;
        RECT 104.025 127.975 107.925 128.655 ;
        RECT 107.935 127.975 109.305 128.755 ;
        RECT 109.315 127.975 112.065 128.785 ;
        RECT 112.075 127.975 113.445 128.785 ;
        RECT 15.155 127.765 15.325 127.975 ;
        RECT 19.755 127.765 19.925 127.955 ;
        RECT 21.135 127.765 21.305 127.955 ;
        RECT 22.515 127.765 22.685 127.955 ;
        RECT 23.895 127.810 24.055 127.920 ;
        RECT 24.630 127.765 24.800 127.955 ;
        RECT 25.735 127.785 25.905 127.975 ;
        RECT 27.115 127.785 27.285 127.975 ;
        RECT 27.630 127.815 27.750 127.925 ;
        RECT 28.035 127.785 28.205 127.975 ;
        RECT 31.255 127.955 31.405 127.975 ;
        RECT 28.550 127.815 28.670 127.925 ;
        RECT 31.255 127.765 31.425 127.955 ;
        RECT 35.120 127.785 35.290 127.975 ;
        RECT 37.235 127.785 37.405 127.975 ;
        RECT 37.970 127.785 38.140 127.975 ;
        RECT 40.915 127.765 41.085 127.955 ;
        RECT 43.215 127.785 43.385 127.975 ;
        RECT 43.675 127.925 43.845 127.975 ;
        RECT 43.675 127.815 43.850 127.925 ;
        RECT 43.675 127.785 43.845 127.815 ;
        RECT 45.975 127.785 46.145 127.955 ;
        RECT 46.435 127.785 46.605 127.955 ;
        RECT 49.250 127.815 49.370 127.925 ;
        RECT 43.215 127.765 43.365 127.785 ;
        RECT 45.975 127.765 46.125 127.785 ;
        RECT 15.015 126.955 16.385 127.765 ;
        RECT 16.395 126.955 20.065 127.765 ;
        RECT 20.085 126.855 21.435 127.765 ;
        RECT 21.455 126.955 22.825 127.765 ;
        RECT 22.845 126.895 23.275 127.680 ;
        RECT 24.215 127.085 28.115 127.765 ;
        RECT 24.215 126.855 25.145 127.085 ;
        RECT 28.815 126.955 31.565 127.765 ;
        RECT 31.945 127.085 41.225 127.765 ;
        RECT 31.945 126.965 34.280 127.085 ;
        RECT 31.945 126.855 32.865 126.965 ;
        RECT 38.945 126.865 39.865 127.085 ;
        RECT 41.435 126.945 43.365 127.765 ;
        RECT 44.195 126.945 46.125 127.765 ;
        RECT 46.455 127.765 46.605 127.785 ;
        RECT 52.415 127.765 52.585 127.955 ;
        RECT 52.930 127.815 53.050 127.925 ;
        RECT 55.175 127.765 55.345 127.955 ;
        RECT 55.635 127.765 55.805 127.955 ;
        RECT 56.740 127.785 56.910 127.975 ;
        RECT 60.880 127.785 61.050 127.975 ;
        RECT 62.535 127.820 62.695 127.930 ;
        RECT 64.375 127.785 64.545 127.975 ;
        RECT 64.835 127.785 65.005 127.975 ;
        RECT 66.215 127.765 66.385 127.955 ;
        RECT 67.595 127.765 67.765 127.955 ;
        RECT 68.515 127.785 68.685 127.975 ;
        RECT 68.975 127.765 69.145 127.955 ;
        RECT 69.710 127.765 69.880 127.955 ;
        RECT 72.380 127.785 72.550 127.975 ;
        RECT 73.115 127.785 73.285 127.975 ;
        RECT 74.035 127.810 74.195 127.920 ;
        RECT 76.795 127.785 76.965 127.955 ;
        RECT 76.795 127.765 76.945 127.785 ;
        RECT 77.255 127.765 77.425 127.955 ;
        RECT 80.935 127.765 81.105 127.955 ;
        RECT 82.830 127.815 82.950 127.925 ;
        RECT 86.455 127.765 86.625 127.955 ;
        RECT 86.640 127.785 86.810 127.975 ;
        RECT 88.315 127.955 88.465 127.975 ;
        RECT 86.915 127.765 87.085 127.955 ;
        RECT 87.890 127.815 88.010 127.925 ;
        RECT 88.295 127.785 88.465 127.955 ;
        RECT 88.755 127.810 88.915 127.920 ;
        RECT 90.595 127.785 90.765 127.975 ;
        RECT 92.620 127.765 92.790 127.955 ;
        RECT 92.895 127.785 93.065 127.975 ;
        RECT 93.375 127.955 93.525 127.975 ;
        RECT 98.415 127.955 98.565 127.975 ;
        RECT 93.355 127.765 93.525 127.955 ;
        RECT 96.115 127.820 96.275 127.930 ;
        RECT 98.140 127.765 98.310 127.955 ;
        RECT 98.415 127.785 98.585 127.955 ;
        RECT 98.875 127.765 99.045 127.955 ;
        RECT 99.335 127.820 99.495 127.930 ;
        RECT 100.715 127.765 100.885 127.955 ;
        RECT 103.200 127.785 103.370 127.975 ;
        RECT 107.340 127.785 107.510 127.975 ;
        RECT 108.075 127.785 108.245 127.975 ;
        RECT 111.295 127.765 111.465 127.955 ;
        RECT 111.755 127.925 111.925 127.975 ;
        RECT 111.755 127.815 111.930 127.925 ;
        RECT 111.755 127.785 111.925 127.815 ;
        RECT 113.135 127.765 113.305 127.975 ;
        RECT 46.455 126.945 48.385 127.765 ;
        RECT 41.435 126.855 42.385 126.945 ;
        RECT 44.195 126.855 45.145 126.945 ;
        RECT 47.435 126.855 48.385 126.945 ;
        RECT 48.605 126.895 49.035 127.680 ;
        RECT 49.515 126.855 52.675 127.765 ;
        RECT 52.735 126.955 55.485 127.765 ;
        RECT 55.495 126.985 56.865 127.765 ;
        RECT 57.245 127.085 66.525 127.765 ;
        RECT 57.245 126.965 59.580 127.085 ;
        RECT 57.245 126.855 58.165 126.965 ;
        RECT 64.245 126.865 65.165 127.085 ;
        RECT 66.535 126.955 67.905 127.765 ;
        RECT 67.915 126.985 69.285 127.765 ;
        RECT 69.295 127.085 73.195 127.765 ;
        RECT 69.295 126.855 70.225 127.085 ;
        RECT 74.365 126.895 74.795 127.680 ;
        RECT 75.015 126.945 76.945 127.765 ;
        RECT 75.015 126.855 75.965 126.945 ;
        RECT 77.125 126.855 78.475 127.765 ;
        RECT 78.495 126.955 81.245 127.765 ;
        RECT 81.255 126.955 86.765 127.765 ;
        RECT 86.785 126.855 88.135 127.765 ;
        RECT 89.305 127.085 93.205 127.765 ;
        RECT 92.275 126.855 93.205 127.085 ;
        RECT 93.225 126.855 94.575 127.765 ;
        RECT 94.825 127.085 98.725 127.765 ;
        RECT 97.795 126.855 98.725 127.085 ;
        RECT 98.745 126.855 100.095 127.765 ;
        RECT 100.125 126.895 100.555 127.680 ;
        RECT 100.585 126.855 101.935 127.765 ;
        RECT 102.325 127.085 111.605 127.765 ;
        RECT 102.325 126.965 104.660 127.085 ;
        RECT 102.325 126.855 103.245 126.965 ;
        RECT 109.325 126.865 110.245 127.085 ;
        RECT 112.075 126.955 113.445 127.765 ;
      LAYER nwell ;
        RECT 14.820 123.735 113.640 126.565 ;
      LAYER pwell ;
        RECT 15.015 122.535 16.385 123.345 ;
        RECT 16.855 122.535 18.685 123.345 ;
        RECT 18.705 122.535 20.055 123.445 ;
        RECT 20.445 123.335 21.365 123.445 ;
        RECT 20.445 123.215 22.780 123.335 ;
        RECT 27.445 123.215 28.365 123.435 ;
        RECT 33.395 123.215 34.325 123.445 ;
        RECT 20.445 122.535 29.725 123.215 ;
        RECT 30.425 122.535 34.325 123.215 ;
        RECT 34.335 122.535 35.705 123.345 ;
        RECT 35.725 122.620 36.155 123.405 ;
        RECT 40.535 123.355 41.485 123.445 ;
        RECT 36.175 122.535 38.005 123.345 ;
        RECT 38.015 122.535 39.385 123.315 ;
        RECT 39.555 122.535 41.485 123.355 ;
        RECT 41.695 123.215 42.625 123.445 ;
        RECT 49.035 123.215 49.965 123.445 ;
        RECT 41.695 122.535 45.595 123.215 ;
        RECT 46.065 122.535 49.965 123.215 ;
        RECT 49.975 122.535 51.805 123.345 ;
        RECT 52.185 123.335 53.105 123.445 ;
        RECT 52.185 123.215 54.520 123.335 ;
        RECT 59.185 123.215 60.105 123.435 ;
        RECT 52.185 122.535 61.465 123.215 ;
        RECT 61.485 122.620 61.915 123.405 ;
        RECT 61.945 122.535 63.295 123.445 ;
        RECT 63.315 122.535 64.685 123.315 ;
        RECT 64.695 122.535 66.525 123.345 ;
        RECT 66.545 122.535 67.895 123.445 ;
        RECT 68.285 123.335 69.205 123.445 ;
        RECT 68.285 123.215 70.620 123.335 ;
        RECT 75.285 123.215 76.205 123.435 ;
        RECT 68.285 122.535 77.565 123.215 ;
        RECT 77.575 122.535 81.245 123.345 ;
        RECT 84.455 123.215 85.385 123.445 ;
        RECT 81.485 122.535 85.385 123.215 ;
        RECT 85.395 122.535 87.225 123.345 ;
        RECT 87.245 122.620 87.675 123.405 ;
        RECT 87.695 122.535 90.445 123.345 ;
        RECT 90.825 123.335 91.745 123.445 ;
        RECT 90.825 123.215 93.160 123.335 ;
        RECT 97.825 123.215 98.745 123.435 ;
        RECT 100.485 123.335 101.405 123.445 ;
        RECT 100.485 123.215 102.820 123.335 ;
        RECT 107.485 123.215 108.405 123.435 ;
        RECT 90.825 122.535 100.105 123.215 ;
        RECT 100.485 122.535 109.765 123.215 ;
        RECT 110.235 122.535 112.065 123.345 ;
        RECT 112.075 122.535 113.445 123.345 ;
        RECT 15.155 122.325 15.325 122.535 ;
        RECT 16.590 122.375 16.710 122.485 ;
        RECT 16.995 122.370 17.155 122.480 ;
        RECT 17.455 122.325 17.625 122.515 ;
        RECT 18.375 122.345 18.545 122.535 ;
        RECT 19.110 122.325 19.280 122.515 ;
        RECT 19.755 122.345 19.925 122.535 ;
        RECT 23.435 122.325 23.605 122.515 ;
        RECT 25.275 122.370 25.435 122.480 ;
        RECT 25.735 122.325 25.905 122.515 ;
        RECT 29.415 122.345 29.585 122.535 ;
        RECT 29.930 122.375 30.050 122.485 ;
        RECT 33.740 122.345 33.910 122.535 ;
        RECT 35.395 122.345 35.565 122.535 ;
        RECT 36.315 122.325 36.485 122.515 ;
        RECT 37.695 122.325 37.865 122.535 ;
        RECT 38.155 122.345 38.325 122.535 ;
        RECT 39.555 122.515 39.705 122.535 ;
        RECT 39.535 122.345 39.705 122.515 ;
        RECT 42.110 122.345 42.280 122.535 ;
        RECT 47.355 122.325 47.525 122.515 ;
        RECT 48.275 122.370 48.435 122.480 ;
        RECT 49.380 122.345 49.550 122.535 ;
        RECT 50.115 122.325 50.285 122.515 ;
        RECT 50.575 122.325 50.745 122.515 ;
        RECT 51.495 122.345 51.665 122.535 ;
        RECT 54.250 122.325 54.420 122.515 ;
        RECT 55.635 122.325 55.805 122.515 ;
        RECT 57.015 122.325 57.185 122.515 ;
        RECT 58.855 122.325 59.025 122.515 ;
        RECT 61.155 122.345 61.325 122.535 ;
        RECT 62.995 122.345 63.165 122.535 ;
        RECT 63.455 122.345 63.625 122.535 ;
        RECT 64.375 122.325 64.545 122.515 ;
        RECT 64.835 122.325 65.005 122.515 ;
        RECT 66.215 122.345 66.385 122.535 ;
        RECT 66.675 122.345 66.845 122.535 ;
        RECT 74.955 122.325 75.125 122.515 ;
        RECT 77.255 122.325 77.425 122.535 ;
        RECT 80.935 122.345 81.105 122.535 ;
        RECT 84.800 122.345 84.970 122.535 ;
        RECT 86.915 122.325 87.085 122.535 ;
        RECT 90.135 122.345 90.305 122.535 ;
        RECT 96.575 122.325 96.745 122.515 ;
        RECT 97.090 122.375 97.210 122.485 ;
        RECT 98.415 122.325 98.585 122.515 ;
        RECT 99.795 122.325 99.965 122.535 ;
        RECT 104.120 122.325 104.290 122.515 ;
        RECT 104.855 122.325 105.025 122.515 ;
        RECT 106.290 122.375 106.410 122.485 ;
        RECT 106.695 122.325 106.865 122.515 ;
        RECT 108.130 122.375 108.250 122.485 ;
        RECT 109.455 122.345 109.625 122.535 ;
        RECT 109.970 122.375 110.090 122.485 ;
        RECT 111.755 122.325 111.925 122.535 ;
        RECT 113.135 122.325 113.305 122.535 ;
        RECT 15.015 121.515 16.385 122.325 ;
        RECT 17.315 121.545 18.685 122.325 ;
        RECT 18.695 121.645 22.595 122.325 ;
        RECT 18.695 121.415 19.625 121.645 ;
        RECT 22.845 121.455 23.275 122.240 ;
        RECT 23.305 121.415 24.655 122.325 ;
        RECT 25.595 121.545 26.965 122.325 ;
        RECT 27.345 121.645 36.625 122.325 ;
        RECT 27.345 121.525 29.680 121.645 ;
        RECT 27.345 121.415 28.265 121.525 ;
        RECT 34.345 121.425 35.265 121.645 ;
        RECT 36.635 121.515 38.005 122.325 ;
        RECT 38.385 121.645 47.665 122.325 ;
        RECT 38.385 121.525 40.720 121.645 ;
        RECT 38.385 121.415 39.305 121.525 ;
        RECT 45.385 121.425 46.305 121.645 ;
        RECT 48.605 121.455 49.035 122.240 ;
        RECT 49.065 121.415 50.415 122.325 ;
        RECT 50.435 121.545 51.805 122.325 ;
        RECT 51.955 121.415 54.565 122.325 ;
        RECT 54.575 121.515 55.945 122.325 ;
        RECT 55.965 121.415 57.315 122.325 ;
        RECT 57.335 121.515 59.165 122.325 ;
        RECT 59.175 121.515 64.685 122.325 ;
        RECT 64.695 121.645 73.975 122.325 ;
        RECT 66.055 121.425 66.975 121.645 ;
        RECT 71.640 121.525 73.975 121.645 ;
        RECT 73.055 121.415 73.975 121.525 ;
        RECT 74.365 121.455 74.795 122.240 ;
        RECT 74.815 121.545 76.185 122.325 ;
        RECT 76.195 121.515 77.565 122.325 ;
        RECT 77.945 121.645 87.225 122.325 ;
        RECT 87.605 121.645 96.885 122.325 ;
        RECT 77.945 121.525 80.280 121.645 ;
        RECT 77.945 121.415 78.865 121.525 ;
        RECT 84.945 121.425 85.865 121.645 ;
        RECT 87.605 121.525 89.940 121.645 ;
        RECT 87.605 121.415 88.525 121.525 ;
        RECT 94.605 121.425 95.525 121.645 ;
        RECT 97.355 121.545 98.725 122.325 ;
        RECT 98.735 121.515 100.105 122.325 ;
        RECT 100.125 121.455 100.555 122.240 ;
        RECT 100.805 121.645 104.705 122.325 ;
        RECT 103.775 121.415 104.705 121.645 ;
        RECT 104.715 121.545 106.085 122.325 ;
        RECT 106.555 121.545 107.925 122.325 ;
        RECT 108.395 121.515 112.065 122.325 ;
        RECT 112.075 121.515 113.445 122.325 ;
      LAYER nwell ;
        RECT 14.820 118.295 113.640 121.125 ;
      LAYER pwell ;
        RECT 15.015 117.095 16.385 117.905 ;
        RECT 16.395 117.095 19.145 117.905 ;
        RECT 19.355 117.775 21.565 118.005 ;
        RECT 24.285 117.775 25.215 117.995 ;
        RECT 19.355 117.095 29.725 117.775 ;
        RECT 30.205 117.095 31.555 118.005 ;
        RECT 31.575 117.095 33.405 117.905 ;
        RECT 33.415 117.095 34.785 117.875 ;
        RECT 35.725 117.180 36.155 117.965 ;
        RECT 36.175 117.095 37.545 117.905 ;
        RECT 37.555 117.095 41.225 117.905 ;
        RECT 41.245 117.095 42.595 118.005 ;
        RECT 44.825 117.895 45.745 118.005 ;
        RECT 43.075 117.095 44.445 117.875 ;
        RECT 44.825 117.775 47.160 117.895 ;
        RECT 51.825 117.775 52.745 117.995 ;
        RECT 44.825 117.095 54.105 117.775 ;
        RECT 54.115 117.095 55.945 117.905 ;
        RECT 55.955 117.095 61.465 117.905 ;
        RECT 61.485 117.180 61.915 117.965 ;
        RECT 61.935 117.095 64.685 117.905 ;
        RECT 64.695 117.095 70.205 117.905 ;
        RECT 70.225 117.095 71.575 118.005 ;
        RECT 74.795 117.775 75.725 118.005 ;
        RECT 71.825 117.095 75.725 117.775 ;
        RECT 75.735 117.095 81.245 117.905 ;
        RECT 81.265 117.095 82.615 118.005 ;
        RECT 83.105 117.095 84.455 118.005 ;
        RECT 84.475 117.095 85.845 117.875 ;
        RECT 85.855 117.095 87.225 117.905 ;
        RECT 87.245 117.180 87.675 117.965 ;
        RECT 88.155 117.095 90.905 117.905 ;
        RECT 90.915 117.095 92.285 117.875 ;
        RECT 92.755 117.095 94.585 117.905 ;
        RECT 94.595 117.095 100.105 117.905 ;
        RECT 100.115 117.095 105.625 117.905 ;
        RECT 105.645 117.095 106.995 118.005 ;
        RECT 107.015 117.095 108.385 117.875 ;
        RECT 108.395 117.095 109.765 117.875 ;
        RECT 110.235 117.095 112.065 117.905 ;
        RECT 112.075 117.095 113.445 117.905 ;
        RECT 15.155 116.885 15.325 117.095 ;
        RECT 16.995 116.930 17.155 117.040 ;
        RECT 18.835 116.905 19.005 117.095 ;
        RECT 22.515 116.885 22.685 117.075 ;
        RECT 29.415 116.905 29.585 117.095 ;
        RECT 29.930 116.935 30.050 117.045 ;
        RECT 30.335 116.905 30.505 117.095 ;
        RECT 33.095 116.905 33.265 117.095 ;
        RECT 33.555 116.885 33.725 117.095 ;
        RECT 34.070 116.935 34.190 117.045 ;
        RECT 35.395 116.885 35.565 117.075 ;
        RECT 35.910 116.935 36.030 117.045 ;
        RECT 37.235 116.905 37.405 117.095 ;
        RECT 40.915 116.905 41.085 117.095 ;
        RECT 41.375 116.885 41.545 117.095 ;
        RECT 42.810 116.935 42.930 117.045 ;
        RECT 43.215 116.905 43.385 117.095 ;
        RECT 46.895 116.885 47.065 117.075 ;
        RECT 47.355 116.885 47.525 117.075 ;
        RECT 50.115 116.885 50.285 117.075 ;
        RECT 53.795 116.905 53.965 117.095 ;
        RECT 55.635 116.885 55.805 117.095 ;
        RECT 56.100 116.885 56.270 117.075 ;
        RECT 61.155 116.905 61.325 117.095 ;
        RECT 63.915 116.885 64.085 117.075 ;
        RECT 64.375 116.905 64.545 117.095 ;
        RECT 69.435 116.885 69.605 117.075 ;
        RECT 69.895 116.905 70.065 117.095 ;
        RECT 70.355 116.905 70.525 117.095 ;
        RECT 70.815 116.885 70.985 117.075 ;
        RECT 71.330 116.935 71.450 117.045 ;
        RECT 71.740 116.885 71.910 117.075 ;
        RECT 75.140 116.905 75.310 117.095 ;
        RECT 77.255 116.885 77.425 117.075 ;
        RECT 77.715 116.885 77.885 117.075 ;
        RECT 79.150 116.935 79.270 117.045 ;
        RECT 80.935 116.905 81.105 117.095 ;
        RECT 82.315 116.905 82.485 117.095 ;
        RECT 82.775 117.045 82.945 117.075 ;
        RECT 82.775 116.935 82.950 117.045 ;
        RECT 82.775 116.885 82.945 116.935 ;
        RECT 83.235 116.905 83.405 117.095 ;
        RECT 84.155 116.885 84.325 117.075 ;
        RECT 84.615 116.905 84.785 117.095 ;
        RECT 85.535 116.885 85.705 117.075 ;
        RECT 86.915 116.905 87.085 117.095 ;
        RECT 87.890 116.935 88.010 117.045 ;
        RECT 89.215 116.885 89.385 117.075 ;
        RECT 89.675 116.885 89.845 117.075 ;
        RECT 90.595 116.905 90.765 117.095 ;
        RECT 91.055 116.905 91.225 117.095 ;
        RECT 92.490 116.935 92.610 117.045 ;
        RECT 94.275 116.885 94.445 117.095 ;
        RECT 94.735 116.885 94.905 117.075 ;
        RECT 98.415 116.885 98.585 117.075 ;
        RECT 98.875 116.885 99.045 117.075 ;
        RECT 99.795 116.905 99.965 117.095 ;
        RECT 101.175 116.930 101.335 117.040 ;
        RECT 101.635 116.885 101.805 117.075 ;
        RECT 105.315 116.905 105.485 117.095 ;
        RECT 105.775 116.905 105.945 117.095 ;
        RECT 107.155 116.905 107.325 117.095 ;
        RECT 109.455 116.905 109.625 117.095 ;
        RECT 109.970 116.935 110.090 117.045 ;
        RECT 111.755 116.905 111.925 117.095 ;
        RECT 113.135 116.885 113.305 117.095 ;
        RECT 15.015 116.075 16.385 116.885 ;
        RECT 17.315 116.075 22.825 116.885 ;
        RECT 22.845 116.015 23.275 116.800 ;
        RECT 23.495 116.205 33.865 116.885 ;
        RECT 23.495 115.975 25.705 116.205 ;
        RECT 28.425 115.985 29.355 116.205 ;
        RECT 34.335 116.105 35.705 116.885 ;
        RECT 36.175 116.075 41.685 116.885 ;
        RECT 41.695 116.075 47.205 116.885 ;
        RECT 47.215 116.105 48.585 116.885 ;
        RECT 48.605 116.015 49.035 116.800 ;
        RECT 49.055 116.075 50.425 116.885 ;
        RECT 50.435 116.075 55.945 116.885 ;
        RECT 55.955 115.975 58.565 116.885 ;
        RECT 58.715 116.075 64.225 116.885 ;
        RECT 64.235 116.075 69.745 116.885 ;
        RECT 69.765 115.975 71.115 116.885 ;
        RECT 71.595 115.975 74.205 116.885 ;
        RECT 74.365 116.015 74.795 116.800 ;
        RECT 74.815 116.075 77.565 116.885 ;
        RECT 77.575 116.105 78.945 116.885 ;
        RECT 79.415 116.075 83.085 116.885 ;
        RECT 83.105 115.975 84.455 116.885 ;
        RECT 84.475 116.075 85.845 116.885 ;
        RECT 85.855 116.075 89.525 116.885 ;
        RECT 89.535 116.105 90.905 116.885 ;
        RECT 90.915 116.075 94.585 116.885 ;
        RECT 94.595 116.105 95.965 116.885 ;
        RECT 95.975 116.075 98.725 116.885 ;
        RECT 98.735 116.105 100.105 116.885 ;
        RECT 100.125 116.015 100.555 116.800 ;
        RECT 101.495 116.205 111.865 116.885 ;
        RECT 106.005 115.985 106.935 116.205 ;
        RECT 109.655 115.975 111.865 116.205 ;
        RECT 112.075 116.075 113.445 116.885 ;
      LAYER nwell ;
        RECT 14.820 112.855 113.640 115.685 ;
      LAYER pwell ;
        RECT 15.015 111.655 16.385 112.465 ;
        RECT 16.855 111.655 22.365 112.465 ;
        RECT 22.375 111.655 23.745 112.435 ;
        RECT 23.755 111.655 25.125 112.435 ;
        RECT 25.335 112.335 27.545 112.565 ;
        RECT 30.265 112.335 31.195 112.555 ;
        RECT 25.335 111.655 35.705 112.335 ;
        RECT 35.725 111.740 36.155 112.525 ;
        RECT 37.105 111.655 38.455 112.565 ;
        RECT 38.475 111.655 40.305 112.465 ;
        RECT 40.315 111.655 41.685 112.435 ;
        RECT 42.155 111.655 43.525 112.435 ;
        RECT 43.735 112.335 45.945 112.565 ;
        RECT 48.665 112.335 49.595 112.555 ;
        RECT 43.735 111.655 54.105 112.335 ;
        RECT 54.115 111.655 55.485 112.435 ;
        RECT 56.425 111.655 57.775 112.565 ;
        RECT 57.805 111.655 59.155 112.565 ;
        RECT 59.635 111.655 61.005 112.435 ;
        RECT 61.485 111.740 61.915 112.525 ;
        RECT 62.855 111.655 64.225 112.435 ;
        RECT 64.435 112.335 66.645 112.565 ;
        RECT 69.365 112.335 70.295 112.555 ;
        RECT 75.015 112.335 77.225 112.565 ;
        RECT 79.945 112.335 80.875 112.555 ;
        RECT 64.435 111.655 74.805 112.335 ;
        RECT 75.015 111.655 85.385 112.335 ;
        RECT 85.395 111.655 86.765 112.435 ;
        RECT 87.245 111.740 87.675 112.525 ;
        RECT 88.815 112.335 91.025 112.565 ;
        RECT 93.745 112.335 94.675 112.555 ;
        RECT 88.815 111.655 99.185 112.335 ;
        RECT 99.195 111.655 100.565 112.435 ;
        RECT 101.695 112.335 103.905 112.565 ;
        RECT 106.625 112.335 107.555 112.555 ;
        RECT 101.695 111.655 112.065 112.335 ;
        RECT 112.075 111.655 113.445 112.465 ;
        RECT 15.155 111.445 15.325 111.655 ;
        RECT 16.590 111.495 16.710 111.605 ;
        RECT 19.755 111.445 19.925 111.635 ;
        RECT 21.135 111.445 21.305 111.635 ;
        RECT 21.595 111.445 21.765 111.635 ;
        RECT 22.055 111.465 22.225 111.655 ;
        RECT 22.515 111.465 22.685 111.655 ;
        RECT 23.435 111.445 23.605 111.635 ;
        RECT 23.895 111.465 24.065 111.655 ;
        RECT 24.815 111.445 24.985 111.635 ;
        RECT 26.195 111.445 26.365 111.635 ;
        RECT 27.575 111.445 27.745 111.635 ;
        RECT 35.395 111.465 35.565 111.655 ;
        RECT 36.775 111.500 36.935 111.610 ;
        RECT 38.155 111.465 38.325 111.655 ;
        RECT 39.995 111.465 40.165 111.655 ;
        RECT 41.375 111.465 41.545 111.655 ;
        RECT 41.890 111.495 42.010 111.605 ;
        RECT 42.295 111.465 42.465 111.655 ;
        RECT 48.275 111.445 48.445 111.635 ;
        RECT 53.795 111.465 53.965 111.655 ;
        RECT 54.255 111.465 54.425 111.655 ;
        RECT 56.095 111.500 56.255 111.610 ;
        RECT 56.555 111.465 56.725 111.655 ;
        RECT 57.935 111.465 58.105 111.655 ;
        RECT 59.315 111.605 59.485 111.635 ;
        RECT 59.315 111.495 59.490 111.605 ;
        RECT 59.315 111.445 59.485 111.495 ;
        RECT 60.695 111.465 60.865 111.655 ;
        RECT 61.210 111.495 61.330 111.605 ;
        RECT 62.535 111.500 62.695 111.610 ;
        RECT 62.995 111.465 63.165 111.655 ;
        RECT 69.895 111.445 70.065 111.635 ;
        RECT 70.410 111.495 70.530 111.605 ;
        RECT 70.815 111.445 70.985 111.635 ;
        RECT 72.195 111.445 72.365 111.635 ;
        RECT 74.035 111.490 74.195 111.600 ;
        RECT 74.495 111.465 74.665 111.655 ;
        RECT 85.075 111.445 85.245 111.655 ;
        RECT 86.455 111.465 86.625 111.655 ;
        RECT 86.970 111.495 87.090 111.605 ;
        RECT 88.295 111.500 88.455 111.610 ;
        RECT 95.655 111.445 95.825 111.635 ;
        RECT 97.035 111.445 97.205 111.635 ;
        RECT 98.415 111.445 98.585 111.635 ;
        RECT 98.875 111.445 99.045 111.655 ;
        RECT 100.255 111.465 100.425 111.655 ;
        RECT 101.175 111.500 101.335 111.610 ;
        RECT 110.835 111.445 111.005 111.635 ;
        RECT 111.755 111.465 111.925 111.655 ;
        RECT 113.135 111.445 113.305 111.655 ;
        RECT 15.015 110.635 16.385 111.445 ;
        RECT 16.395 110.635 20.065 111.445 ;
        RECT 20.085 110.535 21.435 111.445 ;
        RECT 21.465 110.535 22.815 111.445 ;
        RECT 22.845 110.575 23.275 111.360 ;
        RECT 23.305 110.535 24.655 111.445 ;
        RECT 24.685 110.535 26.035 111.445 ;
        RECT 26.055 110.665 27.425 111.445 ;
        RECT 27.435 110.765 37.805 111.445 ;
        RECT 31.945 110.545 32.875 110.765 ;
        RECT 35.595 110.535 37.805 110.765 ;
        RECT 38.215 110.765 48.585 111.445 ;
        RECT 38.215 110.535 40.425 110.765 ;
        RECT 43.145 110.545 44.075 110.765 ;
        RECT 48.605 110.575 49.035 111.360 ;
        RECT 49.255 110.765 59.625 111.445 ;
        RECT 59.835 110.765 70.205 111.445 ;
        RECT 49.255 110.535 51.465 110.765 ;
        RECT 54.185 110.545 55.115 110.765 ;
        RECT 59.835 110.535 62.045 110.765 ;
        RECT 64.765 110.545 65.695 110.765 ;
        RECT 70.675 110.665 72.045 111.445 ;
        RECT 72.055 110.665 73.425 111.445 ;
        RECT 74.365 110.575 74.795 111.360 ;
        RECT 75.015 110.765 85.385 111.445 ;
        RECT 85.595 110.765 95.965 111.445 ;
        RECT 75.015 110.535 77.225 110.765 ;
        RECT 79.945 110.545 80.875 110.765 ;
        RECT 85.595 110.535 87.805 110.765 ;
        RECT 90.525 110.545 91.455 110.765 ;
        RECT 95.985 110.535 97.335 111.445 ;
        RECT 97.365 110.535 98.715 111.445 ;
        RECT 98.745 110.535 100.095 111.445 ;
        RECT 100.125 110.575 100.555 111.360 ;
        RECT 100.775 110.765 111.145 111.445 ;
        RECT 100.775 110.535 102.985 110.765 ;
        RECT 105.705 110.545 106.635 110.765 ;
        RECT 112.075 110.635 113.445 111.445 ;
      LAYER nwell ;
        RECT 14.820 107.415 113.640 110.245 ;
      LAYER pwell ;
        RECT 15.015 106.215 16.385 107.025 ;
        RECT 17.315 106.215 22.825 107.025 ;
        RECT 22.845 106.300 23.275 107.085 ;
        RECT 23.495 106.895 25.705 107.125 ;
        RECT 28.425 106.895 29.355 107.115 ;
        RECT 23.495 106.215 33.865 106.895 ;
        RECT 33.875 106.215 35.705 107.025 ;
        RECT 35.725 106.300 36.155 107.085 ;
        RECT 36.635 106.215 42.145 107.025 ;
        RECT 42.165 106.215 43.515 107.125 ;
        RECT 43.535 106.215 47.205 107.025 ;
        RECT 47.225 106.215 48.575 107.125 ;
        RECT 48.605 106.300 49.035 107.085 ;
        RECT 49.525 106.215 50.875 107.125 ;
        RECT 51.095 106.895 53.305 107.125 ;
        RECT 56.025 106.895 56.955 107.115 ;
        RECT 51.095 106.215 61.465 106.895 ;
        RECT 61.485 106.300 61.915 107.085 ;
        RECT 62.395 106.215 65.145 107.025 ;
        RECT 65.155 106.215 70.665 107.025 ;
        RECT 70.685 106.215 72.035 107.125 ;
        RECT 72.525 106.215 73.875 107.125 ;
        RECT 74.365 106.300 74.795 107.085 ;
        RECT 75.285 106.215 76.635 107.125 ;
        RECT 76.855 106.895 79.065 107.125 ;
        RECT 81.785 106.895 82.715 107.115 ;
        RECT 76.855 106.215 87.225 106.895 ;
        RECT 87.245 106.300 87.675 107.085 ;
        RECT 88.165 106.215 89.515 107.125 ;
        RECT 89.735 106.895 91.945 107.125 ;
        RECT 94.665 106.895 95.595 107.115 ;
        RECT 89.735 106.215 100.105 106.895 ;
        RECT 100.125 106.300 100.555 107.085 ;
        RECT 100.575 106.215 101.945 107.025 ;
        RECT 101.955 106.215 105.625 107.025 ;
        RECT 105.645 106.215 106.995 107.125 ;
        RECT 107.015 106.215 110.685 107.025 ;
        RECT 110.695 106.215 112.065 106.995 ;
        RECT 112.075 106.215 113.445 107.025 ;
        RECT 15.155 106.025 15.325 106.215 ;
        RECT 16.995 106.060 17.155 106.170 ;
        RECT 22.515 106.025 22.685 106.215 ;
        RECT 33.555 106.025 33.725 106.215 ;
        RECT 35.395 106.025 35.565 106.215 ;
        RECT 36.370 106.055 36.490 106.165 ;
        RECT 41.835 106.025 42.005 106.215 ;
        RECT 43.215 106.025 43.385 106.215 ;
        RECT 46.895 106.025 47.065 106.215 ;
        RECT 47.355 106.025 47.525 106.215 ;
        RECT 49.250 106.055 49.370 106.165 ;
        RECT 49.655 106.025 49.825 106.215 ;
        RECT 61.155 106.025 61.325 106.215 ;
        RECT 62.130 106.055 62.250 106.165 ;
        RECT 64.835 106.025 65.005 106.215 ;
        RECT 70.355 106.025 70.525 106.215 ;
        RECT 71.735 106.025 71.905 106.215 ;
        RECT 72.250 106.055 72.370 106.165 ;
        RECT 72.655 106.025 72.825 106.215 ;
        RECT 74.090 106.055 74.210 106.165 ;
        RECT 75.010 106.055 75.130 106.165 ;
        RECT 75.415 106.025 75.585 106.215 ;
        RECT 86.915 106.025 87.085 106.215 ;
        RECT 87.890 106.055 88.010 106.165 ;
        RECT 88.295 106.025 88.465 106.215 ;
        RECT 99.795 106.025 99.965 106.215 ;
        RECT 101.635 106.025 101.805 106.215 ;
        RECT 105.315 106.025 105.485 106.215 ;
        RECT 106.695 106.025 106.865 106.215 ;
        RECT 110.375 106.025 110.545 106.215 ;
        RECT 111.745 106.025 111.915 106.215 ;
        RECT 113.135 106.025 113.305 106.215 ;
      LAYER nwell ;
        RECT 20.485 54.580 29.875 66.420 ;
        RECT 31.685 54.590 41.075 66.430 ;
        RECT 42.905 54.560 52.295 66.400 ;
        RECT 54.155 54.540 63.545 66.380 ;
        RECT 65.375 54.530 74.765 66.370 ;
        RECT 76.615 54.520 86.005 66.360 ;
        RECT 87.865 54.530 97.255 66.370 ;
        RECT 99.145 54.520 108.535 66.360 ;
        RECT 110.415 54.520 119.805 66.360 ;
        RECT 121.665 54.520 131.055 66.360 ;
        RECT 132.415 54.490 139.375 66.330 ;
        RECT 20.655 49.020 23.115 53.210 ;
      LAYER pwell ;
        RECT 20.555 45.340 22.915 48.340 ;
      LAYER nwell ;
        RECT 24.735 45.940 29.125 53.130 ;
        RECT 31.855 49.030 34.315 53.220 ;
      LAYER pwell ;
        RECT 31.755 45.350 34.115 48.350 ;
      LAYER nwell ;
        RECT 35.935 45.950 40.325 53.140 ;
        RECT 43.075 49.000 45.535 53.190 ;
      LAYER pwell ;
        RECT 42.975 45.320 45.335 48.320 ;
      LAYER nwell ;
        RECT 47.155 45.920 51.545 53.110 ;
        RECT 54.325 48.980 56.785 53.170 ;
      LAYER pwell ;
        RECT 54.225 45.300 56.585 48.300 ;
      LAYER nwell ;
        RECT 58.405 45.900 62.795 53.090 ;
        RECT 65.545 48.970 68.005 53.160 ;
      LAYER pwell ;
        RECT 65.445 45.290 67.805 48.290 ;
      LAYER nwell ;
        RECT 69.625 45.890 74.015 53.080 ;
        RECT 76.785 48.960 79.245 53.150 ;
      LAYER pwell ;
        RECT 76.685 45.280 79.045 48.280 ;
      LAYER nwell ;
        RECT 80.865 45.880 85.255 53.070 ;
        RECT 88.035 48.970 90.495 53.160 ;
      LAYER pwell ;
        RECT 87.935 45.290 90.295 48.290 ;
      LAYER nwell ;
        RECT 92.115 45.890 96.505 53.080 ;
        RECT 99.315 48.960 101.775 53.150 ;
      LAYER pwell ;
        RECT 99.215 45.280 101.575 48.280 ;
      LAYER nwell ;
        RECT 103.395 45.880 107.785 53.070 ;
        RECT 110.585 48.960 113.045 53.150 ;
      LAYER pwell ;
        RECT 110.485 45.280 112.845 48.280 ;
      LAYER nwell ;
        RECT 114.665 45.880 119.055 53.070 ;
        RECT 121.835 48.960 124.295 53.150 ;
      LAYER pwell ;
        RECT 121.735 45.280 124.095 48.280 ;
      LAYER nwell ;
        RECT 125.915 45.880 130.305 53.070 ;
        RECT 19.615 32.280 24.005 39.470 ;
      LAYER pwell ;
        RECT 25.825 37.070 28.185 40.070 ;
      LAYER nwell ;
        RECT 25.625 32.200 28.085 36.390 ;
        RECT 30.895 32.280 35.285 39.470 ;
      LAYER pwell ;
        RECT 37.105 37.070 39.465 40.070 ;
      LAYER nwell ;
        RECT 36.905 32.200 39.365 36.390 ;
        RECT 42.185 32.260 46.575 39.450 ;
      LAYER pwell ;
        RECT 48.395 37.050 50.755 40.050 ;
      LAYER nwell ;
        RECT 48.195 32.180 50.655 36.370 ;
        RECT 53.405 32.260 57.795 39.450 ;
      LAYER pwell ;
        RECT 59.615 37.050 61.975 40.050 ;
      LAYER nwell ;
        RECT 59.415 32.180 61.875 36.370 ;
        RECT 64.605 32.260 68.995 39.450 ;
      LAYER pwell ;
        RECT 70.815 37.050 73.175 40.050 ;
      LAYER nwell ;
        RECT 70.615 32.180 73.075 36.370 ;
        RECT 75.895 32.250 80.285 39.440 ;
      LAYER pwell ;
        RECT 82.105 37.040 84.465 40.040 ;
      LAYER nwell ;
        RECT 81.905 32.170 84.365 36.360 ;
        RECT 87.135 32.270 91.525 39.460 ;
      LAYER pwell ;
        RECT 93.345 37.060 95.705 40.060 ;
      LAYER nwell ;
        RECT 93.145 32.190 95.605 36.380 ;
        RECT 98.345 32.290 102.735 39.480 ;
      LAYER pwell ;
        RECT 104.555 37.080 106.915 40.080 ;
      LAYER nwell ;
        RECT 104.355 32.210 106.815 36.400 ;
        RECT 109.545 32.330 113.935 39.520 ;
      LAYER pwell ;
        RECT 115.755 37.120 118.115 40.120 ;
      LAYER nwell ;
        RECT 115.555 32.250 118.015 36.440 ;
        RECT 120.755 32.350 125.145 39.540 ;
      LAYER pwell ;
        RECT 126.965 37.140 129.325 40.140 ;
      LAYER nwell ;
        RECT 126.765 32.270 129.225 36.460 ;
        RECT 18.865 18.990 28.255 30.830 ;
        RECT 30.145 18.990 39.535 30.830 ;
        RECT 41.435 18.970 50.825 30.810 ;
        RECT 52.655 18.970 62.045 30.810 ;
        RECT 63.855 18.970 73.245 30.810 ;
        RECT 75.145 18.960 84.535 30.800 ;
        RECT 86.385 18.980 95.775 30.820 ;
        RECT 97.595 19.000 106.985 30.840 ;
        RECT 108.795 19.040 118.185 30.880 ;
        RECT 120.005 19.060 129.395 30.900 ;
        RECT 131.725 19.030 138.685 30.870 ;
      LAYER li1 ;
        RECT 15.010 203.945 113.450 204.115 ;
        RECT 15.095 203.195 16.305 203.945 ;
        RECT 17.400 203.400 22.745 203.945 ;
        RECT 15.095 202.655 15.615 203.195 ;
        RECT 15.785 202.485 16.305 203.025 ;
        RECT 15.095 201.395 16.305 202.485 ;
        RECT 18.990 201.830 19.340 203.080 ;
        RECT 20.820 202.570 21.160 203.400 ;
        RECT 22.915 203.220 23.205 203.945 ;
        RECT 23.375 203.195 24.585 203.945 ;
        RECT 24.760 203.400 30.105 203.945 ;
        RECT 30.280 203.400 35.625 203.945 ;
        RECT 17.400 201.395 22.745 201.830 ;
        RECT 22.915 201.395 23.205 202.560 ;
        RECT 23.375 202.485 23.895 203.025 ;
        RECT 24.065 202.655 24.585 203.195 ;
        RECT 23.375 201.395 24.585 202.485 ;
        RECT 26.350 201.830 26.700 203.080 ;
        RECT 28.180 202.570 28.520 203.400 ;
        RECT 31.870 201.830 32.220 203.080 ;
        RECT 33.700 202.570 34.040 203.400 ;
        RECT 35.795 203.220 36.085 203.945 ;
        RECT 36.255 203.195 37.465 203.945 ;
        RECT 37.640 203.400 42.985 203.945 ;
        RECT 43.160 203.400 48.505 203.945 ;
        RECT 24.760 201.395 30.105 201.830 ;
        RECT 30.280 201.395 35.625 201.830 ;
        RECT 35.795 201.395 36.085 202.560 ;
        RECT 36.255 202.485 36.775 203.025 ;
        RECT 36.945 202.655 37.465 203.195 ;
        RECT 36.255 201.395 37.465 202.485 ;
        RECT 39.230 201.830 39.580 203.080 ;
        RECT 41.060 202.570 41.400 203.400 ;
        RECT 44.750 201.830 45.100 203.080 ;
        RECT 46.580 202.570 46.920 203.400 ;
        RECT 48.675 203.220 48.965 203.945 ;
        RECT 49.140 203.400 54.485 203.945 ;
        RECT 54.660 203.400 60.005 203.945 ;
        RECT 37.640 201.395 42.985 201.830 ;
        RECT 43.160 201.395 48.505 201.830 ;
        RECT 48.675 201.395 48.965 202.560 ;
        RECT 50.730 201.830 51.080 203.080 ;
        RECT 52.560 202.570 52.900 203.400 ;
        RECT 56.250 201.830 56.600 203.080 ;
        RECT 58.080 202.570 58.420 203.400 ;
        RECT 60.175 203.270 60.435 203.775 ;
        RECT 60.615 203.565 60.945 203.945 ;
        RECT 61.125 203.395 61.295 203.775 ;
        RECT 60.175 202.470 60.345 203.270 ;
        RECT 60.630 203.225 61.295 203.395 ;
        RECT 60.630 202.970 60.800 203.225 ;
        RECT 61.555 203.220 61.845 203.945 ;
        RECT 62.020 203.400 67.365 203.945 ;
        RECT 67.540 203.400 72.885 203.945 ;
        RECT 60.515 202.640 60.800 202.970 ;
        RECT 61.035 202.675 61.365 203.045 ;
        RECT 60.630 202.495 60.800 202.640 ;
        RECT 49.140 201.395 54.485 201.830 ;
        RECT 54.660 201.395 60.005 201.830 ;
        RECT 60.175 201.565 60.445 202.470 ;
        RECT 60.630 202.325 61.295 202.495 ;
        RECT 60.615 201.395 60.945 202.155 ;
        RECT 61.125 201.565 61.295 202.325 ;
        RECT 61.555 201.395 61.845 202.560 ;
        RECT 63.610 201.830 63.960 203.080 ;
        RECT 65.440 202.570 65.780 203.400 ;
        RECT 69.130 201.830 69.480 203.080 ;
        RECT 70.960 202.570 71.300 203.400 ;
        RECT 73.115 203.125 73.325 203.945 ;
        RECT 73.495 203.145 73.825 203.775 ;
        RECT 73.495 202.545 73.745 203.145 ;
        RECT 73.995 203.125 74.225 203.945 ;
        RECT 74.435 203.220 74.725 203.945 ;
        RECT 74.895 203.195 76.105 203.945 ;
        RECT 76.280 203.400 81.625 203.945 ;
        RECT 81.800 203.400 87.145 203.945 ;
        RECT 73.915 202.705 74.245 202.955 ;
        RECT 62.020 201.395 67.365 201.830 ;
        RECT 67.540 201.395 72.885 201.830 ;
        RECT 73.115 201.395 73.325 202.535 ;
        RECT 73.495 201.565 73.825 202.545 ;
        RECT 73.995 201.395 74.225 202.535 ;
        RECT 74.435 201.395 74.725 202.560 ;
        RECT 74.895 202.485 75.415 203.025 ;
        RECT 75.585 202.655 76.105 203.195 ;
        RECT 74.895 201.395 76.105 202.485 ;
        RECT 77.870 201.830 78.220 203.080 ;
        RECT 79.700 202.570 80.040 203.400 ;
        RECT 83.390 201.830 83.740 203.080 ;
        RECT 85.220 202.570 85.560 203.400 ;
        RECT 87.315 203.220 87.605 203.945 ;
        RECT 87.775 203.195 88.985 203.945 ;
        RECT 89.160 203.400 94.505 203.945 ;
        RECT 94.680 203.400 100.025 203.945 ;
        RECT 76.280 201.395 81.625 201.830 ;
        RECT 81.800 201.395 87.145 201.830 ;
        RECT 87.315 201.395 87.605 202.560 ;
        RECT 87.775 202.485 88.295 203.025 ;
        RECT 88.465 202.655 88.985 203.195 ;
        RECT 87.775 201.395 88.985 202.485 ;
        RECT 90.750 201.830 91.100 203.080 ;
        RECT 92.580 202.570 92.920 203.400 ;
        RECT 96.270 201.830 96.620 203.080 ;
        RECT 98.100 202.570 98.440 203.400 ;
        RECT 100.195 203.220 100.485 203.945 ;
        RECT 101.120 203.400 106.465 203.945 ;
        RECT 106.640 203.400 111.985 203.945 ;
        RECT 89.160 201.395 94.505 201.830 ;
        RECT 94.680 201.395 100.025 201.830 ;
        RECT 100.195 201.395 100.485 202.560 ;
        RECT 102.710 201.830 103.060 203.080 ;
        RECT 104.540 202.570 104.880 203.400 ;
        RECT 108.230 201.830 108.580 203.080 ;
        RECT 110.060 202.570 110.400 203.400 ;
        RECT 112.155 203.195 113.365 203.945 ;
        RECT 112.155 202.485 112.675 203.025 ;
        RECT 112.845 202.655 113.365 203.195 ;
        RECT 101.120 201.395 106.465 201.830 ;
        RECT 106.640 201.395 111.985 201.830 ;
        RECT 112.155 201.395 113.365 202.485 ;
        RECT 15.010 201.225 113.450 201.395 ;
        RECT 15.095 200.135 16.305 201.225 ;
        RECT 15.095 199.425 15.615 199.965 ;
        RECT 15.785 199.595 16.305 200.135 ;
        RECT 16.475 200.135 19.065 201.225 ;
        RECT 19.240 200.790 24.585 201.225 ;
        RECT 24.760 200.790 30.105 201.225 ;
        RECT 30.280 200.790 35.625 201.225 ;
        RECT 16.475 199.615 17.685 200.135 ;
        RECT 17.855 199.445 19.065 199.965 ;
        RECT 20.830 199.540 21.180 200.790 ;
        RECT 15.095 198.675 16.305 199.425 ;
        RECT 16.475 198.675 19.065 199.445 ;
        RECT 22.660 199.220 23.000 200.050 ;
        RECT 26.350 199.540 26.700 200.790 ;
        RECT 28.180 199.220 28.520 200.050 ;
        RECT 31.870 199.540 32.220 200.790 ;
        RECT 35.795 200.060 36.085 201.225 ;
        RECT 36.715 200.135 40.225 201.225 ;
        RECT 40.400 200.790 45.745 201.225 ;
        RECT 45.920 200.790 51.265 201.225 ;
        RECT 33.700 199.220 34.040 200.050 ;
        RECT 36.715 199.615 38.405 200.135 ;
        RECT 38.575 199.445 40.225 199.965 ;
        RECT 41.990 199.540 42.340 200.790 ;
        RECT 19.240 198.675 24.585 199.220 ;
        RECT 24.760 198.675 30.105 199.220 ;
        RECT 30.280 198.675 35.625 199.220 ;
        RECT 35.795 198.675 36.085 199.400 ;
        RECT 36.715 198.675 40.225 199.445 ;
        RECT 43.820 199.220 44.160 200.050 ;
        RECT 47.510 199.540 47.860 200.790 ;
        RECT 49.340 199.220 49.680 200.050 ;
        RECT 51.440 200.035 51.695 200.915 ;
        RECT 51.865 200.085 52.170 201.225 ;
        RECT 52.510 200.845 52.840 201.225 ;
        RECT 53.020 200.675 53.190 200.965 ;
        RECT 53.360 200.765 53.610 201.225 ;
        RECT 52.390 200.505 53.190 200.675 ;
        RECT 53.780 200.715 54.650 201.055 ;
        RECT 51.440 199.385 51.650 200.035 ;
        RECT 52.390 199.915 52.560 200.505 ;
        RECT 53.780 200.335 53.950 200.715 ;
        RECT 54.885 200.595 55.055 201.055 ;
        RECT 55.225 200.765 55.595 201.225 ;
        RECT 55.890 200.625 56.060 200.965 ;
        RECT 56.230 200.795 56.560 201.225 ;
        RECT 56.795 200.625 56.965 200.965 ;
        RECT 52.730 200.165 53.950 200.335 ;
        RECT 54.120 200.255 54.580 200.545 ;
        RECT 54.885 200.425 55.445 200.595 ;
        RECT 55.890 200.455 56.965 200.625 ;
        RECT 57.135 200.725 57.815 201.055 ;
        RECT 58.030 200.725 58.280 201.055 ;
        RECT 58.450 200.765 58.700 201.225 ;
        RECT 55.275 200.285 55.445 200.425 ;
        RECT 54.120 200.245 55.085 200.255 ;
        RECT 53.780 200.075 53.950 200.165 ;
        RECT 54.410 200.085 55.085 200.245 ;
        RECT 51.820 199.885 52.560 199.915 ;
        RECT 51.820 199.585 52.735 199.885 ;
        RECT 52.410 199.410 52.735 199.585 ;
        RECT 40.400 198.675 45.745 199.220 ;
        RECT 45.920 198.675 51.265 199.220 ;
        RECT 51.440 198.855 51.695 199.385 ;
        RECT 51.865 198.675 52.170 199.135 ;
        RECT 52.415 199.055 52.735 199.410 ;
        RECT 52.905 199.625 53.445 199.995 ;
        RECT 53.780 199.905 54.185 200.075 ;
        RECT 52.905 199.225 53.145 199.625 ;
        RECT 53.625 199.455 53.845 199.735 ;
        RECT 53.315 199.285 53.845 199.455 ;
        RECT 53.315 199.055 53.485 199.285 ;
        RECT 54.015 199.125 54.185 199.905 ;
        RECT 54.355 199.295 54.705 199.915 ;
        RECT 54.875 199.295 55.085 200.085 ;
        RECT 55.275 200.115 56.775 200.285 ;
        RECT 55.275 199.425 55.445 200.115 ;
        RECT 57.135 199.945 57.305 200.725 ;
        RECT 58.110 200.595 58.280 200.725 ;
        RECT 55.615 199.775 57.305 199.945 ;
        RECT 57.475 200.165 57.940 200.555 ;
        RECT 58.110 200.425 58.505 200.595 ;
        RECT 55.615 199.595 55.785 199.775 ;
        RECT 52.415 198.885 53.485 199.055 ;
        RECT 53.655 198.675 53.845 199.115 ;
        RECT 54.015 198.845 54.965 199.125 ;
        RECT 55.275 199.035 55.535 199.425 ;
        RECT 55.955 199.355 56.745 199.605 ;
        RECT 55.185 198.865 55.535 199.035 ;
        RECT 55.745 198.675 56.075 199.135 ;
        RECT 56.950 199.065 57.120 199.775 ;
        RECT 57.475 199.575 57.645 200.165 ;
        RECT 57.290 199.355 57.645 199.575 ;
        RECT 57.815 199.355 58.165 199.975 ;
        RECT 58.335 199.065 58.505 200.425 ;
        RECT 58.870 200.255 59.195 201.040 ;
        RECT 58.675 199.205 59.135 200.255 ;
        RECT 56.950 198.895 57.805 199.065 ;
        RECT 58.010 198.895 58.505 199.065 ;
        RECT 58.675 198.675 59.005 199.035 ;
        RECT 59.365 198.935 59.535 201.055 ;
        RECT 59.705 200.725 60.035 201.225 ;
        RECT 60.205 200.555 60.460 201.055 ;
        RECT 59.710 200.385 60.460 200.555 ;
        RECT 59.710 199.395 59.940 200.385 ;
        RECT 60.110 199.565 60.460 200.215 ;
        RECT 61.555 200.060 61.845 201.225 ;
        RECT 62.035 200.715 62.335 201.225 ;
        RECT 62.505 200.715 62.885 200.885 ;
        RECT 63.465 200.715 64.095 201.225 ;
        RECT 62.505 200.545 62.675 200.715 ;
        RECT 64.265 200.545 64.595 201.055 ;
        RECT 64.765 200.715 65.065 201.225 ;
        RECT 62.015 200.345 62.675 200.545 ;
        RECT 62.845 200.375 65.065 200.545 ;
        RECT 62.015 199.415 62.185 200.345 ;
        RECT 62.845 200.175 63.015 200.375 ;
        RECT 62.355 200.005 63.015 200.175 ;
        RECT 63.185 200.035 64.725 200.205 ;
        RECT 62.355 199.585 62.525 200.005 ;
        RECT 63.185 199.835 63.355 200.035 ;
        RECT 62.755 199.665 63.355 199.835 ;
        RECT 63.525 199.665 64.220 199.865 ;
        RECT 64.480 199.585 64.725 200.035 ;
        RECT 62.845 199.415 63.755 199.495 ;
        RECT 59.710 199.225 60.460 199.395 ;
        RECT 59.705 198.675 60.035 199.055 ;
        RECT 60.205 198.935 60.460 199.225 ;
        RECT 61.555 198.675 61.845 199.400 ;
        RECT 62.015 198.935 62.335 199.415 ;
        RECT 62.505 199.325 63.755 199.415 ;
        RECT 62.505 199.245 63.015 199.325 ;
        RECT 62.505 198.845 62.735 199.245 ;
        RECT 62.905 198.675 63.255 199.065 ;
        RECT 63.425 198.845 63.755 199.325 ;
        RECT 63.925 198.675 64.095 199.495 ;
        RECT 64.895 199.415 65.065 200.375 ;
        RECT 64.600 198.870 65.065 199.415 ;
        RECT 65.235 200.355 65.510 201.055 ;
        RECT 65.680 200.680 65.935 201.225 ;
        RECT 66.105 200.715 66.585 201.055 ;
        RECT 66.760 200.670 67.365 201.225 ;
        RECT 66.750 200.570 67.365 200.670 ;
        RECT 66.750 200.545 66.935 200.570 ;
        RECT 65.235 199.325 65.405 200.355 ;
        RECT 65.680 200.225 66.435 200.475 ;
        RECT 66.605 200.300 66.935 200.545 ;
        RECT 65.680 200.190 66.450 200.225 ;
        RECT 65.680 200.180 66.465 200.190 ;
        RECT 65.575 200.165 66.470 200.180 ;
        RECT 65.575 200.150 66.490 200.165 ;
        RECT 65.575 200.140 66.510 200.150 ;
        RECT 65.575 200.130 66.535 200.140 ;
        RECT 65.575 200.100 66.605 200.130 ;
        RECT 65.575 200.070 66.625 200.100 ;
        RECT 65.575 200.040 66.645 200.070 ;
        RECT 65.575 200.015 66.675 200.040 ;
        RECT 65.575 199.980 66.710 200.015 ;
        RECT 65.575 199.975 66.740 199.980 ;
        RECT 65.575 199.580 65.805 199.975 ;
        RECT 66.350 199.970 66.740 199.975 ;
        RECT 66.375 199.960 66.740 199.970 ;
        RECT 66.390 199.955 66.740 199.960 ;
        RECT 66.405 199.950 66.740 199.955 ;
        RECT 67.105 199.950 67.365 200.400 ;
        RECT 68.515 200.085 68.725 201.225 ;
        RECT 66.405 199.945 67.365 199.950 ;
        RECT 66.415 199.935 67.365 199.945 ;
        RECT 66.425 199.930 67.365 199.935 ;
        RECT 66.435 199.920 67.365 199.930 ;
        RECT 66.440 199.910 67.365 199.920 ;
        RECT 66.445 199.905 67.365 199.910 ;
        RECT 66.455 199.890 67.365 199.905 ;
        RECT 66.460 199.875 67.365 199.890 ;
        RECT 66.470 199.850 67.365 199.875 ;
        RECT 65.975 199.380 66.305 199.805 ;
        RECT 65.235 198.845 65.495 199.325 ;
        RECT 65.665 198.675 65.915 199.215 ;
        RECT 66.085 198.895 66.305 199.380 ;
        RECT 66.475 199.780 67.365 199.850 ;
        RECT 68.895 200.075 69.225 201.055 ;
        RECT 69.395 200.085 69.625 201.225 ;
        RECT 66.475 199.055 66.645 199.780 ;
        RECT 66.815 199.225 67.365 199.610 ;
        RECT 66.475 198.885 67.365 199.055 ;
        RECT 68.515 198.675 68.725 199.495 ;
        RECT 68.895 199.475 69.145 200.075 ;
        RECT 69.840 200.035 70.095 200.915 ;
        RECT 70.265 200.085 70.570 201.225 ;
        RECT 70.910 200.845 71.240 201.225 ;
        RECT 71.420 200.675 71.590 200.965 ;
        RECT 71.760 200.765 72.010 201.225 ;
        RECT 70.790 200.505 71.590 200.675 ;
        RECT 72.180 200.715 73.050 201.055 ;
        RECT 69.315 199.665 69.645 199.915 ;
        RECT 68.895 198.845 69.225 199.475 ;
        RECT 69.395 198.675 69.625 199.495 ;
        RECT 69.840 199.385 70.050 200.035 ;
        RECT 70.790 199.915 70.960 200.505 ;
        RECT 72.180 200.335 72.350 200.715 ;
        RECT 73.285 200.595 73.455 201.055 ;
        RECT 73.625 200.765 73.995 201.225 ;
        RECT 74.290 200.625 74.460 200.965 ;
        RECT 74.630 200.795 74.960 201.225 ;
        RECT 75.195 200.625 75.365 200.965 ;
        RECT 71.130 200.165 72.350 200.335 ;
        RECT 72.520 200.255 72.980 200.545 ;
        RECT 73.285 200.425 73.845 200.595 ;
        RECT 74.290 200.455 75.365 200.625 ;
        RECT 75.535 200.725 76.215 201.055 ;
        RECT 76.430 200.725 76.680 201.055 ;
        RECT 76.850 200.765 77.100 201.225 ;
        RECT 73.675 200.285 73.845 200.425 ;
        RECT 72.520 200.245 73.485 200.255 ;
        RECT 72.180 200.075 72.350 200.165 ;
        RECT 72.810 200.085 73.485 200.245 ;
        RECT 70.220 199.885 70.960 199.915 ;
        RECT 70.220 199.585 71.135 199.885 ;
        RECT 70.810 199.410 71.135 199.585 ;
        RECT 69.840 198.855 70.095 199.385 ;
        RECT 70.265 198.675 70.570 199.135 ;
        RECT 70.815 199.055 71.135 199.410 ;
        RECT 71.305 199.625 71.845 199.995 ;
        RECT 72.180 199.905 72.585 200.075 ;
        RECT 71.305 199.225 71.545 199.625 ;
        RECT 72.025 199.455 72.245 199.735 ;
        RECT 71.715 199.285 72.245 199.455 ;
        RECT 71.715 199.055 71.885 199.285 ;
        RECT 72.415 199.125 72.585 199.905 ;
        RECT 72.755 199.295 73.105 199.915 ;
        RECT 73.275 199.295 73.485 200.085 ;
        RECT 73.675 200.115 75.175 200.285 ;
        RECT 73.675 199.425 73.845 200.115 ;
        RECT 75.535 199.945 75.705 200.725 ;
        RECT 76.510 200.595 76.680 200.725 ;
        RECT 74.015 199.775 75.705 199.945 ;
        RECT 75.875 200.165 76.340 200.555 ;
        RECT 76.510 200.425 76.905 200.595 ;
        RECT 74.015 199.595 74.185 199.775 ;
        RECT 70.815 198.885 71.885 199.055 ;
        RECT 72.055 198.675 72.245 199.115 ;
        RECT 72.415 198.845 73.365 199.125 ;
        RECT 73.675 199.035 73.935 199.425 ;
        RECT 74.355 199.355 75.145 199.605 ;
        RECT 73.585 198.865 73.935 199.035 ;
        RECT 74.145 198.675 74.475 199.135 ;
        RECT 75.350 199.065 75.520 199.775 ;
        RECT 75.875 199.575 76.045 200.165 ;
        RECT 75.690 199.355 76.045 199.575 ;
        RECT 76.215 199.355 76.565 199.975 ;
        RECT 76.735 199.065 76.905 200.425 ;
        RECT 77.270 200.255 77.595 201.040 ;
        RECT 77.075 199.205 77.535 200.255 ;
        RECT 75.350 198.895 76.205 199.065 ;
        RECT 76.410 198.895 76.905 199.065 ;
        RECT 77.075 198.675 77.405 199.035 ;
        RECT 77.765 198.935 77.935 201.055 ;
        RECT 78.105 200.725 78.435 201.225 ;
        RECT 78.605 200.555 78.860 201.055 ;
        RECT 78.110 200.385 78.860 200.555 ;
        RECT 78.110 199.395 78.340 200.385 ;
        RECT 78.510 199.565 78.860 200.215 ;
        RECT 79.095 200.085 79.305 201.225 ;
        RECT 79.475 200.075 79.805 201.055 ;
        RECT 79.975 200.085 80.205 201.225 ;
        RECT 80.415 200.135 81.625 201.225 ;
        RECT 81.800 200.790 87.145 201.225 ;
        RECT 78.110 199.225 78.860 199.395 ;
        RECT 78.105 198.675 78.435 199.055 ;
        RECT 78.605 198.935 78.860 199.225 ;
        RECT 79.095 198.675 79.305 199.495 ;
        RECT 79.475 199.475 79.725 200.075 ;
        RECT 79.895 199.665 80.225 199.915 ;
        RECT 80.415 199.595 80.935 200.135 ;
        RECT 79.475 198.845 79.805 199.475 ;
        RECT 79.975 198.675 80.205 199.495 ;
        RECT 81.105 199.425 81.625 199.965 ;
        RECT 83.390 199.540 83.740 200.790 ;
        RECT 87.315 200.060 87.605 201.225 ;
        RECT 88.235 200.135 89.905 201.225 ;
        RECT 90.080 200.790 95.425 201.225 ;
        RECT 95.600 200.790 100.945 201.225 ;
        RECT 101.120 200.790 106.465 201.225 ;
        RECT 106.640 200.790 111.985 201.225 ;
        RECT 80.415 198.675 81.625 199.425 ;
        RECT 85.220 199.220 85.560 200.050 ;
        RECT 88.235 199.615 88.985 200.135 ;
        RECT 89.155 199.445 89.905 199.965 ;
        RECT 91.670 199.540 92.020 200.790 ;
        RECT 81.800 198.675 87.145 199.220 ;
        RECT 87.315 198.675 87.605 199.400 ;
        RECT 88.235 198.675 89.905 199.445 ;
        RECT 93.500 199.220 93.840 200.050 ;
        RECT 97.190 199.540 97.540 200.790 ;
        RECT 99.020 199.220 99.360 200.050 ;
        RECT 102.710 199.540 103.060 200.790 ;
        RECT 104.540 199.220 104.880 200.050 ;
        RECT 108.230 199.540 108.580 200.790 ;
        RECT 112.155 200.135 113.365 201.225 ;
        RECT 110.060 199.220 110.400 200.050 ;
        RECT 112.155 199.595 112.675 200.135 ;
        RECT 112.845 199.425 113.365 199.965 ;
        RECT 90.080 198.675 95.425 199.220 ;
        RECT 95.600 198.675 100.945 199.220 ;
        RECT 101.120 198.675 106.465 199.220 ;
        RECT 106.640 198.675 111.985 199.220 ;
        RECT 112.155 198.675 113.365 199.425 ;
        RECT 15.010 198.505 113.450 198.675 ;
        RECT 15.095 197.755 16.305 198.505 ;
        RECT 17.400 197.960 22.745 198.505 ;
        RECT 15.095 197.215 15.615 197.755 ;
        RECT 15.785 197.045 16.305 197.585 ;
        RECT 15.095 195.955 16.305 197.045 ;
        RECT 18.990 196.390 19.340 197.640 ;
        RECT 20.820 197.130 21.160 197.960 ;
        RECT 22.915 197.780 23.205 198.505 ;
        RECT 23.835 197.735 26.425 198.505 ;
        RECT 26.600 197.960 31.945 198.505 ;
        RECT 32.120 197.960 37.465 198.505 ;
        RECT 37.640 197.960 42.985 198.505 ;
        RECT 43.160 197.960 48.505 198.505 ;
        RECT 17.400 195.955 22.745 196.390 ;
        RECT 22.915 195.955 23.205 197.120 ;
        RECT 23.835 197.045 25.045 197.565 ;
        RECT 25.215 197.215 26.425 197.735 ;
        RECT 23.835 195.955 26.425 197.045 ;
        RECT 28.190 196.390 28.540 197.640 ;
        RECT 30.020 197.130 30.360 197.960 ;
        RECT 33.710 196.390 34.060 197.640 ;
        RECT 35.540 197.130 35.880 197.960 ;
        RECT 39.230 196.390 39.580 197.640 ;
        RECT 41.060 197.130 41.400 197.960 ;
        RECT 44.750 196.390 45.100 197.640 ;
        RECT 46.580 197.130 46.920 197.960 ;
        RECT 48.675 197.780 48.965 198.505 ;
        RECT 49.135 197.735 51.725 198.505 ;
        RECT 52.205 198.035 52.375 198.505 ;
        RECT 52.545 197.855 52.875 198.335 ;
        RECT 53.045 198.035 53.215 198.505 ;
        RECT 53.385 197.855 53.715 198.335 ;
        RECT 26.600 195.955 31.945 196.390 ;
        RECT 32.120 195.955 37.465 196.390 ;
        RECT 37.640 195.955 42.985 196.390 ;
        RECT 43.160 195.955 48.505 196.390 ;
        RECT 48.675 195.955 48.965 197.120 ;
        RECT 49.135 197.045 50.345 197.565 ;
        RECT 50.515 197.215 51.725 197.735 ;
        RECT 51.950 197.685 53.715 197.855 ;
        RECT 53.885 197.695 54.055 198.505 ;
        RECT 54.255 198.125 55.325 198.295 ;
        RECT 54.255 197.770 54.575 198.125 ;
        RECT 51.950 197.135 52.360 197.685 ;
        RECT 54.250 197.515 54.575 197.770 ;
        RECT 52.545 197.305 54.575 197.515 ;
        RECT 54.230 197.295 54.575 197.305 ;
        RECT 54.745 197.555 54.985 197.955 ;
        RECT 55.155 197.895 55.325 198.125 ;
        RECT 55.495 198.065 55.685 198.505 ;
        RECT 55.855 198.055 56.805 198.335 ;
        RECT 57.025 198.145 57.375 198.315 ;
        RECT 55.155 197.725 55.685 197.895 ;
        RECT 49.135 195.955 51.725 197.045 ;
        RECT 51.950 196.965 53.675 197.135 ;
        RECT 52.205 195.955 52.375 196.795 ;
        RECT 52.585 196.125 52.835 196.965 ;
        RECT 53.045 195.955 53.215 196.795 ;
        RECT 53.385 196.125 53.675 196.965 ;
        RECT 53.885 195.955 54.055 197.015 ;
        RECT 54.230 196.675 54.400 197.295 ;
        RECT 54.745 197.185 55.285 197.555 ;
        RECT 55.465 197.445 55.685 197.725 ;
        RECT 55.855 197.275 56.025 198.055 ;
        RECT 55.620 197.105 56.025 197.275 ;
        RECT 56.195 197.265 56.545 197.885 ;
        RECT 55.620 197.015 55.790 197.105 ;
        RECT 56.715 197.095 56.925 197.885 ;
        RECT 54.570 196.845 55.790 197.015 ;
        RECT 56.250 196.935 56.925 197.095 ;
        RECT 54.230 196.505 55.030 196.675 ;
        RECT 54.350 195.955 54.680 196.335 ;
        RECT 54.860 196.215 55.030 196.505 ;
        RECT 55.620 196.465 55.790 196.845 ;
        RECT 55.960 196.925 56.925 196.935 ;
        RECT 57.115 197.755 57.375 198.145 ;
        RECT 57.585 198.045 57.915 198.505 ;
        RECT 58.790 198.115 59.645 198.285 ;
        RECT 59.850 198.115 60.345 198.285 ;
        RECT 60.515 198.145 60.845 198.505 ;
        RECT 57.115 197.065 57.285 197.755 ;
        RECT 57.455 197.405 57.625 197.585 ;
        RECT 57.795 197.575 58.585 197.825 ;
        RECT 58.790 197.405 58.960 198.115 ;
        RECT 59.130 197.605 59.485 197.825 ;
        RECT 57.455 197.235 59.145 197.405 ;
        RECT 55.960 196.635 56.420 196.925 ;
        RECT 57.115 196.895 58.615 197.065 ;
        RECT 57.115 196.755 57.285 196.895 ;
        RECT 56.725 196.585 57.285 196.755 ;
        RECT 55.200 195.955 55.450 196.415 ;
        RECT 55.620 196.125 56.490 196.465 ;
        RECT 56.725 196.125 56.895 196.585 ;
        RECT 57.730 196.555 58.805 196.725 ;
        RECT 57.065 195.955 57.435 196.415 ;
        RECT 57.730 196.215 57.900 196.555 ;
        RECT 58.070 195.955 58.400 196.385 ;
        RECT 58.635 196.215 58.805 196.555 ;
        RECT 58.975 196.455 59.145 197.235 ;
        RECT 59.315 197.015 59.485 197.605 ;
        RECT 59.655 197.205 60.005 197.825 ;
        RECT 59.315 196.625 59.780 197.015 ;
        RECT 60.175 196.755 60.345 198.115 ;
        RECT 60.515 196.925 60.975 197.975 ;
        RECT 59.950 196.585 60.345 196.755 ;
        RECT 59.950 196.455 60.120 196.585 ;
        RECT 58.975 196.125 59.655 196.455 ;
        RECT 59.870 196.125 60.120 196.455 ;
        RECT 60.290 195.955 60.540 196.415 ;
        RECT 60.710 196.140 61.035 196.925 ;
        RECT 61.205 196.125 61.375 198.245 ;
        RECT 61.545 198.125 61.875 198.505 ;
        RECT 62.045 197.955 62.300 198.245 ;
        RECT 61.550 197.785 62.300 197.955 ;
        RECT 61.550 196.795 61.780 197.785 ;
        RECT 62.940 197.765 63.275 198.505 ;
        RECT 61.950 196.965 62.300 197.615 ;
        RECT 63.445 197.595 63.660 198.290 ;
        RECT 63.850 197.765 64.200 198.290 ;
        RECT 64.370 197.765 65.065 198.335 ;
        RECT 65.240 197.795 65.495 198.325 ;
        RECT 65.665 198.045 65.970 198.505 ;
        RECT 66.215 198.125 67.285 198.295 ;
        RECT 63.995 197.595 64.200 197.765 ;
        RECT 62.960 197.265 63.245 197.595 ;
        RECT 63.445 197.265 63.825 197.595 ;
        RECT 63.995 197.265 64.305 197.595 ;
        RECT 64.475 197.095 64.645 197.765 ;
        RECT 61.550 196.625 62.300 196.795 ;
        RECT 61.545 195.955 61.875 196.455 ;
        RECT 62.045 196.125 62.300 196.625 ;
        RECT 62.935 195.955 63.195 197.095 ;
        RECT 63.365 196.925 64.645 197.095 ;
        RECT 64.825 196.925 65.065 197.595 ;
        RECT 65.240 197.145 65.450 197.795 ;
        RECT 66.215 197.770 66.535 198.125 ;
        RECT 66.210 197.595 66.535 197.770 ;
        RECT 65.620 197.295 66.535 197.595 ;
        RECT 66.705 197.555 66.945 197.955 ;
        RECT 67.115 197.895 67.285 198.125 ;
        RECT 67.455 198.065 67.645 198.505 ;
        RECT 67.815 198.055 68.765 198.335 ;
        RECT 68.985 198.145 69.335 198.315 ;
        RECT 67.115 197.725 67.645 197.895 ;
        RECT 65.620 197.265 66.360 197.295 ;
        RECT 63.365 196.125 63.695 196.925 ;
        RECT 63.865 195.955 64.035 196.755 ;
        RECT 64.235 196.125 64.565 196.925 ;
        RECT 64.765 195.955 65.045 196.755 ;
        RECT 65.240 196.265 65.495 197.145 ;
        RECT 65.665 195.955 65.970 197.095 ;
        RECT 66.190 196.675 66.360 197.265 ;
        RECT 66.705 197.185 67.245 197.555 ;
        RECT 67.425 197.445 67.645 197.725 ;
        RECT 67.815 197.275 67.985 198.055 ;
        RECT 67.580 197.105 67.985 197.275 ;
        RECT 68.155 197.265 68.505 197.885 ;
        RECT 67.580 197.015 67.750 197.105 ;
        RECT 68.675 197.095 68.885 197.885 ;
        RECT 66.530 196.845 67.750 197.015 ;
        RECT 68.210 196.935 68.885 197.095 ;
        RECT 66.190 196.505 66.990 196.675 ;
        RECT 66.310 195.955 66.640 196.335 ;
        RECT 66.820 196.215 66.990 196.505 ;
        RECT 67.580 196.465 67.750 196.845 ;
        RECT 67.920 196.925 68.885 196.935 ;
        RECT 69.075 197.755 69.335 198.145 ;
        RECT 69.545 198.045 69.875 198.505 ;
        RECT 70.750 198.115 71.605 198.285 ;
        RECT 71.810 198.115 72.305 198.285 ;
        RECT 72.475 198.145 72.805 198.505 ;
        RECT 69.075 197.065 69.245 197.755 ;
        RECT 69.415 197.405 69.585 197.585 ;
        RECT 69.755 197.575 70.545 197.825 ;
        RECT 70.750 197.405 70.920 198.115 ;
        RECT 71.090 197.605 71.445 197.825 ;
        RECT 69.415 197.235 71.105 197.405 ;
        RECT 67.920 196.635 68.380 196.925 ;
        RECT 69.075 196.895 70.575 197.065 ;
        RECT 69.075 196.755 69.245 196.895 ;
        RECT 68.685 196.585 69.245 196.755 ;
        RECT 67.160 195.955 67.410 196.415 ;
        RECT 67.580 196.125 68.450 196.465 ;
        RECT 68.685 196.125 68.855 196.585 ;
        RECT 69.690 196.555 70.765 196.725 ;
        RECT 69.025 195.955 69.395 196.415 ;
        RECT 69.690 196.215 69.860 196.555 ;
        RECT 70.030 195.955 70.360 196.385 ;
        RECT 70.595 196.215 70.765 196.555 ;
        RECT 70.935 196.455 71.105 197.235 ;
        RECT 71.275 197.015 71.445 197.605 ;
        RECT 71.615 197.205 71.965 197.825 ;
        RECT 71.275 196.625 71.740 197.015 ;
        RECT 72.135 196.755 72.305 198.115 ;
        RECT 72.475 196.925 72.935 197.975 ;
        RECT 71.910 196.585 72.305 196.755 ;
        RECT 71.910 196.455 72.080 196.585 ;
        RECT 70.935 196.125 71.615 196.455 ;
        RECT 71.830 196.125 72.080 196.455 ;
        RECT 72.250 195.955 72.500 196.415 ;
        RECT 72.670 196.140 72.995 196.925 ;
        RECT 73.165 196.125 73.335 198.245 ;
        RECT 73.505 198.125 73.835 198.505 ;
        RECT 74.005 197.955 74.260 198.245 ;
        RECT 73.510 197.785 74.260 197.955 ;
        RECT 73.510 196.795 73.740 197.785 ;
        RECT 74.435 197.780 74.725 198.505 ;
        RECT 74.900 197.795 75.155 198.325 ;
        RECT 75.325 198.045 75.630 198.505 ;
        RECT 75.875 198.125 76.945 198.295 ;
        RECT 73.910 196.965 74.260 197.615 ;
        RECT 74.900 197.145 75.110 197.795 ;
        RECT 75.875 197.770 76.195 198.125 ;
        RECT 75.870 197.595 76.195 197.770 ;
        RECT 75.280 197.295 76.195 197.595 ;
        RECT 76.365 197.555 76.605 197.955 ;
        RECT 76.775 197.895 76.945 198.125 ;
        RECT 77.115 198.065 77.305 198.505 ;
        RECT 77.475 198.055 78.425 198.335 ;
        RECT 78.645 198.145 78.995 198.315 ;
        RECT 76.775 197.725 77.305 197.895 ;
        RECT 75.280 197.265 76.020 197.295 ;
        RECT 73.510 196.625 74.260 196.795 ;
        RECT 73.505 195.955 73.835 196.455 ;
        RECT 74.005 196.125 74.260 196.625 ;
        RECT 74.435 195.955 74.725 197.120 ;
        RECT 74.900 196.265 75.155 197.145 ;
        RECT 75.325 195.955 75.630 197.095 ;
        RECT 75.850 196.675 76.020 197.265 ;
        RECT 76.365 197.185 76.905 197.555 ;
        RECT 77.085 197.445 77.305 197.725 ;
        RECT 77.475 197.275 77.645 198.055 ;
        RECT 77.240 197.105 77.645 197.275 ;
        RECT 77.815 197.265 78.165 197.885 ;
        RECT 77.240 197.015 77.410 197.105 ;
        RECT 78.335 197.095 78.545 197.885 ;
        RECT 76.190 196.845 77.410 197.015 ;
        RECT 77.870 196.935 78.545 197.095 ;
        RECT 75.850 196.505 76.650 196.675 ;
        RECT 75.970 195.955 76.300 196.335 ;
        RECT 76.480 196.215 76.650 196.505 ;
        RECT 77.240 196.465 77.410 196.845 ;
        RECT 77.580 196.925 78.545 196.935 ;
        RECT 78.735 197.755 78.995 198.145 ;
        RECT 79.205 198.045 79.535 198.505 ;
        RECT 80.410 198.115 81.265 198.285 ;
        RECT 81.470 198.115 81.965 198.285 ;
        RECT 82.135 198.145 82.465 198.505 ;
        RECT 78.735 197.065 78.905 197.755 ;
        RECT 79.075 197.405 79.245 197.585 ;
        RECT 79.415 197.575 80.205 197.825 ;
        RECT 80.410 197.405 80.580 198.115 ;
        RECT 80.750 197.605 81.105 197.825 ;
        RECT 79.075 197.235 80.765 197.405 ;
        RECT 77.580 196.635 78.040 196.925 ;
        RECT 78.735 196.895 80.235 197.065 ;
        RECT 78.735 196.755 78.905 196.895 ;
        RECT 78.345 196.585 78.905 196.755 ;
        RECT 76.820 195.955 77.070 196.415 ;
        RECT 77.240 196.125 78.110 196.465 ;
        RECT 78.345 196.125 78.515 196.585 ;
        RECT 79.350 196.555 80.425 196.725 ;
        RECT 78.685 195.955 79.055 196.415 ;
        RECT 79.350 196.215 79.520 196.555 ;
        RECT 79.690 195.955 80.020 196.385 ;
        RECT 80.255 196.215 80.425 196.555 ;
        RECT 80.595 196.455 80.765 197.235 ;
        RECT 80.935 197.015 81.105 197.605 ;
        RECT 81.275 197.205 81.625 197.825 ;
        RECT 80.935 196.625 81.400 197.015 ;
        RECT 81.795 196.755 81.965 198.115 ;
        RECT 82.135 196.925 82.595 197.975 ;
        RECT 81.570 196.585 81.965 196.755 ;
        RECT 81.570 196.455 81.740 196.585 ;
        RECT 80.595 196.125 81.275 196.455 ;
        RECT 81.490 196.125 81.740 196.455 ;
        RECT 81.910 195.955 82.160 196.415 ;
        RECT 82.330 196.140 82.655 196.925 ;
        RECT 82.825 196.125 82.995 198.245 ;
        RECT 83.165 198.125 83.495 198.505 ;
        RECT 83.665 197.955 83.920 198.245 ;
        RECT 83.170 197.785 83.920 197.955 ;
        RECT 83.170 196.795 83.400 197.785 ;
        RECT 84.095 197.755 85.305 198.505 ;
        RECT 83.570 196.965 83.920 197.615 ;
        RECT 84.095 197.045 84.615 197.585 ;
        RECT 84.785 197.215 85.305 197.755 ;
        RECT 85.475 197.735 88.985 198.505 ;
        RECT 89.160 197.960 94.505 198.505 ;
        RECT 85.475 197.045 87.165 197.565 ;
        RECT 87.335 197.215 88.985 197.735 ;
        RECT 83.170 196.625 83.920 196.795 ;
        RECT 83.165 195.955 83.495 196.455 ;
        RECT 83.665 196.125 83.920 196.625 ;
        RECT 84.095 195.955 85.305 197.045 ;
        RECT 85.475 195.955 88.985 197.045 ;
        RECT 90.750 196.390 91.100 197.640 ;
        RECT 92.580 197.130 92.920 197.960 ;
        RECT 94.790 197.875 95.075 198.335 ;
        RECT 95.245 198.045 95.515 198.505 ;
        RECT 94.790 197.705 95.745 197.875 ;
        RECT 94.675 196.975 95.365 197.535 ;
        RECT 95.535 196.805 95.745 197.705 ;
        RECT 94.790 196.585 95.745 196.805 ;
        RECT 95.915 197.535 96.315 198.335 ;
        RECT 96.505 197.875 96.785 198.335 ;
        RECT 97.305 198.045 97.630 198.505 ;
        RECT 96.505 197.705 97.630 197.875 ;
        RECT 97.800 197.765 98.185 198.335 ;
        RECT 97.180 197.595 97.630 197.705 ;
        RECT 95.915 196.975 97.010 197.535 ;
        RECT 97.180 197.265 97.735 197.595 ;
        RECT 89.160 195.955 94.505 196.390 ;
        RECT 94.790 196.125 95.075 196.585 ;
        RECT 95.245 195.955 95.515 196.415 ;
        RECT 95.915 196.125 96.315 196.975 ;
        RECT 97.180 196.805 97.630 197.265 ;
        RECT 97.905 197.095 98.185 197.765 ;
        RECT 98.355 197.735 100.025 198.505 ;
        RECT 100.195 197.780 100.485 198.505 ;
        RECT 101.120 197.960 106.465 198.505 ;
        RECT 106.640 197.960 111.985 198.505 ;
        RECT 96.505 196.585 97.630 196.805 ;
        RECT 96.505 196.125 96.785 196.585 ;
        RECT 97.305 195.955 97.630 196.415 ;
        RECT 97.800 196.125 98.185 197.095 ;
        RECT 98.355 197.045 99.105 197.565 ;
        RECT 99.275 197.215 100.025 197.735 ;
        RECT 98.355 195.955 100.025 197.045 ;
        RECT 100.195 195.955 100.485 197.120 ;
        RECT 102.710 196.390 103.060 197.640 ;
        RECT 104.540 197.130 104.880 197.960 ;
        RECT 108.230 196.390 108.580 197.640 ;
        RECT 110.060 197.130 110.400 197.960 ;
        RECT 112.155 197.755 113.365 198.505 ;
        RECT 112.155 197.045 112.675 197.585 ;
        RECT 112.845 197.215 113.365 197.755 ;
        RECT 101.120 195.955 106.465 196.390 ;
        RECT 106.640 195.955 111.985 196.390 ;
        RECT 112.155 195.955 113.365 197.045 ;
        RECT 15.010 195.785 113.450 195.955 ;
        RECT 15.095 194.695 16.305 195.785 ;
        RECT 15.095 193.985 15.615 194.525 ;
        RECT 15.785 194.155 16.305 194.695 ;
        RECT 16.475 194.695 19.065 195.785 ;
        RECT 19.240 195.350 24.585 195.785 ;
        RECT 24.760 195.350 30.105 195.785 ;
        RECT 30.280 195.350 35.625 195.785 ;
        RECT 16.475 194.175 17.685 194.695 ;
        RECT 17.855 194.005 19.065 194.525 ;
        RECT 20.830 194.100 21.180 195.350 ;
        RECT 15.095 193.235 16.305 193.985 ;
        RECT 16.475 193.235 19.065 194.005 ;
        RECT 22.660 193.780 23.000 194.610 ;
        RECT 26.350 194.100 26.700 195.350 ;
        RECT 28.180 193.780 28.520 194.610 ;
        RECT 31.870 194.100 32.220 195.350 ;
        RECT 35.795 194.620 36.085 195.785 ;
        RECT 37.175 194.695 40.685 195.785 ;
        RECT 40.860 195.350 46.205 195.785 ;
        RECT 46.380 195.350 51.725 195.785 ;
        RECT 33.700 193.780 34.040 194.610 ;
        RECT 37.175 194.175 38.865 194.695 ;
        RECT 39.035 194.005 40.685 194.525 ;
        RECT 42.450 194.100 42.800 195.350 ;
        RECT 19.240 193.235 24.585 193.780 ;
        RECT 24.760 193.235 30.105 193.780 ;
        RECT 30.280 193.235 35.625 193.780 ;
        RECT 35.795 193.235 36.085 193.960 ;
        RECT 37.175 193.235 40.685 194.005 ;
        RECT 44.280 193.780 44.620 194.610 ;
        RECT 47.970 194.100 48.320 195.350 ;
        RECT 51.955 194.645 52.165 195.785 ;
        RECT 52.335 194.635 52.665 195.615 ;
        RECT 52.835 194.645 53.065 195.785 ;
        RECT 53.315 194.645 53.545 195.785 ;
        RECT 53.715 194.635 54.045 195.615 ;
        RECT 54.215 194.645 54.425 195.785 ;
        RECT 54.655 194.645 54.915 195.785 ;
        RECT 55.155 195.275 56.770 195.605 ;
        RECT 49.800 193.780 50.140 194.610 ;
        RECT 40.860 193.235 46.205 193.780 ;
        RECT 46.380 193.235 51.725 193.780 ;
        RECT 51.955 193.235 52.165 194.055 ;
        RECT 52.335 194.035 52.585 194.635 ;
        RECT 52.755 194.225 53.085 194.475 ;
        RECT 53.295 194.225 53.625 194.475 ;
        RECT 52.335 193.405 52.665 194.035 ;
        RECT 52.835 193.235 53.065 194.055 ;
        RECT 53.315 193.235 53.545 194.055 ;
        RECT 53.795 194.035 54.045 194.635 ;
        RECT 55.165 194.475 55.335 195.035 ;
        RECT 55.595 194.935 56.770 195.105 ;
        RECT 56.940 194.985 57.220 195.785 ;
        RECT 55.595 194.645 55.925 194.935 ;
        RECT 56.600 194.815 56.770 194.935 ;
        RECT 56.095 194.475 56.340 194.765 ;
        RECT 56.600 194.645 57.260 194.815 ;
        RECT 57.430 194.645 57.705 195.615 ;
        RECT 57.990 195.155 58.275 195.615 ;
        RECT 58.445 195.325 58.715 195.785 ;
        RECT 57.990 194.935 58.945 195.155 ;
        RECT 57.090 194.475 57.260 194.645 ;
        RECT 54.660 194.225 54.995 194.475 ;
        RECT 55.165 194.145 55.880 194.475 ;
        RECT 56.095 194.145 56.920 194.475 ;
        RECT 57.090 194.145 57.365 194.475 ;
        RECT 55.165 194.055 55.415 194.145 ;
        RECT 53.715 193.405 54.045 194.035 ;
        RECT 54.215 193.235 54.425 194.055 ;
        RECT 54.655 193.235 54.915 194.055 ;
        RECT 55.085 193.635 55.415 194.055 ;
        RECT 57.090 193.975 57.260 194.145 ;
        RECT 55.595 193.805 57.260 193.975 ;
        RECT 57.535 193.910 57.705 194.645 ;
        RECT 57.875 194.205 58.565 194.765 ;
        RECT 58.735 194.035 58.945 194.935 ;
        RECT 55.595 193.405 55.855 193.805 ;
        RECT 56.025 193.235 56.355 193.635 ;
        RECT 56.525 193.455 56.695 193.805 ;
        RECT 56.865 193.235 57.240 193.635 ;
        RECT 57.430 193.565 57.705 193.910 ;
        RECT 57.990 193.865 58.945 194.035 ;
        RECT 59.115 194.765 59.515 195.615 ;
        RECT 59.705 195.155 59.985 195.615 ;
        RECT 60.505 195.325 60.830 195.785 ;
        RECT 59.705 194.935 60.830 195.155 ;
        RECT 59.115 194.205 60.210 194.765 ;
        RECT 60.380 194.475 60.830 194.935 ;
        RECT 61.000 194.645 61.385 195.615 ;
        RECT 57.990 193.405 58.275 193.865 ;
        RECT 58.445 193.235 58.715 193.695 ;
        RECT 59.115 193.405 59.515 194.205 ;
        RECT 60.380 194.145 60.935 194.475 ;
        RECT 60.380 194.035 60.830 194.145 ;
        RECT 59.705 193.865 60.830 194.035 ;
        RECT 61.105 193.975 61.385 194.645 ;
        RECT 61.555 194.620 61.845 195.785 ;
        RECT 62.315 195.145 62.645 195.575 ;
        RECT 62.190 194.975 62.645 195.145 ;
        RECT 62.825 195.145 63.075 195.565 ;
        RECT 63.305 195.315 63.635 195.785 ;
        RECT 63.865 195.145 64.115 195.565 ;
        RECT 62.825 194.975 64.115 195.145 ;
        RECT 59.705 193.405 59.985 193.865 ;
        RECT 60.505 193.235 60.830 193.695 ;
        RECT 61.000 193.405 61.385 193.975 ;
        RECT 62.190 193.975 62.360 194.975 ;
        RECT 62.530 194.145 62.775 194.805 ;
        RECT 62.990 194.145 63.255 194.805 ;
        RECT 63.450 194.145 63.735 194.805 ;
        RECT 63.910 194.475 64.125 194.805 ;
        RECT 64.305 194.645 64.555 195.785 ;
        RECT 64.725 194.725 65.055 195.575 ;
        RECT 65.320 195.165 65.495 195.615 ;
        RECT 65.665 195.345 65.995 195.785 ;
        RECT 66.300 195.195 66.470 195.615 ;
        RECT 66.705 195.375 67.375 195.785 ;
        RECT 67.590 195.195 67.760 195.615 ;
        RECT 67.960 195.375 68.290 195.785 ;
        RECT 65.320 194.995 65.950 195.165 ;
        RECT 63.910 194.145 64.215 194.475 ;
        RECT 64.385 194.145 64.695 194.475 ;
        RECT 64.385 193.975 64.555 194.145 ;
        RECT 61.555 193.235 61.845 193.960 ;
        RECT 62.190 193.805 64.555 193.975 ;
        RECT 64.865 193.960 65.055 194.725 ;
        RECT 65.235 194.145 65.600 194.825 ;
        RECT 65.780 194.475 65.950 194.995 ;
        RECT 66.300 195.025 68.315 195.195 ;
        RECT 65.780 194.145 66.130 194.475 ;
        RECT 65.780 193.975 65.950 194.145 ;
        RECT 62.345 193.235 62.675 193.635 ;
        RECT 62.845 193.465 63.175 193.805 ;
        RECT 64.225 193.235 64.555 193.635 ;
        RECT 64.725 193.450 65.055 193.960 ;
        RECT 65.320 193.805 65.950 193.975 ;
        RECT 65.320 193.405 65.495 193.805 ;
        RECT 66.300 193.735 66.470 195.025 ;
        RECT 65.665 193.235 65.995 193.615 ;
        RECT 66.240 193.405 66.470 193.735 ;
        RECT 66.670 193.570 66.950 194.845 ;
        RECT 67.175 194.085 67.445 194.845 ;
        RECT 67.135 193.915 67.445 194.085 ;
        RECT 67.175 193.570 67.445 193.915 ;
        RECT 67.635 193.815 67.975 194.845 ;
        RECT 68.145 194.475 68.315 195.025 ;
        RECT 68.485 194.645 68.745 195.615 ;
        RECT 69.560 194.815 69.950 194.990 ;
        RECT 70.435 194.985 70.765 195.785 ;
        RECT 70.935 194.995 71.470 195.615 ;
        RECT 69.560 194.645 70.985 194.815 ;
        RECT 68.145 194.145 68.405 194.475 ;
        RECT 68.575 193.955 68.745 194.645 ;
        RECT 67.905 193.235 68.235 193.615 ;
        RECT 68.405 193.490 68.745 193.955 ;
        RECT 69.435 193.915 69.790 194.475 ;
        RECT 69.960 193.745 70.130 194.645 ;
        RECT 70.300 193.915 70.565 194.475 ;
        RECT 70.815 194.145 70.985 194.645 ;
        RECT 71.155 193.975 71.470 194.995 ;
        RECT 71.790 195.155 72.075 195.615 ;
        RECT 72.245 195.325 72.515 195.785 ;
        RECT 71.790 194.935 72.745 195.155 ;
        RECT 71.675 194.205 72.365 194.765 ;
        RECT 72.535 194.035 72.745 194.935 ;
        RECT 68.405 193.445 68.740 193.490 ;
        RECT 69.540 193.235 69.780 193.745 ;
        RECT 69.960 193.415 70.240 193.745 ;
        RECT 70.470 193.235 70.685 193.745 ;
        RECT 70.855 193.405 71.470 193.975 ;
        RECT 71.790 193.865 72.745 194.035 ;
        RECT 72.915 194.765 73.315 195.615 ;
        RECT 73.505 195.155 73.785 195.615 ;
        RECT 74.305 195.325 74.630 195.785 ;
        RECT 73.505 194.935 74.630 195.155 ;
        RECT 72.915 194.205 74.010 194.765 ;
        RECT 74.180 194.475 74.630 194.935 ;
        RECT 74.800 194.645 75.185 195.615 ;
        RECT 75.375 195.275 75.675 195.785 ;
        RECT 75.845 195.275 76.225 195.445 ;
        RECT 76.805 195.275 77.435 195.785 ;
        RECT 75.845 195.105 76.015 195.275 ;
        RECT 77.605 195.105 77.935 195.615 ;
        RECT 78.105 195.275 78.405 195.785 ;
        RECT 71.790 193.405 72.075 193.865 ;
        RECT 72.245 193.235 72.515 193.695 ;
        RECT 72.915 193.405 73.315 194.205 ;
        RECT 74.180 194.145 74.735 194.475 ;
        RECT 74.180 194.035 74.630 194.145 ;
        RECT 73.505 193.865 74.630 194.035 ;
        RECT 74.905 193.975 75.185 194.645 ;
        RECT 73.505 193.405 73.785 193.865 ;
        RECT 74.305 193.235 74.630 193.695 ;
        RECT 74.800 193.405 75.185 193.975 ;
        RECT 75.355 194.905 76.015 195.105 ;
        RECT 76.185 194.935 78.405 195.105 ;
        RECT 75.355 193.975 75.525 194.905 ;
        RECT 76.185 194.735 76.355 194.935 ;
        RECT 75.695 194.565 76.355 194.735 ;
        RECT 76.525 194.595 78.065 194.765 ;
        RECT 75.695 194.145 75.865 194.565 ;
        RECT 76.525 194.395 76.695 194.595 ;
        RECT 76.095 194.225 76.695 194.395 ;
        RECT 76.865 194.225 77.560 194.425 ;
        RECT 77.820 194.145 78.065 194.595 ;
        RECT 76.185 193.975 77.095 194.055 ;
        RECT 75.355 193.495 75.675 193.975 ;
        RECT 75.845 193.885 77.095 193.975 ;
        RECT 75.845 193.805 76.355 193.885 ;
        RECT 75.845 193.405 76.075 193.805 ;
        RECT 76.245 193.235 76.595 193.625 ;
        RECT 76.765 193.405 77.095 193.885 ;
        RECT 77.265 193.235 77.435 194.055 ;
        RECT 78.235 193.975 78.405 194.935 ;
        RECT 77.940 193.430 78.405 193.975 ;
        RECT 78.575 194.710 78.845 195.615 ;
        RECT 79.015 195.025 79.345 195.785 ;
        RECT 79.525 194.855 79.695 195.615 ;
        RECT 78.575 193.910 78.745 194.710 ;
        RECT 79.030 194.685 79.695 194.855 ;
        RECT 79.030 194.540 79.200 194.685 ;
        RECT 79.995 194.645 80.225 195.785 ;
        RECT 80.395 194.635 80.725 195.615 ;
        RECT 80.895 194.645 81.105 195.785 ;
        RECT 82.255 194.695 85.765 195.785 ;
        RECT 78.915 194.210 79.200 194.540 ;
        RECT 79.030 193.955 79.200 194.210 ;
        RECT 79.435 194.135 79.765 194.505 ;
        RECT 79.975 194.225 80.305 194.475 ;
        RECT 78.575 193.405 78.835 193.910 ;
        RECT 79.030 193.785 79.695 193.955 ;
        RECT 79.015 193.235 79.345 193.615 ;
        RECT 79.525 193.405 79.695 193.785 ;
        RECT 79.995 193.235 80.225 194.055 ;
        RECT 80.475 194.035 80.725 194.635 ;
        RECT 82.255 194.175 83.945 194.695 ;
        RECT 85.975 194.645 86.205 195.785 ;
        RECT 86.375 194.635 86.705 195.615 ;
        RECT 86.875 194.645 87.085 195.785 ;
        RECT 80.395 193.405 80.725 194.035 ;
        RECT 80.895 193.235 81.105 194.055 ;
        RECT 84.115 194.005 85.765 194.525 ;
        RECT 85.955 194.225 86.285 194.475 ;
        RECT 82.255 193.235 85.765 194.005 ;
        RECT 85.975 193.235 86.205 194.055 ;
        RECT 86.455 194.035 86.705 194.635 ;
        RECT 87.315 194.620 87.605 195.785 ;
        RECT 88.350 195.155 88.635 195.615 ;
        RECT 88.805 195.325 89.075 195.785 ;
        RECT 88.350 194.935 89.305 195.155 ;
        RECT 88.235 194.205 88.925 194.765 ;
        RECT 86.375 193.405 86.705 194.035 ;
        RECT 86.875 193.235 87.085 194.055 ;
        RECT 89.095 194.035 89.305 194.935 ;
        RECT 87.315 193.235 87.605 193.960 ;
        RECT 88.350 193.865 89.305 194.035 ;
        RECT 89.475 194.765 89.875 195.615 ;
        RECT 90.065 195.155 90.345 195.615 ;
        RECT 90.865 195.325 91.190 195.785 ;
        RECT 90.065 194.935 91.190 195.155 ;
        RECT 89.475 194.205 90.570 194.765 ;
        RECT 90.740 194.475 91.190 194.935 ;
        RECT 91.360 194.645 91.745 195.615 ;
        RECT 92.005 194.855 92.175 195.615 ;
        RECT 92.355 195.025 92.685 195.785 ;
        RECT 92.005 194.685 92.670 194.855 ;
        RECT 92.855 194.710 93.125 195.615 ;
        RECT 88.350 193.405 88.635 193.865 ;
        RECT 88.805 193.235 89.075 193.695 ;
        RECT 89.475 193.405 89.875 194.205 ;
        RECT 90.740 194.145 91.295 194.475 ;
        RECT 90.740 194.035 91.190 194.145 ;
        RECT 90.065 193.865 91.190 194.035 ;
        RECT 91.465 193.975 91.745 194.645 ;
        RECT 92.500 194.540 92.670 194.685 ;
        RECT 91.935 194.135 92.265 194.505 ;
        RECT 92.500 194.210 92.785 194.540 ;
        RECT 90.065 193.405 90.345 193.865 ;
        RECT 90.865 193.235 91.190 193.695 ;
        RECT 91.360 193.405 91.745 193.975 ;
        RECT 92.500 193.955 92.670 194.210 ;
        RECT 92.005 193.785 92.670 193.955 ;
        RECT 92.955 193.910 93.125 194.710 ;
        RECT 93.795 194.645 94.025 195.785 ;
        RECT 94.195 194.635 94.525 195.615 ;
        RECT 94.695 194.645 94.905 195.785 ;
        RECT 93.775 194.225 94.105 194.475 ;
        RECT 92.005 193.405 92.175 193.785 ;
        RECT 92.355 193.235 92.685 193.615 ;
        RECT 92.865 193.405 93.125 193.910 ;
        RECT 93.795 193.235 94.025 194.055 ;
        RECT 94.275 194.035 94.525 194.635 ;
        RECT 95.140 194.595 95.395 195.475 ;
        RECT 95.565 194.645 95.870 195.785 ;
        RECT 96.210 195.405 96.540 195.785 ;
        RECT 96.720 195.235 96.890 195.525 ;
        RECT 97.060 195.325 97.310 195.785 ;
        RECT 96.090 195.065 96.890 195.235 ;
        RECT 97.480 195.275 98.350 195.615 ;
        RECT 94.195 193.405 94.525 194.035 ;
        RECT 94.695 193.235 94.905 194.055 ;
        RECT 95.140 193.945 95.350 194.595 ;
        RECT 96.090 194.475 96.260 195.065 ;
        RECT 97.480 194.895 97.650 195.275 ;
        RECT 98.585 195.155 98.755 195.615 ;
        RECT 98.925 195.325 99.295 195.785 ;
        RECT 99.590 195.185 99.760 195.525 ;
        RECT 99.930 195.355 100.260 195.785 ;
        RECT 100.495 195.185 100.665 195.525 ;
        RECT 96.430 194.725 97.650 194.895 ;
        RECT 97.820 194.815 98.280 195.105 ;
        RECT 98.585 194.985 99.145 195.155 ;
        RECT 99.590 195.015 100.665 195.185 ;
        RECT 100.835 195.285 101.515 195.615 ;
        RECT 101.730 195.285 101.980 195.615 ;
        RECT 102.150 195.325 102.400 195.785 ;
        RECT 98.975 194.845 99.145 194.985 ;
        RECT 97.820 194.805 98.785 194.815 ;
        RECT 97.480 194.635 97.650 194.725 ;
        RECT 98.110 194.645 98.785 194.805 ;
        RECT 95.520 194.445 96.260 194.475 ;
        RECT 95.520 194.145 96.435 194.445 ;
        RECT 96.110 193.970 96.435 194.145 ;
        RECT 95.140 193.415 95.395 193.945 ;
        RECT 95.565 193.235 95.870 193.695 ;
        RECT 96.115 193.615 96.435 193.970 ;
        RECT 96.605 194.185 97.145 194.555 ;
        RECT 97.480 194.465 97.885 194.635 ;
        RECT 96.605 193.785 96.845 194.185 ;
        RECT 97.325 194.015 97.545 194.295 ;
        RECT 97.015 193.845 97.545 194.015 ;
        RECT 97.015 193.615 97.185 193.845 ;
        RECT 97.715 193.685 97.885 194.465 ;
        RECT 98.055 193.855 98.405 194.475 ;
        RECT 98.575 193.855 98.785 194.645 ;
        RECT 98.975 194.675 100.475 194.845 ;
        RECT 98.975 193.985 99.145 194.675 ;
        RECT 100.835 194.505 101.005 195.285 ;
        RECT 101.810 195.155 101.980 195.285 ;
        RECT 99.315 194.335 101.005 194.505 ;
        RECT 101.175 194.725 101.640 195.115 ;
        RECT 101.810 194.985 102.205 195.155 ;
        RECT 99.315 194.155 99.485 194.335 ;
        RECT 96.115 193.445 97.185 193.615 ;
        RECT 97.355 193.235 97.545 193.675 ;
        RECT 97.715 193.405 98.665 193.685 ;
        RECT 98.975 193.595 99.235 193.985 ;
        RECT 99.655 193.915 100.445 194.165 ;
        RECT 98.885 193.425 99.235 193.595 ;
        RECT 99.445 193.235 99.775 193.695 ;
        RECT 100.650 193.625 100.820 194.335 ;
        RECT 101.175 194.135 101.345 194.725 ;
        RECT 100.990 193.915 101.345 194.135 ;
        RECT 101.515 193.915 101.865 194.535 ;
        RECT 102.035 193.625 102.205 194.985 ;
        RECT 102.570 194.815 102.895 195.600 ;
        RECT 102.375 193.765 102.835 194.815 ;
        RECT 100.650 193.455 101.505 193.625 ;
        RECT 101.710 193.455 102.205 193.625 ;
        RECT 102.375 193.235 102.705 193.595 ;
        RECT 103.065 193.495 103.235 195.615 ;
        RECT 103.405 195.285 103.735 195.785 ;
        RECT 103.905 195.115 104.160 195.615 ;
        RECT 103.410 194.945 104.160 195.115 ;
        RECT 103.410 193.955 103.640 194.945 ;
        RECT 103.810 194.125 104.160 194.775 ;
        RECT 104.795 194.695 106.465 195.785 ;
        RECT 106.640 195.350 111.985 195.785 ;
        RECT 104.795 194.175 105.545 194.695 ;
        RECT 105.715 194.005 106.465 194.525 ;
        RECT 108.230 194.100 108.580 195.350 ;
        RECT 112.155 194.695 113.365 195.785 ;
        RECT 103.410 193.785 104.160 193.955 ;
        RECT 103.405 193.235 103.735 193.615 ;
        RECT 103.905 193.495 104.160 193.785 ;
        RECT 104.795 193.235 106.465 194.005 ;
        RECT 110.060 193.780 110.400 194.610 ;
        RECT 112.155 194.155 112.675 194.695 ;
        RECT 112.845 193.985 113.365 194.525 ;
        RECT 106.640 193.235 111.985 193.780 ;
        RECT 112.155 193.235 113.365 193.985 ;
        RECT 15.010 193.065 113.450 193.235 ;
        RECT 15.095 192.315 16.305 193.065 ;
        RECT 17.400 192.520 22.745 193.065 ;
        RECT 15.095 191.775 15.615 192.315 ;
        RECT 15.785 191.605 16.305 192.145 ;
        RECT 15.095 190.515 16.305 191.605 ;
        RECT 18.990 190.950 19.340 192.200 ;
        RECT 20.820 191.690 21.160 192.520 ;
        RECT 22.915 192.340 23.205 193.065 ;
        RECT 23.375 192.295 25.045 193.065 ;
        RECT 25.220 192.520 30.565 193.065 ;
        RECT 30.740 192.520 36.085 193.065 ;
        RECT 36.260 192.520 41.605 193.065 ;
        RECT 17.400 190.515 22.745 190.950 ;
        RECT 22.915 190.515 23.205 191.680 ;
        RECT 23.375 191.605 24.125 192.125 ;
        RECT 24.295 191.775 25.045 192.295 ;
        RECT 23.375 190.515 25.045 191.605 ;
        RECT 26.810 190.950 27.160 192.200 ;
        RECT 28.640 191.690 28.980 192.520 ;
        RECT 32.330 190.950 32.680 192.200 ;
        RECT 34.160 191.690 34.500 192.520 ;
        RECT 37.850 190.950 38.200 192.200 ;
        RECT 39.680 191.690 40.020 192.520 ;
        RECT 41.890 192.435 42.175 192.895 ;
        RECT 42.345 192.605 42.615 193.065 ;
        RECT 41.890 192.265 42.845 192.435 ;
        RECT 41.775 191.535 42.465 192.095 ;
        RECT 42.635 191.365 42.845 192.265 ;
        RECT 41.890 191.145 42.845 191.365 ;
        RECT 43.015 192.095 43.415 192.895 ;
        RECT 43.605 192.435 43.885 192.895 ;
        RECT 44.405 192.605 44.730 193.065 ;
        RECT 43.605 192.265 44.730 192.435 ;
        RECT 44.900 192.325 45.285 192.895 ;
        RECT 44.280 192.155 44.730 192.265 ;
        RECT 43.015 191.535 44.110 192.095 ;
        RECT 44.280 191.825 44.835 192.155 ;
        RECT 25.220 190.515 30.565 190.950 ;
        RECT 30.740 190.515 36.085 190.950 ;
        RECT 36.260 190.515 41.605 190.950 ;
        RECT 41.890 190.685 42.175 191.145 ;
        RECT 42.345 190.515 42.615 190.975 ;
        RECT 43.015 190.685 43.415 191.535 ;
        RECT 44.280 191.365 44.730 191.825 ;
        RECT 45.005 191.655 45.285 192.325 ;
        RECT 45.455 192.295 47.125 193.065 ;
        RECT 43.605 191.145 44.730 191.365 ;
        RECT 43.605 190.685 43.885 191.145 ;
        RECT 44.405 190.515 44.730 190.975 ;
        RECT 44.900 190.685 45.285 191.655 ;
        RECT 45.455 191.605 46.205 192.125 ;
        RECT 46.375 191.775 47.125 192.295 ;
        RECT 47.355 192.245 47.565 193.065 ;
        RECT 47.735 192.265 48.065 192.895 ;
        RECT 47.735 191.665 47.985 192.265 ;
        RECT 48.235 192.245 48.465 193.065 ;
        RECT 48.675 192.340 48.965 193.065 ;
        RECT 49.600 192.520 54.945 193.065 ;
        RECT 55.120 192.520 60.465 193.065 ;
        RECT 48.155 191.825 48.485 192.075 ;
        RECT 45.455 190.515 47.125 191.605 ;
        RECT 47.355 190.515 47.565 191.655 ;
        RECT 47.735 190.685 48.065 191.665 ;
        RECT 48.235 190.515 48.465 191.655 ;
        RECT 48.675 190.515 48.965 191.680 ;
        RECT 51.190 190.950 51.540 192.200 ;
        RECT 53.020 191.690 53.360 192.520 ;
        RECT 56.710 190.950 57.060 192.200 ;
        RECT 58.540 191.690 58.880 192.520 ;
        RECT 60.640 192.225 60.900 193.065 ;
        RECT 61.075 192.320 61.330 192.895 ;
        RECT 61.500 192.685 61.830 193.065 ;
        RECT 62.045 192.515 62.215 192.895 ;
        RECT 61.500 192.345 62.215 192.515 ;
        RECT 49.600 190.515 54.945 190.950 ;
        RECT 55.120 190.515 60.465 190.950 ;
        RECT 60.640 190.515 60.900 191.665 ;
        RECT 61.075 191.590 61.245 192.320 ;
        RECT 61.500 192.155 61.670 192.345 ;
        RECT 62.475 192.245 62.735 193.065 ;
        RECT 62.905 192.245 63.235 192.665 ;
        RECT 63.415 192.495 63.675 192.895 ;
        RECT 63.845 192.665 64.175 193.065 ;
        RECT 64.345 192.495 64.515 192.845 ;
        RECT 64.685 192.665 65.060 193.065 ;
        RECT 63.415 192.325 65.080 192.495 ;
        RECT 65.250 192.390 65.525 192.735 ;
        RECT 61.415 191.825 61.670 192.155 ;
        RECT 61.500 191.615 61.670 191.825 ;
        RECT 61.950 191.795 62.305 192.165 ;
        RECT 62.985 192.155 63.235 192.245 ;
        RECT 64.910 192.155 65.080 192.325 ;
        RECT 62.480 191.825 62.815 192.075 ;
        RECT 62.985 191.825 63.700 192.155 ;
        RECT 63.915 191.825 64.740 192.155 ;
        RECT 64.910 191.825 65.185 192.155 ;
        RECT 61.075 190.685 61.330 191.590 ;
        RECT 61.500 191.445 62.215 191.615 ;
        RECT 61.500 190.515 61.830 191.275 ;
        RECT 62.045 190.685 62.215 191.445 ;
        RECT 62.475 190.515 62.735 191.655 ;
        RECT 62.985 191.265 63.155 191.825 ;
        RECT 63.415 191.365 63.745 191.655 ;
        RECT 63.915 191.535 64.160 191.825 ;
        RECT 64.910 191.655 65.080 191.825 ;
        RECT 65.355 191.655 65.525 192.390 ;
        RECT 64.420 191.485 65.080 191.655 ;
        RECT 64.420 191.365 64.590 191.485 ;
        RECT 63.415 191.195 64.590 191.365 ;
        RECT 62.975 190.695 64.590 191.025 ;
        RECT 64.760 190.515 65.040 191.315 ;
        RECT 65.250 190.685 65.525 191.655 ;
        RECT 65.695 192.565 65.955 192.895 ;
        RECT 66.265 192.685 66.595 193.065 ;
        RECT 66.775 192.725 68.255 192.895 ;
        RECT 65.695 191.865 65.865 192.565 ;
        RECT 66.775 192.395 67.175 192.725 ;
        RECT 66.215 192.205 66.425 192.385 ;
        RECT 66.215 192.035 66.835 192.205 ;
        RECT 67.005 191.915 67.175 192.395 ;
        RECT 67.365 192.225 67.915 192.555 ;
        RECT 65.695 191.695 66.825 191.865 ;
        RECT 67.005 191.745 67.575 191.915 ;
        RECT 65.695 191.015 65.865 191.695 ;
        RECT 66.655 191.575 66.825 191.695 ;
        RECT 66.035 191.195 66.385 191.525 ;
        RECT 66.655 191.405 67.235 191.575 ;
        RECT 67.405 191.235 67.575 191.745 ;
        RECT 66.835 191.065 67.575 191.235 ;
        RECT 67.745 191.235 67.915 192.225 ;
        RECT 68.085 191.825 68.255 192.725 ;
        RECT 68.505 192.155 68.690 192.735 ;
        RECT 68.960 192.155 69.155 192.730 ;
        RECT 69.365 192.685 69.695 193.065 ;
        RECT 68.505 191.825 68.735 192.155 ;
        RECT 68.960 191.825 69.215 192.155 ;
        RECT 68.505 191.515 68.690 191.825 ;
        RECT 68.960 191.515 69.155 191.825 ;
        RECT 69.525 191.235 69.695 192.155 ;
        RECT 67.745 191.065 69.695 191.235 ;
        RECT 65.695 190.685 65.955 191.015 ;
        RECT 66.265 190.515 66.595 190.895 ;
        RECT 66.835 190.685 67.025 191.065 ;
        RECT 67.275 190.515 67.605 190.895 ;
        RECT 67.815 190.685 67.985 191.065 ;
        RECT 68.180 190.515 68.510 190.895 ;
        RECT 68.770 190.685 68.940 191.065 ;
        RECT 69.365 190.515 69.695 190.895 ;
        RECT 69.865 190.685 70.125 192.895 ;
        RECT 70.295 192.685 71.185 192.855 ;
        RECT 70.295 192.130 70.845 192.515 ;
        RECT 71.015 191.960 71.185 192.685 ;
        RECT 70.295 191.890 71.185 191.960 ;
        RECT 71.355 192.360 71.575 192.845 ;
        RECT 71.745 192.525 71.995 193.065 ;
        RECT 72.165 192.415 72.425 192.895 ;
        RECT 71.355 191.935 71.685 192.360 ;
        RECT 70.295 191.865 71.190 191.890 ;
        RECT 70.295 191.850 71.200 191.865 ;
        RECT 70.295 191.835 71.205 191.850 ;
        RECT 70.295 191.830 71.215 191.835 ;
        RECT 70.295 191.820 71.220 191.830 ;
        RECT 70.295 191.810 71.225 191.820 ;
        RECT 70.295 191.805 71.235 191.810 ;
        RECT 70.295 191.795 71.245 191.805 ;
        RECT 70.295 191.790 71.255 191.795 ;
        RECT 70.295 191.340 70.555 191.790 ;
        RECT 70.920 191.785 71.255 191.790 ;
        RECT 70.920 191.780 71.270 191.785 ;
        RECT 70.920 191.770 71.285 191.780 ;
        RECT 70.920 191.765 71.310 191.770 ;
        RECT 71.855 191.765 72.085 192.160 ;
        RECT 70.920 191.760 72.085 191.765 ;
        RECT 70.950 191.725 72.085 191.760 ;
        RECT 70.985 191.700 72.085 191.725 ;
        RECT 71.015 191.670 72.085 191.700 ;
        RECT 71.035 191.640 72.085 191.670 ;
        RECT 71.055 191.610 72.085 191.640 ;
        RECT 71.125 191.600 72.085 191.610 ;
        RECT 71.150 191.590 72.085 191.600 ;
        RECT 71.170 191.575 72.085 191.590 ;
        RECT 71.190 191.560 72.085 191.575 ;
        RECT 71.195 191.550 71.980 191.560 ;
        RECT 71.210 191.515 71.980 191.550 ;
        RECT 70.725 191.195 71.055 191.440 ;
        RECT 71.225 191.265 71.980 191.515 ;
        RECT 72.255 191.385 72.425 192.415 ;
        RECT 72.595 192.265 73.290 192.895 ;
        RECT 73.495 192.265 73.805 193.065 ;
        RECT 74.435 192.340 74.725 193.065 ;
        RECT 75.355 192.565 75.615 192.895 ;
        RECT 75.825 192.585 76.100 193.065 ;
        RECT 72.615 191.825 72.950 192.075 ;
        RECT 73.120 191.665 73.290 192.265 ;
        RECT 73.460 191.825 73.795 192.095 ;
        RECT 70.725 191.170 70.910 191.195 ;
        RECT 70.295 191.070 70.910 191.170 ;
        RECT 70.295 190.515 70.900 191.070 ;
        RECT 71.075 190.685 71.555 191.025 ;
        RECT 71.725 190.515 71.980 191.060 ;
        RECT 72.150 190.685 72.425 191.385 ;
        RECT 72.595 190.515 72.855 191.655 ;
        RECT 73.025 190.685 73.355 191.665 ;
        RECT 73.525 190.515 73.805 191.655 ;
        RECT 74.435 190.515 74.725 191.680 ;
        RECT 75.355 191.655 75.525 192.565 ;
        RECT 76.310 192.495 76.515 192.895 ;
        RECT 76.685 192.665 77.020 193.065 ;
        RECT 75.695 191.825 76.055 192.405 ;
        RECT 76.310 192.325 76.995 192.495 ;
        RECT 76.235 191.655 76.485 192.155 ;
        RECT 75.355 191.485 76.485 191.655 ;
        RECT 75.355 190.715 75.625 191.485 ;
        RECT 76.655 191.295 76.995 192.325 ;
        RECT 77.195 192.295 78.865 193.065 ;
        RECT 79.040 192.520 84.385 193.065 ;
        RECT 75.795 190.515 76.125 191.295 ;
        RECT 76.330 191.120 76.995 191.295 ;
        RECT 77.195 191.605 77.945 192.125 ;
        RECT 78.115 191.775 78.865 192.295 ;
        RECT 76.330 190.715 76.515 191.120 ;
        RECT 76.685 190.515 77.020 190.940 ;
        RECT 77.195 190.515 78.865 191.605 ;
        RECT 80.630 190.950 80.980 192.200 ;
        RECT 82.460 191.690 82.800 192.520 ;
        RECT 84.645 192.515 84.815 192.895 ;
        RECT 84.995 192.685 85.325 193.065 ;
        RECT 84.645 192.345 85.310 192.515 ;
        RECT 85.505 192.390 85.765 192.895 ;
        RECT 84.575 191.795 84.905 192.165 ;
        RECT 85.140 192.090 85.310 192.345 ;
        RECT 85.140 191.760 85.425 192.090 ;
        RECT 85.140 191.615 85.310 191.760 ;
        RECT 84.645 191.445 85.310 191.615 ;
        RECT 85.595 191.590 85.765 192.390 ;
        RECT 79.040 190.515 84.385 190.950 ;
        RECT 84.645 190.685 84.815 191.445 ;
        RECT 84.995 190.515 85.325 191.275 ;
        RECT 85.495 190.685 85.765 191.590 ;
        RECT 85.940 192.355 86.195 192.885 ;
        RECT 86.365 192.605 86.670 193.065 ;
        RECT 86.915 192.685 87.985 192.855 ;
        RECT 85.940 191.705 86.150 192.355 ;
        RECT 86.915 192.330 87.235 192.685 ;
        RECT 86.910 192.155 87.235 192.330 ;
        RECT 86.320 191.855 87.235 192.155 ;
        RECT 87.405 192.115 87.645 192.515 ;
        RECT 87.815 192.455 87.985 192.685 ;
        RECT 88.155 192.625 88.345 193.065 ;
        RECT 88.515 192.615 89.465 192.895 ;
        RECT 89.685 192.705 90.035 192.875 ;
        RECT 87.815 192.285 88.345 192.455 ;
        RECT 86.320 191.825 87.060 191.855 ;
        RECT 85.940 190.825 86.195 191.705 ;
        RECT 86.365 190.515 86.670 191.655 ;
        RECT 86.890 191.235 87.060 191.825 ;
        RECT 87.405 191.745 87.945 192.115 ;
        RECT 88.125 192.005 88.345 192.285 ;
        RECT 88.515 191.835 88.685 192.615 ;
        RECT 88.280 191.665 88.685 191.835 ;
        RECT 88.855 191.825 89.205 192.445 ;
        RECT 88.280 191.575 88.450 191.665 ;
        RECT 89.375 191.655 89.585 192.445 ;
        RECT 87.230 191.405 88.450 191.575 ;
        RECT 88.910 191.495 89.585 191.655 ;
        RECT 86.890 191.065 87.690 191.235 ;
        RECT 87.010 190.515 87.340 190.895 ;
        RECT 87.520 190.775 87.690 191.065 ;
        RECT 88.280 191.025 88.450 191.405 ;
        RECT 88.620 191.485 89.585 191.495 ;
        RECT 89.775 192.315 90.035 192.705 ;
        RECT 90.245 192.605 90.575 193.065 ;
        RECT 91.450 192.675 92.305 192.845 ;
        RECT 92.510 192.675 93.005 192.845 ;
        RECT 93.175 192.705 93.505 193.065 ;
        RECT 89.775 191.625 89.945 192.315 ;
        RECT 90.115 191.965 90.285 192.145 ;
        RECT 90.455 192.135 91.245 192.385 ;
        RECT 91.450 191.965 91.620 192.675 ;
        RECT 91.790 192.165 92.145 192.385 ;
        RECT 90.115 191.795 91.805 191.965 ;
        RECT 88.620 191.195 89.080 191.485 ;
        RECT 89.775 191.455 91.275 191.625 ;
        RECT 89.775 191.315 89.945 191.455 ;
        RECT 89.385 191.145 89.945 191.315 ;
        RECT 87.860 190.515 88.110 190.975 ;
        RECT 88.280 190.685 89.150 191.025 ;
        RECT 89.385 190.685 89.555 191.145 ;
        RECT 90.390 191.115 91.465 191.285 ;
        RECT 89.725 190.515 90.095 190.975 ;
        RECT 90.390 190.775 90.560 191.115 ;
        RECT 90.730 190.515 91.060 190.945 ;
        RECT 91.295 190.775 91.465 191.115 ;
        RECT 91.635 191.015 91.805 191.795 ;
        RECT 91.975 191.575 92.145 192.165 ;
        RECT 92.315 191.765 92.665 192.385 ;
        RECT 91.975 191.185 92.440 191.575 ;
        RECT 92.835 191.315 93.005 192.675 ;
        RECT 93.175 191.485 93.635 192.535 ;
        RECT 92.610 191.145 93.005 191.315 ;
        RECT 92.610 191.015 92.780 191.145 ;
        RECT 91.635 190.685 92.315 191.015 ;
        RECT 92.530 190.685 92.780 191.015 ;
        RECT 92.950 190.515 93.200 190.975 ;
        RECT 93.370 190.700 93.695 191.485 ;
        RECT 93.865 190.685 94.035 192.805 ;
        RECT 94.205 192.685 94.535 193.065 ;
        RECT 94.705 192.515 94.960 192.805 ;
        RECT 94.210 192.345 94.960 192.515 ;
        RECT 94.210 191.355 94.440 192.345 ;
        RECT 96.330 192.255 96.575 192.860 ;
        RECT 96.795 192.530 97.305 193.065 ;
        RECT 94.610 191.525 94.960 192.175 ;
        RECT 96.055 192.085 97.285 192.255 ;
        RECT 94.210 191.185 94.960 191.355 ;
        RECT 94.205 190.515 94.535 191.015 ;
        RECT 94.705 190.685 94.960 191.185 ;
        RECT 96.055 191.275 96.395 192.085 ;
        RECT 96.565 191.520 97.315 191.710 ;
        RECT 96.055 190.865 96.570 191.275 ;
        RECT 96.805 190.515 96.975 191.275 ;
        RECT 97.145 190.855 97.315 191.520 ;
        RECT 97.485 191.535 97.675 192.895 ;
        RECT 97.845 192.725 98.120 192.895 ;
        RECT 97.845 192.555 98.125 192.725 ;
        RECT 97.845 191.735 98.120 192.555 ;
        RECT 98.310 192.530 98.840 192.895 ;
        RECT 99.265 192.665 99.595 193.065 ;
        RECT 98.665 192.495 98.840 192.530 ;
        RECT 98.325 191.535 98.495 192.335 ;
        RECT 97.485 191.365 98.495 191.535 ;
        RECT 98.665 192.325 99.595 192.495 ;
        RECT 99.765 192.325 100.020 192.895 ;
        RECT 100.195 192.340 100.485 193.065 ;
        RECT 100.660 192.355 100.915 192.885 ;
        RECT 101.085 192.605 101.390 193.065 ;
        RECT 101.635 192.685 102.705 192.855 ;
        RECT 98.665 191.195 98.835 192.325 ;
        RECT 99.425 192.155 99.595 192.325 ;
        RECT 97.710 191.025 98.835 191.195 ;
        RECT 99.005 191.825 99.200 192.155 ;
        RECT 99.425 191.825 99.680 192.155 ;
        RECT 99.005 190.855 99.175 191.825 ;
        RECT 99.850 191.655 100.020 192.325 ;
        RECT 100.660 191.705 100.870 192.355 ;
        RECT 101.635 192.330 101.955 192.685 ;
        RECT 101.630 192.155 101.955 192.330 ;
        RECT 101.040 191.855 101.955 192.155 ;
        RECT 102.125 192.115 102.365 192.515 ;
        RECT 102.535 192.455 102.705 192.685 ;
        RECT 102.875 192.625 103.065 193.065 ;
        RECT 103.235 192.615 104.185 192.895 ;
        RECT 104.405 192.705 104.755 192.875 ;
        RECT 102.535 192.285 103.065 192.455 ;
        RECT 101.040 191.825 101.780 191.855 ;
        RECT 97.145 190.685 99.175 190.855 ;
        RECT 99.345 190.515 99.515 191.655 ;
        RECT 99.685 190.685 100.020 191.655 ;
        RECT 100.195 190.515 100.485 191.680 ;
        RECT 100.660 190.825 100.915 191.705 ;
        RECT 101.085 190.515 101.390 191.655 ;
        RECT 101.610 191.235 101.780 191.825 ;
        RECT 102.125 191.745 102.665 192.115 ;
        RECT 102.845 192.005 103.065 192.285 ;
        RECT 103.235 191.835 103.405 192.615 ;
        RECT 103.000 191.665 103.405 191.835 ;
        RECT 103.575 191.825 103.925 192.445 ;
        RECT 103.000 191.575 103.170 191.665 ;
        RECT 104.095 191.655 104.305 192.445 ;
        RECT 101.950 191.405 103.170 191.575 ;
        RECT 103.630 191.495 104.305 191.655 ;
        RECT 101.610 191.065 102.410 191.235 ;
        RECT 101.730 190.515 102.060 190.895 ;
        RECT 102.240 190.775 102.410 191.065 ;
        RECT 103.000 191.025 103.170 191.405 ;
        RECT 103.340 191.485 104.305 191.495 ;
        RECT 104.495 192.315 104.755 192.705 ;
        RECT 104.965 192.605 105.295 193.065 ;
        RECT 106.170 192.675 107.025 192.845 ;
        RECT 107.230 192.675 107.725 192.845 ;
        RECT 107.895 192.705 108.225 193.065 ;
        RECT 104.495 191.625 104.665 192.315 ;
        RECT 104.835 191.965 105.005 192.145 ;
        RECT 105.175 192.135 105.965 192.385 ;
        RECT 106.170 191.965 106.340 192.675 ;
        RECT 106.510 192.165 106.865 192.385 ;
        RECT 104.835 191.795 106.525 191.965 ;
        RECT 103.340 191.195 103.800 191.485 ;
        RECT 104.495 191.455 105.995 191.625 ;
        RECT 104.495 191.315 104.665 191.455 ;
        RECT 104.105 191.145 104.665 191.315 ;
        RECT 102.580 190.515 102.830 190.975 ;
        RECT 103.000 190.685 103.870 191.025 ;
        RECT 104.105 190.685 104.275 191.145 ;
        RECT 105.110 191.115 106.185 191.285 ;
        RECT 104.445 190.515 104.815 190.975 ;
        RECT 105.110 190.775 105.280 191.115 ;
        RECT 105.450 190.515 105.780 190.945 ;
        RECT 106.015 190.775 106.185 191.115 ;
        RECT 106.355 191.015 106.525 191.795 ;
        RECT 106.695 191.575 106.865 192.165 ;
        RECT 107.035 191.765 107.385 192.385 ;
        RECT 106.695 191.185 107.160 191.575 ;
        RECT 107.555 191.315 107.725 192.675 ;
        RECT 107.895 191.485 108.355 192.535 ;
        RECT 107.330 191.145 107.725 191.315 ;
        RECT 107.330 191.015 107.500 191.145 ;
        RECT 106.355 190.685 107.035 191.015 ;
        RECT 107.250 190.685 107.500 191.015 ;
        RECT 107.670 190.515 107.920 190.975 ;
        RECT 108.090 190.700 108.415 191.485 ;
        RECT 108.585 190.685 108.755 192.805 ;
        RECT 108.925 192.685 109.255 193.065 ;
        RECT 109.425 192.515 109.680 192.805 ;
        RECT 108.930 192.345 109.680 192.515 ;
        RECT 108.930 191.355 109.160 192.345 ;
        RECT 110.315 192.295 111.985 193.065 ;
        RECT 112.155 192.315 113.365 193.065 ;
        RECT 109.330 191.525 109.680 192.175 ;
        RECT 110.315 191.605 111.065 192.125 ;
        RECT 111.235 191.775 111.985 192.295 ;
        RECT 112.155 191.605 112.675 192.145 ;
        RECT 112.845 191.775 113.365 192.315 ;
        RECT 108.930 191.185 109.680 191.355 ;
        RECT 108.925 190.515 109.255 191.015 ;
        RECT 109.425 190.685 109.680 191.185 ;
        RECT 110.315 190.515 111.985 191.605 ;
        RECT 112.155 190.515 113.365 191.605 ;
        RECT 15.010 190.345 113.450 190.515 ;
        RECT 15.095 189.255 16.305 190.345 ;
        RECT 15.095 188.545 15.615 189.085 ;
        RECT 15.785 188.715 16.305 189.255 ;
        RECT 16.475 189.255 17.685 190.345 ;
        RECT 17.860 189.910 23.205 190.345 ;
        RECT 23.380 189.910 28.725 190.345 ;
        RECT 28.900 189.910 34.245 190.345 ;
        RECT 16.475 188.715 16.995 189.255 ;
        RECT 17.165 188.545 17.685 189.085 ;
        RECT 19.450 188.660 19.800 189.910 ;
        RECT 15.095 187.795 16.305 188.545 ;
        RECT 16.475 187.795 17.685 188.545 ;
        RECT 21.280 188.340 21.620 189.170 ;
        RECT 24.970 188.660 25.320 189.910 ;
        RECT 26.800 188.340 27.140 189.170 ;
        RECT 30.490 188.660 30.840 189.910 ;
        RECT 34.455 189.205 34.685 190.345 ;
        RECT 34.855 189.195 35.185 190.175 ;
        RECT 35.355 189.205 35.565 190.345 ;
        RECT 32.320 188.340 32.660 189.170 ;
        RECT 34.435 188.785 34.765 189.035 ;
        RECT 17.860 187.795 23.205 188.340 ;
        RECT 23.380 187.795 28.725 188.340 ;
        RECT 28.900 187.795 34.245 188.340 ;
        RECT 34.455 187.795 34.685 188.615 ;
        RECT 34.935 188.595 35.185 189.195 ;
        RECT 35.795 189.180 36.085 190.345 ;
        RECT 36.715 189.255 38.385 190.345 ;
        RECT 38.645 189.415 38.815 190.175 ;
        RECT 38.995 189.585 39.325 190.345 ;
        RECT 36.715 188.735 37.465 189.255 ;
        RECT 38.645 189.245 39.310 189.415 ;
        RECT 39.495 189.270 39.765 190.175 ;
        RECT 39.140 189.100 39.310 189.245 ;
        RECT 34.855 187.965 35.185 188.595 ;
        RECT 35.355 187.795 35.565 188.615 ;
        RECT 37.635 188.565 38.385 189.085 ;
        RECT 38.575 188.695 38.905 189.065 ;
        RECT 39.140 188.770 39.425 189.100 ;
        RECT 35.795 187.795 36.085 188.520 ;
        RECT 36.715 187.795 38.385 188.565 ;
        RECT 39.140 188.515 39.310 188.770 ;
        RECT 38.645 188.345 39.310 188.515 ;
        RECT 39.595 188.470 39.765 189.270 ;
        RECT 39.935 189.585 40.450 189.995 ;
        RECT 40.685 189.585 40.855 190.345 ;
        RECT 41.025 190.005 43.055 190.175 ;
        RECT 39.935 188.775 40.275 189.585 ;
        RECT 41.025 189.340 41.195 190.005 ;
        RECT 41.590 189.665 42.715 189.835 ;
        RECT 40.445 189.150 41.195 189.340 ;
        RECT 41.365 189.325 42.375 189.495 ;
        RECT 39.935 188.605 41.165 188.775 ;
        RECT 38.645 187.965 38.815 188.345 ;
        RECT 38.995 187.795 39.325 188.175 ;
        RECT 39.505 187.965 39.765 188.470 ;
        RECT 40.210 188.000 40.455 188.605 ;
        RECT 40.675 187.795 41.185 188.330 ;
        RECT 41.365 187.965 41.555 189.325 ;
        RECT 41.725 188.305 42.000 189.125 ;
        RECT 42.205 188.525 42.375 189.325 ;
        RECT 42.545 188.535 42.715 189.665 ;
        RECT 42.885 189.035 43.055 190.005 ;
        RECT 43.225 189.205 43.395 190.345 ;
        RECT 43.565 189.205 43.900 190.175 ;
        RECT 42.885 188.705 43.080 189.035 ;
        RECT 43.305 188.705 43.560 189.035 ;
        RECT 43.305 188.535 43.475 188.705 ;
        RECT 43.730 188.535 43.900 189.205 ;
        RECT 42.545 188.365 43.475 188.535 ;
        RECT 42.545 188.330 42.720 188.365 ;
        RECT 41.725 188.135 42.005 188.305 ;
        RECT 41.725 187.965 42.000 188.135 ;
        RECT 42.190 187.965 42.720 188.330 ;
        RECT 43.145 187.795 43.475 188.195 ;
        RECT 43.645 187.965 43.900 188.535 ;
        RECT 44.080 189.155 44.335 190.035 ;
        RECT 44.505 189.205 44.810 190.345 ;
        RECT 45.150 189.965 45.480 190.345 ;
        RECT 45.660 189.795 45.830 190.085 ;
        RECT 46.000 189.885 46.250 190.345 ;
        RECT 45.030 189.625 45.830 189.795 ;
        RECT 46.420 189.835 47.290 190.175 ;
        RECT 44.080 188.505 44.290 189.155 ;
        RECT 45.030 189.035 45.200 189.625 ;
        RECT 46.420 189.455 46.590 189.835 ;
        RECT 47.525 189.715 47.695 190.175 ;
        RECT 47.865 189.885 48.235 190.345 ;
        RECT 48.530 189.745 48.700 190.085 ;
        RECT 48.870 189.915 49.200 190.345 ;
        RECT 49.435 189.745 49.605 190.085 ;
        RECT 45.370 189.285 46.590 189.455 ;
        RECT 46.760 189.375 47.220 189.665 ;
        RECT 47.525 189.545 48.085 189.715 ;
        RECT 48.530 189.575 49.605 189.745 ;
        RECT 49.775 189.845 50.455 190.175 ;
        RECT 50.670 189.845 50.920 190.175 ;
        RECT 51.090 189.885 51.340 190.345 ;
        RECT 47.915 189.405 48.085 189.545 ;
        RECT 46.760 189.365 47.725 189.375 ;
        RECT 46.420 189.195 46.590 189.285 ;
        RECT 47.050 189.205 47.725 189.365 ;
        RECT 44.460 189.005 45.200 189.035 ;
        RECT 44.460 188.705 45.375 189.005 ;
        RECT 45.050 188.530 45.375 188.705 ;
        RECT 44.080 187.975 44.335 188.505 ;
        RECT 44.505 187.795 44.810 188.255 ;
        RECT 45.055 188.175 45.375 188.530 ;
        RECT 45.545 188.745 46.085 189.115 ;
        RECT 46.420 189.025 46.825 189.195 ;
        RECT 45.545 188.345 45.785 188.745 ;
        RECT 46.265 188.575 46.485 188.855 ;
        RECT 45.955 188.405 46.485 188.575 ;
        RECT 45.955 188.175 46.125 188.405 ;
        RECT 46.655 188.245 46.825 189.025 ;
        RECT 46.995 188.415 47.345 189.035 ;
        RECT 47.515 188.415 47.725 189.205 ;
        RECT 47.915 189.235 49.415 189.405 ;
        RECT 47.915 188.545 48.085 189.235 ;
        RECT 49.775 189.065 49.945 189.845 ;
        RECT 50.750 189.715 50.920 189.845 ;
        RECT 48.255 188.895 49.945 189.065 ;
        RECT 50.115 189.285 50.580 189.675 ;
        RECT 50.750 189.545 51.145 189.715 ;
        RECT 48.255 188.715 48.425 188.895 ;
        RECT 45.055 188.005 46.125 188.175 ;
        RECT 46.295 187.795 46.485 188.235 ;
        RECT 46.655 187.965 47.605 188.245 ;
        RECT 47.915 188.155 48.175 188.545 ;
        RECT 48.595 188.475 49.385 188.725 ;
        RECT 47.825 187.985 48.175 188.155 ;
        RECT 48.385 187.795 48.715 188.255 ;
        RECT 49.590 188.185 49.760 188.895 ;
        RECT 50.115 188.695 50.285 189.285 ;
        RECT 49.930 188.475 50.285 188.695 ;
        RECT 50.455 188.475 50.805 189.095 ;
        RECT 50.975 188.185 51.145 189.545 ;
        RECT 51.510 189.375 51.835 190.160 ;
        RECT 51.315 188.325 51.775 189.375 ;
        RECT 49.590 188.015 50.445 188.185 ;
        RECT 50.650 188.015 51.145 188.185 ;
        RECT 51.315 187.795 51.645 188.155 ;
        RECT 52.005 188.055 52.175 190.175 ;
        RECT 52.345 189.845 52.675 190.345 ;
        RECT 52.845 189.675 53.100 190.175 ;
        RECT 52.350 189.505 53.100 189.675 ;
        RECT 52.350 188.515 52.580 189.505 ;
        RECT 52.750 188.685 53.100 189.335 ;
        RECT 53.275 189.255 54.485 190.345 ;
        RECT 54.745 189.415 54.915 190.175 ;
        RECT 55.095 189.585 55.425 190.345 ;
        RECT 53.275 188.715 53.795 189.255 ;
        RECT 54.745 189.245 55.410 189.415 ;
        RECT 55.595 189.270 55.865 190.175 ;
        RECT 56.040 189.910 61.385 190.345 ;
        RECT 55.240 189.100 55.410 189.245 ;
        RECT 53.965 188.545 54.485 189.085 ;
        RECT 54.675 188.695 55.005 189.065 ;
        RECT 55.240 188.770 55.525 189.100 ;
        RECT 52.350 188.345 53.100 188.515 ;
        RECT 52.345 187.795 52.675 188.175 ;
        RECT 52.845 188.055 53.100 188.345 ;
        RECT 53.275 187.795 54.485 188.545 ;
        RECT 55.240 188.515 55.410 188.770 ;
        RECT 54.745 188.345 55.410 188.515 ;
        RECT 55.695 188.470 55.865 189.270 ;
        RECT 57.630 188.660 57.980 189.910 ;
        RECT 61.555 189.180 61.845 190.345 ;
        RECT 62.935 189.255 66.445 190.345 ;
        RECT 66.620 189.920 66.955 190.345 ;
        RECT 67.125 189.740 67.310 190.145 ;
        RECT 66.645 189.565 67.310 189.740 ;
        RECT 67.515 189.565 67.845 190.345 ;
        RECT 54.745 187.965 54.915 188.345 ;
        RECT 55.095 187.795 55.425 188.175 ;
        RECT 55.605 187.965 55.865 188.470 ;
        RECT 59.460 188.340 59.800 189.170 ;
        RECT 62.935 188.735 64.625 189.255 ;
        RECT 64.795 188.565 66.445 189.085 ;
        RECT 56.040 187.795 61.385 188.340 ;
        RECT 61.555 187.795 61.845 188.520 ;
        RECT 62.935 187.795 66.445 188.565 ;
        RECT 66.645 188.535 66.985 189.565 ;
        RECT 68.015 189.375 68.285 190.145 ;
        RECT 67.155 189.205 68.285 189.375 ;
        RECT 67.155 188.705 67.405 189.205 ;
        RECT 66.645 188.365 67.330 188.535 ;
        RECT 67.585 188.455 67.945 189.035 ;
        RECT 66.620 187.795 66.955 188.195 ;
        RECT 67.125 187.965 67.330 188.365 ;
        RECT 68.115 188.295 68.285 189.205 ;
        RECT 68.455 189.255 71.965 190.345 ;
        RECT 72.140 189.910 77.485 190.345 ;
        RECT 68.455 188.735 70.145 189.255 ;
        RECT 70.315 188.565 71.965 189.085 ;
        RECT 73.730 188.660 74.080 189.910 ;
        RECT 78.030 189.365 78.285 190.035 ;
        RECT 78.465 189.545 78.750 190.345 ;
        RECT 78.930 189.625 79.260 190.135 ;
        RECT 67.540 187.795 67.815 188.275 ;
        RECT 68.025 187.965 68.285 188.295 ;
        RECT 68.455 187.795 71.965 188.565 ;
        RECT 75.560 188.340 75.900 189.170 ;
        RECT 78.030 188.505 78.210 189.365 ;
        RECT 78.930 189.035 79.180 189.625 ;
        RECT 79.530 189.475 79.700 190.085 ;
        RECT 79.870 189.655 80.200 190.345 ;
        RECT 80.430 189.795 80.670 190.085 ;
        RECT 80.870 189.965 81.290 190.345 ;
        RECT 81.470 189.875 82.100 190.125 ;
        RECT 82.570 189.965 82.900 190.345 ;
        RECT 81.470 189.795 81.640 189.875 ;
        RECT 83.070 189.795 83.240 190.085 ;
        RECT 83.420 189.965 83.800 190.345 ;
        RECT 84.040 189.960 84.870 190.130 ;
        RECT 80.430 189.625 81.640 189.795 ;
        RECT 78.380 188.705 79.180 189.035 ;
        RECT 72.140 187.795 77.485 188.340 ;
        RECT 78.030 188.305 78.285 188.505 ;
        RECT 77.945 188.135 78.285 188.305 ;
        RECT 78.030 187.975 78.285 188.135 ;
        RECT 78.465 187.795 78.750 188.255 ;
        RECT 78.930 188.055 79.180 188.705 ;
        RECT 79.380 189.455 79.700 189.475 ;
        RECT 79.380 189.285 81.300 189.455 ;
        RECT 79.380 188.390 79.570 189.285 ;
        RECT 81.470 189.115 81.640 189.625 ;
        RECT 81.810 189.365 82.330 189.675 ;
        RECT 79.740 188.945 81.640 189.115 ;
        RECT 79.740 188.885 80.070 188.945 ;
        RECT 80.220 188.715 80.550 188.775 ;
        RECT 79.890 188.445 80.550 188.715 ;
        RECT 79.380 188.060 79.700 188.390 ;
        RECT 79.880 187.795 80.540 188.275 ;
        RECT 80.740 188.185 80.910 188.945 ;
        RECT 81.810 188.775 81.990 189.185 ;
        RECT 81.080 188.605 81.410 188.725 ;
        RECT 82.160 188.605 82.330 189.365 ;
        RECT 81.080 188.435 82.330 188.605 ;
        RECT 82.500 189.545 83.870 189.795 ;
        RECT 82.500 188.775 82.690 189.545 ;
        RECT 83.620 189.285 83.870 189.545 ;
        RECT 82.860 189.115 83.110 189.275 ;
        RECT 84.040 189.115 84.210 189.960 ;
        RECT 85.105 189.675 85.275 190.175 ;
        RECT 85.445 189.845 85.775 190.345 ;
        RECT 84.380 189.285 84.880 189.665 ;
        RECT 85.105 189.505 85.800 189.675 ;
        RECT 82.860 188.945 84.210 189.115 ;
        RECT 83.790 188.905 84.210 188.945 ;
        RECT 82.500 188.435 82.920 188.775 ;
        RECT 83.210 188.445 83.620 188.775 ;
        RECT 80.740 188.015 81.590 188.185 ;
        RECT 82.150 187.795 82.470 188.255 ;
        RECT 82.670 188.005 82.920 188.435 ;
        RECT 83.210 187.795 83.620 188.235 ;
        RECT 83.790 188.175 83.960 188.905 ;
        RECT 84.130 188.355 84.480 188.725 ;
        RECT 84.660 188.415 84.880 189.285 ;
        RECT 85.050 188.715 85.460 189.335 ;
        RECT 85.630 188.535 85.800 189.505 ;
        RECT 85.105 188.345 85.800 188.535 ;
        RECT 83.790 187.975 84.805 188.175 ;
        RECT 85.105 188.015 85.275 188.345 ;
        RECT 85.445 187.795 85.775 188.175 ;
        RECT 85.990 188.055 86.215 190.175 ;
        RECT 86.385 189.845 86.715 190.345 ;
        RECT 86.885 189.675 87.055 190.175 ;
        RECT 86.390 189.505 87.055 189.675 ;
        RECT 86.390 188.515 86.620 189.505 ;
        RECT 86.790 188.685 87.140 189.335 ;
        RECT 87.315 189.180 87.605 190.345 ;
        RECT 87.775 189.585 88.290 189.995 ;
        RECT 88.525 189.585 88.695 190.345 ;
        RECT 88.865 190.005 90.895 190.175 ;
        RECT 87.775 188.775 88.115 189.585 ;
        RECT 88.865 189.340 89.035 190.005 ;
        RECT 89.430 189.665 90.555 189.835 ;
        RECT 88.285 189.150 89.035 189.340 ;
        RECT 89.205 189.325 90.215 189.495 ;
        RECT 87.775 188.605 89.005 188.775 ;
        RECT 86.390 188.345 87.055 188.515 ;
        RECT 86.385 187.795 86.715 188.175 ;
        RECT 86.885 188.055 87.055 188.345 ;
        RECT 87.315 187.795 87.605 188.520 ;
        RECT 88.050 188.000 88.295 188.605 ;
        RECT 88.515 187.795 89.025 188.330 ;
        RECT 89.205 187.965 89.395 189.325 ;
        RECT 89.565 188.305 89.840 189.125 ;
        RECT 90.045 188.525 90.215 189.325 ;
        RECT 90.385 188.535 90.555 189.665 ;
        RECT 90.725 189.035 90.895 190.005 ;
        RECT 91.065 189.205 91.235 190.345 ;
        RECT 91.405 189.205 91.740 190.175 ;
        RECT 90.725 188.705 90.920 189.035 ;
        RECT 91.145 188.705 91.400 189.035 ;
        RECT 91.145 188.535 91.315 188.705 ;
        RECT 91.570 188.535 91.740 189.205 ;
        RECT 91.915 189.255 93.585 190.345 ;
        RECT 91.915 188.735 92.665 189.255 ;
        RECT 93.755 189.205 94.140 190.175 ;
        RECT 94.310 189.885 94.635 190.345 ;
        RECT 95.155 189.715 95.435 190.175 ;
        RECT 94.310 189.495 95.435 189.715 ;
        RECT 92.835 188.565 93.585 189.085 ;
        RECT 90.385 188.365 91.315 188.535 ;
        RECT 90.385 188.330 90.560 188.365 ;
        RECT 89.565 188.135 89.845 188.305 ;
        RECT 89.565 187.965 89.840 188.135 ;
        RECT 90.030 187.965 90.560 188.330 ;
        RECT 90.985 187.795 91.315 188.195 ;
        RECT 91.485 187.965 91.740 188.535 ;
        RECT 91.915 187.795 93.585 188.565 ;
        RECT 93.755 188.535 94.035 189.205 ;
        RECT 94.310 189.035 94.760 189.495 ;
        RECT 95.625 189.325 96.025 190.175 ;
        RECT 96.425 189.885 96.695 190.345 ;
        RECT 96.865 189.715 97.150 190.175 ;
        RECT 94.205 188.705 94.760 189.035 ;
        RECT 94.930 188.765 96.025 189.325 ;
        RECT 94.310 188.595 94.760 188.705 ;
        RECT 93.755 187.965 94.140 188.535 ;
        RECT 94.310 188.425 95.435 188.595 ;
        RECT 94.310 187.795 94.635 188.255 ;
        RECT 95.155 187.965 95.435 188.425 ;
        RECT 95.625 187.965 96.025 188.765 ;
        RECT 96.195 189.495 97.150 189.715 ;
        RECT 96.195 188.595 96.405 189.495 ;
        RECT 97.985 189.415 98.155 190.175 ;
        RECT 98.335 189.585 98.665 190.345 ;
        RECT 96.575 188.765 97.265 189.325 ;
        RECT 97.985 189.245 98.650 189.415 ;
        RECT 98.835 189.270 99.105 190.175 ;
        RECT 98.480 189.100 98.650 189.245 ;
        RECT 97.915 188.695 98.245 189.065 ;
        RECT 98.480 188.770 98.765 189.100 ;
        RECT 96.195 188.425 97.150 188.595 ;
        RECT 98.480 188.515 98.650 188.770 ;
        RECT 96.425 187.795 96.695 188.255 ;
        RECT 96.865 187.965 97.150 188.425 ;
        RECT 97.985 188.345 98.650 188.515 ;
        RECT 98.935 188.470 99.105 189.270 ;
        RECT 99.275 189.585 99.790 189.995 ;
        RECT 100.025 189.585 100.195 190.345 ;
        RECT 100.365 190.005 102.395 190.175 ;
        RECT 99.275 188.775 99.615 189.585 ;
        RECT 100.365 189.340 100.535 190.005 ;
        RECT 100.930 189.665 102.055 189.835 ;
        RECT 99.785 189.150 100.535 189.340 ;
        RECT 100.705 189.325 101.715 189.495 ;
        RECT 99.275 188.605 100.505 188.775 ;
        RECT 97.985 187.965 98.155 188.345 ;
        RECT 98.335 187.795 98.665 188.175 ;
        RECT 98.845 187.965 99.105 188.470 ;
        RECT 99.550 188.000 99.795 188.605 ;
        RECT 100.015 187.795 100.525 188.330 ;
        RECT 100.705 187.965 100.895 189.325 ;
        RECT 101.065 188.305 101.340 189.125 ;
        RECT 101.545 188.525 101.715 189.325 ;
        RECT 101.885 188.535 102.055 189.665 ;
        RECT 102.225 189.035 102.395 190.005 ;
        RECT 102.565 189.205 102.735 190.345 ;
        RECT 102.905 189.205 103.240 190.175 ;
        RECT 102.225 188.705 102.420 189.035 ;
        RECT 102.645 188.705 102.900 189.035 ;
        RECT 102.645 188.535 102.815 188.705 ;
        RECT 103.070 188.535 103.240 189.205 ;
        RECT 101.885 188.365 102.815 188.535 ;
        RECT 101.885 188.330 102.060 188.365 ;
        RECT 101.065 188.135 101.345 188.305 ;
        RECT 101.065 187.965 101.340 188.135 ;
        RECT 101.530 187.965 102.060 188.330 ;
        RECT 102.485 187.795 102.815 188.195 ;
        RECT 102.985 187.965 103.240 188.535 ;
        RECT 103.415 189.205 103.800 190.175 ;
        RECT 103.970 189.885 104.295 190.345 ;
        RECT 104.815 189.715 105.095 190.175 ;
        RECT 103.970 189.495 105.095 189.715 ;
        RECT 103.415 188.535 103.695 189.205 ;
        RECT 103.970 189.035 104.420 189.495 ;
        RECT 105.285 189.325 105.685 190.175 ;
        RECT 106.085 189.885 106.355 190.345 ;
        RECT 106.525 189.715 106.810 190.175 ;
        RECT 103.865 188.705 104.420 189.035 ;
        RECT 104.590 188.765 105.685 189.325 ;
        RECT 103.970 188.595 104.420 188.705 ;
        RECT 103.415 187.965 103.800 188.535 ;
        RECT 103.970 188.425 105.095 188.595 ;
        RECT 103.970 187.795 104.295 188.255 ;
        RECT 104.815 187.965 105.095 188.425 ;
        RECT 105.285 187.965 105.685 188.765 ;
        RECT 105.855 189.495 106.810 189.715 ;
        RECT 105.855 188.595 106.065 189.495 ;
        RECT 106.235 188.765 106.925 189.325 ;
        RECT 107.155 189.205 107.365 190.345 ;
        RECT 107.535 189.195 107.865 190.175 ;
        RECT 108.035 189.205 108.265 190.345 ;
        RECT 108.475 189.270 108.745 190.175 ;
        RECT 108.915 189.585 109.245 190.345 ;
        RECT 109.425 189.415 109.595 190.175 ;
        RECT 105.855 188.425 106.810 188.595 ;
        RECT 106.085 187.795 106.355 188.255 ;
        RECT 106.525 187.965 106.810 188.425 ;
        RECT 107.155 187.795 107.365 188.615 ;
        RECT 107.535 188.595 107.785 189.195 ;
        RECT 107.955 188.785 108.285 189.035 ;
        RECT 107.535 187.965 107.865 188.595 ;
        RECT 108.035 187.795 108.265 188.615 ;
        RECT 108.475 188.470 108.645 189.270 ;
        RECT 108.930 189.245 109.595 189.415 ;
        RECT 110.315 189.255 111.985 190.345 ;
        RECT 112.155 189.255 113.365 190.345 ;
        RECT 108.930 189.100 109.100 189.245 ;
        RECT 108.815 188.770 109.100 189.100 ;
        RECT 108.930 188.515 109.100 188.770 ;
        RECT 109.335 188.695 109.665 189.065 ;
        RECT 110.315 188.735 111.065 189.255 ;
        RECT 111.235 188.565 111.985 189.085 ;
        RECT 112.155 188.715 112.675 189.255 ;
        RECT 108.475 187.965 108.735 188.470 ;
        RECT 108.930 188.345 109.595 188.515 ;
        RECT 108.915 187.795 109.245 188.175 ;
        RECT 109.425 187.965 109.595 188.345 ;
        RECT 110.315 187.795 111.985 188.565 ;
        RECT 112.845 188.545 113.365 189.085 ;
        RECT 112.155 187.795 113.365 188.545 ;
        RECT 15.010 187.625 113.450 187.795 ;
        RECT 15.095 186.875 16.305 187.625 ;
        RECT 16.475 186.875 17.685 187.625 ;
        RECT 15.095 186.335 15.615 186.875 ;
        RECT 15.785 186.165 16.305 186.705 ;
        RECT 15.095 185.075 16.305 186.165 ;
        RECT 16.475 186.165 16.995 186.705 ;
        RECT 17.165 186.335 17.685 186.875 ;
        RECT 17.855 186.855 21.365 187.625 ;
        RECT 17.855 186.165 19.545 186.685 ;
        RECT 19.715 186.335 21.365 186.855 ;
        RECT 21.575 186.805 21.805 187.625 ;
        RECT 21.975 186.825 22.305 187.455 ;
        RECT 21.555 186.385 21.885 186.635 ;
        RECT 22.055 186.225 22.305 186.825 ;
        RECT 22.475 186.805 22.685 187.625 ;
        RECT 22.915 186.900 23.205 187.625 ;
        RECT 23.465 187.075 23.635 187.455 ;
        RECT 23.815 187.245 24.145 187.625 ;
        RECT 23.465 186.905 24.130 187.075 ;
        RECT 24.325 186.950 24.585 187.455 ;
        RECT 23.395 186.355 23.725 186.725 ;
        RECT 23.960 186.650 24.130 186.905 ;
        RECT 23.960 186.320 24.245 186.650 ;
        RECT 16.475 185.075 17.685 186.165 ;
        RECT 17.855 185.075 21.365 186.165 ;
        RECT 21.575 185.075 21.805 186.215 ;
        RECT 21.975 185.245 22.305 186.225 ;
        RECT 22.475 185.075 22.685 186.215 ;
        RECT 22.915 185.075 23.205 186.240 ;
        RECT 23.960 186.175 24.130 186.320 ;
        RECT 23.465 186.005 24.130 186.175 ;
        RECT 24.415 186.150 24.585 186.950 ;
        RECT 24.870 186.995 25.155 187.455 ;
        RECT 25.325 187.165 25.595 187.625 ;
        RECT 24.870 186.825 25.825 186.995 ;
        RECT 23.465 185.245 23.635 186.005 ;
        RECT 23.815 185.075 24.145 185.835 ;
        RECT 24.315 185.245 24.585 186.150 ;
        RECT 24.755 186.095 25.445 186.655 ;
        RECT 25.615 185.925 25.825 186.825 ;
        RECT 24.870 185.705 25.825 185.925 ;
        RECT 25.995 186.655 26.395 187.455 ;
        RECT 26.585 186.995 26.865 187.455 ;
        RECT 27.385 187.165 27.710 187.625 ;
        RECT 26.585 186.825 27.710 186.995 ;
        RECT 27.880 186.885 28.265 187.455 ;
        RECT 27.260 186.715 27.710 186.825 ;
        RECT 25.995 186.095 27.090 186.655 ;
        RECT 27.260 186.385 27.815 186.715 ;
        RECT 24.870 185.245 25.155 185.705 ;
        RECT 25.325 185.075 25.595 185.535 ;
        RECT 25.995 185.245 26.395 186.095 ;
        RECT 27.260 185.925 27.710 186.385 ;
        RECT 27.985 186.215 28.265 186.885 ;
        RECT 28.710 186.815 28.955 187.420 ;
        RECT 29.175 187.090 29.685 187.625 ;
        RECT 26.585 185.705 27.710 185.925 ;
        RECT 26.585 185.245 26.865 185.705 ;
        RECT 27.385 185.075 27.710 185.535 ;
        RECT 27.880 185.245 28.265 186.215 ;
        RECT 28.435 186.645 29.665 186.815 ;
        RECT 28.435 185.835 28.775 186.645 ;
        RECT 28.945 186.080 29.695 186.270 ;
        RECT 28.435 185.425 28.950 185.835 ;
        RECT 29.185 185.075 29.355 185.835 ;
        RECT 29.525 185.415 29.695 186.080 ;
        RECT 29.865 186.095 30.055 187.455 ;
        RECT 30.225 186.945 30.500 187.455 ;
        RECT 30.690 187.090 31.220 187.455 ;
        RECT 31.645 187.225 31.975 187.625 ;
        RECT 31.045 187.055 31.220 187.090 ;
        RECT 30.225 186.775 30.505 186.945 ;
        RECT 30.225 186.295 30.500 186.775 ;
        RECT 30.705 186.095 30.875 186.895 ;
        RECT 29.865 185.925 30.875 186.095 ;
        RECT 31.045 186.885 31.975 187.055 ;
        RECT 32.145 186.885 32.400 187.455 ;
        RECT 31.045 185.755 31.215 186.885 ;
        RECT 31.805 186.715 31.975 186.885 ;
        RECT 30.090 185.585 31.215 185.755 ;
        RECT 31.385 186.385 31.580 186.715 ;
        RECT 31.805 186.385 32.060 186.715 ;
        RECT 31.385 185.415 31.555 186.385 ;
        RECT 32.230 186.215 32.400 186.885 ;
        RECT 29.525 185.245 31.555 185.415 ;
        RECT 31.725 185.075 31.895 186.215 ;
        RECT 32.065 185.245 32.400 186.215 ;
        RECT 32.950 186.915 33.205 187.445 ;
        RECT 33.385 187.165 33.670 187.625 ;
        RECT 32.950 186.055 33.130 186.915 ;
        RECT 33.850 186.715 34.100 187.365 ;
        RECT 33.300 186.385 34.100 186.715 ;
        RECT 32.950 185.585 33.205 186.055 ;
        RECT 32.865 185.415 33.205 185.585 ;
        RECT 32.950 185.385 33.205 185.415 ;
        RECT 33.385 185.075 33.670 185.875 ;
        RECT 33.850 185.795 34.100 186.385 ;
        RECT 34.300 187.030 34.620 187.360 ;
        RECT 34.800 187.145 35.460 187.625 ;
        RECT 35.660 187.235 36.510 187.405 ;
        RECT 34.300 186.135 34.490 187.030 ;
        RECT 34.810 186.705 35.470 186.975 ;
        RECT 35.140 186.645 35.470 186.705 ;
        RECT 34.660 186.475 34.990 186.535 ;
        RECT 35.660 186.475 35.830 187.235 ;
        RECT 37.070 187.165 37.390 187.625 ;
        RECT 37.590 186.985 37.840 187.415 ;
        RECT 38.130 187.185 38.540 187.625 ;
        RECT 38.710 187.245 39.725 187.445 ;
        RECT 36.000 186.815 37.250 186.985 ;
        RECT 36.000 186.695 36.330 186.815 ;
        RECT 34.660 186.305 36.560 186.475 ;
        RECT 34.300 185.965 36.220 186.135 ;
        RECT 34.300 185.945 34.620 185.965 ;
        RECT 33.850 185.285 34.180 185.795 ;
        RECT 34.450 185.335 34.620 185.945 ;
        RECT 36.390 185.795 36.560 186.305 ;
        RECT 36.730 186.235 36.910 186.645 ;
        RECT 37.080 186.055 37.250 186.815 ;
        RECT 34.790 185.075 35.120 185.765 ;
        RECT 35.350 185.625 36.560 185.795 ;
        RECT 36.730 185.745 37.250 186.055 ;
        RECT 37.420 186.645 37.840 186.985 ;
        RECT 38.130 186.645 38.540 186.975 ;
        RECT 37.420 185.875 37.610 186.645 ;
        RECT 38.710 186.515 38.880 187.245 ;
        RECT 40.025 187.075 40.195 187.405 ;
        RECT 40.365 187.245 40.695 187.625 ;
        RECT 39.050 186.695 39.400 187.065 ;
        RECT 38.710 186.475 39.130 186.515 ;
        RECT 37.780 186.305 39.130 186.475 ;
        RECT 37.780 186.145 38.030 186.305 ;
        RECT 38.540 185.875 38.790 186.135 ;
        RECT 37.420 185.625 38.790 185.875 ;
        RECT 35.350 185.335 35.590 185.625 ;
        RECT 36.390 185.545 36.560 185.625 ;
        RECT 35.790 185.075 36.210 185.455 ;
        RECT 36.390 185.295 37.020 185.545 ;
        RECT 37.490 185.075 37.820 185.455 ;
        RECT 37.990 185.335 38.160 185.625 ;
        RECT 38.960 185.460 39.130 186.305 ;
        RECT 39.580 186.135 39.800 187.005 ;
        RECT 40.025 186.885 40.720 187.075 ;
        RECT 39.300 185.755 39.800 186.135 ;
        RECT 39.970 186.085 40.380 186.705 ;
        RECT 40.550 185.915 40.720 186.885 ;
        RECT 40.025 185.745 40.720 185.915 ;
        RECT 38.340 185.075 38.720 185.455 ;
        RECT 38.960 185.290 39.790 185.460 ;
        RECT 40.025 185.245 40.195 185.745 ;
        RECT 40.365 185.075 40.695 185.575 ;
        RECT 40.910 185.245 41.135 187.365 ;
        RECT 41.305 187.245 41.635 187.625 ;
        RECT 41.805 187.075 41.975 187.365 ;
        RECT 41.310 186.905 41.975 187.075 ;
        RECT 43.245 187.075 43.415 187.455 ;
        RECT 43.595 187.245 43.925 187.625 ;
        RECT 43.245 186.905 43.910 187.075 ;
        RECT 44.105 186.950 44.365 187.455 ;
        RECT 41.310 185.915 41.540 186.905 ;
        RECT 41.710 186.085 42.060 186.735 ;
        RECT 43.175 186.355 43.505 186.725 ;
        RECT 43.740 186.650 43.910 186.905 ;
        RECT 43.740 186.320 44.025 186.650 ;
        RECT 43.740 186.175 43.910 186.320 ;
        RECT 43.245 186.005 43.910 186.175 ;
        RECT 44.195 186.150 44.365 186.950 ;
        RECT 44.810 186.815 45.055 187.420 ;
        RECT 45.275 187.090 45.785 187.625 ;
        RECT 41.310 185.745 41.975 185.915 ;
        RECT 41.305 185.075 41.635 185.575 ;
        RECT 41.805 185.245 41.975 185.745 ;
        RECT 43.245 185.245 43.415 186.005 ;
        RECT 43.595 185.075 43.925 185.835 ;
        RECT 44.095 185.245 44.365 186.150 ;
        RECT 44.535 186.645 45.765 186.815 ;
        RECT 44.535 185.835 44.875 186.645 ;
        RECT 45.045 186.080 45.795 186.270 ;
        RECT 44.535 185.425 45.050 185.835 ;
        RECT 45.285 185.075 45.455 185.835 ;
        RECT 45.625 185.415 45.795 186.080 ;
        RECT 45.965 186.095 46.155 187.455 ;
        RECT 46.325 186.945 46.600 187.455 ;
        RECT 46.790 187.090 47.320 187.455 ;
        RECT 47.745 187.225 48.075 187.625 ;
        RECT 47.145 187.055 47.320 187.090 ;
        RECT 46.325 186.775 46.605 186.945 ;
        RECT 46.325 186.295 46.600 186.775 ;
        RECT 46.805 186.095 46.975 186.895 ;
        RECT 45.965 185.925 46.975 186.095 ;
        RECT 47.145 186.885 48.075 187.055 ;
        RECT 48.245 186.885 48.500 187.455 ;
        RECT 48.675 186.900 48.965 187.625 ;
        RECT 49.600 186.915 49.855 187.445 ;
        RECT 50.025 187.165 50.330 187.625 ;
        RECT 50.575 187.245 51.645 187.415 ;
        RECT 47.145 185.755 47.315 186.885 ;
        RECT 47.905 186.715 48.075 186.885 ;
        RECT 46.190 185.585 47.315 185.755 ;
        RECT 47.485 186.385 47.680 186.715 ;
        RECT 47.905 186.385 48.160 186.715 ;
        RECT 47.485 185.415 47.655 186.385 ;
        RECT 48.330 186.215 48.500 186.885 ;
        RECT 49.600 186.265 49.810 186.915 ;
        RECT 50.575 186.890 50.895 187.245 ;
        RECT 50.570 186.715 50.895 186.890 ;
        RECT 49.980 186.415 50.895 186.715 ;
        RECT 51.065 186.675 51.305 187.075 ;
        RECT 51.475 187.015 51.645 187.245 ;
        RECT 51.815 187.185 52.005 187.625 ;
        RECT 52.175 187.175 53.125 187.455 ;
        RECT 53.345 187.265 53.695 187.435 ;
        RECT 51.475 186.845 52.005 187.015 ;
        RECT 49.980 186.385 50.720 186.415 ;
        RECT 45.625 185.245 47.655 185.415 ;
        RECT 47.825 185.075 47.995 186.215 ;
        RECT 48.165 185.245 48.500 186.215 ;
        RECT 48.675 185.075 48.965 186.240 ;
        RECT 49.600 185.385 49.855 186.265 ;
        RECT 50.025 185.075 50.330 186.215 ;
        RECT 50.550 185.795 50.720 186.385 ;
        RECT 51.065 186.305 51.605 186.675 ;
        RECT 51.785 186.565 52.005 186.845 ;
        RECT 52.175 186.395 52.345 187.175 ;
        RECT 51.940 186.225 52.345 186.395 ;
        RECT 52.515 186.385 52.865 187.005 ;
        RECT 51.940 186.135 52.110 186.225 ;
        RECT 53.035 186.215 53.245 187.005 ;
        RECT 50.890 185.965 52.110 186.135 ;
        RECT 52.570 186.055 53.245 186.215 ;
        RECT 50.550 185.625 51.350 185.795 ;
        RECT 50.670 185.075 51.000 185.455 ;
        RECT 51.180 185.335 51.350 185.625 ;
        RECT 51.940 185.585 52.110 185.965 ;
        RECT 52.280 186.045 53.245 186.055 ;
        RECT 53.435 186.875 53.695 187.265 ;
        RECT 53.905 187.165 54.235 187.625 ;
        RECT 55.110 187.235 55.965 187.405 ;
        RECT 56.170 187.235 56.665 187.405 ;
        RECT 56.835 187.265 57.165 187.625 ;
        RECT 53.435 186.185 53.605 186.875 ;
        RECT 53.775 186.525 53.945 186.705 ;
        RECT 54.115 186.695 54.905 186.945 ;
        RECT 55.110 186.525 55.280 187.235 ;
        RECT 55.450 186.725 55.805 186.945 ;
        RECT 53.775 186.355 55.465 186.525 ;
        RECT 52.280 185.755 52.740 186.045 ;
        RECT 53.435 186.015 54.935 186.185 ;
        RECT 53.435 185.875 53.605 186.015 ;
        RECT 53.045 185.705 53.605 185.875 ;
        RECT 51.520 185.075 51.770 185.535 ;
        RECT 51.940 185.245 52.810 185.585 ;
        RECT 53.045 185.245 53.215 185.705 ;
        RECT 54.050 185.675 55.125 185.845 ;
        RECT 53.385 185.075 53.755 185.535 ;
        RECT 54.050 185.335 54.220 185.675 ;
        RECT 54.390 185.075 54.720 185.505 ;
        RECT 54.955 185.335 55.125 185.675 ;
        RECT 55.295 185.575 55.465 186.355 ;
        RECT 55.635 186.135 55.805 186.725 ;
        RECT 55.975 186.325 56.325 186.945 ;
        RECT 55.635 185.745 56.100 186.135 ;
        RECT 56.495 185.875 56.665 187.235 ;
        RECT 56.835 186.045 57.295 187.095 ;
        RECT 56.270 185.705 56.665 185.875 ;
        RECT 56.270 185.575 56.440 185.705 ;
        RECT 55.295 185.245 55.975 185.575 ;
        RECT 56.190 185.245 56.440 185.575 ;
        RECT 56.610 185.075 56.860 185.535 ;
        RECT 57.030 185.260 57.355 186.045 ;
        RECT 57.525 185.245 57.695 187.365 ;
        RECT 57.865 187.245 58.195 187.625 ;
        RECT 58.365 187.075 58.620 187.365 ;
        RECT 57.870 186.905 58.620 187.075 ;
        RECT 57.870 185.915 58.100 186.905 ;
        RECT 59.255 186.855 62.765 187.625 ;
        RECT 63.205 187.230 63.535 187.625 ;
        RECT 63.705 187.055 63.905 187.410 ;
        RECT 64.075 187.225 64.405 187.625 ;
        RECT 64.575 187.055 64.775 187.400 ;
        RECT 58.270 186.085 58.620 186.735 ;
        RECT 59.255 186.165 60.945 186.685 ;
        RECT 61.115 186.335 62.765 186.855 ;
        RECT 62.935 186.885 64.775 187.055 ;
        RECT 64.945 186.885 65.275 187.625 ;
        RECT 65.510 187.055 65.680 187.305 ;
        RECT 65.510 186.885 65.985 187.055 ;
        RECT 57.870 185.745 58.620 185.915 ;
        RECT 57.865 185.075 58.195 185.575 ;
        RECT 58.365 185.245 58.620 185.745 ;
        RECT 59.255 185.075 62.765 186.165 ;
        RECT 62.935 185.260 63.195 186.885 ;
        RECT 63.375 185.915 63.595 186.715 ;
        RECT 63.835 186.095 64.135 186.715 ;
        RECT 64.305 186.095 64.635 186.715 ;
        RECT 64.805 186.095 65.125 186.715 ;
        RECT 65.295 186.095 65.645 186.715 ;
        RECT 65.815 185.915 65.985 186.885 ;
        RECT 66.155 186.855 68.745 187.625 ;
        RECT 68.920 187.080 74.265 187.625 ;
        RECT 63.375 185.705 65.985 185.915 ;
        RECT 66.155 186.165 67.365 186.685 ;
        RECT 67.535 186.335 68.745 186.855 ;
        RECT 64.945 185.075 65.275 185.525 ;
        RECT 66.155 185.075 68.745 186.165 ;
        RECT 70.510 185.510 70.860 186.760 ;
        RECT 72.340 186.250 72.680 187.080 ;
        RECT 74.435 186.900 74.725 187.625 ;
        RECT 74.895 186.875 76.105 187.625 ;
        RECT 68.920 185.075 74.265 185.510 ;
        RECT 74.435 185.075 74.725 186.240 ;
        RECT 74.895 186.165 75.415 186.705 ;
        RECT 75.585 186.335 76.105 186.875 ;
        RECT 76.315 186.805 76.545 187.625 ;
        RECT 76.715 186.825 77.045 187.455 ;
        RECT 76.295 186.385 76.625 186.635 ;
        RECT 76.795 186.225 77.045 186.825 ;
        RECT 77.215 186.805 77.425 187.625 ;
        RECT 77.930 186.815 78.175 187.420 ;
        RECT 78.395 187.090 78.905 187.625 ;
        RECT 74.895 185.075 76.105 186.165 ;
        RECT 76.315 185.075 76.545 186.215 ;
        RECT 76.715 185.245 77.045 186.225 ;
        RECT 77.655 186.645 78.885 186.815 ;
        RECT 77.215 185.075 77.425 186.215 ;
        RECT 77.655 185.835 77.995 186.645 ;
        RECT 78.165 186.080 78.915 186.270 ;
        RECT 77.655 185.425 78.170 185.835 ;
        RECT 78.405 185.075 78.575 185.835 ;
        RECT 78.745 185.415 78.915 186.080 ;
        RECT 79.085 186.095 79.275 187.455 ;
        RECT 79.445 186.945 79.720 187.455 ;
        RECT 79.910 187.090 80.440 187.455 ;
        RECT 80.865 187.225 81.195 187.625 ;
        RECT 80.265 187.055 80.440 187.090 ;
        RECT 79.445 186.775 79.725 186.945 ;
        RECT 79.445 186.295 79.720 186.775 ;
        RECT 79.925 186.095 80.095 186.895 ;
        RECT 79.085 185.925 80.095 186.095 ;
        RECT 80.265 186.885 81.195 187.055 ;
        RECT 81.365 186.885 81.620 187.455 ;
        RECT 80.265 185.755 80.435 186.885 ;
        RECT 81.025 186.715 81.195 186.885 ;
        RECT 79.310 185.585 80.435 185.755 ;
        RECT 80.605 186.385 80.800 186.715 ;
        RECT 81.025 186.385 81.280 186.715 ;
        RECT 80.605 185.415 80.775 186.385 ;
        RECT 81.450 186.215 81.620 186.885 ;
        RECT 78.745 185.245 80.775 185.415 ;
        RECT 80.945 185.075 81.115 186.215 ;
        RECT 81.285 185.245 81.620 186.215 ;
        RECT 81.795 186.950 82.055 187.455 ;
        RECT 82.235 187.245 82.565 187.625 ;
        RECT 82.745 187.075 82.915 187.455 ;
        RECT 81.795 186.150 81.965 186.950 ;
        RECT 82.250 186.905 82.915 187.075 ;
        RECT 82.250 186.650 82.420 186.905 ;
        RECT 83.635 186.885 84.020 187.455 ;
        RECT 84.190 187.165 84.515 187.625 ;
        RECT 85.035 186.995 85.315 187.455 ;
        RECT 82.135 186.320 82.420 186.650 ;
        RECT 82.655 186.355 82.985 186.725 ;
        RECT 82.250 186.175 82.420 186.320 ;
        RECT 83.635 186.215 83.915 186.885 ;
        RECT 84.190 186.825 85.315 186.995 ;
        RECT 84.190 186.715 84.640 186.825 ;
        RECT 84.085 186.385 84.640 186.715 ;
        RECT 85.505 186.655 85.905 187.455 ;
        RECT 86.305 187.165 86.575 187.625 ;
        RECT 86.745 186.995 87.030 187.455 ;
        RECT 81.795 185.245 82.065 186.150 ;
        RECT 82.250 186.005 82.915 186.175 ;
        RECT 82.235 185.075 82.565 185.835 ;
        RECT 82.745 185.245 82.915 186.005 ;
        RECT 83.635 185.245 84.020 186.215 ;
        RECT 84.190 185.925 84.640 186.385 ;
        RECT 84.810 186.095 85.905 186.655 ;
        RECT 84.190 185.705 85.315 185.925 ;
        RECT 84.190 185.075 84.515 185.535 ;
        RECT 85.035 185.245 85.315 185.705 ;
        RECT 85.505 185.245 85.905 186.095 ;
        RECT 86.075 186.825 87.030 186.995 ;
        RECT 86.075 185.925 86.285 186.825 ;
        RECT 87.375 186.805 87.585 187.625 ;
        RECT 87.755 186.825 88.085 187.455 ;
        RECT 86.455 186.095 87.145 186.655 ;
        RECT 87.755 186.225 88.005 186.825 ;
        RECT 88.255 186.805 88.485 187.625 ;
        RECT 89.730 186.995 90.015 187.455 ;
        RECT 90.185 187.165 90.455 187.625 ;
        RECT 89.730 186.825 90.685 186.995 ;
        RECT 88.175 186.385 88.505 186.635 ;
        RECT 86.075 185.705 87.030 185.925 ;
        RECT 86.305 185.075 86.575 185.535 ;
        RECT 86.745 185.245 87.030 185.705 ;
        RECT 87.375 185.075 87.585 186.215 ;
        RECT 87.755 185.245 88.085 186.225 ;
        RECT 88.255 185.075 88.485 186.215 ;
        RECT 89.615 186.095 90.305 186.655 ;
        RECT 90.475 185.925 90.685 186.825 ;
        RECT 89.730 185.705 90.685 185.925 ;
        RECT 90.855 186.655 91.255 187.455 ;
        RECT 91.445 186.995 91.725 187.455 ;
        RECT 92.245 187.165 92.570 187.625 ;
        RECT 91.445 186.825 92.570 186.995 ;
        RECT 92.740 186.885 93.125 187.455 ;
        RECT 92.120 186.715 92.570 186.825 ;
        RECT 90.855 186.095 91.950 186.655 ;
        RECT 92.120 186.385 92.675 186.715 ;
        RECT 89.730 185.245 90.015 185.705 ;
        RECT 90.185 185.075 90.455 185.535 ;
        RECT 90.855 185.245 91.255 186.095 ;
        RECT 92.120 185.925 92.570 186.385 ;
        RECT 92.845 186.215 93.125 186.885 ;
        RECT 91.445 185.705 92.570 185.925 ;
        RECT 91.445 185.245 91.725 185.705 ;
        RECT 92.245 185.075 92.570 185.535 ;
        RECT 92.740 185.245 93.125 186.215 ;
        RECT 93.300 186.885 93.555 187.455 ;
        RECT 93.725 187.225 94.055 187.625 ;
        RECT 94.480 187.090 95.010 187.455 ;
        RECT 94.480 187.055 94.655 187.090 ;
        RECT 93.725 186.885 94.655 187.055 ;
        RECT 93.300 186.215 93.470 186.885 ;
        RECT 93.725 186.715 93.895 186.885 ;
        RECT 93.640 186.385 93.895 186.715 ;
        RECT 94.120 186.385 94.315 186.715 ;
        RECT 93.300 185.245 93.635 186.215 ;
        RECT 93.805 185.075 93.975 186.215 ;
        RECT 94.145 185.415 94.315 186.385 ;
        RECT 94.485 185.755 94.655 186.885 ;
        RECT 94.825 186.095 94.995 186.895 ;
        RECT 95.200 186.605 95.475 187.455 ;
        RECT 95.195 186.435 95.475 186.605 ;
        RECT 95.200 186.295 95.475 186.435 ;
        RECT 95.645 186.095 95.835 187.455 ;
        RECT 96.015 187.090 96.525 187.625 ;
        RECT 96.745 186.815 96.990 187.420 ;
        RECT 97.435 186.855 100.025 187.625 ;
        RECT 100.195 186.900 100.485 187.625 ;
        RECT 96.035 186.645 97.265 186.815 ;
        RECT 94.825 185.925 95.835 186.095 ;
        RECT 96.005 186.080 96.755 186.270 ;
        RECT 94.485 185.585 95.610 185.755 ;
        RECT 96.005 185.415 96.175 186.080 ;
        RECT 96.925 185.835 97.265 186.645 ;
        RECT 94.145 185.245 96.175 185.415 ;
        RECT 96.345 185.075 96.515 185.835 ;
        RECT 96.750 185.425 97.265 185.835 ;
        RECT 97.435 186.165 98.645 186.685 ;
        RECT 98.815 186.335 100.025 186.855 ;
        RECT 100.695 186.805 100.925 187.625 ;
        RECT 101.095 186.825 101.425 187.455 ;
        RECT 100.675 186.385 101.005 186.635 ;
        RECT 97.435 185.075 100.025 186.165 ;
        RECT 100.195 185.075 100.485 186.240 ;
        RECT 101.175 186.225 101.425 186.825 ;
        RECT 101.595 186.805 101.805 187.625 ;
        RECT 102.040 186.915 102.295 187.445 ;
        RECT 102.465 187.165 102.770 187.625 ;
        RECT 103.015 187.245 104.085 187.415 ;
        RECT 100.695 185.075 100.925 186.215 ;
        RECT 101.095 185.245 101.425 186.225 ;
        RECT 102.040 186.265 102.250 186.915 ;
        RECT 103.015 186.890 103.335 187.245 ;
        RECT 103.010 186.715 103.335 186.890 ;
        RECT 102.420 186.415 103.335 186.715 ;
        RECT 103.505 186.675 103.745 187.075 ;
        RECT 103.915 187.015 104.085 187.245 ;
        RECT 104.255 187.185 104.445 187.625 ;
        RECT 104.615 187.175 105.565 187.455 ;
        RECT 105.785 187.265 106.135 187.435 ;
        RECT 103.915 186.845 104.445 187.015 ;
        RECT 102.420 186.385 103.160 186.415 ;
        RECT 101.595 185.075 101.805 186.215 ;
        RECT 102.040 185.385 102.295 186.265 ;
        RECT 102.465 185.075 102.770 186.215 ;
        RECT 102.990 185.795 103.160 186.385 ;
        RECT 103.505 186.305 104.045 186.675 ;
        RECT 104.225 186.565 104.445 186.845 ;
        RECT 104.615 186.395 104.785 187.175 ;
        RECT 104.380 186.225 104.785 186.395 ;
        RECT 104.955 186.385 105.305 187.005 ;
        RECT 104.380 186.135 104.550 186.225 ;
        RECT 105.475 186.215 105.685 187.005 ;
        RECT 103.330 185.965 104.550 186.135 ;
        RECT 105.010 186.055 105.685 186.215 ;
        RECT 102.990 185.625 103.790 185.795 ;
        RECT 103.110 185.075 103.440 185.455 ;
        RECT 103.620 185.335 103.790 185.625 ;
        RECT 104.380 185.585 104.550 185.965 ;
        RECT 104.720 186.045 105.685 186.055 ;
        RECT 105.875 186.875 106.135 187.265 ;
        RECT 106.345 187.165 106.675 187.625 ;
        RECT 107.550 187.235 108.405 187.405 ;
        RECT 108.610 187.235 109.105 187.405 ;
        RECT 109.275 187.265 109.605 187.625 ;
        RECT 105.875 186.185 106.045 186.875 ;
        RECT 106.215 186.525 106.385 186.705 ;
        RECT 106.555 186.695 107.345 186.945 ;
        RECT 107.550 186.525 107.720 187.235 ;
        RECT 107.890 186.725 108.245 186.945 ;
        RECT 106.215 186.355 107.905 186.525 ;
        RECT 104.720 185.755 105.180 186.045 ;
        RECT 105.875 186.015 107.375 186.185 ;
        RECT 105.875 185.875 106.045 186.015 ;
        RECT 105.485 185.705 106.045 185.875 ;
        RECT 103.960 185.075 104.210 185.535 ;
        RECT 104.380 185.245 105.250 185.585 ;
        RECT 105.485 185.245 105.655 185.705 ;
        RECT 106.490 185.675 107.565 185.845 ;
        RECT 105.825 185.075 106.195 185.535 ;
        RECT 106.490 185.335 106.660 185.675 ;
        RECT 106.830 185.075 107.160 185.505 ;
        RECT 107.395 185.335 107.565 185.675 ;
        RECT 107.735 185.575 107.905 186.355 ;
        RECT 108.075 186.135 108.245 186.725 ;
        RECT 108.415 186.325 108.765 186.945 ;
        RECT 108.075 185.745 108.540 186.135 ;
        RECT 108.935 185.875 109.105 187.235 ;
        RECT 109.275 186.045 109.735 187.095 ;
        RECT 108.710 185.705 109.105 185.875 ;
        RECT 108.710 185.575 108.880 185.705 ;
        RECT 107.735 185.245 108.415 185.575 ;
        RECT 108.630 185.245 108.880 185.575 ;
        RECT 109.050 185.075 109.300 185.535 ;
        RECT 109.470 185.260 109.795 186.045 ;
        RECT 109.965 185.245 110.135 187.365 ;
        RECT 110.305 187.245 110.635 187.625 ;
        RECT 110.805 187.075 111.060 187.365 ;
        RECT 110.310 186.905 111.060 187.075 ;
        RECT 110.310 185.915 110.540 186.905 ;
        RECT 112.155 186.875 113.365 187.625 ;
        RECT 110.710 186.085 111.060 186.735 ;
        RECT 112.155 186.165 112.675 186.705 ;
        RECT 112.845 186.335 113.365 186.875 ;
        RECT 110.310 185.745 111.060 185.915 ;
        RECT 110.305 185.075 110.635 185.575 ;
        RECT 110.805 185.245 111.060 185.745 ;
        RECT 112.155 185.075 113.365 186.165 ;
        RECT 15.010 184.905 113.450 185.075 ;
        RECT 15.095 183.815 16.305 184.905 ;
        RECT 15.095 183.105 15.615 183.645 ;
        RECT 15.785 183.275 16.305 183.815 ;
        RECT 16.935 183.815 20.445 184.905 ;
        RECT 16.935 183.295 18.625 183.815 ;
        RECT 20.615 183.765 21.000 184.735 ;
        RECT 21.170 184.445 21.495 184.905 ;
        RECT 22.015 184.275 22.295 184.735 ;
        RECT 21.170 184.055 22.295 184.275 ;
        RECT 18.795 183.125 20.445 183.645 ;
        RECT 15.095 182.355 16.305 183.105 ;
        RECT 16.935 182.355 20.445 183.125 ;
        RECT 20.615 183.095 20.895 183.765 ;
        RECT 21.170 183.595 21.620 184.055 ;
        RECT 22.485 183.885 22.885 184.735 ;
        RECT 23.285 184.445 23.555 184.905 ;
        RECT 23.725 184.275 24.010 184.735 ;
        RECT 21.065 183.265 21.620 183.595 ;
        RECT 21.790 183.325 22.885 183.885 ;
        RECT 21.170 183.155 21.620 183.265 ;
        RECT 20.615 182.525 21.000 183.095 ;
        RECT 21.170 182.985 22.295 183.155 ;
        RECT 21.170 182.355 21.495 182.815 ;
        RECT 22.015 182.525 22.295 182.985 ;
        RECT 22.485 182.525 22.885 183.325 ;
        RECT 23.055 184.055 24.010 184.275 ;
        RECT 24.300 184.235 24.555 184.735 ;
        RECT 24.725 184.405 25.055 184.905 ;
        RECT 24.300 184.065 25.050 184.235 ;
        RECT 23.055 183.155 23.265 184.055 ;
        RECT 23.435 183.325 24.125 183.885 ;
        RECT 24.300 183.245 24.650 183.895 ;
        RECT 23.055 182.985 24.010 183.155 ;
        RECT 24.820 183.075 25.050 184.065 ;
        RECT 23.285 182.355 23.555 182.815 ;
        RECT 23.725 182.525 24.010 182.985 ;
        RECT 24.300 182.905 25.050 183.075 ;
        RECT 24.300 182.615 24.555 182.905 ;
        RECT 24.725 182.355 25.055 182.735 ;
        RECT 25.225 182.615 25.395 184.735 ;
        RECT 25.565 183.935 25.890 184.720 ;
        RECT 26.060 184.445 26.310 184.905 ;
        RECT 26.480 184.405 26.730 184.735 ;
        RECT 26.945 184.405 27.625 184.735 ;
        RECT 26.480 184.275 26.650 184.405 ;
        RECT 26.255 184.105 26.650 184.275 ;
        RECT 25.625 182.885 26.085 183.935 ;
        RECT 26.255 182.745 26.425 184.105 ;
        RECT 26.820 183.845 27.285 184.235 ;
        RECT 26.595 183.035 26.945 183.655 ;
        RECT 27.115 183.255 27.285 183.845 ;
        RECT 27.455 183.625 27.625 184.405 ;
        RECT 27.795 184.305 27.965 184.645 ;
        RECT 28.200 184.475 28.530 184.905 ;
        RECT 28.700 184.305 28.870 184.645 ;
        RECT 29.165 184.445 29.535 184.905 ;
        RECT 27.795 184.135 28.870 184.305 ;
        RECT 29.705 184.275 29.875 184.735 ;
        RECT 30.110 184.395 30.980 184.735 ;
        RECT 31.150 184.445 31.400 184.905 ;
        RECT 29.315 184.105 29.875 184.275 ;
        RECT 29.315 183.965 29.485 184.105 ;
        RECT 27.985 183.795 29.485 183.965 ;
        RECT 30.180 183.935 30.640 184.225 ;
        RECT 27.455 183.455 29.145 183.625 ;
        RECT 27.115 183.035 27.470 183.255 ;
        RECT 27.640 182.745 27.810 183.455 ;
        RECT 28.015 183.035 28.805 183.285 ;
        RECT 28.975 183.275 29.145 183.455 ;
        RECT 29.315 183.105 29.485 183.795 ;
        RECT 25.755 182.355 26.085 182.715 ;
        RECT 26.255 182.575 26.750 182.745 ;
        RECT 26.955 182.575 27.810 182.745 ;
        RECT 28.685 182.355 29.015 182.815 ;
        RECT 29.225 182.715 29.485 183.105 ;
        RECT 29.675 183.925 30.640 183.935 ;
        RECT 30.810 184.015 30.980 184.395 ;
        RECT 31.570 184.355 31.740 184.645 ;
        RECT 31.920 184.525 32.250 184.905 ;
        RECT 31.570 184.185 32.370 184.355 ;
        RECT 29.675 183.765 30.350 183.925 ;
        RECT 30.810 183.845 32.030 184.015 ;
        RECT 29.675 182.975 29.885 183.765 ;
        RECT 30.810 183.755 30.980 183.845 ;
        RECT 30.055 182.975 30.405 183.595 ;
        RECT 30.575 183.585 30.980 183.755 ;
        RECT 30.575 182.805 30.745 183.585 ;
        RECT 30.915 183.135 31.135 183.415 ;
        RECT 31.315 183.305 31.855 183.675 ;
        RECT 32.200 183.595 32.370 184.185 ;
        RECT 32.590 183.765 32.895 184.905 ;
        RECT 33.065 183.715 33.320 184.595 ;
        RECT 34.455 183.765 34.685 184.905 ;
        RECT 34.855 183.755 35.185 184.735 ;
        RECT 35.355 183.765 35.565 184.905 ;
        RECT 32.200 183.565 32.940 183.595 ;
        RECT 30.915 182.965 31.445 183.135 ;
        RECT 29.225 182.545 29.575 182.715 ;
        RECT 29.795 182.525 30.745 182.805 ;
        RECT 30.915 182.355 31.105 182.795 ;
        RECT 31.275 182.735 31.445 182.965 ;
        RECT 31.615 182.905 31.855 183.305 ;
        RECT 32.025 183.265 32.940 183.565 ;
        RECT 32.025 183.090 32.350 183.265 ;
        RECT 32.025 182.735 32.345 183.090 ;
        RECT 33.110 183.065 33.320 183.715 ;
        RECT 34.435 183.345 34.765 183.595 ;
        RECT 31.275 182.565 32.345 182.735 ;
        RECT 32.590 182.355 32.895 182.815 ;
        RECT 33.065 182.535 33.320 183.065 ;
        RECT 34.455 182.355 34.685 183.175 ;
        RECT 34.935 183.155 35.185 183.755 ;
        RECT 35.795 183.740 36.085 184.905 ;
        RECT 36.255 183.815 37.925 184.905 ;
        RECT 38.185 183.975 38.355 184.735 ;
        RECT 38.535 184.145 38.865 184.905 ;
        RECT 36.255 183.295 37.005 183.815 ;
        RECT 38.185 183.805 38.850 183.975 ;
        RECT 39.035 183.830 39.305 184.735 ;
        RECT 38.680 183.660 38.850 183.805 ;
        RECT 34.855 182.525 35.185 183.155 ;
        RECT 35.355 182.355 35.565 183.175 ;
        RECT 37.175 183.125 37.925 183.645 ;
        RECT 38.115 183.255 38.445 183.625 ;
        RECT 38.680 183.330 38.965 183.660 ;
        RECT 35.795 182.355 36.085 183.080 ;
        RECT 36.255 182.355 37.925 183.125 ;
        RECT 38.680 183.075 38.850 183.330 ;
        RECT 38.185 182.905 38.850 183.075 ;
        RECT 39.135 183.030 39.305 183.830 ;
        RECT 38.185 182.525 38.355 182.905 ;
        RECT 38.535 182.355 38.865 182.735 ;
        RECT 39.045 182.525 39.305 183.030 ;
        RECT 39.480 183.765 39.815 184.735 ;
        RECT 39.985 183.765 40.155 184.905 ;
        RECT 40.325 184.565 42.355 184.735 ;
        RECT 39.480 183.095 39.650 183.765 ;
        RECT 40.325 183.595 40.495 184.565 ;
        RECT 39.820 183.265 40.075 183.595 ;
        RECT 40.300 183.265 40.495 183.595 ;
        RECT 40.665 184.225 41.790 184.395 ;
        RECT 39.905 183.095 40.075 183.265 ;
        RECT 40.665 183.095 40.835 184.225 ;
        RECT 39.480 182.525 39.735 183.095 ;
        RECT 39.905 182.925 40.835 183.095 ;
        RECT 41.005 183.885 42.015 184.055 ;
        RECT 41.005 183.085 41.175 183.885 ;
        RECT 40.660 182.890 40.835 182.925 ;
        RECT 39.905 182.355 40.235 182.755 ;
        RECT 40.660 182.525 41.190 182.890 ;
        RECT 41.380 182.865 41.655 183.685 ;
        RECT 41.375 182.695 41.655 182.865 ;
        RECT 41.380 182.525 41.655 182.695 ;
        RECT 41.825 182.525 42.015 183.885 ;
        RECT 42.185 183.900 42.355 184.565 ;
        RECT 42.525 184.145 42.695 184.905 ;
        RECT 42.930 184.145 43.445 184.555 ;
        RECT 42.185 183.710 42.935 183.900 ;
        RECT 43.105 183.335 43.445 184.145 ;
        RECT 42.215 183.165 43.445 183.335 ;
        RECT 43.620 183.715 43.875 184.595 ;
        RECT 44.045 183.765 44.350 184.905 ;
        RECT 44.690 184.525 45.020 184.905 ;
        RECT 45.200 184.355 45.370 184.645 ;
        RECT 45.540 184.445 45.790 184.905 ;
        RECT 44.570 184.185 45.370 184.355 ;
        RECT 45.960 184.395 46.830 184.735 ;
        RECT 42.195 182.355 42.705 182.890 ;
        RECT 42.925 182.560 43.170 183.165 ;
        RECT 43.620 183.065 43.830 183.715 ;
        RECT 44.570 183.595 44.740 184.185 ;
        RECT 45.960 184.015 46.130 184.395 ;
        RECT 47.065 184.275 47.235 184.735 ;
        RECT 47.405 184.445 47.775 184.905 ;
        RECT 48.070 184.305 48.240 184.645 ;
        RECT 48.410 184.475 48.740 184.905 ;
        RECT 48.975 184.305 49.145 184.645 ;
        RECT 44.910 183.845 46.130 184.015 ;
        RECT 46.300 183.935 46.760 184.225 ;
        RECT 47.065 184.105 47.625 184.275 ;
        RECT 48.070 184.135 49.145 184.305 ;
        RECT 49.315 184.405 49.995 184.735 ;
        RECT 50.210 184.405 50.460 184.735 ;
        RECT 50.630 184.445 50.880 184.905 ;
        RECT 47.455 183.965 47.625 184.105 ;
        RECT 46.300 183.925 47.265 183.935 ;
        RECT 45.960 183.755 46.130 183.845 ;
        RECT 46.590 183.765 47.265 183.925 ;
        RECT 44.000 183.565 44.740 183.595 ;
        RECT 44.000 183.265 44.915 183.565 ;
        RECT 44.590 183.090 44.915 183.265 ;
        RECT 43.620 182.535 43.875 183.065 ;
        RECT 44.045 182.355 44.350 182.815 ;
        RECT 44.595 182.735 44.915 183.090 ;
        RECT 45.085 183.305 45.625 183.675 ;
        RECT 45.960 183.585 46.365 183.755 ;
        RECT 45.085 182.905 45.325 183.305 ;
        RECT 45.805 183.135 46.025 183.415 ;
        RECT 45.495 182.965 46.025 183.135 ;
        RECT 45.495 182.735 45.665 182.965 ;
        RECT 46.195 182.805 46.365 183.585 ;
        RECT 46.535 182.975 46.885 183.595 ;
        RECT 47.055 182.975 47.265 183.765 ;
        RECT 47.455 183.795 48.955 183.965 ;
        RECT 47.455 183.105 47.625 183.795 ;
        RECT 49.315 183.625 49.485 184.405 ;
        RECT 50.290 184.275 50.460 184.405 ;
        RECT 47.795 183.455 49.485 183.625 ;
        RECT 49.655 183.845 50.120 184.235 ;
        RECT 50.290 184.105 50.685 184.275 ;
        RECT 47.795 183.275 47.965 183.455 ;
        RECT 44.595 182.565 45.665 182.735 ;
        RECT 45.835 182.355 46.025 182.795 ;
        RECT 46.195 182.525 47.145 182.805 ;
        RECT 47.455 182.715 47.715 183.105 ;
        RECT 48.135 183.035 48.925 183.285 ;
        RECT 47.365 182.545 47.715 182.715 ;
        RECT 47.925 182.355 48.255 182.815 ;
        RECT 49.130 182.745 49.300 183.455 ;
        RECT 49.655 183.255 49.825 183.845 ;
        RECT 49.470 183.035 49.825 183.255 ;
        RECT 49.995 183.035 50.345 183.655 ;
        RECT 50.515 182.745 50.685 184.105 ;
        RECT 51.050 183.935 51.375 184.720 ;
        RECT 50.855 182.885 51.315 183.935 ;
        RECT 49.130 182.575 49.985 182.745 ;
        RECT 50.190 182.575 50.685 182.745 ;
        RECT 50.855 182.355 51.185 182.715 ;
        RECT 51.545 182.615 51.715 184.735 ;
        RECT 51.885 184.405 52.215 184.905 ;
        RECT 52.385 184.235 52.640 184.735 ;
        RECT 51.890 184.065 52.640 184.235 ;
        RECT 52.930 184.275 53.215 184.735 ;
        RECT 53.385 184.445 53.655 184.905 ;
        RECT 51.890 183.075 52.120 184.065 ;
        RECT 52.930 184.055 53.885 184.275 ;
        RECT 52.290 183.245 52.640 183.895 ;
        RECT 52.815 183.325 53.505 183.885 ;
        RECT 53.675 183.155 53.885 184.055 ;
        RECT 51.890 182.905 52.640 183.075 ;
        RECT 51.885 182.355 52.215 182.735 ;
        RECT 52.385 182.615 52.640 182.905 ;
        RECT 52.930 182.985 53.885 183.155 ;
        RECT 54.055 183.885 54.455 184.735 ;
        RECT 54.645 184.275 54.925 184.735 ;
        RECT 55.445 184.445 55.770 184.905 ;
        RECT 54.645 184.055 55.770 184.275 ;
        RECT 54.055 183.325 55.150 183.885 ;
        RECT 55.320 183.595 55.770 184.055 ;
        RECT 55.940 183.765 56.325 184.735 ;
        RECT 56.555 183.765 56.765 184.905 ;
        RECT 52.930 182.525 53.215 182.985 ;
        RECT 53.385 182.355 53.655 182.815 ;
        RECT 54.055 182.525 54.455 183.325 ;
        RECT 55.320 183.265 55.875 183.595 ;
        RECT 55.320 183.155 55.770 183.265 ;
        RECT 54.645 182.985 55.770 183.155 ;
        RECT 56.045 183.095 56.325 183.765 ;
        RECT 56.935 183.755 57.265 184.735 ;
        RECT 57.435 183.765 57.665 184.905 ;
        RECT 59.045 184.455 59.375 184.905 ;
        RECT 58.335 184.065 60.945 184.275 ;
        RECT 54.645 182.525 54.925 182.985 ;
        RECT 55.445 182.355 55.770 182.815 ;
        RECT 55.940 182.525 56.325 183.095 ;
        RECT 56.555 182.355 56.765 183.175 ;
        RECT 56.935 183.155 57.185 183.755 ;
        RECT 57.355 183.345 57.685 183.595 ;
        RECT 56.935 182.525 57.265 183.155 ;
        RECT 57.435 182.355 57.665 183.175 ;
        RECT 58.335 183.095 58.505 184.065 ;
        RECT 58.675 183.265 59.025 183.885 ;
        RECT 59.195 183.265 59.515 183.885 ;
        RECT 59.685 183.265 60.015 183.885 ;
        RECT 60.185 183.265 60.485 183.885 ;
        RECT 60.725 183.265 60.945 184.065 ;
        RECT 61.125 183.095 61.385 184.720 ;
        RECT 61.555 183.740 61.845 184.905 ;
        RECT 62.015 183.815 64.605 184.905 ;
        RECT 64.775 184.405 65.035 184.735 ;
        RECT 65.345 184.525 65.675 184.905 ;
        RECT 62.015 183.295 63.225 183.815 ;
        RECT 64.775 183.725 64.945 184.405 ;
        RECT 65.915 184.355 66.105 184.735 ;
        RECT 66.355 184.525 66.685 184.905 ;
        RECT 66.895 184.355 67.065 184.735 ;
        RECT 67.260 184.525 67.590 184.905 ;
        RECT 67.850 184.355 68.020 184.735 ;
        RECT 68.445 184.525 68.775 184.905 ;
        RECT 65.115 183.895 65.465 184.225 ;
        RECT 65.915 184.185 66.655 184.355 ;
        RECT 65.735 183.845 66.315 184.015 ;
        RECT 65.735 183.725 65.905 183.845 ;
        RECT 63.395 183.125 64.605 183.645 ;
        RECT 58.335 182.925 58.810 183.095 ;
        RECT 58.640 182.675 58.810 182.925 ;
        RECT 59.045 182.355 59.375 183.095 ;
        RECT 59.545 182.925 61.385 183.095 ;
        RECT 59.545 182.580 59.745 182.925 ;
        RECT 59.915 182.355 60.245 182.755 ;
        RECT 60.415 182.570 60.615 182.925 ;
        RECT 60.785 182.355 61.115 182.750 ;
        RECT 61.555 182.355 61.845 183.080 ;
        RECT 62.015 182.355 64.605 183.125 ;
        RECT 64.775 183.555 65.905 183.725 ;
        RECT 66.485 183.675 66.655 184.185 ;
        RECT 64.775 182.855 64.945 183.555 ;
        RECT 66.085 183.505 66.655 183.675 ;
        RECT 66.825 184.185 68.775 184.355 ;
        RECT 65.295 183.215 65.915 183.385 ;
        RECT 65.295 183.035 65.505 183.215 ;
        RECT 66.085 183.025 66.255 183.505 ;
        RECT 66.825 183.195 66.995 184.185 ;
        RECT 67.585 183.595 67.770 183.905 ;
        RECT 68.040 183.595 68.235 183.905 ;
        RECT 64.775 182.525 65.035 182.855 ;
        RECT 65.345 182.355 65.675 182.735 ;
        RECT 65.855 182.695 66.255 183.025 ;
        RECT 66.445 182.865 66.995 183.195 ;
        RECT 67.165 182.695 67.335 183.595 ;
        RECT 65.855 182.525 67.335 182.695 ;
        RECT 67.585 183.265 67.815 183.595 ;
        RECT 68.040 183.265 68.295 183.595 ;
        RECT 68.605 183.265 68.775 184.185 ;
        RECT 67.585 182.685 67.770 183.265 ;
        RECT 68.040 182.690 68.235 183.265 ;
        RECT 68.445 182.355 68.775 182.735 ;
        RECT 68.945 182.525 69.205 184.735 ;
        RECT 69.375 183.095 69.635 184.720 ;
        RECT 71.385 184.455 71.715 184.905 ;
        RECT 73.890 184.565 74.145 184.595 ;
        RECT 73.805 184.395 74.145 184.565 ;
        RECT 69.815 184.065 72.425 184.275 ;
        RECT 69.815 183.265 70.035 184.065 ;
        RECT 70.275 183.265 70.575 183.885 ;
        RECT 70.745 183.265 71.075 183.885 ;
        RECT 71.245 183.265 71.565 183.885 ;
        RECT 71.735 183.265 72.085 183.885 ;
        RECT 72.255 183.095 72.425 184.065 ;
        RECT 69.375 182.925 71.215 183.095 ;
        RECT 69.645 182.355 69.975 182.750 ;
        RECT 70.145 182.570 70.345 182.925 ;
        RECT 70.515 182.355 70.845 182.755 ;
        RECT 71.015 182.580 71.215 182.925 ;
        RECT 71.385 182.355 71.715 183.095 ;
        RECT 71.950 182.925 72.425 183.095 ;
        RECT 73.890 183.925 74.145 184.395 ;
        RECT 74.325 184.105 74.610 184.905 ;
        RECT 74.790 184.185 75.120 184.695 ;
        RECT 73.890 183.065 74.070 183.925 ;
        RECT 74.790 183.595 75.040 184.185 ;
        RECT 75.390 184.035 75.560 184.645 ;
        RECT 75.730 184.215 76.060 184.905 ;
        RECT 76.290 184.355 76.530 184.645 ;
        RECT 76.730 184.525 77.150 184.905 ;
        RECT 77.330 184.435 77.960 184.685 ;
        RECT 78.430 184.525 78.760 184.905 ;
        RECT 77.330 184.355 77.500 184.435 ;
        RECT 78.930 184.355 79.100 184.645 ;
        RECT 79.280 184.525 79.660 184.905 ;
        RECT 79.900 184.520 80.730 184.690 ;
        RECT 76.290 184.185 77.500 184.355 ;
        RECT 74.240 183.265 75.040 183.595 ;
        RECT 71.950 182.675 72.120 182.925 ;
        RECT 73.890 182.535 74.145 183.065 ;
        RECT 74.325 182.355 74.610 182.815 ;
        RECT 74.790 182.615 75.040 183.265 ;
        RECT 75.240 184.015 75.560 184.035 ;
        RECT 75.240 183.845 77.160 184.015 ;
        RECT 75.240 182.950 75.430 183.845 ;
        RECT 77.330 183.675 77.500 184.185 ;
        RECT 77.670 183.925 78.190 184.235 ;
        RECT 75.600 183.505 77.500 183.675 ;
        RECT 75.600 183.445 75.930 183.505 ;
        RECT 76.080 183.275 76.410 183.335 ;
        RECT 75.750 183.005 76.410 183.275 ;
        RECT 75.240 182.620 75.560 182.950 ;
        RECT 75.740 182.355 76.400 182.835 ;
        RECT 76.600 182.745 76.770 183.505 ;
        RECT 77.670 183.335 77.850 183.745 ;
        RECT 76.940 183.165 77.270 183.285 ;
        RECT 78.020 183.165 78.190 183.925 ;
        RECT 76.940 182.995 78.190 183.165 ;
        RECT 78.360 184.105 79.730 184.355 ;
        RECT 78.360 183.335 78.550 184.105 ;
        RECT 79.480 183.845 79.730 184.105 ;
        RECT 78.720 183.675 78.970 183.835 ;
        RECT 79.900 183.675 80.070 184.520 ;
        RECT 80.965 184.235 81.135 184.735 ;
        RECT 81.305 184.405 81.635 184.905 ;
        RECT 80.240 183.845 80.740 184.225 ;
        RECT 80.965 184.065 81.660 184.235 ;
        RECT 78.720 183.505 80.070 183.675 ;
        RECT 79.650 183.465 80.070 183.505 ;
        RECT 78.360 182.995 78.780 183.335 ;
        RECT 79.070 183.005 79.480 183.335 ;
        RECT 76.600 182.575 77.450 182.745 ;
        RECT 78.010 182.355 78.330 182.815 ;
        RECT 78.530 182.565 78.780 182.995 ;
        RECT 79.070 182.355 79.480 182.795 ;
        RECT 79.650 182.735 79.820 183.465 ;
        RECT 79.990 182.915 80.340 183.285 ;
        RECT 80.520 182.975 80.740 183.845 ;
        RECT 80.910 183.275 81.320 183.895 ;
        RECT 81.490 183.095 81.660 184.065 ;
        RECT 80.965 182.905 81.660 183.095 ;
        RECT 79.650 182.535 80.665 182.735 ;
        RECT 80.965 182.575 81.135 182.905 ;
        RECT 81.305 182.355 81.635 182.735 ;
        RECT 81.850 182.615 82.075 184.735 ;
        RECT 82.245 184.405 82.575 184.905 ;
        RECT 82.745 184.235 82.915 184.735 ;
        RECT 82.250 184.065 82.915 184.235 ;
        RECT 83.175 184.145 83.690 184.555 ;
        RECT 83.925 184.145 84.095 184.905 ;
        RECT 84.265 184.565 86.295 184.735 ;
        RECT 82.250 183.075 82.480 184.065 ;
        RECT 82.650 183.245 83.000 183.895 ;
        RECT 83.175 183.335 83.515 184.145 ;
        RECT 84.265 183.900 84.435 184.565 ;
        RECT 84.830 184.225 85.955 184.395 ;
        RECT 83.685 183.710 84.435 183.900 ;
        RECT 84.605 183.885 85.615 184.055 ;
        RECT 83.175 183.165 84.405 183.335 ;
        RECT 82.250 182.905 82.915 183.075 ;
        RECT 82.245 182.355 82.575 182.735 ;
        RECT 82.745 182.615 82.915 182.905 ;
        RECT 83.450 182.560 83.695 183.165 ;
        RECT 83.915 182.355 84.425 182.890 ;
        RECT 84.605 182.525 84.795 183.885 ;
        RECT 84.965 183.545 85.240 183.685 ;
        RECT 84.965 183.375 85.245 183.545 ;
        RECT 84.965 182.525 85.240 183.375 ;
        RECT 85.445 183.085 85.615 183.885 ;
        RECT 85.785 183.095 85.955 184.225 ;
        RECT 86.125 183.595 86.295 184.565 ;
        RECT 86.465 183.765 86.635 184.905 ;
        RECT 86.805 183.765 87.140 184.735 ;
        RECT 86.125 183.265 86.320 183.595 ;
        RECT 86.545 183.265 86.800 183.595 ;
        RECT 86.545 183.095 86.715 183.265 ;
        RECT 86.970 183.095 87.140 183.765 ;
        RECT 87.315 183.740 87.605 184.905 ;
        RECT 87.815 183.765 88.045 184.905 ;
        RECT 88.215 183.755 88.545 184.735 ;
        RECT 88.715 183.765 88.925 184.905 ;
        RECT 87.795 183.345 88.125 183.595 ;
        RECT 85.785 182.925 86.715 183.095 ;
        RECT 85.785 182.890 85.960 182.925 ;
        RECT 85.430 182.525 85.960 182.890 ;
        RECT 86.385 182.355 86.715 182.755 ;
        RECT 86.885 182.525 87.140 183.095 ;
        RECT 87.315 182.355 87.605 183.080 ;
        RECT 87.815 182.355 88.045 183.175 ;
        RECT 88.295 183.155 88.545 183.755 ;
        RECT 89.160 183.715 89.415 184.595 ;
        RECT 89.585 183.765 89.890 184.905 ;
        RECT 90.230 184.525 90.560 184.905 ;
        RECT 90.740 184.355 90.910 184.645 ;
        RECT 91.080 184.445 91.330 184.905 ;
        RECT 90.110 184.185 90.910 184.355 ;
        RECT 91.500 184.395 92.370 184.735 ;
        RECT 88.215 182.525 88.545 183.155 ;
        RECT 88.715 182.355 88.925 183.175 ;
        RECT 89.160 183.065 89.370 183.715 ;
        RECT 90.110 183.595 90.280 184.185 ;
        RECT 91.500 184.015 91.670 184.395 ;
        RECT 92.605 184.275 92.775 184.735 ;
        RECT 92.945 184.445 93.315 184.905 ;
        RECT 93.610 184.305 93.780 184.645 ;
        RECT 93.950 184.475 94.280 184.905 ;
        RECT 94.515 184.305 94.685 184.645 ;
        RECT 90.450 183.845 91.670 184.015 ;
        RECT 91.840 183.935 92.300 184.225 ;
        RECT 92.605 184.105 93.165 184.275 ;
        RECT 93.610 184.135 94.685 184.305 ;
        RECT 94.855 184.405 95.535 184.735 ;
        RECT 95.750 184.405 96.000 184.735 ;
        RECT 96.170 184.445 96.420 184.905 ;
        RECT 92.995 183.965 93.165 184.105 ;
        RECT 91.840 183.925 92.805 183.935 ;
        RECT 91.500 183.755 91.670 183.845 ;
        RECT 92.130 183.765 92.805 183.925 ;
        RECT 89.540 183.565 90.280 183.595 ;
        RECT 89.540 183.265 90.455 183.565 ;
        RECT 90.130 183.090 90.455 183.265 ;
        RECT 89.160 182.535 89.415 183.065 ;
        RECT 89.585 182.355 89.890 182.815 ;
        RECT 90.135 182.735 90.455 183.090 ;
        RECT 90.625 183.305 91.165 183.675 ;
        RECT 91.500 183.585 91.905 183.755 ;
        RECT 90.625 182.905 90.865 183.305 ;
        RECT 91.345 183.135 91.565 183.415 ;
        RECT 91.035 182.965 91.565 183.135 ;
        RECT 91.035 182.735 91.205 182.965 ;
        RECT 91.735 182.805 91.905 183.585 ;
        RECT 92.075 182.975 92.425 183.595 ;
        RECT 92.595 182.975 92.805 183.765 ;
        RECT 92.995 183.795 94.495 183.965 ;
        RECT 92.995 183.105 93.165 183.795 ;
        RECT 94.855 183.625 95.025 184.405 ;
        RECT 95.830 184.275 96.000 184.405 ;
        RECT 93.335 183.455 95.025 183.625 ;
        RECT 95.195 183.845 95.660 184.235 ;
        RECT 95.830 184.105 96.225 184.275 ;
        RECT 93.335 183.275 93.505 183.455 ;
        RECT 90.135 182.565 91.205 182.735 ;
        RECT 91.375 182.355 91.565 182.795 ;
        RECT 91.735 182.525 92.685 182.805 ;
        RECT 92.995 182.715 93.255 183.105 ;
        RECT 93.675 183.035 94.465 183.285 ;
        RECT 92.905 182.545 93.255 182.715 ;
        RECT 93.465 182.355 93.795 182.815 ;
        RECT 94.670 182.745 94.840 183.455 ;
        RECT 95.195 183.255 95.365 183.845 ;
        RECT 95.010 183.035 95.365 183.255 ;
        RECT 95.535 183.035 95.885 183.655 ;
        RECT 96.055 182.745 96.225 184.105 ;
        RECT 96.590 183.935 96.915 184.720 ;
        RECT 96.395 182.885 96.855 183.935 ;
        RECT 94.670 182.575 95.525 182.745 ;
        RECT 95.730 182.575 96.225 182.745 ;
        RECT 96.395 182.355 96.725 182.715 ;
        RECT 97.085 182.615 97.255 184.735 ;
        RECT 97.425 184.405 97.755 184.905 ;
        RECT 97.925 184.235 98.180 184.735 ;
        RECT 97.430 184.065 98.180 184.235 ;
        RECT 97.430 183.075 97.660 184.065 ;
        RECT 97.830 183.245 98.180 183.895 ;
        RECT 99.280 183.715 99.535 184.595 ;
        RECT 99.705 183.765 100.010 184.905 ;
        RECT 100.350 184.525 100.680 184.905 ;
        RECT 100.860 184.355 101.030 184.645 ;
        RECT 101.200 184.445 101.450 184.905 ;
        RECT 100.230 184.185 101.030 184.355 ;
        RECT 101.620 184.395 102.490 184.735 ;
        RECT 97.430 182.905 98.180 183.075 ;
        RECT 97.425 182.355 97.755 182.735 ;
        RECT 97.925 182.615 98.180 182.905 ;
        RECT 99.280 183.065 99.490 183.715 ;
        RECT 100.230 183.595 100.400 184.185 ;
        RECT 101.620 184.015 101.790 184.395 ;
        RECT 102.725 184.275 102.895 184.735 ;
        RECT 103.065 184.445 103.435 184.905 ;
        RECT 103.730 184.305 103.900 184.645 ;
        RECT 104.070 184.475 104.400 184.905 ;
        RECT 104.635 184.305 104.805 184.645 ;
        RECT 100.570 183.845 101.790 184.015 ;
        RECT 101.960 183.935 102.420 184.225 ;
        RECT 102.725 184.105 103.285 184.275 ;
        RECT 103.730 184.135 104.805 184.305 ;
        RECT 104.975 184.405 105.655 184.735 ;
        RECT 105.870 184.405 106.120 184.735 ;
        RECT 106.290 184.445 106.540 184.905 ;
        RECT 103.115 183.965 103.285 184.105 ;
        RECT 101.960 183.925 102.925 183.935 ;
        RECT 101.620 183.755 101.790 183.845 ;
        RECT 102.250 183.765 102.925 183.925 ;
        RECT 99.660 183.565 100.400 183.595 ;
        RECT 99.660 183.265 100.575 183.565 ;
        RECT 100.250 183.090 100.575 183.265 ;
        RECT 99.280 182.535 99.535 183.065 ;
        RECT 99.705 182.355 100.010 182.815 ;
        RECT 100.255 182.735 100.575 183.090 ;
        RECT 100.745 183.305 101.285 183.675 ;
        RECT 101.620 183.585 102.025 183.755 ;
        RECT 100.745 182.905 100.985 183.305 ;
        RECT 101.465 183.135 101.685 183.415 ;
        RECT 101.155 182.965 101.685 183.135 ;
        RECT 101.155 182.735 101.325 182.965 ;
        RECT 101.855 182.805 102.025 183.585 ;
        RECT 102.195 182.975 102.545 183.595 ;
        RECT 102.715 182.975 102.925 183.765 ;
        RECT 103.115 183.795 104.615 183.965 ;
        RECT 103.115 183.105 103.285 183.795 ;
        RECT 104.975 183.625 105.145 184.405 ;
        RECT 105.950 184.275 106.120 184.405 ;
        RECT 103.455 183.455 105.145 183.625 ;
        RECT 105.315 183.845 105.780 184.235 ;
        RECT 105.950 184.105 106.345 184.275 ;
        RECT 103.455 183.275 103.625 183.455 ;
        RECT 100.255 182.565 101.325 182.735 ;
        RECT 101.495 182.355 101.685 182.795 ;
        RECT 101.855 182.525 102.805 182.805 ;
        RECT 103.115 182.715 103.375 183.105 ;
        RECT 103.795 183.035 104.585 183.285 ;
        RECT 103.025 182.545 103.375 182.715 ;
        RECT 103.585 182.355 103.915 182.815 ;
        RECT 104.790 182.745 104.960 183.455 ;
        RECT 105.315 183.255 105.485 183.845 ;
        RECT 105.130 183.035 105.485 183.255 ;
        RECT 105.655 183.035 106.005 183.655 ;
        RECT 106.175 182.745 106.345 184.105 ;
        RECT 106.710 183.935 107.035 184.720 ;
        RECT 106.515 182.885 106.975 183.935 ;
        RECT 104.790 182.575 105.645 182.745 ;
        RECT 105.850 182.575 106.345 182.745 ;
        RECT 106.515 182.355 106.845 182.715 ;
        RECT 107.205 182.615 107.375 184.735 ;
        RECT 107.545 184.405 107.875 184.905 ;
        RECT 108.045 184.235 108.300 184.735 ;
        RECT 107.550 184.065 108.300 184.235 ;
        RECT 107.550 183.075 107.780 184.065 ;
        RECT 107.950 183.245 108.300 183.895 ;
        RECT 108.515 183.765 108.745 184.905 ;
        RECT 108.915 183.755 109.245 184.735 ;
        RECT 109.415 183.765 109.625 184.905 ;
        RECT 110.315 183.815 111.985 184.905 ;
        RECT 112.155 183.815 113.365 184.905 ;
        RECT 108.495 183.345 108.825 183.595 ;
        RECT 107.550 182.905 108.300 183.075 ;
        RECT 107.545 182.355 107.875 182.735 ;
        RECT 108.045 182.615 108.300 182.905 ;
        RECT 108.515 182.355 108.745 183.175 ;
        RECT 108.995 183.155 109.245 183.755 ;
        RECT 110.315 183.295 111.065 183.815 ;
        RECT 108.915 182.525 109.245 183.155 ;
        RECT 109.415 182.355 109.625 183.175 ;
        RECT 111.235 183.125 111.985 183.645 ;
        RECT 112.155 183.275 112.675 183.815 ;
        RECT 110.315 182.355 111.985 183.125 ;
        RECT 112.845 183.105 113.365 183.645 ;
        RECT 112.155 182.355 113.365 183.105 ;
        RECT 15.010 182.185 113.450 182.355 ;
        RECT 15.095 181.435 16.305 182.185 ;
        RECT 16.475 181.435 17.685 182.185 ;
        RECT 15.095 180.895 15.615 181.435 ;
        RECT 15.785 180.725 16.305 181.265 ;
        RECT 15.095 179.635 16.305 180.725 ;
        RECT 16.475 180.725 16.995 181.265 ;
        RECT 17.165 180.895 17.685 181.435 ;
        RECT 17.915 181.365 18.125 182.185 ;
        RECT 18.295 181.385 18.625 182.015 ;
        RECT 18.295 180.785 18.545 181.385 ;
        RECT 18.795 181.365 19.025 182.185 ;
        RECT 19.350 181.555 19.635 182.015 ;
        RECT 19.805 181.725 20.075 182.185 ;
        RECT 19.350 181.385 20.305 181.555 ;
        RECT 18.715 180.945 19.045 181.195 ;
        RECT 16.475 179.635 17.685 180.725 ;
        RECT 17.915 179.635 18.125 180.775 ;
        RECT 18.295 179.805 18.625 180.785 ;
        RECT 18.795 179.635 19.025 180.775 ;
        RECT 19.235 180.655 19.925 181.215 ;
        RECT 20.095 180.485 20.305 181.385 ;
        RECT 19.350 180.265 20.305 180.485 ;
        RECT 20.475 181.215 20.875 182.015 ;
        RECT 21.065 181.555 21.345 182.015 ;
        RECT 21.865 181.725 22.190 182.185 ;
        RECT 21.065 181.385 22.190 181.555 ;
        RECT 22.360 181.445 22.745 182.015 ;
        RECT 22.915 181.460 23.205 182.185 ;
        RECT 23.465 181.635 23.635 182.015 ;
        RECT 23.815 181.805 24.145 182.185 ;
        RECT 23.465 181.465 24.130 181.635 ;
        RECT 24.325 181.510 24.585 182.015 ;
        RECT 21.740 181.275 22.190 181.385 ;
        RECT 20.475 180.655 21.570 181.215 ;
        RECT 21.740 180.945 22.295 181.275 ;
        RECT 19.350 179.805 19.635 180.265 ;
        RECT 19.805 179.635 20.075 180.095 ;
        RECT 20.475 179.805 20.875 180.655 ;
        RECT 21.740 180.485 22.190 180.945 ;
        RECT 22.465 180.775 22.745 181.445 ;
        RECT 23.395 180.915 23.725 181.285 ;
        RECT 23.960 181.210 24.130 181.465 ;
        RECT 23.960 180.880 24.245 181.210 ;
        RECT 21.065 180.265 22.190 180.485 ;
        RECT 21.065 179.805 21.345 180.265 ;
        RECT 21.865 179.635 22.190 180.095 ;
        RECT 22.360 179.805 22.745 180.775 ;
        RECT 22.915 179.635 23.205 180.800 ;
        RECT 23.960 180.735 24.130 180.880 ;
        RECT 23.465 180.565 24.130 180.735 ;
        RECT 24.415 180.710 24.585 181.510 ;
        RECT 24.870 181.555 25.155 182.015 ;
        RECT 25.325 181.725 25.595 182.185 ;
        RECT 24.870 181.385 25.825 181.555 ;
        RECT 23.465 179.805 23.635 180.565 ;
        RECT 23.815 179.635 24.145 180.395 ;
        RECT 24.315 179.805 24.585 180.710 ;
        RECT 24.755 180.655 25.445 181.215 ;
        RECT 25.615 180.485 25.825 181.385 ;
        RECT 24.870 180.265 25.825 180.485 ;
        RECT 25.995 181.215 26.395 182.015 ;
        RECT 26.585 181.555 26.865 182.015 ;
        RECT 27.385 181.725 27.710 182.185 ;
        RECT 26.585 181.385 27.710 181.555 ;
        RECT 27.880 181.445 28.265 182.015 ;
        RECT 27.260 181.275 27.710 181.385 ;
        RECT 25.995 180.655 27.090 181.215 ;
        RECT 27.260 180.945 27.815 181.275 ;
        RECT 24.870 179.805 25.155 180.265 ;
        RECT 25.325 179.635 25.595 180.095 ;
        RECT 25.995 179.805 26.395 180.655 ;
        RECT 27.260 180.485 27.710 180.945 ;
        RECT 27.985 180.775 28.265 181.445 ;
        RECT 26.585 180.265 27.710 180.485 ;
        RECT 26.585 179.805 26.865 180.265 ;
        RECT 27.385 179.635 27.710 180.095 ;
        RECT 27.880 179.805 28.265 180.775 ;
        RECT 28.440 181.445 28.695 182.015 ;
        RECT 28.865 181.785 29.195 182.185 ;
        RECT 29.620 181.650 30.150 182.015 ;
        RECT 29.620 181.615 29.795 181.650 ;
        RECT 28.865 181.445 29.795 181.615 ;
        RECT 30.340 181.505 30.615 182.015 ;
        RECT 28.440 180.775 28.610 181.445 ;
        RECT 28.865 181.275 29.035 181.445 ;
        RECT 28.780 180.945 29.035 181.275 ;
        RECT 29.260 180.945 29.455 181.275 ;
        RECT 28.440 179.805 28.775 180.775 ;
        RECT 28.945 179.635 29.115 180.775 ;
        RECT 29.285 179.975 29.455 180.945 ;
        RECT 29.625 180.315 29.795 181.445 ;
        RECT 29.965 180.655 30.135 181.455 ;
        RECT 30.335 181.335 30.615 181.505 ;
        RECT 30.340 180.855 30.615 181.335 ;
        RECT 30.785 180.655 30.975 182.015 ;
        RECT 31.155 181.650 31.665 182.185 ;
        RECT 31.885 181.375 32.130 181.980 ;
        RECT 33.040 181.475 33.295 182.005 ;
        RECT 33.465 181.725 33.770 182.185 ;
        RECT 34.015 181.805 35.085 181.975 ;
        RECT 31.175 181.205 32.405 181.375 ;
        RECT 29.965 180.485 30.975 180.655 ;
        RECT 31.145 180.640 31.895 180.830 ;
        RECT 29.625 180.145 30.750 180.315 ;
        RECT 31.145 179.975 31.315 180.640 ;
        RECT 32.065 180.395 32.405 181.205 ;
        RECT 29.285 179.805 31.315 179.975 ;
        RECT 31.485 179.635 31.655 180.395 ;
        RECT 31.890 179.985 32.405 180.395 ;
        RECT 33.040 180.825 33.250 181.475 ;
        RECT 34.015 181.450 34.335 181.805 ;
        RECT 34.010 181.275 34.335 181.450 ;
        RECT 33.420 180.975 34.335 181.275 ;
        RECT 34.505 181.235 34.745 181.635 ;
        RECT 34.915 181.575 35.085 181.805 ;
        RECT 35.255 181.745 35.445 182.185 ;
        RECT 35.615 181.735 36.565 182.015 ;
        RECT 36.785 181.825 37.135 181.995 ;
        RECT 34.915 181.405 35.445 181.575 ;
        RECT 33.420 180.945 34.160 180.975 ;
        RECT 33.040 179.945 33.295 180.825 ;
        RECT 33.465 179.635 33.770 180.775 ;
        RECT 33.990 180.355 34.160 180.945 ;
        RECT 34.505 180.865 35.045 181.235 ;
        RECT 35.225 181.125 35.445 181.405 ;
        RECT 35.615 180.955 35.785 181.735 ;
        RECT 35.380 180.785 35.785 180.955 ;
        RECT 35.955 180.945 36.305 181.565 ;
        RECT 35.380 180.695 35.550 180.785 ;
        RECT 36.475 180.775 36.685 181.565 ;
        RECT 34.330 180.525 35.550 180.695 ;
        RECT 36.010 180.615 36.685 180.775 ;
        RECT 33.990 180.185 34.790 180.355 ;
        RECT 34.110 179.635 34.440 180.015 ;
        RECT 34.620 179.895 34.790 180.185 ;
        RECT 35.380 180.145 35.550 180.525 ;
        RECT 35.720 180.605 36.685 180.615 ;
        RECT 36.875 181.435 37.135 181.825 ;
        RECT 37.345 181.725 37.675 182.185 ;
        RECT 38.550 181.795 39.405 181.965 ;
        RECT 39.610 181.795 40.105 181.965 ;
        RECT 40.275 181.825 40.605 182.185 ;
        RECT 36.875 180.745 37.045 181.435 ;
        RECT 37.215 181.085 37.385 181.265 ;
        RECT 37.555 181.255 38.345 181.505 ;
        RECT 38.550 181.085 38.720 181.795 ;
        RECT 38.890 181.285 39.245 181.505 ;
        RECT 37.215 180.915 38.905 181.085 ;
        RECT 35.720 180.315 36.180 180.605 ;
        RECT 36.875 180.575 38.375 180.745 ;
        RECT 36.875 180.435 37.045 180.575 ;
        RECT 36.485 180.265 37.045 180.435 ;
        RECT 34.960 179.635 35.210 180.095 ;
        RECT 35.380 179.805 36.250 180.145 ;
        RECT 36.485 179.805 36.655 180.265 ;
        RECT 37.490 180.235 38.565 180.405 ;
        RECT 36.825 179.635 37.195 180.095 ;
        RECT 37.490 179.895 37.660 180.235 ;
        RECT 37.830 179.635 38.160 180.065 ;
        RECT 38.395 179.895 38.565 180.235 ;
        RECT 38.735 180.135 38.905 180.915 ;
        RECT 39.075 180.695 39.245 181.285 ;
        RECT 39.415 180.885 39.765 181.505 ;
        RECT 39.075 180.305 39.540 180.695 ;
        RECT 39.935 180.435 40.105 181.795 ;
        RECT 40.275 180.605 40.735 181.655 ;
        RECT 39.710 180.265 40.105 180.435 ;
        RECT 39.710 180.135 39.880 180.265 ;
        RECT 38.735 179.805 39.415 180.135 ;
        RECT 39.630 179.805 39.880 180.135 ;
        RECT 40.050 179.635 40.300 180.095 ;
        RECT 40.470 179.820 40.795 180.605 ;
        RECT 40.965 179.805 41.135 181.925 ;
        RECT 41.305 181.805 41.635 182.185 ;
        RECT 41.805 181.635 42.060 181.925 ;
        RECT 41.310 181.465 42.060 181.635 ;
        RECT 41.310 180.475 41.540 181.465 ;
        RECT 42.235 181.435 43.445 182.185 ;
        RECT 41.710 180.645 42.060 181.295 ;
        RECT 42.235 180.725 42.755 181.265 ;
        RECT 42.925 180.895 43.445 181.435 ;
        RECT 43.675 181.365 43.885 182.185 ;
        RECT 44.055 181.385 44.385 182.015 ;
        RECT 44.055 180.785 44.305 181.385 ;
        RECT 44.555 181.365 44.785 182.185 ;
        RECT 45.110 181.555 45.395 182.015 ;
        RECT 45.565 181.725 45.835 182.185 ;
        RECT 45.110 181.385 46.065 181.555 ;
        RECT 44.475 180.945 44.805 181.195 ;
        RECT 41.310 180.305 42.060 180.475 ;
        RECT 41.305 179.635 41.635 180.135 ;
        RECT 41.805 179.805 42.060 180.305 ;
        RECT 42.235 179.635 43.445 180.725 ;
        RECT 43.675 179.635 43.885 180.775 ;
        RECT 44.055 179.805 44.385 180.785 ;
        RECT 44.555 179.635 44.785 180.775 ;
        RECT 44.995 180.655 45.685 181.215 ;
        RECT 45.855 180.485 46.065 181.385 ;
        RECT 45.110 180.265 46.065 180.485 ;
        RECT 46.235 181.215 46.635 182.015 ;
        RECT 46.825 181.555 47.105 182.015 ;
        RECT 47.625 181.725 47.950 182.185 ;
        RECT 46.825 181.385 47.950 181.555 ;
        RECT 48.120 181.445 48.505 182.015 ;
        RECT 48.675 181.460 48.965 182.185 ;
        RECT 47.500 181.275 47.950 181.385 ;
        RECT 46.235 180.655 47.330 181.215 ;
        RECT 47.500 180.945 48.055 181.275 ;
        RECT 45.110 179.805 45.395 180.265 ;
        RECT 45.565 179.635 45.835 180.095 ;
        RECT 46.235 179.805 46.635 180.655 ;
        RECT 47.500 180.485 47.950 180.945 ;
        RECT 48.225 180.775 48.505 181.445 ;
        RECT 49.135 181.445 49.520 182.015 ;
        RECT 49.690 181.725 50.015 182.185 ;
        RECT 50.535 181.555 50.815 182.015 ;
        RECT 46.825 180.265 47.950 180.485 ;
        RECT 46.825 179.805 47.105 180.265 ;
        RECT 47.625 179.635 47.950 180.095 ;
        RECT 48.120 179.805 48.505 180.775 ;
        RECT 48.675 179.635 48.965 180.800 ;
        RECT 49.135 180.775 49.415 181.445 ;
        RECT 49.690 181.385 50.815 181.555 ;
        RECT 49.690 181.275 50.140 181.385 ;
        RECT 49.585 180.945 50.140 181.275 ;
        RECT 51.005 181.215 51.405 182.015 ;
        RECT 51.805 181.725 52.075 182.185 ;
        RECT 52.245 181.555 52.530 182.015 ;
        RECT 49.135 179.805 49.520 180.775 ;
        RECT 49.690 180.485 50.140 180.945 ;
        RECT 50.310 180.655 51.405 181.215 ;
        RECT 49.690 180.265 50.815 180.485 ;
        RECT 49.690 179.635 50.015 180.095 ;
        RECT 50.535 179.805 50.815 180.265 ;
        RECT 51.005 179.805 51.405 180.655 ;
        RECT 51.575 181.385 52.530 181.555 ;
        RECT 51.575 180.485 51.785 181.385 ;
        RECT 52.875 181.365 53.085 182.185 ;
        RECT 53.255 181.385 53.585 182.015 ;
        RECT 51.955 180.655 52.645 181.215 ;
        RECT 53.255 180.785 53.505 181.385 ;
        RECT 53.755 181.365 53.985 182.185 ;
        RECT 54.195 181.510 54.455 182.015 ;
        RECT 54.635 181.805 54.965 182.185 ;
        RECT 55.145 181.635 55.315 182.015 ;
        RECT 53.675 180.945 54.005 181.195 ;
        RECT 51.575 180.265 52.530 180.485 ;
        RECT 51.805 179.635 52.075 180.095 ;
        RECT 52.245 179.805 52.530 180.265 ;
        RECT 52.875 179.635 53.085 180.775 ;
        RECT 53.255 179.805 53.585 180.785 ;
        RECT 53.755 179.635 53.985 180.775 ;
        RECT 54.195 180.710 54.365 181.510 ;
        RECT 54.650 181.465 55.315 181.635 ;
        RECT 54.650 181.210 54.820 181.465 ;
        RECT 55.575 181.415 57.245 182.185 ;
        RECT 54.535 180.880 54.820 181.210 ;
        RECT 55.055 180.915 55.385 181.285 ;
        RECT 54.650 180.735 54.820 180.880 ;
        RECT 54.195 179.805 54.465 180.710 ;
        RECT 54.650 180.565 55.315 180.735 ;
        RECT 54.635 179.635 54.965 180.395 ;
        RECT 55.145 179.805 55.315 180.565 ;
        RECT 55.575 180.725 56.325 181.245 ;
        RECT 56.495 180.895 57.245 181.415 ;
        RECT 57.505 181.535 57.675 182.015 ;
        RECT 57.855 181.705 58.095 182.185 ;
        RECT 58.345 181.535 58.515 182.015 ;
        RECT 58.685 181.705 59.015 182.185 ;
        RECT 59.185 181.535 59.355 182.015 ;
        RECT 57.505 181.365 58.140 181.535 ;
        RECT 58.345 181.365 59.355 181.535 ;
        RECT 59.525 181.385 59.855 182.185 ;
        RECT 60.215 181.365 60.445 182.185 ;
        RECT 60.615 181.385 60.945 182.015 ;
        RECT 57.970 181.195 58.140 181.365 ;
        RECT 58.855 181.335 59.355 181.365 ;
        RECT 57.420 180.955 57.800 181.195 ;
        RECT 57.970 181.025 58.470 181.195 ;
        RECT 57.970 180.785 58.140 181.025 ;
        RECT 58.860 180.825 59.355 181.335 ;
        RECT 60.195 180.945 60.525 181.195 ;
        RECT 55.575 179.635 57.245 180.725 ;
        RECT 57.425 180.615 58.140 180.785 ;
        RECT 58.345 180.655 59.355 180.825 ;
        RECT 60.695 180.785 60.945 181.385 ;
        RECT 61.115 181.365 61.325 182.185 ;
        RECT 61.645 181.635 61.815 182.015 ;
        RECT 62.030 181.805 62.360 182.185 ;
        RECT 61.645 181.465 62.360 181.635 ;
        RECT 61.555 180.915 61.910 181.285 ;
        RECT 62.190 181.275 62.360 181.465 ;
        RECT 62.530 181.440 62.785 182.015 ;
        RECT 62.190 180.945 62.445 181.275 ;
        RECT 57.425 179.805 57.755 180.615 ;
        RECT 57.925 179.635 58.165 180.435 ;
        RECT 58.345 179.805 58.515 180.655 ;
        RECT 58.685 179.635 59.015 180.435 ;
        RECT 59.185 179.805 59.355 180.655 ;
        RECT 59.525 179.635 59.855 180.785 ;
        RECT 60.215 179.635 60.445 180.775 ;
        RECT 60.615 179.805 60.945 180.785 ;
        RECT 61.115 179.635 61.325 180.775 ;
        RECT 62.190 180.735 62.360 180.945 ;
        RECT 61.645 180.565 62.360 180.735 ;
        RECT 62.615 180.710 62.785 181.440 ;
        RECT 62.960 181.345 63.220 182.185 ;
        RECT 63.665 181.790 63.995 182.185 ;
        RECT 64.165 181.615 64.365 181.970 ;
        RECT 64.535 181.785 64.865 182.185 ;
        RECT 65.035 181.615 65.235 181.960 ;
        RECT 63.395 181.445 65.235 181.615 ;
        RECT 65.405 181.445 65.735 182.185 ;
        RECT 65.970 181.615 66.140 181.865 ;
        RECT 65.970 181.445 66.445 181.615 ;
        RECT 61.645 179.805 61.815 180.565 ;
        RECT 62.030 179.635 62.360 180.395 ;
        RECT 62.530 179.805 62.785 180.710 ;
        RECT 62.960 179.635 63.220 180.785 ;
        RECT 63.395 179.820 63.655 181.445 ;
        RECT 63.835 180.475 64.055 181.275 ;
        RECT 64.295 180.655 64.595 181.275 ;
        RECT 64.765 180.655 65.095 181.275 ;
        RECT 65.265 180.655 65.585 181.275 ;
        RECT 65.755 180.655 66.105 181.275 ;
        RECT 66.275 180.475 66.445 181.445 ;
        RECT 66.730 181.555 67.015 182.015 ;
        RECT 67.185 181.725 67.455 182.185 ;
        RECT 66.730 181.385 67.685 181.555 ;
        RECT 66.615 180.655 67.305 181.215 ;
        RECT 67.475 180.485 67.685 181.385 ;
        RECT 63.835 180.265 66.445 180.475 ;
        RECT 66.730 180.265 67.685 180.485 ;
        RECT 67.855 181.215 68.255 182.015 ;
        RECT 68.445 181.555 68.725 182.015 ;
        RECT 69.245 181.725 69.570 182.185 ;
        RECT 68.445 181.385 69.570 181.555 ;
        RECT 69.740 181.445 70.125 182.015 ;
        RECT 69.120 181.275 69.570 181.385 ;
        RECT 67.855 180.655 68.950 181.215 ;
        RECT 69.120 180.945 69.675 181.275 ;
        RECT 65.405 179.635 65.735 180.085 ;
        RECT 66.730 179.805 67.015 180.265 ;
        RECT 67.185 179.635 67.455 180.095 ;
        RECT 67.855 179.805 68.255 180.655 ;
        RECT 69.120 180.485 69.570 180.945 ;
        RECT 69.845 180.775 70.125 181.445 ;
        RECT 70.570 181.375 70.815 181.980 ;
        RECT 71.035 181.650 71.545 182.185 ;
        RECT 68.445 180.265 69.570 180.485 ;
        RECT 68.445 179.805 68.725 180.265 ;
        RECT 69.245 179.635 69.570 180.095 ;
        RECT 69.740 179.805 70.125 180.775 ;
        RECT 70.295 181.205 71.525 181.375 ;
        RECT 70.295 180.395 70.635 181.205 ;
        RECT 70.805 180.640 71.555 180.830 ;
        RECT 70.295 179.985 70.810 180.395 ;
        RECT 71.045 179.635 71.215 180.395 ;
        RECT 71.385 179.975 71.555 180.640 ;
        RECT 71.725 180.655 71.915 182.015 ;
        RECT 72.085 181.505 72.360 182.015 ;
        RECT 72.550 181.650 73.080 182.015 ;
        RECT 73.505 181.785 73.835 182.185 ;
        RECT 72.905 181.615 73.080 181.650 ;
        RECT 72.085 181.335 72.365 181.505 ;
        RECT 72.085 180.855 72.360 181.335 ;
        RECT 72.565 180.655 72.735 181.455 ;
        RECT 71.725 180.485 72.735 180.655 ;
        RECT 72.905 181.445 73.835 181.615 ;
        RECT 74.005 181.445 74.260 182.015 ;
        RECT 74.435 181.460 74.725 182.185 ;
        RECT 74.900 181.475 75.155 182.005 ;
        RECT 75.325 181.725 75.630 182.185 ;
        RECT 75.875 181.805 76.945 181.975 ;
        RECT 72.905 180.315 73.075 181.445 ;
        RECT 73.665 181.275 73.835 181.445 ;
        RECT 71.950 180.145 73.075 180.315 ;
        RECT 73.245 180.945 73.440 181.275 ;
        RECT 73.665 180.945 73.920 181.275 ;
        RECT 73.245 179.975 73.415 180.945 ;
        RECT 74.090 180.775 74.260 181.445 ;
        RECT 74.900 180.825 75.110 181.475 ;
        RECT 75.875 181.450 76.195 181.805 ;
        RECT 75.870 181.275 76.195 181.450 ;
        RECT 75.280 180.975 76.195 181.275 ;
        RECT 76.365 181.235 76.605 181.635 ;
        RECT 76.775 181.575 76.945 181.805 ;
        RECT 77.115 181.745 77.305 182.185 ;
        RECT 77.475 181.735 78.425 182.015 ;
        RECT 78.645 181.825 78.995 181.995 ;
        RECT 76.775 181.405 77.305 181.575 ;
        RECT 75.280 180.945 76.020 180.975 ;
        RECT 71.385 179.805 73.415 179.975 ;
        RECT 73.585 179.635 73.755 180.775 ;
        RECT 73.925 179.805 74.260 180.775 ;
        RECT 74.435 179.635 74.725 180.800 ;
        RECT 74.900 179.945 75.155 180.825 ;
        RECT 75.325 179.635 75.630 180.775 ;
        RECT 75.850 180.355 76.020 180.945 ;
        RECT 76.365 180.865 76.905 181.235 ;
        RECT 77.085 181.125 77.305 181.405 ;
        RECT 77.475 180.955 77.645 181.735 ;
        RECT 77.240 180.785 77.645 180.955 ;
        RECT 77.815 180.945 78.165 181.565 ;
        RECT 77.240 180.695 77.410 180.785 ;
        RECT 78.335 180.775 78.545 181.565 ;
        RECT 76.190 180.525 77.410 180.695 ;
        RECT 77.870 180.615 78.545 180.775 ;
        RECT 75.850 180.185 76.650 180.355 ;
        RECT 75.970 179.635 76.300 180.015 ;
        RECT 76.480 179.895 76.650 180.185 ;
        RECT 77.240 180.145 77.410 180.525 ;
        RECT 77.580 180.605 78.545 180.615 ;
        RECT 78.735 181.435 78.995 181.825 ;
        RECT 79.205 181.725 79.535 182.185 ;
        RECT 80.410 181.795 81.265 181.965 ;
        RECT 81.470 181.795 81.965 181.965 ;
        RECT 82.135 181.825 82.465 182.185 ;
        RECT 78.735 180.745 78.905 181.435 ;
        RECT 79.075 181.085 79.245 181.265 ;
        RECT 79.415 181.255 80.205 181.505 ;
        RECT 80.410 181.085 80.580 181.795 ;
        RECT 80.750 181.285 81.105 181.505 ;
        RECT 79.075 180.915 80.765 181.085 ;
        RECT 77.580 180.315 78.040 180.605 ;
        RECT 78.735 180.575 80.235 180.745 ;
        RECT 78.735 180.435 78.905 180.575 ;
        RECT 78.345 180.265 78.905 180.435 ;
        RECT 76.820 179.635 77.070 180.095 ;
        RECT 77.240 179.805 78.110 180.145 ;
        RECT 78.345 179.805 78.515 180.265 ;
        RECT 79.350 180.235 80.425 180.405 ;
        RECT 78.685 179.635 79.055 180.095 ;
        RECT 79.350 179.895 79.520 180.235 ;
        RECT 79.690 179.635 80.020 180.065 ;
        RECT 80.255 179.895 80.425 180.235 ;
        RECT 80.595 180.135 80.765 180.915 ;
        RECT 80.935 180.695 81.105 181.285 ;
        RECT 81.275 180.885 81.625 181.505 ;
        RECT 80.935 180.305 81.400 180.695 ;
        RECT 81.795 180.435 81.965 181.795 ;
        RECT 82.135 180.605 82.595 181.655 ;
        RECT 81.570 180.265 81.965 180.435 ;
        RECT 81.570 180.135 81.740 180.265 ;
        RECT 80.595 179.805 81.275 180.135 ;
        RECT 81.490 179.805 81.740 180.135 ;
        RECT 81.910 179.635 82.160 180.095 ;
        RECT 82.330 179.820 82.655 180.605 ;
        RECT 82.825 179.805 82.995 181.925 ;
        RECT 83.165 181.805 83.495 182.185 ;
        RECT 83.665 181.635 83.920 181.925 ;
        RECT 83.170 181.465 83.920 181.635 ;
        RECT 84.100 181.475 84.355 182.005 ;
        RECT 84.525 181.725 84.830 182.185 ;
        RECT 85.075 181.805 86.145 181.975 ;
        RECT 83.170 180.475 83.400 181.465 ;
        RECT 83.570 180.645 83.920 181.295 ;
        RECT 84.100 180.825 84.310 181.475 ;
        RECT 85.075 181.450 85.395 181.805 ;
        RECT 85.070 181.275 85.395 181.450 ;
        RECT 84.480 180.975 85.395 181.275 ;
        RECT 85.565 181.235 85.805 181.635 ;
        RECT 85.975 181.575 86.145 181.805 ;
        RECT 86.315 181.745 86.505 182.185 ;
        RECT 86.675 181.735 87.625 182.015 ;
        RECT 87.845 181.825 88.195 181.995 ;
        RECT 85.975 181.405 86.505 181.575 ;
        RECT 84.480 180.945 85.220 180.975 ;
        RECT 83.170 180.305 83.920 180.475 ;
        RECT 83.165 179.635 83.495 180.135 ;
        RECT 83.665 179.805 83.920 180.305 ;
        RECT 84.100 179.945 84.355 180.825 ;
        RECT 84.525 179.635 84.830 180.775 ;
        RECT 85.050 180.355 85.220 180.945 ;
        RECT 85.565 180.865 86.105 181.235 ;
        RECT 86.285 181.125 86.505 181.405 ;
        RECT 86.675 180.955 86.845 181.735 ;
        RECT 86.440 180.785 86.845 180.955 ;
        RECT 87.015 180.945 87.365 181.565 ;
        RECT 86.440 180.695 86.610 180.785 ;
        RECT 87.535 180.775 87.745 181.565 ;
        RECT 85.390 180.525 86.610 180.695 ;
        RECT 87.070 180.615 87.745 180.775 ;
        RECT 85.050 180.185 85.850 180.355 ;
        RECT 85.170 179.635 85.500 180.015 ;
        RECT 85.680 179.895 85.850 180.185 ;
        RECT 86.440 180.145 86.610 180.525 ;
        RECT 86.780 180.605 87.745 180.615 ;
        RECT 87.935 181.435 88.195 181.825 ;
        RECT 88.405 181.725 88.735 182.185 ;
        RECT 89.610 181.795 90.465 181.965 ;
        RECT 90.670 181.795 91.165 181.965 ;
        RECT 91.335 181.825 91.665 182.185 ;
        RECT 87.935 180.745 88.105 181.435 ;
        RECT 88.275 181.085 88.445 181.265 ;
        RECT 88.615 181.255 89.405 181.505 ;
        RECT 89.610 181.085 89.780 181.795 ;
        RECT 89.950 181.285 90.305 181.505 ;
        RECT 88.275 180.915 89.965 181.085 ;
        RECT 86.780 180.315 87.240 180.605 ;
        RECT 87.935 180.575 89.435 180.745 ;
        RECT 87.935 180.435 88.105 180.575 ;
        RECT 87.545 180.265 88.105 180.435 ;
        RECT 86.020 179.635 86.270 180.095 ;
        RECT 86.440 179.805 87.310 180.145 ;
        RECT 87.545 179.805 87.715 180.265 ;
        RECT 88.550 180.235 89.625 180.405 ;
        RECT 87.885 179.635 88.255 180.095 ;
        RECT 88.550 179.895 88.720 180.235 ;
        RECT 88.890 179.635 89.220 180.065 ;
        RECT 89.455 179.895 89.625 180.235 ;
        RECT 89.795 180.135 89.965 180.915 ;
        RECT 90.135 180.695 90.305 181.285 ;
        RECT 90.475 180.885 90.825 181.505 ;
        RECT 90.135 180.305 90.600 180.695 ;
        RECT 90.995 180.435 91.165 181.795 ;
        RECT 91.335 180.605 91.795 181.655 ;
        RECT 90.770 180.265 91.165 180.435 ;
        RECT 90.770 180.135 90.940 180.265 ;
        RECT 89.795 179.805 90.475 180.135 ;
        RECT 90.690 179.805 90.940 180.135 ;
        RECT 91.110 179.635 91.360 180.095 ;
        RECT 91.530 179.820 91.855 180.605 ;
        RECT 92.025 179.805 92.195 181.925 ;
        RECT 92.365 181.805 92.695 182.185 ;
        RECT 92.865 181.635 93.120 181.925 ;
        RECT 92.370 181.465 93.120 181.635 ;
        RECT 93.295 181.510 93.555 182.015 ;
        RECT 93.735 181.805 94.065 182.185 ;
        RECT 94.245 181.635 94.415 182.015 ;
        RECT 92.370 180.475 92.600 181.465 ;
        RECT 92.770 180.645 93.120 181.295 ;
        RECT 93.295 180.710 93.465 181.510 ;
        RECT 93.750 181.465 94.415 181.635 ;
        RECT 94.765 181.635 94.935 182.015 ;
        RECT 95.115 181.805 95.445 182.185 ;
        RECT 94.765 181.465 95.430 181.635 ;
        RECT 95.625 181.510 95.885 182.015 ;
        RECT 93.750 181.210 93.920 181.465 ;
        RECT 93.635 180.880 93.920 181.210 ;
        RECT 94.155 180.915 94.485 181.285 ;
        RECT 94.695 180.915 95.025 181.285 ;
        RECT 95.260 181.210 95.430 181.465 ;
        RECT 93.750 180.735 93.920 180.880 ;
        RECT 95.260 180.880 95.545 181.210 ;
        RECT 95.260 180.735 95.430 180.880 ;
        RECT 92.370 180.305 93.120 180.475 ;
        RECT 92.365 179.635 92.695 180.135 ;
        RECT 92.865 179.805 93.120 180.305 ;
        RECT 93.295 179.805 93.565 180.710 ;
        RECT 93.750 180.565 94.415 180.735 ;
        RECT 93.735 179.635 94.065 180.395 ;
        RECT 94.245 179.805 94.415 180.565 ;
        RECT 94.765 180.565 95.430 180.735 ;
        RECT 95.715 180.710 95.885 181.510 ;
        RECT 96.330 181.375 96.575 181.980 ;
        RECT 96.795 181.650 97.305 182.185 ;
        RECT 94.765 179.805 94.935 180.565 ;
        RECT 95.115 179.635 95.445 180.395 ;
        RECT 95.615 179.805 95.885 180.710 ;
        RECT 96.055 181.205 97.285 181.375 ;
        RECT 96.055 180.395 96.395 181.205 ;
        RECT 96.565 180.640 97.315 180.830 ;
        RECT 96.055 179.985 96.570 180.395 ;
        RECT 96.805 179.635 96.975 180.395 ;
        RECT 97.145 179.975 97.315 180.640 ;
        RECT 97.485 180.655 97.675 182.015 ;
        RECT 97.845 181.165 98.120 182.015 ;
        RECT 98.310 181.650 98.840 182.015 ;
        RECT 99.265 181.785 99.595 182.185 ;
        RECT 98.665 181.615 98.840 181.650 ;
        RECT 97.845 180.995 98.125 181.165 ;
        RECT 97.845 180.855 98.120 180.995 ;
        RECT 98.325 180.655 98.495 181.455 ;
        RECT 97.485 180.485 98.495 180.655 ;
        RECT 98.665 181.445 99.595 181.615 ;
        RECT 99.765 181.445 100.020 182.015 ;
        RECT 100.195 181.460 100.485 182.185 ;
        RECT 98.665 180.315 98.835 181.445 ;
        RECT 99.425 181.275 99.595 181.445 ;
        RECT 97.710 180.145 98.835 180.315 ;
        RECT 99.005 180.945 99.200 181.275 ;
        RECT 99.425 180.945 99.680 181.275 ;
        RECT 99.005 179.975 99.175 180.945 ;
        RECT 99.850 180.775 100.020 181.445 ;
        RECT 100.930 181.375 101.175 181.980 ;
        RECT 101.395 181.650 101.905 182.185 ;
        RECT 100.655 181.205 101.885 181.375 ;
        RECT 97.145 179.805 99.175 179.975 ;
        RECT 99.345 179.635 99.515 180.775 ;
        RECT 99.685 179.805 100.020 180.775 ;
        RECT 100.195 179.635 100.485 180.800 ;
        RECT 100.655 180.395 100.995 181.205 ;
        RECT 101.165 180.640 101.915 180.830 ;
        RECT 100.655 179.985 101.170 180.395 ;
        RECT 101.405 179.635 101.575 180.395 ;
        RECT 101.745 179.975 101.915 180.640 ;
        RECT 102.085 180.655 102.275 182.015 ;
        RECT 102.445 181.845 102.720 182.015 ;
        RECT 102.445 181.675 102.725 181.845 ;
        RECT 102.445 180.855 102.720 181.675 ;
        RECT 102.910 181.650 103.440 182.015 ;
        RECT 103.865 181.785 104.195 182.185 ;
        RECT 103.265 181.615 103.440 181.650 ;
        RECT 102.925 180.655 103.095 181.455 ;
        RECT 102.085 180.485 103.095 180.655 ;
        RECT 103.265 181.445 104.195 181.615 ;
        RECT 104.365 181.445 104.620 182.015 ;
        RECT 103.265 180.315 103.435 181.445 ;
        RECT 104.025 181.275 104.195 181.445 ;
        RECT 102.310 180.145 103.435 180.315 ;
        RECT 103.605 180.945 103.800 181.275 ;
        RECT 104.025 180.945 104.280 181.275 ;
        RECT 103.605 179.975 103.775 180.945 ;
        RECT 104.450 180.775 104.620 181.445 ;
        RECT 101.745 179.805 103.775 179.975 ;
        RECT 103.945 179.635 104.115 180.775 ;
        RECT 104.285 179.805 104.620 180.775 ;
        RECT 104.795 181.445 105.180 182.015 ;
        RECT 105.350 181.725 105.675 182.185 ;
        RECT 106.195 181.555 106.475 182.015 ;
        RECT 104.795 180.775 105.075 181.445 ;
        RECT 105.350 181.385 106.475 181.555 ;
        RECT 105.350 181.275 105.800 181.385 ;
        RECT 105.245 180.945 105.800 181.275 ;
        RECT 106.665 181.215 107.065 182.015 ;
        RECT 107.465 181.725 107.735 182.185 ;
        RECT 107.905 181.555 108.190 182.015 ;
        RECT 104.795 179.805 105.180 180.775 ;
        RECT 105.350 180.485 105.800 180.945 ;
        RECT 105.970 180.655 107.065 181.215 ;
        RECT 105.350 180.265 106.475 180.485 ;
        RECT 105.350 179.635 105.675 180.095 ;
        RECT 106.195 179.805 106.475 180.265 ;
        RECT 106.665 179.805 107.065 180.655 ;
        RECT 107.235 181.385 108.190 181.555 ;
        RECT 108.475 181.445 108.860 182.015 ;
        RECT 109.030 181.725 109.355 182.185 ;
        RECT 109.875 181.555 110.155 182.015 ;
        RECT 107.235 180.485 107.445 181.385 ;
        RECT 107.615 180.655 108.305 181.215 ;
        RECT 108.475 180.775 108.755 181.445 ;
        RECT 109.030 181.385 110.155 181.555 ;
        RECT 109.030 181.275 109.480 181.385 ;
        RECT 108.925 180.945 109.480 181.275 ;
        RECT 110.345 181.215 110.745 182.015 ;
        RECT 111.145 181.725 111.415 182.185 ;
        RECT 111.585 181.555 111.870 182.015 ;
        RECT 107.235 180.265 108.190 180.485 ;
        RECT 107.465 179.635 107.735 180.095 ;
        RECT 107.905 179.805 108.190 180.265 ;
        RECT 108.475 179.805 108.860 180.775 ;
        RECT 109.030 180.485 109.480 180.945 ;
        RECT 109.650 180.655 110.745 181.215 ;
        RECT 109.030 180.265 110.155 180.485 ;
        RECT 109.030 179.635 109.355 180.095 ;
        RECT 109.875 179.805 110.155 180.265 ;
        RECT 110.345 179.805 110.745 180.655 ;
        RECT 110.915 181.385 111.870 181.555 ;
        RECT 112.155 181.435 113.365 182.185 ;
        RECT 110.915 180.485 111.125 181.385 ;
        RECT 111.295 180.655 111.985 181.215 ;
        RECT 112.155 180.725 112.675 181.265 ;
        RECT 112.845 180.895 113.365 181.435 ;
        RECT 110.915 180.265 111.870 180.485 ;
        RECT 111.145 179.635 111.415 180.095 ;
        RECT 111.585 179.805 111.870 180.265 ;
        RECT 112.155 179.635 113.365 180.725 ;
        RECT 15.010 179.465 113.450 179.635 ;
        RECT 15.095 178.375 16.305 179.465 ;
        RECT 15.095 177.665 15.615 178.205 ;
        RECT 15.785 177.835 16.305 178.375 ;
        RECT 16.475 178.375 18.145 179.465 ;
        RECT 18.430 178.835 18.715 179.295 ;
        RECT 18.885 179.005 19.155 179.465 ;
        RECT 18.430 178.615 19.385 178.835 ;
        RECT 16.475 177.855 17.225 178.375 ;
        RECT 17.395 177.685 18.145 178.205 ;
        RECT 18.315 177.885 19.005 178.445 ;
        RECT 19.175 177.715 19.385 178.615 ;
        RECT 15.095 176.915 16.305 177.665 ;
        RECT 16.475 176.915 18.145 177.685 ;
        RECT 18.430 177.545 19.385 177.715 ;
        RECT 19.555 178.445 19.955 179.295 ;
        RECT 20.145 178.835 20.425 179.295 ;
        RECT 20.945 179.005 21.270 179.465 ;
        RECT 20.145 178.615 21.270 178.835 ;
        RECT 19.555 177.885 20.650 178.445 ;
        RECT 20.820 178.155 21.270 178.615 ;
        RECT 21.440 178.325 21.825 179.295 ;
        RECT 18.430 177.085 18.715 177.545 ;
        RECT 18.885 176.915 19.155 177.375 ;
        RECT 19.555 177.085 19.955 177.885 ;
        RECT 20.820 177.825 21.375 178.155 ;
        RECT 20.820 177.715 21.270 177.825 ;
        RECT 20.145 177.545 21.270 177.715 ;
        RECT 21.545 177.655 21.825 178.325 ;
        RECT 20.145 177.085 20.425 177.545 ;
        RECT 20.945 176.915 21.270 177.375 ;
        RECT 21.440 177.085 21.825 177.655 ;
        RECT 22.000 178.275 22.255 179.155 ;
        RECT 22.425 178.325 22.730 179.465 ;
        RECT 23.070 179.085 23.400 179.465 ;
        RECT 23.580 178.915 23.750 179.205 ;
        RECT 23.920 179.005 24.170 179.465 ;
        RECT 22.950 178.745 23.750 178.915 ;
        RECT 24.340 178.955 25.210 179.295 ;
        RECT 22.000 177.625 22.210 178.275 ;
        RECT 22.950 178.155 23.120 178.745 ;
        RECT 24.340 178.575 24.510 178.955 ;
        RECT 25.445 178.835 25.615 179.295 ;
        RECT 25.785 179.005 26.155 179.465 ;
        RECT 26.450 178.865 26.620 179.205 ;
        RECT 26.790 179.035 27.120 179.465 ;
        RECT 27.355 178.865 27.525 179.205 ;
        RECT 23.290 178.405 24.510 178.575 ;
        RECT 24.680 178.495 25.140 178.785 ;
        RECT 25.445 178.665 26.005 178.835 ;
        RECT 26.450 178.695 27.525 178.865 ;
        RECT 27.695 178.965 28.375 179.295 ;
        RECT 28.590 178.965 28.840 179.295 ;
        RECT 29.010 179.005 29.260 179.465 ;
        RECT 25.835 178.525 26.005 178.665 ;
        RECT 24.680 178.485 25.645 178.495 ;
        RECT 24.340 178.315 24.510 178.405 ;
        RECT 24.970 178.325 25.645 178.485 ;
        RECT 22.380 178.125 23.120 178.155 ;
        RECT 22.380 177.825 23.295 178.125 ;
        RECT 22.970 177.650 23.295 177.825 ;
        RECT 22.000 177.095 22.255 177.625 ;
        RECT 22.425 176.915 22.730 177.375 ;
        RECT 22.975 177.295 23.295 177.650 ;
        RECT 23.465 177.865 24.005 178.235 ;
        RECT 24.340 178.145 24.745 178.315 ;
        RECT 23.465 177.465 23.705 177.865 ;
        RECT 24.185 177.695 24.405 177.975 ;
        RECT 23.875 177.525 24.405 177.695 ;
        RECT 23.875 177.295 24.045 177.525 ;
        RECT 24.575 177.365 24.745 178.145 ;
        RECT 24.915 177.535 25.265 178.155 ;
        RECT 25.435 177.535 25.645 178.325 ;
        RECT 25.835 178.355 27.335 178.525 ;
        RECT 25.835 177.665 26.005 178.355 ;
        RECT 27.695 178.185 27.865 178.965 ;
        RECT 28.670 178.835 28.840 178.965 ;
        RECT 26.175 178.015 27.865 178.185 ;
        RECT 28.035 178.405 28.500 178.795 ;
        RECT 28.670 178.665 29.065 178.835 ;
        RECT 26.175 177.835 26.345 178.015 ;
        RECT 22.975 177.125 24.045 177.295 ;
        RECT 24.215 176.915 24.405 177.355 ;
        RECT 24.575 177.085 25.525 177.365 ;
        RECT 25.835 177.275 26.095 177.665 ;
        RECT 26.515 177.595 27.305 177.845 ;
        RECT 25.745 177.105 26.095 177.275 ;
        RECT 26.305 176.915 26.635 177.375 ;
        RECT 27.510 177.305 27.680 178.015 ;
        RECT 28.035 177.815 28.205 178.405 ;
        RECT 27.850 177.595 28.205 177.815 ;
        RECT 28.375 177.595 28.725 178.215 ;
        RECT 28.895 177.305 29.065 178.665 ;
        RECT 29.430 178.495 29.755 179.280 ;
        RECT 29.235 177.445 29.695 178.495 ;
        RECT 27.510 177.135 28.365 177.305 ;
        RECT 28.570 177.135 29.065 177.305 ;
        RECT 29.235 176.915 29.565 177.275 ;
        RECT 29.925 177.175 30.095 179.295 ;
        RECT 30.265 178.965 30.595 179.465 ;
        RECT 30.765 178.795 31.020 179.295 ;
        RECT 30.270 178.625 31.020 178.795 ;
        RECT 30.270 177.635 30.500 178.625 ;
        RECT 30.670 177.805 31.020 178.455 ;
        RECT 31.660 178.325 31.995 179.295 ;
        RECT 32.165 178.325 32.335 179.465 ;
        RECT 32.505 179.125 34.535 179.295 ;
        RECT 31.660 177.655 31.830 178.325 ;
        RECT 32.505 178.155 32.675 179.125 ;
        RECT 32.000 177.825 32.255 178.155 ;
        RECT 32.480 177.825 32.675 178.155 ;
        RECT 32.845 178.785 33.970 178.955 ;
        RECT 32.085 177.655 32.255 177.825 ;
        RECT 32.845 177.655 33.015 178.785 ;
        RECT 30.270 177.465 31.020 177.635 ;
        RECT 30.265 176.915 30.595 177.295 ;
        RECT 30.765 177.175 31.020 177.465 ;
        RECT 31.660 177.085 31.915 177.655 ;
        RECT 32.085 177.485 33.015 177.655 ;
        RECT 33.185 178.445 34.195 178.615 ;
        RECT 33.185 177.645 33.355 178.445 ;
        RECT 32.840 177.450 33.015 177.485 ;
        RECT 32.085 176.915 32.415 177.315 ;
        RECT 32.840 177.085 33.370 177.450 ;
        RECT 33.560 177.425 33.835 178.245 ;
        RECT 33.555 177.255 33.835 177.425 ;
        RECT 33.560 177.085 33.835 177.255 ;
        RECT 34.005 177.085 34.195 178.445 ;
        RECT 34.365 178.460 34.535 179.125 ;
        RECT 34.705 178.705 34.875 179.465 ;
        RECT 35.110 178.705 35.625 179.115 ;
        RECT 34.365 178.270 35.115 178.460 ;
        RECT 35.285 177.895 35.625 178.705 ;
        RECT 35.795 178.300 36.085 179.465 ;
        RECT 36.255 178.375 37.465 179.465 ;
        RECT 37.840 178.495 38.170 179.295 ;
        RECT 38.340 178.665 38.670 179.465 ;
        RECT 38.970 178.495 39.300 179.295 ;
        RECT 39.945 178.665 40.195 179.465 ;
        RECT 34.395 177.725 35.625 177.895 ;
        RECT 36.255 177.835 36.775 178.375 ;
        RECT 37.840 178.325 40.275 178.495 ;
        RECT 40.465 178.325 40.635 179.465 ;
        RECT 40.805 178.325 41.145 179.295 ;
        RECT 41.520 178.495 41.850 179.295 ;
        RECT 42.020 178.665 42.350 179.465 ;
        RECT 42.650 178.495 42.980 179.295 ;
        RECT 43.625 178.665 43.875 179.465 ;
        RECT 41.520 178.325 43.955 178.495 ;
        RECT 44.145 178.325 44.315 179.465 ;
        RECT 44.485 178.325 44.825 179.295 ;
        RECT 34.375 176.915 34.885 177.450 ;
        RECT 35.105 177.120 35.350 177.725 ;
        RECT 36.945 177.665 37.465 178.205 ;
        RECT 37.635 177.905 37.985 178.155 ;
        RECT 38.170 177.695 38.340 178.325 ;
        RECT 38.510 177.905 38.840 178.105 ;
        RECT 39.010 177.905 39.340 178.105 ;
        RECT 39.510 177.905 39.930 178.105 ;
        RECT 40.105 178.075 40.275 178.325 ;
        RECT 40.105 177.905 40.800 178.075 ;
        RECT 35.795 176.915 36.085 177.640 ;
        RECT 36.255 176.915 37.465 177.665 ;
        RECT 37.840 177.085 38.340 177.695 ;
        RECT 38.970 177.565 40.195 177.735 ;
        RECT 40.970 177.715 41.145 178.325 ;
        RECT 41.315 177.905 41.665 178.155 ;
        RECT 38.970 177.085 39.300 177.565 ;
        RECT 39.470 176.915 39.695 177.375 ;
        RECT 39.865 177.085 40.195 177.565 ;
        RECT 40.385 176.915 40.635 177.715 ;
        RECT 40.805 177.085 41.145 177.715 ;
        RECT 41.850 177.695 42.020 178.325 ;
        RECT 42.190 177.905 42.520 178.105 ;
        RECT 42.690 177.905 43.020 178.105 ;
        RECT 43.190 177.905 43.610 178.105 ;
        RECT 43.785 178.075 43.955 178.325 ;
        RECT 44.595 178.275 44.825 178.325 ;
        RECT 43.785 177.905 44.480 178.075 ;
        RECT 41.520 177.085 42.020 177.695 ;
        RECT 42.650 177.565 43.875 177.735 ;
        RECT 44.650 177.715 44.825 178.275 ;
        RECT 42.650 177.085 42.980 177.565 ;
        RECT 43.150 176.915 43.375 177.375 ;
        RECT 43.545 177.085 43.875 177.565 ;
        RECT 44.065 176.915 44.315 177.715 ;
        RECT 44.485 177.085 44.825 177.715 ;
        RECT 45.000 178.325 45.335 179.295 ;
        RECT 45.505 178.325 45.675 179.465 ;
        RECT 45.845 179.125 47.875 179.295 ;
        RECT 45.000 177.655 45.170 178.325 ;
        RECT 45.845 178.155 46.015 179.125 ;
        RECT 45.340 177.825 45.595 178.155 ;
        RECT 45.820 177.825 46.015 178.155 ;
        RECT 46.185 178.785 47.310 178.955 ;
        RECT 45.425 177.655 45.595 177.825 ;
        RECT 46.185 177.655 46.355 178.785 ;
        RECT 45.000 177.085 45.255 177.655 ;
        RECT 45.425 177.485 46.355 177.655 ;
        RECT 46.525 178.445 47.535 178.615 ;
        RECT 46.525 177.645 46.695 178.445 ;
        RECT 46.180 177.450 46.355 177.485 ;
        RECT 45.425 176.915 45.755 177.315 ;
        RECT 46.180 177.085 46.710 177.450 ;
        RECT 46.900 177.425 47.175 178.245 ;
        RECT 46.895 177.255 47.175 177.425 ;
        RECT 46.900 177.085 47.175 177.255 ;
        RECT 47.345 177.085 47.535 178.445 ;
        RECT 47.705 178.460 47.875 179.125 ;
        RECT 48.045 178.705 48.215 179.465 ;
        RECT 48.450 178.705 48.965 179.115 ;
        RECT 47.705 178.270 48.455 178.460 ;
        RECT 48.625 177.895 48.965 178.705 ;
        RECT 47.735 177.725 48.965 177.895 ;
        RECT 49.135 178.705 49.650 179.115 ;
        RECT 49.885 178.705 50.055 179.465 ;
        RECT 50.225 179.125 52.255 179.295 ;
        RECT 49.135 177.895 49.475 178.705 ;
        RECT 50.225 178.460 50.395 179.125 ;
        RECT 50.790 178.785 51.915 178.955 ;
        RECT 49.645 178.270 50.395 178.460 ;
        RECT 50.565 178.445 51.575 178.615 ;
        RECT 49.135 177.725 50.365 177.895 ;
        RECT 47.715 176.915 48.225 177.450 ;
        RECT 48.445 177.120 48.690 177.725 ;
        RECT 49.410 177.120 49.655 177.725 ;
        RECT 49.875 176.915 50.385 177.450 ;
        RECT 50.565 177.085 50.755 178.445 ;
        RECT 50.925 177.425 51.200 178.245 ;
        RECT 51.405 177.645 51.575 178.445 ;
        RECT 51.745 177.655 51.915 178.785 ;
        RECT 52.085 178.155 52.255 179.125 ;
        RECT 52.425 178.325 52.595 179.465 ;
        RECT 52.765 178.325 53.100 179.295 ;
        RECT 52.085 177.825 52.280 178.155 ;
        RECT 52.505 177.825 52.760 178.155 ;
        RECT 52.505 177.655 52.675 177.825 ;
        RECT 52.930 177.655 53.100 178.325 ;
        RECT 53.275 178.705 53.790 179.115 ;
        RECT 54.025 178.705 54.195 179.465 ;
        RECT 54.365 179.125 56.395 179.295 ;
        RECT 53.275 177.895 53.615 178.705 ;
        RECT 54.365 178.460 54.535 179.125 ;
        RECT 54.930 178.785 56.055 178.955 ;
        RECT 53.785 178.270 54.535 178.460 ;
        RECT 54.705 178.445 55.715 178.615 ;
        RECT 53.275 177.725 54.505 177.895 ;
        RECT 51.745 177.485 52.675 177.655 ;
        RECT 51.745 177.450 51.920 177.485 ;
        RECT 50.925 177.255 51.205 177.425 ;
        RECT 50.925 177.085 51.200 177.255 ;
        RECT 51.390 177.085 51.920 177.450 ;
        RECT 52.345 176.915 52.675 177.315 ;
        RECT 52.845 177.085 53.100 177.655 ;
        RECT 53.550 177.120 53.795 177.725 ;
        RECT 54.015 176.915 54.525 177.450 ;
        RECT 54.705 177.085 54.895 178.445 ;
        RECT 55.065 178.105 55.340 178.245 ;
        RECT 55.065 177.935 55.345 178.105 ;
        RECT 55.065 177.085 55.340 177.935 ;
        RECT 55.545 177.645 55.715 178.445 ;
        RECT 55.885 177.655 56.055 178.785 ;
        RECT 56.225 178.155 56.395 179.125 ;
        RECT 56.565 178.325 56.735 179.465 ;
        RECT 56.905 178.325 57.240 179.295 ;
        RECT 57.470 178.595 57.755 179.465 ;
        RECT 57.925 178.835 58.185 179.295 ;
        RECT 58.360 179.005 58.615 179.465 ;
        RECT 58.785 178.835 59.045 179.295 ;
        RECT 57.925 178.665 59.045 178.835 ;
        RECT 59.215 178.665 59.525 179.465 ;
        RECT 57.925 178.415 58.185 178.665 ;
        RECT 59.695 178.495 60.005 179.295 ;
        RECT 56.225 177.825 56.420 178.155 ;
        RECT 56.645 177.825 56.900 178.155 ;
        RECT 56.645 177.655 56.815 177.825 ;
        RECT 57.070 177.655 57.240 178.325 ;
        RECT 55.885 177.485 56.815 177.655 ;
        RECT 55.885 177.450 56.060 177.485 ;
        RECT 55.530 177.085 56.060 177.450 ;
        RECT 56.485 176.915 56.815 177.315 ;
        RECT 56.985 177.085 57.240 177.655 ;
        RECT 57.430 178.245 58.185 178.415 ;
        RECT 58.975 178.325 60.005 178.495 ;
        RECT 57.430 177.735 57.835 178.245 ;
        RECT 58.975 178.075 59.145 178.325 ;
        RECT 58.005 177.905 59.145 178.075 ;
        RECT 57.430 177.565 59.080 177.735 ;
        RECT 59.315 177.585 59.665 178.155 ;
        RECT 57.475 176.915 57.755 177.395 ;
        RECT 57.925 177.175 58.185 177.565 ;
        RECT 58.360 176.915 58.615 177.395 ;
        RECT 58.785 177.175 59.080 177.565 ;
        RECT 59.835 177.415 60.005 178.325 ;
        RECT 59.260 176.915 59.535 177.395 ;
        RECT 59.705 177.085 60.005 177.415 ;
        RECT 60.175 178.390 60.445 179.295 ;
        RECT 60.615 178.705 60.945 179.465 ;
        RECT 61.125 178.535 61.295 179.295 ;
        RECT 60.175 177.590 60.345 178.390 ;
        RECT 60.630 178.365 61.295 178.535 ;
        RECT 60.630 178.220 60.800 178.365 ;
        RECT 61.555 178.300 61.845 179.465 ;
        RECT 62.020 178.315 62.280 179.465 ;
        RECT 62.455 178.390 62.710 179.295 ;
        RECT 62.880 178.705 63.210 179.465 ;
        RECT 63.425 178.535 63.595 179.295 ;
        RECT 60.515 177.890 60.800 178.220 ;
        RECT 60.630 177.635 60.800 177.890 ;
        RECT 61.035 177.815 61.365 178.185 ;
        RECT 60.175 177.085 60.435 177.590 ;
        RECT 60.630 177.465 61.295 177.635 ;
        RECT 60.615 176.915 60.945 177.295 ;
        RECT 61.125 177.085 61.295 177.465 ;
        RECT 61.555 176.915 61.845 177.640 ;
        RECT 62.020 176.915 62.280 177.755 ;
        RECT 62.455 177.660 62.625 178.390 ;
        RECT 62.880 178.365 63.595 178.535 ;
        RECT 63.945 178.535 64.115 179.295 ;
        RECT 64.330 178.705 64.660 179.465 ;
        RECT 63.945 178.365 64.660 178.535 ;
        RECT 64.830 178.390 65.085 179.295 ;
        RECT 62.880 178.155 63.050 178.365 ;
        RECT 62.795 177.825 63.050 178.155 ;
        RECT 62.455 177.085 62.710 177.660 ;
        RECT 62.880 177.635 63.050 177.825 ;
        RECT 63.330 177.815 63.685 178.185 ;
        RECT 63.855 177.815 64.210 178.185 ;
        RECT 64.490 178.155 64.660 178.365 ;
        RECT 64.490 177.825 64.745 178.155 ;
        RECT 64.490 177.635 64.660 177.825 ;
        RECT 64.915 177.660 65.085 178.390 ;
        RECT 65.260 178.315 65.520 179.465 ;
        RECT 65.705 178.405 66.035 179.465 ;
        RECT 66.215 178.155 66.385 179.080 ;
        RECT 66.555 178.875 66.885 179.275 ;
        RECT 67.055 179.105 67.385 179.465 ;
        RECT 67.585 178.875 68.285 179.295 ;
        RECT 66.555 178.645 68.285 178.875 ;
        RECT 66.555 178.425 66.885 178.645 ;
        RECT 67.080 178.155 67.405 178.445 ;
        RECT 65.695 177.825 66.005 178.155 ;
        RECT 66.215 177.825 66.590 178.155 ;
        RECT 66.910 177.825 67.405 178.155 ;
        RECT 67.580 177.905 67.910 178.445 ;
        RECT 68.080 177.765 68.285 178.645 ;
        RECT 62.880 177.465 63.595 177.635 ;
        RECT 62.880 176.915 63.210 177.295 ;
        RECT 63.425 177.085 63.595 177.465 ;
        RECT 63.945 177.465 64.660 177.635 ;
        RECT 63.945 177.085 64.115 177.465 ;
        RECT 64.330 176.915 64.660 177.295 ;
        RECT 64.830 177.085 65.085 177.660 ;
        RECT 65.260 176.915 65.520 177.755 ;
        RECT 68.055 177.675 68.285 177.765 ;
        RECT 65.705 177.445 67.065 177.655 ;
        RECT 65.705 177.085 66.035 177.445 ;
        RECT 66.205 176.915 66.535 177.275 ;
        RECT 66.735 177.085 67.065 177.445 ;
        RECT 67.575 177.085 68.285 177.675 ;
        RECT 68.915 178.495 69.225 179.295 ;
        RECT 69.395 178.665 69.705 179.465 ;
        RECT 69.875 178.835 70.135 179.295 ;
        RECT 70.305 179.005 70.560 179.465 ;
        RECT 70.735 178.835 70.995 179.295 ;
        RECT 69.875 178.665 70.995 178.835 ;
        RECT 68.915 178.325 69.945 178.495 ;
        RECT 68.915 177.415 69.085 178.325 ;
        RECT 69.255 177.585 69.605 178.155 ;
        RECT 69.775 178.075 69.945 178.325 ;
        RECT 70.735 178.415 70.995 178.665 ;
        RECT 71.165 178.595 71.450 179.465 ;
        RECT 70.735 178.245 71.490 178.415 ;
        RECT 69.775 177.905 70.915 178.075 ;
        RECT 71.085 177.735 71.490 178.245 ;
        RECT 69.840 177.565 71.490 177.735 ;
        RECT 71.675 178.325 72.015 179.295 ;
        RECT 72.185 178.325 72.355 179.465 ;
        RECT 72.625 178.665 72.875 179.465 ;
        RECT 73.520 178.495 73.850 179.295 ;
        RECT 74.150 178.665 74.480 179.465 ;
        RECT 74.650 178.495 74.980 179.295 ;
        RECT 72.545 178.325 74.980 178.495 ;
        RECT 75.415 178.325 75.625 179.465 ;
        RECT 71.675 177.715 71.850 178.325 ;
        RECT 72.545 178.075 72.715 178.325 ;
        RECT 72.020 177.905 72.715 178.075 ;
        RECT 72.890 177.905 73.310 178.105 ;
        RECT 73.480 177.905 73.810 178.105 ;
        RECT 73.980 177.905 74.310 178.105 ;
        RECT 68.915 177.085 69.215 177.415 ;
        RECT 69.385 176.915 69.660 177.395 ;
        RECT 69.840 177.175 70.135 177.565 ;
        RECT 70.305 176.915 70.560 177.395 ;
        RECT 70.735 177.175 70.995 177.565 ;
        RECT 71.165 176.915 71.445 177.395 ;
        RECT 71.675 177.085 72.015 177.715 ;
        RECT 72.185 176.915 72.435 177.715 ;
        RECT 72.625 177.565 73.850 177.735 ;
        RECT 72.625 177.085 72.955 177.565 ;
        RECT 73.125 176.915 73.350 177.375 ;
        RECT 73.520 177.085 73.850 177.565 ;
        RECT 74.480 177.695 74.650 178.325 ;
        RECT 75.795 178.315 76.125 179.295 ;
        RECT 76.295 178.325 76.525 179.465 ;
        RECT 76.735 178.705 77.250 179.115 ;
        RECT 77.485 178.705 77.655 179.465 ;
        RECT 77.825 179.125 79.855 179.295 ;
        RECT 74.835 177.905 75.185 178.155 ;
        RECT 74.480 177.085 74.980 177.695 ;
        RECT 75.415 176.915 75.625 177.735 ;
        RECT 75.795 177.715 76.045 178.315 ;
        RECT 76.215 177.905 76.545 178.155 ;
        RECT 76.735 177.895 77.075 178.705 ;
        RECT 77.825 178.460 77.995 179.125 ;
        RECT 78.390 178.785 79.515 178.955 ;
        RECT 77.245 178.270 77.995 178.460 ;
        RECT 78.165 178.445 79.175 178.615 ;
        RECT 75.795 177.085 76.125 177.715 ;
        RECT 76.295 176.915 76.525 177.735 ;
        RECT 76.735 177.725 77.965 177.895 ;
        RECT 77.010 177.120 77.255 177.725 ;
        RECT 77.475 176.915 77.985 177.450 ;
        RECT 78.165 177.085 78.355 178.445 ;
        RECT 78.525 178.105 78.800 178.245 ;
        RECT 78.525 177.935 78.805 178.105 ;
        RECT 78.525 177.085 78.800 177.935 ;
        RECT 79.005 177.645 79.175 178.445 ;
        RECT 79.345 177.655 79.515 178.785 ;
        RECT 79.685 178.155 79.855 179.125 ;
        RECT 80.025 178.325 80.195 179.465 ;
        RECT 80.365 178.325 80.700 179.295 ;
        RECT 79.685 177.825 79.880 178.155 ;
        RECT 80.105 177.825 80.360 178.155 ;
        RECT 80.105 177.655 80.275 177.825 ;
        RECT 80.530 177.655 80.700 178.325 ;
        RECT 79.345 177.485 80.275 177.655 ;
        RECT 79.345 177.450 79.520 177.485 ;
        RECT 78.990 177.085 79.520 177.450 ;
        RECT 79.945 176.915 80.275 177.315 ;
        RECT 80.445 177.085 80.700 177.655 ;
        RECT 80.875 178.325 81.260 179.295 ;
        RECT 81.430 179.005 81.755 179.465 ;
        RECT 82.275 178.835 82.555 179.295 ;
        RECT 81.430 178.615 82.555 178.835 ;
        RECT 80.875 177.655 81.155 178.325 ;
        RECT 81.430 178.155 81.880 178.615 ;
        RECT 82.745 178.445 83.145 179.295 ;
        RECT 83.545 179.005 83.815 179.465 ;
        RECT 83.985 178.835 84.270 179.295 ;
        RECT 81.325 177.825 81.880 178.155 ;
        RECT 82.050 177.885 83.145 178.445 ;
        RECT 81.430 177.715 81.880 177.825 ;
        RECT 80.875 177.085 81.260 177.655 ;
        RECT 81.430 177.545 82.555 177.715 ;
        RECT 81.430 176.915 81.755 177.375 ;
        RECT 82.275 177.085 82.555 177.545 ;
        RECT 82.745 177.085 83.145 177.885 ;
        RECT 83.315 178.615 84.270 178.835 ;
        RECT 83.315 177.715 83.525 178.615 ;
        RECT 84.565 178.485 84.895 179.295 ;
        RECT 85.065 178.665 85.305 179.465 ;
        RECT 83.695 177.885 84.385 178.445 ;
        RECT 84.565 178.315 85.280 178.485 ;
        RECT 84.560 177.905 84.940 178.145 ;
        RECT 85.110 178.075 85.280 178.315 ;
        RECT 85.485 178.445 85.655 179.295 ;
        RECT 85.825 178.665 86.155 179.465 ;
        RECT 86.325 178.445 86.495 179.295 ;
        RECT 85.485 178.275 86.495 178.445 ;
        RECT 86.665 178.315 86.995 179.465 ;
        RECT 87.315 178.300 87.605 179.465 ;
        RECT 88.695 178.325 89.035 179.295 ;
        RECT 89.205 178.325 89.375 179.465 ;
        RECT 89.645 178.665 89.895 179.465 ;
        RECT 90.540 178.495 90.870 179.295 ;
        RECT 91.170 178.665 91.500 179.465 ;
        RECT 91.670 178.495 92.000 179.295 ;
        RECT 89.565 178.325 92.000 178.495 ;
        RECT 92.435 178.325 92.645 179.465 ;
        RECT 85.110 177.905 85.610 178.075 ;
        RECT 85.110 177.735 85.280 177.905 ;
        RECT 86.000 177.765 86.495 178.275 ;
        RECT 85.995 177.735 86.495 177.765 ;
        RECT 83.315 177.545 84.270 177.715 ;
        RECT 83.545 176.915 83.815 177.375 ;
        RECT 83.985 177.085 84.270 177.545 ;
        RECT 84.645 177.565 85.280 177.735 ;
        RECT 85.485 177.565 86.495 177.735 ;
        RECT 88.695 177.715 88.870 178.325 ;
        RECT 89.565 178.075 89.735 178.325 ;
        RECT 89.040 177.905 89.735 178.075 ;
        RECT 89.905 177.935 90.330 178.105 ;
        RECT 89.910 177.905 90.330 177.935 ;
        RECT 90.500 177.905 90.830 178.105 ;
        RECT 91.000 177.905 91.330 178.105 ;
        RECT 84.645 177.085 84.815 177.565 ;
        RECT 84.995 176.915 85.235 177.395 ;
        RECT 85.485 177.085 85.655 177.565 ;
        RECT 85.825 176.915 86.155 177.395 ;
        RECT 86.325 177.085 86.495 177.565 ;
        RECT 86.665 176.915 86.995 177.715 ;
        RECT 87.315 176.915 87.605 177.640 ;
        RECT 88.695 177.085 89.035 177.715 ;
        RECT 89.205 176.915 89.455 177.715 ;
        RECT 89.645 177.565 90.870 177.735 ;
        RECT 89.645 177.085 89.975 177.565 ;
        RECT 90.145 176.915 90.370 177.375 ;
        RECT 90.540 177.085 90.870 177.565 ;
        RECT 91.500 177.695 91.670 178.325 ;
        RECT 92.815 178.315 93.145 179.295 ;
        RECT 93.315 178.325 93.545 179.465 ;
        RECT 93.755 178.325 94.095 179.295 ;
        RECT 94.265 178.325 94.435 179.465 ;
        RECT 94.705 178.665 94.955 179.465 ;
        RECT 95.600 178.495 95.930 179.295 ;
        RECT 96.230 178.665 96.560 179.465 ;
        RECT 96.730 178.495 97.060 179.295 ;
        RECT 94.625 178.325 97.060 178.495 ;
        RECT 97.435 178.375 99.105 179.465 ;
        RECT 91.855 177.905 92.205 178.155 ;
        RECT 91.500 177.085 92.000 177.695 ;
        RECT 92.435 176.915 92.645 177.735 ;
        RECT 92.815 177.715 93.065 178.315 ;
        RECT 93.235 177.905 93.565 178.155 ;
        RECT 92.815 177.085 93.145 177.715 ;
        RECT 93.315 176.915 93.545 177.735 ;
        RECT 93.755 177.715 93.930 178.325 ;
        RECT 94.625 178.075 94.795 178.325 ;
        RECT 94.100 177.905 94.795 178.075 ;
        RECT 94.970 177.905 95.390 178.105 ;
        RECT 95.560 177.905 95.890 178.105 ;
        RECT 96.060 177.905 96.390 178.105 ;
        RECT 93.755 177.085 94.095 177.715 ;
        RECT 94.265 176.915 94.515 177.715 ;
        RECT 94.705 177.565 95.930 177.735 ;
        RECT 94.705 177.085 95.035 177.565 ;
        RECT 95.205 176.915 95.430 177.375 ;
        RECT 95.600 177.085 95.930 177.565 ;
        RECT 96.560 177.695 96.730 178.325 ;
        RECT 96.915 177.905 97.265 178.155 ;
        RECT 97.435 177.855 98.185 178.375 ;
        RECT 99.275 178.325 99.660 179.295 ;
        RECT 99.830 179.005 100.155 179.465 ;
        RECT 100.675 178.835 100.955 179.295 ;
        RECT 99.830 178.615 100.955 178.835 ;
        RECT 96.560 177.085 97.060 177.695 ;
        RECT 98.355 177.685 99.105 178.205 ;
        RECT 97.435 176.915 99.105 177.685 ;
        RECT 99.275 177.655 99.555 178.325 ;
        RECT 99.830 178.155 100.280 178.615 ;
        RECT 101.145 178.445 101.545 179.295 ;
        RECT 101.945 179.005 102.215 179.465 ;
        RECT 102.385 178.835 102.670 179.295 ;
        RECT 99.725 177.825 100.280 178.155 ;
        RECT 100.450 177.885 101.545 178.445 ;
        RECT 99.830 177.715 100.280 177.825 ;
        RECT 99.275 177.085 99.660 177.655 ;
        RECT 99.830 177.545 100.955 177.715 ;
        RECT 99.830 176.915 100.155 177.375 ;
        RECT 100.675 177.085 100.955 177.545 ;
        RECT 101.145 177.085 101.545 177.885 ;
        RECT 101.715 178.615 102.670 178.835 ;
        RECT 101.715 177.715 101.925 178.615 ;
        RECT 102.095 177.885 102.785 178.445 ;
        RECT 102.955 178.325 103.295 179.295 ;
        RECT 103.465 178.325 103.635 179.465 ;
        RECT 103.905 178.665 104.155 179.465 ;
        RECT 104.800 178.495 105.130 179.295 ;
        RECT 105.430 178.665 105.760 179.465 ;
        RECT 105.930 178.495 106.260 179.295 ;
        RECT 103.825 178.325 106.260 178.495 ;
        RECT 106.635 178.390 106.905 179.295 ;
        RECT 107.075 178.705 107.405 179.465 ;
        RECT 107.585 178.535 107.755 179.295 ;
        RECT 102.955 177.765 103.130 178.325 ;
        RECT 103.825 178.075 103.995 178.325 ;
        RECT 103.300 177.905 103.995 178.075 ;
        RECT 104.170 177.905 104.590 178.105 ;
        RECT 104.760 177.905 105.090 178.105 ;
        RECT 105.260 177.905 105.590 178.105 ;
        RECT 102.955 177.715 103.185 177.765 ;
        RECT 101.715 177.545 102.670 177.715 ;
        RECT 101.945 176.915 102.215 177.375 ;
        RECT 102.385 177.085 102.670 177.545 ;
        RECT 102.955 177.085 103.295 177.715 ;
        RECT 103.465 176.915 103.715 177.715 ;
        RECT 103.905 177.565 105.130 177.735 ;
        RECT 103.905 177.085 104.235 177.565 ;
        RECT 104.405 176.915 104.630 177.375 ;
        RECT 104.800 177.085 105.130 177.565 ;
        RECT 105.760 177.695 105.930 178.325 ;
        RECT 106.115 177.905 106.465 178.155 ;
        RECT 105.760 177.085 106.260 177.695 ;
        RECT 106.635 177.590 106.805 178.390 ;
        RECT 107.090 178.365 107.755 178.535 ;
        RECT 108.105 178.535 108.275 179.295 ;
        RECT 108.455 178.705 108.785 179.465 ;
        RECT 108.105 178.365 108.770 178.535 ;
        RECT 108.955 178.390 109.225 179.295 ;
        RECT 107.090 178.220 107.260 178.365 ;
        RECT 106.975 177.890 107.260 178.220 ;
        RECT 108.600 178.220 108.770 178.365 ;
        RECT 107.090 177.635 107.260 177.890 ;
        RECT 107.495 177.815 107.825 178.185 ;
        RECT 108.035 177.815 108.365 178.185 ;
        RECT 108.600 177.890 108.885 178.220 ;
        RECT 108.600 177.635 108.770 177.890 ;
        RECT 106.635 177.085 106.895 177.590 ;
        RECT 107.090 177.465 107.755 177.635 ;
        RECT 107.075 176.915 107.405 177.295 ;
        RECT 107.585 177.085 107.755 177.465 ;
        RECT 108.105 177.465 108.770 177.635 ;
        RECT 109.055 177.590 109.225 178.390 ;
        RECT 109.395 178.375 111.985 179.465 ;
        RECT 112.155 178.375 113.365 179.465 ;
        RECT 109.395 177.855 110.605 178.375 ;
        RECT 110.775 177.685 111.985 178.205 ;
        RECT 112.155 177.835 112.675 178.375 ;
        RECT 108.105 177.085 108.275 177.465 ;
        RECT 108.455 176.915 108.785 177.295 ;
        RECT 108.965 177.085 109.225 177.590 ;
        RECT 109.395 176.915 111.985 177.685 ;
        RECT 112.845 177.665 113.365 178.205 ;
        RECT 112.155 176.915 113.365 177.665 ;
        RECT 15.010 176.745 113.450 176.915 ;
        RECT 15.095 175.995 16.305 176.745 ;
        RECT 15.095 175.455 15.615 175.995 ;
        RECT 16.475 175.975 19.065 176.745 ;
        RECT 15.785 175.285 16.305 175.825 ;
        RECT 15.095 174.195 16.305 175.285 ;
        RECT 16.475 175.285 17.685 175.805 ;
        RECT 17.855 175.455 19.065 175.975 ;
        RECT 19.350 176.115 19.635 176.575 ;
        RECT 19.805 176.285 20.075 176.745 ;
        RECT 19.350 175.945 20.305 176.115 ;
        RECT 16.475 174.195 19.065 175.285 ;
        RECT 19.235 175.215 19.925 175.775 ;
        RECT 20.095 175.045 20.305 175.945 ;
        RECT 19.350 174.825 20.305 175.045 ;
        RECT 20.475 175.775 20.875 176.575 ;
        RECT 21.065 176.115 21.345 176.575 ;
        RECT 21.865 176.285 22.190 176.745 ;
        RECT 21.065 175.945 22.190 176.115 ;
        RECT 22.360 176.005 22.745 176.575 ;
        RECT 22.915 176.020 23.205 176.745 ;
        RECT 21.740 175.835 22.190 175.945 ;
        RECT 20.475 175.215 21.570 175.775 ;
        RECT 21.740 175.505 22.295 175.835 ;
        RECT 19.350 174.365 19.635 174.825 ;
        RECT 19.805 174.195 20.075 174.655 ;
        RECT 20.475 174.365 20.875 175.215 ;
        RECT 21.740 175.045 22.190 175.505 ;
        RECT 22.465 175.335 22.745 176.005 ;
        RECT 23.375 175.975 25.045 176.745 ;
        RECT 21.065 174.825 22.190 175.045 ;
        RECT 21.065 174.365 21.345 174.825 ;
        RECT 21.865 174.195 22.190 174.655 ;
        RECT 22.360 174.365 22.745 175.335 ;
        RECT 22.915 174.195 23.205 175.360 ;
        RECT 23.375 175.285 24.125 175.805 ;
        RECT 24.295 175.455 25.045 175.975 ;
        RECT 25.255 175.925 25.485 176.745 ;
        RECT 25.655 175.945 25.985 176.575 ;
        RECT 25.235 175.505 25.565 175.755 ;
        RECT 25.735 175.345 25.985 175.945 ;
        RECT 26.155 175.925 26.365 176.745 ;
        RECT 26.600 176.035 26.855 176.565 ;
        RECT 27.025 176.285 27.330 176.745 ;
        RECT 27.575 176.365 28.645 176.535 ;
        RECT 23.375 174.195 25.045 175.285 ;
        RECT 25.255 174.195 25.485 175.335 ;
        RECT 25.655 174.365 25.985 175.345 ;
        RECT 26.600 175.385 26.810 176.035 ;
        RECT 27.575 176.010 27.895 176.365 ;
        RECT 27.570 175.835 27.895 176.010 ;
        RECT 26.980 175.535 27.895 175.835 ;
        RECT 28.065 175.795 28.305 176.195 ;
        RECT 28.475 176.135 28.645 176.365 ;
        RECT 28.815 176.305 29.005 176.745 ;
        RECT 29.175 176.295 30.125 176.575 ;
        RECT 30.345 176.385 30.695 176.555 ;
        RECT 28.475 175.965 29.005 176.135 ;
        RECT 26.980 175.505 27.720 175.535 ;
        RECT 26.155 174.195 26.365 175.335 ;
        RECT 26.600 174.505 26.855 175.385 ;
        RECT 27.025 174.195 27.330 175.335 ;
        RECT 27.550 174.915 27.720 175.505 ;
        RECT 28.065 175.425 28.605 175.795 ;
        RECT 28.785 175.685 29.005 175.965 ;
        RECT 29.175 175.515 29.345 176.295 ;
        RECT 28.940 175.345 29.345 175.515 ;
        RECT 29.515 175.505 29.865 176.125 ;
        RECT 28.940 175.255 29.110 175.345 ;
        RECT 30.035 175.335 30.245 176.125 ;
        RECT 27.890 175.085 29.110 175.255 ;
        RECT 29.570 175.175 30.245 175.335 ;
        RECT 27.550 174.745 28.350 174.915 ;
        RECT 27.670 174.195 28.000 174.575 ;
        RECT 28.180 174.455 28.350 174.745 ;
        RECT 28.940 174.705 29.110 175.085 ;
        RECT 29.280 175.165 30.245 175.175 ;
        RECT 30.435 175.995 30.695 176.385 ;
        RECT 30.905 176.285 31.235 176.745 ;
        RECT 32.110 176.355 32.965 176.525 ;
        RECT 33.170 176.355 33.665 176.525 ;
        RECT 33.835 176.385 34.165 176.745 ;
        RECT 30.435 175.305 30.605 175.995 ;
        RECT 30.775 175.645 30.945 175.825 ;
        RECT 31.115 175.815 31.905 176.065 ;
        RECT 32.110 175.645 32.280 176.355 ;
        RECT 32.450 175.845 32.805 176.065 ;
        RECT 30.775 175.475 32.465 175.645 ;
        RECT 29.280 174.875 29.740 175.165 ;
        RECT 30.435 175.135 31.935 175.305 ;
        RECT 30.435 174.995 30.605 175.135 ;
        RECT 30.045 174.825 30.605 174.995 ;
        RECT 28.520 174.195 28.770 174.655 ;
        RECT 28.940 174.365 29.810 174.705 ;
        RECT 30.045 174.365 30.215 174.825 ;
        RECT 31.050 174.795 32.125 174.965 ;
        RECT 30.385 174.195 30.755 174.655 ;
        RECT 31.050 174.455 31.220 174.795 ;
        RECT 31.390 174.195 31.720 174.625 ;
        RECT 31.955 174.455 32.125 174.795 ;
        RECT 32.295 174.695 32.465 175.475 ;
        RECT 32.635 175.255 32.805 175.845 ;
        RECT 32.975 175.445 33.325 176.065 ;
        RECT 32.635 174.865 33.100 175.255 ;
        RECT 33.495 174.995 33.665 176.355 ;
        RECT 33.835 175.165 34.295 176.215 ;
        RECT 33.270 174.825 33.665 174.995 ;
        RECT 33.270 174.695 33.440 174.825 ;
        RECT 32.295 174.365 32.975 174.695 ;
        RECT 33.190 174.365 33.440 174.695 ;
        RECT 33.610 174.195 33.860 174.655 ;
        RECT 34.030 174.380 34.355 175.165 ;
        RECT 34.525 174.365 34.695 176.485 ;
        RECT 34.865 176.365 35.195 176.745 ;
        RECT 35.365 176.195 35.620 176.485 ;
        RECT 34.870 176.025 35.620 176.195 ;
        RECT 35.795 176.070 36.055 176.575 ;
        RECT 36.235 176.365 36.565 176.745 ;
        RECT 36.745 176.195 36.915 176.575 ;
        RECT 34.870 175.035 35.100 176.025 ;
        RECT 35.270 175.205 35.620 175.855 ;
        RECT 35.795 175.270 35.965 176.070 ;
        RECT 36.250 176.025 36.915 176.195 ;
        RECT 36.250 175.770 36.420 176.025 ;
        RECT 37.840 175.965 38.340 176.575 ;
        RECT 36.135 175.440 36.420 175.770 ;
        RECT 36.655 175.475 36.985 175.845 ;
        RECT 37.635 175.505 37.985 175.755 ;
        RECT 36.250 175.295 36.420 175.440 ;
        RECT 38.170 175.335 38.340 175.965 ;
        RECT 38.970 176.095 39.300 176.575 ;
        RECT 39.470 176.285 39.695 176.745 ;
        RECT 39.865 176.095 40.195 176.575 ;
        RECT 38.970 175.925 40.195 176.095 ;
        RECT 40.385 175.945 40.635 176.745 ;
        RECT 40.805 175.945 41.145 176.575 ;
        RECT 41.430 176.115 41.715 176.575 ;
        RECT 41.885 176.285 42.155 176.745 ;
        RECT 41.430 175.945 42.385 176.115 ;
        RECT 38.510 175.555 38.840 175.755 ;
        RECT 39.010 175.555 39.340 175.755 ;
        RECT 39.510 175.555 39.930 175.755 ;
        RECT 40.105 175.585 40.800 175.755 ;
        RECT 40.105 175.335 40.275 175.585 ;
        RECT 40.970 175.335 41.145 175.945 ;
        RECT 34.870 174.865 35.620 175.035 ;
        RECT 34.865 174.195 35.195 174.695 ;
        RECT 35.365 174.365 35.620 174.865 ;
        RECT 35.795 174.365 36.065 175.270 ;
        RECT 36.250 175.125 36.915 175.295 ;
        RECT 36.235 174.195 36.565 174.955 ;
        RECT 36.745 174.365 36.915 175.125 ;
        RECT 37.840 175.165 40.275 175.335 ;
        RECT 37.840 174.365 38.170 175.165 ;
        RECT 38.340 174.195 38.670 174.995 ;
        RECT 38.970 174.365 39.300 175.165 ;
        RECT 39.945 174.195 40.195 174.995 ;
        RECT 40.465 174.195 40.635 175.335 ;
        RECT 40.805 174.365 41.145 175.335 ;
        RECT 41.315 175.215 42.005 175.775 ;
        RECT 42.175 175.045 42.385 175.945 ;
        RECT 41.430 174.825 42.385 175.045 ;
        RECT 42.555 175.775 42.955 176.575 ;
        RECT 43.145 176.115 43.425 176.575 ;
        RECT 43.945 176.285 44.270 176.745 ;
        RECT 43.145 175.945 44.270 176.115 ;
        RECT 44.440 176.005 44.825 176.575 ;
        RECT 43.820 175.835 44.270 175.945 ;
        RECT 42.555 175.215 43.650 175.775 ;
        RECT 43.820 175.505 44.375 175.835 ;
        RECT 41.430 174.365 41.715 174.825 ;
        RECT 41.885 174.195 42.155 174.655 ;
        RECT 42.555 174.365 42.955 175.215 ;
        RECT 43.820 175.045 44.270 175.505 ;
        RECT 44.545 175.335 44.825 176.005 ;
        RECT 43.145 174.825 44.270 175.045 ;
        RECT 43.145 174.365 43.425 174.825 ;
        RECT 43.945 174.195 44.270 174.655 ;
        RECT 44.440 174.365 44.825 175.335 ;
        RECT 44.995 175.945 45.335 176.575 ;
        RECT 45.505 175.945 45.755 176.745 ;
        RECT 45.945 176.095 46.275 176.575 ;
        RECT 46.445 176.285 46.670 176.745 ;
        RECT 46.840 176.095 47.170 176.575 ;
        RECT 44.995 175.335 45.170 175.945 ;
        RECT 45.945 175.925 47.170 176.095 ;
        RECT 47.800 175.965 48.300 176.575 ;
        RECT 48.675 176.020 48.965 176.745 ;
        RECT 49.140 176.035 49.395 176.565 ;
        RECT 49.565 176.285 49.870 176.745 ;
        RECT 50.115 176.365 51.185 176.535 ;
        RECT 45.340 175.585 46.035 175.755 ;
        RECT 45.865 175.335 46.035 175.585 ;
        RECT 46.210 175.555 46.630 175.755 ;
        RECT 46.800 175.555 47.130 175.755 ;
        RECT 47.300 175.555 47.630 175.755 ;
        RECT 47.800 175.335 47.970 175.965 ;
        RECT 48.155 175.505 48.505 175.755 ;
        RECT 49.140 175.385 49.350 176.035 ;
        RECT 50.115 176.010 50.435 176.365 ;
        RECT 50.110 175.835 50.435 176.010 ;
        RECT 49.520 175.535 50.435 175.835 ;
        RECT 50.605 175.795 50.845 176.195 ;
        RECT 51.015 176.135 51.185 176.365 ;
        RECT 51.355 176.305 51.545 176.745 ;
        RECT 51.715 176.295 52.665 176.575 ;
        RECT 52.885 176.385 53.235 176.555 ;
        RECT 51.015 175.965 51.545 176.135 ;
        RECT 49.520 175.505 50.260 175.535 ;
        RECT 44.995 174.365 45.335 175.335 ;
        RECT 45.505 174.195 45.675 175.335 ;
        RECT 45.865 175.165 48.300 175.335 ;
        RECT 45.945 174.195 46.195 174.995 ;
        RECT 46.840 174.365 47.170 175.165 ;
        RECT 47.470 174.195 47.800 174.995 ;
        RECT 47.970 174.365 48.300 175.165 ;
        RECT 48.675 174.195 48.965 175.360 ;
        RECT 49.140 174.505 49.395 175.385 ;
        RECT 49.565 174.195 49.870 175.335 ;
        RECT 50.090 174.915 50.260 175.505 ;
        RECT 50.605 175.425 51.145 175.795 ;
        RECT 51.325 175.685 51.545 175.965 ;
        RECT 51.715 175.515 51.885 176.295 ;
        RECT 51.480 175.345 51.885 175.515 ;
        RECT 52.055 175.505 52.405 176.125 ;
        RECT 51.480 175.255 51.650 175.345 ;
        RECT 52.575 175.335 52.785 176.125 ;
        RECT 50.430 175.085 51.650 175.255 ;
        RECT 52.110 175.175 52.785 175.335 ;
        RECT 50.090 174.745 50.890 174.915 ;
        RECT 50.210 174.195 50.540 174.575 ;
        RECT 50.720 174.455 50.890 174.745 ;
        RECT 51.480 174.705 51.650 175.085 ;
        RECT 51.820 175.165 52.785 175.175 ;
        RECT 52.975 175.995 53.235 176.385 ;
        RECT 53.445 176.285 53.775 176.745 ;
        RECT 54.650 176.355 55.505 176.525 ;
        RECT 55.710 176.355 56.205 176.525 ;
        RECT 56.375 176.385 56.705 176.745 ;
        RECT 52.975 175.305 53.145 175.995 ;
        RECT 53.315 175.645 53.485 175.825 ;
        RECT 53.655 175.815 54.445 176.065 ;
        RECT 54.650 175.645 54.820 176.355 ;
        RECT 54.990 175.845 55.345 176.065 ;
        RECT 53.315 175.475 55.005 175.645 ;
        RECT 51.820 174.875 52.280 175.165 ;
        RECT 52.975 175.135 54.475 175.305 ;
        RECT 52.975 174.995 53.145 175.135 ;
        RECT 52.585 174.825 53.145 174.995 ;
        RECT 51.060 174.195 51.310 174.655 ;
        RECT 51.480 174.365 52.350 174.705 ;
        RECT 52.585 174.365 52.755 174.825 ;
        RECT 53.590 174.795 54.665 174.965 ;
        RECT 52.925 174.195 53.295 174.655 ;
        RECT 53.590 174.455 53.760 174.795 ;
        RECT 53.930 174.195 54.260 174.625 ;
        RECT 54.495 174.455 54.665 174.795 ;
        RECT 54.835 174.695 55.005 175.475 ;
        RECT 55.175 175.255 55.345 175.845 ;
        RECT 55.515 175.445 55.865 176.065 ;
        RECT 55.175 174.865 55.640 175.255 ;
        RECT 56.035 174.995 56.205 176.355 ;
        RECT 56.375 175.165 56.835 176.215 ;
        RECT 55.810 174.825 56.205 174.995 ;
        RECT 55.810 174.695 55.980 174.825 ;
        RECT 54.835 174.365 55.515 174.695 ;
        RECT 55.730 174.365 55.980 174.695 ;
        RECT 56.150 174.195 56.400 174.655 ;
        RECT 56.570 174.380 56.895 175.165 ;
        RECT 57.065 174.365 57.235 176.485 ;
        RECT 57.405 176.365 57.735 176.745 ;
        RECT 57.905 176.195 58.160 176.485 ;
        RECT 57.410 176.025 58.160 176.195 ;
        RECT 58.450 176.115 58.735 176.575 ;
        RECT 58.905 176.285 59.175 176.745 ;
        RECT 57.410 175.035 57.640 176.025 ;
        RECT 58.450 175.945 59.405 176.115 ;
        RECT 57.810 175.205 58.160 175.855 ;
        RECT 58.335 175.215 59.025 175.775 ;
        RECT 59.195 175.045 59.405 175.945 ;
        RECT 57.410 174.865 58.160 175.035 ;
        RECT 57.405 174.195 57.735 174.695 ;
        RECT 57.905 174.365 58.160 174.865 ;
        RECT 58.450 174.825 59.405 175.045 ;
        RECT 59.575 175.775 59.975 176.575 ;
        RECT 60.165 176.115 60.445 176.575 ;
        RECT 60.965 176.285 61.290 176.745 ;
        RECT 60.165 175.945 61.290 176.115 ;
        RECT 61.460 176.005 61.845 176.575 ;
        RECT 62.565 176.195 62.735 176.575 ;
        RECT 62.950 176.365 63.280 176.745 ;
        RECT 62.565 176.025 63.280 176.195 ;
        RECT 60.840 175.835 61.290 175.945 ;
        RECT 59.575 175.215 60.670 175.775 ;
        RECT 60.840 175.505 61.395 175.835 ;
        RECT 58.450 174.365 58.735 174.825 ;
        RECT 58.905 174.195 59.175 174.655 ;
        RECT 59.575 174.365 59.975 175.215 ;
        RECT 60.840 175.045 61.290 175.505 ;
        RECT 61.565 175.335 61.845 176.005 ;
        RECT 62.475 175.475 62.830 175.845 ;
        RECT 63.110 175.835 63.280 176.025 ;
        RECT 63.450 176.000 63.705 176.575 ;
        RECT 63.110 175.505 63.365 175.835 ;
        RECT 60.165 174.825 61.290 175.045 ;
        RECT 60.165 174.365 60.445 174.825 ;
        RECT 60.965 174.195 61.290 174.655 ;
        RECT 61.460 174.365 61.845 175.335 ;
        RECT 63.110 175.295 63.280 175.505 ;
        RECT 62.565 175.125 63.280 175.295 ;
        RECT 63.535 175.270 63.705 176.000 ;
        RECT 63.880 175.905 64.140 176.745 ;
        RECT 64.320 175.905 64.580 176.745 ;
        RECT 64.755 176.000 65.010 176.575 ;
        RECT 65.180 176.365 65.510 176.745 ;
        RECT 65.725 176.195 65.895 176.575 ;
        RECT 65.180 176.025 65.895 176.195 ;
        RECT 62.565 174.365 62.735 175.125 ;
        RECT 62.950 174.195 63.280 174.955 ;
        RECT 63.450 174.365 63.705 175.270 ;
        RECT 63.880 174.195 64.140 175.345 ;
        RECT 64.320 174.195 64.580 175.345 ;
        RECT 64.755 175.270 64.925 176.000 ;
        RECT 65.180 175.835 65.350 176.025 ;
        RECT 67.075 175.945 67.415 176.575 ;
        RECT 67.585 175.945 67.835 176.745 ;
        RECT 68.025 176.095 68.355 176.575 ;
        RECT 68.525 176.285 68.750 176.745 ;
        RECT 68.920 176.095 69.250 176.575 ;
        RECT 65.095 175.505 65.350 175.835 ;
        RECT 65.180 175.295 65.350 175.505 ;
        RECT 65.630 175.475 65.985 175.845 ;
        RECT 67.075 175.335 67.250 175.945 ;
        RECT 68.025 175.925 69.250 176.095 ;
        RECT 69.880 175.965 70.380 176.575 ;
        RECT 67.420 175.585 68.115 175.755 ;
        RECT 67.945 175.335 68.115 175.585 ;
        RECT 68.290 175.555 68.710 175.755 ;
        RECT 68.880 175.555 69.210 175.755 ;
        RECT 69.380 175.555 69.710 175.755 ;
        RECT 69.880 175.335 70.050 175.965 ;
        RECT 70.755 175.945 71.095 176.575 ;
        RECT 71.265 175.945 71.515 176.745 ;
        RECT 71.705 176.095 72.035 176.575 ;
        RECT 72.205 176.285 72.430 176.745 ;
        RECT 72.600 176.095 72.930 176.575 ;
        RECT 70.235 175.505 70.585 175.755 ;
        RECT 70.755 175.335 70.930 175.945 ;
        RECT 71.705 175.925 72.930 176.095 ;
        RECT 73.560 175.965 74.060 176.575 ;
        RECT 74.435 176.020 74.725 176.745 ;
        RECT 71.100 175.585 71.795 175.755 ;
        RECT 71.625 175.335 71.795 175.585 ;
        RECT 71.970 175.555 72.390 175.755 ;
        RECT 72.560 175.555 72.890 175.755 ;
        RECT 73.060 175.555 73.390 175.755 ;
        RECT 73.560 175.335 73.730 175.965 ;
        RECT 74.895 175.945 75.235 176.575 ;
        RECT 75.405 175.945 75.655 176.745 ;
        RECT 75.845 176.095 76.175 176.575 ;
        RECT 76.345 176.285 76.570 176.745 ;
        RECT 76.740 176.095 77.070 176.575 ;
        RECT 73.915 175.505 74.265 175.755 ;
        RECT 64.755 174.365 65.010 175.270 ;
        RECT 65.180 175.125 65.895 175.295 ;
        RECT 65.180 174.195 65.510 174.955 ;
        RECT 65.725 174.365 65.895 175.125 ;
        RECT 67.075 174.365 67.415 175.335 ;
        RECT 67.585 174.195 67.755 175.335 ;
        RECT 67.945 175.165 70.380 175.335 ;
        RECT 68.025 174.195 68.275 174.995 ;
        RECT 68.920 174.365 69.250 175.165 ;
        RECT 69.550 174.195 69.880 174.995 ;
        RECT 70.050 174.365 70.380 175.165 ;
        RECT 70.755 174.365 71.095 175.335 ;
        RECT 71.265 174.195 71.435 175.335 ;
        RECT 71.625 175.165 74.060 175.335 ;
        RECT 71.705 174.195 71.955 174.995 ;
        RECT 72.600 174.365 72.930 175.165 ;
        RECT 73.230 174.195 73.560 174.995 ;
        RECT 73.730 174.365 74.060 175.165 ;
        RECT 74.435 174.195 74.725 175.360 ;
        RECT 74.895 175.335 75.070 175.945 ;
        RECT 75.845 175.925 77.070 176.095 ;
        RECT 77.700 175.965 78.200 176.575 ;
        RECT 78.690 176.115 78.975 176.575 ;
        RECT 79.145 176.285 79.415 176.745 ;
        RECT 75.240 175.585 75.935 175.755 ;
        RECT 75.765 175.335 75.935 175.585 ;
        RECT 76.110 175.555 76.530 175.755 ;
        RECT 76.700 175.555 77.030 175.755 ;
        RECT 77.200 175.555 77.530 175.755 ;
        RECT 77.700 175.335 77.870 175.965 ;
        RECT 78.690 175.945 79.645 176.115 ;
        RECT 78.055 175.505 78.405 175.755 ;
        RECT 74.895 174.365 75.235 175.335 ;
        RECT 75.405 174.195 75.575 175.335 ;
        RECT 75.765 175.165 78.200 175.335 ;
        RECT 78.575 175.215 79.265 175.775 ;
        RECT 75.845 174.195 76.095 174.995 ;
        RECT 76.740 174.365 77.070 175.165 ;
        RECT 77.370 174.195 77.700 174.995 ;
        RECT 77.870 174.365 78.200 175.165 ;
        RECT 79.435 175.045 79.645 175.945 ;
        RECT 78.690 174.825 79.645 175.045 ;
        RECT 79.815 175.775 80.215 176.575 ;
        RECT 80.405 176.115 80.685 176.575 ;
        RECT 81.205 176.285 81.530 176.745 ;
        RECT 80.405 175.945 81.530 176.115 ;
        RECT 81.700 176.005 82.085 176.575 ;
        RECT 82.260 176.195 82.515 176.485 ;
        RECT 82.685 176.365 83.015 176.745 ;
        RECT 82.260 176.025 83.010 176.195 ;
        RECT 81.080 175.835 81.530 175.945 ;
        RECT 79.815 175.215 80.910 175.775 ;
        RECT 81.080 175.505 81.635 175.835 ;
        RECT 78.690 174.365 78.975 174.825 ;
        RECT 79.145 174.195 79.415 174.655 ;
        RECT 79.815 174.365 80.215 175.215 ;
        RECT 81.080 175.045 81.530 175.505 ;
        RECT 81.805 175.335 82.085 176.005 ;
        RECT 80.405 174.825 81.530 175.045 ;
        RECT 80.405 174.365 80.685 174.825 ;
        RECT 81.205 174.195 81.530 174.655 ;
        RECT 81.700 174.365 82.085 175.335 ;
        RECT 82.260 175.205 82.610 175.855 ;
        RECT 82.780 175.035 83.010 176.025 ;
        RECT 82.260 174.865 83.010 175.035 ;
        RECT 82.260 174.365 82.515 174.865 ;
        RECT 82.685 174.195 83.015 174.695 ;
        RECT 83.185 174.365 83.355 176.485 ;
        RECT 83.715 176.385 84.045 176.745 ;
        RECT 84.215 176.355 84.710 176.525 ;
        RECT 84.915 176.355 85.770 176.525 ;
        RECT 83.585 175.165 84.045 176.215 ;
        RECT 83.525 174.380 83.850 175.165 ;
        RECT 84.215 174.995 84.385 176.355 ;
        RECT 84.555 175.445 84.905 176.065 ;
        RECT 85.075 175.845 85.430 176.065 ;
        RECT 85.075 175.255 85.245 175.845 ;
        RECT 85.600 175.645 85.770 176.355 ;
        RECT 86.645 176.285 86.975 176.745 ;
        RECT 87.185 176.385 87.535 176.555 ;
        RECT 85.975 175.815 86.765 176.065 ;
        RECT 87.185 175.995 87.445 176.385 ;
        RECT 87.755 176.295 88.705 176.575 ;
        RECT 88.875 176.305 89.065 176.745 ;
        RECT 89.235 176.365 90.305 176.535 ;
        RECT 86.935 175.645 87.105 175.825 ;
        RECT 84.215 174.825 84.610 174.995 ;
        RECT 84.780 174.865 85.245 175.255 ;
        RECT 85.415 175.475 87.105 175.645 ;
        RECT 84.440 174.695 84.610 174.825 ;
        RECT 85.415 174.695 85.585 175.475 ;
        RECT 87.275 175.305 87.445 175.995 ;
        RECT 85.945 175.135 87.445 175.305 ;
        RECT 87.635 175.335 87.845 176.125 ;
        RECT 88.015 175.505 88.365 176.125 ;
        RECT 88.535 175.515 88.705 176.295 ;
        RECT 89.235 176.135 89.405 176.365 ;
        RECT 88.875 175.965 89.405 176.135 ;
        RECT 88.875 175.685 89.095 175.965 ;
        RECT 89.575 175.795 89.815 176.195 ;
        RECT 88.535 175.345 88.940 175.515 ;
        RECT 89.275 175.425 89.815 175.795 ;
        RECT 89.985 176.010 90.305 176.365 ;
        RECT 90.550 176.285 90.855 176.745 ;
        RECT 91.025 176.035 91.280 176.565 ;
        RECT 89.985 175.835 90.310 176.010 ;
        RECT 89.985 175.535 90.900 175.835 ;
        RECT 90.160 175.505 90.900 175.535 ;
        RECT 87.635 175.175 88.310 175.335 ;
        RECT 88.770 175.255 88.940 175.345 ;
        RECT 87.635 175.165 88.600 175.175 ;
        RECT 87.275 174.995 87.445 175.135 ;
        RECT 84.020 174.195 84.270 174.655 ;
        RECT 84.440 174.365 84.690 174.695 ;
        RECT 84.905 174.365 85.585 174.695 ;
        RECT 85.755 174.795 86.830 174.965 ;
        RECT 87.275 174.825 87.835 174.995 ;
        RECT 88.140 174.875 88.600 175.165 ;
        RECT 88.770 175.085 89.990 175.255 ;
        RECT 85.755 174.455 85.925 174.795 ;
        RECT 86.160 174.195 86.490 174.625 ;
        RECT 86.660 174.455 86.830 174.795 ;
        RECT 87.125 174.195 87.495 174.655 ;
        RECT 87.665 174.365 87.835 174.825 ;
        RECT 88.770 174.705 88.940 175.085 ;
        RECT 90.160 174.915 90.330 175.505 ;
        RECT 91.070 175.385 91.280 176.035 ;
        RECT 88.070 174.365 88.940 174.705 ;
        RECT 89.530 174.745 90.330 174.915 ;
        RECT 89.110 174.195 89.360 174.655 ;
        RECT 89.530 174.455 89.700 174.745 ;
        RECT 89.880 174.195 90.210 174.575 ;
        RECT 90.550 174.195 90.855 175.335 ;
        RECT 91.025 174.505 91.280 175.385 ;
        RECT 91.455 176.070 91.715 176.575 ;
        RECT 91.895 176.365 92.225 176.745 ;
        RECT 92.405 176.195 92.575 176.575 ;
        RECT 91.455 175.270 91.625 176.070 ;
        RECT 91.910 176.025 92.575 176.195 ;
        RECT 91.910 175.770 92.080 176.025 ;
        RECT 93.755 175.945 94.095 176.575 ;
        RECT 94.265 175.945 94.515 176.745 ;
        RECT 94.705 176.095 95.035 176.575 ;
        RECT 95.205 176.285 95.430 176.745 ;
        RECT 95.600 176.095 95.930 176.575 ;
        RECT 91.795 175.440 92.080 175.770 ;
        RECT 92.315 175.475 92.645 175.845 ;
        RECT 91.910 175.295 92.080 175.440 ;
        RECT 93.755 175.335 93.930 175.945 ;
        RECT 94.705 175.925 95.930 176.095 ;
        RECT 96.560 175.965 97.060 176.575 ;
        RECT 97.435 175.975 100.025 176.745 ;
        RECT 100.195 176.020 100.485 176.745 ;
        RECT 100.655 175.975 102.325 176.745 ;
        RECT 94.100 175.585 94.795 175.755 ;
        RECT 94.625 175.335 94.795 175.585 ;
        RECT 94.970 175.555 95.390 175.755 ;
        RECT 95.560 175.555 95.890 175.755 ;
        RECT 96.060 175.555 96.390 175.755 ;
        RECT 96.560 175.335 96.730 175.965 ;
        RECT 96.915 175.505 97.265 175.755 ;
        RECT 91.455 174.365 91.725 175.270 ;
        RECT 91.910 175.125 92.575 175.295 ;
        RECT 91.895 174.195 92.225 174.955 ;
        RECT 92.405 174.365 92.575 175.125 ;
        RECT 93.755 174.365 94.095 175.335 ;
        RECT 94.265 174.195 94.435 175.335 ;
        RECT 94.625 175.165 97.060 175.335 ;
        RECT 94.705 174.195 94.955 174.995 ;
        RECT 95.600 174.365 95.930 175.165 ;
        RECT 96.230 174.195 96.560 174.995 ;
        RECT 96.730 174.365 97.060 175.165 ;
        RECT 97.435 175.285 98.645 175.805 ;
        RECT 98.815 175.455 100.025 175.975 ;
        RECT 97.435 174.195 100.025 175.285 ;
        RECT 100.195 174.195 100.485 175.360 ;
        RECT 100.655 175.285 101.405 175.805 ;
        RECT 101.575 175.455 102.325 175.975 ;
        RECT 102.500 176.035 102.755 176.565 ;
        RECT 102.925 176.285 103.230 176.745 ;
        RECT 103.475 176.365 104.545 176.535 ;
        RECT 102.500 175.385 102.710 176.035 ;
        RECT 103.475 176.010 103.795 176.365 ;
        RECT 103.470 175.835 103.795 176.010 ;
        RECT 102.880 175.535 103.795 175.835 ;
        RECT 103.965 175.795 104.205 176.195 ;
        RECT 104.375 176.135 104.545 176.365 ;
        RECT 104.715 176.305 104.905 176.745 ;
        RECT 105.075 176.295 106.025 176.575 ;
        RECT 106.245 176.385 106.595 176.555 ;
        RECT 104.375 175.965 104.905 176.135 ;
        RECT 102.880 175.505 103.620 175.535 ;
        RECT 100.655 174.195 102.325 175.285 ;
        RECT 102.500 174.505 102.755 175.385 ;
        RECT 102.925 174.195 103.230 175.335 ;
        RECT 103.450 174.915 103.620 175.505 ;
        RECT 103.965 175.425 104.505 175.795 ;
        RECT 104.685 175.685 104.905 175.965 ;
        RECT 105.075 175.515 105.245 176.295 ;
        RECT 104.840 175.345 105.245 175.515 ;
        RECT 105.415 175.505 105.765 176.125 ;
        RECT 104.840 175.255 105.010 175.345 ;
        RECT 105.935 175.335 106.145 176.125 ;
        RECT 103.790 175.085 105.010 175.255 ;
        RECT 105.470 175.175 106.145 175.335 ;
        RECT 103.450 174.745 104.250 174.915 ;
        RECT 103.570 174.195 103.900 174.575 ;
        RECT 104.080 174.455 104.250 174.745 ;
        RECT 104.840 174.705 105.010 175.085 ;
        RECT 105.180 175.165 106.145 175.175 ;
        RECT 106.335 175.995 106.595 176.385 ;
        RECT 106.805 176.285 107.135 176.745 ;
        RECT 108.010 176.355 108.865 176.525 ;
        RECT 109.070 176.355 109.565 176.525 ;
        RECT 109.735 176.385 110.065 176.745 ;
        RECT 106.335 175.305 106.505 175.995 ;
        RECT 106.675 175.645 106.845 175.825 ;
        RECT 107.015 175.815 107.805 176.065 ;
        RECT 108.010 175.645 108.180 176.355 ;
        RECT 108.350 175.845 108.705 176.065 ;
        RECT 106.675 175.475 108.365 175.645 ;
        RECT 105.180 174.875 105.640 175.165 ;
        RECT 106.335 175.135 107.835 175.305 ;
        RECT 106.335 174.995 106.505 175.135 ;
        RECT 105.945 174.825 106.505 174.995 ;
        RECT 104.420 174.195 104.670 174.655 ;
        RECT 104.840 174.365 105.710 174.705 ;
        RECT 105.945 174.365 106.115 174.825 ;
        RECT 106.950 174.795 108.025 174.965 ;
        RECT 106.285 174.195 106.655 174.655 ;
        RECT 106.950 174.455 107.120 174.795 ;
        RECT 107.290 174.195 107.620 174.625 ;
        RECT 107.855 174.455 108.025 174.795 ;
        RECT 108.195 174.695 108.365 175.475 ;
        RECT 108.535 175.255 108.705 175.845 ;
        RECT 108.875 175.445 109.225 176.065 ;
        RECT 108.535 174.865 109.000 175.255 ;
        RECT 109.395 174.995 109.565 176.355 ;
        RECT 109.735 175.165 110.195 176.215 ;
        RECT 109.170 174.825 109.565 174.995 ;
        RECT 109.170 174.695 109.340 174.825 ;
        RECT 108.195 174.365 108.875 174.695 ;
        RECT 109.090 174.365 109.340 174.695 ;
        RECT 109.510 174.195 109.760 174.655 ;
        RECT 109.930 174.380 110.255 175.165 ;
        RECT 110.425 174.365 110.595 176.485 ;
        RECT 110.765 176.365 111.095 176.745 ;
        RECT 111.265 176.195 111.520 176.485 ;
        RECT 110.770 176.025 111.520 176.195 ;
        RECT 110.770 175.035 111.000 176.025 ;
        RECT 112.155 175.995 113.365 176.745 ;
        RECT 111.170 175.205 111.520 175.855 ;
        RECT 112.155 175.285 112.675 175.825 ;
        RECT 112.845 175.455 113.365 175.995 ;
        RECT 110.770 174.865 111.520 175.035 ;
        RECT 110.765 174.195 111.095 174.695 ;
        RECT 111.265 174.365 111.520 174.865 ;
        RECT 112.155 174.195 113.365 175.285 ;
        RECT 15.010 174.025 113.450 174.195 ;
        RECT 15.095 172.935 16.305 174.025 ;
        RECT 16.590 173.395 16.875 173.855 ;
        RECT 17.045 173.565 17.315 174.025 ;
        RECT 16.590 173.175 17.545 173.395 ;
        RECT 15.095 172.225 15.615 172.765 ;
        RECT 15.785 172.395 16.305 172.935 ;
        RECT 16.475 172.445 17.165 173.005 ;
        RECT 17.335 172.275 17.545 173.175 ;
        RECT 15.095 171.475 16.305 172.225 ;
        RECT 16.590 172.105 17.545 172.275 ;
        RECT 17.715 173.005 18.115 173.855 ;
        RECT 18.305 173.395 18.585 173.855 ;
        RECT 19.105 173.565 19.430 174.025 ;
        RECT 18.305 173.175 19.430 173.395 ;
        RECT 17.715 172.445 18.810 173.005 ;
        RECT 18.980 172.715 19.430 173.175 ;
        RECT 19.600 172.885 19.985 173.855 ;
        RECT 16.590 171.645 16.875 172.105 ;
        RECT 17.045 171.475 17.315 171.935 ;
        RECT 17.715 171.645 18.115 172.445 ;
        RECT 18.980 172.385 19.535 172.715 ;
        RECT 18.980 172.275 19.430 172.385 ;
        RECT 18.305 172.105 19.430 172.275 ;
        RECT 19.705 172.215 19.985 172.885 ;
        RECT 18.305 171.645 18.585 172.105 ;
        RECT 19.105 171.475 19.430 171.935 ;
        RECT 19.600 171.645 19.985 172.215 ;
        RECT 20.160 172.835 20.415 173.715 ;
        RECT 20.585 172.885 20.890 174.025 ;
        RECT 21.230 173.645 21.560 174.025 ;
        RECT 21.740 173.475 21.910 173.765 ;
        RECT 22.080 173.565 22.330 174.025 ;
        RECT 21.110 173.305 21.910 173.475 ;
        RECT 22.500 173.515 23.370 173.855 ;
        RECT 20.160 172.185 20.370 172.835 ;
        RECT 21.110 172.715 21.280 173.305 ;
        RECT 22.500 173.135 22.670 173.515 ;
        RECT 23.605 173.395 23.775 173.855 ;
        RECT 23.945 173.565 24.315 174.025 ;
        RECT 24.610 173.425 24.780 173.765 ;
        RECT 24.950 173.595 25.280 174.025 ;
        RECT 25.515 173.425 25.685 173.765 ;
        RECT 21.450 172.965 22.670 173.135 ;
        RECT 22.840 173.055 23.300 173.345 ;
        RECT 23.605 173.225 24.165 173.395 ;
        RECT 24.610 173.255 25.685 173.425 ;
        RECT 25.855 173.525 26.535 173.855 ;
        RECT 26.750 173.525 27.000 173.855 ;
        RECT 27.170 173.565 27.420 174.025 ;
        RECT 23.995 173.085 24.165 173.225 ;
        RECT 22.840 173.045 23.805 173.055 ;
        RECT 22.500 172.875 22.670 172.965 ;
        RECT 23.130 172.885 23.805 173.045 ;
        RECT 20.540 172.685 21.280 172.715 ;
        RECT 20.540 172.385 21.455 172.685 ;
        RECT 21.130 172.210 21.455 172.385 ;
        RECT 20.160 171.655 20.415 172.185 ;
        RECT 20.585 171.475 20.890 171.935 ;
        RECT 21.135 171.855 21.455 172.210 ;
        RECT 21.625 172.425 22.165 172.795 ;
        RECT 22.500 172.705 22.905 172.875 ;
        RECT 21.625 172.025 21.865 172.425 ;
        RECT 22.345 172.255 22.565 172.535 ;
        RECT 22.035 172.085 22.565 172.255 ;
        RECT 22.035 171.855 22.205 172.085 ;
        RECT 22.735 171.925 22.905 172.705 ;
        RECT 23.075 172.095 23.425 172.715 ;
        RECT 23.595 172.095 23.805 172.885 ;
        RECT 23.995 172.915 25.495 173.085 ;
        RECT 23.995 172.225 24.165 172.915 ;
        RECT 25.855 172.745 26.025 173.525 ;
        RECT 26.830 173.395 27.000 173.525 ;
        RECT 24.335 172.575 26.025 172.745 ;
        RECT 26.195 172.965 26.660 173.355 ;
        RECT 26.830 173.225 27.225 173.395 ;
        RECT 24.335 172.395 24.505 172.575 ;
        RECT 21.135 171.685 22.205 171.855 ;
        RECT 22.375 171.475 22.565 171.915 ;
        RECT 22.735 171.645 23.685 171.925 ;
        RECT 23.995 171.835 24.255 172.225 ;
        RECT 24.675 172.155 25.465 172.405 ;
        RECT 23.905 171.665 24.255 171.835 ;
        RECT 24.465 171.475 24.795 171.935 ;
        RECT 25.670 171.865 25.840 172.575 ;
        RECT 26.195 172.375 26.365 172.965 ;
        RECT 26.010 172.155 26.365 172.375 ;
        RECT 26.535 172.155 26.885 172.775 ;
        RECT 27.055 171.865 27.225 173.225 ;
        RECT 27.590 173.055 27.915 173.840 ;
        RECT 27.395 172.005 27.855 173.055 ;
        RECT 25.670 171.695 26.525 171.865 ;
        RECT 26.730 171.695 27.225 171.865 ;
        RECT 27.395 171.475 27.725 171.835 ;
        RECT 28.085 171.735 28.255 173.855 ;
        RECT 28.425 173.525 28.755 174.025 ;
        RECT 28.925 173.355 29.180 173.855 ;
        RECT 28.430 173.185 29.180 173.355 ;
        RECT 28.430 172.195 28.660 173.185 ;
        RECT 28.830 172.365 29.180 173.015 ;
        RECT 29.360 172.885 29.695 173.855 ;
        RECT 29.865 172.885 30.035 174.025 ;
        RECT 30.205 173.685 32.235 173.855 ;
        RECT 29.360 172.215 29.530 172.885 ;
        RECT 30.205 172.715 30.375 173.685 ;
        RECT 29.700 172.385 29.955 172.715 ;
        RECT 30.180 172.385 30.375 172.715 ;
        RECT 30.545 173.345 31.670 173.515 ;
        RECT 29.785 172.215 29.955 172.385 ;
        RECT 30.545 172.215 30.715 173.345 ;
        RECT 28.430 172.025 29.180 172.195 ;
        RECT 28.425 171.475 28.755 171.855 ;
        RECT 28.925 171.735 29.180 172.025 ;
        RECT 29.360 171.645 29.615 172.215 ;
        RECT 29.785 172.045 30.715 172.215 ;
        RECT 30.885 173.005 31.895 173.175 ;
        RECT 30.885 172.205 31.055 173.005 ;
        RECT 30.540 172.010 30.715 172.045 ;
        RECT 29.785 171.475 30.115 171.875 ;
        RECT 30.540 171.645 31.070 172.010 ;
        RECT 31.260 171.985 31.535 172.805 ;
        RECT 31.255 171.815 31.535 171.985 ;
        RECT 31.260 171.645 31.535 171.815 ;
        RECT 31.705 171.645 31.895 173.005 ;
        RECT 32.065 173.020 32.235 173.685 ;
        RECT 32.405 173.265 32.575 174.025 ;
        RECT 32.810 173.265 33.325 173.675 ;
        RECT 32.065 172.830 32.815 173.020 ;
        RECT 32.985 172.455 33.325 173.265 ;
        RECT 32.095 172.285 33.325 172.455 ;
        RECT 33.955 172.935 35.625 174.025 ;
        RECT 33.955 172.415 34.705 172.935 ;
        RECT 35.795 172.860 36.085 174.025 ;
        RECT 36.315 172.885 36.525 174.025 ;
        RECT 36.695 172.875 37.025 173.855 ;
        RECT 37.195 172.885 37.425 174.025 ;
        RECT 37.635 172.885 37.975 173.855 ;
        RECT 38.145 172.885 38.315 174.025 ;
        RECT 38.585 173.225 38.835 174.025 ;
        RECT 39.480 173.055 39.810 173.855 ;
        RECT 40.110 173.225 40.440 174.025 ;
        RECT 40.610 173.055 40.940 173.855 ;
        RECT 38.505 172.885 40.940 173.055 ;
        RECT 41.315 172.885 41.655 173.855 ;
        RECT 41.825 172.885 41.995 174.025 ;
        RECT 42.265 173.225 42.515 174.025 ;
        RECT 43.160 173.055 43.490 173.855 ;
        RECT 43.790 173.225 44.120 174.025 ;
        RECT 44.290 173.055 44.620 173.855 ;
        RECT 42.185 172.885 44.620 173.055 ;
        RECT 45.200 173.055 45.530 173.855 ;
        RECT 45.700 173.225 46.030 174.025 ;
        RECT 46.330 173.055 46.660 173.855 ;
        RECT 47.305 173.225 47.555 174.025 ;
        RECT 45.200 172.885 47.635 173.055 ;
        RECT 47.825 172.885 47.995 174.025 ;
        RECT 48.165 172.885 48.505 173.855 ;
        RECT 48.790 173.395 49.075 173.855 ;
        RECT 49.245 173.565 49.515 174.025 ;
        RECT 48.790 173.175 49.745 173.395 ;
        RECT 32.075 171.475 32.585 172.010 ;
        RECT 32.805 171.680 33.050 172.285 ;
        RECT 34.875 172.245 35.625 172.765 ;
        RECT 33.955 171.475 35.625 172.245 ;
        RECT 35.795 171.475 36.085 172.200 ;
        RECT 36.315 171.475 36.525 172.295 ;
        RECT 36.695 172.275 36.945 172.875 ;
        RECT 37.115 172.465 37.445 172.715 ;
        RECT 36.695 171.645 37.025 172.275 ;
        RECT 37.195 171.475 37.425 172.295 ;
        RECT 37.635 172.275 37.810 172.885 ;
        RECT 38.505 172.635 38.675 172.885 ;
        RECT 37.980 172.465 38.675 172.635 ;
        RECT 38.850 172.465 39.270 172.665 ;
        RECT 39.440 172.465 39.770 172.665 ;
        RECT 39.940 172.465 40.270 172.665 ;
        RECT 37.635 171.645 37.975 172.275 ;
        RECT 38.145 171.475 38.395 172.275 ;
        RECT 38.585 172.125 39.810 172.295 ;
        RECT 38.585 171.645 38.915 172.125 ;
        RECT 39.085 171.475 39.310 171.935 ;
        RECT 39.480 171.645 39.810 172.125 ;
        RECT 40.440 172.255 40.610 172.885 ;
        RECT 40.795 172.465 41.145 172.715 ;
        RECT 41.315 172.275 41.490 172.885 ;
        RECT 42.185 172.635 42.355 172.885 ;
        RECT 41.660 172.465 42.355 172.635 ;
        RECT 42.530 172.465 42.950 172.665 ;
        RECT 43.120 172.465 43.450 172.665 ;
        RECT 43.620 172.465 43.950 172.665 ;
        RECT 40.440 171.645 40.940 172.255 ;
        RECT 41.315 171.645 41.655 172.275 ;
        RECT 41.825 171.475 42.075 172.275 ;
        RECT 42.265 172.125 43.490 172.295 ;
        RECT 42.265 171.645 42.595 172.125 ;
        RECT 42.765 171.475 42.990 171.935 ;
        RECT 43.160 171.645 43.490 172.125 ;
        RECT 44.120 172.255 44.290 172.885 ;
        RECT 44.475 172.465 44.825 172.715 ;
        RECT 44.995 172.465 45.345 172.715 ;
        RECT 45.530 172.255 45.700 172.885 ;
        RECT 45.870 172.465 46.200 172.665 ;
        RECT 46.370 172.465 46.700 172.665 ;
        RECT 46.870 172.465 47.290 172.665 ;
        RECT 47.465 172.635 47.635 172.885 ;
        RECT 47.465 172.465 48.160 172.635 ;
        RECT 44.120 171.645 44.620 172.255 ;
        RECT 45.200 171.645 45.700 172.255 ;
        RECT 46.330 172.125 47.555 172.295 ;
        RECT 48.330 172.275 48.505 172.885 ;
        RECT 48.675 172.445 49.365 173.005 ;
        RECT 49.535 172.275 49.745 173.175 ;
        RECT 46.330 171.645 46.660 172.125 ;
        RECT 46.830 171.475 47.055 171.935 ;
        RECT 47.225 171.645 47.555 172.125 ;
        RECT 47.745 171.475 47.995 172.275 ;
        RECT 48.165 171.645 48.505 172.275 ;
        RECT 48.790 172.105 49.745 172.275 ;
        RECT 49.915 173.005 50.315 173.855 ;
        RECT 50.505 173.395 50.785 173.855 ;
        RECT 51.305 173.565 51.630 174.025 ;
        RECT 50.505 173.175 51.630 173.395 ;
        RECT 49.915 172.445 51.010 173.005 ;
        RECT 51.180 172.715 51.630 173.175 ;
        RECT 51.800 172.885 52.185 173.855 ;
        RECT 48.790 171.645 49.075 172.105 ;
        RECT 49.245 171.475 49.515 171.935 ;
        RECT 49.915 171.645 50.315 172.445 ;
        RECT 51.180 172.385 51.735 172.715 ;
        RECT 51.180 172.275 51.630 172.385 ;
        RECT 50.505 172.105 51.630 172.275 ;
        RECT 51.905 172.215 52.185 172.885 ;
        RECT 50.505 171.645 50.785 172.105 ;
        RECT 51.305 171.475 51.630 171.935 ;
        RECT 51.800 171.645 52.185 172.215 ;
        RECT 52.360 172.835 52.615 173.715 ;
        RECT 52.785 172.885 53.090 174.025 ;
        RECT 53.430 173.645 53.760 174.025 ;
        RECT 53.940 173.475 54.110 173.765 ;
        RECT 54.280 173.565 54.530 174.025 ;
        RECT 53.310 173.305 54.110 173.475 ;
        RECT 54.700 173.515 55.570 173.855 ;
        RECT 52.360 172.185 52.570 172.835 ;
        RECT 53.310 172.715 53.480 173.305 ;
        RECT 54.700 173.135 54.870 173.515 ;
        RECT 55.805 173.395 55.975 173.855 ;
        RECT 56.145 173.565 56.515 174.025 ;
        RECT 56.810 173.425 56.980 173.765 ;
        RECT 57.150 173.595 57.480 174.025 ;
        RECT 57.715 173.425 57.885 173.765 ;
        RECT 53.650 172.965 54.870 173.135 ;
        RECT 55.040 173.055 55.500 173.345 ;
        RECT 55.805 173.225 56.365 173.395 ;
        RECT 56.810 173.255 57.885 173.425 ;
        RECT 58.055 173.525 58.735 173.855 ;
        RECT 58.950 173.525 59.200 173.855 ;
        RECT 59.370 173.565 59.620 174.025 ;
        RECT 56.195 173.085 56.365 173.225 ;
        RECT 55.040 173.045 56.005 173.055 ;
        RECT 54.700 172.875 54.870 172.965 ;
        RECT 55.330 172.885 56.005 173.045 ;
        RECT 52.740 172.685 53.480 172.715 ;
        RECT 52.740 172.385 53.655 172.685 ;
        RECT 53.330 172.210 53.655 172.385 ;
        RECT 52.360 171.655 52.615 172.185 ;
        RECT 52.785 171.475 53.090 171.935 ;
        RECT 53.335 171.855 53.655 172.210 ;
        RECT 53.825 172.425 54.365 172.795 ;
        RECT 54.700 172.705 55.105 172.875 ;
        RECT 53.825 172.025 54.065 172.425 ;
        RECT 54.545 172.255 54.765 172.535 ;
        RECT 54.235 172.085 54.765 172.255 ;
        RECT 54.235 171.855 54.405 172.085 ;
        RECT 54.935 171.925 55.105 172.705 ;
        RECT 55.275 172.095 55.625 172.715 ;
        RECT 55.795 172.095 56.005 172.885 ;
        RECT 56.195 172.915 57.695 173.085 ;
        RECT 56.195 172.225 56.365 172.915 ;
        RECT 58.055 172.745 58.225 173.525 ;
        RECT 59.030 173.395 59.200 173.525 ;
        RECT 56.535 172.575 58.225 172.745 ;
        RECT 58.395 172.965 58.860 173.355 ;
        RECT 59.030 173.225 59.425 173.395 ;
        RECT 56.535 172.395 56.705 172.575 ;
        RECT 53.335 171.685 54.405 171.855 ;
        RECT 54.575 171.475 54.765 171.915 ;
        RECT 54.935 171.645 55.885 171.925 ;
        RECT 56.195 171.835 56.455 172.225 ;
        RECT 56.875 172.155 57.665 172.405 ;
        RECT 56.105 171.665 56.455 171.835 ;
        RECT 56.665 171.475 56.995 171.935 ;
        RECT 57.870 171.865 58.040 172.575 ;
        RECT 58.395 172.375 58.565 172.965 ;
        RECT 58.210 172.155 58.565 172.375 ;
        RECT 58.735 172.155 59.085 172.775 ;
        RECT 59.255 171.865 59.425 173.225 ;
        RECT 59.790 173.055 60.115 173.840 ;
        RECT 59.595 172.005 60.055 173.055 ;
        RECT 57.870 171.695 58.725 171.865 ;
        RECT 58.930 171.695 59.425 171.865 ;
        RECT 59.595 171.475 59.925 171.835 ;
        RECT 60.285 171.735 60.455 173.855 ;
        RECT 60.625 173.525 60.955 174.025 ;
        RECT 61.125 173.355 61.380 173.855 ;
        RECT 60.630 173.185 61.380 173.355 ;
        RECT 60.630 172.195 60.860 173.185 ;
        RECT 61.030 172.365 61.380 173.015 ;
        RECT 61.555 172.860 61.845 174.025 ;
        RECT 62.015 172.950 62.285 173.855 ;
        RECT 62.455 173.265 62.785 174.025 ;
        RECT 62.965 173.095 63.135 173.855 ;
        RECT 60.630 172.025 61.380 172.195 ;
        RECT 60.625 171.475 60.955 171.855 ;
        RECT 61.125 171.735 61.380 172.025 ;
        RECT 61.555 171.475 61.845 172.200 ;
        RECT 62.015 172.150 62.185 172.950 ;
        RECT 62.470 172.925 63.135 173.095 ;
        RECT 62.470 172.780 62.640 172.925 ;
        RECT 64.320 172.875 64.580 174.025 ;
        RECT 64.755 172.950 65.010 173.855 ;
        RECT 65.180 173.265 65.510 174.025 ;
        RECT 65.725 173.095 65.895 173.855 ;
        RECT 66.620 173.590 71.965 174.025 ;
        RECT 62.355 172.450 62.640 172.780 ;
        RECT 62.470 172.195 62.640 172.450 ;
        RECT 62.875 172.375 63.205 172.745 ;
        RECT 62.015 171.645 62.275 172.150 ;
        RECT 62.470 172.025 63.135 172.195 ;
        RECT 62.455 171.475 62.785 171.855 ;
        RECT 62.965 171.645 63.135 172.025 ;
        RECT 64.320 171.475 64.580 172.315 ;
        RECT 64.755 172.220 64.925 172.950 ;
        RECT 65.180 172.925 65.895 173.095 ;
        RECT 65.180 172.715 65.350 172.925 ;
        RECT 65.095 172.385 65.350 172.715 ;
        RECT 64.755 171.645 65.010 172.220 ;
        RECT 65.180 172.195 65.350 172.385 ;
        RECT 65.630 172.375 65.985 172.745 ;
        RECT 68.210 172.340 68.560 173.590 ;
        RECT 72.225 173.355 72.395 173.855 ;
        RECT 72.565 173.525 72.895 174.025 ;
        RECT 72.225 173.185 72.890 173.355 ;
        RECT 65.180 172.025 65.895 172.195 ;
        RECT 65.180 171.475 65.510 171.855 ;
        RECT 65.725 171.645 65.895 172.025 ;
        RECT 70.040 172.020 70.380 172.850 ;
        RECT 72.140 172.365 72.490 173.015 ;
        RECT 72.660 172.195 72.890 173.185 ;
        RECT 72.225 172.025 72.890 172.195 ;
        RECT 66.620 171.475 71.965 172.020 ;
        RECT 72.225 171.735 72.395 172.025 ;
        RECT 72.565 171.475 72.895 171.855 ;
        RECT 73.065 171.735 73.290 173.855 ;
        RECT 73.505 173.525 73.835 174.025 ;
        RECT 74.005 173.355 74.175 173.855 ;
        RECT 74.410 173.640 75.240 173.810 ;
        RECT 75.480 173.645 75.860 174.025 ;
        RECT 73.480 173.185 74.175 173.355 ;
        RECT 73.480 172.215 73.650 173.185 ;
        RECT 73.820 172.395 74.230 173.015 ;
        RECT 74.400 172.965 74.900 173.345 ;
        RECT 73.480 172.025 74.175 172.215 ;
        RECT 74.400 172.095 74.620 172.965 ;
        RECT 75.070 172.795 75.240 173.640 ;
        RECT 76.040 173.475 76.210 173.765 ;
        RECT 76.380 173.645 76.710 174.025 ;
        RECT 77.180 173.555 77.810 173.805 ;
        RECT 77.990 173.645 78.410 174.025 ;
        RECT 77.640 173.475 77.810 173.555 ;
        RECT 78.610 173.475 78.850 173.765 ;
        RECT 75.410 173.225 76.780 173.475 ;
        RECT 75.410 172.965 75.660 173.225 ;
        RECT 76.170 172.795 76.420 172.955 ;
        RECT 75.070 172.625 76.420 172.795 ;
        RECT 75.070 172.585 75.490 172.625 ;
        RECT 74.800 172.035 75.150 172.405 ;
        RECT 73.505 171.475 73.835 171.855 ;
        RECT 74.005 171.695 74.175 172.025 ;
        RECT 75.320 171.855 75.490 172.585 ;
        RECT 76.590 172.455 76.780 173.225 ;
        RECT 75.660 172.125 76.070 172.455 ;
        RECT 76.360 172.115 76.780 172.455 ;
        RECT 76.950 173.045 77.470 173.355 ;
        RECT 77.640 173.305 78.850 173.475 ;
        RECT 79.080 173.335 79.410 174.025 ;
        RECT 76.950 172.285 77.120 173.045 ;
        RECT 77.290 172.455 77.470 172.865 ;
        RECT 77.640 172.795 77.810 173.305 ;
        RECT 79.580 173.155 79.750 173.765 ;
        RECT 80.020 173.305 80.350 173.815 ;
        RECT 79.580 173.135 79.900 173.155 ;
        RECT 77.980 172.965 79.900 173.135 ;
        RECT 77.640 172.625 79.540 172.795 ;
        RECT 77.870 172.285 78.200 172.405 ;
        RECT 76.950 172.115 78.200 172.285 ;
        RECT 74.475 171.655 75.490 171.855 ;
        RECT 75.660 171.475 76.070 171.915 ;
        RECT 76.360 171.685 76.610 172.115 ;
        RECT 76.810 171.475 77.130 171.935 ;
        RECT 78.370 171.865 78.540 172.625 ;
        RECT 79.210 172.565 79.540 172.625 ;
        RECT 78.730 172.395 79.060 172.455 ;
        RECT 78.730 172.125 79.390 172.395 ;
        RECT 79.710 172.070 79.900 172.965 ;
        RECT 77.690 171.695 78.540 171.865 ;
        RECT 78.740 171.475 79.400 171.955 ;
        RECT 79.580 171.740 79.900 172.070 ;
        RECT 80.100 172.715 80.350 173.305 ;
        RECT 80.530 173.225 80.815 174.025 ;
        RECT 80.995 173.045 81.250 173.715 ;
        RECT 80.100 172.385 80.900 172.715 ;
        RECT 80.100 171.735 80.350 172.385 ;
        RECT 81.070 172.185 81.250 173.045 ;
        RECT 81.835 172.885 82.065 174.025 ;
        RECT 82.235 172.875 82.565 173.855 ;
        RECT 82.735 172.885 82.945 174.025 ;
        RECT 83.175 173.265 83.690 173.675 ;
        RECT 83.925 173.265 84.095 174.025 ;
        RECT 84.265 173.685 86.295 173.855 ;
        RECT 81.815 172.465 82.145 172.715 ;
        RECT 80.995 171.985 81.250 172.185 ;
        RECT 80.530 171.475 80.815 171.935 ;
        RECT 80.995 171.815 81.335 171.985 ;
        RECT 80.995 171.655 81.250 171.815 ;
        RECT 81.835 171.475 82.065 172.295 ;
        RECT 82.315 172.275 82.565 172.875 ;
        RECT 83.175 172.455 83.515 173.265 ;
        RECT 84.265 173.020 84.435 173.685 ;
        RECT 84.830 173.345 85.955 173.515 ;
        RECT 83.685 172.830 84.435 173.020 ;
        RECT 84.605 173.005 85.615 173.175 ;
        RECT 82.235 171.645 82.565 172.275 ;
        RECT 82.735 171.475 82.945 172.295 ;
        RECT 83.175 172.285 84.405 172.455 ;
        RECT 83.450 171.680 83.695 172.285 ;
        RECT 83.915 171.475 84.425 172.010 ;
        RECT 84.605 171.645 84.795 173.005 ;
        RECT 84.965 171.985 85.240 172.805 ;
        RECT 85.445 172.205 85.615 173.005 ;
        RECT 85.785 172.215 85.955 173.345 ;
        RECT 86.125 172.715 86.295 173.685 ;
        RECT 86.465 172.885 86.635 174.025 ;
        RECT 86.805 172.885 87.140 173.855 ;
        RECT 86.125 172.385 86.320 172.715 ;
        RECT 86.545 172.385 86.800 172.715 ;
        RECT 86.545 172.215 86.715 172.385 ;
        RECT 86.970 172.215 87.140 172.885 ;
        RECT 87.315 172.860 87.605 174.025 ;
        RECT 87.775 172.885 88.160 173.855 ;
        RECT 88.330 173.565 88.655 174.025 ;
        RECT 89.175 173.395 89.455 173.855 ;
        RECT 88.330 173.175 89.455 173.395 ;
        RECT 85.785 172.045 86.715 172.215 ;
        RECT 85.785 172.010 85.960 172.045 ;
        RECT 84.965 171.815 85.245 171.985 ;
        RECT 84.965 171.645 85.240 171.815 ;
        RECT 85.430 171.645 85.960 172.010 ;
        RECT 86.385 171.475 86.715 171.875 ;
        RECT 86.885 171.645 87.140 172.215 ;
        RECT 87.775 172.215 88.055 172.885 ;
        RECT 88.330 172.715 88.780 173.175 ;
        RECT 89.645 173.005 90.045 173.855 ;
        RECT 90.445 173.565 90.715 174.025 ;
        RECT 90.885 173.395 91.170 173.855 ;
        RECT 88.225 172.385 88.780 172.715 ;
        RECT 88.950 172.445 90.045 173.005 ;
        RECT 88.330 172.275 88.780 172.385 ;
        RECT 87.315 171.475 87.605 172.200 ;
        RECT 87.775 171.645 88.160 172.215 ;
        RECT 88.330 172.105 89.455 172.275 ;
        RECT 88.330 171.475 88.655 171.935 ;
        RECT 89.175 171.645 89.455 172.105 ;
        RECT 89.645 171.645 90.045 172.445 ;
        RECT 90.215 173.175 91.170 173.395 ;
        RECT 90.215 172.275 90.425 173.175 ;
        RECT 91.660 173.055 91.990 173.855 ;
        RECT 92.160 173.225 92.490 174.025 ;
        RECT 92.790 173.055 93.120 173.855 ;
        RECT 93.765 173.225 94.015 174.025 ;
        RECT 90.595 172.445 91.285 173.005 ;
        RECT 91.660 172.885 94.095 173.055 ;
        RECT 94.285 172.885 94.455 174.025 ;
        RECT 94.625 172.885 94.965 173.855 ;
        RECT 91.455 172.465 91.805 172.715 ;
        RECT 90.215 172.105 91.170 172.275 ;
        RECT 91.990 172.255 92.160 172.885 ;
        RECT 92.330 172.465 92.660 172.665 ;
        RECT 92.830 172.465 93.160 172.665 ;
        RECT 93.330 172.465 93.750 172.665 ;
        RECT 93.925 172.635 94.095 172.885 ;
        RECT 93.925 172.465 94.620 172.635 ;
        RECT 94.790 172.325 94.965 172.885 ;
        RECT 90.445 171.475 90.715 171.935 ;
        RECT 90.885 171.645 91.170 172.105 ;
        RECT 91.660 171.645 92.160 172.255 ;
        RECT 92.790 172.125 94.015 172.295 ;
        RECT 94.735 172.275 94.965 172.325 ;
        RECT 92.790 171.645 93.120 172.125 ;
        RECT 93.290 171.475 93.515 171.935 ;
        RECT 93.685 171.645 94.015 172.125 ;
        RECT 94.205 171.475 94.455 172.275 ;
        RECT 94.625 171.645 94.965 172.275 ;
        RECT 95.135 172.885 95.475 173.855 ;
        RECT 95.645 172.885 95.815 174.025 ;
        RECT 96.085 173.225 96.335 174.025 ;
        RECT 96.980 173.055 97.310 173.855 ;
        RECT 97.610 173.225 97.940 174.025 ;
        RECT 98.110 173.055 98.440 173.855 ;
        RECT 96.005 172.885 98.440 173.055 ;
        RECT 99.315 172.885 99.545 174.025 ;
        RECT 95.135 172.835 95.365 172.885 ;
        RECT 95.135 172.275 95.310 172.835 ;
        RECT 96.005 172.635 96.175 172.885 ;
        RECT 95.480 172.465 96.175 172.635 ;
        RECT 96.350 172.465 96.770 172.665 ;
        RECT 96.940 172.465 97.270 172.665 ;
        RECT 97.440 172.465 97.770 172.665 ;
        RECT 95.135 171.645 95.475 172.275 ;
        RECT 95.645 171.475 95.895 172.275 ;
        RECT 96.085 172.125 97.310 172.295 ;
        RECT 96.085 171.645 96.415 172.125 ;
        RECT 96.585 171.475 96.810 171.935 ;
        RECT 96.980 171.645 97.310 172.125 ;
        RECT 97.940 172.255 98.110 172.885 ;
        RECT 99.715 172.875 100.045 173.855 ;
        RECT 100.215 172.885 100.425 174.025 ;
        RECT 100.695 172.885 100.925 174.025 ;
        RECT 101.095 172.875 101.425 173.855 ;
        RECT 101.595 172.885 101.805 174.025 ;
        RECT 98.295 172.465 98.645 172.715 ;
        RECT 99.295 172.465 99.625 172.715 ;
        RECT 97.940 171.645 98.440 172.255 ;
        RECT 99.315 171.475 99.545 172.295 ;
        RECT 99.795 172.275 100.045 172.875 ;
        RECT 100.675 172.465 101.005 172.715 ;
        RECT 99.715 171.645 100.045 172.275 ;
        RECT 100.215 171.475 100.425 172.295 ;
        RECT 100.695 171.475 100.925 172.295 ;
        RECT 101.175 172.275 101.425 172.875 ;
        RECT 102.040 172.835 102.295 173.715 ;
        RECT 102.465 172.885 102.770 174.025 ;
        RECT 103.110 173.645 103.440 174.025 ;
        RECT 103.620 173.475 103.790 173.765 ;
        RECT 103.960 173.565 104.210 174.025 ;
        RECT 102.990 173.305 103.790 173.475 ;
        RECT 104.380 173.515 105.250 173.855 ;
        RECT 101.095 171.645 101.425 172.275 ;
        RECT 101.595 171.475 101.805 172.295 ;
        RECT 102.040 172.185 102.250 172.835 ;
        RECT 102.990 172.715 103.160 173.305 ;
        RECT 104.380 173.135 104.550 173.515 ;
        RECT 105.485 173.395 105.655 173.855 ;
        RECT 105.825 173.565 106.195 174.025 ;
        RECT 106.490 173.425 106.660 173.765 ;
        RECT 106.830 173.595 107.160 174.025 ;
        RECT 107.395 173.425 107.565 173.765 ;
        RECT 103.330 172.965 104.550 173.135 ;
        RECT 104.720 173.055 105.180 173.345 ;
        RECT 105.485 173.225 106.045 173.395 ;
        RECT 106.490 173.255 107.565 173.425 ;
        RECT 107.735 173.525 108.415 173.855 ;
        RECT 108.630 173.525 108.880 173.855 ;
        RECT 109.050 173.565 109.300 174.025 ;
        RECT 105.875 173.085 106.045 173.225 ;
        RECT 104.720 173.045 105.685 173.055 ;
        RECT 104.380 172.875 104.550 172.965 ;
        RECT 105.010 172.885 105.685 173.045 ;
        RECT 102.420 172.685 103.160 172.715 ;
        RECT 102.420 172.385 103.335 172.685 ;
        RECT 103.010 172.210 103.335 172.385 ;
        RECT 102.040 171.655 102.295 172.185 ;
        RECT 102.465 171.475 102.770 171.935 ;
        RECT 103.015 171.855 103.335 172.210 ;
        RECT 103.505 172.425 104.045 172.795 ;
        RECT 104.380 172.705 104.785 172.875 ;
        RECT 103.505 172.025 103.745 172.425 ;
        RECT 104.225 172.255 104.445 172.535 ;
        RECT 103.915 172.085 104.445 172.255 ;
        RECT 103.915 171.855 104.085 172.085 ;
        RECT 104.615 171.925 104.785 172.705 ;
        RECT 104.955 172.095 105.305 172.715 ;
        RECT 105.475 172.095 105.685 172.885 ;
        RECT 105.875 172.915 107.375 173.085 ;
        RECT 105.875 172.225 106.045 172.915 ;
        RECT 107.735 172.745 107.905 173.525 ;
        RECT 108.710 173.395 108.880 173.525 ;
        RECT 106.215 172.575 107.905 172.745 ;
        RECT 108.075 172.965 108.540 173.355 ;
        RECT 108.710 173.225 109.105 173.395 ;
        RECT 106.215 172.395 106.385 172.575 ;
        RECT 103.015 171.685 104.085 171.855 ;
        RECT 104.255 171.475 104.445 171.915 ;
        RECT 104.615 171.645 105.565 171.925 ;
        RECT 105.875 171.835 106.135 172.225 ;
        RECT 106.555 172.155 107.345 172.405 ;
        RECT 105.785 171.665 106.135 171.835 ;
        RECT 106.345 171.475 106.675 171.935 ;
        RECT 107.550 171.865 107.720 172.575 ;
        RECT 108.075 172.375 108.245 172.965 ;
        RECT 107.890 172.155 108.245 172.375 ;
        RECT 108.415 172.155 108.765 172.775 ;
        RECT 108.935 171.865 109.105 173.225 ;
        RECT 109.470 173.055 109.795 173.840 ;
        RECT 109.275 172.005 109.735 173.055 ;
        RECT 107.550 171.695 108.405 171.865 ;
        RECT 108.610 171.695 109.105 171.865 ;
        RECT 109.275 171.475 109.605 171.835 ;
        RECT 109.965 171.735 110.135 173.855 ;
        RECT 110.305 173.525 110.635 174.025 ;
        RECT 110.805 173.355 111.060 173.855 ;
        RECT 110.310 173.185 111.060 173.355 ;
        RECT 110.310 172.195 110.540 173.185 ;
        RECT 110.710 172.365 111.060 173.015 ;
        RECT 112.155 172.935 113.365 174.025 ;
        RECT 112.155 172.395 112.675 172.935 ;
        RECT 112.845 172.225 113.365 172.765 ;
        RECT 110.310 172.025 111.060 172.195 ;
        RECT 110.305 171.475 110.635 171.855 ;
        RECT 110.805 171.735 111.060 172.025 ;
        RECT 112.155 171.475 113.365 172.225 ;
        RECT 15.010 171.305 113.450 171.475 ;
        RECT 15.095 170.555 16.305 171.305 ;
        RECT 16.475 170.555 17.685 171.305 ;
        RECT 15.095 170.015 15.615 170.555 ;
        RECT 15.785 169.845 16.305 170.385 ;
        RECT 15.095 168.755 16.305 169.845 ;
        RECT 16.475 169.845 16.995 170.385 ;
        RECT 17.165 170.015 17.685 170.555 ;
        RECT 17.915 170.485 18.125 171.305 ;
        RECT 18.295 170.505 18.625 171.135 ;
        RECT 18.295 169.905 18.545 170.505 ;
        RECT 18.795 170.485 19.025 171.305 ;
        RECT 19.350 170.675 19.635 171.135 ;
        RECT 19.805 170.845 20.075 171.305 ;
        RECT 19.350 170.505 20.305 170.675 ;
        RECT 18.715 170.065 19.045 170.315 ;
        RECT 16.475 168.755 17.685 169.845 ;
        RECT 17.915 168.755 18.125 169.895 ;
        RECT 18.295 168.925 18.625 169.905 ;
        RECT 18.795 168.755 19.025 169.895 ;
        RECT 19.235 169.775 19.925 170.335 ;
        RECT 20.095 169.605 20.305 170.505 ;
        RECT 19.350 169.385 20.305 169.605 ;
        RECT 20.475 170.335 20.875 171.135 ;
        RECT 21.065 170.675 21.345 171.135 ;
        RECT 21.865 170.845 22.190 171.305 ;
        RECT 21.065 170.505 22.190 170.675 ;
        RECT 22.360 170.565 22.745 171.135 ;
        RECT 22.915 170.580 23.205 171.305 ;
        RECT 21.740 170.395 22.190 170.505 ;
        RECT 20.475 169.775 21.570 170.335 ;
        RECT 21.740 170.065 22.295 170.395 ;
        RECT 19.350 168.925 19.635 169.385 ;
        RECT 19.805 168.755 20.075 169.215 ;
        RECT 20.475 168.925 20.875 169.775 ;
        RECT 21.740 169.605 22.190 170.065 ;
        RECT 22.465 169.895 22.745 170.565 ;
        RECT 23.835 170.535 25.505 171.305 ;
        RECT 21.065 169.385 22.190 169.605 ;
        RECT 21.065 168.925 21.345 169.385 ;
        RECT 21.865 168.755 22.190 169.215 ;
        RECT 22.360 168.925 22.745 169.895 ;
        RECT 22.915 168.755 23.205 169.920 ;
        RECT 23.835 169.845 24.585 170.365 ;
        RECT 24.755 170.015 25.505 170.535 ;
        RECT 25.790 170.675 26.075 171.135 ;
        RECT 26.245 170.845 26.515 171.305 ;
        RECT 25.790 170.505 26.745 170.675 ;
        RECT 23.835 168.755 25.505 169.845 ;
        RECT 25.675 169.775 26.365 170.335 ;
        RECT 26.535 169.605 26.745 170.505 ;
        RECT 25.790 169.385 26.745 169.605 ;
        RECT 26.915 170.335 27.315 171.135 ;
        RECT 27.505 170.675 27.785 171.135 ;
        RECT 28.305 170.845 28.630 171.305 ;
        RECT 27.505 170.505 28.630 170.675 ;
        RECT 28.800 170.565 29.185 171.135 ;
        RECT 28.180 170.395 28.630 170.505 ;
        RECT 26.915 169.775 28.010 170.335 ;
        RECT 28.180 170.065 28.735 170.395 ;
        RECT 25.790 168.925 26.075 169.385 ;
        RECT 26.245 168.755 26.515 169.215 ;
        RECT 26.915 168.925 27.315 169.775 ;
        RECT 28.180 169.605 28.630 170.065 ;
        RECT 28.905 169.895 29.185 170.565 ;
        RECT 27.505 169.385 28.630 169.605 ;
        RECT 27.505 168.925 27.785 169.385 ;
        RECT 28.305 168.755 28.630 169.215 ;
        RECT 28.800 168.925 29.185 169.895 ;
        RECT 30.275 170.505 30.615 171.135 ;
        RECT 30.785 170.505 31.035 171.305 ;
        RECT 31.225 170.655 31.555 171.135 ;
        RECT 31.725 170.845 31.950 171.305 ;
        RECT 32.120 170.655 32.450 171.135 ;
        RECT 30.275 169.895 30.450 170.505 ;
        RECT 31.225 170.485 32.450 170.655 ;
        RECT 33.080 170.525 33.580 171.135 ;
        RECT 30.620 170.145 31.315 170.315 ;
        RECT 31.145 169.895 31.315 170.145 ;
        RECT 31.490 170.115 31.910 170.315 ;
        RECT 32.080 170.115 32.410 170.315 ;
        RECT 32.580 170.115 32.910 170.315 ;
        RECT 33.080 169.895 33.250 170.525 ;
        RECT 33.955 170.505 34.295 171.135 ;
        RECT 34.465 170.505 34.715 171.305 ;
        RECT 34.905 170.655 35.235 171.135 ;
        RECT 35.405 170.845 35.630 171.305 ;
        RECT 35.800 170.655 36.130 171.135 ;
        RECT 33.435 170.065 33.785 170.315 ;
        RECT 33.955 169.945 34.130 170.505 ;
        RECT 34.905 170.485 36.130 170.655 ;
        RECT 36.760 170.525 37.260 171.135 ;
        RECT 34.300 170.145 34.995 170.315 ;
        RECT 33.955 169.895 34.185 169.945 ;
        RECT 34.825 169.895 34.995 170.145 ;
        RECT 35.170 170.115 35.590 170.315 ;
        RECT 35.760 170.115 36.090 170.315 ;
        RECT 36.260 170.115 36.590 170.315 ;
        RECT 36.760 169.895 36.930 170.525 ;
        RECT 37.635 170.505 37.975 171.135 ;
        RECT 38.145 170.505 38.395 171.305 ;
        RECT 38.585 170.655 38.915 171.135 ;
        RECT 39.085 170.845 39.310 171.305 ;
        RECT 39.480 170.655 39.810 171.135 ;
        RECT 37.115 170.065 37.465 170.315 ;
        RECT 37.635 169.895 37.810 170.505 ;
        RECT 38.585 170.485 39.810 170.655 ;
        RECT 40.440 170.525 40.940 171.135 ;
        RECT 41.315 170.630 41.575 171.135 ;
        RECT 41.755 170.925 42.085 171.305 ;
        RECT 42.265 170.755 42.435 171.135 ;
        RECT 37.980 170.145 38.675 170.315 ;
        RECT 38.505 169.895 38.675 170.145 ;
        RECT 38.850 170.115 39.270 170.315 ;
        RECT 39.440 170.115 39.770 170.315 ;
        RECT 39.940 170.115 40.270 170.315 ;
        RECT 40.440 169.895 40.610 170.525 ;
        RECT 40.795 170.065 41.145 170.315 ;
        RECT 30.275 168.925 30.615 169.895 ;
        RECT 30.785 168.755 30.955 169.895 ;
        RECT 31.145 169.725 33.580 169.895 ;
        RECT 31.225 168.755 31.475 169.555 ;
        RECT 32.120 168.925 32.450 169.725 ;
        RECT 32.750 168.755 33.080 169.555 ;
        RECT 33.250 168.925 33.580 169.725 ;
        RECT 33.955 168.925 34.295 169.895 ;
        RECT 34.465 168.755 34.635 169.895 ;
        RECT 34.825 169.725 37.260 169.895 ;
        RECT 34.905 168.755 35.155 169.555 ;
        RECT 35.800 168.925 36.130 169.725 ;
        RECT 36.430 168.755 36.760 169.555 ;
        RECT 36.930 168.925 37.260 169.725 ;
        RECT 37.635 168.925 37.975 169.895 ;
        RECT 38.145 168.755 38.315 169.895 ;
        RECT 38.505 169.725 40.940 169.895 ;
        RECT 38.585 168.755 38.835 169.555 ;
        RECT 39.480 168.925 39.810 169.725 ;
        RECT 40.110 168.755 40.440 169.555 ;
        RECT 40.610 168.925 40.940 169.725 ;
        RECT 41.315 169.830 41.485 170.630 ;
        RECT 41.770 170.585 42.435 170.755 ;
        RECT 41.770 170.330 41.940 170.585 ;
        RECT 42.695 170.535 44.365 171.305 ;
        RECT 41.655 170.000 41.940 170.330 ;
        RECT 42.175 170.035 42.505 170.405 ;
        RECT 41.770 169.855 41.940 170.000 ;
        RECT 41.315 168.925 41.585 169.830 ;
        RECT 41.770 169.685 42.435 169.855 ;
        RECT 41.755 168.755 42.085 169.515 ;
        RECT 42.265 168.925 42.435 169.685 ;
        RECT 42.695 169.845 43.445 170.365 ;
        RECT 43.615 170.015 44.365 170.535 ;
        RECT 44.540 170.565 44.795 171.135 ;
        RECT 44.965 170.905 45.295 171.305 ;
        RECT 45.720 170.770 46.250 171.135 ;
        RECT 45.720 170.735 45.895 170.770 ;
        RECT 44.965 170.565 45.895 170.735 ;
        RECT 44.540 169.895 44.710 170.565 ;
        RECT 44.965 170.395 45.135 170.565 ;
        RECT 44.880 170.065 45.135 170.395 ;
        RECT 45.360 170.065 45.555 170.395 ;
        RECT 42.695 168.755 44.365 169.845 ;
        RECT 44.540 168.925 44.875 169.895 ;
        RECT 45.045 168.755 45.215 169.895 ;
        RECT 45.385 169.095 45.555 170.065 ;
        RECT 45.725 169.435 45.895 170.565 ;
        RECT 46.065 169.775 46.235 170.575 ;
        RECT 46.440 170.285 46.715 171.135 ;
        RECT 46.435 170.115 46.715 170.285 ;
        RECT 46.440 169.975 46.715 170.115 ;
        RECT 46.885 169.775 47.075 171.135 ;
        RECT 47.255 170.770 47.765 171.305 ;
        RECT 47.985 170.495 48.230 171.100 ;
        RECT 48.675 170.580 48.965 171.305 ;
        RECT 49.645 170.845 49.950 171.305 ;
        RECT 50.120 170.675 50.450 171.135 ;
        RECT 50.620 170.845 50.790 171.305 ;
        RECT 50.960 170.675 51.290 171.135 ;
        RECT 51.460 170.845 51.630 171.305 ;
        RECT 51.800 170.675 52.130 171.135 ;
        RECT 52.300 170.845 52.470 171.305 ;
        RECT 52.640 170.675 52.970 171.135 ;
        RECT 53.140 170.845 53.395 171.305 ;
        RECT 47.275 170.325 48.505 170.495 ;
        RECT 46.065 169.605 47.075 169.775 ;
        RECT 47.245 169.760 47.995 169.950 ;
        RECT 45.725 169.265 46.850 169.435 ;
        RECT 47.245 169.095 47.415 169.760 ;
        RECT 48.165 169.515 48.505 170.325 ;
        RECT 49.595 170.485 53.565 170.675 ;
        RECT 53.735 170.535 57.245 171.305 ;
        RECT 45.385 168.925 47.415 169.095 ;
        RECT 47.585 168.755 47.755 169.515 ;
        RECT 47.990 169.105 48.505 169.515 ;
        RECT 48.675 168.755 48.965 169.920 ;
        RECT 49.595 169.895 49.915 170.485 ;
        RECT 50.115 170.285 52.970 170.315 ;
        RECT 50.115 170.115 53.045 170.285 ;
        RECT 50.115 170.065 52.970 170.115 ;
        RECT 53.220 169.895 53.565 170.485 ;
        RECT 49.595 169.725 53.565 169.895 ;
        RECT 53.735 169.845 55.425 170.365 ;
        RECT 55.595 170.015 57.245 170.535 ;
        RECT 57.475 170.485 57.685 171.305 ;
        RECT 57.855 170.505 58.185 171.135 ;
        RECT 57.855 169.905 58.105 170.505 ;
        RECT 58.355 170.485 58.585 171.305 ;
        RECT 59.255 170.535 62.765 171.305 ;
        RECT 58.275 170.065 58.605 170.315 ;
        RECT 49.650 168.755 49.950 169.555 ;
        RECT 50.120 168.925 50.450 169.725 ;
        RECT 50.620 168.755 50.790 169.555 ;
        RECT 50.960 168.925 51.290 169.725 ;
        RECT 51.460 168.755 51.630 169.555 ;
        RECT 51.800 168.925 52.130 169.725 ;
        RECT 52.300 168.755 52.470 169.555 ;
        RECT 52.640 168.925 52.970 169.725 ;
        RECT 53.140 168.755 53.395 169.555 ;
        RECT 53.735 168.755 57.245 169.845 ;
        RECT 57.475 168.755 57.685 169.895 ;
        RECT 57.855 168.925 58.185 169.905 ;
        RECT 58.355 168.755 58.585 169.895 ;
        RECT 59.255 169.845 60.945 170.365 ;
        RECT 61.115 170.015 62.765 170.535 ;
        RECT 62.940 170.465 63.200 171.305 ;
        RECT 63.375 170.560 63.630 171.135 ;
        RECT 63.800 170.925 64.130 171.305 ;
        RECT 64.345 170.755 64.515 171.135 ;
        RECT 63.800 170.585 64.515 170.755 ;
        RECT 64.775 170.805 65.075 171.135 ;
        RECT 65.245 170.825 65.520 171.305 ;
        RECT 59.255 168.755 62.765 169.845 ;
        RECT 62.940 168.755 63.200 169.905 ;
        RECT 63.375 169.830 63.545 170.560 ;
        RECT 63.800 170.395 63.970 170.585 ;
        RECT 63.715 170.065 63.970 170.395 ;
        RECT 63.800 169.855 63.970 170.065 ;
        RECT 64.250 170.035 64.605 170.405 ;
        RECT 64.775 169.895 64.945 170.805 ;
        RECT 65.700 170.655 65.995 171.045 ;
        RECT 66.165 170.825 66.420 171.305 ;
        RECT 66.595 170.655 66.855 171.045 ;
        RECT 67.025 170.825 67.305 171.305 ;
        RECT 65.115 170.065 65.465 170.635 ;
        RECT 65.700 170.485 67.350 170.655 ;
        RECT 67.595 170.485 67.805 171.305 ;
        RECT 67.975 170.505 68.305 171.135 ;
        RECT 65.635 170.145 66.775 170.315 ;
        RECT 65.635 169.895 65.805 170.145 ;
        RECT 66.945 169.975 67.350 170.485 ;
        RECT 63.375 168.925 63.630 169.830 ;
        RECT 63.800 169.685 64.515 169.855 ;
        RECT 63.800 168.755 64.130 169.515 ;
        RECT 64.345 168.925 64.515 169.685 ;
        RECT 64.775 169.725 65.805 169.895 ;
        RECT 66.595 169.805 67.350 169.975 ;
        RECT 67.975 169.905 68.225 170.505 ;
        RECT 68.475 170.485 68.705 171.305 ;
        RECT 69.005 170.755 69.175 171.135 ;
        RECT 69.355 170.925 69.685 171.305 ;
        RECT 69.005 170.585 69.670 170.755 ;
        RECT 69.865 170.630 70.125 171.135 ;
        RECT 68.395 170.065 68.725 170.315 ;
        RECT 68.935 170.035 69.265 170.405 ;
        RECT 69.500 170.330 69.670 170.585 ;
        RECT 69.500 170.000 69.785 170.330 ;
        RECT 64.775 168.925 65.085 169.725 ;
        RECT 66.595 169.555 66.855 169.805 ;
        RECT 65.255 168.755 65.565 169.555 ;
        RECT 65.735 169.385 66.855 169.555 ;
        RECT 65.735 168.925 65.995 169.385 ;
        RECT 66.165 168.755 66.420 169.215 ;
        RECT 66.595 168.925 66.855 169.385 ;
        RECT 67.025 168.755 67.310 169.625 ;
        RECT 67.595 168.755 67.805 169.895 ;
        RECT 67.975 168.925 68.305 169.905 ;
        RECT 68.475 168.755 68.705 169.895 ;
        RECT 69.500 169.855 69.670 170.000 ;
        RECT 69.005 169.685 69.670 169.855 ;
        RECT 69.955 169.830 70.125 170.630 ;
        RECT 69.005 168.925 69.175 169.685 ;
        RECT 69.355 168.755 69.685 169.515 ;
        RECT 69.855 168.925 70.125 169.830 ;
        RECT 70.300 170.565 70.555 171.135 ;
        RECT 70.725 170.905 71.055 171.305 ;
        RECT 71.480 170.770 72.010 171.135 ;
        RECT 71.480 170.735 71.655 170.770 ;
        RECT 70.725 170.565 71.655 170.735 ;
        RECT 70.300 169.895 70.470 170.565 ;
        RECT 70.725 170.395 70.895 170.565 ;
        RECT 70.640 170.065 70.895 170.395 ;
        RECT 71.120 170.065 71.315 170.395 ;
        RECT 70.300 168.925 70.635 169.895 ;
        RECT 70.805 168.755 70.975 169.895 ;
        RECT 71.145 169.095 71.315 170.065 ;
        RECT 71.485 169.435 71.655 170.565 ;
        RECT 71.825 169.775 71.995 170.575 ;
        RECT 72.200 170.285 72.475 171.135 ;
        RECT 72.195 170.115 72.475 170.285 ;
        RECT 72.200 169.975 72.475 170.115 ;
        RECT 72.645 169.775 72.835 171.135 ;
        RECT 73.015 170.770 73.525 171.305 ;
        RECT 73.745 170.495 73.990 171.100 ;
        RECT 74.435 170.580 74.725 171.305 ;
        RECT 75.005 170.825 75.175 171.305 ;
        RECT 75.345 170.655 75.675 171.130 ;
        RECT 75.845 170.825 76.015 171.305 ;
        RECT 76.185 170.655 76.515 171.130 ;
        RECT 76.685 170.825 76.855 171.305 ;
        RECT 77.025 170.655 77.355 171.130 ;
        RECT 77.525 170.825 77.695 171.305 ;
        RECT 77.865 170.655 78.195 171.130 ;
        RECT 78.365 170.825 78.535 171.305 ;
        RECT 78.705 170.655 79.035 171.130 ;
        RECT 79.205 170.825 79.375 171.305 ;
        RECT 79.625 171.130 79.795 171.135 ;
        RECT 79.545 170.655 79.875 171.130 ;
        RECT 80.045 170.825 80.215 171.305 ;
        RECT 80.465 171.130 80.635 171.135 ;
        RECT 80.385 170.655 80.715 171.130 ;
        RECT 80.885 170.825 81.055 171.305 ;
        RECT 81.305 171.130 81.555 171.135 ;
        RECT 81.225 170.655 81.555 171.130 ;
        RECT 81.725 170.825 81.895 171.305 ;
        RECT 82.065 170.655 82.395 171.130 ;
        RECT 82.565 170.825 82.735 171.305 ;
        RECT 82.905 170.655 83.235 171.130 ;
        RECT 83.405 170.825 83.575 171.305 ;
        RECT 83.745 170.655 84.075 171.130 ;
        RECT 84.245 170.825 84.415 171.305 ;
        RECT 84.585 170.655 84.915 171.130 ;
        RECT 85.085 170.825 85.255 171.305 ;
        RECT 85.425 170.655 85.755 171.130 ;
        RECT 73.035 170.325 74.265 170.495 ;
        RECT 71.825 169.605 72.835 169.775 ;
        RECT 73.005 169.760 73.755 169.950 ;
        RECT 71.485 169.265 72.610 169.435 ;
        RECT 73.005 169.095 73.175 169.760 ;
        RECT 73.925 169.515 74.265 170.325 ;
        RECT 74.895 170.485 81.555 170.655 ;
        RECT 81.725 170.485 84.075 170.655 ;
        RECT 84.245 170.485 85.755 170.655 ;
        RECT 85.935 170.535 87.605 171.305 ;
        RECT 74.895 169.945 75.170 170.485 ;
        RECT 81.725 170.315 81.900 170.485 ;
        RECT 84.245 170.315 84.415 170.485 ;
        RECT 75.340 170.115 81.900 170.315 ;
        RECT 82.105 170.115 84.415 170.315 ;
        RECT 84.585 170.115 85.760 170.315 ;
        RECT 81.725 169.945 81.900 170.115 ;
        RECT 84.245 169.945 84.415 170.115 ;
        RECT 71.145 168.925 73.175 169.095 ;
        RECT 73.345 168.755 73.515 169.515 ;
        RECT 73.750 169.105 74.265 169.515 ;
        RECT 74.435 168.755 74.725 169.920 ;
        RECT 74.895 169.775 81.555 169.945 ;
        RECT 81.725 169.775 84.075 169.945 ;
        RECT 84.245 169.775 85.755 169.945 ;
        RECT 75.005 168.755 75.175 169.555 ;
        RECT 75.345 168.925 75.675 169.775 ;
        RECT 75.845 168.755 76.015 169.555 ;
        RECT 76.185 168.925 76.515 169.775 ;
        RECT 76.685 168.755 76.855 169.555 ;
        RECT 77.025 168.925 77.355 169.775 ;
        RECT 77.525 168.755 77.695 169.555 ;
        RECT 77.865 168.925 78.195 169.775 ;
        RECT 78.365 168.755 78.535 169.555 ;
        RECT 78.705 168.925 79.035 169.775 ;
        RECT 79.205 168.755 79.375 169.555 ;
        RECT 79.545 168.925 79.875 169.775 ;
        RECT 80.045 168.755 80.215 169.555 ;
        RECT 80.385 168.925 80.715 169.775 ;
        RECT 80.885 168.755 81.055 169.555 ;
        RECT 81.225 168.925 81.555 169.775 ;
        RECT 81.725 168.755 81.895 169.555 ;
        RECT 82.065 168.925 82.395 169.775 ;
        RECT 82.565 168.755 82.735 169.555 ;
        RECT 82.905 168.925 83.235 169.775 ;
        RECT 83.405 168.755 83.575 169.555 ;
        RECT 83.745 168.925 84.075 169.775 ;
        RECT 84.245 168.755 84.415 169.605 ;
        RECT 84.585 168.925 84.915 169.775 ;
        RECT 85.085 168.755 85.255 169.605 ;
        RECT 85.425 168.925 85.755 169.775 ;
        RECT 85.935 169.845 86.685 170.365 ;
        RECT 86.855 170.015 87.605 170.535 ;
        RECT 87.775 170.630 88.035 171.135 ;
        RECT 88.215 170.925 88.545 171.305 ;
        RECT 88.725 170.755 88.895 171.135 ;
        RECT 89.160 170.760 94.505 171.305 ;
        RECT 85.935 168.755 87.605 169.845 ;
        RECT 87.775 169.830 87.945 170.630 ;
        RECT 88.230 170.585 88.895 170.755 ;
        RECT 88.230 170.330 88.400 170.585 ;
        RECT 88.115 170.000 88.400 170.330 ;
        RECT 88.635 170.035 88.965 170.405 ;
        RECT 88.230 169.855 88.400 170.000 ;
        RECT 87.775 168.925 88.045 169.830 ;
        RECT 88.230 169.685 88.895 169.855 ;
        RECT 88.215 168.755 88.545 169.515 ;
        RECT 88.725 168.925 88.895 169.685 ;
        RECT 90.750 169.190 91.100 170.440 ;
        RECT 92.580 169.930 92.920 170.760 ;
        RECT 94.715 170.485 94.945 171.305 ;
        RECT 95.115 170.505 95.445 171.135 ;
        RECT 94.695 170.065 95.025 170.315 ;
        RECT 95.195 169.905 95.445 170.505 ;
        RECT 95.615 170.485 95.825 171.305 ;
        RECT 96.330 170.495 96.575 171.100 ;
        RECT 96.795 170.770 97.305 171.305 ;
        RECT 89.160 168.755 94.505 169.190 ;
        RECT 94.715 168.755 94.945 169.895 ;
        RECT 95.115 168.925 95.445 169.905 ;
        RECT 96.055 170.325 97.285 170.495 ;
        RECT 95.615 168.755 95.825 169.895 ;
        RECT 96.055 169.515 96.395 170.325 ;
        RECT 96.565 169.760 97.315 169.950 ;
        RECT 96.055 169.105 96.570 169.515 ;
        RECT 96.805 168.755 96.975 169.515 ;
        RECT 97.145 169.095 97.315 169.760 ;
        RECT 97.485 169.775 97.675 171.135 ;
        RECT 97.845 170.965 98.120 171.135 ;
        RECT 97.845 170.795 98.125 170.965 ;
        RECT 97.845 169.975 98.120 170.795 ;
        RECT 98.310 170.770 98.840 171.135 ;
        RECT 99.265 170.905 99.595 171.305 ;
        RECT 98.665 170.735 98.840 170.770 ;
        RECT 98.325 169.775 98.495 170.575 ;
        RECT 97.485 169.605 98.495 169.775 ;
        RECT 98.665 170.565 99.595 170.735 ;
        RECT 99.765 170.565 100.020 171.135 ;
        RECT 100.195 170.580 100.485 171.305 ;
        RECT 98.665 169.435 98.835 170.565 ;
        RECT 99.425 170.395 99.595 170.565 ;
        RECT 97.710 169.265 98.835 169.435 ;
        RECT 99.005 170.065 99.200 170.395 ;
        RECT 99.425 170.065 99.680 170.395 ;
        RECT 99.005 169.095 99.175 170.065 ;
        RECT 99.850 169.895 100.020 170.565 ;
        RECT 101.850 170.495 102.095 171.100 ;
        RECT 102.315 170.770 102.825 171.305 ;
        RECT 101.575 170.325 102.805 170.495 ;
        RECT 97.145 168.925 99.175 169.095 ;
        RECT 99.345 168.755 99.515 169.895 ;
        RECT 99.685 168.925 100.020 169.895 ;
        RECT 100.195 168.755 100.485 169.920 ;
        RECT 101.575 169.515 101.915 170.325 ;
        RECT 102.085 169.760 102.835 169.950 ;
        RECT 101.575 169.105 102.090 169.515 ;
        RECT 102.325 168.755 102.495 169.515 ;
        RECT 102.665 169.095 102.835 169.760 ;
        RECT 103.005 169.775 103.195 171.135 ;
        RECT 103.365 170.625 103.640 171.135 ;
        RECT 103.830 170.770 104.360 171.135 ;
        RECT 104.785 170.905 105.115 171.305 ;
        RECT 104.185 170.735 104.360 170.770 ;
        RECT 103.365 170.455 103.645 170.625 ;
        RECT 103.365 169.975 103.640 170.455 ;
        RECT 103.845 169.775 104.015 170.575 ;
        RECT 103.005 169.605 104.015 169.775 ;
        RECT 104.185 170.565 105.115 170.735 ;
        RECT 105.285 170.565 105.540 171.135 ;
        RECT 105.805 170.755 105.975 171.135 ;
        RECT 106.155 170.925 106.485 171.305 ;
        RECT 105.805 170.585 106.470 170.755 ;
        RECT 106.665 170.630 106.925 171.135 ;
        RECT 104.185 169.435 104.355 170.565 ;
        RECT 104.945 170.395 105.115 170.565 ;
        RECT 103.230 169.265 104.355 169.435 ;
        RECT 104.525 170.065 104.720 170.395 ;
        RECT 104.945 170.065 105.200 170.395 ;
        RECT 104.525 169.095 104.695 170.065 ;
        RECT 105.370 169.895 105.540 170.565 ;
        RECT 105.735 170.035 106.065 170.405 ;
        RECT 106.300 170.330 106.470 170.585 ;
        RECT 102.665 168.925 104.695 169.095 ;
        RECT 104.865 168.755 105.035 169.895 ;
        RECT 105.205 168.925 105.540 169.895 ;
        RECT 106.300 170.000 106.585 170.330 ;
        RECT 106.300 169.855 106.470 170.000 ;
        RECT 105.805 169.685 106.470 169.855 ;
        RECT 106.755 169.830 106.925 170.630 ;
        RECT 107.185 170.755 107.355 171.135 ;
        RECT 107.535 170.925 107.865 171.305 ;
        RECT 107.185 170.585 107.850 170.755 ;
        RECT 108.045 170.630 108.305 171.135 ;
        RECT 107.115 170.035 107.445 170.405 ;
        RECT 107.680 170.330 107.850 170.585 ;
        RECT 107.680 170.000 107.965 170.330 ;
        RECT 107.680 169.855 107.850 170.000 ;
        RECT 105.805 168.925 105.975 169.685 ;
        RECT 106.155 168.755 106.485 169.515 ;
        RECT 106.655 168.925 106.925 169.830 ;
        RECT 107.185 169.685 107.850 169.855 ;
        RECT 108.135 169.830 108.305 170.630 ;
        RECT 108.475 170.535 111.985 171.305 ;
        RECT 112.155 170.555 113.365 171.305 ;
        RECT 107.185 168.925 107.355 169.685 ;
        RECT 107.535 168.755 107.865 169.515 ;
        RECT 108.035 168.925 108.305 169.830 ;
        RECT 108.475 169.845 110.165 170.365 ;
        RECT 110.335 170.015 111.985 170.535 ;
        RECT 112.155 169.845 112.675 170.385 ;
        RECT 112.845 170.015 113.365 170.555 ;
        RECT 108.475 168.755 111.985 169.845 ;
        RECT 112.155 168.755 113.365 169.845 ;
        RECT 15.010 168.585 113.450 168.755 ;
        RECT 15.095 167.495 16.305 168.585 ;
        RECT 15.095 166.785 15.615 167.325 ;
        RECT 15.785 166.955 16.305 167.495 ;
        RECT 17.400 167.395 17.655 168.275 ;
        RECT 17.825 167.445 18.130 168.585 ;
        RECT 18.470 168.205 18.800 168.585 ;
        RECT 18.980 168.035 19.150 168.325 ;
        RECT 19.320 168.125 19.570 168.585 ;
        RECT 18.350 167.865 19.150 168.035 ;
        RECT 19.740 168.075 20.610 168.415 ;
        RECT 15.095 166.035 16.305 166.785 ;
        RECT 17.400 166.745 17.610 167.395 ;
        RECT 18.350 167.275 18.520 167.865 ;
        RECT 19.740 167.695 19.910 168.075 ;
        RECT 20.845 167.955 21.015 168.415 ;
        RECT 21.185 168.125 21.555 168.585 ;
        RECT 21.850 167.985 22.020 168.325 ;
        RECT 22.190 168.155 22.520 168.585 ;
        RECT 22.755 167.985 22.925 168.325 ;
        RECT 18.690 167.525 19.910 167.695 ;
        RECT 20.080 167.615 20.540 167.905 ;
        RECT 20.845 167.785 21.405 167.955 ;
        RECT 21.850 167.815 22.925 167.985 ;
        RECT 23.095 168.085 23.775 168.415 ;
        RECT 23.990 168.085 24.240 168.415 ;
        RECT 24.410 168.125 24.660 168.585 ;
        RECT 21.235 167.645 21.405 167.785 ;
        RECT 20.080 167.605 21.045 167.615 ;
        RECT 19.740 167.435 19.910 167.525 ;
        RECT 20.370 167.445 21.045 167.605 ;
        RECT 17.780 167.245 18.520 167.275 ;
        RECT 17.780 166.945 18.695 167.245 ;
        RECT 18.370 166.770 18.695 166.945 ;
        RECT 17.400 166.215 17.655 166.745 ;
        RECT 17.825 166.035 18.130 166.495 ;
        RECT 18.375 166.415 18.695 166.770 ;
        RECT 18.865 166.985 19.405 167.355 ;
        RECT 19.740 167.265 20.145 167.435 ;
        RECT 18.865 166.585 19.105 166.985 ;
        RECT 19.585 166.815 19.805 167.095 ;
        RECT 19.275 166.645 19.805 166.815 ;
        RECT 19.275 166.415 19.445 166.645 ;
        RECT 19.975 166.485 20.145 167.265 ;
        RECT 20.315 166.655 20.665 167.275 ;
        RECT 20.835 166.655 21.045 167.445 ;
        RECT 21.235 167.475 22.735 167.645 ;
        RECT 21.235 166.785 21.405 167.475 ;
        RECT 23.095 167.305 23.265 168.085 ;
        RECT 24.070 167.955 24.240 168.085 ;
        RECT 21.575 167.135 23.265 167.305 ;
        RECT 23.435 167.525 23.900 167.915 ;
        RECT 24.070 167.785 24.465 167.955 ;
        RECT 21.575 166.955 21.745 167.135 ;
        RECT 18.375 166.245 19.445 166.415 ;
        RECT 19.615 166.035 19.805 166.475 ;
        RECT 19.975 166.205 20.925 166.485 ;
        RECT 21.235 166.395 21.495 166.785 ;
        RECT 21.915 166.715 22.705 166.965 ;
        RECT 21.145 166.225 21.495 166.395 ;
        RECT 21.705 166.035 22.035 166.495 ;
        RECT 22.910 166.425 23.080 167.135 ;
        RECT 23.435 166.935 23.605 167.525 ;
        RECT 23.250 166.715 23.605 166.935 ;
        RECT 23.775 166.715 24.125 167.335 ;
        RECT 24.295 166.425 24.465 167.785 ;
        RECT 24.830 167.615 25.155 168.400 ;
        RECT 24.635 166.565 25.095 167.615 ;
        RECT 22.910 166.255 23.765 166.425 ;
        RECT 23.970 166.255 24.465 166.425 ;
        RECT 24.635 166.035 24.965 166.395 ;
        RECT 25.325 166.295 25.495 168.415 ;
        RECT 25.665 168.085 25.995 168.585 ;
        RECT 26.165 167.915 26.420 168.415 ;
        RECT 25.670 167.745 26.420 167.915 ;
        RECT 25.670 166.755 25.900 167.745 ;
        RECT 26.070 166.925 26.420 167.575 ;
        RECT 26.600 167.395 26.855 168.275 ;
        RECT 27.025 167.445 27.330 168.585 ;
        RECT 27.670 168.205 28.000 168.585 ;
        RECT 28.180 168.035 28.350 168.325 ;
        RECT 28.520 168.125 28.770 168.585 ;
        RECT 27.550 167.865 28.350 168.035 ;
        RECT 28.940 168.075 29.810 168.415 ;
        RECT 25.670 166.585 26.420 166.755 ;
        RECT 25.665 166.035 25.995 166.415 ;
        RECT 26.165 166.295 26.420 166.585 ;
        RECT 26.600 166.745 26.810 167.395 ;
        RECT 27.550 167.275 27.720 167.865 ;
        RECT 28.940 167.695 29.110 168.075 ;
        RECT 30.045 167.955 30.215 168.415 ;
        RECT 30.385 168.125 30.755 168.585 ;
        RECT 31.050 167.985 31.220 168.325 ;
        RECT 31.390 168.155 31.720 168.585 ;
        RECT 31.955 167.985 32.125 168.325 ;
        RECT 27.890 167.525 29.110 167.695 ;
        RECT 29.280 167.615 29.740 167.905 ;
        RECT 30.045 167.785 30.605 167.955 ;
        RECT 31.050 167.815 32.125 167.985 ;
        RECT 32.295 168.085 32.975 168.415 ;
        RECT 33.190 168.085 33.440 168.415 ;
        RECT 33.610 168.125 33.860 168.585 ;
        RECT 30.435 167.645 30.605 167.785 ;
        RECT 29.280 167.605 30.245 167.615 ;
        RECT 28.940 167.435 29.110 167.525 ;
        RECT 29.570 167.445 30.245 167.605 ;
        RECT 26.980 167.245 27.720 167.275 ;
        RECT 26.980 166.945 27.895 167.245 ;
        RECT 27.570 166.770 27.895 166.945 ;
        RECT 26.600 166.215 26.855 166.745 ;
        RECT 27.025 166.035 27.330 166.495 ;
        RECT 27.575 166.415 27.895 166.770 ;
        RECT 28.065 166.985 28.605 167.355 ;
        RECT 28.940 167.265 29.345 167.435 ;
        RECT 28.065 166.585 28.305 166.985 ;
        RECT 28.785 166.815 29.005 167.095 ;
        RECT 28.475 166.645 29.005 166.815 ;
        RECT 28.475 166.415 28.645 166.645 ;
        RECT 29.175 166.485 29.345 167.265 ;
        RECT 29.515 166.655 29.865 167.275 ;
        RECT 30.035 166.655 30.245 167.445 ;
        RECT 30.435 167.475 31.935 167.645 ;
        RECT 30.435 166.785 30.605 167.475 ;
        RECT 32.295 167.305 32.465 168.085 ;
        RECT 33.270 167.955 33.440 168.085 ;
        RECT 30.775 167.135 32.465 167.305 ;
        RECT 32.635 167.525 33.100 167.915 ;
        RECT 33.270 167.785 33.665 167.955 ;
        RECT 30.775 166.955 30.945 167.135 ;
        RECT 27.575 166.245 28.645 166.415 ;
        RECT 28.815 166.035 29.005 166.475 ;
        RECT 29.175 166.205 30.125 166.485 ;
        RECT 30.435 166.395 30.695 166.785 ;
        RECT 31.115 166.715 31.905 166.965 ;
        RECT 30.345 166.225 30.695 166.395 ;
        RECT 30.905 166.035 31.235 166.495 ;
        RECT 32.110 166.425 32.280 167.135 ;
        RECT 32.635 166.935 32.805 167.525 ;
        RECT 32.450 166.715 32.805 166.935 ;
        RECT 32.975 166.715 33.325 167.335 ;
        RECT 33.495 166.425 33.665 167.785 ;
        RECT 34.030 167.615 34.355 168.400 ;
        RECT 33.835 166.565 34.295 167.615 ;
        RECT 32.110 166.255 32.965 166.425 ;
        RECT 33.170 166.255 33.665 166.425 ;
        RECT 33.835 166.035 34.165 166.395 ;
        RECT 34.525 166.295 34.695 168.415 ;
        RECT 34.865 168.085 35.195 168.585 ;
        RECT 35.365 167.915 35.620 168.415 ;
        RECT 34.870 167.745 35.620 167.915 ;
        RECT 34.870 166.755 35.100 167.745 ;
        RECT 35.270 166.925 35.620 167.575 ;
        RECT 35.795 167.420 36.085 168.585 ;
        RECT 36.255 167.750 36.640 168.585 ;
        RECT 36.810 167.580 37.070 168.385 ;
        RECT 37.240 167.750 37.500 168.585 ;
        RECT 37.670 167.580 37.925 168.385 ;
        RECT 38.100 167.750 38.360 168.585 ;
        RECT 38.530 167.580 38.785 168.385 ;
        RECT 38.960 167.750 39.305 168.585 ;
        RECT 39.590 167.955 39.875 168.415 ;
        RECT 40.045 168.125 40.315 168.585 ;
        RECT 39.590 167.735 40.545 167.955 ;
        RECT 36.255 167.410 39.285 167.580 ;
        RECT 36.255 166.845 36.555 167.410 ;
        RECT 36.730 167.015 38.945 167.240 ;
        RECT 39.115 166.845 39.285 167.410 ;
        RECT 39.475 167.005 40.165 167.565 ;
        RECT 34.870 166.585 35.620 166.755 ;
        RECT 34.865 166.035 35.195 166.415 ;
        RECT 35.365 166.295 35.620 166.585 ;
        RECT 35.795 166.035 36.085 166.760 ;
        RECT 36.255 166.675 39.285 166.845 ;
        RECT 40.335 166.835 40.545 167.735 ;
        RECT 36.775 166.035 37.075 166.505 ;
        RECT 37.245 166.230 37.500 166.675 ;
        RECT 37.670 166.035 37.930 166.505 ;
        RECT 38.100 166.230 38.360 166.675 ;
        RECT 39.590 166.665 40.545 166.835 ;
        RECT 40.715 167.565 41.115 168.415 ;
        RECT 41.305 167.955 41.585 168.415 ;
        RECT 42.105 168.125 42.430 168.585 ;
        RECT 41.305 167.735 42.430 167.955 ;
        RECT 40.715 167.005 41.810 167.565 ;
        RECT 41.980 167.275 42.430 167.735 ;
        RECT 42.600 167.445 42.985 168.415 ;
        RECT 43.215 167.445 43.425 168.585 ;
        RECT 38.530 166.035 38.825 166.505 ;
        RECT 39.590 166.205 39.875 166.665 ;
        RECT 40.045 166.035 40.315 166.495 ;
        RECT 40.715 166.205 41.115 167.005 ;
        RECT 41.980 166.945 42.535 167.275 ;
        RECT 41.980 166.835 42.430 166.945 ;
        RECT 41.305 166.665 42.430 166.835 ;
        RECT 42.705 166.775 42.985 167.445 ;
        RECT 43.595 167.435 43.925 168.415 ;
        RECT 44.095 167.445 44.325 168.585 ;
        RECT 44.545 167.775 44.840 168.585 ;
        RECT 41.305 166.205 41.585 166.665 ;
        RECT 42.105 166.035 42.430 166.495 ;
        RECT 42.600 166.205 42.985 166.775 ;
        RECT 43.215 166.035 43.425 166.855 ;
        RECT 43.595 166.835 43.845 167.435 ;
        RECT 45.020 167.275 45.265 168.415 ;
        RECT 45.440 167.775 45.700 168.585 ;
        RECT 46.300 168.580 52.575 168.585 ;
        RECT 45.880 167.275 46.130 168.410 ;
        RECT 46.300 167.785 46.560 168.580 ;
        RECT 46.730 167.685 46.990 168.410 ;
        RECT 47.160 167.855 47.420 168.580 ;
        RECT 47.590 167.685 47.850 168.410 ;
        RECT 48.020 167.855 48.280 168.580 ;
        RECT 48.450 167.685 48.710 168.410 ;
        RECT 48.880 167.855 49.140 168.580 ;
        RECT 49.310 167.685 49.570 168.410 ;
        RECT 49.740 167.855 49.985 168.580 ;
        RECT 50.155 167.685 50.415 168.410 ;
        RECT 50.600 167.855 50.845 168.580 ;
        RECT 51.015 167.685 51.275 168.410 ;
        RECT 51.460 167.855 51.705 168.580 ;
        RECT 51.875 167.685 52.135 168.410 ;
        RECT 52.320 167.855 52.575 168.580 ;
        RECT 46.730 167.670 52.135 167.685 ;
        RECT 52.745 167.670 53.035 168.410 ;
        RECT 53.205 167.840 53.475 168.585 ;
        RECT 46.730 167.565 53.475 167.670 ;
        RECT 46.730 167.445 53.505 167.565 ;
        RECT 52.310 167.395 53.505 167.445 ;
        RECT 53.885 167.435 54.215 168.585 ;
        RECT 54.385 167.565 54.555 168.415 ;
        RECT 54.725 167.785 55.055 168.585 ;
        RECT 55.225 167.565 55.395 168.415 ;
        RECT 55.575 167.785 55.815 168.585 ;
        RECT 55.985 167.605 56.315 168.415 ;
        RECT 54.385 167.395 55.395 167.565 ;
        RECT 55.600 167.435 56.315 167.605 ;
        RECT 56.535 167.445 56.765 168.585 ;
        RECT 56.935 167.435 57.265 168.415 ;
        RECT 57.435 167.445 57.645 168.585 ;
        RECT 58.850 167.715 59.135 168.585 ;
        RECT 59.305 167.955 59.565 168.415 ;
        RECT 59.740 168.125 59.995 168.585 ;
        RECT 60.165 167.955 60.425 168.415 ;
        RECT 59.305 167.785 60.425 167.955 ;
        RECT 60.595 167.785 60.905 168.585 ;
        RECT 59.305 167.535 59.565 167.785 ;
        RECT 61.075 167.615 61.385 168.415 ;
        RECT 44.015 167.025 44.345 167.275 ;
        RECT 43.595 166.205 43.925 166.835 ;
        RECT 44.095 166.035 44.325 166.855 ;
        RECT 44.535 166.715 44.850 167.275 ;
        RECT 45.020 167.025 52.140 167.275 ;
        RECT 44.535 166.035 44.840 166.545 ;
        RECT 45.020 166.215 45.270 167.025 ;
        RECT 45.440 166.035 45.700 166.560 ;
        RECT 45.880 166.215 46.130 167.025 ;
        RECT 52.310 166.855 53.475 167.395 ;
        RECT 46.730 166.685 53.475 166.855 ;
        RECT 54.385 167.225 54.880 167.395 ;
        RECT 54.385 167.055 54.885 167.225 ;
        RECT 55.600 167.195 55.770 167.435 ;
        RECT 54.385 166.855 54.880 167.055 ;
        RECT 55.270 167.025 55.770 167.195 ;
        RECT 55.940 167.025 56.320 167.265 ;
        RECT 56.515 167.025 56.845 167.275 ;
        RECT 55.600 166.855 55.770 167.025 ;
        RECT 46.300 166.035 46.560 166.595 ;
        RECT 46.730 166.230 46.990 166.685 ;
        RECT 47.160 166.035 47.420 166.515 ;
        RECT 47.590 166.230 47.850 166.685 ;
        RECT 48.020 166.035 48.280 166.515 ;
        RECT 48.450 166.230 48.710 166.685 ;
        RECT 48.880 166.035 49.125 166.515 ;
        RECT 49.295 166.230 49.570 166.685 ;
        RECT 49.740 166.035 49.985 166.515 ;
        RECT 50.155 166.230 50.415 166.685 ;
        RECT 50.595 166.035 50.845 166.515 ;
        RECT 51.015 166.230 51.275 166.685 ;
        RECT 51.455 166.035 51.705 166.515 ;
        RECT 51.875 166.230 52.135 166.685 ;
        RECT 52.315 166.035 52.575 166.515 ;
        RECT 52.745 166.230 53.005 166.685 ;
        RECT 53.175 166.035 53.475 166.515 ;
        RECT 53.885 166.035 54.215 166.835 ;
        RECT 54.385 166.685 55.395 166.855 ;
        RECT 55.600 166.685 56.235 166.855 ;
        RECT 54.385 166.205 54.555 166.685 ;
        RECT 54.725 166.035 55.055 166.515 ;
        RECT 55.225 166.205 55.395 166.685 ;
        RECT 55.645 166.035 55.885 166.515 ;
        RECT 56.065 166.205 56.235 166.685 ;
        RECT 56.535 166.035 56.765 166.855 ;
        RECT 57.015 166.835 57.265 167.435 ;
        RECT 58.810 167.365 59.565 167.535 ;
        RECT 60.355 167.445 61.385 167.615 ;
        RECT 58.810 166.855 59.215 167.365 ;
        RECT 60.355 167.195 60.525 167.445 ;
        RECT 59.385 167.025 60.525 167.195 ;
        RECT 56.935 166.205 57.265 166.835 ;
        RECT 57.435 166.035 57.645 166.855 ;
        RECT 58.810 166.685 60.460 166.855 ;
        RECT 60.695 166.705 61.045 167.275 ;
        RECT 58.855 166.035 59.135 166.515 ;
        RECT 59.305 166.295 59.565 166.685 ;
        RECT 59.740 166.035 59.995 166.515 ;
        RECT 60.165 166.295 60.460 166.685 ;
        RECT 61.215 166.535 61.385 167.445 ;
        RECT 61.555 167.420 61.845 168.585 ;
        RECT 62.015 167.495 63.685 168.585 ;
        RECT 63.855 167.995 64.555 168.415 ;
        RECT 64.755 168.225 65.085 168.585 ;
        RECT 65.255 167.995 65.585 168.395 ;
        RECT 63.855 167.765 65.585 167.995 ;
        RECT 62.015 166.975 62.765 167.495 ;
        RECT 62.935 166.805 63.685 167.325 ;
        RECT 60.640 166.035 60.915 166.515 ;
        RECT 61.085 166.205 61.385 166.535 ;
        RECT 61.555 166.035 61.845 166.760 ;
        RECT 62.015 166.035 63.685 166.805 ;
        RECT 63.855 166.795 64.060 167.765 ;
        RECT 64.230 167.025 64.560 167.565 ;
        RECT 64.735 167.275 65.060 167.565 ;
        RECT 65.255 167.545 65.585 167.765 ;
        RECT 65.755 167.275 65.925 168.245 ;
        RECT 66.105 167.525 66.435 168.585 ;
        RECT 66.615 167.495 68.285 168.585 ;
        RECT 68.830 167.605 69.085 168.275 ;
        RECT 69.265 167.785 69.550 168.585 ;
        RECT 69.730 167.865 70.060 168.375 ;
        RECT 64.735 166.945 65.230 167.275 ;
        RECT 65.550 166.945 65.925 167.275 ;
        RECT 66.135 166.945 66.445 167.275 ;
        RECT 66.615 166.975 67.365 167.495 ;
        RECT 67.535 166.805 68.285 167.325 ;
        RECT 68.830 167.225 69.010 167.605 ;
        RECT 69.730 167.275 69.980 167.865 ;
        RECT 70.330 167.715 70.500 168.325 ;
        RECT 70.670 167.895 71.000 168.585 ;
        RECT 71.230 168.035 71.470 168.325 ;
        RECT 71.670 168.205 72.090 168.585 ;
        RECT 72.270 168.115 72.900 168.365 ;
        RECT 73.370 168.205 73.700 168.585 ;
        RECT 72.270 168.035 72.440 168.115 ;
        RECT 73.870 168.035 74.040 168.325 ;
        RECT 74.220 168.205 74.600 168.585 ;
        RECT 74.840 168.200 75.670 168.370 ;
        RECT 71.230 167.865 72.440 168.035 ;
        RECT 68.745 167.055 69.010 167.225 ;
        RECT 63.855 166.205 64.565 166.795 ;
        RECT 65.075 166.565 66.435 166.775 ;
        RECT 65.075 166.205 65.405 166.565 ;
        RECT 65.605 166.035 65.935 166.395 ;
        RECT 66.105 166.205 66.435 166.565 ;
        RECT 66.615 166.035 68.285 166.805 ;
        RECT 68.830 166.745 69.010 167.055 ;
        RECT 69.180 166.945 69.980 167.275 ;
        RECT 68.830 166.215 69.085 166.745 ;
        RECT 69.265 166.035 69.550 166.495 ;
        RECT 69.730 166.295 69.980 166.945 ;
        RECT 70.180 167.695 70.500 167.715 ;
        RECT 70.180 167.525 72.100 167.695 ;
        RECT 70.180 166.630 70.370 167.525 ;
        RECT 72.270 167.355 72.440 167.865 ;
        RECT 72.610 167.605 73.130 167.915 ;
        RECT 70.540 167.185 72.440 167.355 ;
        RECT 70.540 167.125 70.870 167.185 ;
        RECT 71.020 166.955 71.350 167.015 ;
        RECT 70.690 166.685 71.350 166.955 ;
        RECT 70.180 166.300 70.500 166.630 ;
        RECT 70.680 166.035 71.340 166.515 ;
        RECT 71.540 166.425 71.710 167.185 ;
        RECT 72.610 167.015 72.790 167.425 ;
        RECT 71.880 166.845 72.210 166.965 ;
        RECT 72.960 166.845 73.130 167.605 ;
        RECT 71.880 166.675 73.130 166.845 ;
        RECT 73.300 167.785 74.670 168.035 ;
        RECT 73.300 167.015 73.490 167.785 ;
        RECT 74.420 167.525 74.670 167.785 ;
        RECT 73.660 167.355 73.910 167.515 ;
        RECT 74.840 167.355 75.010 168.200 ;
        RECT 75.905 167.915 76.075 168.415 ;
        RECT 76.245 168.085 76.575 168.585 ;
        RECT 75.180 167.525 75.680 167.905 ;
        RECT 75.905 167.745 76.600 167.915 ;
        RECT 73.660 167.185 75.010 167.355 ;
        RECT 74.590 167.145 75.010 167.185 ;
        RECT 73.300 166.675 73.720 167.015 ;
        RECT 74.010 166.685 74.420 167.015 ;
        RECT 71.540 166.255 72.390 166.425 ;
        RECT 72.950 166.035 73.270 166.495 ;
        RECT 73.470 166.245 73.720 166.675 ;
        RECT 74.010 166.035 74.420 166.475 ;
        RECT 74.590 166.415 74.760 167.145 ;
        RECT 74.930 166.595 75.280 166.965 ;
        RECT 75.460 166.655 75.680 167.525 ;
        RECT 75.850 166.955 76.260 167.575 ;
        RECT 76.430 166.775 76.600 167.745 ;
        RECT 75.905 166.585 76.600 166.775 ;
        RECT 74.590 166.215 75.605 166.415 ;
        RECT 75.905 166.255 76.075 166.585 ;
        RECT 76.245 166.035 76.575 166.415 ;
        RECT 76.790 166.295 77.015 168.415 ;
        RECT 77.185 168.085 77.515 168.585 ;
        RECT 77.685 167.915 77.855 168.415 ;
        RECT 77.190 167.745 77.855 167.915 ;
        RECT 78.125 167.775 78.420 168.585 ;
        RECT 77.190 166.755 77.420 167.745 ;
        RECT 77.590 166.925 77.940 167.575 ;
        RECT 78.600 167.275 78.845 168.415 ;
        RECT 79.020 167.775 79.280 168.585 ;
        RECT 79.880 168.580 86.155 168.585 ;
        RECT 79.460 167.275 79.710 168.410 ;
        RECT 79.880 167.785 80.140 168.580 ;
        RECT 80.310 167.685 80.570 168.410 ;
        RECT 80.740 167.855 81.000 168.580 ;
        RECT 81.170 167.685 81.430 168.410 ;
        RECT 81.600 167.855 81.860 168.580 ;
        RECT 82.030 167.685 82.290 168.410 ;
        RECT 82.460 167.855 82.720 168.580 ;
        RECT 82.890 167.685 83.150 168.410 ;
        RECT 83.320 167.855 83.565 168.580 ;
        RECT 83.735 167.685 83.995 168.410 ;
        RECT 84.180 167.855 84.425 168.580 ;
        RECT 84.595 167.685 84.855 168.410 ;
        RECT 85.040 167.855 85.285 168.580 ;
        RECT 85.455 167.685 85.715 168.410 ;
        RECT 85.900 167.855 86.155 168.580 ;
        RECT 80.310 167.670 85.715 167.685 ;
        RECT 86.325 167.670 86.615 168.410 ;
        RECT 86.785 167.840 87.055 168.585 ;
        RECT 80.310 167.445 87.055 167.670 ;
        RECT 77.190 166.585 77.855 166.755 ;
        RECT 78.115 166.715 78.430 167.275 ;
        RECT 78.600 167.025 85.720 167.275 ;
        RECT 77.185 166.035 77.515 166.415 ;
        RECT 77.685 166.295 77.855 166.585 ;
        RECT 78.115 166.035 78.420 166.545 ;
        RECT 78.600 166.215 78.850 167.025 ;
        RECT 79.020 166.035 79.280 166.560 ;
        RECT 79.460 166.215 79.710 167.025 ;
        RECT 85.890 166.855 87.055 167.445 ;
        RECT 87.315 167.420 87.605 168.585 ;
        RECT 87.775 167.510 88.045 168.415 ;
        RECT 88.215 167.825 88.545 168.585 ;
        RECT 88.725 167.655 88.895 168.415 ;
        RECT 80.310 166.685 87.055 166.855 ;
        RECT 79.880 166.035 80.140 166.595 ;
        RECT 80.310 166.230 80.570 166.685 ;
        RECT 80.740 166.035 81.000 166.515 ;
        RECT 81.170 166.230 81.430 166.685 ;
        RECT 81.600 166.035 81.860 166.515 ;
        RECT 82.030 166.230 82.290 166.685 ;
        RECT 82.460 166.035 82.705 166.515 ;
        RECT 82.875 166.230 83.150 166.685 ;
        RECT 83.320 166.035 83.565 166.515 ;
        RECT 83.735 166.230 83.995 166.685 ;
        RECT 84.175 166.035 84.425 166.515 ;
        RECT 84.595 166.230 84.855 166.685 ;
        RECT 85.035 166.035 85.285 166.515 ;
        RECT 85.455 166.230 85.715 166.685 ;
        RECT 85.895 166.035 86.155 166.515 ;
        RECT 86.325 166.230 86.585 166.685 ;
        RECT 86.755 166.035 87.055 166.515 ;
        RECT 87.315 166.035 87.605 166.760 ;
        RECT 87.775 166.710 87.945 167.510 ;
        RECT 88.230 167.485 88.895 167.655 ;
        RECT 88.230 167.340 88.400 167.485 ;
        RECT 89.195 167.445 89.425 168.585 ;
        RECT 89.595 167.435 89.925 168.415 ;
        RECT 90.095 167.445 90.305 168.585 ;
        RECT 91.085 167.655 91.255 168.415 ;
        RECT 91.435 167.825 91.765 168.585 ;
        RECT 91.085 167.485 91.750 167.655 ;
        RECT 91.935 167.510 92.205 168.415 ;
        RECT 88.115 167.010 88.400 167.340 ;
        RECT 88.230 166.755 88.400 167.010 ;
        RECT 88.635 166.935 88.965 167.305 ;
        RECT 89.175 167.025 89.505 167.275 ;
        RECT 87.775 166.205 88.035 166.710 ;
        RECT 88.230 166.585 88.895 166.755 ;
        RECT 88.215 166.035 88.545 166.415 ;
        RECT 88.725 166.205 88.895 166.585 ;
        RECT 89.195 166.035 89.425 166.855 ;
        RECT 89.675 166.835 89.925 167.435 ;
        RECT 91.580 167.340 91.750 167.485 ;
        RECT 91.015 166.935 91.345 167.305 ;
        RECT 91.580 167.010 91.865 167.340 ;
        RECT 89.595 166.205 89.925 166.835 ;
        RECT 90.095 166.035 90.305 166.855 ;
        RECT 91.580 166.755 91.750 167.010 ;
        RECT 91.085 166.585 91.750 166.755 ;
        RECT 92.035 166.710 92.205 167.510 ;
        RECT 91.085 166.205 91.255 166.585 ;
        RECT 91.435 166.035 91.765 166.415 ;
        RECT 91.945 166.205 92.205 166.710 ;
        RECT 92.380 167.395 92.635 168.275 ;
        RECT 92.805 167.445 93.110 168.585 ;
        RECT 93.450 168.205 93.780 168.585 ;
        RECT 93.960 168.035 94.130 168.325 ;
        RECT 94.300 168.125 94.550 168.585 ;
        RECT 93.330 167.865 94.130 168.035 ;
        RECT 94.720 168.075 95.590 168.415 ;
        RECT 92.380 166.745 92.590 167.395 ;
        RECT 93.330 167.275 93.500 167.865 ;
        RECT 94.720 167.695 94.890 168.075 ;
        RECT 95.825 167.955 95.995 168.415 ;
        RECT 96.165 168.125 96.535 168.585 ;
        RECT 96.830 167.985 97.000 168.325 ;
        RECT 97.170 168.155 97.500 168.585 ;
        RECT 97.735 167.985 97.905 168.325 ;
        RECT 93.670 167.525 94.890 167.695 ;
        RECT 95.060 167.615 95.520 167.905 ;
        RECT 95.825 167.785 96.385 167.955 ;
        RECT 96.830 167.815 97.905 167.985 ;
        RECT 98.075 168.085 98.755 168.415 ;
        RECT 98.970 168.085 99.220 168.415 ;
        RECT 99.390 168.125 99.640 168.585 ;
        RECT 96.215 167.645 96.385 167.785 ;
        RECT 95.060 167.605 96.025 167.615 ;
        RECT 94.720 167.435 94.890 167.525 ;
        RECT 95.350 167.445 96.025 167.605 ;
        RECT 92.760 167.245 93.500 167.275 ;
        RECT 92.760 166.945 93.675 167.245 ;
        RECT 93.350 166.770 93.675 166.945 ;
        RECT 92.380 166.215 92.635 166.745 ;
        RECT 92.805 166.035 93.110 166.495 ;
        RECT 93.355 166.415 93.675 166.770 ;
        RECT 93.845 166.985 94.385 167.355 ;
        RECT 94.720 167.265 95.125 167.435 ;
        RECT 93.845 166.585 94.085 166.985 ;
        RECT 94.565 166.815 94.785 167.095 ;
        RECT 94.255 166.645 94.785 166.815 ;
        RECT 94.255 166.415 94.425 166.645 ;
        RECT 94.955 166.485 95.125 167.265 ;
        RECT 95.295 166.655 95.645 167.275 ;
        RECT 95.815 166.655 96.025 167.445 ;
        RECT 96.215 167.475 97.715 167.645 ;
        RECT 96.215 166.785 96.385 167.475 ;
        RECT 98.075 167.305 98.245 168.085 ;
        RECT 99.050 167.955 99.220 168.085 ;
        RECT 96.555 167.135 98.245 167.305 ;
        RECT 98.415 167.525 98.880 167.915 ;
        RECT 99.050 167.785 99.445 167.955 ;
        RECT 96.555 166.955 96.725 167.135 ;
        RECT 93.355 166.245 94.425 166.415 ;
        RECT 94.595 166.035 94.785 166.475 ;
        RECT 94.955 166.205 95.905 166.485 ;
        RECT 96.215 166.395 96.475 166.785 ;
        RECT 96.895 166.715 97.685 166.965 ;
        RECT 96.125 166.225 96.475 166.395 ;
        RECT 96.685 166.035 97.015 166.495 ;
        RECT 97.890 166.425 98.060 167.135 ;
        RECT 98.415 166.935 98.585 167.525 ;
        RECT 98.230 166.715 98.585 166.935 ;
        RECT 98.755 166.715 99.105 167.335 ;
        RECT 99.275 166.425 99.445 167.785 ;
        RECT 99.810 167.615 100.135 168.400 ;
        RECT 99.615 166.565 100.075 167.615 ;
        RECT 97.890 166.255 98.745 166.425 ;
        RECT 98.950 166.255 99.445 166.425 ;
        RECT 99.615 166.035 99.945 166.395 ;
        RECT 100.305 166.295 100.475 168.415 ;
        RECT 100.645 168.085 100.975 168.585 ;
        RECT 101.145 167.915 101.400 168.415 ;
        RECT 100.650 167.745 101.400 167.915 ;
        RECT 101.690 167.955 101.975 168.415 ;
        RECT 102.145 168.125 102.415 168.585 ;
        RECT 100.650 166.755 100.880 167.745 ;
        RECT 101.690 167.735 102.645 167.955 ;
        RECT 101.050 166.925 101.400 167.575 ;
        RECT 101.575 167.005 102.265 167.565 ;
        RECT 102.435 166.835 102.645 167.735 ;
        RECT 100.650 166.585 101.400 166.755 ;
        RECT 100.645 166.035 100.975 166.415 ;
        RECT 101.145 166.295 101.400 166.585 ;
        RECT 101.690 166.665 102.645 166.835 ;
        RECT 102.815 167.565 103.215 168.415 ;
        RECT 103.405 167.955 103.685 168.415 ;
        RECT 104.205 168.125 104.530 168.585 ;
        RECT 103.405 167.735 104.530 167.955 ;
        RECT 102.815 167.005 103.910 167.565 ;
        RECT 104.080 167.275 104.530 167.735 ;
        RECT 104.700 167.445 105.085 168.415 ;
        RECT 101.690 166.205 101.975 166.665 ;
        RECT 102.145 166.035 102.415 166.495 ;
        RECT 102.815 166.205 103.215 167.005 ;
        RECT 104.080 166.945 104.635 167.275 ;
        RECT 104.080 166.835 104.530 166.945 ;
        RECT 103.405 166.665 104.530 166.835 ;
        RECT 104.805 166.775 105.085 167.445 ;
        RECT 105.255 167.495 106.465 168.585 ;
        RECT 106.725 167.655 106.895 168.415 ;
        RECT 107.075 167.825 107.405 168.585 ;
        RECT 105.255 166.955 105.775 167.495 ;
        RECT 106.725 167.485 107.390 167.655 ;
        RECT 107.575 167.510 107.845 168.415 ;
        RECT 108.020 168.160 108.355 168.585 ;
        RECT 108.525 167.980 108.710 168.385 ;
        RECT 107.220 167.340 107.390 167.485 ;
        RECT 105.945 166.785 106.465 167.325 ;
        RECT 106.655 166.935 106.985 167.305 ;
        RECT 107.220 167.010 107.505 167.340 ;
        RECT 103.405 166.205 103.685 166.665 ;
        RECT 104.205 166.035 104.530 166.495 ;
        RECT 104.700 166.205 105.085 166.775 ;
        RECT 105.255 166.035 106.465 166.785 ;
        RECT 107.220 166.755 107.390 167.010 ;
        RECT 106.725 166.585 107.390 166.755 ;
        RECT 107.675 166.710 107.845 167.510 ;
        RECT 106.725 166.205 106.895 166.585 ;
        RECT 107.075 166.035 107.405 166.415 ;
        RECT 107.585 166.205 107.845 166.710 ;
        RECT 108.045 167.805 108.710 167.980 ;
        RECT 108.915 167.805 109.245 168.585 ;
        RECT 108.045 166.775 108.385 167.805 ;
        RECT 109.415 167.615 109.685 168.385 ;
        RECT 108.555 167.445 109.685 167.615 ;
        RECT 108.555 166.945 108.805 167.445 ;
        RECT 108.045 166.605 108.730 166.775 ;
        RECT 108.985 166.695 109.345 167.275 ;
        RECT 108.020 166.035 108.355 166.435 ;
        RECT 108.525 166.205 108.730 166.605 ;
        RECT 109.515 166.535 109.685 167.445 ;
        RECT 110.315 167.495 111.985 168.585 ;
        RECT 112.155 167.495 113.365 168.585 ;
        RECT 110.315 166.975 111.065 167.495 ;
        RECT 111.235 166.805 111.985 167.325 ;
        RECT 112.155 166.955 112.675 167.495 ;
        RECT 108.940 166.035 109.215 166.515 ;
        RECT 109.425 166.205 109.685 166.535 ;
        RECT 110.315 166.035 111.985 166.805 ;
        RECT 112.845 166.785 113.365 167.325 ;
        RECT 112.155 166.035 113.365 166.785 ;
        RECT 15.010 165.865 113.450 166.035 ;
        RECT 15.095 165.115 16.305 165.865 ;
        RECT 15.095 164.575 15.615 165.115 ;
        RECT 17.455 165.045 17.665 165.865 ;
        RECT 17.835 165.065 18.165 165.695 ;
        RECT 15.785 164.405 16.305 164.945 ;
        RECT 17.835 164.465 18.085 165.065 ;
        RECT 18.335 165.045 18.565 165.865 ;
        RECT 19.050 165.055 19.295 165.660 ;
        RECT 19.515 165.330 20.025 165.865 ;
        RECT 18.775 164.885 20.005 165.055 ;
        RECT 18.255 164.625 18.585 164.875 ;
        RECT 15.095 163.315 16.305 164.405 ;
        RECT 17.455 163.315 17.665 164.455 ;
        RECT 17.835 163.485 18.165 164.465 ;
        RECT 18.335 163.315 18.565 164.455 ;
        RECT 18.775 164.075 19.115 164.885 ;
        RECT 19.285 164.320 20.035 164.510 ;
        RECT 18.775 163.665 19.290 164.075 ;
        RECT 19.525 163.315 19.695 164.075 ;
        RECT 19.865 163.655 20.035 164.320 ;
        RECT 20.205 164.335 20.395 165.695 ;
        RECT 20.565 164.845 20.840 165.695 ;
        RECT 21.030 165.330 21.560 165.695 ;
        RECT 21.985 165.465 22.315 165.865 ;
        RECT 21.385 165.295 21.560 165.330 ;
        RECT 20.565 164.675 20.845 164.845 ;
        RECT 20.565 164.535 20.840 164.675 ;
        RECT 21.045 164.335 21.215 165.135 ;
        RECT 20.205 164.165 21.215 164.335 ;
        RECT 21.385 165.125 22.315 165.295 ;
        RECT 22.485 165.125 22.740 165.695 ;
        RECT 22.915 165.140 23.205 165.865 ;
        RECT 23.925 165.315 24.095 165.695 ;
        RECT 24.275 165.485 24.605 165.865 ;
        RECT 23.925 165.145 24.590 165.315 ;
        RECT 24.785 165.190 25.045 165.695 ;
        RECT 21.385 163.995 21.555 165.125 ;
        RECT 22.145 164.955 22.315 165.125 ;
        RECT 20.430 163.825 21.555 163.995 ;
        RECT 21.725 164.625 21.920 164.955 ;
        RECT 22.145 164.625 22.400 164.955 ;
        RECT 21.725 163.655 21.895 164.625 ;
        RECT 22.570 164.455 22.740 165.125 ;
        RECT 23.855 164.595 24.185 164.965 ;
        RECT 24.420 164.890 24.590 165.145 ;
        RECT 24.420 164.560 24.705 164.890 ;
        RECT 19.865 163.485 21.895 163.655 ;
        RECT 22.065 163.315 22.235 164.455 ;
        RECT 22.405 163.485 22.740 164.455 ;
        RECT 22.915 163.315 23.205 164.480 ;
        RECT 24.420 164.415 24.590 164.560 ;
        RECT 23.925 164.245 24.590 164.415 ;
        RECT 24.875 164.390 25.045 165.190 ;
        RECT 23.925 163.485 24.095 164.245 ;
        RECT 24.275 163.315 24.605 164.075 ;
        RECT 24.775 163.485 25.045 164.390 ;
        RECT 25.215 165.190 25.475 165.695 ;
        RECT 25.655 165.485 25.985 165.865 ;
        RECT 26.165 165.315 26.335 165.695 ;
        RECT 25.215 164.390 25.385 165.190 ;
        RECT 25.670 165.145 26.335 165.315 ;
        RECT 26.710 165.235 26.995 165.695 ;
        RECT 27.165 165.405 27.435 165.865 ;
        RECT 25.670 164.890 25.840 165.145 ;
        RECT 26.710 165.065 27.665 165.235 ;
        RECT 25.555 164.560 25.840 164.890 ;
        RECT 26.075 164.595 26.405 164.965 ;
        RECT 25.670 164.415 25.840 164.560 ;
        RECT 25.215 163.485 25.485 164.390 ;
        RECT 25.670 164.245 26.335 164.415 ;
        RECT 26.595 164.335 27.285 164.895 ;
        RECT 25.655 163.315 25.985 164.075 ;
        RECT 26.165 163.485 26.335 164.245 ;
        RECT 27.455 164.165 27.665 165.065 ;
        RECT 26.710 163.945 27.665 164.165 ;
        RECT 27.835 164.895 28.235 165.695 ;
        RECT 28.425 165.235 28.705 165.695 ;
        RECT 29.225 165.405 29.550 165.865 ;
        RECT 28.425 165.065 29.550 165.235 ;
        RECT 29.720 165.125 30.105 165.695 ;
        RECT 30.365 165.385 30.665 165.865 ;
        RECT 30.835 165.215 31.095 165.670 ;
        RECT 31.265 165.385 31.525 165.865 ;
        RECT 31.705 165.215 31.965 165.670 ;
        RECT 32.135 165.385 32.385 165.865 ;
        RECT 32.565 165.215 32.825 165.670 ;
        RECT 32.995 165.385 33.245 165.865 ;
        RECT 33.425 165.215 33.685 165.670 ;
        RECT 33.855 165.385 34.100 165.865 ;
        RECT 34.270 165.215 34.545 165.670 ;
        RECT 34.715 165.385 34.960 165.865 ;
        RECT 35.130 165.215 35.390 165.670 ;
        RECT 35.560 165.385 35.820 165.865 ;
        RECT 35.990 165.215 36.250 165.670 ;
        RECT 36.420 165.385 36.680 165.865 ;
        RECT 36.850 165.215 37.110 165.670 ;
        RECT 37.280 165.305 37.540 165.865 ;
        RECT 30.365 165.185 37.110 165.215 ;
        RECT 29.100 164.955 29.550 165.065 ;
        RECT 27.835 164.335 28.930 164.895 ;
        RECT 29.100 164.625 29.655 164.955 ;
        RECT 26.710 163.485 26.995 163.945 ;
        RECT 27.165 163.315 27.435 163.775 ;
        RECT 27.835 163.485 28.235 164.335 ;
        RECT 29.100 164.165 29.550 164.625 ;
        RECT 29.825 164.455 30.105 165.125 ;
        RECT 30.335 165.045 37.110 165.185 ;
        RECT 30.335 165.015 31.530 165.045 ;
        RECT 28.425 163.945 29.550 164.165 ;
        RECT 28.425 163.485 28.705 163.945 ;
        RECT 29.225 163.315 29.550 163.775 ;
        RECT 29.720 163.485 30.105 164.455 ;
        RECT 30.365 164.455 31.530 165.015 ;
        RECT 37.710 164.875 37.960 165.685 ;
        RECT 38.140 165.340 38.400 165.865 ;
        RECT 38.570 164.875 38.820 165.685 ;
        RECT 39.000 165.355 39.305 165.865 ;
        RECT 31.700 164.625 38.820 164.875 ;
        RECT 38.990 164.625 39.305 165.185 ;
        RECT 39.480 165.155 39.735 165.685 ;
        RECT 39.905 165.405 40.210 165.865 ;
        RECT 40.455 165.485 41.525 165.655 ;
        RECT 30.365 164.230 37.110 164.455 ;
        RECT 30.365 163.315 30.635 164.060 ;
        RECT 30.805 163.490 31.095 164.230 ;
        RECT 31.705 164.215 37.110 164.230 ;
        RECT 31.265 163.320 31.520 164.045 ;
        RECT 31.705 163.490 31.965 164.215 ;
        RECT 32.135 163.320 32.380 164.045 ;
        RECT 32.565 163.490 32.825 164.215 ;
        RECT 32.995 163.320 33.240 164.045 ;
        RECT 33.425 163.490 33.685 164.215 ;
        RECT 33.855 163.320 34.100 164.045 ;
        RECT 34.270 163.490 34.530 164.215 ;
        RECT 34.700 163.320 34.960 164.045 ;
        RECT 35.130 163.490 35.390 164.215 ;
        RECT 35.560 163.320 35.820 164.045 ;
        RECT 35.990 163.490 36.250 164.215 ;
        RECT 36.420 163.320 36.680 164.045 ;
        RECT 36.850 163.490 37.110 164.215 ;
        RECT 37.280 163.320 37.540 164.115 ;
        RECT 37.710 163.490 37.960 164.625 ;
        RECT 31.265 163.315 37.540 163.320 ;
        RECT 38.140 163.315 38.400 164.125 ;
        RECT 38.575 163.485 38.820 164.625 ;
        RECT 39.480 164.505 39.690 165.155 ;
        RECT 40.455 165.130 40.775 165.485 ;
        RECT 40.450 164.955 40.775 165.130 ;
        RECT 39.860 164.655 40.775 164.955 ;
        RECT 40.945 164.915 41.185 165.315 ;
        RECT 41.355 165.255 41.525 165.485 ;
        RECT 41.695 165.425 41.885 165.865 ;
        RECT 42.055 165.415 43.005 165.695 ;
        RECT 43.225 165.505 43.575 165.675 ;
        RECT 41.355 165.085 41.885 165.255 ;
        RECT 39.860 164.625 40.600 164.655 ;
        RECT 39.000 163.315 39.295 164.125 ;
        RECT 39.480 163.625 39.735 164.505 ;
        RECT 39.905 163.315 40.210 164.455 ;
        RECT 40.430 164.035 40.600 164.625 ;
        RECT 40.945 164.545 41.485 164.915 ;
        RECT 41.665 164.805 41.885 165.085 ;
        RECT 42.055 164.635 42.225 165.415 ;
        RECT 41.820 164.465 42.225 164.635 ;
        RECT 42.395 164.625 42.745 165.245 ;
        RECT 41.820 164.375 41.990 164.465 ;
        RECT 42.915 164.455 43.125 165.245 ;
        RECT 40.770 164.205 41.990 164.375 ;
        RECT 42.450 164.295 43.125 164.455 ;
        RECT 40.430 163.865 41.230 164.035 ;
        RECT 40.550 163.315 40.880 163.695 ;
        RECT 41.060 163.575 41.230 163.865 ;
        RECT 41.820 163.825 41.990 164.205 ;
        RECT 42.160 164.285 43.125 164.295 ;
        RECT 43.315 165.115 43.575 165.505 ;
        RECT 43.785 165.405 44.115 165.865 ;
        RECT 44.990 165.475 45.845 165.645 ;
        RECT 46.050 165.475 46.545 165.645 ;
        RECT 46.715 165.505 47.045 165.865 ;
        RECT 43.315 164.425 43.485 165.115 ;
        RECT 43.655 164.765 43.825 164.945 ;
        RECT 43.995 164.935 44.785 165.185 ;
        RECT 44.990 164.765 45.160 165.475 ;
        RECT 45.330 164.965 45.685 165.185 ;
        RECT 43.655 164.595 45.345 164.765 ;
        RECT 42.160 163.995 42.620 164.285 ;
        RECT 43.315 164.255 44.815 164.425 ;
        RECT 43.315 164.115 43.485 164.255 ;
        RECT 42.925 163.945 43.485 164.115 ;
        RECT 41.400 163.315 41.650 163.775 ;
        RECT 41.820 163.485 42.690 163.825 ;
        RECT 42.925 163.485 43.095 163.945 ;
        RECT 43.930 163.915 45.005 164.085 ;
        RECT 43.265 163.315 43.635 163.775 ;
        RECT 43.930 163.575 44.100 163.915 ;
        RECT 44.270 163.315 44.600 163.745 ;
        RECT 44.835 163.575 45.005 163.915 ;
        RECT 45.175 163.815 45.345 164.595 ;
        RECT 45.515 164.375 45.685 164.965 ;
        RECT 45.855 164.565 46.205 165.185 ;
        RECT 45.515 163.985 45.980 164.375 ;
        RECT 46.375 164.115 46.545 165.475 ;
        RECT 46.715 164.285 47.175 165.335 ;
        RECT 46.150 163.945 46.545 164.115 ;
        RECT 46.150 163.815 46.320 163.945 ;
        RECT 45.175 163.485 45.855 163.815 ;
        RECT 46.070 163.485 46.320 163.815 ;
        RECT 46.490 163.315 46.740 163.775 ;
        RECT 46.910 163.500 47.235 164.285 ;
        RECT 47.405 163.485 47.575 165.605 ;
        RECT 47.745 165.485 48.075 165.865 ;
        RECT 48.245 165.315 48.500 165.605 ;
        RECT 47.750 165.145 48.500 165.315 ;
        RECT 47.750 164.155 47.980 165.145 ;
        RECT 48.675 165.140 48.965 165.865 ;
        RECT 50.060 165.155 50.315 165.685 ;
        RECT 50.485 165.405 50.790 165.865 ;
        RECT 51.035 165.485 52.105 165.655 ;
        RECT 48.150 164.325 48.500 164.975 ;
        RECT 50.060 164.505 50.270 165.155 ;
        RECT 51.035 165.130 51.355 165.485 ;
        RECT 51.030 164.955 51.355 165.130 ;
        RECT 50.440 164.655 51.355 164.955 ;
        RECT 51.525 164.915 51.765 165.315 ;
        RECT 51.935 165.255 52.105 165.485 ;
        RECT 52.275 165.425 52.465 165.865 ;
        RECT 52.635 165.415 53.585 165.695 ;
        RECT 53.805 165.505 54.155 165.675 ;
        RECT 51.935 165.085 52.465 165.255 ;
        RECT 50.440 164.625 51.180 164.655 ;
        RECT 47.750 163.985 48.500 164.155 ;
        RECT 47.745 163.315 48.075 163.815 ;
        RECT 48.245 163.485 48.500 163.985 ;
        RECT 48.675 163.315 48.965 164.480 ;
        RECT 50.060 163.625 50.315 164.505 ;
        RECT 50.485 163.315 50.790 164.455 ;
        RECT 51.010 164.035 51.180 164.625 ;
        RECT 51.525 164.545 52.065 164.915 ;
        RECT 52.245 164.805 52.465 165.085 ;
        RECT 52.635 164.635 52.805 165.415 ;
        RECT 52.400 164.465 52.805 164.635 ;
        RECT 52.975 164.625 53.325 165.245 ;
        RECT 52.400 164.375 52.570 164.465 ;
        RECT 53.495 164.455 53.705 165.245 ;
        RECT 51.350 164.205 52.570 164.375 ;
        RECT 53.030 164.295 53.705 164.455 ;
        RECT 51.010 163.865 51.810 164.035 ;
        RECT 51.130 163.315 51.460 163.695 ;
        RECT 51.640 163.575 51.810 163.865 ;
        RECT 52.400 163.825 52.570 164.205 ;
        RECT 52.740 164.285 53.705 164.295 ;
        RECT 53.895 165.115 54.155 165.505 ;
        RECT 54.365 165.405 54.695 165.865 ;
        RECT 55.570 165.475 56.425 165.645 ;
        RECT 56.630 165.475 57.125 165.645 ;
        RECT 57.295 165.505 57.625 165.865 ;
        RECT 53.895 164.425 54.065 165.115 ;
        RECT 54.235 164.765 54.405 164.945 ;
        RECT 54.575 164.935 55.365 165.185 ;
        RECT 55.570 164.765 55.740 165.475 ;
        RECT 55.910 164.965 56.265 165.185 ;
        RECT 54.235 164.595 55.925 164.765 ;
        RECT 52.740 163.995 53.200 164.285 ;
        RECT 53.895 164.255 55.395 164.425 ;
        RECT 53.895 164.115 54.065 164.255 ;
        RECT 53.505 163.945 54.065 164.115 ;
        RECT 51.980 163.315 52.230 163.775 ;
        RECT 52.400 163.485 53.270 163.825 ;
        RECT 53.505 163.485 53.675 163.945 ;
        RECT 54.510 163.915 55.585 164.085 ;
        RECT 53.845 163.315 54.215 163.775 ;
        RECT 54.510 163.575 54.680 163.915 ;
        RECT 54.850 163.315 55.180 163.745 ;
        RECT 55.415 163.575 55.585 163.915 ;
        RECT 55.755 163.815 55.925 164.595 ;
        RECT 56.095 164.375 56.265 164.965 ;
        RECT 56.435 164.565 56.785 165.185 ;
        RECT 56.095 163.985 56.560 164.375 ;
        RECT 56.955 164.115 57.125 165.475 ;
        RECT 57.295 164.285 57.755 165.335 ;
        RECT 56.730 163.945 57.125 164.115 ;
        RECT 56.730 163.815 56.900 163.945 ;
        RECT 55.755 163.485 56.435 163.815 ;
        RECT 56.650 163.485 56.900 163.815 ;
        RECT 57.070 163.315 57.320 163.775 ;
        RECT 57.490 163.500 57.815 164.285 ;
        RECT 57.985 163.485 58.155 165.605 ;
        RECT 58.325 165.485 58.655 165.865 ;
        RECT 58.825 165.315 59.080 165.605 ;
        RECT 58.330 165.145 59.080 165.315 ;
        RECT 58.330 164.155 58.560 165.145 ;
        RECT 59.405 165.065 59.735 165.865 ;
        RECT 59.905 165.215 60.075 165.695 ;
        RECT 60.245 165.385 60.575 165.865 ;
        RECT 60.745 165.215 60.915 165.695 ;
        RECT 61.165 165.385 61.405 165.865 ;
        RECT 61.585 165.215 61.755 165.695 ;
        RECT 62.075 165.385 62.355 165.865 ;
        RECT 62.525 165.215 62.785 165.605 ;
        RECT 62.960 165.385 63.215 165.865 ;
        RECT 63.385 165.215 63.680 165.605 ;
        RECT 63.860 165.385 64.135 165.865 ;
        RECT 64.305 165.365 64.605 165.695 ;
        RECT 59.905 165.045 60.915 165.215 ;
        RECT 61.120 165.045 61.755 165.215 ;
        RECT 62.030 165.045 63.680 165.215 ;
        RECT 58.730 164.325 59.080 164.975 ;
        RECT 59.905 164.505 60.400 165.045 ;
        RECT 61.120 164.875 61.290 165.045 ;
        RECT 60.790 164.705 61.290 164.875 ;
        RECT 58.330 163.985 59.080 164.155 ;
        RECT 58.325 163.315 58.655 163.815 ;
        RECT 58.825 163.485 59.080 163.985 ;
        RECT 59.405 163.315 59.735 164.465 ;
        RECT 59.905 164.335 60.915 164.505 ;
        RECT 59.905 163.485 60.075 164.335 ;
        RECT 60.245 163.315 60.575 164.115 ;
        RECT 60.745 163.485 60.915 164.335 ;
        RECT 61.120 164.465 61.290 164.705 ;
        RECT 61.460 164.635 61.840 164.875 ;
        RECT 62.030 164.535 62.435 165.045 ;
        RECT 62.605 164.705 63.745 164.875 ;
        RECT 61.120 164.295 61.835 164.465 ;
        RECT 62.030 164.365 62.785 164.535 ;
        RECT 61.095 163.315 61.335 164.115 ;
        RECT 61.505 163.485 61.835 164.295 ;
        RECT 62.070 163.315 62.355 164.185 ;
        RECT 62.525 164.115 62.785 164.365 ;
        RECT 63.575 164.455 63.745 164.705 ;
        RECT 63.915 164.625 64.265 165.195 ;
        RECT 64.435 164.455 64.605 165.365 ;
        RECT 64.780 165.320 70.125 165.865 ;
        RECT 63.575 164.285 64.605 164.455 ;
        RECT 62.525 163.945 63.645 164.115 ;
        RECT 62.525 163.485 62.785 163.945 ;
        RECT 62.960 163.315 63.215 163.775 ;
        RECT 63.385 163.485 63.645 163.945 ;
        RECT 63.815 163.315 64.125 164.115 ;
        RECT 64.295 163.485 64.605 164.285 ;
        RECT 66.370 163.750 66.720 165.000 ;
        RECT 68.200 164.490 68.540 165.320 ;
        RECT 70.570 165.055 70.815 165.660 ;
        RECT 71.035 165.330 71.545 165.865 ;
        RECT 70.295 164.885 71.525 165.055 ;
        RECT 70.295 164.075 70.635 164.885 ;
        RECT 70.805 164.320 71.555 164.510 ;
        RECT 64.780 163.315 70.125 163.750 ;
        RECT 70.295 163.665 70.810 164.075 ;
        RECT 71.045 163.315 71.215 164.075 ;
        RECT 71.385 163.655 71.555 164.320 ;
        RECT 71.725 164.335 71.915 165.695 ;
        RECT 72.085 165.185 72.360 165.695 ;
        RECT 72.550 165.330 73.080 165.695 ;
        RECT 73.505 165.465 73.835 165.865 ;
        RECT 72.905 165.295 73.080 165.330 ;
        RECT 72.085 165.015 72.365 165.185 ;
        RECT 72.085 164.535 72.360 165.015 ;
        RECT 72.565 164.335 72.735 165.135 ;
        RECT 71.725 164.165 72.735 164.335 ;
        RECT 72.905 165.125 73.835 165.295 ;
        RECT 74.005 165.125 74.260 165.695 ;
        RECT 74.435 165.140 74.725 165.865 ;
        RECT 74.985 165.315 75.155 165.695 ;
        RECT 75.335 165.485 75.665 165.865 ;
        RECT 74.985 165.145 75.650 165.315 ;
        RECT 75.845 165.190 76.105 165.695 ;
        RECT 72.905 163.995 73.075 165.125 ;
        RECT 73.665 164.955 73.835 165.125 ;
        RECT 71.950 163.825 73.075 163.995 ;
        RECT 73.245 164.625 73.440 164.955 ;
        RECT 73.665 164.625 73.920 164.955 ;
        RECT 73.245 163.655 73.415 164.625 ;
        RECT 74.090 164.455 74.260 165.125 ;
        RECT 74.915 164.595 75.245 164.965 ;
        RECT 75.480 164.890 75.650 165.145 ;
        RECT 75.480 164.560 75.765 164.890 ;
        RECT 71.385 163.485 73.415 163.655 ;
        RECT 73.585 163.315 73.755 164.455 ;
        RECT 73.925 163.485 74.260 164.455 ;
        RECT 74.435 163.315 74.725 164.480 ;
        RECT 75.480 164.415 75.650 164.560 ;
        RECT 74.985 164.245 75.650 164.415 ;
        RECT 75.935 164.390 76.105 165.190 ;
        RECT 76.795 165.045 77.005 165.865 ;
        RECT 77.175 165.065 77.505 165.695 ;
        RECT 77.175 164.465 77.425 165.065 ;
        RECT 77.675 165.045 77.905 165.865 ;
        RECT 78.175 165.045 78.385 165.865 ;
        RECT 78.555 165.065 78.885 165.695 ;
        RECT 77.595 164.625 77.925 164.875 ;
        RECT 78.555 164.465 78.805 165.065 ;
        RECT 79.055 165.045 79.285 165.865 ;
        RECT 79.870 165.155 80.125 165.685 ;
        RECT 80.305 165.405 80.590 165.865 ;
        RECT 78.975 164.625 79.305 164.875 ;
        RECT 74.985 163.485 75.155 164.245 ;
        RECT 75.335 163.315 75.665 164.075 ;
        RECT 75.835 163.485 76.105 164.390 ;
        RECT 76.795 163.315 77.005 164.455 ;
        RECT 77.175 163.485 77.505 164.465 ;
        RECT 77.675 163.315 77.905 164.455 ;
        RECT 78.175 163.315 78.385 164.455 ;
        RECT 78.555 163.485 78.885 164.465 ;
        RECT 79.055 163.315 79.285 164.455 ;
        RECT 79.870 164.295 80.050 165.155 ;
        RECT 80.770 164.955 81.020 165.605 ;
        RECT 80.220 164.625 81.020 164.955 ;
        RECT 79.870 164.165 80.125 164.295 ;
        RECT 79.785 163.995 80.125 164.165 ;
        RECT 79.870 163.625 80.125 163.995 ;
        RECT 80.305 163.315 80.590 164.115 ;
        RECT 80.770 164.035 81.020 164.625 ;
        RECT 81.220 165.270 81.540 165.600 ;
        RECT 81.720 165.385 82.380 165.865 ;
        RECT 82.580 165.475 83.430 165.645 ;
        RECT 81.220 164.375 81.410 165.270 ;
        RECT 81.730 164.945 82.390 165.215 ;
        RECT 82.060 164.885 82.390 164.945 ;
        RECT 81.580 164.715 81.910 164.775 ;
        RECT 82.580 164.715 82.750 165.475 ;
        RECT 83.990 165.405 84.310 165.865 ;
        RECT 84.510 165.225 84.760 165.655 ;
        RECT 85.050 165.425 85.460 165.865 ;
        RECT 85.630 165.485 86.645 165.685 ;
        RECT 82.920 165.055 84.170 165.225 ;
        RECT 82.920 164.935 83.250 165.055 ;
        RECT 81.580 164.545 83.480 164.715 ;
        RECT 81.220 164.205 83.140 164.375 ;
        RECT 81.220 164.185 81.540 164.205 ;
        RECT 80.770 163.525 81.100 164.035 ;
        RECT 81.370 163.575 81.540 164.185 ;
        RECT 83.310 164.035 83.480 164.545 ;
        RECT 83.650 164.475 83.830 164.885 ;
        RECT 84.000 164.295 84.170 165.055 ;
        RECT 81.710 163.315 82.040 164.005 ;
        RECT 82.270 163.865 83.480 164.035 ;
        RECT 83.650 163.985 84.170 164.295 ;
        RECT 84.340 164.885 84.760 165.225 ;
        RECT 85.050 164.885 85.460 165.215 ;
        RECT 84.340 164.115 84.530 164.885 ;
        RECT 85.630 164.755 85.800 165.485 ;
        RECT 86.945 165.315 87.115 165.645 ;
        RECT 87.285 165.485 87.615 165.865 ;
        RECT 85.970 164.935 86.320 165.305 ;
        RECT 85.630 164.715 86.050 164.755 ;
        RECT 84.700 164.545 86.050 164.715 ;
        RECT 84.700 164.385 84.950 164.545 ;
        RECT 85.460 164.115 85.710 164.375 ;
        RECT 84.340 163.865 85.710 164.115 ;
        RECT 82.270 163.575 82.510 163.865 ;
        RECT 83.310 163.785 83.480 163.865 ;
        RECT 82.710 163.315 83.130 163.695 ;
        RECT 83.310 163.535 83.940 163.785 ;
        RECT 84.410 163.315 84.740 163.695 ;
        RECT 84.910 163.575 85.080 163.865 ;
        RECT 85.880 163.700 86.050 164.545 ;
        RECT 86.500 164.375 86.720 165.245 ;
        RECT 86.945 165.125 87.640 165.315 ;
        RECT 86.220 163.995 86.720 164.375 ;
        RECT 86.890 164.325 87.300 164.945 ;
        RECT 87.470 164.155 87.640 165.125 ;
        RECT 86.945 163.985 87.640 164.155 ;
        RECT 85.260 163.315 85.640 163.695 ;
        RECT 85.880 163.530 86.710 163.700 ;
        RECT 86.945 163.485 87.115 163.985 ;
        RECT 87.285 163.315 87.615 163.815 ;
        RECT 87.830 163.485 88.055 165.605 ;
        RECT 88.225 165.485 88.555 165.865 ;
        RECT 88.725 165.315 88.895 165.605 ;
        RECT 88.230 165.145 88.895 165.315 ;
        RECT 89.530 165.155 89.785 165.685 ;
        RECT 89.965 165.405 90.250 165.865 ;
        RECT 88.230 164.155 88.460 165.145 ;
        RECT 88.630 164.325 88.980 164.975 ;
        RECT 89.530 164.295 89.710 165.155 ;
        RECT 90.430 164.955 90.680 165.605 ;
        RECT 89.880 164.625 90.680 164.955 ;
        RECT 88.230 163.985 88.895 164.155 ;
        RECT 88.225 163.315 88.555 163.815 ;
        RECT 88.725 163.485 88.895 163.985 ;
        RECT 89.530 163.825 89.785 164.295 ;
        RECT 89.445 163.655 89.785 163.825 ;
        RECT 89.530 163.625 89.785 163.655 ;
        RECT 89.965 163.315 90.250 164.115 ;
        RECT 90.430 164.035 90.680 164.625 ;
        RECT 90.880 165.270 91.200 165.600 ;
        RECT 91.380 165.385 92.040 165.865 ;
        RECT 92.240 165.475 93.090 165.645 ;
        RECT 90.880 164.375 91.070 165.270 ;
        RECT 91.390 164.945 92.050 165.215 ;
        RECT 91.720 164.885 92.050 164.945 ;
        RECT 91.240 164.715 91.570 164.775 ;
        RECT 92.240 164.715 92.410 165.475 ;
        RECT 93.650 165.405 93.970 165.865 ;
        RECT 94.170 165.225 94.420 165.655 ;
        RECT 94.710 165.425 95.120 165.865 ;
        RECT 95.290 165.485 96.305 165.685 ;
        RECT 92.580 165.055 93.830 165.225 ;
        RECT 92.580 164.935 92.910 165.055 ;
        RECT 91.240 164.545 93.140 164.715 ;
        RECT 90.880 164.205 92.800 164.375 ;
        RECT 90.880 164.185 91.200 164.205 ;
        RECT 90.430 163.525 90.760 164.035 ;
        RECT 91.030 163.575 91.200 164.185 ;
        RECT 92.970 164.035 93.140 164.545 ;
        RECT 93.310 164.475 93.490 164.885 ;
        RECT 93.660 164.295 93.830 165.055 ;
        RECT 91.370 163.315 91.700 164.005 ;
        RECT 91.930 163.865 93.140 164.035 ;
        RECT 93.310 163.985 93.830 164.295 ;
        RECT 94.000 164.885 94.420 165.225 ;
        RECT 94.710 164.885 95.120 165.215 ;
        RECT 94.000 164.115 94.190 164.885 ;
        RECT 95.290 164.755 95.460 165.485 ;
        RECT 96.605 165.315 96.775 165.645 ;
        RECT 96.945 165.485 97.275 165.865 ;
        RECT 95.630 164.935 95.980 165.305 ;
        RECT 95.290 164.715 95.710 164.755 ;
        RECT 94.360 164.545 95.710 164.715 ;
        RECT 94.360 164.385 94.610 164.545 ;
        RECT 95.120 164.115 95.370 164.375 ;
        RECT 94.000 163.865 95.370 164.115 ;
        RECT 91.930 163.575 92.170 163.865 ;
        RECT 92.970 163.785 93.140 163.865 ;
        RECT 92.370 163.315 92.790 163.695 ;
        RECT 92.970 163.535 93.600 163.785 ;
        RECT 94.070 163.315 94.400 163.695 ;
        RECT 94.570 163.575 94.740 163.865 ;
        RECT 95.540 163.700 95.710 164.545 ;
        RECT 96.160 164.375 96.380 165.245 ;
        RECT 96.605 165.125 97.300 165.315 ;
        RECT 95.880 163.995 96.380 164.375 ;
        RECT 96.550 164.325 96.960 164.945 ;
        RECT 97.130 164.155 97.300 165.125 ;
        RECT 96.605 163.985 97.300 164.155 ;
        RECT 94.920 163.315 95.300 163.695 ;
        RECT 95.540 163.530 96.370 163.700 ;
        RECT 96.605 163.485 96.775 163.985 ;
        RECT 96.945 163.315 97.275 163.815 ;
        RECT 97.490 163.485 97.715 165.605 ;
        RECT 97.885 165.485 98.215 165.865 ;
        RECT 98.385 165.315 98.555 165.605 ;
        RECT 97.890 165.145 98.555 165.315 ;
        RECT 98.905 165.315 99.075 165.695 ;
        RECT 99.255 165.485 99.585 165.865 ;
        RECT 98.905 165.145 99.570 165.315 ;
        RECT 99.765 165.190 100.025 165.695 ;
        RECT 97.890 164.155 98.120 165.145 ;
        RECT 98.290 164.325 98.640 164.975 ;
        RECT 98.835 164.595 99.165 164.965 ;
        RECT 99.400 164.890 99.570 165.145 ;
        RECT 99.400 164.560 99.685 164.890 ;
        RECT 99.400 164.415 99.570 164.560 ;
        RECT 98.905 164.245 99.570 164.415 ;
        RECT 99.855 164.390 100.025 165.190 ;
        RECT 100.195 165.140 100.485 165.865 ;
        RECT 100.695 165.045 100.925 165.865 ;
        RECT 101.095 165.065 101.425 165.695 ;
        RECT 100.675 164.625 101.005 164.875 ;
        RECT 97.890 163.985 98.555 164.155 ;
        RECT 97.885 163.315 98.215 163.815 ;
        RECT 98.385 163.485 98.555 163.985 ;
        RECT 98.905 163.485 99.075 164.245 ;
        RECT 99.255 163.315 99.585 164.075 ;
        RECT 99.755 163.485 100.025 164.390 ;
        RECT 100.195 163.315 100.485 164.480 ;
        RECT 101.175 164.465 101.425 165.065 ;
        RECT 101.595 165.045 101.805 165.865 ;
        RECT 102.040 165.155 102.295 165.685 ;
        RECT 102.465 165.405 102.770 165.865 ;
        RECT 103.015 165.485 104.085 165.655 ;
        RECT 100.695 163.315 100.925 164.455 ;
        RECT 101.095 163.485 101.425 164.465 ;
        RECT 102.040 164.505 102.250 165.155 ;
        RECT 103.015 165.130 103.335 165.485 ;
        RECT 103.010 164.955 103.335 165.130 ;
        RECT 102.420 164.655 103.335 164.955 ;
        RECT 103.505 164.915 103.745 165.315 ;
        RECT 103.915 165.255 104.085 165.485 ;
        RECT 104.255 165.425 104.445 165.865 ;
        RECT 104.615 165.415 105.565 165.695 ;
        RECT 105.785 165.505 106.135 165.675 ;
        RECT 103.915 165.085 104.445 165.255 ;
        RECT 102.420 164.625 103.160 164.655 ;
        RECT 101.595 163.315 101.805 164.455 ;
        RECT 102.040 163.625 102.295 164.505 ;
        RECT 102.465 163.315 102.770 164.455 ;
        RECT 102.990 164.035 103.160 164.625 ;
        RECT 103.505 164.545 104.045 164.915 ;
        RECT 104.225 164.805 104.445 165.085 ;
        RECT 104.615 164.635 104.785 165.415 ;
        RECT 104.380 164.465 104.785 164.635 ;
        RECT 104.955 164.625 105.305 165.245 ;
        RECT 104.380 164.375 104.550 164.465 ;
        RECT 105.475 164.455 105.685 165.245 ;
        RECT 103.330 164.205 104.550 164.375 ;
        RECT 105.010 164.295 105.685 164.455 ;
        RECT 102.990 163.865 103.790 164.035 ;
        RECT 103.110 163.315 103.440 163.695 ;
        RECT 103.620 163.575 103.790 163.865 ;
        RECT 104.380 163.825 104.550 164.205 ;
        RECT 104.720 164.285 105.685 164.295 ;
        RECT 105.875 165.115 106.135 165.505 ;
        RECT 106.345 165.405 106.675 165.865 ;
        RECT 107.550 165.475 108.405 165.645 ;
        RECT 108.610 165.475 109.105 165.645 ;
        RECT 109.275 165.505 109.605 165.865 ;
        RECT 105.875 164.425 106.045 165.115 ;
        RECT 106.215 164.765 106.385 164.945 ;
        RECT 106.555 164.935 107.345 165.185 ;
        RECT 107.550 164.765 107.720 165.475 ;
        RECT 107.890 164.965 108.245 165.185 ;
        RECT 106.215 164.595 107.905 164.765 ;
        RECT 104.720 163.995 105.180 164.285 ;
        RECT 105.875 164.255 107.375 164.425 ;
        RECT 105.875 164.115 106.045 164.255 ;
        RECT 105.485 163.945 106.045 164.115 ;
        RECT 103.960 163.315 104.210 163.775 ;
        RECT 104.380 163.485 105.250 163.825 ;
        RECT 105.485 163.485 105.655 163.945 ;
        RECT 106.490 163.915 107.565 164.085 ;
        RECT 105.825 163.315 106.195 163.775 ;
        RECT 106.490 163.575 106.660 163.915 ;
        RECT 106.830 163.315 107.160 163.745 ;
        RECT 107.395 163.575 107.565 163.915 ;
        RECT 107.735 163.815 107.905 164.595 ;
        RECT 108.075 164.375 108.245 164.965 ;
        RECT 108.415 164.565 108.765 165.185 ;
        RECT 108.075 163.985 108.540 164.375 ;
        RECT 108.935 164.115 109.105 165.475 ;
        RECT 109.275 164.285 109.735 165.335 ;
        RECT 108.710 163.945 109.105 164.115 ;
        RECT 108.710 163.815 108.880 163.945 ;
        RECT 107.735 163.485 108.415 163.815 ;
        RECT 108.630 163.485 108.880 163.815 ;
        RECT 109.050 163.315 109.300 163.775 ;
        RECT 109.470 163.500 109.795 164.285 ;
        RECT 109.965 163.485 110.135 165.605 ;
        RECT 110.305 165.485 110.635 165.865 ;
        RECT 110.805 165.315 111.060 165.605 ;
        RECT 110.310 165.145 111.060 165.315 ;
        RECT 110.310 164.155 110.540 165.145 ;
        RECT 112.155 165.115 113.365 165.865 ;
        RECT 110.710 164.325 111.060 164.975 ;
        RECT 112.155 164.405 112.675 164.945 ;
        RECT 112.845 164.575 113.365 165.115 ;
        RECT 110.310 163.985 111.060 164.155 ;
        RECT 110.305 163.315 110.635 163.815 ;
        RECT 110.805 163.485 111.060 163.985 ;
        RECT 112.155 163.315 113.365 164.405 ;
        RECT 15.010 163.145 113.450 163.315 ;
        RECT 15.095 162.055 16.305 163.145 ;
        RECT 15.095 161.345 15.615 161.885 ;
        RECT 15.785 161.515 16.305 162.055 ;
        RECT 16.850 162.165 17.105 162.835 ;
        RECT 17.285 162.345 17.570 163.145 ;
        RECT 17.750 162.425 18.080 162.935 ;
        RECT 15.095 160.595 16.305 161.345 ;
        RECT 16.850 161.305 17.030 162.165 ;
        RECT 17.750 161.835 18.000 162.425 ;
        RECT 18.350 162.275 18.520 162.885 ;
        RECT 18.690 162.455 19.020 163.145 ;
        RECT 19.250 162.595 19.490 162.885 ;
        RECT 19.690 162.765 20.110 163.145 ;
        RECT 20.290 162.675 20.920 162.925 ;
        RECT 21.390 162.765 21.720 163.145 ;
        RECT 20.290 162.595 20.460 162.675 ;
        RECT 21.890 162.595 22.060 162.885 ;
        RECT 22.240 162.765 22.620 163.145 ;
        RECT 22.860 162.760 23.690 162.930 ;
        RECT 19.250 162.425 20.460 162.595 ;
        RECT 17.200 161.505 18.000 161.835 ;
        RECT 16.850 161.105 17.105 161.305 ;
        RECT 16.765 160.935 17.105 161.105 ;
        RECT 16.850 160.775 17.105 160.935 ;
        RECT 17.285 160.595 17.570 161.055 ;
        RECT 17.750 160.855 18.000 161.505 ;
        RECT 18.200 162.255 18.520 162.275 ;
        RECT 18.200 162.085 20.120 162.255 ;
        RECT 18.200 161.190 18.390 162.085 ;
        RECT 20.290 161.915 20.460 162.425 ;
        RECT 20.630 162.165 21.150 162.475 ;
        RECT 18.560 161.745 20.460 161.915 ;
        RECT 18.560 161.685 18.890 161.745 ;
        RECT 19.040 161.515 19.370 161.575 ;
        RECT 18.710 161.245 19.370 161.515 ;
        RECT 18.200 160.860 18.520 161.190 ;
        RECT 18.700 160.595 19.360 161.075 ;
        RECT 19.560 160.985 19.730 161.745 ;
        RECT 20.630 161.575 20.810 161.985 ;
        RECT 19.900 161.405 20.230 161.525 ;
        RECT 20.980 161.405 21.150 162.165 ;
        RECT 19.900 161.235 21.150 161.405 ;
        RECT 21.320 162.345 22.690 162.595 ;
        RECT 21.320 161.575 21.510 162.345 ;
        RECT 22.440 162.085 22.690 162.345 ;
        RECT 21.680 161.915 21.930 162.075 ;
        RECT 22.860 161.915 23.030 162.760 ;
        RECT 23.925 162.475 24.095 162.975 ;
        RECT 24.265 162.645 24.595 163.145 ;
        RECT 23.200 162.085 23.700 162.465 ;
        RECT 23.925 162.305 24.620 162.475 ;
        RECT 21.680 161.745 23.030 161.915 ;
        RECT 22.610 161.705 23.030 161.745 ;
        RECT 21.320 161.235 21.740 161.575 ;
        RECT 22.030 161.245 22.440 161.575 ;
        RECT 19.560 160.815 20.410 160.985 ;
        RECT 20.970 160.595 21.290 161.055 ;
        RECT 21.490 160.805 21.740 161.235 ;
        RECT 22.030 160.595 22.440 161.035 ;
        RECT 22.610 160.975 22.780 161.705 ;
        RECT 22.950 161.155 23.300 161.525 ;
        RECT 23.480 161.215 23.700 162.085 ;
        RECT 23.870 161.515 24.280 162.135 ;
        RECT 24.450 161.335 24.620 162.305 ;
        RECT 23.925 161.145 24.620 161.335 ;
        RECT 22.610 160.775 23.625 160.975 ;
        RECT 23.925 160.815 24.095 161.145 ;
        RECT 24.265 160.595 24.595 160.975 ;
        RECT 24.810 160.855 25.035 162.975 ;
        RECT 25.205 162.645 25.535 163.145 ;
        RECT 25.705 162.475 25.875 162.975 ;
        RECT 25.210 162.305 25.875 162.475 ;
        RECT 25.210 161.315 25.440 162.305 ;
        RECT 25.610 161.485 25.960 162.135 ;
        RECT 26.140 162.005 26.475 162.975 ;
        RECT 26.645 162.005 26.815 163.145 ;
        RECT 26.985 162.805 29.015 162.975 ;
        RECT 26.140 161.335 26.310 162.005 ;
        RECT 26.985 161.835 27.155 162.805 ;
        RECT 26.480 161.505 26.735 161.835 ;
        RECT 26.960 161.505 27.155 161.835 ;
        RECT 27.325 162.465 28.450 162.635 ;
        RECT 26.565 161.335 26.735 161.505 ;
        RECT 27.325 161.335 27.495 162.465 ;
        RECT 25.210 161.145 25.875 161.315 ;
        RECT 25.205 160.595 25.535 160.975 ;
        RECT 25.705 160.855 25.875 161.145 ;
        RECT 26.140 160.765 26.395 161.335 ;
        RECT 26.565 161.165 27.495 161.335 ;
        RECT 27.665 162.125 28.675 162.295 ;
        RECT 27.665 161.325 27.835 162.125 ;
        RECT 27.320 161.130 27.495 161.165 ;
        RECT 26.565 160.595 26.895 160.995 ;
        RECT 27.320 160.765 27.850 161.130 ;
        RECT 28.040 161.105 28.315 161.925 ;
        RECT 28.035 160.935 28.315 161.105 ;
        RECT 28.040 160.765 28.315 160.935 ;
        RECT 28.485 160.765 28.675 162.125 ;
        RECT 28.845 162.140 29.015 162.805 ;
        RECT 29.185 162.385 29.355 163.145 ;
        RECT 29.590 162.385 30.105 162.795 ;
        RECT 28.845 161.950 29.595 162.140 ;
        RECT 29.765 161.575 30.105 162.385 ;
        RECT 30.315 162.005 30.545 163.145 ;
        RECT 30.715 161.995 31.045 162.975 ;
        RECT 31.215 162.005 31.425 163.145 ;
        RECT 31.655 162.385 32.170 162.795 ;
        RECT 32.405 162.385 32.575 163.145 ;
        RECT 32.745 162.805 34.775 162.975 ;
        RECT 30.295 161.585 30.625 161.835 ;
        RECT 28.875 161.405 30.105 161.575 ;
        RECT 28.855 160.595 29.365 161.130 ;
        RECT 29.585 160.800 29.830 161.405 ;
        RECT 30.315 160.595 30.545 161.415 ;
        RECT 30.795 161.395 31.045 161.995 ;
        RECT 31.655 161.575 31.995 162.385 ;
        RECT 32.745 162.140 32.915 162.805 ;
        RECT 33.310 162.465 34.435 162.635 ;
        RECT 32.165 161.950 32.915 162.140 ;
        RECT 33.085 162.125 34.095 162.295 ;
        RECT 30.715 160.765 31.045 161.395 ;
        RECT 31.215 160.595 31.425 161.415 ;
        RECT 31.655 161.405 32.885 161.575 ;
        RECT 31.930 160.800 32.175 161.405 ;
        RECT 32.395 160.595 32.905 161.130 ;
        RECT 33.085 160.765 33.275 162.125 ;
        RECT 33.445 161.785 33.720 161.925 ;
        RECT 33.445 161.615 33.725 161.785 ;
        RECT 33.445 160.765 33.720 161.615 ;
        RECT 33.925 161.325 34.095 162.125 ;
        RECT 34.265 161.335 34.435 162.465 ;
        RECT 34.605 161.835 34.775 162.805 ;
        RECT 34.945 162.005 35.115 163.145 ;
        RECT 35.285 162.005 35.620 162.975 ;
        RECT 34.605 161.505 34.800 161.835 ;
        RECT 35.025 161.505 35.280 161.835 ;
        RECT 35.025 161.335 35.195 161.505 ;
        RECT 35.450 161.335 35.620 162.005 ;
        RECT 35.795 161.980 36.085 163.145 ;
        RECT 36.715 162.055 39.305 163.145 ;
        RECT 39.475 162.385 39.990 162.795 ;
        RECT 40.225 162.385 40.395 163.145 ;
        RECT 40.565 162.805 42.595 162.975 ;
        RECT 36.715 161.535 37.925 162.055 ;
        RECT 38.095 161.365 39.305 161.885 ;
        RECT 39.475 161.575 39.815 162.385 ;
        RECT 40.565 162.140 40.735 162.805 ;
        RECT 41.130 162.465 42.255 162.635 ;
        RECT 39.985 161.950 40.735 162.140 ;
        RECT 40.905 162.125 41.915 162.295 ;
        RECT 39.475 161.405 40.705 161.575 ;
        RECT 34.265 161.165 35.195 161.335 ;
        RECT 34.265 161.130 34.440 161.165 ;
        RECT 33.910 160.765 34.440 161.130 ;
        RECT 34.865 160.595 35.195 160.995 ;
        RECT 35.365 160.765 35.620 161.335 ;
        RECT 35.795 160.595 36.085 161.320 ;
        RECT 36.715 160.595 39.305 161.365 ;
        RECT 39.750 160.800 39.995 161.405 ;
        RECT 40.215 160.595 40.725 161.130 ;
        RECT 40.905 160.765 41.095 162.125 ;
        RECT 41.265 161.785 41.540 161.925 ;
        RECT 41.265 161.615 41.545 161.785 ;
        RECT 41.265 160.765 41.540 161.615 ;
        RECT 41.745 161.325 41.915 162.125 ;
        RECT 42.085 161.335 42.255 162.465 ;
        RECT 42.425 161.835 42.595 162.805 ;
        RECT 42.765 162.005 42.935 163.145 ;
        RECT 43.105 162.005 43.440 162.975 ;
        RECT 44.625 162.215 44.795 162.975 ;
        RECT 44.975 162.385 45.305 163.145 ;
        RECT 44.625 162.045 45.290 162.215 ;
        RECT 45.475 162.070 45.745 162.975 ;
        RECT 46.030 162.515 46.315 162.975 ;
        RECT 46.485 162.685 46.755 163.145 ;
        RECT 46.030 162.295 46.985 162.515 ;
        RECT 42.425 161.505 42.620 161.835 ;
        RECT 42.845 161.505 43.100 161.835 ;
        RECT 42.845 161.335 43.015 161.505 ;
        RECT 43.270 161.335 43.440 162.005 ;
        RECT 45.120 161.900 45.290 162.045 ;
        RECT 44.555 161.495 44.885 161.865 ;
        RECT 45.120 161.570 45.405 161.900 ;
        RECT 42.085 161.165 43.015 161.335 ;
        RECT 42.085 161.130 42.260 161.165 ;
        RECT 41.730 160.765 42.260 161.130 ;
        RECT 42.685 160.595 43.015 160.995 ;
        RECT 43.185 160.765 43.440 161.335 ;
        RECT 45.120 161.315 45.290 161.570 ;
        RECT 44.625 161.145 45.290 161.315 ;
        RECT 45.575 161.270 45.745 162.070 ;
        RECT 45.915 161.565 46.605 162.125 ;
        RECT 46.775 161.395 46.985 162.295 ;
        RECT 44.625 160.765 44.795 161.145 ;
        RECT 44.975 160.595 45.305 160.975 ;
        RECT 45.485 160.765 45.745 161.270 ;
        RECT 46.030 161.225 46.985 161.395 ;
        RECT 47.155 162.125 47.555 162.975 ;
        RECT 47.745 162.515 48.025 162.975 ;
        RECT 48.545 162.685 48.870 163.145 ;
        RECT 47.745 162.295 48.870 162.515 ;
        RECT 47.155 161.565 48.250 162.125 ;
        RECT 48.420 161.835 48.870 162.295 ;
        RECT 49.040 162.005 49.425 162.975 ;
        RECT 46.030 160.765 46.315 161.225 ;
        RECT 46.485 160.595 46.755 161.055 ;
        RECT 47.155 160.765 47.555 161.565 ;
        RECT 48.420 161.505 48.975 161.835 ;
        RECT 48.420 161.395 48.870 161.505 ;
        RECT 47.745 161.225 48.870 161.395 ;
        RECT 49.145 161.335 49.425 162.005 ;
        RECT 49.595 162.385 50.110 162.795 ;
        RECT 50.345 162.385 50.515 163.145 ;
        RECT 50.685 162.805 52.715 162.975 ;
        RECT 49.595 161.575 49.935 162.385 ;
        RECT 50.685 162.140 50.855 162.805 ;
        RECT 51.250 162.465 52.375 162.635 ;
        RECT 50.105 161.950 50.855 162.140 ;
        RECT 51.025 162.125 52.035 162.295 ;
        RECT 49.595 161.405 50.825 161.575 ;
        RECT 47.745 160.765 48.025 161.225 ;
        RECT 48.545 160.595 48.870 161.055 ;
        RECT 49.040 160.765 49.425 161.335 ;
        RECT 49.870 160.800 50.115 161.405 ;
        RECT 50.335 160.595 50.845 161.130 ;
        RECT 51.025 160.765 51.215 162.125 ;
        RECT 51.385 161.785 51.660 161.925 ;
        RECT 51.385 161.615 51.665 161.785 ;
        RECT 51.385 160.765 51.660 161.615 ;
        RECT 51.865 161.325 52.035 162.125 ;
        RECT 52.205 161.335 52.375 162.465 ;
        RECT 52.545 161.835 52.715 162.805 ;
        RECT 52.885 162.005 53.055 163.145 ;
        RECT 53.225 162.005 53.560 162.975 ;
        RECT 54.745 162.215 54.915 162.975 ;
        RECT 55.095 162.385 55.425 163.145 ;
        RECT 54.745 162.045 55.410 162.215 ;
        RECT 55.595 162.070 55.865 162.975 ;
        RECT 52.545 161.505 52.740 161.835 ;
        RECT 52.965 161.505 53.220 161.835 ;
        RECT 52.965 161.335 53.135 161.505 ;
        RECT 53.390 161.335 53.560 162.005 ;
        RECT 55.240 161.900 55.410 162.045 ;
        RECT 54.675 161.495 55.005 161.865 ;
        RECT 55.240 161.570 55.525 161.900 ;
        RECT 52.205 161.165 53.135 161.335 ;
        RECT 52.205 161.130 52.380 161.165 ;
        RECT 51.850 160.765 52.380 161.130 ;
        RECT 52.805 160.595 53.135 160.995 ;
        RECT 53.305 160.765 53.560 161.335 ;
        RECT 55.240 161.315 55.410 161.570 ;
        RECT 54.745 161.145 55.410 161.315 ;
        RECT 55.695 161.270 55.865 162.070 ;
        RECT 56.035 162.055 57.705 163.145 ;
        RECT 56.035 161.535 56.785 162.055 ;
        RECT 57.880 161.995 58.140 163.145 ;
        RECT 58.315 162.070 58.570 162.975 ;
        RECT 58.740 162.385 59.070 163.145 ;
        RECT 59.285 162.215 59.455 162.975 ;
        RECT 56.955 161.365 57.705 161.885 ;
        RECT 54.745 160.765 54.915 161.145 ;
        RECT 55.095 160.595 55.425 160.975 ;
        RECT 55.605 160.765 55.865 161.270 ;
        RECT 56.035 160.595 57.705 161.365 ;
        RECT 57.880 160.595 58.140 161.435 ;
        RECT 58.315 161.340 58.485 162.070 ;
        RECT 58.740 162.045 59.455 162.215 ;
        RECT 59.805 162.215 59.975 162.975 ;
        RECT 60.190 162.385 60.520 163.145 ;
        RECT 59.805 162.045 60.520 162.215 ;
        RECT 60.690 162.070 60.945 162.975 ;
        RECT 58.740 161.835 58.910 162.045 ;
        RECT 58.655 161.505 58.910 161.835 ;
        RECT 58.315 160.765 58.570 161.340 ;
        RECT 58.740 161.315 58.910 161.505 ;
        RECT 59.190 161.495 59.545 161.865 ;
        RECT 59.715 161.495 60.070 161.865 ;
        RECT 60.350 161.835 60.520 162.045 ;
        RECT 60.350 161.505 60.605 161.835 ;
        RECT 60.350 161.315 60.520 161.505 ;
        RECT 60.775 161.340 60.945 162.070 ;
        RECT 61.120 161.995 61.380 163.145 ;
        RECT 61.555 161.980 61.845 163.145 ;
        RECT 62.015 162.055 63.225 163.145 ;
        RECT 63.485 162.215 63.655 162.975 ;
        RECT 63.870 162.385 64.200 163.145 ;
        RECT 62.015 161.515 62.535 162.055 ;
        RECT 63.485 162.045 64.200 162.215 ;
        RECT 64.370 162.070 64.625 162.975 ;
        RECT 58.740 161.145 59.455 161.315 ;
        RECT 58.740 160.595 59.070 160.975 ;
        RECT 59.285 160.765 59.455 161.145 ;
        RECT 59.805 161.145 60.520 161.315 ;
        RECT 59.805 160.765 59.975 161.145 ;
        RECT 60.190 160.595 60.520 160.975 ;
        RECT 60.690 160.765 60.945 161.340 ;
        RECT 61.120 160.595 61.380 161.435 ;
        RECT 62.705 161.345 63.225 161.885 ;
        RECT 63.395 161.495 63.750 161.865 ;
        RECT 64.030 161.835 64.200 162.045 ;
        RECT 64.030 161.505 64.285 161.835 ;
        RECT 61.555 160.595 61.845 161.320 ;
        RECT 62.015 160.595 63.225 161.345 ;
        RECT 64.030 161.315 64.200 161.505 ;
        RECT 64.455 161.340 64.625 162.070 ;
        RECT 64.800 161.995 65.060 163.145 ;
        RECT 65.325 162.215 65.495 162.975 ;
        RECT 65.710 162.385 66.040 163.145 ;
        RECT 65.325 162.045 66.040 162.215 ;
        RECT 66.210 162.070 66.465 162.975 ;
        RECT 65.235 161.495 65.590 161.865 ;
        RECT 65.870 161.835 66.040 162.045 ;
        RECT 65.870 161.505 66.125 161.835 ;
        RECT 63.485 161.145 64.200 161.315 ;
        RECT 63.485 160.765 63.655 161.145 ;
        RECT 63.870 160.595 64.200 160.975 ;
        RECT 64.370 160.765 64.625 161.340 ;
        RECT 64.800 160.595 65.060 161.435 ;
        RECT 65.870 161.315 66.040 161.505 ;
        RECT 66.295 161.340 66.465 162.070 ;
        RECT 66.640 161.995 66.900 163.145 ;
        RECT 67.165 162.215 67.335 162.975 ;
        RECT 67.550 162.385 67.880 163.145 ;
        RECT 67.165 162.045 67.880 162.215 ;
        RECT 68.050 162.070 68.305 162.975 ;
        RECT 67.075 161.495 67.430 161.865 ;
        RECT 67.710 161.835 67.880 162.045 ;
        RECT 67.710 161.505 67.965 161.835 ;
        RECT 65.325 161.145 66.040 161.315 ;
        RECT 65.325 160.765 65.495 161.145 ;
        RECT 65.710 160.595 66.040 160.975 ;
        RECT 66.210 160.765 66.465 161.340 ;
        RECT 66.640 160.595 66.900 161.435 ;
        RECT 67.710 161.315 67.880 161.505 ;
        RECT 68.135 161.340 68.305 162.070 ;
        RECT 68.480 161.995 68.740 163.145 ;
        RECT 68.915 162.385 69.430 162.795 ;
        RECT 69.665 162.385 69.835 163.145 ;
        RECT 70.005 162.805 72.035 162.975 ;
        RECT 68.915 161.575 69.255 162.385 ;
        RECT 70.005 162.140 70.175 162.805 ;
        RECT 70.570 162.465 71.695 162.635 ;
        RECT 69.425 161.950 70.175 162.140 ;
        RECT 70.345 162.125 71.355 162.295 ;
        RECT 67.165 161.145 67.880 161.315 ;
        RECT 67.165 160.765 67.335 161.145 ;
        RECT 67.550 160.595 67.880 160.975 ;
        RECT 68.050 160.765 68.305 161.340 ;
        RECT 68.480 160.595 68.740 161.435 ;
        RECT 68.915 161.405 70.145 161.575 ;
        RECT 69.190 160.800 69.435 161.405 ;
        RECT 69.655 160.595 70.165 161.130 ;
        RECT 70.345 160.765 70.535 162.125 ;
        RECT 70.705 161.445 70.980 161.925 ;
        RECT 70.705 161.275 70.985 161.445 ;
        RECT 71.185 161.325 71.355 162.125 ;
        RECT 71.525 161.335 71.695 162.465 ;
        RECT 71.865 161.835 72.035 162.805 ;
        RECT 72.205 162.005 72.375 163.145 ;
        RECT 72.545 162.005 72.880 162.975 ;
        RECT 71.865 161.505 72.060 161.835 ;
        RECT 72.285 161.505 72.540 161.835 ;
        RECT 72.285 161.335 72.455 161.505 ;
        RECT 72.710 161.335 72.880 162.005 ;
        RECT 73.430 162.165 73.685 162.835 ;
        RECT 73.865 162.345 74.150 163.145 ;
        RECT 74.330 162.425 74.660 162.935 ;
        RECT 73.430 161.445 73.610 162.165 ;
        RECT 74.330 161.835 74.580 162.425 ;
        RECT 74.930 162.275 75.100 162.885 ;
        RECT 75.270 162.455 75.600 163.145 ;
        RECT 75.830 162.595 76.070 162.885 ;
        RECT 76.270 162.765 76.690 163.145 ;
        RECT 76.870 162.675 77.500 162.925 ;
        RECT 77.970 162.765 78.300 163.145 ;
        RECT 76.870 162.595 77.040 162.675 ;
        RECT 78.470 162.595 78.640 162.885 ;
        RECT 78.820 162.765 79.200 163.145 ;
        RECT 79.440 162.760 80.270 162.930 ;
        RECT 75.830 162.425 77.040 162.595 ;
        RECT 73.780 161.505 74.580 161.835 ;
        RECT 70.705 160.765 70.980 161.275 ;
        RECT 71.525 161.165 72.455 161.335 ;
        RECT 71.525 161.130 71.700 161.165 ;
        RECT 71.170 160.765 71.700 161.130 ;
        RECT 72.125 160.595 72.455 160.995 ;
        RECT 72.625 160.765 72.880 161.335 ;
        RECT 73.345 161.305 73.610 161.445 ;
        RECT 73.345 161.275 73.685 161.305 ;
        RECT 73.430 160.775 73.685 161.275 ;
        RECT 73.865 160.595 74.150 161.055 ;
        RECT 74.330 160.855 74.580 161.505 ;
        RECT 74.780 162.255 75.100 162.275 ;
        RECT 74.780 162.085 76.700 162.255 ;
        RECT 74.780 161.190 74.970 162.085 ;
        RECT 76.870 161.915 77.040 162.425 ;
        RECT 77.210 162.165 77.730 162.475 ;
        RECT 75.140 161.745 77.040 161.915 ;
        RECT 75.140 161.685 75.470 161.745 ;
        RECT 75.620 161.515 75.950 161.575 ;
        RECT 75.290 161.245 75.950 161.515 ;
        RECT 74.780 160.860 75.100 161.190 ;
        RECT 75.280 160.595 75.940 161.075 ;
        RECT 76.140 160.985 76.310 161.745 ;
        RECT 77.210 161.575 77.390 161.985 ;
        RECT 76.480 161.405 76.810 161.525 ;
        RECT 77.560 161.405 77.730 162.165 ;
        RECT 76.480 161.235 77.730 161.405 ;
        RECT 77.900 162.345 79.270 162.595 ;
        RECT 77.900 161.575 78.090 162.345 ;
        RECT 79.020 162.085 79.270 162.345 ;
        RECT 78.260 161.915 78.510 162.075 ;
        RECT 79.440 161.915 79.610 162.760 ;
        RECT 80.505 162.475 80.675 162.975 ;
        RECT 80.845 162.645 81.175 163.145 ;
        RECT 79.780 162.085 80.280 162.465 ;
        RECT 80.505 162.305 81.200 162.475 ;
        RECT 78.260 161.745 79.610 161.915 ;
        RECT 79.190 161.705 79.610 161.745 ;
        RECT 77.900 161.235 78.320 161.575 ;
        RECT 78.610 161.245 79.020 161.575 ;
        RECT 76.140 160.815 76.990 160.985 ;
        RECT 77.550 160.595 77.870 161.055 ;
        RECT 78.070 160.805 78.320 161.235 ;
        RECT 78.610 160.595 79.020 161.035 ;
        RECT 79.190 160.975 79.360 161.705 ;
        RECT 79.530 161.155 79.880 161.525 ;
        RECT 80.060 161.215 80.280 162.085 ;
        RECT 80.450 161.515 80.860 162.135 ;
        RECT 81.030 161.335 81.200 162.305 ;
        RECT 80.505 161.145 81.200 161.335 ;
        RECT 79.190 160.775 80.205 160.975 ;
        RECT 80.505 160.815 80.675 161.145 ;
        RECT 80.845 160.595 81.175 160.975 ;
        RECT 81.390 160.855 81.615 162.975 ;
        RECT 81.785 162.645 82.115 163.145 ;
        RECT 82.285 162.475 82.455 162.975 ;
        RECT 81.790 162.305 82.455 162.475 ;
        RECT 83.175 162.385 83.690 162.795 ;
        RECT 83.925 162.385 84.095 163.145 ;
        RECT 84.265 162.805 86.295 162.975 ;
        RECT 81.790 161.315 82.020 162.305 ;
        RECT 82.190 161.485 82.540 162.135 ;
        RECT 83.175 161.575 83.515 162.385 ;
        RECT 84.265 162.140 84.435 162.805 ;
        RECT 84.830 162.465 85.955 162.635 ;
        RECT 83.685 161.950 84.435 162.140 ;
        RECT 84.605 162.125 85.615 162.295 ;
        RECT 83.175 161.405 84.405 161.575 ;
        RECT 81.790 161.145 82.455 161.315 ;
        RECT 81.785 160.595 82.115 160.975 ;
        RECT 82.285 160.855 82.455 161.145 ;
        RECT 83.450 160.800 83.695 161.405 ;
        RECT 83.915 160.595 84.425 161.130 ;
        RECT 84.605 160.765 84.795 162.125 ;
        RECT 84.965 161.105 85.240 161.925 ;
        RECT 85.445 161.325 85.615 162.125 ;
        RECT 85.785 161.335 85.955 162.465 ;
        RECT 86.125 161.835 86.295 162.805 ;
        RECT 86.465 162.005 86.635 163.145 ;
        RECT 86.805 162.005 87.140 162.975 ;
        RECT 86.125 161.505 86.320 161.835 ;
        RECT 86.545 161.505 86.800 161.835 ;
        RECT 86.545 161.335 86.715 161.505 ;
        RECT 86.970 161.335 87.140 162.005 ;
        RECT 87.315 161.980 87.605 163.145 ;
        RECT 87.830 162.345 88.130 163.145 ;
        RECT 88.300 162.175 88.630 162.975 ;
        RECT 88.800 162.345 88.970 163.145 ;
        RECT 89.140 162.175 89.470 162.975 ;
        RECT 89.640 162.345 89.810 163.145 ;
        RECT 89.980 162.175 90.310 162.975 ;
        RECT 90.480 162.345 90.650 163.145 ;
        RECT 90.820 162.175 91.150 162.975 ;
        RECT 91.320 162.345 91.575 163.145 ;
        RECT 87.775 162.005 91.745 162.175 ;
        RECT 85.785 161.165 86.715 161.335 ;
        RECT 85.785 161.130 85.960 161.165 ;
        RECT 84.965 160.935 85.245 161.105 ;
        RECT 84.965 160.765 85.240 160.935 ;
        RECT 85.430 160.765 85.960 161.130 ;
        RECT 86.385 160.595 86.715 160.995 ;
        RECT 86.885 160.765 87.140 161.335 ;
        RECT 87.775 161.415 88.095 162.005 ;
        RECT 88.295 161.585 91.150 161.835 ;
        RECT 91.400 161.415 91.745 162.005 ;
        RECT 87.315 160.595 87.605 161.320 ;
        RECT 87.775 161.225 91.745 161.415 ;
        RECT 91.920 162.005 92.255 162.975 ;
        RECT 92.425 162.005 92.595 163.145 ;
        RECT 92.765 162.805 94.795 162.975 ;
        RECT 91.920 161.335 92.090 162.005 ;
        RECT 92.765 161.835 92.935 162.805 ;
        RECT 92.260 161.505 92.515 161.835 ;
        RECT 92.740 161.505 92.935 161.835 ;
        RECT 93.105 162.465 94.230 162.635 ;
        RECT 92.345 161.335 92.515 161.505 ;
        RECT 93.105 161.335 93.275 162.465 ;
        RECT 87.825 160.595 88.130 161.055 ;
        RECT 88.300 160.765 88.630 161.225 ;
        RECT 88.800 160.595 88.970 161.055 ;
        RECT 89.140 160.765 89.470 161.225 ;
        RECT 89.640 160.595 89.810 161.055 ;
        RECT 89.980 160.765 90.310 161.225 ;
        RECT 90.480 160.595 90.650 161.055 ;
        RECT 90.820 160.765 91.150 161.225 ;
        RECT 91.320 160.595 91.575 161.055 ;
        RECT 91.920 160.765 92.175 161.335 ;
        RECT 92.345 161.165 93.275 161.335 ;
        RECT 93.445 162.125 94.455 162.295 ;
        RECT 93.445 161.325 93.615 162.125 ;
        RECT 93.100 161.130 93.275 161.165 ;
        RECT 92.345 160.595 92.675 160.995 ;
        RECT 93.100 160.765 93.630 161.130 ;
        RECT 93.820 161.105 94.095 161.925 ;
        RECT 93.815 160.935 94.095 161.105 ;
        RECT 93.820 160.765 94.095 160.935 ;
        RECT 94.265 160.765 94.455 162.125 ;
        RECT 94.625 162.140 94.795 162.805 ;
        RECT 94.965 162.385 95.135 163.145 ;
        RECT 95.370 162.385 95.885 162.795 ;
        RECT 94.625 161.950 95.375 162.140 ;
        RECT 95.545 161.575 95.885 162.385 ;
        RECT 94.655 161.405 95.885 161.575 ;
        RECT 96.055 162.385 96.570 162.795 ;
        RECT 96.805 162.385 96.975 163.145 ;
        RECT 97.145 162.805 99.175 162.975 ;
        RECT 96.055 161.575 96.395 162.385 ;
        RECT 97.145 162.140 97.315 162.805 ;
        RECT 97.710 162.465 98.835 162.635 ;
        RECT 96.565 161.950 97.315 162.140 ;
        RECT 97.485 162.125 98.495 162.295 ;
        RECT 96.055 161.405 97.285 161.575 ;
        RECT 94.635 160.595 95.145 161.130 ;
        RECT 95.365 160.800 95.610 161.405 ;
        RECT 96.330 160.800 96.575 161.405 ;
        RECT 96.795 160.595 97.305 161.130 ;
        RECT 97.485 160.765 97.675 162.125 ;
        RECT 97.845 161.105 98.120 161.925 ;
        RECT 98.325 161.325 98.495 162.125 ;
        RECT 98.665 161.335 98.835 162.465 ;
        RECT 99.005 161.835 99.175 162.805 ;
        RECT 99.345 162.005 99.515 163.145 ;
        RECT 99.685 162.005 100.020 162.975 ;
        RECT 99.005 161.505 99.200 161.835 ;
        RECT 99.425 161.505 99.680 161.835 ;
        RECT 99.425 161.335 99.595 161.505 ;
        RECT 99.850 161.335 100.020 162.005 ;
        RECT 101.115 162.385 101.630 162.795 ;
        RECT 101.865 162.385 102.035 163.145 ;
        RECT 102.205 162.805 104.235 162.975 ;
        RECT 101.115 161.575 101.455 162.385 ;
        RECT 102.205 162.140 102.375 162.805 ;
        RECT 102.770 162.465 103.895 162.635 ;
        RECT 101.625 161.950 102.375 162.140 ;
        RECT 102.545 162.125 103.555 162.295 ;
        RECT 101.115 161.405 102.345 161.575 ;
        RECT 98.665 161.165 99.595 161.335 ;
        RECT 98.665 161.130 98.840 161.165 ;
        RECT 97.845 160.935 98.125 161.105 ;
        RECT 97.845 160.765 98.120 160.935 ;
        RECT 98.310 160.765 98.840 161.130 ;
        RECT 99.265 160.595 99.595 160.995 ;
        RECT 99.765 160.765 100.020 161.335 ;
        RECT 101.390 160.800 101.635 161.405 ;
        RECT 101.855 160.595 102.365 161.130 ;
        RECT 102.545 160.765 102.735 162.125 ;
        RECT 102.905 161.785 103.180 161.925 ;
        RECT 102.905 161.615 103.185 161.785 ;
        RECT 102.905 160.765 103.180 161.615 ;
        RECT 103.385 161.325 103.555 162.125 ;
        RECT 103.725 161.335 103.895 162.465 ;
        RECT 104.065 161.835 104.235 162.805 ;
        RECT 104.405 162.005 104.575 163.145 ;
        RECT 104.745 162.005 105.080 162.975 ;
        RECT 104.065 161.505 104.260 161.835 ;
        RECT 104.485 161.505 104.740 161.835 ;
        RECT 104.485 161.335 104.655 161.505 ;
        RECT 104.910 161.335 105.080 162.005 ;
        RECT 103.725 161.165 104.655 161.335 ;
        RECT 103.725 161.130 103.900 161.165 ;
        RECT 103.370 160.765 103.900 161.130 ;
        RECT 104.325 160.595 104.655 160.995 ;
        RECT 104.825 160.765 105.080 161.335 ;
        RECT 105.255 162.005 105.640 162.975 ;
        RECT 105.810 162.685 106.135 163.145 ;
        RECT 106.655 162.515 106.935 162.975 ;
        RECT 105.810 162.295 106.935 162.515 ;
        RECT 105.255 161.335 105.535 162.005 ;
        RECT 105.810 161.835 106.260 162.295 ;
        RECT 107.125 162.125 107.525 162.975 ;
        RECT 107.925 162.685 108.195 163.145 ;
        RECT 108.365 162.515 108.650 162.975 ;
        RECT 105.705 161.505 106.260 161.835 ;
        RECT 106.430 161.565 107.525 162.125 ;
        RECT 105.810 161.395 106.260 161.505 ;
        RECT 105.255 160.765 105.640 161.335 ;
        RECT 105.810 161.225 106.935 161.395 ;
        RECT 105.810 160.595 106.135 161.055 ;
        RECT 106.655 160.765 106.935 161.225 ;
        RECT 107.125 160.765 107.525 161.565 ;
        RECT 107.695 162.295 108.650 162.515 ;
        RECT 107.695 161.395 107.905 162.295 ;
        RECT 108.945 162.165 109.275 162.975 ;
        RECT 109.445 162.345 109.685 163.145 ;
        RECT 108.075 161.565 108.765 162.125 ;
        RECT 108.945 161.995 109.660 162.165 ;
        RECT 108.940 161.585 109.320 161.825 ;
        RECT 109.490 161.755 109.660 161.995 ;
        RECT 109.865 162.125 110.035 162.975 ;
        RECT 110.205 162.345 110.535 163.145 ;
        RECT 110.705 162.125 110.875 162.975 ;
        RECT 109.865 161.955 110.875 162.125 ;
        RECT 111.045 161.995 111.375 163.145 ;
        RECT 112.155 162.055 113.365 163.145 ;
        RECT 109.490 161.585 109.990 161.755 ;
        RECT 109.490 161.415 109.660 161.585 ;
        RECT 110.380 161.415 110.875 161.955 ;
        RECT 112.155 161.515 112.675 162.055 ;
        RECT 107.695 161.225 108.650 161.395 ;
        RECT 107.925 160.595 108.195 161.055 ;
        RECT 108.365 160.765 108.650 161.225 ;
        RECT 109.025 161.245 109.660 161.415 ;
        RECT 109.865 161.245 110.875 161.415 ;
        RECT 109.025 160.765 109.195 161.245 ;
        RECT 109.375 160.595 109.615 161.075 ;
        RECT 109.865 160.765 110.035 161.245 ;
        RECT 110.205 160.595 110.535 161.075 ;
        RECT 110.705 160.765 110.875 161.245 ;
        RECT 111.045 160.595 111.375 161.395 ;
        RECT 112.845 161.345 113.365 161.885 ;
        RECT 112.155 160.595 113.365 161.345 ;
        RECT 15.010 160.425 113.450 160.595 ;
        RECT 15.095 159.675 16.305 160.425 ;
        RECT 15.095 159.135 15.615 159.675 ;
        RECT 17.455 159.605 17.665 160.425 ;
        RECT 17.835 159.625 18.165 160.255 ;
        RECT 15.785 158.965 16.305 159.505 ;
        RECT 17.835 159.025 18.085 159.625 ;
        RECT 18.335 159.605 18.565 160.425 ;
        RECT 19.050 159.615 19.295 160.220 ;
        RECT 19.515 159.890 20.025 160.425 ;
        RECT 18.775 159.445 20.005 159.615 ;
        RECT 18.255 159.185 18.585 159.435 ;
        RECT 15.095 157.875 16.305 158.965 ;
        RECT 17.455 157.875 17.665 159.015 ;
        RECT 17.835 158.045 18.165 159.025 ;
        RECT 18.335 157.875 18.565 159.015 ;
        RECT 18.775 158.635 19.115 159.445 ;
        RECT 19.285 158.880 20.035 159.070 ;
        RECT 18.775 158.225 19.290 158.635 ;
        RECT 19.525 157.875 19.695 158.635 ;
        RECT 19.865 158.215 20.035 158.880 ;
        RECT 20.205 158.895 20.395 160.255 ;
        RECT 20.565 159.405 20.840 160.255 ;
        RECT 21.030 159.890 21.560 160.255 ;
        RECT 21.985 160.025 22.315 160.425 ;
        RECT 21.385 159.855 21.560 159.890 ;
        RECT 20.565 159.235 20.845 159.405 ;
        RECT 20.565 159.095 20.840 159.235 ;
        RECT 21.045 158.895 21.215 159.695 ;
        RECT 20.205 158.725 21.215 158.895 ;
        RECT 21.385 159.685 22.315 159.855 ;
        RECT 22.485 159.685 22.740 160.255 ;
        RECT 22.915 159.700 23.205 160.425 ;
        RECT 23.465 159.875 23.635 160.255 ;
        RECT 23.815 160.045 24.145 160.425 ;
        RECT 23.465 159.705 24.130 159.875 ;
        RECT 24.325 159.750 24.585 160.255 ;
        RECT 21.385 158.555 21.555 159.685 ;
        RECT 22.145 159.515 22.315 159.685 ;
        RECT 20.430 158.385 21.555 158.555 ;
        RECT 21.725 159.185 21.920 159.515 ;
        RECT 22.145 159.185 22.400 159.515 ;
        RECT 21.725 158.215 21.895 159.185 ;
        RECT 22.570 159.015 22.740 159.685 ;
        RECT 23.395 159.155 23.725 159.525 ;
        RECT 23.960 159.450 24.130 159.705 ;
        RECT 23.960 159.120 24.245 159.450 ;
        RECT 19.865 158.045 21.895 158.215 ;
        RECT 22.065 157.875 22.235 159.015 ;
        RECT 22.405 158.045 22.740 159.015 ;
        RECT 22.915 157.875 23.205 159.040 ;
        RECT 23.960 158.975 24.130 159.120 ;
        RECT 23.465 158.805 24.130 158.975 ;
        RECT 24.415 158.950 24.585 159.750 ;
        RECT 25.215 159.655 28.725 160.425 ;
        RECT 23.465 158.045 23.635 158.805 ;
        RECT 23.815 157.875 24.145 158.635 ;
        RECT 24.315 158.045 24.585 158.950 ;
        RECT 25.215 158.965 26.905 159.485 ;
        RECT 27.075 159.135 28.725 159.655 ;
        RECT 29.270 159.715 29.525 160.245 ;
        RECT 29.705 159.965 29.990 160.425 ;
        RECT 25.215 157.875 28.725 158.965 ;
        RECT 29.270 158.855 29.450 159.715 ;
        RECT 30.170 159.515 30.420 160.165 ;
        RECT 29.620 159.185 30.420 159.515 ;
        RECT 29.270 158.385 29.525 158.855 ;
        RECT 29.185 158.215 29.525 158.385 ;
        RECT 29.270 158.185 29.525 158.215 ;
        RECT 29.705 157.875 29.990 158.675 ;
        RECT 30.170 158.595 30.420 159.185 ;
        RECT 30.620 159.830 30.940 160.160 ;
        RECT 31.120 159.945 31.780 160.425 ;
        RECT 31.980 160.035 32.830 160.205 ;
        RECT 30.620 158.935 30.810 159.830 ;
        RECT 31.130 159.505 31.790 159.775 ;
        RECT 31.460 159.445 31.790 159.505 ;
        RECT 30.980 159.275 31.310 159.335 ;
        RECT 31.980 159.275 32.150 160.035 ;
        RECT 33.390 159.965 33.710 160.425 ;
        RECT 33.910 159.785 34.160 160.215 ;
        RECT 34.450 159.985 34.860 160.425 ;
        RECT 35.030 160.045 36.045 160.245 ;
        RECT 32.320 159.615 33.570 159.785 ;
        RECT 32.320 159.495 32.650 159.615 ;
        RECT 30.980 159.105 32.880 159.275 ;
        RECT 30.620 158.765 32.540 158.935 ;
        RECT 30.620 158.745 30.940 158.765 ;
        RECT 30.170 158.085 30.500 158.595 ;
        RECT 30.770 158.135 30.940 158.745 ;
        RECT 32.710 158.595 32.880 159.105 ;
        RECT 33.050 159.035 33.230 159.445 ;
        RECT 33.400 158.855 33.570 159.615 ;
        RECT 31.110 157.875 31.440 158.565 ;
        RECT 31.670 158.425 32.880 158.595 ;
        RECT 33.050 158.545 33.570 158.855 ;
        RECT 33.740 159.445 34.160 159.785 ;
        RECT 34.450 159.445 34.860 159.775 ;
        RECT 33.740 158.675 33.930 159.445 ;
        RECT 35.030 159.315 35.200 160.045 ;
        RECT 36.345 159.875 36.515 160.205 ;
        RECT 36.685 160.045 37.015 160.425 ;
        RECT 35.370 159.495 35.720 159.865 ;
        RECT 35.030 159.275 35.450 159.315 ;
        RECT 34.100 159.105 35.450 159.275 ;
        RECT 34.100 158.945 34.350 159.105 ;
        RECT 34.860 158.675 35.110 158.935 ;
        RECT 33.740 158.425 35.110 158.675 ;
        RECT 31.670 158.135 31.910 158.425 ;
        RECT 32.710 158.345 32.880 158.425 ;
        RECT 32.110 157.875 32.530 158.255 ;
        RECT 32.710 158.095 33.340 158.345 ;
        RECT 33.810 157.875 34.140 158.255 ;
        RECT 34.310 158.135 34.480 158.425 ;
        RECT 35.280 158.260 35.450 159.105 ;
        RECT 35.900 158.935 36.120 159.805 ;
        RECT 36.345 159.685 37.040 159.875 ;
        RECT 35.620 158.555 36.120 158.935 ;
        RECT 36.290 158.885 36.700 159.505 ;
        RECT 36.870 158.715 37.040 159.685 ;
        RECT 36.345 158.545 37.040 158.715 ;
        RECT 34.660 157.875 35.040 158.255 ;
        RECT 35.280 158.090 36.110 158.260 ;
        RECT 36.345 158.045 36.515 158.545 ;
        RECT 36.685 157.875 37.015 158.375 ;
        RECT 37.230 158.045 37.455 160.165 ;
        RECT 37.625 160.045 37.955 160.425 ;
        RECT 38.125 159.875 38.295 160.165 ;
        RECT 37.630 159.705 38.295 159.875 ;
        RECT 38.555 159.750 38.815 160.255 ;
        RECT 38.995 160.045 39.325 160.425 ;
        RECT 39.505 159.875 39.675 160.255 ;
        RECT 37.630 158.715 37.860 159.705 ;
        RECT 38.030 158.885 38.380 159.535 ;
        RECT 38.555 158.950 38.725 159.750 ;
        RECT 39.010 159.705 39.675 159.875 ;
        RECT 39.010 159.450 39.180 159.705 ;
        RECT 39.935 159.675 41.145 160.425 ;
        RECT 38.895 159.120 39.180 159.450 ;
        RECT 39.415 159.155 39.745 159.525 ;
        RECT 39.010 158.975 39.180 159.120 ;
        RECT 37.630 158.545 38.295 158.715 ;
        RECT 37.625 157.875 37.955 158.375 ;
        RECT 38.125 158.045 38.295 158.545 ;
        RECT 38.555 158.045 38.825 158.950 ;
        RECT 39.010 158.805 39.675 158.975 ;
        RECT 38.995 157.875 39.325 158.635 ;
        RECT 39.505 158.045 39.675 158.805 ;
        RECT 39.935 158.965 40.455 159.505 ;
        RECT 40.625 159.135 41.145 159.675 ;
        RECT 41.315 159.625 41.655 160.255 ;
        RECT 41.825 159.625 42.075 160.425 ;
        RECT 42.265 159.775 42.595 160.255 ;
        RECT 42.765 159.965 42.990 160.425 ;
        RECT 43.160 159.775 43.490 160.255 ;
        RECT 41.315 159.015 41.490 159.625 ;
        RECT 42.265 159.605 43.490 159.775 ;
        RECT 44.120 159.645 44.620 160.255 ;
        RECT 45.200 159.645 45.700 160.255 ;
        RECT 41.660 159.265 42.355 159.435 ;
        RECT 42.185 159.015 42.355 159.265 ;
        RECT 42.530 159.235 42.950 159.435 ;
        RECT 43.120 159.235 43.450 159.435 ;
        RECT 43.620 159.235 43.950 159.435 ;
        RECT 44.120 159.015 44.290 159.645 ;
        RECT 44.475 159.185 44.825 159.435 ;
        RECT 44.995 159.185 45.345 159.435 ;
        RECT 45.530 159.015 45.700 159.645 ;
        RECT 46.330 159.775 46.660 160.255 ;
        RECT 46.830 159.965 47.055 160.425 ;
        RECT 47.225 159.775 47.555 160.255 ;
        RECT 46.330 159.605 47.555 159.775 ;
        RECT 47.745 159.625 47.995 160.425 ;
        RECT 48.165 159.625 48.505 160.255 ;
        RECT 48.675 159.700 48.965 160.425 ;
        RECT 49.135 159.675 50.345 160.425 ;
        RECT 45.870 159.235 46.200 159.435 ;
        RECT 46.370 159.235 46.700 159.435 ;
        RECT 46.870 159.235 47.290 159.435 ;
        RECT 47.465 159.265 48.160 159.435 ;
        RECT 47.465 159.015 47.635 159.265 ;
        RECT 48.330 159.015 48.505 159.625 ;
        RECT 39.935 157.875 41.145 158.965 ;
        RECT 41.315 158.045 41.655 159.015 ;
        RECT 41.825 157.875 41.995 159.015 ;
        RECT 42.185 158.845 44.620 159.015 ;
        RECT 42.265 157.875 42.515 158.675 ;
        RECT 43.160 158.045 43.490 158.845 ;
        RECT 43.790 157.875 44.120 158.675 ;
        RECT 44.290 158.045 44.620 158.845 ;
        RECT 45.200 158.845 47.635 159.015 ;
        RECT 45.200 158.045 45.530 158.845 ;
        RECT 45.700 157.875 46.030 158.675 ;
        RECT 46.330 158.045 46.660 158.845 ;
        RECT 47.305 157.875 47.555 158.675 ;
        RECT 47.825 157.875 47.995 159.015 ;
        RECT 48.165 158.045 48.505 159.015 ;
        RECT 48.675 157.875 48.965 159.040 ;
        RECT 49.135 158.965 49.655 159.505 ;
        RECT 49.825 159.135 50.345 159.675 ;
        RECT 50.630 159.795 50.915 160.255 ;
        RECT 51.085 159.965 51.355 160.425 ;
        RECT 50.630 159.625 51.585 159.795 ;
        RECT 49.135 157.875 50.345 158.965 ;
        RECT 50.515 158.895 51.205 159.455 ;
        RECT 51.375 158.725 51.585 159.625 ;
        RECT 50.630 158.505 51.585 158.725 ;
        RECT 51.755 159.455 52.155 160.255 ;
        RECT 52.345 159.795 52.625 160.255 ;
        RECT 53.145 159.965 53.470 160.425 ;
        RECT 52.345 159.625 53.470 159.795 ;
        RECT 53.640 159.685 54.025 160.255 ;
        RECT 53.020 159.515 53.470 159.625 ;
        RECT 51.755 158.895 52.850 159.455 ;
        RECT 53.020 159.185 53.575 159.515 ;
        RECT 50.630 158.045 50.915 158.505 ;
        RECT 51.085 157.875 51.355 158.335 ;
        RECT 51.755 158.045 52.155 158.895 ;
        RECT 53.020 158.725 53.470 159.185 ;
        RECT 53.745 159.015 54.025 159.685 ;
        RECT 54.345 159.625 54.675 160.425 ;
        RECT 54.845 159.775 55.015 160.255 ;
        RECT 55.185 159.945 55.515 160.425 ;
        RECT 55.685 159.775 55.855 160.255 ;
        RECT 56.105 159.945 56.345 160.425 ;
        RECT 56.525 159.775 56.695 160.255 ;
        RECT 54.845 159.605 55.855 159.775 ;
        RECT 56.060 159.605 56.695 159.775 ;
        RECT 57.015 159.605 57.225 160.425 ;
        RECT 57.395 159.625 57.725 160.255 ;
        RECT 54.845 159.575 55.345 159.605 ;
        RECT 54.845 159.065 55.340 159.575 ;
        RECT 56.060 159.435 56.230 159.605 ;
        RECT 55.730 159.265 56.230 159.435 ;
        RECT 52.345 158.505 53.470 158.725 ;
        RECT 52.345 158.045 52.625 158.505 ;
        RECT 53.145 157.875 53.470 158.335 ;
        RECT 53.640 158.045 54.025 159.015 ;
        RECT 54.345 157.875 54.675 159.025 ;
        RECT 54.845 158.895 55.855 159.065 ;
        RECT 54.845 158.045 55.015 158.895 ;
        RECT 55.185 157.875 55.515 158.675 ;
        RECT 55.685 158.045 55.855 158.895 ;
        RECT 56.060 159.025 56.230 159.265 ;
        RECT 56.400 159.195 56.780 159.435 ;
        RECT 57.395 159.025 57.645 159.625 ;
        RECT 57.895 159.605 58.125 160.425 ;
        RECT 58.340 159.585 58.600 160.425 ;
        RECT 58.775 159.680 59.030 160.255 ;
        RECT 59.200 160.045 59.530 160.425 ;
        RECT 59.745 159.875 59.915 160.255 ;
        RECT 59.200 159.705 59.915 159.875 ;
        RECT 57.815 159.185 58.145 159.435 ;
        RECT 56.060 158.855 56.775 159.025 ;
        RECT 56.035 157.875 56.275 158.675 ;
        RECT 56.445 158.045 56.775 158.855 ;
        RECT 57.015 157.875 57.225 159.015 ;
        RECT 57.395 158.045 57.725 159.025 ;
        RECT 57.895 157.875 58.125 159.015 ;
        RECT 58.340 157.875 58.600 159.025 ;
        RECT 58.775 158.950 58.945 159.680 ;
        RECT 59.200 159.515 59.370 159.705 ;
        RECT 60.180 159.585 60.440 160.425 ;
        RECT 60.615 159.680 60.870 160.255 ;
        RECT 61.040 160.045 61.370 160.425 ;
        RECT 61.585 159.875 61.755 160.255 ;
        RECT 61.040 159.705 61.755 159.875 ;
        RECT 59.115 159.185 59.370 159.515 ;
        RECT 59.200 158.975 59.370 159.185 ;
        RECT 59.650 159.155 60.005 159.525 ;
        RECT 58.775 158.045 59.030 158.950 ;
        RECT 59.200 158.805 59.915 158.975 ;
        RECT 59.200 157.875 59.530 158.635 ;
        RECT 59.745 158.045 59.915 158.805 ;
        RECT 60.180 157.875 60.440 159.025 ;
        RECT 60.615 158.950 60.785 159.680 ;
        RECT 61.040 159.515 61.210 159.705 ;
        RECT 62.480 159.585 62.740 160.425 ;
        RECT 62.915 159.680 63.170 160.255 ;
        RECT 63.340 160.045 63.670 160.425 ;
        RECT 63.885 159.875 64.055 160.255 ;
        RECT 63.340 159.705 64.055 159.875 ;
        RECT 60.955 159.185 61.210 159.515 ;
        RECT 61.040 158.975 61.210 159.185 ;
        RECT 61.490 159.155 61.845 159.525 ;
        RECT 60.615 158.045 60.870 158.950 ;
        RECT 61.040 158.805 61.755 158.975 ;
        RECT 61.040 157.875 61.370 158.635 ;
        RECT 61.585 158.045 61.755 158.805 ;
        RECT 62.480 157.875 62.740 159.025 ;
        RECT 62.915 158.950 63.085 159.680 ;
        RECT 63.340 159.515 63.510 159.705 ;
        RECT 65.440 159.645 65.940 160.255 ;
        RECT 63.255 159.185 63.510 159.515 ;
        RECT 63.340 158.975 63.510 159.185 ;
        RECT 63.790 159.155 64.145 159.525 ;
        RECT 65.235 159.185 65.585 159.435 ;
        RECT 65.770 159.015 65.940 159.645 ;
        RECT 66.570 159.775 66.900 160.255 ;
        RECT 67.070 159.965 67.295 160.425 ;
        RECT 67.465 159.775 67.795 160.255 ;
        RECT 66.570 159.605 67.795 159.775 ;
        RECT 67.985 159.625 68.235 160.425 ;
        RECT 68.405 159.625 68.745 160.255 ;
        RECT 66.110 159.235 66.440 159.435 ;
        RECT 66.610 159.235 66.940 159.435 ;
        RECT 67.110 159.235 67.530 159.435 ;
        RECT 67.705 159.265 68.400 159.435 ;
        RECT 67.705 159.015 67.875 159.265 ;
        RECT 68.570 159.015 68.745 159.625 ;
        RECT 62.915 158.045 63.170 158.950 ;
        RECT 63.340 158.805 64.055 158.975 ;
        RECT 63.340 157.875 63.670 158.635 ;
        RECT 63.885 158.045 64.055 158.805 ;
        RECT 65.440 158.845 67.875 159.015 ;
        RECT 65.440 158.045 65.770 158.845 ;
        RECT 65.940 157.875 66.270 158.675 ;
        RECT 66.570 158.045 66.900 158.845 ;
        RECT 67.545 157.875 67.795 158.675 ;
        RECT 68.065 157.875 68.235 159.015 ;
        RECT 68.405 158.045 68.745 159.015 ;
        RECT 68.915 159.625 69.255 160.255 ;
        RECT 69.425 159.625 69.675 160.425 ;
        RECT 69.865 159.775 70.195 160.255 ;
        RECT 70.365 159.965 70.590 160.425 ;
        RECT 70.760 159.775 71.090 160.255 ;
        RECT 68.915 159.015 69.090 159.625 ;
        RECT 69.865 159.605 71.090 159.775 ;
        RECT 71.720 159.645 72.220 160.255 ;
        RECT 72.595 159.655 74.265 160.425 ;
        RECT 74.435 159.700 74.725 160.425 ;
        RECT 74.895 159.655 78.405 160.425 ;
        RECT 78.665 159.875 78.835 160.255 ;
        RECT 79.015 160.045 79.345 160.425 ;
        RECT 78.665 159.705 79.330 159.875 ;
        RECT 79.525 159.750 79.785 160.255 ;
        RECT 69.260 159.265 69.955 159.435 ;
        RECT 69.785 159.015 69.955 159.265 ;
        RECT 70.130 159.235 70.550 159.435 ;
        RECT 70.720 159.235 71.050 159.435 ;
        RECT 71.220 159.235 71.550 159.435 ;
        RECT 71.720 159.015 71.890 159.645 ;
        RECT 72.075 159.185 72.425 159.435 ;
        RECT 68.915 158.045 69.255 159.015 ;
        RECT 69.425 157.875 69.595 159.015 ;
        RECT 69.785 158.845 72.220 159.015 ;
        RECT 69.865 157.875 70.115 158.675 ;
        RECT 70.760 158.045 71.090 158.845 ;
        RECT 71.390 157.875 71.720 158.675 ;
        RECT 71.890 158.045 72.220 158.845 ;
        RECT 72.595 158.965 73.345 159.485 ;
        RECT 73.515 159.135 74.265 159.655 ;
        RECT 72.595 157.875 74.265 158.965 ;
        RECT 74.435 157.875 74.725 159.040 ;
        RECT 74.895 158.965 76.585 159.485 ;
        RECT 76.755 159.135 78.405 159.655 ;
        RECT 78.595 159.155 78.925 159.525 ;
        RECT 79.160 159.450 79.330 159.705 ;
        RECT 79.160 159.120 79.445 159.450 ;
        RECT 79.160 158.975 79.330 159.120 ;
        RECT 74.895 157.875 78.405 158.965 ;
        RECT 78.665 158.805 79.330 158.975 ;
        RECT 79.615 158.950 79.785 159.750 ;
        RECT 80.455 159.605 80.685 160.425 ;
        RECT 80.855 159.625 81.185 160.255 ;
        RECT 80.435 159.185 80.765 159.435 ;
        RECT 80.935 159.025 81.185 159.625 ;
        RECT 81.355 159.605 81.565 160.425 ;
        RECT 81.795 159.915 82.100 160.425 ;
        RECT 81.795 159.185 82.110 159.745 ;
        RECT 82.280 159.435 82.530 160.245 ;
        RECT 82.700 159.900 82.960 160.425 ;
        RECT 83.140 159.435 83.390 160.245 ;
        RECT 83.560 159.865 83.820 160.425 ;
        RECT 83.990 159.775 84.250 160.230 ;
        RECT 84.420 159.945 84.680 160.425 ;
        RECT 84.850 159.775 85.110 160.230 ;
        RECT 85.280 159.945 85.540 160.425 ;
        RECT 85.710 159.775 85.970 160.230 ;
        RECT 86.140 159.945 86.385 160.425 ;
        RECT 86.555 159.775 86.830 160.230 ;
        RECT 87.000 159.945 87.245 160.425 ;
        RECT 87.415 159.775 87.675 160.230 ;
        RECT 87.855 159.945 88.105 160.425 ;
        RECT 88.275 159.775 88.535 160.230 ;
        RECT 88.715 159.945 88.965 160.425 ;
        RECT 89.135 159.775 89.395 160.230 ;
        RECT 89.575 159.945 89.835 160.425 ;
        RECT 90.005 159.775 90.265 160.230 ;
        RECT 90.435 159.945 90.735 160.425 ;
        RECT 91.110 159.795 91.395 160.255 ;
        RECT 91.565 159.965 91.835 160.425 ;
        RECT 83.990 159.605 90.735 159.775 ;
        RECT 91.110 159.625 92.065 159.795 ;
        RECT 82.280 159.185 89.400 159.435 ;
        RECT 78.665 158.045 78.835 158.805 ;
        RECT 79.015 157.875 79.345 158.635 ;
        RECT 79.515 158.045 79.785 158.950 ;
        RECT 80.455 157.875 80.685 159.015 ;
        RECT 80.855 158.045 81.185 159.025 ;
        RECT 81.355 157.875 81.565 159.015 ;
        RECT 81.805 157.875 82.100 158.685 ;
        RECT 82.280 158.045 82.525 159.185 ;
        RECT 82.700 157.875 82.960 158.685 ;
        RECT 83.140 158.050 83.390 159.185 ;
        RECT 89.570 159.015 90.735 159.605 ;
        RECT 83.990 158.790 90.735 159.015 ;
        RECT 90.995 158.895 91.685 159.455 ;
        RECT 83.990 158.775 89.395 158.790 ;
        RECT 83.560 157.880 83.820 158.675 ;
        RECT 83.990 158.050 84.250 158.775 ;
        RECT 84.420 157.880 84.680 158.605 ;
        RECT 84.850 158.050 85.110 158.775 ;
        RECT 85.280 157.880 85.540 158.605 ;
        RECT 85.710 158.050 85.970 158.775 ;
        RECT 86.140 157.880 86.400 158.605 ;
        RECT 86.570 158.050 86.830 158.775 ;
        RECT 87.000 157.880 87.245 158.605 ;
        RECT 87.415 158.050 87.675 158.775 ;
        RECT 87.860 157.880 88.105 158.605 ;
        RECT 88.275 158.050 88.535 158.775 ;
        RECT 88.720 157.880 88.965 158.605 ;
        RECT 89.135 158.050 89.395 158.775 ;
        RECT 89.580 157.880 89.835 158.605 ;
        RECT 90.005 158.050 90.295 158.790 ;
        RECT 91.855 158.725 92.065 159.625 ;
        RECT 83.560 157.875 89.835 157.880 ;
        RECT 90.465 157.875 90.735 158.620 ;
        RECT 91.110 158.505 92.065 158.725 ;
        RECT 92.235 159.455 92.635 160.255 ;
        RECT 92.825 159.795 93.105 160.255 ;
        RECT 93.625 159.965 93.950 160.425 ;
        RECT 92.825 159.625 93.950 159.795 ;
        RECT 94.120 159.685 94.505 160.255 ;
        RECT 93.500 159.515 93.950 159.625 ;
        RECT 92.235 158.895 93.330 159.455 ;
        RECT 93.500 159.185 94.055 159.515 ;
        RECT 91.110 158.045 91.395 158.505 ;
        RECT 91.565 157.875 91.835 158.335 ;
        RECT 92.235 158.045 92.635 158.895 ;
        RECT 93.500 158.725 93.950 159.185 ;
        RECT 94.225 159.015 94.505 159.685 ;
        RECT 94.675 159.655 96.345 160.425 ;
        RECT 92.825 158.505 93.950 158.725 ;
        RECT 92.825 158.045 93.105 158.505 ;
        RECT 93.625 157.875 93.950 158.335 ;
        RECT 94.120 158.045 94.505 159.015 ;
        RECT 94.675 158.965 95.425 159.485 ;
        RECT 95.595 159.135 96.345 159.655 ;
        RECT 96.515 159.625 96.855 160.255 ;
        RECT 97.025 159.625 97.275 160.425 ;
        RECT 97.465 159.775 97.795 160.255 ;
        RECT 97.965 159.965 98.190 160.425 ;
        RECT 98.360 159.775 98.690 160.255 ;
        RECT 96.515 159.015 96.690 159.625 ;
        RECT 97.465 159.605 98.690 159.775 ;
        RECT 99.320 159.645 99.820 160.255 ;
        RECT 100.195 159.700 100.485 160.425 ;
        RECT 96.860 159.265 97.555 159.435 ;
        RECT 97.385 159.015 97.555 159.265 ;
        RECT 97.730 159.235 98.150 159.435 ;
        RECT 98.320 159.235 98.650 159.435 ;
        RECT 98.820 159.235 99.150 159.435 ;
        RECT 99.320 159.015 99.490 159.645 ;
        RECT 100.655 159.625 100.995 160.255 ;
        RECT 101.165 159.625 101.415 160.425 ;
        RECT 101.605 159.775 101.935 160.255 ;
        RECT 102.105 159.965 102.330 160.425 ;
        RECT 102.500 159.775 102.830 160.255 ;
        RECT 99.675 159.185 100.025 159.435 ;
        RECT 100.655 159.065 100.830 159.625 ;
        RECT 101.605 159.605 102.830 159.775 ;
        RECT 103.460 159.645 103.960 160.255 ;
        RECT 104.335 159.685 104.720 160.255 ;
        RECT 104.890 159.965 105.215 160.425 ;
        RECT 105.735 159.795 106.015 160.255 ;
        RECT 101.000 159.265 101.695 159.435 ;
        RECT 94.675 157.875 96.345 158.965 ;
        RECT 96.515 158.045 96.855 159.015 ;
        RECT 97.025 157.875 97.195 159.015 ;
        RECT 97.385 158.845 99.820 159.015 ;
        RECT 97.465 157.875 97.715 158.675 ;
        RECT 98.360 158.045 98.690 158.845 ;
        RECT 98.990 157.875 99.320 158.675 ;
        RECT 99.490 158.045 99.820 158.845 ;
        RECT 100.195 157.875 100.485 159.040 ;
        RECT 100.655 159.015 100.885 159.065 ;
        RECT 101.525 159.015 101.695 159.265 ;
        RECT 101.870 159.235 102.290 159.435 ;
        RECT 102.460 159.235 102.790 159.435 ;
        RECT 102.960 159.235 103.290 159.435 ;
        RECT 103.460 159.015 103.630 159.645 ;
        RECT 103.815 159.185 104.165 159.435 ;
        RECT 104.335 159.015 104.615 159.685 ;
        RECT 104.890 159.625 106.015 159.795 ;
        RECT 104.890 159.515 105.340 159.625 ;
        RECT 104.785 159.185 105.340 159.515 ;
        RECT 106.205 159.455 106.605 160.255 ;
        RECT 107.005 159.965 107.275 160.425 ;
        RECT 107.445 159.795 107.730 160.255 ;
        RECT 100.655 158.045 100.995 159.015 ;
        RECT 101.165 157.875 101.335 159.015 ;
        RECT 101.525 158.845 103.960 159.015 ;
        RECT 101.605 157.875 101.855 158.675 ;
        RECT 102.500 158.045 102.830 158.845 ;
        RECT 103.130 157.875 103.460 158.675 ;
        RECT 103.630 158.045 103.960 158.845 ;
        RECT 104.335 158.045 104.720 159.015 ;
        RECT 104.890 158.725 105.340 159.185 ;
        RECT 105.510 158.895 106.605 159.455 ;
        RECT 104.890 158.505 106.015 158.725 ;
        RECT 104.890 157.875 105.215 158.335 ;
        RECT 105.735 158.045 106.015 158.505 ;
        RECT 106.205 158.045 106.605 158.895 ;
        RECT 106.775 159.625 107.730 159.795 ;
        RECT 108.165 159.625 108.495 160.425 ;
        RECT 108.665 159.775 108.835 160.255 ;
        RECT 109.005 159.945 109.335 160.425 ;
        RECT 109.505 159.775 109.675 160.255 ;
        RECT 109.925 159.945 110.165 160.425 ;
        RECT 110.345 159.775 110.515 160.255 ;
        RECT 106.775 158.725 106.985 159.625 ;
        RECT 108.665 159.605 109.675 159.775 ;
        RECT 109.880 159.605 110.515 159.775 ;
        RECT 110.815 159.605 111.045 160.425 ;
        RECT 111.215 159.625 111.545 160.255 ;
        RECT 107.155 158.895 107.845 159.455 ;
        RECT 108.665 159.405 109.160 159.605 ;
        RECT 109.880 159.435 110.050 159.605 ;
        RECT 108.665 159.235 109.165 159.405 ;
        RECT 109.550 159.265 110.050 159.435 ;
        RECT 108.665 159.065 109.160 159.235 ;
        RECT 106.775 158.505 107.730 158.725 ;
        RECT 107.005 157.875 107.275 158.335 ;
        RECT 107.445 158.045 107.730 158.505 ;
        RECT 108.165 157.875 108.495 159.025 ;
        RECT 108.665 158.895 109.675 159.065 ;
        RECT 108.665 158.045 108.835 158.895 ;
        RECT 109.005 157.875 109.335 158.675 ;
        RECT 109.505 158.045 109.675 158.895 ;
        RECT 109.880 159.025 110.050 159.265 ;
        RECT 110.220 159.195 110.600 159.435 ;
        RECT 110.795 159.185 111.125 159.435 ;
        RECT 111.295 159.025 111.545 159.625 ;
        RECT 111.715 159.605 111.925 160.425 ;
        RECT 112.155 159.675 113.365 160.425 ;
        RECT 109.880 158.855 110.595 159.025 ;
        RECT 109.855 157.875 110.095 158.675 ;
        RECT 110.265 158.045 110.595 158.855 ;
        RECT 110.815 157.875 111.045 159.015 ;
        RECT 111.215 158.045 111.545 159.025 ;
        RECT 111.715 157.875 111.925 159.015 ;
        RECT 112.155 158.965 112.675 159.505 ;
        RECT 112.845 159.135 113.365 159.675 ;
        RECT 112.155 157.875 113.365 158.965 ;
        RECT 15.010 157.705 113.450 157.875 ;
        RECT 15.095 156.615 16.305 157.705 ;
        RECT 16.850 156.725 17.105 157.395 ;
        RECT 17.285 156.905 17.570 157.705 ;
        RECT 17.750 156.985 18.080 157.495 ;
        RECT 16.850 156.685 17.030 156.725 ;
        RECT 15.095 155.905 15.615 156.445 ;
        RECT 15.785 156.075 16.305 156.615 ;
        RECT 16.765 156.515 17.030 156.685 ;
        RECT 15.095 155.155 16.305 155.905 ;
        RECT 16.850 155.865 17.030 156.515 ;
        RECT 17.750 156.395 18.000 156.985 ;
        RECT 18.350 156.835 18.520 157.445 ;
        RECT 18.690 157.015 19.020 157.705 ;
        RECT 19.250 157.155 19.490 157.445 ;
        RECT 19.690 157.325 20.110 157.705 ;
        RECT 20.290 157.235 20.920 157.485 ;
        RECT 21.390 157.325 21.720 157.705 ;
        RECT 20.290 157.155 20.460 157.235 ;
        RECT 21.890 157.155 22.060 157.445 ;
        RECT 22.240 157.325 22.620 157.705 ;
        RECT 22.860 157.320 23.690 157.490 ;
        RECT 19.250 156.985 20.460 157.155 ;
        RECT 17.200 156.065 18.000 156.395 ;
        RECT 16.850 155.335 17.105 155.865 ;
        RECT 17.285 155.155 17.570 155.615 ;
        RECT 17.750 155.415 18.000 156.065 ;
        RECT 18.200 156.815 18.520 156.835 ;
        RECT 18.200 156.645 20.120 156.815 ;
        RECT 18.200 155.750 18.390 156.645 ;
        RECT 20.290 156.475 20.460 156.985 ;
        RECT 20.630 156.725 21.150 157.035 ;
        RECT 18.560 156.305 20.460 156.475 ;
        RECT 18.560 156.245 18.890 156.305 ;
        RECT 19.040 156.075 19.370 156.135 ;
        RECT 18.710 155.805 19.370 156.075 ;
        RECT 18.200 155.420 18.520 155.750 ;
        RECT 18.700 155.155 19.360 155.635 ;
        RECT 19.560 155.545 19.730 156.305 ;
        RECT 20.630 156.135 20.810 156.545 ;
        RECT 19.900 155.965 20.230 156.085 ;
        RECT 20.980 155.965 21.150 156.725 ;
        RECT 19.900 155.795 21.150 155.965 ;
        RECT 21.320 156.905 22.690 157.155 ;
        RECT 21.320 156.135 21.510 156.905 ;
        RECT 22.440 156.645 22.690 156.905 ;
        RECT 21.680 156.475 21.930 156.635 ;
        RECT 22.860 156.475 23.030 157.320 ;
        RECT 23.925 157.035 24.095 157.535 ;
        RECT 24.265 157.205 24.595 157.705 ;
        RECT 23.200 156.645 23.700 157.025 ;
        RECT 23.925 156.865 24.620 157.035 ;
        RECT 21.680 156.305 23.030 156.475 ;
        RECT 22.610 156.265 23.030 156.305 ;
        RECT 21.320 155.795 21.740 156.135 ;
        RECT 22.030 155.805 22.440 156.135 ;
        RECT 19.560 155.375 20.410 155.545 ;
        RECT 20.970 155.155 21.290 155.615 ;
        RECT 21.490 155.365 21.740 155.795 ;
        RECT 22.030 155.155 22.440 155.595 ;
        RECT 22.610 155.535 22.780 156.265 ;
        RECT 22.950 155.715 23.300 156.085 ;
        RECT 23.480 155.775 23.700 156.645 ;
        RECT 23.870 156.075 24.280 156.695 ;
        RECT 24.450 155.895 24.620 156.865 ;
        RECT 23.925 155.705 24.620 155.895 ;
        RECT 22.610 155.335 23.625 155.535 ;
        RECT 23.925 155.375 24.095 155.705 ;
        RECT 24.265 155.155 24.595 155.535 ;
        RECT 24.810 155.415 25.035 157.535 ;
        RECT 25.205 157.205 25.535 157.705 ;
        RECT 25.705 157.035 25.875 157.535 ;
        RECT 25.210 156.865 25.875 157.035 ;
        RECT 25.210 155.875 25.440 156.865 ;
        RECT 25.610 156.045 25.960 156.695 ;
        RECT 26.595 156.615 28.265 157.705 ;
        RECT 26.595 156.095 27.345 156.615 ;
        RECT 28.435 156.565 28.775 157.535 ;
        RECT 28.945 156.565 29.115 157.705 ;
        RECT 29.385 156.905 29.635 157.705 ;
        RECT 30.280 156.735 30.610 157.535 ;
        RECT 30.910 156.905 31.240 157.705 ;
        RECT 31.410 156.735 31.740 157.535 ;
        RECT 29.305 156.565 31.740 156.735 ;
        RECT 32.320 156.735 32.650 157.535 ;
        RECT 32.820 156.905 33.150 157.705 ;
        RECT 33.450 156.735 33.780 157.535 ;
        RECT 34.425 156.905 34.675 157.705 ;
        RECT 32.320 156.565 34.755 156.735 ;
        RECT 34.945 156.565 35.115 157.705 ;
        RECT 35.285 156.565 35.625 157.535 ;
        RECT 27.515 155.925 28.265 156.445 ;
        RECT 25.210 155.705 25.875 155.875 ;
        RECT 25.205 155.155 25.535 155.535 ;
        RECT 25.705 155.415 25.875 155.705 ;
        RECT 26.595 155.155 28.265 155.925 ;
        RECT 28.435 155.955 28.610 156.565 ;
        RECT 29.305 156.315 29.475 156.565 ;
        RECT 28.780 156.145 29.475 156.315 ;
        RECT 29.650 156.145 30.070 156.345 ;
        RECT 30.240 156.145 30.570 156.345 ;
        RECT 30.740 156.145 31.070 156.345 ;
        RECT 28.435 155.325 28.775 155.955 ;
        RECT 28.945 155.155 29.195 155.955 ;
        RECT 29.385 155.805 30.610 155.975 ;
        RECT 29.385 155.325 29.715 155.805 ;
        RECT 29.885 155.155 30.110 155.615 ;
        RECT 30.280 155.325 30.610 155.805 ;
        RECT 31.240 155.935 31.410 156.565 ;
        RECT 31.595 156.145 31.945 156.395 ;
        RECT 32.115 156.145 32.465 156.395 ;
        RECT 32.650 155.935 32.820 156.565 ;
        RECT 32.990 156.145 33.320 156.345 ;
        RECT 33.490 156.145 33.820 156.345 ;
        RECT 33.990 156.145 34.410 156.345 ;
        RECT 34.585 156.315 34.755 156.565 ;
        RECT 34.585 156.145 35.280 156.315 ;
        RECT 31.240 155.325 31.740 155.935 ;
        RECT 32.320 155.325 32.820 155.935 ;
        RECT 33.450 155.805 34.675 155.975 ;
        RECT 35.450 155.955 35.625 156.565 ;
        RECT 35.795 156.540 36.085 157.705 ;
        RECT 37.380 156.735 37.710 157.535 ;
        RECT 37.880 156.905 38.210 157.705 ;
        RECT 38.510 156.735 38.840 157.535 ;
        RECT 39.485 156.905 39.735 157.705 ;
        RECT 37.380 156.565 39.815 156.735 ;
        RECT 40.005 156.565 40.175 157.705 ;
        RECT 40.345 156.565 40.685 157.535 ;
        RECT 41.060 156.735 41.390 157.535 ;
        RECT 41.560 156.905 41.890 157.705 ;
        RECT 42.190 156.735 42.520 157.535 ;
        RECT 43.165 156.905 43.415 157.705 ;
        RECT 41.060 156.565 43.495 156.735 ;
        RECT 43.685 156.565 43.855 157.705 ;
        RECT 44.025 156.565 44.365 157.535 ;
        RECT 37.175 156.145 37.525 156.395 ;
        RECT 33.450 155.325 33.780 155.805 ;
        RECT 33.950 155.155 34.175 155.615 ;
        RECT 34.345 155.325 34.675 155.805 ;
        RECT 34.865 155.155 35.115 155.955 ;
        RECT 35.285 155.325 35.625 155.955 ;
        RECT 37.710 155.935 37.880 156.565 ;
        RECT 38.050 156.145 38.380 156.345 ;
        RECT 38.550 156.145 38.880 156.345 ;
        RECT 39.050 156.145 39.470 156.345 ;
        RECT 39.645 156.315 39.815 156.565 ;
        RECT 39.645 156.145 40.340 156.315 ;
        RECT 40.510 156.005 40.685 156.565 ;
        RECT 40.855 156.145 41.205 156.395 ;
        RECT 35.795 155.155 36.085 155.880 ;
        RECT 37.380 155.325 37.880 155.935 ;
        RECT 38.510 155.805 39.735 155.975 ;
        RECT 40.455 155.955 40.685 156.005 ;
        RECT 38.510 155.325 38.840 155.805 ;
        RECT 39.010 155.155 39.235 155.615 ;
        RECT 39.405 155.325 39.735 155.805 ;
        RECT 39.925 155.155 40.175 155.955 ;
        RECT 40.345 155.325 40.685 155.955 ;
        RECT 41.390 155.935 41.560 156.565 ;
        RECT 41.730 156.145 42.060 156.345 ;
        RECT 42.230 156.145 42.560 156.345 ;
        RECT 42.730 156.145 43.150 156.345 ;
        RECT 43.325 156.315 43.495 156.565 ;
        RECT 43.325 156.145 44.020 156.315 ;
        RECT 41.060 155.325 41.560 155.935 ;
        RECT 42.190 155.805 43.415 155.975 ;
        RECT 44.190 155.955 44.365 156.565 ;
        RECT 44.535 156.615 46.205 157.705 ;
        RECT 46.380 157.270 51.725 157.705 ;
        RECT 44.535 156.095 45.285 156.615 ;
        RECT 42.190 155.325 42.520 155.805 ;
        RECT 42.690 155.155 42.915 155.615 ;
        RECT 43.085 155.325 43.415 155.805 ;
        RECT 43.605 155.155 43.855 155.955 ;
        RECT 44.025 155.325 44.365 155.955 ;
        RECT 45.455 155.925 46.205 156.445 ;
        RECT 47.970 156.020 48.320 157.270 ;
        RECT 52.270 156.725 52.525 157.395 ;
        RECT 52.705 156.905 52.990 157.705 ;
        RECT 53.170 156.985 53.500 157.495 ;
        RECT 44.535 155.155 46.205 155.925 ;
        RECT 49.800 155.700 50.140 156.530 ;
        RECT 52.270 155.865 52.450 156.725 ;
        RECT 53.170 156.395 53.420 156.985 ;
        RECT 53.770 156.835 53.940 157.445 ;
        RECT 54.110 157.015 54.440 157.705 ;
        RECT 54.670 157.155 54.910 157.445 ;
        RECT 55.110 157.325 55.530 157.705 ;
        RECT 55.710 157.235 56.340 157.485 ;
        RECT 56.810 157.325 57.140 157.705 ;
        RECT 55.710 157.155 55.880 157.235 ;
        RECT 57.310 157.155 57.480 157.445 ;
        RECT 57.660 157.325 58.040 157.705 ;
        RECT 58.280 157.320 59.110 157.490 ;
        RECT 54.670 156.985 55.880 157.155 ;
        RECT 52.620 156.065 53.420 156.395 ;
        RECT 46.380 155.155 51.725 155.700 ;
        RECT 52.270 155.665 52.525 155.865 ;
        RECT 52.185 155.495 52.525 155.665 ;
        RECT 52.270 155.335 52.525 155.495 ;
        RECT 52.705 155.155 52.990 155.615 ;
        RECT 53.170 155.415 53.420 156.065 ;
        RECT 53.620 156.815 53.940 156.835 ;
        RECT 53.620 156.645 55.540 156.815 ;
        RECT 53.620 155.750 53.810 156.645 ;
        RECT 55.710 156.475 55.880 156.985 ;
        RECT 56.050 156.725 56.570 157.035 ;
        RECT 53.980 156.305 55.880 156.475 ;
        RECT 53.980 156.245 54.310 156.305 ;
        RECT 54.460 156.075 54.790 156.135 ;
        RECT 54.130 155.805 54.790 156.075 ;
        RECT 53.620 155.420 53.940 155.750 ;
        RECT 54.120 155.155 54.780 155.635 ;
        RECT 54.980 155.545 55.150 156.305 ;
        RECT 56.050 156.135 56.230 156.545 ;
        RECT 55.320 155.965 55.650 156.085 ;
        RECT 56.400 155.965 56.570 156.725 ;
        RECT 55.320 155.795 56.570 155.965 ;
        RECT 56.740 156.905 58.110 157.155 ;
        RECT 56.740 156.135 56.930 156.905 ;
        RECT 57.860 156.645 58.110 156.905 ;
        RECT 57.100 156.475 57.350 156.635 ;
        RECT 58.280 156.475 58.450 157.320 ;
        RECT 59.345 157.035 59.515 157.535 ;
        RECT 59.685 157.205 60.015 157.705 ;
        RECT 58.620 156.645 59.120 157.025 ;
        RECT 59.345 156.865 60.040 157.035 ;
        RECT 57.100 156.305 58.450 156.475 ;
        RECT 58.030 156.265 58.450 156.305 ;
        RECT 56.740 155.795 57.160 156.135 ;
        RECT 57.450 155.805 57.860 156.135 ;
        RECT 54.980 155.375 55.830 155.545 ;
        RECT 56.390 155.155 56.710 155.615 ;
        RECT 56.910 155.365 57.160 155.795 ;
        RECT 57.450 155.155 57.860 155.595 ;
        RECT 58.030 155.535 58.200 156.265 ;
        RECT 58.370 155.715 58.720 156.085 ;
        RECT 58.900 155.775 59.120 156.645 ;
        RECT 59.290 156.075 59.700 156.695 ;
        RECT 59.870 155.895 60.040 156.865 ;
        RECT 59.345 155.705 60.040 155.895 ;
        RECT 58.030 155.335 59.045 155.535 ;
        RECT 59.345 155.375 59.515 155.705 ;
        RECT 59.685 155.155 60.015 155.535 ;
        RECT 60.230 155.415 60.455 157.535 ;
        RECT 60.625 157.205 60.955 157.705 ;
        RECT 61.125 157.035 61.295 157.535 ;
        RECT 60.630 156.865 61.295 157.035 ;
        RECT 60.630 155.875 60.860 156.865 ;
        RECT 61.030 156.045 61.380 156.695 ;
        RECT 61.555 156.540 61.845 157.705 ;
        RECT 62.015 156.855 62.275 157.535 ;
        RECT 62.445 156.925 62.695 157.705 ;
        RECT 62.945 157.155 63.195 157.535 ;
        RECT 63.365 157.325 63.720 157.705 ;
        RECT 64.725 157.315 65.060 157.535 ;
        RECT 64.325 157.155 64.555 157.195 ;
        RECT 62.945 156.955 64.555 157.155 ;
        RECT 62.945 156.945 63.780 156.955 ;
        RECT 64.370 156.865 64.555 156.955 ;
        RECT 60.630 155.705 61.295 155.875 ;
        RECT 60.625 155.155 60.955 155.535 ;
        RECT 61.125 155.415 61.295 155.705 ;
        RECT 61.555 155.155 61.845 155.880 ;
        RECT 62.015 155.655 62.185 156.855 ;
        RECT 63.885 156.755 64.215 156.785 ;
        RECT 62.415 156.695 64.215 156.755 ;
        RECT 64.805 156.695 65.060 157.315 ;
        RECT 62.355 156.585 65.060 156.695 ;
        RECT 62.355 156.550 62.555 156.585 ;
        RECT 62.355 155.975 62.525 156.550 ;
        RECT 63.885 156.525 65.060 156.585 ;
        RECT 65.900 156.735 66.230 157.535 ;
        RECT 66.400 156.905 66.730 157.705 ;
        RECT 67.030 156.735 67.360 157.535 ;
        RECT 68.005 156.905 68.255 157.705 ;
        RECT 65.900 156.565 68.335 156.735 ;
        RECT 68.525 156.565 68.695 157.705 ;
        RECT 68.865 156.565 69.205 157.535 ;
        RECT 62.755 156.110 63.165 156.415 ;
        RECT 63.335 156.145 63.665 156.355 ;
        RECT 62.355 155.855 62.625 155.975 ;
        RECT 62.355 155.810 63.200 155.855 ;
        RECT 62.445 155.685 63.200 155.810 ;
        RECT 63.455 155.745 63.665 156.145 ;
        RECT 63.910 156.145 64.385 156.355 ;
        RECT 64.575 156.145 65.065 156.345 ;
        RECT 65.695 156.145 66.045 156.395 ;
        RECT 63.910 155.745 64.130 156.145 ;
        RECT 66.230 155.935 66.400 156.565 ;
        RECT 66.570 156.145 66.900 156.345 ;
        RECT 67.070 156.145 67.400 156.345 ;
        RECT 67.570 156.145 67.990 156.345 ;
        RECT 68.165 156.315 68.335 156.565 ;
        RECT 68.165 156.145 68.860 156.315 ;
        RECT 69.030 156.005 69.205 156.565 ;
        RECT 62.015 155.325 62.275 155.655 ;
        RECT 63.030 155.535 63.200 155.685 ;
        RECT 62.445 155.155 62.775 155.515 ;
        RECT 63.030 155.325 64.330 155.535 ;
        RECT 64.605 155.155 65.060 155.920 ;
        RECT 65.900 155.325 66.400 155.935 ;
        RECT 67.030 155.805 68.255 155.975 ;
        RECT 68.975 155.955 69.205 156.005 ;
        RECT 67.030 155.325 67.360 155.805 ;
        RECT 67.530 155.155 67.755 155.615 ;
        RECT 67.925 155.325 68.255 155.805 ;
        RECT 68.445 155.155 68.695 155.955 ;
        RECT 68.865 155.325 69.205 155.955 ;
        RECT 69.375 156.565 69.715 157.535 ;
        RECT 69.885 156.565 70.055 157.705 ;
        RECT 70.325 156.905 70.575 157.705 ;
        RECT 71.220 156.735 71.550 157.535 ;
        RECT 71.850 156.905 72.180 157.705 ;
        RECT 72.350 156.735 72.680 157.535 ;
        RECT 70.245 156.565 72.680 156.735 ;
        RECT 73.055 156.615 74.265 157.705 ;
        RECT 74.435 156.615 77.945 157.705 ;
        RECT 78.120 157.270 83.465 157.705 ;
        RECT 69.375 155.955 69.550 156.565 ;
        RECT 70.245 156.315 70.415 156.565 ;
        RECT 69.720 156.145 70.415 156.315 ;
        RECT 70.590 156.145 71.010 156.345 ;
        RECT 71.180 156.145 71.510 156.345 ;
        RECT 71.680 156.145 72.010 156.345 ;
        RECT 69.375 155.325 69.715 155.955 ;
        RECT 69.885 155.155 70.135 155.955 ;
        RECT 70.325 155.805 71.550 155.975 ;
        RECT 70.325 155.325 70.655 155.805 ;
        RECT 70.825 155.155 71.050 155.615 ;
        RECT 71.220 155.325 71.550 155.805 ;
        RECT 72.180 155.935 72.350 156.565 ;
        RECT 72.535 156.145 72.885 156.395 ;
        RECT 73.055 156.075 73.575 156.615 ;
        RECT 72.180 155.325 72.680 155.935 ;
        RECT 73.745 155.905 74.265 156.445 ;
        RECT 74.435 156.095 76.125 156.615 ;
        RECT 76.295 155.925 77.945 156.445 ;
        RECT 79.710 156.020 80.060 157.270 ;
        RECT 83.840 156.735 84.170 157.535 ;
        RECT 84.340 156.905 84.670 157.705 ;
        RECT 84.970 156.735 85.300 157.535 ;
        RECT 85.945 156.905 86.195 157.705 ;
        RECT 83.840 156.565 86.275 156.735 ;
        RECT 86.465 156.565 86.635 157.705 ;
        RECT 86.805 156.565 87.145 157.535 ;
        RECT 73.055 155.155 74.265 155.905 ;
        RECT 74.435 155.155 77.945 155.925 ;
        RECT 81.540 155.700 81.880 156.530 ;
        RECT 83.635 156.145 83.985 156.395 ;
        RECT 84.170 155.935 84.340 156.565 ;
        RECT 84.510 156.145 84.840 156.345 ;
        RECT 85.010 156.145 85.340 156.345 ;
        RECT 85.510 156.145 85.930 156.345 ;
        RECT 86.105 156.315 86.275 156.565 ;
        RECT 86.105 156.145 86.800 156.315 ;
        RECT 78.120 155.155 83.465 155.700 ;
        RECT 83.840 155.325 84.340 155.935 ;
        RECT 84.970 155.805 86.195 155.975 ;
        RECT 86.970 155.955 87.145 156.565 ;
        RECT 87.315 156.540 87.605 157.705 ;
        RECT 88.235 156.615 89.905 157.705 ;
        RECT 90.280 156.735 90.610 157.535 ;
        RECT 90.780 156.905 91.110 157.705 ;
        RECT 91.410 156.735 91.740 157.535 ;
        RECT 92.385 156.905 92.635 157.705 ;
        RECT 88.235 156.095 88.985 156.615 ;
        RECT 90.280 156.565 92.715 156.735 ;
        RECT 92.905 156.565 93.075 157.705 ;
        RECT 93.245 156.565 93.585 157.535 ;
        RECT 84.970 155.325 85.300 155.805 ;
        RECT 85.470 155.155 85.695 155.615 ;
        RECT 85.865 155.325 86.195 155.805 ;
        RECT 86.385 155.155 86.635 155.955 ;
        RECT 86.805 155.325 87.145 155.955 ;
        RECT 89.155 155.925 89.905 156.445 ;
        RECT 90.075 156.145 90.425 156.395 ;
        RECT 90.610 155.935 90.780 156.565 ;
        RECT 90.950 156.145 91.280 156.345 ;
        RECT 91.450 156.145 91.780 156.345 ;
        RECT 91.950 156.145 92.370 156.345 ;
        RECT 92.545 156.315 92.715 156.565 ;
        RECT 92.545 156.145 93.240 156.315 ;
        RECT 87.315 155.155 87.605 155.880 ;
        RECT 88.235 155.155 89.905 155.925 ;
        RECT 90.280 155.325 90.780 155.935 ;
        RECT 91.410 155.805 92.635 155.975 ;
        RECT 93.410 155.955 93.585 156.565 ;
        RECT 91.410 155.325 91.740 155.805 ;
        RECT 91.910 155.155 92.135 155.615 ;
        RECT 92.305 155.325 92.635 155.805 ;
        RECT 92.825 155.155 93.075 155.955 ;
        RECT 93.245 155.325 93.585 155.955 ;
        RECT 93.755 156.565 94.095 157.535 ;
        RECT 94.265 156.565 94.435 157.705 ;
        RECT 94.705 156.905 94.955 157.705 ;
        RECT 95.600 156.735 95.930 157.535 ;
        RECT 96.230 156.905 96.560 157.705 ;
        RECT 96.730 156.735 97.060 157.535 ;
        RECT 94.625 156.565 97.060 156.735 ;
        RECT 97.435 156.615 99.105 157.705 ;
        RECT 99.390 157.075 99.675 157.535 ;
        RECT 99.845 157.245 100.115 157.705 ;
        RECT 99.390 156.855 100.345 157.075 ;
        RECT 93.755 156.005 93.930 156.565 ;
        RECT 94.625 156.315 94.795 156.565 ;
        RECT 94.100 156.145 94.795 156.315 ;
        RECT 94.970 156.145 95.390 156.345 ;
        RECT 95.560 156.145 95.890 156.345 ;
        RECT 96.060 156.145 96.390 156.345 ;
        RECT 93.755 155.955 93.985 156.005 ;
        RECT 93.755 155.325 94.095 155.955 ;
        RECT 94.265 155.155 94.515 155.955 ;
        RECT 94.705 155.805 95.930 155.975 ;
        RECT 94.705 155.325 95.035 155.805 ;
        RECT 95.205 155.155 95.430 155.615 ;
        RECT 95.600 155.325 95.930 155.805 ;
        RECT 96.560 155.935 96.730 156.565 ;
        RECT 96.915 156.145 97.265 156.395 ;
        RECT 97.435 156.095 98.185 156.615 ;
        RECT 96.560 155.325 97.060 155.935 ;
        RECT 98.355 155.925 99.105 156.445 ;
        RECT 99.275 156.125 99.965 156.685 ;
        RECT 100.135 155.955 100.345 156.855 ;
        RECT 97.435 155.155 99.105 155.925 ;
        RECT 99.390 155.785 100.345 155.955 ;
        RECT 100.515 156.685 100.915 157.535 ;
        RECT 101.105 157.075 101.385 157.535 ;
        RECT 101.905 157.245 102.230 157.705 ;
        RECT 101.105 156.855 102.230 157.075 ;
        RECT 100.515 156.125 101.610 156.685 ;
        RECT 101.780 156.395 102.230 156.855 ;
        RECT 102.400 156.565 102.785 157.535 ;
        RECT 99.390 155.325 99.675 155.785 ;
        RECT 99.845 155.155 100.115 155.615 ;
        RECT 100.515 155.325 100.915 156.125 ;
        RECT 101.780 156.065 102.335 156.395 ;
        RECT 101.780 155.955 102.230 156.065 ;
        RECT 101.105 155.785 102.230 155.955 ;
        RECT 102.505 155.895 102.785 156.565 ;
        RECT 101.105 155.325 101.385 155.785 ;
        RECT 101.905 155.155 102.230 155.615 ;
        RECT 102.400 155.325 102.785 155.895 ;
        RECT 102.960 156.515 103.215 157.395 ;
        RECT 103.385 156.565 103.690 157.705 ;
        RECT 104.030 157.325 104.360 157.705 ;
        RECT 104.540 157.155 104.710 157.445 ;
        RECT 104.880 157.245 105.130 157.705 ;
        RECT 103.910 156.985 104.710 157.155 ;
        RECT 105.300 157.195 106.170 157.535 ;
        RECT 102.960 155.865 103.170 156.515 ;
        RECT 103.910 156.395 104.080 156.985 ;
        RECT 105.300 156.815 105.470 157.195 ;
        RECT 106.405 157.075 106.575 157.535 ;
        RECT 106.745 157.245 107.115 157.705 ;
        RECT 107.410 157.105 107.580 157.445 ;
        RECT 107.750 157.275 108.080 157.705 ;
        RECT 108.315 157.105 108.485 157.445 ;
        RECT 104.250 156.645 105.470 156.815 ;
        RECT 105.640 156.735 106.100 157.025 ;
        RECT 106.405 156.905 106.965 157.075 ;
        RECT 107.410 156.935 108.485 157.105 ;
        RECT 108.655 157.205 109.335 157.535 ;
        RECT 109.550 157.205 109.800 157.535 ;
        RECT 109.970 157.245 110.220 157.705 ;
        RECT 106.795 156.765 106.965 156.905 ;
        RECT 105.640 156.725 106.605 156.735 ;
        RECT 105.300 156.555 105.470 156.645 ;
        RECT 105.930 156.565 106.605 156.725 ;
        RECT 103.340 156.365 104.080 156.395 ;
        RECT 103.340 156.065 104.255 156.365 ;
        RECT 103.930 155.890 104.255 156.065 ;
        RECT 102.960 155.335 103.215 155.865 ;
        RECT 103.385 155.155 103.690 155.615 ;
        RECT 103.935 155.535 104.255 155.890 ;
        RECT 104.425 156.105 104.965 156.475 ;
        RECT 105.300 156.385 105.705 156.555 ;
        RECT 104.425 155.705 104.665 156.105 ;
        RECT 105.145 155.935 105.365 156.215 ;
        RECT 104.835 155.765 105.365 155.935 ;
        RECT 104.835 155.535 105.005 155.765 ;
        RECT 105.535 155.605 105.705 156.385 ;
        RECT 105.875 155.775 106.225 156.395 ;
        RECT 106.395 155.775 106.605 156.565 ;
        RECT 106.795 156.595 108.295 156.765 ;
        RECT 106.795 155.905 106.965 156.595 ;
        RECT 108.655 156.425 108.825 157.205 ;
        RECT 109.630 157.075 109.800 157.205 ;
        RECT 107.135 156.255 108.825 156.425 ;
        RECT 108.995 156.645 109.460 157.035 ;
        RECT 109.630 156.905 110.025 157.075 ;
        RECT 107.135 156.075 107.305 156.255 ;
        RECT 103.935 155.365 105.005 155.535 ;
        RECT 105.175 155.155 105.365 155.595 ;
        RECT 105.535 155.325 106.485 155.605 ;
        RECT 106.795 155.515 107.055 155.905 ;
        RECT 107.475 155.835 108.265 156.085 ;
        RECT 106.705 155.345 107.055 155.515 ;
        RECT 107.265 155.155 107.595 155.615 ;
        RECT 108.470 155.545 108.640 156.255 ;
        RECT 108.995 156.055 109.165 156.645 ;
        RECT 108.810 155.835 109.165 156.055 ;
        RECT 109.335 155.835 109.685 156.455 ;
        RECT 109.855 155.545 110.025 156.905 ;
        RECT 110.390 156.735 110.715 157.520 ;
        RECT 110.195 155.685 110.655 156.735 ;
        RECT 108.470 155.375 109.325 155.545 ;
        RECT 109.530 155.375 110.025 155.545 ;
        RECT 110.195 155.155 110.525 155.515 ;
        RECT 110.885 155.415 111.055 157.535 ;
        RECT 111.225 157.205 111.555 157.705 ;
        RECT 111.725 157.035 111.980 157.535 ;
        RECT 111.230 156.865 111.980 157.035 ;
        RECT 111.230 155.875 111.460 156.865 ;
        RECT 111.630 156.045 111.980 156.695 ;
        RECT 112.155 156.615 113.365 157.705 ;
        RECT 112.155 156.075 112.675 156.615 ;
        RECT 112.845 155.905 113.365 156.445 ;
        RECT 111.230 155.705 111.980 155.875 ;
        RECT 111.225 155.155 111.555 155.535 ;
        RECT 111.725 155.415 111.980 155.705 ;
        RECT 112.155 155.155 113.365 155.905 ;
        RECT 15.010 154.985 113.450 155.155 ;
        RECT 15.095 154.235 16.305 154.985 ;
        RECT 15.095 153.695 15.615 154.235 ;
        RECT 16.935 154.215 18.605 154.985 ;
        RECT 15.785 153.525 16.305 154.065 ;
        RECT 15.095 152.435 16.305 153.525 ;
        RECT 16.935 153.525 17.685 154.045 ;
        RECT 17.855 153.695 18.605 154.215 ;
        RECT 18.780 154.245 19.035 154.815 ;
        RECT 19.205 154.585 19.535 154.985 ;
        RECT 19.960 154.450 20.490 154.815 ;
        RECT 19.960 154.415 20.135 154.450 ;
        RECT 19.205 154.245 20.135 154.415 ;
        RECT 20.680 154.305 20.955 154.815 ;
        RECT 18.780 153.575 18.950 154.245 ;
        RECT 19.205 154.075 19.375 154.245 ;
        RECT 19.120 153.745 19.375 154.075 ;
        RECT 19.600 153.745 19.795 154.075 ;
        RECT 16.935 152.435 18.605 153.525 ;
        RECT 18.780 152.605 19.115 153.575 ;
        RECT 19.285 152.435 19.455 153.575 ;
        RECT 19.625 152.775 19.795 153.745 ;
        RECT 19.965 153.115 20.135 154.245 ;
        RECT 20.305 153.455 20.475 154.255 ;
        RECT 20.675 154.135 20.955 154.305 ;
        RECT 20.680 153.655 20.955 154.135 ;
        RECT 21.125 153.455 21.315 154.815 ;
        RECT 21.495 154.450 22.005 154.985 ;
        RECT 22.225 154.175 22.470 154.780 ;
        RECT 22.915 154.260 23.205 154.985 ;
        RECT 23.840 154.245 24.095 154.815 ;
        RECT 24.265 154.585 24.595 154.985 ;
        RECT 25.020 154.450 25.550 154.815 ;
        RECT 25.020 154.415 25.195 154.450 ;
        RECT 24.265 154.245 25.195 154.415 ;
        RECT 21.515 154.005 22.745 154.175 ;
        RECT 20.305 153.285 21.315 153.455 ;
        RECT 21.485 153.440 22.235 153.630 ;
        RECT 19.965 152.945 21.090 153.115 ;
        RECT 21.485 152.775 21.655 153.440 ;
        RECT 22.405 153.195 22.745 154.005 ;
        RECT 19.625 152.605 21.655 152.775 ;
        RECT 21.825 152.435 21.995 153.195 ;
        RECT 22.230 152.785 22.745 153.195 ;
        RECT 22.915 152.435 23.205 153.600 ;
        RECT 23.840 153.575 24.010 154.245 ;
        RECT 24.265 154.075 24.435 154.245 ;
        RECT 24.180 153.745 24.435 154.075 ;
        RECT 24.660 153.745 24.855 154.075 ;
        RECT 23.840 152.605 24.175 153.575 ;
        RECT 24.345 152.435 24.515 153.575 ;
        RECT 24.685 152.775 24.855 153.745 ;
        RECT 25.025 153.115 25.195 154.245 ;
        RECT 25.365 153.455 25.535 154.255 ;
        RECT 25.740 153.965 26.015 154.815 ;
        RECT 25.735 153.795 26.015 153.965 ;
        RECT 25.740 153.655 26.015 153.795 ;
        RECT 26.185 153.455 26.375 154.815 ;
        RECT 26.555 154.450 27.065 154.985 ;
        RECT 27.285 154.175 27.530 154.780 ;
        RECT 28.435 154.215 31.025 154.985 ;
        RECT 26.575 154.005 27.805 154.175 ;
        RECT 25.365 153.285 26.375 153.455 ;
        RECT 26.545 153.440 27.295 153.630 ;
        RECT 25.025 152.945 26.150 153.115 ;
        RECT 26.545 152.775 26.715 153.440 ;
        RECT 27.465 153.195 27.805 154.005 ;
        RECT 24.685 152.605 26.715 152.775 ;
        RECT 26.885 152.435 27.055 153.195 ;
        RECT 27.290 152.785 27.805 153.195 ;
        RECT 28.435 153.525 29.645 154.045 ;
        RECT 29.815 153.695 31.025 154.215 ;
        RECT 31.195 154.185 31.535 154.815 ;
        RECT 31.705 154.185 31.955 154.985 ;
        RECT 32.145 154.335 32.475 154.815 ;
        RECT 32.645 154.525 32.870 154.985 ;
        RECT 33.040 154.335 33.370 154.815 ;
        RECT 31.195 153.575 31.370 154.185 ;
        RECT 32.145 154.165 33.370 154.335 ;
        RECT 34.000 154.205 34.500 154.815 ;
        RECT 35.080 154.205 35.580 154.815 ;
        RECT 31.540 153.825 32.235 153.995 ;
        RECT 32.065 153.575 32.235 153.825 ;
        RECT 32.410 153.795 32.830 153.995 ;
        RECT 33.000 153.795 33.330 153.995 ;
        RECT 33.500 153.795 33.830 153.995 ;
        RECT 34.000 153.575 34.170 154.205 ;
        RECT 34.355 153.745 34.705 153.995 ;
        RECT 34.875 153.745 35.225 153.995 ;
        RECT 35.410 153.575 35.580 154.205 ;
        RECT 36.210 154.335 36.540 154.815 ;
        RECT 36.710 154.525 36.935 154.985 ;
        RECT 37.105 154.335 37.435 154.815 ;
        RECT 36.210 154.165 37.435 154.335 ;
        RECT 37.625 154.185 37.875 154.985 ;
        RECT 38.045 154.185 38.385 154.815 ;
        RECT 38.760 154.205 39.260 154.815 ;
        RECT 35.750 153.795 36.080 153.995 ;
        RECT 36.250 153.795 36.580 153.995 ;
        RECT 36.750 153.795 37.170 153.995 ;
        RECT 37.345 153.825 38.040 153.995 ;
        RECT 37.345 153.575 37.515 153.825 ;
        RECT 38.210 153.625 38.385 154.185 ;
        RECT 38.555 153.745 38.905 153.995 ;
        RECT 38.155 153.575 38.385 153.625 ;
        RECT 39.090 153.575 39.260 154.205 ;
        RECT 39.890 154.335 40.220 154.815 ;
        RECT 40.390 154.525 40.615 154.985 ;
        RECT 40.785 154.335 41.115 154.815 ;
        RECT 39.890 154.165 41.115 154.335 ;
        RECT 41.305 154.185 41.555 154.985 ;
        RECT 41.725 154.185 42.065 154.815 ;
        RECT 42.235 154.235 43.445 154.985 ;
        RECT 39.430 153.795 39.760 153.995 ;
        RECT 39.930 153.795 40.260 153.995 ;
        RECT 40.430 153.795 40.850 153.995 ;
        RECT 41.025 153.825 41.720 153.995 ;
        RECT 41.025 153.575 41.195 153.825 ;
        RECT 41.890 153.575 42.065 154.185 ;
        RECT 28.435 152.435 31.025 153.525 ;
        RECT 31.195 152.605 31.535 153.575 ;
        RECT 31.705 152.435 31.875 153.575 ;
        RECT 32.065 153.405 34.500 153.575 ;
        RECT 32.145 152.435 32.395 153.235 ;
        RECT 33.040 152.605 33.370 153.405 ;
        RECT 33.670 152.435 34.000 153.235 ;
        RECT 34.170 152.605 34.500 153.405 ;
        RECT 35.080 153.405 37.515 153.575 ;
        RECT 35.080 152.605 35.410 153.405 ;
        RECT 35.580 152.435 35.910 153.235 ;
        RECT 36.210 152.605 36.540 153.405 ;
        RECT 37.185 152.435 37.435 153.235 ;
        RECT 37.705 152.435 37.875 153.575 ;
        RECT 38.045 152.605 38.385 153.575 ;
        RECT 38.760 153.405 41.195 153.575 ;
        RECT 38.760 152.605 39.090 153.405 ;
        RECT 39.260 152.435 39.590 153.235 ;
        RECT 39.890 152.605 40.220 153.405 ;
        RECT 40.865 152.435 41.115 153.235 ;
        RECT 41.385 152.435 41.555 153.575 ;
        RECT 41.725 152.605 42.065 153.575 ;
        RECT 42.235 153.525 42.755 154.065 ;
        RECT 42.925 153.695 43.445 154.235 ;
        RECT 43.615 154.215 47.125 154.985 ;
        RECT 43.615 153.525 45.305 154.045 ;
        RECT 45.475 153.695 47.125 154.215 ;
        RECT 47.335 154.165 47.565 154.985 ;
        RECT 47.735 154.185 48.065 154.815 ;
        RECT 47.315 153.745 47.645 153.995 ;
        RECT 47.815 153.585 48.065 154.185 ;
        RECT 48.235 154.165 48.445 154.985 ;
        RECT 48.675 154.260 48.965 154.985 ;
        RECT 49.140 154.275 49.395 154.805 ;
        RECT 49.565 154.525 49.870 154.985 ;
        RECT 50.115 154.605 51.185 154.775 ;
        RECT 49.140 153.625 49.350 154.275 ;
        RECT 50.115 154.250 50.435 154.605 ;
        RECT 50.110 154.075 50.435 154.250 ;
        RECT 49.520 153.775 50.435 154.075 ;
        RECT 50.605 154.035 50.845 154.435 ;
        RECT 51.015 154.375 51.185 154.605 ;
        RECT 51.355 154.545 51.545 154.985 ;
        RECT 51.715 154.535 52.665 154.815 ;
        RECT 52.885 154.625 53.235 154.795 ;
        RECT 51.015 154.205 51.545 154.375 ;
        RECT 49.520 153.745 50.260 153.775 ;
        RECT 42.235 152.435 43.445 153.525 ;
        RECT 43.615 152.435 47.125 153.525 ;
        RECT 47.335 152.435 47.565 153.575 ;
        RECT 47.735 152.605 48.065 153.585 ;
        RECT 48.235 152.435 48.445 153.575 ;
        RECT 48.675 152.435 48.965 153.600 ;
        RECT 49.140 152.745 49.395 153.625 ;
        RECT 49.565 152.435 49.870 153.575 ;
        RECT 50.090 153.155 50.260 153.745 ;
        RECT 50.605 153.665 51.145 154.035 ;
        RECT 51.325 153.925 51.545 154.205 ;
        RECT 51.715 153.755 51.885 154.535 ;
        RECT 51.480 153.585 51.885 153.755 ;
        RECT 52.055 153.745 52.405 154.365 ;
        RECT 51.480 153.495 51.650 153.585 ;
        RECT 52.575 153.575 52.785 154.365 ;
        RECT 50.430 153.325 51.650 153.495 ;
        RECT 52.110 153.415 52.785 153.575 ;
        RECT 50.090 152.985 50.890 153.155 ;
        RECT 50.210 152.435 50.540 152.815 ;
        RECT 50.720 152.695 50.890 152.985 ;
        RECT 51.480 152.945 51.650 153.325 ;
        RECT 51.820 153.405 52.785 153.415 ;
        RECT 52.975 154.235 53.235 154.625 ;
        RECT 53.445 154.525 53.775 154.985 ;
        RECT 54.650 154.595 55.505 154.765 ;
        RECT 55.710 154.595 56.205 154.765 ;
        RECT 56.375 154.625 56.705 154.985 ;
        RECT 52.975 153.545 53.145 154.235 ;
        RECT 53.315 153.885 53.485 154.065 ;
        RECT 53.655 154.055 54.445 154.305 ;
        RECT 54.650 153.885 54.820 154.595 ;
        RECT 54.990 154.085 55.345 154.305 ;
        RECT 53.315 153.715 55.005 153.885 ;
        RECT 51.820 153.115 52.280 153.405 ;
        RECT 52.975 153.375 54.475 153.545 ;
        RECT 52.975 153.235 53.145 153.375 ;
        RECT 52.585 153.065 53.145 153.235 ;
        RECT 51.060 152.435 51.310 152.895 ;
        RECT 51.480 152.605 52.350 152.945 ;
        RECT 52.585 152.605 52.755 153.065 ;
        RECT 53.590 153.035 54.665 153.205 ;
        RECT 52.925 152.435 53.295 152.895 ;
        RECT 53.590 152.695 53.760 153.035 ;
        RECT 53.930 152.435 54.260 152.865 ;
        RECT 54.495 152.695 54.665 153.035 ;
        RECT 54.835 152.935 55.005 153.715 ;
        RECT 55.175 153.495 55.345 154.085 ;
        RECT 55.515 153.685 55.865 154.305 ;
        RECT 55.175 153.105 55.640 153.495 ;
        RECT 56.035 153.235 56.205 154.595 ;
        RECT 56.375 153.405 56.835 154.455 ;
        RECT 55.810 153.065 56.205 153.235 ;
        RECT 55.810 152.935 55.980 153.065 ;
        RECT 54.835 152.605 55.515 152.935 ;
        RECT 55.730 152.605 55.980 152.935 ;
        RECT 56.150 152.435 56.400 152.895 ;
        RECT 56.570 152.620 56.895 153.405 ;
        RECT 57.065 152.605 57.235 154.725 ;
        RECT 57.405 154.605 57.735 154.985 ;
        RECT 57.905 154.435 58.160 154.725 ;
        RECT 57.410 154.265 58.160 154.435 ;
        RECT 58.450 154.355 58.735 154.815 ;
        RECT 58.905 154.525 59.175 154.985 ;
        RECT 57.410 153.275 57.640 154.265 ;
        RECT 58.450 154.185 59.405 154.355 ;
        RECT 57.810 153.445 58.160 154.095 ;
        RECT 58.335 153.455 59.025 154.015 ;
        RECT 59.195 153.285 59.405 154.185 ;
        RECT 57.410 153.105 58.160 153.275 ;
        RECT 57.405 152.435 57.735 152.935 ;
        RECT 57.905 152.605 58.160 153.105 ;
        RECT 58.450 153.065 59.405 153.285 ;
        RECT 59.575 154.015 59.975 154.815 ;
        RECT 60.165 154.355 60.445 154.815 ;
        RECT 60.965 154.525 61.290 154.985 ;
        RECT 60.165 154.185 61.290 154.355 ;
        RECT 61.460 154.245 61.845 154.815 ;
        RECT 60.840 154.075 61.290 154.185 ;
        RECT 59.575 153.455 60.670 154.015 ;
        RECT 60.840 153.745 61.395 154.075 ;
        RECT 58.450 152.605 58.735 153.065 ;
        RECT 58.905 152.435 59.175 152.895 ;
        RECT 59.575 152.605 59.975 153.455 ;
        RECT 60.840 153.285 61.290 153.745 ;
        RECT 61.565 153.575 61.845 154.245 ;
        RECT 60.165 153.065 61.290 153.285 ;
        RECT 60.165 152.605 60.445 153.065 ;
        RECT 60.965 152.435 61.290 152.895 ;
        RECT 61.460 152.605 61.845 153.575 ;
        RECT 62.015 154.185 62.355 154.815 ;
        RECT 62.525 154.185 62.775 154.985 ;
        RECT 62.965 154.335 63.295 154.815 ;
        RECT 63.465 154.525 63.690 154.985 ;
        RECT 63.860 154.335 64.190 154.815 ;
        RECT 62.015 153.575 62.190 154.185 ;
        RECT 62.965 154.165 64.190 154.335 ;
        RECT 64.820 154.205 65.320 154.815 ;
        RECT 65.755 154.505 66.035 154.985 ;
        RECT 66.205 154.335 66.465 154.725 ;
        RECT 66.640 154.505 66.895 154.985 ;
        RECT 67.065 154.335 67.360 154.725 ;
        RECT 67.540 154.505 67.815 154.985 ;
        RECT 67.985 154.485 68.285 154.815 ;
        RECT 62.360 153.825 63.055 153.995 ;
        RECT 62.885 153.575 63.055 153.825 ;
        RECT 63.230 153.795 63.650 153.995 ;
        RECT 63.820 153.795 64.150 153.995 ;
        RECT 64.320 153.795 64.650 153.995 ;
        RECT 64.820 153.575 64.990 154.205 ;
        RECT 65.710 154.165 67.360 154.335 ;
        RECT 65.175 153.745 65.525 153.995 ;
        RECT 65.710 153.655 66.115 154.165 ;
        RECT 66.285 153.825 67.425 153.995 ;
        RECT 62.015 152.605 62.355 153.575 ;
        RECT 62.525 152.435 62.695 153.575 ;
        RECT 62.885 153.405 65.320 153.575 ;
        RECT 65.710 153.485 66.465 153.655 ;
        RECT 62.965 152.435 63.215 153.235 ;
        RECT 63.860 152.605 64.190 153.405 ;
        RECT 64.490 152.435 64.820 153.235 ;
        RECT 64.990 152.605 65.320 153.405 ;
        RECT 65.750 152.435 66.035 153.305 ;
        RECT 66.205 153.235 66.465 153.485 ;
        RECT 67.255 153.575 67.425 153.825 ;
        RECT 67.595 153.745 67.945 154.315 ;
        RECT 68.115 153.575 68.285 154.485 ;
        RECT 67.255 153.405 68.285 153.575 ;
        RECT 66.205 153.065 67.325 153.235 ;
        RECT 66.205 152.605 66.465 153.065 ;
        RECT 66.640 152.435 66.895 152.895 ;
        RECT 67.065 152.605 67.325 153.065 ;
        RECT 67.495 152.435 67.805 153.235 ;
        RECT 67.975 152.605 68.285 153.405 ;
        RECT 68.455 154.225 69.165 154.815 ;
        RECT 69.675 154.455 70.005 154.815 ;
        RECT 70.205 154.625 70.535 154.985 ;
        RECT 70.705 154.455 71.035 154.815 ;
        RECT 69.675 154.245 71.035 154.455 ;
        RECT 71.305 154.435 71.475 154.815 ;
        RECT 71.690 154.605 72.020 154.985 ;
        RECT 71.305 154.265 72.020 154.435 ;
        RECT 68.455 154.135 68.685 154.225 ;
        RECT 68.455 153.255 68.660 154.135 ;
        RECT 68.830 153.455 69.160 153.995 ;
        RECT 69.335 153.745 69.830 154.075 ;
        RECT 70.150 153.745 70.525 154.075 ;
        RECT 70.735 153.745 71.045 154.075 ;
        RECT 69.335 153.455 69.660 153.745 ;
        RECT 69.855 153.255 70.185 153.475 ;
        RECT 68.455 153.025 70.185 153.255 ;
        RECT 68.455 152.605 69.155 153.025 ;
        RECT 69.355 152.435 69.685 152.795 ;
        RECT 69.855 152.625 70.185 153.025 ;
        RECT 70.355 152.775 70.525 153.745 ;
        RECT 71.215 153.715 71.570 154.085 ;
        RECT 71.850 154.075 72.020 154.265 ;
        RECT 72.190 154.240 72.445 154.815 ;
        RECT 71.850 153.745 72.105 154.075 ;
        RECT 71.850 153.535 72.020 153.745 ;
        RECT 70.705 152.435 71.035 153.495 ;
        RECT 71.305 153.365 72.020 153.535 ;
        RECT 72.275 153.510 72.445 154.240 ;
        RECT 72.620 154.145 72.880 154.985 ;
        RECT 73.055 154.235 74.265 154.985 ;
        RECT 74.435 154.260 74.725 154.985 ;
        RECT 71.305 152.605 71.475 153.365 ;
        RECT 71.690 152.435 72.020 153.195 ;
        RECT 72.190 152.605 72.445 153.510 ;
        RECT 72.620 152.435 72.880 153.585 ;
        RECT 73.055 153.525 73.575 154.065 ;
        RECT 73.745 153.695 74.265 154.235 ;
        RECT 75.355 154.215 77.025 154.985 ;
        RECT 73.055 152.435 74.265 153.525 ;
        RECT 74.435 152.435 74.725 153.600 ;
        RECT 75.355 153.525 76.105 154.045 ;
        RECT 76.275 153.695 77.025 154.215 ;
        RECT 77.255 154.165 77.465 154.985 ;
        RECT 77.635 154.185 77.965 154.815 ;
        RECT 77.635 153.585 77.885 154.185 ;
        RECT 78.135 154.165 78.365 154.985 ;
        RECT 78.635 154.165 78.845 154.985 ;
        RECT 79.015 154.185 79.345 154.815 ;
        RECT 78.055 153.745 78.385 153.995 ;
        RECT 79.015 153.585 79.265 154.185 ;
        RECT 79.515 154.165 79.745 154.985 ;
        RECT 80.965 154.435 81.135 154.815 ;
        RECT 81.315 154.605 81.645 154.985 ;
        RECT 80.965 154.265 81.630 154.435 ;
        RECT 81.825 154.310 82.085 154.815 ;
        RECT 79.435 153.745 79.765 153.995 ;
        RECT 80.895 153.715 81.225 154.085 ;
        RECT 81.460 154.010 81.630 154.265 ;
        RECT 81.460 153.680 81.745 154.010 ;
        RECT 75.355 152.435 77.025 153.525 ;
        RECT 77.255 152.435 77.465 153.575 ;
        RECT 77.635 152.605 77.965 153.585 ;
        RECT 78.135 152.435 78.365 153.575 ;
        RECT 78.635 152.435 78.845 153.575 ;
        RECT 79.015 152.605 79.345 153.585 ;
        RECT 79.515 152.435 79.745 153.575 ;
        RECT 81.460 153.535 81.630 153.680 ;
        RECT 80.965 153.365 81.630 153.535 ;
        RECT 81.915 153.510 82.085 154.310 ;
        RECT 83.180 154.435 83.435 154.725 ;
        RECT 83.605 154.605 83.935 154.985 ;
        RECT 83.180 154.265 83.930 154.435 ;
        RECT 80.965 152.605 81.135 153.365 ;
        RECT 81.315 152.435 81.645 153.195 ;
        RECT 81.815 152.605 82.085 153.510 ;
        RECT 83.180 153.445 83.530 154.095 ;
        RECT 83.700 153.275 83.930 154.265 ;
        RECT 83.180 153.105 83.930 153.275 ;
        RECT 83.180 152.605 83.435 153.105 ;
        RECT 83.605 152.435 83.935 152.935 ;
        RECT 84.105 152.605 84.275 154.725 ;
        RECT 84.635 154.625 84.965 154.985 ;
        RECT 85.135 154.595 85.630 154.765 ;
        RECT 85.835 154.595 86.690 154.765 ;
        RECT 84.505 153.405 84.965 154.455 ;
        RECT 84.445 152.620 84.770 153.405 ;
        RECT 85.135 153.235 85.305 154.595 ;
        RECT 85.475 153.685 85.825 154.305 ;
        RECT 85.995 154.085 86.350 154.305 ;
        RECT 85.995 153.495 86.165 154.085 ;
        RECT 86.520 153.885 86.690 154.595 ;
        RECT 87.565 154.525 87.895 154.985 ;
        RECT 88.105 154.625 88.455 154.795 ;
        RECT 86.895 154.055 87.685 154.305 ;
        RECT 88.105 154.235 88.365 154.625 ;
        RECT 88.675 154.535 89.625 154.815 ;
        RECT 89.795 154.545 89.985 154.985 ;
        RECT 90.155 154.605 91.225 154.775 ;
        RECT 87.855 153.885 88.025 154.065 ;
        RECT 85.135 153.065 85.530 153.235 ;
        RECT 85.700 153.105 86.165 153.495 ;
        RECT 86.335 153.715 88.025 153.885 ;
        RECT 85.360 152.935 85.530 153.065 ;
        RECT 86.335 152.935 86.505 153.715 ;
        RECT 88.195 153.545 88.365 154.235 ;
        RECT 86.865 153.375 88.365 153.545 ;
        RECT 88.555 153.575 88.765 154.365 ;
        RECT 88.935 153.745 89.285 154.365 ;
        RECT 89.455 153.755 89.625 154.535 ;
        RECT 90.155 154.375 90.325 154.605 ;
        RECT 89.795 154.205 90.325 154.375 ;
        RECT 89.795 153.925 90.015 154.205 ;
        RECT 90.495 154.035 90.735 154.435 ;
        RECT 89.455 153.585 89.860 153.755 ;
        RECT 90.195 153.665 90.735 154.035 ;
        RECT 90.905 154.250 91.225 154.605 ;
        RECT 91.470 154.525 91.775 154.985 ;
        RECT 91.945 154.275 92.200 154.805 ;
        RECT 90.905 154.075 91.230 154.250 ;
        RECT 90.905 153.775 91.820 154.075 ;
        RECT 91.080 153.745 91.820 153.775 ;
        RECT 88.555 153.415 89.230 153.575 ;
        RECT 89.690 153.495 89.860 153.585 ;
        RECT 88.555 153.405 89.520 153.415 ;
        RECT 88.195 153.235 88.365 153.375 ;
        RECT 84.940 152.435 85.190 152.895 ;
        RECT 85.360 152.605 85.610 152.935 ;
        RECT 85.825 152.605 86.505 152.935 ;
        RECT 86.675 153.035 87.750 153.205 ;
        RECT 88.195 153.065 88.755 153.235 ;
        RECT 89.060 153.115 89.520 153.405 ;
        RECT 89.690 153.325 90.910 153.495 ;
        RECT 86.675 152.695 86.845 153.035 ;
        RECT 87.080 152.435 87.410 152.865 ;
        RECT 87.580 152.695 87.750 153.035 ;
        RECT 88.045 152.435 88.415 152.895 ;
        RECT 88.585 152.605 88.755 153.065 ;
        RECT 89.690 152.945 89.860 153.325 ;
        RECT 91.080 153.155 91.250 153.745 ;
        RECT 91.990 153.625 92.200 154.275 ;
        RECT 88.990 152.605 89.860 152.945 ;
        RECT 90.450 152.985 91.250 153.155 ;
        RECT 90.030 152.435 90.280 152.895 ;
        RECT 90.450 152.695 90.620 152.985 ;
        RECT 90.800 152.435 91.130 152.815 ;
        RECT 91.470 152.435 91.775 153.575 ;
        RECT 91.945 152.745 92.200 153.625 ;
        RECT 92.375 154.245 92.760 154.815 ;
        RECT 92.930 154.525 93.255 154.985 ;
        RECT 93.775 154.355 94.055 154.815 ;
        RECT 92.375 153.575 92.655 154.245 ;
        RECT 92.930 154.185 94.055 154.355 ;
        RECT 92.930 154.075 93.380 154.185 ;
        RECT 92.825 153.745 93.380 154.075 ;
        RECT 94.245 154.015 94.645 154.815 ;
        RECT 95.045 154.525 95.315 154.985 ;
        RECT 95.485 154.355 95.770 154.815 ;
        RECT 92.375 152.605 92.760 153.575 ;
        RECT 92.930 153.285 93.380 153.745 ;
        RECT 93.550 153.455 94.645 154.015 ;
        RECT 92.930 153.065 94.055 153.285 ;
        RECT 92.930 152.435 93.255 152.895 ;
        RECT 93.775 152.605 94.055 153.065 ;
        RECT 94.245 152.605 94.645 153.455 ;
        RECT 94.815 154.185 95.770 154.355 ;
        RECT 96.055 154.185 96.395 154.815 ;
        RECT 96.565 154.185 96.815 154.985 ;
        RECT 97.005 154.335 97.335 154.815 ;
        RECT 97.505 154.525 97.730 154.985 ;
        RECT 97.900 154.335 98.230 154.815 ;
        RECT 94.815 153.285 95.025 154.185 ;
        RECT 95.195 153.455 95.885 154.015 ;
        RECT 96.055 153.575 96.230 154.185 ;
        RECT 97.005 154.165 98.230 154.335 ;
        RECT 98.860 154.205 99.360 154.815 ;
        RECT 100.195 154.260 100.485 154.985 ;
        RECT 100.655 154.215 102.325 154.985 ;
        RECT 96.400 153.825 97.095 153.995 ;
        RECT 96.925 153.575 97.095 153.825 ;
        RECT 97.270 153.795 97.690 153.995 ;
        RECT 97.860 153.795 98.190 153.995 ;
        RECT 98.360 153.795 98.690 153.995 ;
        RECT 98.860 153.575 99.030 154.205 ;
        RECT 99.215 153.745 99.565 153.995 ;
        RECT 94.815 153.065 95.770 153.285 ;
        RECT 95.045 152.435 95.315 152.895 ;
        RECT 95.485 152.605 95.770 153.065 ;
        RECT 96.055 152.605 96.395 153.575 ;
        RECT 96.565 152.435 96.735 153.575 ;
        RECT 96.925 153.405 99.360 153.575 ;
        RECT 97.005 152.435 97.255 153.235 ;
        RECT 97.900 152.605 98.230 153.405 ;
        RECT 98.530 152.435 98.860 153.235 ;
        RECT 99.030 152.605 99.360 153.405 ;
        RECT 100.195 152.435 100.485 153.600 ;
        RECT 100.655 153.525 101.405 154.045 ;
        RECT 101.575 153.695 102.325 154.215 ;
        RECT 102.770 154.175 103.015 154.780 ;
        RECT 103.235 154.450 103.745 154.985 ;
        RECT 102.495 154.005 103.725 154.175 ;
        RECT 100.655 152.435 102.325 153.525 ;
        RECT 102.495 153.195 102.835 154.005 ;
        RECT 103.005 153.440 103.755 153.630 ;
        RECT 102.495 152.785 103.010 153.195 ;
        RECT 103.245 152.435 103.415 153.195 ;
        RECT 103.585 152.775 103.755 153.440 ;
        RECT 103.925 153.455 104.115 154.815 ;
        RECT 104.285 154.305 104.560 154.815 ;
        RECT 104.750 154.450 105.280 154.815 ;
        RECT 105.705 154.585 106.035 154.985 ;
        RECT 105.105 154.415 105.280 154.450 ;
        RECT 104.285 154.135 104.565 154.305 ;
        RECT 104.285 153.655 104.560 154.135 ;
        RECT 104.765 153.455 104.935 154.255 ;
        RECT 103.925 153.285 104.935 153.455 ;
        RECT 105.105 154.245 106.035 154.415 ;
        RECT 106.205 154.245 106.460 154.815 ;
        RECT 105.105 153.115 105.275 154.245 ;
        RECT 105.865 154.075 106.035 154.245 ;
        RECT 104.150 152.945 105.275 153.115 ;
        RECT 105.445 153.745 105.640 154.075 ;
        RECT 105.865 153.745 106.120 154.075 ;
        RECT 105.445 152.775 105.615 153.745 ;
        RECT 106.290 153.575 106.460 154.245 ;
        RECT 106.635 154.235 107.845 154.985 ;
        RECT 108.105 154.435 108.275 154.815 ;
        RECT 108.455 154.605 108.785 154.985 ;
        RECT 108.105 154.265 108.770 154.435 ;
        RECT 108.965 154.310 109.225 154.815 ;
        RECT 103.585 152.605 105.615 152.775 ;
        RECT 105.785 152.435 105.955 153.575 ;
        RECT 106.125 152.605 106.460 153.575 ;
        RECT 106.635 153.525 107.155 154.065 ;
        RECT 107.325 153.695 107.845 154.235 ;
        RECT 108.035 153.715 108.365 154.085 ;
        RECT 108.600 154.010 108.770 154.265 ;
        RECT 108.600 153.680 108.885 154.010 ;
        RECT 108.600 153.535 108.770 153.680 ;
        RECT 106.635 152.435 107.845 153.525 ;
        RECT 108.105 153.365 108.770 153.535 ;
        RECT 109.055 153.510 109.225 154.310 ;
        RECT 109.395 154.215 111.985 154.985 ;
        RECT 112.155 154.235 113.365 154.985 ;
        RECT 108.105 152.605 108.275 153.365 ;
        RECT 108.455 152.435 108.785 153.195 ;
        RECT 108.955 152.605 109.225 153.510 ;
        RECT 109.395 153.525 110.605 154.045 ;
        RECT 110.775 153.695 111.985 154.215 ;
        RECT 112.155 153.525 112.675 154.065 ;
        RECT 112.845 153.695 113.365 154.235 ;
        RECT 109.395 152.435 111.985 153.525 ;
        RECT 112.155 152.435 113.365 153.525 ;
        RECT 15.010 152.265 113.450 152.435 ;
        RECT 15.095 151.175 16.305 152.265 ;
        RECT 17.770 151.925 18.025 151.955 ;
        RECT 17.685 151.755 18.025 151.925 ;
        RECT 15.095 150.465 15.615 151.005 ;
        RECT 15.785 150.635 16.305 151.175 ;
        RECT 17.770 151.285 18.025 151.755 ;
        RECT 18.205 151.465 18.490 152.265 ;
        RECT 18.670 151.545 19.000 152.055 ;
        RECT 15.095 149.715 16.305 150.465 ;
        RECT 17.770 150.425 17.950 151.285 ;
        RECT 18.670 150.955 18.920 151.545 ;
        RECT 19.270 151.395 19.440 152.005 ;
        RECT 19.610 151.575 19.940 152.265 ;
        RECT 20.170 151.715 20.410 152.005 ;
        RECT 20.610 151.885 21.030 152.265 ;
        RECT 21.210 151.795 21.840 152.045 ;
        RECT 22.310 151.885 22.640 152.265 ;
        RECT 21.210 151.715 21.380 151.795 ;
        RECT 22.810 151.715 22.980 152.005 ;
        RECT 23.160 151.885 23.540 152.265 ;
        RECT 23.780 151.880 24.610 152.050 ;
        RECT 20.170 151.545 21.380 151.715 ;
        RECT 18.120 150.625 18.920 150.955 ;
        RECT 17.770 149.895 18.025 150.425 ;
        RECT 18.205 149.715 18.490 150.175 ;
        RECT 18.670 149.975 18.920 150.625 ;
        RECT 19.120 151.375 19.440 151.395 ;
        RECT 19.120 151.205 21.040 151.375 ;
        RECT 19.120 150.310 19.310 151.205 ;
        RECT 21.210 151.035 21.380 151.545 ;
        RECT 21.550 151.285 22.070 151.595 ;
        RECT 19.480 150.865 21.380 151.035 ;
        RECT 19.480 150.805 19.810 150.865 ;
        RECT 19.960 150.635 20.290 150.695 ;
        RECT 19.630 150.365 20.290 150.635 ;
        RECT 19.120 149.980 19.440 150.310 ;
        RECT 19.620 149.715 20.280 150.195 ;
        RECT 20.480 150.105 20.650 150.865 ;
        RECT 21.550 150.695 21.730 151.105 ;
        RECT 20.820 150.525 21.150 150.645 ;
        RECT 21.900 150.525 22.070 151.285 ;
        RECT 20.820 150.355 22.070 150.525 ;
        RECT 22.240 151.465 23.610 151.715 ;
        RECT 22.240 150.695 22.430 151.465 ;
        RECT 23.360 151.205 23.610 151.465 ;
        RECT 22.600 151.035 22.850 151.195 ;
        RECT 23.780 151.035 23.950 151.880 ;
        RECT 24.845 151.595 25.015 152.095 ;
        RECT 25.185 151.765 25.515 152.265 ;
        RECT 24.120 151.205 24.620 151.585 ;
        RECT 24.845 151.425 25.540 151.595 ;
        RECT 22.600 150.865 23.950 151.035 ;
        RECT 23.530 150.825 23.950 150.865 ;
        RECT 22.240 150.355 22.660 150.695 ;
        RECT 22.950 150.365 23.360 150.695 ;
        RECT 20.480 149.935 21.330 150.105 ;
        RECT 21.890 149.715 22.210 150.175 ;
        RECT 22.410 149.925 22.660 150.355 ;
        RECT 22.950 149.715 23.360 150.155 ;
        RECT 23.530 150.095 23.700 150.825 ;
        RECT 23.870 150.275 24.220 150.645 ;
        RECT 24.400 150.335 24.620 151.205 ;
        RECT 24.790 150.635 25.200 151.255 ;
        RECT 25.370 150.455 25.540 151.425 ;
        RECT 24.845 150.265 25.540 150.455 ;
        RECT 23.530 149.895 24.545 150.095 ;
        RECT 24.845 149.935 25.015 150.265 ;
        RECT 25.185 149.715 25.515 150.095 ;
        RECT 25.730 149.975 25.955 152.095 ;
        RECT 26.125 151.765 26.455 152.265 ;
        RECT 26.625 151.595 26.795 152.095 ;
        RECT 26.130 151.425 26.795 151.595 ;
        RECT 26.130 150.435 26.360 151.425 ;
        RECT 26.530 150.605 26.880 151.255 ;
        RECT 27.515 151.125 27.785 152.095 ;
        RECT 27.995 151.465 28.275 152.265 ;
        RECT 28.445 151.755 30.100 152.045 ;
        RECT 28.510 151.415 30.100 151.585 ;
        RECT 28.510 151.295 28.680 151.415 ;
        RECT 27.955 151.125 28.680 151.295 ;
        RECT 26.130 150.265 26.795 150.435 ;
        RECT 26.125 149.715 26.455 150.095 ;
        RECT 26.625 149.975 26.795 150.265 ;
        RECT 27.515 150.390 27.685 151.125 ;
        RECT 27.955 150.955 28.125 151.125 ;
        RECT 27.855 150.625 28.125 150.955 ;
        RECT 28.295 150.625 28.700 150.955 ;
        RECT 28.870 150.625 29.580 151.245 ;
        RECT 29.780 151.125 30.100 151.415 ;
        RECT 30.275 151.505 30.790 151.915 ;
        RECT 31.025 151.505 31.195 152.265 ;
        RECT 31.365 151.925 33.395 152.095 ;
        RECT 27.955 150.455 28.125 150.625 ;
        RECT 27.515 150.045 27.785 150.390 ;
        RECT 27.955 150.285 29.565 150.455 ;
        RECT 29.750 150.385 30.100 150.955 ;
        RECT 30.275 150.695 30.615 151.505 ;
        RECT 31.365 151.260 31.535 151.925 ;
        RECT 31.930 151.585 33.055 151.755 ;
        RECT 30.785 151.070 31.535 151.260 ;
        RECT 31.705 151.245 32.715 151.415 ;
        RECT 30.275 150.525 31.505 150.695 ;
        RECT 27.975 149.715 28.355 150.115 ;
        RECT 28.525 149.935 28.695 150.285 ;
        RECT 28.865 149.715 29.195 150.115 ;
        RECT 29.395 149.935 29.565 150.285 ;
        RECT 29.765 149.715 30.095 150.215 ;
        RECT 30.550 149.920 30.795 150.525 ;
        RECT 31.015 149.715 31.525 150.250 ;
        RECT 31.705 149.885 31.895 151.245 ;
        RECT 32.065 150.905 32.340 151.045 ;
        RECT 32.065 150.735 32.345 150.905 ;
        RECT 32.065 149.885 32.340 150.735 ;
        RECT 32.545 150.445 32.715 151.245 ;
        RECT 32.885 150.455 33.055 151.585 ;
        RECT 33.225 150.955 33.395 151.925 ;
        RECT 33.565 151.125 33.735 152.265 ;
        RECT 33.905 151.125 34.240 152.095 ;
        RECT 33.225 150.625 33.420 150.955 ;
        RECT 33.645 150.625 33.900 150.955 ;
        RECT 33.645 150.455 33.815 150.625 ;
        RECT 34.070 150.455 34.240 151.125 ;
        RECT 32.885 150.285 33.815 150.455 ;
        RECT 32.885 150.250 33.060 150.285 ;
        RECT 32.530 149.885 33.060 150.250 ;
        RECT 33.485 149.715 33.815 150.115 ;
        RECT 33.985 149.885 34.240 150.455 ;
        RECT 34.415 151.190 34.685 152.095 ;
        RECT 34.855 151.505 35.185 152.265 ;
        RECT 35.365 151.335 35.535 152.095 ;
        RECT 34.415 150.390 34.585 151.190 ;
        RECT 34.870 151.165 35.535 151.335 ;
        RECT 34.870 151.020 35.040 151.165 ;
        RECT 35.795 151.100 36.085 152.265 ;
        RECT 36.255 151.125 36.595 152.095 ;
        RECT 36.765 151.125 36.935 152.265 ;
        RECT 37.205 151.465 37.455 152.265 ;
        RECT 38.100 151.295 38.430 152.095 ;
        RECT 38.730 151.465 39.060 152.265 ;
        RECT 39.230 151.295 39.560 152.095 ;
        RECT 37.125 151.125 39.560 151.295 ;
        RECT 40.855 151.125 41.195 152.095 ;
        RECT 41.365 151.125 41.535 152.265 ;
        RECT 41.805 151.465 42.055 152.265 ;
        RECT 42.700 151.295 43.030 152.095 ;
        RECT 43.330 151.465 43.660 152.265 ;
        RECT 43.830 151.295 44.160 152.095 ;
        RECT 44.650 151.635 44.935 152.095 ;
        RECT 45.105 151.805 45.375 152.265 ;
        RECT 44.650 151.415 45.605 151.635 ;
        RECT 41.725 151.125 44.160 151.295 ;
        RECT 34.755 150.690 35.040 151.020 ;
        RECT 34.870 150.435 35.040 150.690 ;
        RECT 35.275 150.615 35.605 150.985 ;
        RECT 36.255 150.515 36.430 151.125 ;
        RECT 37.125 150.875 37.295 151.125 ;
        RECT 36.600 150.705 37.295 150.875 ;
        RECT 37.470 150.705 37.890 150.905 ;
        RECT 38.060 150.705 38.390 150.905 ;
        RECT 38.560 150.705 38.890 150.905 ;
        RECT 34.415 149.885 34.675 150.390 ;
        RECT 34.870 150.265 35.535 150.435 ;
        RECT 34.855 149.715 35.185 150.095 ;
        RECT 35.365 149.885 35.535 150.265 ;
        RECT 35.795 149.715 36.085 150.440 ;
        RECT 36.255 149.885 36.595 150.515 ;
        RECT 36.765 149.715 37.015 150.515 ;
        RECT 37.205 150.365 38.430 150.535 ;
        RECT 37.205 149.885 37.535 150.365 ;
        RECT 37.705 149.715 37.930 150.175 ;
        RECT 38.100 149.885 38.430 150.365 ;
        RECT 39.060 150.495 39.230 151.125 ;
        RECT 39.415 150.705 39.765 150.955 ;
        RECT 40.855 150.515 41.030 151.125 ;
        RECT 41.725 150.875 41.895 151.125 ;
        RECT 41.200 150.705 41.895 150.875 ;
        RECT 42.070 150.705 42.490 150.905 ;
        RECT 42.660 150.705 42.990 150.905 ;
        RECT 43.160 150.705 43.490 150.905 ;
        RECT 39.060 149.885 39.560 150.495 ;
        RECT 40.855 149.885 41.195 150.515 ;
        RECT 41.365 149.715 41.615 150.515 ;
        RECT 41.805 150.365 43.030 150.535 ;
        RECT 41.805 149.885 42.135 150.365 ;
        RECT 42.305 149.715 42.530 150.175 ;
        RECT 42.700 149.885 43.030 150.365 ;
        RECT 43.660 150.495 43.830 151.125 ;
        RECT 44.015 150.705 44.365 150.955 ;
        RECT 44.535 150.685 45.225 151.245 ;
        RECT 45.395 150.515 45.605 151.415 ;
        RECT 43.660 149.885 44.160 150.495 ;
        RECT 44.650 150.345 45.605 150.515 ;
        RECT 45.775 151.245 46.175 152.095 ;
        RECT 46.365 151.635 46.645 152.095 ;
        RECT 47.165 151.805 47.490 152.265 ;
        RECT 46.365 151.415 47.490 151.635 ;
        RECT 45.775 150.685 46.870 151.245 ;
        RECT 47.040 150.955 47.490 151.415 ;
        RECT 47.660 151.125 48.045 152.095 ;
        RECT 44.650 149.885 44.935 150.345 ;
        RECT 45.105 149.715 45.375 150.175 ;
        RECT 45.775 149.885 46.175 150.685 ;
        RECT 47.040 150.625 47.595 150.955 ;
        RECT 47.040 150.515 47.490 150.625 ;
        RECT 46.365 150.345 47.490 150.515 ;
        RECT 47.765 150.455 48.045 151.125 ;
        RECT 48.215 151.505 48.730 151.915 ;
        RECT 48.965 151.505 49.135 152.265 ;
        RECT 49.305 151.925 51.335 152.095 ;
        RECT 48.215 150.695 48.555 151.505 ;
        RECT 49.305 151.260 49.475 151.925 ;
        RECT 49.870 151.585 50.995 151.755 ;
        RECT 48.725 151.070 49.475 151.260 ;
        RECT 49.645 151.245 50.655 151.415 ;
        RECT 48.215 150.525 49.445 150.695 ;
        RECT 46.365 149.885 46.645 150.345 ;
        RECT 47.165 149.715 47.490 150.175 ;
        RECT 47.660 149.885 48.045 150.455 ;
        RECT 48.490 149.920 48.735 150.525 ;
        RECT 48.955 149.715 49.465 150.250 ;
        RECT 49.645 149.885 49.835 151.245 ;
        RECT 50.005 150.905 50.280 151.045 ;
        RECT 50.005 150.735 50.285 150.905 ;
        RECT 50.005 149.885 50.280 150.735 ;
        RECT 50.485 150.445 50.655 151.245 ;
        RECT 50.825 150.455 50.995 151.585 ;
        RECT 51.165 150.955 51.335 151.925 ;
        RECT 51.505 151.125 51.675 152.265 ;
        RECT 51.845 151.125 52.180 152.095 ;
        RECT 52.445 151.520 52.715 152.265 ;
        RECT 53.345 152.260 59.620 152.265 ;
        RECT 52.885 151.350 53.175 152.090 ;
        RECT 53.345 151.535 53.600 152.260 ;
        RECT 53.785 151.365 54.045 152.090 ;
        RECT 54.215 151.535 54.460 152.260 ;
        RECT 54.645 151.365 54.905 152.090 ;
        RECT 55.075 151.535 55.320 152.260 ;
        RECT 55.505 151.365 55.765 152.090 ;
        RECT 55.935 151.535 56.180 152.260 ;
        RECT 56.350 151.365 56.610 152.090 ;
        RECT 56.780 151.535 57.040 152.260 ;
        RECT 57.210 151.365 57.470 152.090 ;
        RECT 57.640 151.535 57.900 152.260 ;
        RECT 58.070 151.365 58.330 152.090 ;
        RECT 58.500 151.535 58.760 152.260 ;
        RECT 58.930 151.365 59.190 152.090 ;
        RECT 59.360 151.465 59.620 152.260 ;
        RECT 53.785 151.350 59.190 151.365 ;
        RECT 51.165 150.625 51.360 150.955 ;
        RECT 51.585 150.625 51.840 150.955 ;
        RECT 51.585 150.455 51.755 150.625 ;
        RECT 52.010 150.455 52.180 151.125 ;
        RECT 52.445 151.125 59.190 151.350 ;
        RECT 52.445 150.565 53.610 151.125 ;
        RECT 59.790 150.955 60.040 152.090 ;
        RECT 60.220 151.455 60.480 152.265 ;
        RECT 60.655 150.955 60.900 152.095 ;
        RECT 61.080 151.455 61.375 152.265 ;
        RECT 61.555 151.100 61.845 152.265 ;
        RECT 62.015 151.125 62.355 152.095 ;
        RECT 62.525 151.125 62.695 152.265 ;
        RECT 62.965 151.465 63.215 152.265 ;
        RECT 63.860 151.295 64.190 152.095 ;
        RECT 64.490 151.465 64.820 152.265 ;
        RECT 64.990 151.295 65.320 152.095 ;
        RECT 66.210 151.395 66.495 152.265 ;
        RECT 66.665 151.635 66.925 152.095 ;
        RECT 67.100 151.805 67.355 152.265 ;
        RECT 67.525 151.635 67.785 152.095 ;
        RECT 66.665 151.465 67.785 151.635 ;
        RECT 67.955 151.465 68.265 152.265 ;
        RECT 62.885 151.125 65.320 151.295 ;
        RECT 66.665 151.215 66.925 151.465 ;
        RECT 68.435 151.295 68.745 152.095 ;
        RECT 53.780 150.705 60.900 150.955 ;
        RECT 50.825 150.285 51.755 150.455 ;
        RECT 50.825 150.250 51.000 150.285 ;
        RECT 50.470 149.885 51.000 150.250 ;
        RECT 51.425 149.715 51.755 150.115 ;
        RECT 51.925 149.885 52.180 150.455 ;
        RECT 52.415 150.535 53.610 150.565 ;
        RECT 52.415 150.395 59.190 150.535 ;
        RECT 52.445 150.365 59.190 150.395 ;
        RECT 52.445 149.715 52.745 150.195 ;
        RECT 52.915 149.910 53.175 150.365 ;
        RECT 53.345 149.715 53.605 150.195 ;
        RECT 53.785 149.910 54.045 150.365 ;
        RECT 54.215 149.715 54.465 150.195 ;
        RECT 54.645 149.910 54.905 150.365 ;
        RECT 55.075 149.715 55.325 150.195 ;
        RECT 55.505 149.910 55.765 150.365 ;
        RECT 55.935 149.715 56.180 150.195 ;
        RECT 56.350 149.910 56.625 150.365 ;
        RECT 56.795 149.715 57.040 150.195 ;
        RECT 57.210 149.910 57.470 150.365 ;
        RECT 57.640 149.715 57.900 150.195 ;
        RECT 58.070 149.910 58.330 150.365 ;
        RECT 58.500 149.715 58.760 150.195 ;
        RECT 58.930 149.910 59.190 150.365 ;
        RECT 59.360 149.715 59.620 150.275 ;
        RECT 59.790 149.895 60.040 150.705 ;
        RECT 60.220 149.715 60.480 150.240 ;
        RECT 60.650 149.895 60.900 150.705 ;
        RECT 61.070 150.395 61.385 150.955 ;
        RECT 62.015 150.515 62.190 151.125 ;
        RECT 62.885 150.875 63.055 151.125 ;
        RECT 62.360 150.705 63.055 150.875 ;
        RECT 63.230 150.705 63.650 150.905 ;
        RECT 63.820 150.705 64.150 150.905 ;
        RECT 64.320 150.705 64.650 150.905 ;
        RECT 61.080 149.715 61.385 150.225 ;
        RECT 61.555 149.715 61.845 150.440 ;
        RECT 62.015 149.885 62.355 150.515 ;
        RECT 62.525 149.715 62.775 150.515 ;
        RECT 62.965 150.365 64.190 150.535 ;
        RECT 62.965 149.885 63.295 150.365 ;
        RECT 63.465 149.715 63.690 150.175 ;
        RECT 63.860 149.885 64.190 150.365 ;
        RECT 64.820 150.495 64.990 151.125 ;
        RECT 66.170 151.045 66.925 151.215 ;
        RECT 67.715 151.125 68.745 151.295 ;
        RECT 65.175 150.705 65.525 150.955 ;
        RECT 66.170 150.535 66.575 151.045 ;
        RECT 67.715 150.875 67.885 151.125 ;
        RECT 66.745 150.705 67.885 150.875 ;
        RECT 64.820 149.885 65.320 150.495 ;
        RECT 66.170 150.365 67.820 150.535 ;
        RECT 68.055 150.385 68.405 150.955 ;
        RECT 66.215 149.715 66.495 150.195 ;
        RECT 66.665 149.975 66.925 150.365 ;
        RECT 67.100 149.715 67.355 150.195 ;
        RECT 67.525 149.975 67.820 150.365 ;
        RECT 68.575 150.215 68.745 151.125 ;
        RECT 68.000 149.715 68.275 150.195 ;
        RECT 68.445 149.885 68.745 150.215 ;
        RECT 68.915 151.125 69.185 152.095 ;
        RECT 69.395 151.465 69.675 152.265 ;
        RECT 69.845 151.755 71.500 152.045 ;
        RECT 69.910 151.415 71.500 151.585 ;
        RECT 69.910 151.295 70.080 151.415 ;
        RECT 69.355 151.125 70.080 151.295 ;
        RECT 68.915 150.390 69.085 151.125 ;
        RECT 69.355 150.955 69.525 151.125 ;
        RECT 70.270 151.075 70.985 151.245 ;
        RECT 71.180 151.125 71.500 151.415 ;
        RECT 71.675 151.125 72.015 152.095 ;
        RECT 72.185 151.125 72.355 152.265 ;
        RECT 72.625 151.465 72.875 152.265 ;
        RECT 73.520 151.295 73.850 152.095 ;
        RECT 74.150 151.465 74.480 152.265 ;
        RECT 74.650 151.295 74.980 152.095 ;
        RECT 72.545 151.125 74.980 151.295 ;
        RECT 75.730 151.285 75.985 151.955 ;
        RECT 76.165 151.465 76.450 152.265 ;
        RECT 76.630 151.545 76.960 152.055 ;
        RECT 69.255 150.625 69.525 150.955 ;
        RECT 69.695 150.625 70.100 150.955 ;
        RECT 70.270 150.625 70.980 151.075 ;
        RECT 69.355 150.455 69.525 150.625 ;
        RECT 68.915 150.045 69.185 150.390 ;
        RECT 69.355 150.285 70.965 150.455 ;
        RECT 71.150 150.385 71.500 150.955 ;
        RECT 71.675 150.565 71.850 151.125 ;
        RECT 72.545 150.875 72.715 151.125 ;
        RECT 72.020 150.705 72.715 150.875 ;
        RECT 72.890 150.705 73.310 150.905 ;
        RECT 73.480 150.705 73.810 150.905 ;
        RECT 73.980 150.705 74.310 150.905 ;
        RECT 71.675 150.515 71.905 150.565 ;
        RECT 69.375 149.715 69.755 150.115 ;
        RECT 69.925 149.935 70.095 150.285 ;
        RECT 70.265 149.715 70.595 150.115 ;
        RECT 70.795 149.935 70.965 150.285 ;
        RECT 71.165 149.715 71.495 150.215 ;
        RECT 71.675 149.885 72.015 150.515 ;
        RECT 72.185 149.715 72.435 150.515 ;
        RECT 72.625 150.365 73.850 150.535 ;
        RECT 72.625 149.885 72.955 150.365 ;
        RECT 73.125 149.715 73.350 150.175 ;
        RECT 73.520 149.885 73.850 150.365 ;
        RECT 74.480 150.495 74.650 151.125 ;
        RECT 74.835 150.705 75.185 150.955 ;
        RECT 74.480 149.885 74.980 150.495 ;
        RECT 75.730 150.425 75.910 151.285 ;
        RECT 76.630 150.955 76.880 151.545 ;
        RECT 77.230 151.395 77.400 152.005 ;
        RECT 77.570 151.575 77.900 152.265 ;
        RECT 78.130 151.715 78.370 152.005 ;
        RECT 78.570 151.885 78.990 152.265 ;
        RECT 79.170 151.795 79.800 152.045 ;
        RECT 80.270 151.885 80.600 152.265 ;
        RECT 79.170 151.715 79.340 151.795 ;
        RECT 80.770 151.715 80.940 152.005 ;
        RECT 81.120 151.885 81.500 152.265 ;
        RECT 81.740 151.880 82.570 152.050 ;
        RECT 78.130 151.545 79.340 151.715 ;
        RECT 76.080 150.625 76.880 150.955 ;
        RECT 75.730 150.225 75.985 150.425 ;
        RECT 75.645 150.055 75.985 150.225 ;
        RECT 75.730 149.895 75.985 150.055 ;
        RECT 76.165 149.715 76.450 150.175 ;
        RECT 76.630 149.975 76.880 150.625 ;
        RECT 77.080 151.375 77.400 151.395 ;
        RECT 77.080 151.205 79.000 151.375 ;
        RECT 77.080 150.310 77.270 151.205 ;
        RECT 79.170 151.035 79.340 151.545 ;
        RECT 79.510 151.285 80.030 151.595 ;
        RECT 77.440 150.865 79.340 151.035 ;
        RECT 77.440 150.805 77.770 150.865 ;
        RECT 77.920 150.635 78.250 150.695 ;
        RECT 77.590 150.365 78.250 150.635 ;
        RECT 77.080 149.980 77.400 150.310 ;
        RECT 77.580 149.715 78.240 150.195 ;
        RECT 78.440 150.105 78.610 150.865 ;
        RECT 79.510 150.695 79.690 151.105 ;
        RECT 78.780 150.525 79.110 150.645 ;
        RECT 79.860 150.525 80.030 151.285 ;
        RECT 78.780 150.355 80.030 150.525 ;
        RECT 80.200 151.465 81.570 151.715 ;
        RECT 80.200 150.695 80.390 151.465 ;
        RECT 81.320 151.205 81.570 151.465 ;
        RECT 80.560 151.035 80.810 151.195 ;
        RECT 81.740 151.035 81.910 151.880 ;
        RECT 82.805 151.595 82.975 152.095 ;
        RECT 83.145 151.765 83.475 152.265 ;
        RECT 82.080 151.205 82.580 151.585 ;
        RECT 82.805 151.425 83.500 151.595 ;
        RECT 80.560 150.865 81.910 151.035 ;
        RECT 81.490 150.825 81.910 150.865 ;
        RECT 80.200 150.355 80.620 150.695 ;
        RECT 80.910 150.365 81.320 150.695 ;
        RECT 78.440 149.935 79.290 150.105 ;
        RECT 79.850 149.715 80.170 150.175 ;
        RECT 80.370 149.925 80.620 150.355 ;
        RECT 80.910 149.715 81.320 150.155 ;
        RECT 81.490 150.095 81.660 150.825 ;
        RECT 81.830 150.275 82.180 150.645 ;
        RECT 82.360 150.335 82.580 151.205 ;
        RECT 82.750 150.635 83.160 151.255 ;
        RECT 83.330 150.455 83.500 151.425 ;
        RECT 82.805 150.265 83.500 150.455 ;
        RECT 81.490 149.895 82.505 150.095 ;
        RECT 82.805 149.935 82.975 150.265 ;
        RECT 83.145 149.715 83.475 150.095 ;
        RECT 83.690 149.975 83.915 152.095 ;
        RECT 84.085 151.765 84.415 152.265 ;
        RECT 84.585 151.595 84.755 152.095 ;
        RECT 84.090 151.425 84.755 151.595 ;
        RECT 84.090 150.435 84.320 151.425 ;
        RECT 84.490 150.605 84.840 151.255 ;
        RECT 85.975 151.125 86.205 152.265 ;
        RECT 86.375 151.115 86.705 152.095 ;
        RECT 86.875 151.125 87.085 152.265 ;
        RECT 85.955 150.705 86.285 150.955 ;
        RECT 84.090 150.265 84.755 150.435 ;
        RECT 84.085 149.715 84.415 150.095 ;
        RECT 84.585 149.975 84.755 150.265 ;
        RECT 85.975 149.715 86.205 150.535 ;
        RECT 86.455 150.515 86.705 151.115 ;
        RECT 87.315 151.100 87.605 152.265 ;
        RECT 88.235 151.190 88.505 152.095 ;
        RECT 88.675 151.505 89.005 152.265 ;
        RECT 89.185 151.335 89.355 152.095 ;
        RECT 86.375 149.885 86.705 150.515 ;
        RECT 86.875 149.715 87.085 150.535 ;
        RECT 87.315 149.715 87.605 150.440 ;
        RECT 88.235 150.390 88.405 151.190 ;
        RECT 88.690 151.165 89.355 151.335 ;
        RECT 88.690 151.020 88.860 151.165 ;
        RECT 88.575 150.690 88.860 151.020 ;
        RECT 89.615 151.125 89.885 152.095 ;
        RECT 90.095 151.465 90.375 152.265 ;
        RECT 90.545 151.755 92.200 152.045 ;
        RECT 90.610 151.415 92.200 151.585 ;
        RECT 90.610 151.295 90.780 151.415 ;
        RECT 90.055 151.125 90.780 151.295 ;
        RECT 88.690 150.435 88.860 150.690 ;
        RECT 89.095 150.615 89.425 150.985 ;
        RECT 88.235 149.885 88.495 150.390 ;
        RECT 88.690 150.265 89.355 150.435 ;
        RECT 88.675 149.715 89.005 150.095 ;
        RECT 89.185 149.885 89.355 150.265 ;
        RECT 89.615 150.390 89.785 151.125 ;
        RECT 90.055 150.955 90.225 151.125 ;
        RECT 89.955 150.625 90.225 150.955 ;
        RECT 90.395 150.625 90.800 150.955 ;
        RECT 90.970 150.625 91.680 151.245 ;
        RECT 91.880 151.125 92.200 151.415 ;
        RECT 92.375 151.125 92.645 152.095 ;
        RECT 92.855 151.465 93.135 152.265 ;
        RECT 93.305 151.755 94.960 152.045 ;
        RECT 93.370 151.415 94.960 151.585 ;
        RECT 93.370 151.295 93.540 151.415 ;
        RECT 92.815 151.125 93.540 151.295 ;
        RECT 90.055 150.455 90.225 150.625 ;
        RECT 89.615 150.045 89.885 150.390 ;
        RECT 90.055 150.285 91.665 150.455 ;
        RECT 91.850 150.385 92.200 150.955 ;
        RECT 92.375 150.390 92.545 151.125 ;
        RECT 92.815 150.955 92.985 151.125 ;
        RECT 93.730 151.075 94.445 151.245 ;
        RECT 94.640 151.125 94.960 151.415 ;
        RECT 95.135 151.125 95.475 152.095 ;
        RECT 95.645 151.125 95.815 152.265 ;
        RECT 96.085 151.465 96.335 152.265 ;
        RECT 96.980 151.295 97.310 152.095 ;
        RECT 97.610 151.465 97.940 152.265 ;
        RECT 98.110 151.295 98.440 152.095 ;
        RECT 96.005 151.125 98.440 151.295 ;
        RECT 98.815 151.125 99.155 152.095 ;
        RECT 99.325 151.125 99.495 152.265 ;
        RECT 99.765 151.465 100.015 152.265 ;
        RECT 100.660 151.295 100.990 152.095 ;
        RECT 101.290 151.465 101.620 152.265 ;
        RECT 101.790 151.295 102.120 152.095 ;
        RECT 99.685 151.125 102.120 151.295 ;
        RECT 103.415 151.505 103.930 151.915 ;
        RECT 104.165 151.505 104.335 152.265 ;
        RECT 104.505 151.925 106.535 152.095 ;
        RECT 92.715 150.625 92.985 150.955 ;
        RECT 93.155 150.625 93.560 150.955 ;
        RECT 93.730 150.625 94.440 151.075 ;
        RECT 92.815 150.455 92.985 150.625 ;
        RECT 90.075 149.715 90.455 150.115 ;
        RECT 90.625 149.935 90.795 150.285 ;
        RECT 90.965 149.715 91.295 150.115 ;
        RECT 91.495 149.935 91.665 150.285 ;
        RECT 91.865 149.715 92.195 150.215 ;
        RECT 92.375 150.045 92.645 150.390 ;
        RECT 92.815 150.285 94.425 150.455 ;
        RECT 94.610 150.385 94.960 150.955 ;
        RECT 95.135 150.565 95.310 151.125 ;
        RECT 96.005 150.875 96.175 151.125 ;
        RECT 95.480 150.705 96.175 150.875 ;
        RECT 96.350 150.705 96.770 150.905 ;
        RECT 96.940 150.705 97.270 150.905 ;
        RECT 97.440 150.705 97.770 150.905 ;
        RECT 95.135 150.515 95.365 150.565 ;
        RECT 92.835 149.715 93.215 150.115 ;
        RECT 93.385 149.935 93.555 150.285 ;
        RECT 93.725 149.715 94.055 150.115 ;
        RECT 94.255 149.935 94.425 150.285 ;
        RECT 94.625 149.715 94.955 150.215 ;
        RECT 95.135 149.885 95.475 150.515 ;
        RECT 95.645 149.715 95.895 150.515 ;
        RECT 96.085 150.365 97.310 150.535 ;
        RECT 96.085 149.885 96.415 150.365 ;
        RECT 96.585 149.715 96.810 150.175 ;
        RECT 96.980 149.885 97.310 150.365 ;
        RECT 97.940 150.495 98.110 151.125 ;
        RECT 98.295 150.705 98.645 150.955 ;
        RECT 98.815 150.515 98.990 151.125 ;
        RECT 99.685 150.875 99.855 151.125 ;
        RECT 99.160 150.705 99.855 150.875 ;
        RECT 100.030 150.705 100.450 150.905 ;
        RECT 100.620 150.705 100.950 150.905 ;
        RECT 101.120 150.705 101.450 150.905 ;
        RECT 97.940 149.885 98.440 150.495 ;
        RECT 98.815 149.885 99.155 150.515 ;
        RECT 99.325 149.715 99.575 150.515 ;
        RECT 99.765 150.365 100.990 150.535 ;
        RECT 99.765 149.885 100.095 150.365 ;
        RECT 100.265 149.715 100.490 150.175 ;
        RECT 100.660 149.885 100.990 150.365 ;
        RECT 101.620 150.495 101.790 151.125 ;
        RECT 101.975 150.705 102.325 150.955 ;
        RECT 103.415 150.695 103.755 151.505 ;
        RECT 104.505 151.260 104.675 151.925 ;
        RECT 105.070 151.585 106.195 151.755 ;
        RECT 103.925 151.070 104.675 151.260 ;
        RECT 104.845 151.245 105.855 151.415 ;
        RECT 103.415 150.525 104.645 150.695 ;
        RECT 101.620 149.885 102.120 150.495 ;
        RECT 103.690 149.920 103.935 150.525 ;
        RECT 104.155 149.715 104.665 150.250 ;
        RECT 104.845 149.885 105.035 151.245 ;
        RECT 105.205 150.905 105.480 151.045 ;
        RECT 105.205 150.735 105.485 150.905 ;
        RECT 105.205 149.885 105.480 150.735 ;
        RECT 105.685 150.445 105.855 151.245 ;
        RECT 106.025 150.455 106.195 151.585 ;
        RECT 106.365 150.955 106.535 151.925 ;
        RECT 106.705 151.125 106.875 152.265 ;
        RECT 107.045 151.125 107.380 152.095 ;
        RECT 108.565 151.335 108.735 152.095 ;
        RECT 108.915 151.505 109.245 152.265 ;
        RECT 108.565 151.165 109.230 151.335 ;
        RECT 109.415 151.190 109.685 152.095 ;
        RECT 106.365 150.625 106.560 150.955 ;
        RECT 106.785 150.625 107.040 150.955 ;
        RECT 106.785 150.455 106.955 150.625 ;
        RECT 107.210 150.455 107.380 151.125 ;
        RECT 109.060 151.020 109.230 151.165 ;
        RECT 108.495 150.615 108.825 150.985 ;
        RECT 109.060 150.690 109.345 151.020 ;
        RECT 106.025 150.285 106.955 150.455 ;
        RECT 106.025 150.250 106.200 150.285 ;
        RECT 105.670 149.885 106.200 150.250 ;
        RECT 106.625 149.715 106.955 150.115 ;
        RECT 107.125 149.885 107.380 150.455 ;
        RECT 109.060 150.435 109.230 150.690 ;
        RECT 108.565 150.265 109.230 150.435 ;
        RECT 109.515 150.390 109.685 151.190 ;
        RECT 110.315 151.175 111.985 152.265 ;
        RECT 112.155 151.175 113.365 152.265 ;
        RECT 110.315 150.655 111.065 151.175 ;
        RECT 111.235 150.485 111.985 151.005 ;
        RECT 112.155 150.635 112.675 151.175 ;
        RECT 108.565 149.885 108.735 150.265 ;
        RECT 108.915 149.715 109.245 150.095 ;
        RECT 109.425 149.885 109.685 150.390 ;
        RECT 110.315 149.715 111.985 150.485 ;
        RECT 112.845 150.465 113.365 151.005 ;
        RECT 112.155 149.715 113.365 150.465 ;
        RECT 15.010 149.545 113.450 149.715 ;
        RECT 15.095 148.795 16.305 149.545 ;
        RECT 15.095 148.255 15.615 148.795 ;
        RECT 16.475 148.775 18.145 149.545 ;
        RECT 15.785 148.085 16.305 148.625 ;
        RECT 15.095 146.995 16.305 148.085 ;
        RECT 16.475 148.085 17.225 148.605 ;
        RECT 17.395 148.255 18.145 148.775 ;
        RECT 18.355 148.725 18.585 149.545 ;
        RECT 18.755 148.745 19.085 149.375 ;
        RECT 18.335 148.305 18.665 148.555 ;
        RECT 18.835 148.145 19.085 148.745 ;
        RECT 19.255 148.725 19.465 149.545 ;
        RECT 19.785 148.995 19.955 149.375 ;
        RECT 20.135 149.165 20.465 149.545 ;
        RECT 19.785 148.825 20.450 148.995 ;
        RECT 20.645 148.870 20.905 149.375 ;
        RECT 19.715 148.275 20.045 148.645 ;
        RECT 20.280 148.570 20.450 148.825 ;
        RECT 16.475 146.995 18.145 148.085 ;
        RECT 18.355 146.995 18.585 148.135 ;
        RECT 18.755 147.165 19.085 148.145 ;
        RECT 20.280 148.240 20.565 148.570 ;
        RECT 19.255 146.995 19.465 148.135 ;
        RECT 20.280 148.095 20.450 148.240 ;
        RECT 19.785 147.925 20.450 148.095 ;
        RECT 20.735 148.070 20.905 148.870 ;
        RECT 21.135 148.725 21.345 149.545 ;
        RECT 21.515 148.745 21.845 149.375 ;
        RECT 21.515 148.145 21.765 148.745 ;
        RECT 22.015 148.725 22.245 149.545 ;
        RECT 22.915 148.820 23.205 149.545 ;
        RECT 23.925 148.995 24.095 149.375 ;
        RECT 24.275 149.165 24.605 149.545 ;
        RECT 23.925 148.825 24.590 148.995 ;
        RECT 24.785 148.870 25.045 149.375 ;
        RECT 25.590 149.205 25.845 149.365 ;
        RECT 25.505 149.035 25.845 149.205 ;
        RECT 26.025 149.085 26.310 149.545 ;
        RECT 21.935 148.305 22.265 148.555 ;
        RECT 23.855 148.275 24.185 148.645 ;
        RECT 24.420 148.570 24.590 148.825 ;
        RECT 24.420 148.240 24.705 148.570 ;
        RECT 19.785 147.165 19.955 147.925 ;
        RECT 20.135 146.995 20.465 147.755 ;
        RECT 20.635 147.165 20.905 148.070 ;
        RECT 21.135 146.995 21.345 148.135 ;
        RECT 21.515 147.165 21.845 148.145 ;
        RECT 22.015 146.995 22.245 148.135 ;
        RECT 22.915 146.995 23.205 148.160 ;
        RECT 24.420 148.095 24.590 148.240 ;
        RECT 23.925 147.925 24.590 148.095 ;
        RECT 24.875 148.070 25.045 148.870 ;
        RECT 23.925 147.165 24.095 147.925 ;
        RECT 24.275 146.995 24.605 147.755 ;
        RECT 24.775 147.165 25.045 148.070 ;
        RECT 25.590 148.835 25.845 149.035 ;
        RECT 25.590 147.975 25.770 148.835 ;
        RECT 26.490 148.635 26.740 149.285 ;
        RECT 25.940 148.305 26.740 148.635 ;
        RECT 25.590 147.305 25.845 147.975 ;
        RECT 26.025 146.995 26.310 147.795 ;
        RECT 26.490 147.715 26.740 148.305 ;
        RECT 26.940 148.950 27.260 149.280 ;
        RECT 27.440 149.065 28.100 149.545 ;
        RECT 28.300 149.155 29.150 149.325 ;
        RECT 26.940 148.055 27.130 148.950 ;
        RECT 27.450 148.625 28.110 148.895 ;
        RECT 27.780 148.565 28.110 148.625 ;
        RECT 27.300 148.395 27.630 148.455 ;
        RECT 28.300 148.395 28.470 149.155 ;
        RECT 29.710 149.085 30.030 149.545 ;
        RECT 30.230 148.905 30.480 149.335 ;
        RECT 30.770 149.105 31.180 149.545 ;
        RECT 31.350 149.165 32.365 149.365 ;
        RECT 28.640 148.735 29.890 148.905 ;
        RECT 28.640 148.615 28.970 148.735 ;
        RECT 27.300 148.225 29.200 148.395 ;
        RECT 26.940 147.885 28.860 148.055 ;
        RECT 26.940 147.865 27.260 147.885 ;
        RECT 26.490 147.205 26.820 147.715 ;
        RECT 27.090 147.255 27.260 147.865 ;
        RECT 29.030 147.715 29.200 148.225 ;
        RECT 29.370 148.155 29.550 148.565 ;
        RECT 29.720 147.975 29.890 148.735 ;
        RECT 27.430 146.995 27.760 147.685 ;
        RECT 27.990 147.545 29.200 147.715 ;
        RECT 29.370 147.665 29.890 147.975 ;
        RECT 30.060 148.565 30.480 148.905 ;
        RECT 30.770 148.565 31.180 148.895 ;
        RECT 30.060 147.795 30.250 148.565 ;
        RECT 31.350 148.435 31.520 149.165 ;
        RECT 32.665 148.995 32.835 149.325 ;
        RECT 33.005 149.165 33.335 149.545 ;
        RECT 31.690 148.615 32.040 148.985 ;
        RECT 31.350 148.395 31.770 148.435 ;
        RECT 30.420 148.225 31.770 148.395 ;
        RECT 30.420 148.065 30.670 148.225 ;
        RECT 31.180 147.795 31.430 148.055 ;
        RECT 30.060 147.545 31.430 147.795 ;
        RECT 27.990 147.255 28.230 147.545 ;
        RECT 29.030 147.465 29.200 147.545 ;
        RECT 28.430 146.995 28.850 147.375 ;
        RECT 29.030 147.215 29.660 147.465 ;
        RECT 30.130 146.995 30.460 147.375 ;
        RECT 30.630 147.255 30.800 147.545 ;
        RECT 31.600 147.380 31.770 148.225 ;
        RECT 32.220 148.055 32.440 148.925 ;
        RECT 32.665 148.805 33.360 148.995 ;
        RECT 31.940 147.675 32.440 148.055 ;
        RECT 32.610 148.005 33.020 148.625 ;
        RECT 33.190 147.835 33.360 148.805 ;
        RECT 32.665 147.665 33.360 147.835 ;
        RECT 30.980 146.995 31.360 147.375 ;
        RECT 31.600 147.210 32.430 147.380 ;
        RECT 32.665 147.165 32.835 147.665 ;
        RECT 33.005 146.995 33.335 147.495 ;
        RECT 33.550 147.165 33.775 149.285 ;
        RECT 33.945 149.165 34.275 149.545 ;
        RECT 34.445 148.995 34.615 149.285 ;
        RECT 33.950 148.825 34.615 148.995 ;
        RECT 33.950 147.835 34.180 148.825 ;
        RECT 34.875 148.795 36.085 149.545 ;
        RECT 34.350 148.005 34.700 148.655 ;
        RECT 34.875 148.085 35.395 148.625 ;
        RECT 35.565 148.255 36.085 148.795 ;
        RECT 36.255 148.870 36.525 149.215 ;
        RECT 36.715 149.145 37.095 149.545 ;
        RECT 37.265 148.975 37.435 149.325 ;
        RECT 37.605 149.145 37.935 149.545 ;
        RECT 38.135 148.975 38.305 149.325 ;
        RECT 38.505 149.045 38.835 149.545 ;
        RECT 36.255 148.135 36.425 148.870 ;
        RECT 36.695 148.805 38.305 148.975 ;
        RECT 36.695 148.635 36.865 148.805 ;
        RECT 36.595 148.305 36.865 148.635 ;
        RECT 37.035 148.305 37.440 148.635 ;
        RECT 36.695 148.135 36.865 148.305 ;
        RECT 37.610 148.185 38.320 148.635 ;
        RECT 38.490 148.305 38.840 148.875 ;
        RECT 39.015 148.870 39.285 149.215 ;
        RECT 39.475 149.145 39.855 149.545 ;
        RECT 40.025 148.975 40.195 149.325 ;
        RECT 40.365 149.145 40.695 149.545 ;
        RECT 40.895 148.975 41.065 149.325 ;
        RECT 41.265 149.045 41.595 149.545 ;
        RECT 41.785 149.045 42.115 149.545 ;
        RECT 33.950 147.665 34.615 147.835 ;
        RECT 33.945 146.995 34.275 147.495 ;
        RECT 34.445 147.165 34.615 147.665 ;
        RECT 34.875 146.995 36.085 148.085 ;
        RECT 36.255 147.165 36.525 148.135 ;
        RECT 36.695 147.965 37.420 148.135 ;
        RECT 37.610 148.015 38.325 148.185 ;
        RECT 39.015 148.135 39.185 148.870 ;
        RECT 39.455 148.805 41.065 148.975 ;
        RECT 42.315 148.975 42.485 149.325 ;
        RECT 42.685 149.145 43.015 149.545 ;
        RECT 43.185 148.975 43.355 149.325 ;
        RECT 43.525 149.145 43.905 149.545 ;
        RECT 39.455 148.635 39.625 148.805 ;
        RECT 39.355 148.305 39.625 148.635 ;
        RECT 39.795 148.305 40.200 148.635 ;
        RECT 39.455 148.135 39.625 148.305 ;
        RECT 37.250 147.845 37.420 147.965 ;
        RECT 38.520 147.845 38.840 148.135 ;
        RECT 36.735 146.995 37.015 147.795 ;
        RECT 37.250 147.675 38.840 147.845 ;
        RECT 37.185 147.215 38.840 147.505 ;
        RECT 39.015 147.165 39.285 148.135 ;
        RECT 39.455 147.965 40.180 148.135 ;
        RECT 40.370 148.015 41.080 148.635 ;
        RECT 41.250 148.305 41.600 148.875 ;
        RECT 41.780 148.305 42.130 148.875 ;
        RECT 42.315 148.805 43.925 148.975 ;
        RECT 44.095 148.870 44.365 149.215 ;
        RECT 43.755 148.635 43.925 148.805 ;
        RECT 42.300 148.185 43.010 148.635 ;
        RECT 43.180 148.305 43.585 148.635 ;
        RECT 43.755 148.305 44.025 148.635 ;
        RECT 40.010 147.845 40.180 147.965 ;
        RECT 41.280 147.845 41.600 148.135 ;
        RECT 39.495 146.995 39.775 147.795 ;
        RECT 40.010 147.675 41.600 147.845 ;
        RECT 41.780 147.845 42.100 148.135 ;
        RECT 42.295 148.015 43.010 148.185 ;
        RECT 43.755 148.135 43.925 148.305 ;
        RECT 44.195 148.135 44.365 148.870 ;
        RECT 44.810 148.735 45.055 149.340 ;
        RECT 45.275 149.010 45.785 149.545 ;
        RECT 43.200 147.965 43.925 148.135 ;
        RECT 43.200 147.845 43.370 147.965 ;
        RECT 41.780 147.675 43.370 147.845 ;
        RECT 39.945 147.215 41.600 147.505 ;
        RECT 41.780 147.215 43.435 147.505 ;
        RECT 43.605 146.995 43.885 147.795 ;
        RECT 44.095 147.165 44.365 148.135 ;
        RECT 44.535 148.565 45.765 148.735 ;
        RECT 44.535 147.755 44.875 148.565 ;
        RECT 45.045 148.000 45.795 148.190 ;
        RECT 44.535 147.345 45.050 147.755 ;
        RECT 45.285 146.995 45.455 147.755 ;
        RECT 45.625 147.335 45.795 148.000 ;
        RECT 45.965 148.015 46.155 149.375 ;
        RECT 46.325 149.205 46.600 149.375 ;
        RECT 46.325 149.035 46.605 149.205 ;
        RECT 46.325 148.215 46.600 149.035 ;
        RECT 46.790 149.010 47.320 149.375 ;
        RECT 47.745 149.145 48.075 149.545 ;
        RECT 47.145 148.975 47.320 149.010 ;
        RECT 46.805 148.015 46.975 148.815 ;
        RECT 45.965 147.845 46.975 148.015 ;
        RECT 47.145 148.805 48.075 148.975 ;
        RECT 48.245 148.805 48.500 149.375 ;
        RECT 48.675 148.820 48.965 149.545 ;
        RECT 47.145 147.675 47.315 148.805 ;
        RECT 47.905 148.635 48.075 148.805 ;
        RECT 46.190 147.505 47.315 147.675 ;
        RECT 47.485 148.305 47.680 148.635 ;
        RECT 47.905 148.305 48.160 148.635 ;
        RECT 47.485 147.335 47.655 148.305 ;
        RECT 48.330 148.135 48.500 148.805 ;
        RECT 49.135 148.795 50.345 149.545 ;
        RECT 50.520 149.000 55.865 149.545 ;
        RECT 45.625 147.165 47.655 147.335 ;
        RECT 47.825 146.995 47.995 148.135 ;
        RECT 48.165 147.165 48.500 148.135 ;
        RECT 48.675 146.995 48.965 148.160 ;
        RECT 49.135 148.085 49.655 148.625 ;
        RECT 49.825 148.255 50.345 148.795 ;
        RECT 49.135 146.995 50.345 148.085 ;
        RECT 52.110 147.430 52.460 148.680 ;
        RECT 53.940 148.170 54.280 149.000 ;
        RECT 56.125 148.995 56.295 149.375 ;
        RECT 56.475 149.165 56.805 149.545 ;
        RECT 56.125 148.825 56.790 148.995 ;
        RECT 56.985 148.870 57.245 149.375 ;
        RECT 56.055 148.275 56.385 148.645 ;
        RECT 56.620 148.570 56.790 148.825 ;
        RECT 56.620 148.240 56.905 148.570 ;
        RECT 56.620 148.095 56.790 148.240 ;
        RECT 56.125 147.925 56.790 148.095 ;
        RECT 57.075 148.070 57.245 148.870 ;
        RECT 57.415 148.795 58.625 149.545 ;
        RECT 59.170 149.205 59.425 149.365 ;
        RECT 59.085 149.035 59.425 149.205 ;
        RECT 59.605 149.085 59.890 149.545 ;
        RECT 50.520 146.995 55.865 147.430 ;
        RECT 56.125 147.165 56.295 147.925 ;
        RECT 56.475 146.995 56.805 147.755 ;
        RECT 56.975 147.165 57.245 148.070 ;
        RECT 57.415 148.085 57.935 148.625 ;
        RECT 58.105 148.255 58.625 148.795 ;
        RECT 59.170 148.835 59.425 149.035 ;
        RECT 57.415 146.995 58.625 148.085 ;
        RECT 59.170 147.975 59.350 148.835 ;
        RECT 60.070 148.635 60.320 149.285 ;
        RECT 59.520 148.305 60.320 148.635 ;
        RECT 59.170 147.305 59.425 147.975 ;
        RECT 59.605 146.995 59.890 147.795 ;
        RECT 60.070 147.715 60.320 148.305 ;
        RECT 60.520 148.950 60.840 149.280 ;
        RECT 61.020 149.065 61.680 149.545 ;
        RECT 61.880 149.155 62.730 149.325 ;
        RECT 60.520 148.055 60.710 148.950 ;
        RECT 61.030 148.625 61.690 148.895 ;
        RECT 61.360 148.565 61.690 148.625 ;
        RECT 60.880 148.395 61.210 148.455 ;
        RECT 61.880 148.395 62.050 149.155 ;
        RECT 63.290 149.085 63.610 149.545 ;
        RECT 63.810 148.905 64.060 149.335 ;
        RECT 64.350 149.105 64.760 149.545 ;
        RECT 64.930 149.165 65.945 149.365 ;
        RECT 62.220 148.735 63.470 148.905 ;
        RECT 62.220 148.615 62.550 148.735 ;
        RECT 60.880 148.225 62.780 148.395 ;
        RECT 60.520 147.885 62.440 148.055 ;
        RECT 60.520 147.865 60.840 147.885 ;
        RECT 60.070 147.205 60.400 147.715 ;
        RECT 60.670 147.255 60.840 147.865 ;
        RECT 62.610 147.715 62.780 148.225 ;
        RECT 62.950 148.155 63.130 148.565 ;
        RECT 63.300 147.975 63.470 148.735 ;
        RECT 61.010 146.995 61.340 147.685 ;
        RECT 61.570 147.545 62.780 147.715 ;
        RECT 62.950 147.665 63.470 147.975 ;
        RECT 63.640 148.565 64.060 148.905 ;
        RECT 64.350 148.565 64.760 148.895 ;
        RECT 63.640 147.795 63.830 148.565 ;
        RECT 64.930 148.435 65.100 149.165 ;
        RECT 66.245 148.995 66.415 149.325 ;
        RECT 66.585 149.165 66.915 149.545 ;
        RECT 65.270 148.615 65.620 148.985 ;
        RECT 64.930 148.395 65.350 148.435 ;
        RECT 64.000 148.225 65.350 148.395 ;
        RECT 64.000 148.065 64.250 148.225 ;
        RECT 64.760 147.795 65.010 148.055 ;
        RECT 63.640 147.545 65.010 147.795 ;
        RECT 61.570 147.255 61.810 147.545 ;
        RECT 62.610 147.465 62.780 147.545 ;
        RECT 62.010 146.995 62.430 147.375 ;
        RECT 62.610 147.215 63.240 147.465 ;
        RECT 63.710 146.995 64.040 147.375 ;
        RECT 64.210 147.255 64.380 147.545 ;
        RECT 65.180 147.380 65.350 148.225 ;
        RECT 65.800 148.055 66.020 148.925 ;
        RECT 66.245 148.805 66.940 148.995 ;
        RECT 65.520 147.675 66.020 148.055 ;
        RECT 66.190 148.005 66.600 148.625 ;
        RECT 66.770 147.835 66.940 148.805 ;
        RECT 66.245 147.665 66.940 147.835 ;
        RECT 64.560 146.995 64.940 147.375 ;
        RECT 65.180 147.210 66.010 147.380 ;
        RECT 66.245 147.165 66.415 147.665 ;
        RECT 66.585 146.995 66.915 147.495 ;
        RECT 67.130 147.165 67.355 149.285 ;
        RECT 67.525 149.165 67.855 149.545 ;
        RECT 68.025 148.995 68.195 149.285 ;
        RECT 67.530 148.825 68.195 148.995 ;
        RECT 68.545 148.995 68.715 149.375 ;
        RECT 68.930 149.165 69.260 149.545 ;
        RECT 68.545 148.825 69.260 148.995 ;
        RECT 67.530 147.835 67.760 148.825 ;
        RECT 67.930 148.005 68.280 148.655 ;
        RECT 68.455 148.275 68.810 148.645 ;
        RECT 69.090 148.635 69.260 148.825 ;
        RECT 69.430 148.800 69.685 149.375 ;
        RECT 69.090 148.305 69.345 148.635 ;
        RECT 69.090 148.095 69.260 148.305 ;
        RECT 68.545 147.925 69.260 148.095 ;
        RECT 69.515 148.070 69.685 148.800 ;
        RECT 69.860 148.705 70.120 149.545 ;
        RECT 70.755 148.745 71.095 149.375 ;
        RECT 71.265 148.745 71.515 149.545 ;
        RECT 71.705 148.895 72.035 149.375 ;
        RECT 72.205 149.085 72.430 149.545 ;
        RECT 72.600 148.895 72.930 149.375 ;
        RECT 67.530 147.665 68.195 147.835 ;
        RECT 67.525 146.995 67.855 147.495 ;
        RECT 68.025 147.165 68.195 147.665 ;
        RECT 68.545 147.165 68.715 147.925 ;
        RECT 68.930 146.995 69.260 147.755 ;
        RECT 69.430 147.165 69.685 148.070 ;
        RECT 69.860 146.995 70.120 148.145 ;
        RECT 70.755 148.135 70.930 148.745 ;
        RECT 71.705 148.725 72.930 148.895 ;
        RECT 73.560 148.765 74.060 149.375 ;
        RECT 74.435 148.820 74.725 149.545 ;
        RECT 71.100 148.385 71.795 148.555 ;
        RECT 71.625 148.135 71.795 148.385 ;
        RECT 71.970 148.355 72.390 148.555 ;
        RECT 72.560 148.355 72.890 148.555 ;
        RECT 73.060 148.355 73.390 148.555 ;
        RECT 73.560 148.135 73.730 148.765 ;
        RECT 75.630 148.735 75.875 149.340 ;
        RECT 76.095 149.010 76.605 149.545 ;
        RECT 75.355 148.565 76.585 148.735 ;
        RECT 73.915 148.305 74.265 148.555 ;
        RECT 70.755 147.165 71.095 148.135 ;
        RECT 71.265 146.995 71.435 148.135 ;
        RECT 71.625 147.965 74.060 148.135 ;
        RECT 71.705 146.995 71.955 147.795 ;
        RECT 72.600 147.165 72.930 147.965 ;
        RECT 73.230 146.995 73.560 147.795 ;
        RECT 73.730 147.165 74.060 147.965 ;
        RECT 74.435 146.995 74.725 148.160 ;
        RECT 75.355 147.755 75.695 148.565 ;
        RECT 75.865 148.000 76.615 148.190 ;
        RECT 75.355 147.345 75.870 147.755 ;
        RECT 76.105 146.995 76.275 147.755 ;
        RECT 76.445 147.335 76.615 148.000 ;
        RECT 76.785 148.015 76.975 149.375 ;
        RECT 77.145 149.205 77.420 149.375 ;
        RECT 77.145 149.035 77.425 149.205 ;
        RECT 77.145 148.215 77.420 149.035 ;
        RECT 77.610 149.010 78.140 149.375 ;
        RECT 78.565 149.145 78.895 149.545 ;
        RECT 77.965 148.975 78.140 149.010 ;
        RECT 77.625 148.015 77.795 148.815 ;
        RECT 76.785 147.845 77.795 148.015 ;
        RECT 77.965 148.805 78.895 148.975 ;
        RECT 79.065 148.805 79.320 149.375 ;
        RECT 77.965 147.675 78.135 148.805 ;
        RECT 78.725 148.635 78.895 148.805 ;
        RECT 77.010 147.505 78.135 147.675 ;
        RECT 78.305 148.305 78.500 148.635 ;
        RECT 78.725 148.305 78.980 148.635 ;
        RECT 78.305 147.335 78.475 148.305 ;
        RECT 79.150 148.135 79.320 148.805 ;
        RECT 76.445 147.165 78.475 147.335 ;
        RECT 78.645 146.995 78.815 148.135 ;
        RECT 78.985 147.165 79.320 148.135 ;
        RECT 79.500 148.805 79.755 149.375 ;
        RECT 79.925 149.145 80.255 149.545 ;
        RECT 80.680 149.010 81.210 149.375 ;
        RECT 80.680 148.975 80.855 149.010 ;
        RECT 79.925 148.805 80.855 148.975 ;
        RECT 79.500 148.135 79.670 148.805 ;
        RECT 79.925 148.635 80.095 148.805 ;
        RECT 79.840 148.305 80.095 148.635 ;
        RECT 80.320 148.305 80.515 148.635 ;
        RECT 79.500 147.165 79.835 148.135 ;
        RECT 80.005 146.995 80.175 148.135 ;
        RECT 80.345 147.335 80.515 148.305 ;
        RECT 80.685 147.675 80.855 148.805 ;
        RECT 81.025 148.015 81.195 148.815 ;
        RECT 81.400 148.525 81.675 149.375 ;
        RECT 81.395 148.355 81.675 148.525 ;
        RECT 81.400 148.215 81.675 148.355 ;
        RECT 81.845 148.015 82.035 149.375 ;
        RECT 82.215 149.010 82.725 149.545 ;
        RECT 82.945 148.735 83.190 149.340 ;
        RECT 83.910 148.735 84.155 149.340 ;
        RECT 84.375 149.010 84.885 149.545 ;
        RECT 82.235 148.565 83.465 148.735 ;
        RECT 81.025 147.845 82.035 148.015 ;
        RECT 82.205 148.000 82.955 148.190 ;
        RECT 80.685 147.505 81.810 147.675 ;
        RECT 82.205 147.335 82.375 148.000 ;
        RECT 83.125 147.755 83.465 148.565 ;
        RECT 80.345 147.165 82.375 147.335 ;
        RECT 82.545 146.995 82.715 147.755 ;
        RECT 82.950 147.345 83.465 147.755 ;
        RECT 83.635 148.565 84.865 148.735 ;
        RECT 83.635 147.755 83.975 148.565 ;
        RECT 84.145 148.000 84.895 148.190 ;
        RECT 83.635 147.345 84.150 147.755 ;
        RECT 84.385 146.995 84.555 147.755 ;
        RECT 84.725 147.335 84.895 148.000 ;
        RECT 85.065 148.015 85.255 149.375 ;
        RECT 85.425 148.865 85.700 149.375 ;
        RECT 85.890 149.010 86.420 149.375 ;
        RECT 86.845 149.145 87.175 149.545 ;
        RECT 86.245 148.975 86.420 149.010 ;
        RECT 85.425 148.695 85.705 148.865 ;
        RECT 85.425 148.215 85.700 148.695 ;
        RECT 85.905 148.015 86.075 148.815 ;
        RECT 85.065 147.845 86.075 148.015 ;
        RECT 86.245 148.805 87.175 148.975 ;
        RECT 87.345 148.805 87.600 149.375 ;
        RECT 88.240 149.000 93.585 149.545 ;
        RECT 86.245 147.675 86.415 148.805 ;
        RECT 87.005 148.635 87.175 148.805 ;
        RECT 85.290 147.505 86.415 147.675 ;
        RECT 86.585 148.305 86.780 148.635 ;
        RECT 87.005 148.305 87.260 148.635 ;
        RECT 86.585 147.335 86.755 148.305 ;
        RECT 87.430 148.135 87.600 148.805 ;
        RECT 84.725 147.165 86.755 147.335 ;
        RECT 86.925 146.995 87.095 148.135 ;
        RECT 87.265 147.165 87.600 148.135 ;
        RECT 89.830 147.430 90.180 148.680 ;
        RECT 91.660 148.170 92.000 149.000 ;
        RECT 93.755 148.870 94.025 149.215 ;
        RECT 94.215 149.145 94.595 149.545 ;
        RECT 94.765 148.975 94.935 149.325 ;
        RECT 95.105 149.145 95.435 149.545 ;
        RECT 95.635 148.975 95.805 149.325 ;
        RECT 96.005 149.045 96.335 149.545 ;
        RECT 93.755 148.135 93.925 148.870 ;
        RECT 94.195 148.805 95.805 148.975 ;
        RECT 94.195 148.635 94.365 148.805 ;
        RECT 94.095 148.305 94.365 148.635 ;
        RECT 94.535 148.305 94.940 148.635 ;
        RECT 94.195 148.135 94.365 148.305 ;
        RECT 95.110 148.185 95.820 148.635 ;
        RECT 95.990 148.305 96.340 148.875 ;
        RECT 96.515 148.745 96.855 149.375 ;
        RECT 97.025 148.745 97.275 149.545 ;
        RECT 97.465 148.895 97.795 149.375 ;
        RECT 97.965 149.085 98.190 149.545 ;
        RECT 98.360 148.895 98.690 149.375 ;
        RECT 96.515 148.695 96.745 148.745 ;
        RECT 97.465 148.725 98.690 148.895 ;
        RECT 99.320 148.765 99.820 149.375 ;
        RECT 100.195 148.820 100.485 149.545 ;
        RECT 88.240 146.995 93.585 147.430 ;
        RECT 93.755 147.165 94.025 148.135 ;
        RECT 94.195 147.965 94.920 148.135 ;
        RECT 95.110 148.015 95.825 148.185 ;
        RECT 96.515 148.135 96.690 148.695 ;
        RECT 96.860 148.385 97.555 148.555 ;
        RECT 97.385 148.135 97.555 148.385 ;
        RECT 97.730 148.355 98.150 148.555 ;
        RECT 98.320 148.355 98.650 148.555 ;
        RECT 98.820 148.355 99.150 148.555 ;
        RECT 99.320 148.135 99.490 148.765 ;
        RECT 101.155 148.725 101.385 149.545 ;
        RECT 101.555 148.745 101.885 149.375 ;
        RECT 99.675 148.305 100.025 148.555 ;
        RECT 101.135 148.305 101.465 148.555 ;
        RECT 94.750 147.845 94.920 147.965 ;
        RECT 96.020 147.845 96.340 148.135 ;
        RECT 94.235 146.995 94.515 147.795 ;
        RECT 94.750 147.675 96.340 147.845 ;
        RECT 94.685 147.215 96.340 147.505 ;
        RECT 96.515 147.165 96.855 148.135 ;
        RECT 97.025 146.995 97.195 148.135 ;
        RECT 97.385 147.965 99.820 148.135 ;
        RECT 97.465 146.995 97.715 147.795 ;
        RECT 98.360 147.165 98.690 147.965 ;
        RECT 98.990 146.995 99.320 147.795 ;
        RECT 99.490 147.165 99.820 147.965 ;
        RECT 100.195 146.995 100.485 148.160 ;
        RECT 101.635 148.145 101.885 148.745 ;
        RECT 102.055 148.725 102.265 149.545 ;
        RECT 102.870 148.835 103.125 149.365 ;
        RECT 103.305 149.085 103.590 149.545 ;
        RECT 101.155 146.995 101.385 148.135 ;
        RECT 101.555 147.165 101.885 148.145 ;
        RECT 102.055 146.995 102.265 148.135 ;
        RECT 102.870 147.975 103.050 148.835 ;
        RECT 103.770 148.635 104.020 149.285 ;
        RECT 103.220 148.305 104.020 148.635 ;
        RECT 102.870 147.505 103.125 147.975 ;
        RECT 102.785 147.335 103.125 147.505 ;
        RECT 102.870 147.305 103.125 147.335 ;
        RECT 103.305 146.995 103.590 147.795 ;
        RECT 103.770 147.715 104.020 148.305 ;
        RECT 104.220 148.950 104.540 149.280 ;
        RECT 104.720 149.065 105.380 149.545 ;
        RECT 105.580 149.155 106.430 149.325 ;
        RECT 104.220 148.055 104.410 148.950 ;
        RECT 104.730 148.625 105.390 148.895 ;
        RECT 105.060 148.565 105.390 148.625 ;
        RECT 104.580 148.395 104.910 148.455 ;
        RECT 105.580 148.395 105.750 149.155 ;
        RECT 106.990 149.085 107.310 149.545 ;
        RECT 107.510 148.905 107.760 149.335 ;
        RECT 108.050 149.105 108.460 149.545 ;
        RECT 108.630 149.165 109.645 149.365 ;
        RECT 105.920 148.735 107.170 148.905 ;
        RECT 105.920 148.615 106.250 148.735 ;
        RECT 104.580 148.225 106.480 148.395 ;
        RECT 104.220 147.885 106.140 148.055 ;
        RECT 104.220 147.865 104.540 147.885 ;
        RECT 103.770 147.205 104.100 147.715 ;
        RECT 104.370 147.255 104.540 147.865 ;
        RECT 106.310 147.715 106.480 148.225 ;
        RECT 106.650 148.155 106.830 148.565 ;
        RECT 107.000 147.975 107.170 148.735 ;
        RECT 104.710 146.995 105.040 147.685 ;
        RECT 105.270 147.545 106.480 147.715 ;
        RECT 106.650 147.665 107.170 147.975 ;
        RECT 107.340 148.565 107.760 148.905 ;
        RECT 108.050 148.565 108.460 148.895 ;
        RECT 107.340 147.795 107.530 148.565 ;
        RECT 108.630 148.435 108.800 149.165 ;
        RECT 109.945 148.995 110.115 149.325 ;
        RECT 110.285 149.165 110.615 149.545 ;
        RECT 108.970 148.615 109.320 148.985 ;
        RECT 108.630 148.395 109.050 148.435 ;
        RECT 107.700 148.225 109.050 148.395 ;
        RECT 107.700 148.065 107.950 148.225 ;
        RECT 108.460 147.795 108.710 148.055 ;
        RECT 107.340 147.545 108.710 147.795 ;
        RECT 105.270 147.255 105.510 147.545 ;
        RECT 106.310 147.465 106.480 147.545 ;
        RECT 105.710 146.995 106.130 147.375 ;
        RECT 106.310 147.215 106.940 147.465 ;
        RECT 107.410 146.995 107.740 147.375 ;
        RECT 107.910 147.255 108.080 147.545 ;
        RECT 108.880 147.380 109.050 148.225 ;
        RECT 109.500 148.055 109.720 148.925 ;
        RECT 109.945 148.805 110.640 148.995 ;
        RECT 109.220 147.675 109.720 148.055 ;
        RECT 109.890 148.005 110.300 148.625 ;
        RECT 110.470 147.835 110.640 148.805 ;
        RECT 109.945 147.665 110.640 147.835 ;
        RECT 108.260 146.995 108.640 147.375 ;
        RECT 108.880 147.210 109.710 147.380 ;
        RECT 109.945 147.165 110.115 147.665 ;
        RECT 110.285 146.995 110.615 147.495 ;
        RECT 110.830 147.165 111.055 149.285 ;
        RECT 111.225 149.165 111.555 149.545 ;
        RECT 111.725 148.995 111.895 149.285 ;
        RECT 111.230 148.825 111.895 148.995 ;
        RECT 111.230 147.835 111.460 148.825 ;
        RECT 112.155 148.795 113.365 149.545 ;
        RECT 111.630 148.005 111.980 148.655 ;
        RECT 112.155 148.085 112.675 148.625 ;
        RECT 112.845 148.255 113.365 148.795 ;
        RECT 111.230 147.665 111.895 147.835 ;
        RECT 111.225 146.995 111.555 147.495 ;
        RECT 111.725 147.165 111.895 147.665 ;
        RECT 112.155 146.995 113.365 148.085 ;
        RECT 15.010 146.825 113.450 146.995 ;
        RECT 15.095 145.735 16.305 146.825 ;
        RECT 17.400 146.390 22.745 146.825 ;
        RECT 22.920 146.390 28.265 146.825 ;
        RECT 15.095 145.025 15.615 145.565 ;
        RECT 15.785 145.195 16.305 145.735 ;
        RECT 18.990 145.140 19.340 146.390 ;
        RECT 15.095 144.275 16.305 145.025 ;
        RECT 20.820 144.820 21.160 145.650 ;
        RECT 24.510 145.140 24.860 146.390 ;
        RECT 28.475 145.685 28.705 146.825 ;
        RECT 28.875 145.675 29.205 146.655 ;
        RECT 29.375 145.685 29.585 146.825 ;
        RECT 30.280 146.390 35.625 146.825 ;
        RECT 26.340 144.820 26.680 145.650 ;
        RECT 28.455 145.265 28.785 145.515 ;
        RECT 17.400 144.275 22.745 144.820 ;
        RECT 22.920 144.275 28.265 144.820 ;
        RECT 28.475 144.275 28.705 145.095 ;
        RECT 28.955 145.075 29.205 145.675 ;
        RECT 31.870 145.140 32.220 146.390 ;
        RECT 35.795 145.660 36.085 146.825 ;
        RECT 36.255 145.735 37.925 146.825 ;
        RECT 28.875 144.445 29.205 145.075 ;
        RECT 29.375 144.275 29.585 145.095 ;
        RECT 33.700 144.820 34.040 145.650 ;
        RECT 36.255 145.215 37.005 145.735 ;
        RECT 38.095 145.685 38.435 146.655 ;
        RECT 38.605 145.685 38.775 146.825 ;
        RECT 39.045 146.025 39.295 146.825 ;
        RECT 39.940 145.855 40.270 146.655 ;
        RECT 40.570 146.025 40.900 146.825 ;
        RECT 41.070 145.855 41.400 146.655 ;
        RECT 38.965 145.685 41.400 145.855 ;
        RECT 42.150 145.845 42.405 146.515 ;
        RECT 42.585 146.025 42.870 146.825 ;
        RECT 43.050 146.105 43.380 146.615 ;
        RECT 38.095 145.635 38.325 145.685 ;
        RECT 37.175 145.045 37.925 145.565 ;
        RECT 30.280 144.275 35.625 144.820 ;
        RECT 35.795 144.275 36.085 145.000 ;
        RECT 36.255 144.275 37.925 145.045 ;
        RECT 38.095 145.075 38.270 145.635 ;
        RECT 38.965 145.435 39.135 145.685 ;
        RECT 38.440 145.265 39.135 145.435 ;
        RECT 39.310 145.265 39.730 145.465 ;
        RECT 39.900 145.265 40.230 145.465 ;
        RECT 40.400 145.265 40.730 145.465 ;
        RECT 38.095 144.445 38.435 145.075 ;
        RECT 38.605 144.275 38.855 145.075 ;
        RECT 39.045 144.925 40.270 145.095 ;
        RECT 39.045 144.445 39.375 144.925 ;
        RECT 39.545 144.275 39.770 144.735 ;
        RECT 39.940 144.445 40.270 144.925 ;
        RECT 40.900 145.055 41.070 145.685 ;
        RECT 41.255 145.265 41.605 145.515 ;
        RECT 40.900 144.445 41.400 145.055 ;
        RECT 42.150 144.985 42.330 145.845 ;
        RECT 43.050 145.515 43.300 146.105 ;
        RECT 43.650 145.955 43.820 146.565 ;
        RECT 43.990 146.135 44.320 146.825 ;
        RECT 44.550 146.275 44.790 146.565 ;
        RECT 44.990 146.445 45.410 146.825 ;
        RECT 45.590 146.355 46.220 146.605 ;
        RECT 46.690 146.445 47.020 146.825 ;
        RECT 45.590 146.275 45.760 146.355 ;
        RECT 47.190 146.275 47.360 146.565 ;
        RECT 47.540 146.445 47.920 146.825 ;
        RECT 48.160 146.440 48.990 146.610 ;
        RECT 44.550 146.105 45.760 146.275 ;
        RECT 42.500 145.185 43.300 145.515 ;
        RECT 42.150 144.785 42.405 144.985 ;
        RECT 42.065 144.615 42.405 144.785 ;
        RECT 42.150 144.455 42.405 144.615 ;
        RECT 42.585 144.275 42.870 144.735 ;
        RECT 43.050 144.535 43.300 145.185 ;
        RECT 43.500 145.935 43.820 145.955 ;
        RECT 43.500 145.765 45.420 145.935 ;
        RECT 43.500 144.870 43.690 145.765 ;
        RECT 45.590 145.595 45.760 146.105 ;
        RECT 45.930 145.845 46.450 146.155 ;
        RECT 43.860 145.425 45.760 145.595 ;
        RECT 43.860 145.365 44.190 145.425 ;
        RECT 44.340 145.195 44.670 145.255 ;
        RECT 44.010 144.925 44.670 145.195 ;
        RECT 43.500 144.540 43.820 144.870 ;
        RECT 44.000 144.275 44.660 144.755 ;
        RECT 44.860 144.665 45.030 145.425 ;
        RECT 45.930 145.255 46.110 145.665 ;
        RECT 45.200 145.085 45.530 145.205 ;
        RECT 46.280 145.085 46.450 145.845 ;
        RECT 45.200 144.915 46.450 145.085 ;
        RECT 46.620 146.025 47.990 146.275 ;
        RECT 46.620 145.255 46.810 146.025 ;
        RECT 47.740 145.765 47.990 146.025 ;
        RECT 46.980 145.595 47.230 145.755 ;
        RECT 48.160 145.595 48.330 146.440 ;
        RECT 49.225 146.155 49.395 146.655 ;
        RECT 49.565 146.325 49.895 146.825 ;
        RECT 48.500 145.765 49.000 146.145 ;
        RECT 49.225 145.985 49.920 146.155 ;
        RECT 46.980 145.425 48.330 145.595 ;
        RECT 47.910 145.385 48.330 145.425 ;
        RECT 46.620 144.915 47.040 145.255 ;
        RECT 47.330 144.925 47.740 145.255 ;
        RECT 44.860 144.495 45.710 144.665 ;
        RECT 46.270 144.275 46.590 144.735 ;
        RECT 46.790 144.485 47.040 144.915 ;
        RECT 47.330 144.275 47.740 144.715 ;
        RECT 47.910 144.655 48.080 145.385 ;
        RECT 48.250 144.835 48.600 145.205 ;
        RECT 48.780 144.895 49.000 145.765 ;
        RECT 49.170 145.195 49.580 145.815 ;
        RECT 49.750 145.015 49.920 145.985 ;
        RECT 49.225 144.825 49.920 145.015 ;
        RECT 47.910 144.455 48.925 144.655 ;
        RECT 49.225 144.495 49.395 144.825 ;
        RECT 49.565 144.275 49.895 144.655 ;
        RECT 50.110 144.535 50.335 146.655 ;
        RECT 50.505 146.325 50.835 146.825 ;
        RECT 51.005 146.155 51.175 146.655 ;
        RECT 50.510 145.985 51.175 146.155 ;
        RECT 50.510 144.995 50.740 145.985 ;
        RECT 50.910 145.165 51.260 145.815 ;
        RECT 51.435 145.750 51.705 146.655 ;
        RECT 51.875 146.065 52.205 146.825 ;
        RECT 52.385 145.895 52.555 146.655 ;
        RECT 50.510 144.825 51.175 144.995 ;
        RECT 50.505 144.275 50.835 144.655 ;
        RECT 51.005 144.535 51.175 144.825 ;
        RECT 51.435 144.950 51.605 145.750 ;
        RECT 51.890 145.725 52.555 145.895 ;
        RECT 53.735 145.735 57.245 146.825 ;
        RECT 57.415 146.065 57.930 146.475 ;
        RECT 58.165 146.065 58.335 146.825 ;
        RECT 58.505 146.485 60.535 146.655 ;
        RECT 51.890 145.580 52.060 145.725 ;
        RECT 51.775 145.250 52.060 145.580 ;
        RECT 51.890 144.995 52.060 145.250 ;
        RECT 52.295 145.175 52.625 145.545 ;
        RECT 53.735 145.215 55.425 145.735 ;
        RECT 55.595 145.045 57.245 145.565 ;
        RECT 57.415 145.255 57.755 146.065 ;
        RECT 58.505 145.820 58.675 146.485 ;
        RECT 59.070 146.145 60.195 146.315 ;
        RECT 57.925 145.630 58.675 145.820 ;
        RECT 58.845 145.805 59.855 145.975 ;
        RECT 57.415 145.085 58.645 145.255 ;
        RECT 51.435 144.445 51.695 144.950 ;
        RECT 51.890 144.825 52.555 144.995 ;
        RECT 51.875 144.275 52.205 144.655 ;
        RECT 52.385 144.445 52.555 144.825 ;
        RECT 53.735 144.275 57.245 145.045 ;
        RECT 57.690 144.480 57.935 145.085 ;
        RECT 58.155 144.275 58.665 144.810 ;
        RECT 58.845 144.445 59.035 145.805 ;
        RECT 59.205 144.785 59.480 145.605 ;
        RECT 59.685 145.005 59.855 145.805 ;
        RECT 60.025 145.015 60.195 146.145 ;
        RECT 60.365 145.515 60.535 146.485 ;
        RECT 60.705 145.685 60.875 146.825 ;
        RECT 61.045 145.685 61.380 146.655 ;
        RECT 60.365 145.185 60.560 145.515 ;
        RECT 60.785 145.185 61.040 145.515 ;
        RECT 60.785 145.015 60.955 145.185 ;
        RECT 61.210 145.015 61.380 145.685 ;
        RECT 61.555 145.660 61.845 146.825 ;
        RECT 62.055 145.685 62.285 146.825 ;
        RECT 62.455 145.675 62.785 146.655 ;
        RECT 62.955 145.685 63.165 146.825 ;
        RECT 64.405 145.895 64.575 146.655 ;
        RECT 64.790 146.065 65.120 146.825 ;
        RECT 64.405 145.725 65.120 145.895 ;
        RECT 65.290 145.750 65.545 146.655 ;
        RECT 62.035 145.265 62.365 145.515 ;
        RECT 60.025 144.845 60.955 145.015 ;
        RECT 60.025 144.810 60.200 144.845 ;
        RECT 59.205 144.615 59.485 144.785 ;
        RECT 59.205 144.445 59.480 144.615 ;
        RECT 59.670 144.445 60.200 144.810 ;
        RECT 60.625 144.275 60.955 144.675 ;
        RECT 61.125 144.445 61.380 145.015 ;
        RECT 61.555 144.275 61.845 145.000 ;
        RECT 62.055 144.275 62.285 145.095 ;
        RECT 62.535 145.075 62.785 145.675 ;
        RECT 64.315 145.175 64.670 145.545 ;
        RECT 64.950 145.515 65.120 145.725 ;
        RECT 64.950 145.185 65.205 145.515 ;
        RECT 62.455 144.445 62.785 145.075 ;
        RECT 62.955 144.275 63.165 145.095 ;
        RECT 64.950 144.995 65.120 145.185 ;
        RECT 65.375 145.020 65.545 145.750 ;
        RECT 65.720 145.675 65.980 146.825 ;
        RECT 66.245 145.895 66.415 146.655 ;
        RECT 66.595 146.065 66.925 146.825 ;
        RECT 66.245 145.725 66.910 145.895 ;
        RECT 67.095 145.750 67.365 146.655 ;
        RECT 66.740 145.580 66.910 145.725 ;
        RECT 66.175 145.175 66.505 145.545 ;
        RECT 66.740 145.250 67.025 145.580 ;
        RECT 64.405 144.825 65.120 144.995 ;
        RECT 64.405 144.445 64.575 144.825 ;
        RECT 64.790 144.275 65.120 144.655 ;
        RECT 65.290 144.445 65.545 145.020 ;
        RECT 65.720 144.275 65.980 145.115 ;
        RECT 66.740 144.995 66.910 145.250 ;
        RECT 66.245 144.825 66.910 144.995 ;
        RECT 67.195 144.950 67.365 145.750 ;
        RECT 67.535 145.735 69.205 146.825 ;
        RECT 67.535 145.215 68.285 145.735 ;
        RECT 69.375 145.685 69.645 146.655 ;
        RECT 69.855 146.025 70.135 146.825 ;
        RECT 70.305 146.315 71.960 146.605 ;
        RECT 70.370 145.975 71.960 146.145 ;
        RECT 70.370 145.855 70.540 145.975 ;
        RECT 69.815 145.685 70.540 145.855 ;
        RECT 68.455 145.045 69.205 145.565 ;
        RECT 66.245 144.445 66.415 144.825 ;
        RECT 66.595 144.275 66.925 144.655 ;
        RECT 67.105 144.445 67.365 144.950 ;
        RECT 67.535 144.275 69.205 145.045 ;
        RECT 69.375 144.950 69.545 145.685 ;
        RECT 69.815 145.515 69.985 145.685 ;
        RECT 69.715 145.185 69.985 145.515 ;
        RECT 70.155 145.185 70.560 145.515 ;
        RECT 70.730 145.185 71.440 145.805 ;
        RECT 71.640 145.685 71.960 145.975 ;
        RECT 72.135 145.735 73.805 146.825 ;
        RECT 74.350 146.485 74.605 146.515 ;
        RECT 74.265 146.315 74.605 146.485 ;
        RECT 74.350 145.845 74.605 146.315 ;
        RECT 74.785 146.025 75.070 146.825 ;
        RECT 75.250 146.105 75.580 146.615 ;
        RECT 69.815 145.015 69.985 145.185 ;
        RECT 69.375 144.605 69.645 144.950 ;
        RECT 69.815 144.845 71.425 145.015 ;
        RECT 71.610 144.945 71.960 145.515 ;
        RECT 72.135 145.215 72.885 145.735 ;
        RECT 73.055 145.045 73.805 145.565 ;
        RECT 69.835 144.275 70.215 144.675 ;
        RECT 70.385 144.495 70.555 144.845 ;
        RECT 70.725 144.275 71.055 144.675 ;
        RECT 71.255 144.495 71.425 144.845 ;
        RECT 71.625 144.275 71.955 144.775 ;
        RECT 72.135 144.275 73.805 145.045 ;
        RECT 74.350 144.985 74.530 145.845 ;
        RECT 75.250 145.515 75.500 146.105 ;
        RECT 75.850 145.955 76.020 146.565 ;
        RECT 76.190 146.135 76.520 146.825 ;
        RECT 76.750 146.275 76.990 146.565 ;
        RECT 77.190 146.445 77.610 146.825 ;
        RECT 77.790 146.355 78.420 146.605 ;
        RECT 78.890 146.445 79.220 146.825 ;
        RECT 77.790 146.275 77.960 146.355 ;
        RECT 79.390 146.275 79.560 146.565 ;
        RECT 79.740 146.445 80.120 146.825 ;
        RECT 80.360 146.440 81.190 146.610 ;
        RECT 76.750 146.105 77.960 146.275 ;
        RECT 74.700 145.185 75.500 145.515 ;
        RECT 74.350 144.455 74.605 144.985 ;
        RECT 74.785 144.275 75.070 144.735 ;
        RECT 75.250 144.535 75.500 145.185 ;
        RECT 75.700 145.935 76.020 145.955 ;
        RECT 75.700 145.765 77.620 145.935 ;
        RECT 75.700 144.870 75.890 145.765 ;
        RECT 77.790 145.595 77.960 146.105 ;
        RECT 78.130 145.845 78.650 146.155 ;
        RECT 76.060 145.425 77.960 145.595 ;
        RECT 76.060 145.365 76.390 145.425 ;
        RECT 76.540 145.195 76.870 145.255 ;
        RECT 76.210 144.925 76.870 145.195 ;
        RECT 75.700 144.540 76.020 144.870 ;
        RECT 76.200 144.275 76.860 144.755 ;
        RECT 77.060 144.665 77.230 145.425 ;
        RECT 78.130 145.255 78.310 145.665 ;
        RECT 77.400 145.085 77.730 145.205 ;
        RECT 78.480 145.085 78.650 145.845 ;
        RECT 77.400 144.915 78.650 145.085 ;
        RECT 78.820 146.025 80.190 146.275 ;
        RECT 78.820 145.255 79.010 146.025 ;
        RECT 79.940 145.765 80.190 146.025 ;
        RECT 79.180 145.595 79.430 145.755 ;
        RECT 80.360 145.595 80.530 146.440 ;
        RECT 81.425 146.155 81.595 146.655 ;
        RECT 81.765 146.325 82.095 146.825 ;
        RECT 80.700 145.765 81.200 146.145 ;
        RECT 81.425 145.985 82.120 146.155 ;
        RECT 79.180 145.425 80.530 145.595 ;
        RECT 80.110 145.385 80.530 145.425 ;
        RECT 78.820 144.915 79.240 145.255 ;
        RECT 79.530 144.925 79.940 145.255 ;
        RECT 77.060 144.495 77.910 144.665 ;
        RECT 78.470 144.275 78.790 144.735 ;
        RECT 78.990 144.485 79.240 144.915 ;
        RECT 79.530 144.275 79.940 144.715 ;
        RECT 80.110 144.655 80.280 145.385 ;
        RECT 80.450 144.835 80.800 145.205 ;
        RECT 80.980 144.895 81.200 145.765 ;
        RECT 81.370 145.195 81.780 145.815 ;
        RECT 81.950 145.015 82.120 145.985 ;
        RECT 81.425 144.825 82.120 145.015 ;
        RECT 80.110 144.455 81.125 144.655 ;
        RECT 81.425 144.495 81.595 144.825 ;
        RECT 81.765 144.275 82.095 144.655 ;
        RECT 82.310 144.535 82.535 146.655 ;
        RECT 82.705 146.325 83.035 146.825 ;
        RECT 83.205 146.155 83.375 146.655 ;
        RECT 82.710 145.985 83.375 146.155 ;
        RECT 82.710 144.995 82.940 145.985 ;
        RECT 83.110 145.165 83.460 145.815 ;
        RECT 83.635 145.735 87.145 146.825 ;
        RECT 83.635 145.215 85.325 145.735 ;
        RECT 87.315 145.660 87.605 146.825 ;
        RECT 87.775 145.685 88.045 146.655 ;
        RECT 88.255 146.025 88.535 146.825 ;
        RECT 88.705 146.315 90.360 146.605 ;
        RECT 88.770 145.975 90.360 146.145 ;
        RECT 88.770 145.855 88.940 145.975 ;
        RECT 88.215 145.685 88.940 145.855 ;
        RECT 85.495 145.045 87.145 145.565 ;
        RECT 82.710 144.825 83.375 144.995 ;
        RECT 82.705 144.275 83.035 144.655 ;
        RECT 83.205 144.535 83.375 144.825 ;
        RECT 83.635 144.275 87.145 145.045 ;
        RECT 87.315 144.275 87.605 145.000 ;
        RECT 87.775 144.950 87.945 145.685 ;
        RECT 88.215 145.515 88.385 145.685 ;
        RECT 89.130 145.635 89.845 145.805 ;
        RECT 90.040 145.685 90.360 145.975 ;
        RECT 90.535 145.735 91.745 146.825 ;
        RECT 91.920 146.390 97.265 146.825 ;
        RECT 88.115 145.185 88.385 145.515 ;
        RECT 88.555 145.185 88.960 145.515 ;
        RECT 89.130 145.185 89.840 145.635 ;
        RECT 88.215 145.015 88.385 145.185 ;
        RECT 87.775 144.605 88.045 144.950 ;
        RECT 88.215 144.845 89.825 145.015 ;
        RECT 90.010 144.945 90.360 145.515 ;
        RECT 90.535 145.195 91.055 145.735 ;
        RECT 91.225 145.025 91.745 145.565 ;
        RECT 93.510 145.140 93.860 146.390 ;
        RECT 97.435 145.685 97.775 146.655 ;
        RECT 97.945 145.685 98.115 146.825 ;
        RECT 98.385 146.025 98.635 146.825 ;
        RECT 99.280 145.855 99.610 146.655 ;
        RECT 99.910 146.025 100.240 146.825 ;
        RECT 100.410 145.855 100.740 146.655 ;
        RECT 98.305 145.685 100.740 145.855 ;
        RECT 101.115 145.735 102.785 146.825 ;
        RECT 102.955 146.065 103.470 146.475 ;
        RECT 103.705 146.065 103.875 146.825 ;
        RECT 104.045 146.485 106.075 146.655 ;
        RECT 88.235 144.275 88.615 144.675 ;
        RECT 88.785 144.495 88.955 144.845 ;
        RECT 89.125 144.275 89.455 144.675 ;
        RECT 89.655 144.495 89.825 144.845 ;
        RECT 90.025 144.275 90.355 144.775 ;
        RECT 90.535 144.275 91.745 145.025 ;
        RECT 95.340 144.820 95.680 145.650 ;
        RECT 97.435 145.075 97.610 145.685 ;
        RECT 98.305 145.435 98.475 145.685 ;
        RECT 97.780 145.265 98.475 145.435 ;
        RECT 98.650 145.265 99.070 145.465 ;
        RECT 99.240 145.265 99.570 145.465 ;
        RECT 99.740 145.265 100.070 145.465 ;
        RECT 91.920 144.275 97.265 144.820 ;
        RECT 97.435 144.445 97.775 145.075 ;
        RECT 97.945 144.275 98.195 145.075 ;
        RECT 98.385 144.925 99.610 145.095 ;
        RECT 98.385 144.445 98.715 144.925 ;
        RECT 98.885 144.275 99.110 144.735 ;
        RECT 99.280 144.445 99.610 144.925 ;
        RECT 100.240 145.055 100.410 145.685 ;
        RECT 100.595 145.265 100.945 145.515 ;
        RECT 101.115 145.215 101.865 145.735 ;
        RECT 100.240 144.445 100.740 145.055 ;
        RECT 102.035 145.045 102.785 145.565 ;
        RECT 102.955 145.255 103.295 146.065 ;
        RECT 104.045 145.820 104.215 146.485 ;
        RECT 104.610 146.145 105.735 146.315 ;
        RECT 103.465 145.630 104.215 145.820 ;
        RECT 104.385 145.805 105.395 145.975 ;
        RECT 102.955 145.085 104.185 145.255 ;
        RECT 101.115 144.275 102.785 145.045 ;
        RECT 103.230 144.480 103.475 145.085 ;
        RECT 103.695 144.275 104.205 144.810 ;
        RECT 104.385 144.445 104.575 145.805 ;
        RECT 104.745 145.465 105.020 145.605 ;
        RECT 104.745 145.295 105.025 145.465 ;
        RECT 104.745 144.445 105.020 145.295 ;
        RECT 105.225 145.005 105.395 145.805 ;
        RECT 105.565 145.015 105.735 146.145 ;
        RECT 105.905 145.515 106.075 146.485 ;
        RECT 106.245 145.685 106.415 146.825 ;
        RECT 106.585 145.685 106.920 146.655 ;
        RECT 107.155 145.685 107.365 146.825 ;
        RECT 105.905 145.185 106.100 145.515 ;
        RECT 106.325 145.185 106.580 145.515 ;
        RECT 106.325 145.015 106.495 145.185 ;
        RECT 106.750 145.015 106.920 145.685 ;
        RECT 107.535 145.675 107.865 146.655 ;
        RECT 108.035 145.685 108.265 146.825 ;
        RECT 108.475 145.735 111.985 146.825 ;
        RECT 112.155 145.735 113.365 146.825 ;
        RECT 105.565 144.845 106.495 145.015 ;
        RECT 105.565 144.810 105.740 144.845 ;
        RECT 105.210 144.445 105.740 144.810 ;
        RECT 106.165 144.275 106.495 144.675 ;
        RECT 106.665 144.445 106.920 145.015 ;
        RECT 107.155 144.275 107.365 145.095 ;
        RECT 107.535 145.075 107.785 145.675 ;
        RECT 107.955 145.265 108.285 145.515 ;
        RECT 108.475 145.215 110.165 145.735 ;
        RECT 107.535 144.445 107.865 145.075 ;
        RECT 108.035 144.275 108.265 145.095 ;
        RECT 110.335 145.045 111.985 145.565 ;
        RECT 112.155 145.195 112.675 145.735 ;
        RECT 108.475 144.275 111.985 145.045 ;
        RECT 112.845 145.025 113.365 145.565 ;
        RECT 112.155 144.275 113.365 145.025 ;
        RECT 15.010 144.105 113.450 144.275 ;
        RECT 15.095 143.355 16.305 144.105 ;
        RECT 17.400 143.560 22.745 144.105 ;
        RECT 15.095 142.815 15.615 143.355 ;
        RECT 15.785 142.645 16.305 143.185 ;
        RECT 15.095 141.555 16.305 142.645 ;
        RECT 18.990 141.990 19.340 143.240 ;
        RECT 20.820 142.730 21.160 143.560 ;
        RECT 22.915 143.380 23.205 144.105 ;
        RECT 23.415 143.285 23.645 144.105 ;
        RECT 23.815 143.305 24.145 143.935 ;
        RECT 23.395 142.865 23.725 143.115 ;
        RECT 17.400 141.555 22.745 141.990 ;
        RECT 22.915 141.555 23.205 142.720 ;
        RECT 23.895 142.705 24.145 143.305 ;
        RECT 24.315 143.285 24.525 144.105 ;
        RECT 24.760 143.560 30.105 144.105 ;
        RECT 23.415 141.555 23.645 142.695 ;
        RECT 23.815 141.725 24.145 142.705 ;
        RECT 24.315 141.555 24.525 142.695 ;
        RECT 26.350 141.990 26.700 143.240 ;
        RECT 28.180 142.730 28.520 143.560 ;
        RECT 30.275 143.430 30.545 143.775 ;
        RECT 30.735 143.705 31.115 144.105 ;
        RECT 31.285 143.535 31.455 143.885 ;
        RECT 31.625 143.705 31.955 144.105 ;
        RECT 32.155 143.535 32.325 143.885 ;
        RECT 32.525 143.605 32.855 144.105 ;
        RECT 30.275 142.695 30.445 143.430 ;
        RECT 30.715 143.365 32.325 143.535 ;
        RECT 30.715 143.195 30.885 143.365 ;
        RECT 30.615 142.865 30.885 143.195 ;
        RECT 31.055 142.865 31.460 143.195 ;
        RECT 30.715 142.695 30.885 142.865 ;
        RECT 24.760 141.555 30.105 141.990 ;
        RECT 30.275 141.725 30.545 142.695 ;
        RECT 30.715 142.525 31.440 142.695 ;
        RECT 31.630 142.575 32.340 143.195 ;
        RECT 32.510 142.865 32.860 143.435 ;
        RECT 33.035 143.430 33.305 143.775 ;
        RECT 33.495 143.705 33.875 144.105 ;
        RECT 34.045 143.535 34.215 143.885 ;
        RECT 34.385 143.705 34.715 144.105 ;
        RECT 34.915 143.535 35.085 143.885 ;
        RECT 35.285 143.605 35.615 144.105 ;
        RECT 33.035 142.695 33.205 143.430 ;
        RECT 33.475 143.365 35.085 143.535 ;
        RECT 33.475 143.195 33.645 143.365 ;
        RECT 33.375 142.865 33.645 143.195 ;
        RECT 33.815 142.865 34.220 143.195 ;
        RECT 33.475 142.695 33.645 142.865 ;
        RECT 31.270 142.405 31.440 142.525 ;
        RECT 32.540 142.405 32.860 142.695 ;
        RECT 30.755 141.555 31.035 142.355 ;
        RECT 31.270 142.235 32.860 142.405 ;
        RECT 31.205 141.775 32.860 142.065 ;
        RECT 33.035 141.725 33.305 142.695 ;
        RECT 33.475 142.525 34.200 142.695 ;
        RECT 34.390 142.575 35.100 143.195 ;
        RECT 35.270 142.865 35.620 143.435 ;
        RECT 36.255 143.335 38.845 144.105 ;
        RECT 34.030 142.405 34.200 142.525 ;
        RECT 35.300 142.405 35.620 142.695 ;
        RECT 33.515 141.555 33.795 142.355 ;
        RECT 34.030 142.235 35.620 142.405 ;
        RECT 36.255 142.645 37.465 143.165 ;
        RECT 37.635 142.815 38.845 143.335 ;
        RECT 39.055 143.285 39.285 144.105 ;
        RECT 39.455 143.305 39.785 143.935 ;
        RECT 39.035 142.865 39.365 143.115 ;
        RECT 39.535 142.705 39.785 143.305 ;
        RECT 39.955 143.285 40.165 144.105 ;
        RECT 40.395 143.335 42.065 144.105 ;
        RECT 33.965 141.775 35.620 142.065 ;
        RECT 36.255 141.555 38.845 142.645 ;
        RECT 39.055 141.555 39.285 142.695 ;
        RECT 39.455 141.725 39.785 142.705 ;
        RECT 39.955 141.555 40.165 142.695 ;
        RECT 40.395 142.645 41.145 143.165 ;
        RECT 41.315 142.815 42.065 143.335 ;
        RECT 42.275 143.285 42.505 144.105 ;
        RECT 42.675 143.305 43.005 143.935 ;
        RECT 42.255 142.865 42.585 143.115 ;
        RECT 42.755 142.705 43.005 143.305 ;
        RECT 43.175 143.285 43.385 144.105 ;
        RECT 43.890 143.295 44.135 143.900 ;
        RECT 44.355 143.570 44.865 144.105 ;
        RECT 40.395 141.555 42.065 142.645 ;
        RECT 42.275 141.555 42.505 142.695 ;
        RECT 42.675 141.725 43.005 142.705 ;
        RECT 43.615 143.125 44.845 143.295 ;
        RECT 43.175 141.555 43.385 142.695 ;
        RECT 43.615 142.315 43.955 143.125 ;
        RECT 44.125 142.560 44.875 142.750 ;
        RECT 43.615 141.905 44.130 142.315 ;
        RECT 44.365 141.555 44.535 142.315 ;
        RECT 44.705 141.895 44.875 142.560 ;
        RECT 45.045 142.575 45.235 143.935 ;
        RECT 45.405 143.765 45.680 143.935 ;
        RECT 45.405 143.595 45.685 143.765 ;
        RECT 45.405 142.775 45.680 143.595 ;
        RECT 45.870 143.570 46.400 143.935 ;
        RECT 46.825 143.705 47.155 144.105 ;
        RECT 46.225 143.535 46.400 143.570 ;
        RECT 45.885 142.575 46.055 143.375 ;
        RECT 45.045 142.405 46.055 142.575 ;
        RECT 46.225 143.365 47.155 143.535 ;
        RECT 47.325 143.365 47.580 143.935 ;
        RECT 48.675 143.380 48.965 144.105 ;
        RECT 49.145 143.605 49.475 144.105 ;
        RECT 49.675 143.535 49.845 143.885 ;
        RECT 50.045 143.705 50.375 144.105 ;
        RECT 50.545 143.535 50.715 143.885 ;
        RECT 50.885 143.705 51.265 144.105 ;
        RECT 46.225 142.235 46.395 143.365 ;
        RECT 46.985 143.195 47.155 143.365 ;
        RECT 45.270 142.065 46.395 142.235 ;
        RECT 46.565 142.865 46.760 143.195 ;
        RECT 46.985 142.865 47.240 143.195 ;
        RECT 46.565 141.895 46.735 142.865 ;
        RECT 47.410 142.695 47.580 143.365 ;
        RECT 49.140 142.865 49.490 143.435 ;
        RECT 49.675 143.365 51.285 143.535 ;
        RECT 51.455 143.430 51.725 143.775 ;
        RECT 51.115 143.195 51.285 143.365 ;
        RECT 44.705 141.725 46.735 141.895 ;
        RECT 46.905 141.555 47.075 142.695 ;
        RECT 47.245 141.725 47.580 142.695 ;
        RECT 48.675 141.555 48.965 142.720 ;
        RECT 49.140 142.405 49.460 142.695 ;
        RECT 49.660 142.575 50.370 143.195 ;
        RECT 50.540 142.865 50.945 143.195 ;
        RECT 51.115 142.865 51.385 143.195 ;
        RECT 51.115 142.695 51.285 142.865 ;
        RECT 51.555 142.695 51.725 143.430 ;
        RECT 50.560 142.525 51.285 142.695 ;
        RECT 50.560 142.405 50.730 142.525 ;
        RECT 49.140 142.235 50.730 142.405 ;
        RECT 49.140 141.775 50.795 142.065 ;
        RECT 50.965 141.555 51.245 142.355 ;
        RECT 51.455 141.725 51.725 142.695 ;
        RECT 51.895 143.305 52.235 143.935 ;
        RECT 52.405 143.305 52.655 144.105 ;
        RECT 52.845 143.455 53.175 143.935 ;
        RECT 53.345 143.645 53.570 144.105 ;
        RECT 53.740 143.455 54.070 143.935 ;
        RECT 51.895 142.695 52.070 143.305 ;
        RECT 52.845 143.285 54.070 143.455 ;
        RECT 54.700 143.325 55.200 143.935 ;
        RECT 52.240 142.945 52.935 143.115 ;
        RECT 52.765 142.695 52.935 142.945 ;
        RECT 53.110 142.915 53.530 143.115 ;
        RECT 53.700 142.915 54.030 143.115 ;
        RECT 54.200 142.915 54.530 143.115 ;
        RECT 54.700 142.695 54.870 143.325 ;
        RECT 55.575 143.305 55.915 143.935 ;
        RECT 56.085 143.305 56.335 144.105 ;
        RECT 56.525 143.455 56.855 143.935 ;
        RECT 57.025 143.645 57.250 144.105 ;
        RECT 57.420 143.455 57.750 143.935 ;
        RECT 55.055 142.865 55.405 143.115 ;
        RECT 55.575 142.695 55.750 143.305 ;
        RECT 56.525 143.285 57.750 143.455 ;
        RECT 58.380 143.325 58.880 143.935 ;
        RECT 59.630 143.395 59.885 143.925 ;
        RECT 60.065 143.645 60.350 144.105 ;
        RECT 55.920 142.945 56.615 143.115 ;
        RECT 56.445 142.695 56.615 142.945 ;
        RECT 56.790 142.915 57.210 143.115 ;
        RECT 57.380 142.915 57.710 143.115 ;
        RECT 57.880 142.915 58.210 143.115 ;
        RECT 58.380 142.695 58.550 143.325 ;
        RECT 58.735 142.865 59.085 143.115 ;
        RECT 51.895 141.725 52.235 142.695 ;
        RECT 52.405 141.555 52.575 142.695 ;
        RECT 52.765 142.525 55.200 142.695 ;
        RECT 52.845 141.555 53.095 142.355 ;
        RECT 53.740 141.725 54.070 142.525 ;
        RECT 54.370 141.555 54.700 142.355 ;
        RECT 54.870 141.725 55.200 142.525 ;
        RECT 55.575 141.725 55.915 142.695 ;
        RECT 56.085 141.555 56.255 142.695 ;
        RECT 56.445 142.525 58.880 142.695 ;
        RECT 56.525 141.555 56.775 142.355 ;
        RECT 57.420 141.725 57.750 142.525 ;
        RECT 58.050 141.555 58.380 142.355 ;
        RECT 58.550 141.725 58.880 142.525 ;
        RECT 59.630 142.535 59.810 143.395 ;
        RECT 60.530 143.195 60.780 143.845 ;
        RECT 59.980 142.865 60.780 143.195 ;
        RECT 59.630 142.065 59.885 142.535 ;
        RECT 59.545 141.895 59.885 142.065 ;
        RECT 59.630 141.865 59.885 141.895 ;
        RECT 60.065 141.555 60.350 142.355 ;
        RECT 60.530 142.275 60.780 142.865 ;
        RECT 60.980 143.510 61.300 143.840 ;
        RECT 61.480 143.625 62.140 144.105 ;
        RECT 62.340 143.715 63.190 143.885 ;
        RECT 60.980 142.615 61.170 143.510 ;
        RECT 61.490 143.185 62.150 143.455 ;
        RECT 61.820 143.125 62.150 143.185 ;
        RECT 61.340 142.955 61.670 143.015 ;
        RECT 62.340 142.955 62.510 143.715 ;
        RECT 63.750 143.645 64.070 144.105 ;
        RECT 64.270 143.465 64.520 143.895 ;
        RECT 64.810 143.665 65.220 144.105 ;
        RECT 65.390 143.725 66.405 143.925 ;
        RECT 62.680 143.295 63.930 143.465 ;
        RECT 62.680 143.175 63.010 143.295 ;
        RECT 61.340 142.785 63.240 142.955 ;
        RECT 60.980 142.445 62.900 142.615 ;
        RECT 60.980 142.425 61.300 142.445 ;
        RECT 60.530 141.765 60.860 142.275 ;
        RECT 61.130 141.815 61.300 142.425 ;
        RECT 63.070 142.275 63.240 142.785 ;
        RECT 63.410 142.715 63.590 143.125 ;
        RECT 63.760 142.535 63.930 143.295 ;
        RECT 61.470 141.555 61.800 142.245 ;
        RECT 62.030 142.105 63.240 142.275 ;
        RECT 63.410 142.225 63.930 142.535 ;
        RECT 64.100 143.125 64.520 143.465 ;
        RECT 64.810 143.125 65.220 143.455 ;
        RECT 64.100 142.355 64.290 143.125 ;
        RECT 65.390 142.995 65.560 143.725 ;
        RECT 66.705 143.555 66.875 143.885 ;
        RECT 67.045 143.725 67.375 144.105 ;
        RECT 65.730 143.175 66.080 143.545 ;
        RECT 65.390 142.955 65.810 142.995 ;
        RECT 64.460 142.785 65.810 142.955 ;
        RECT 64.460 142.625 64.710 142.785 ;
        RECT 65.220 142.355 65.470 142.615 ;
        RECT 64.100 142.105 65.470 142.355 ;
        RECT 62.030 141.815 62.270 142.105 ;
        RECT 63.070 142.025 63.240 142.105 ;
        RECT 62.470 141.555 62.890 141.935 ;
        RECT 63.070 141.775 63.700 142.025 ;
        RECT 64.170 141.555 64.500 141.935 ;
        RECT 64.670 141.815 64.840 142.105 ;
        RECT 65.640 141.940 65.810 142.785 ;
        RECT 66.260 142.615 66.480 143.485 ;
        RECT 66.705 143.365 67.400 143.555 ;
        RECT 65.980 142.235 66.480 142.615 ;
        RECT 66.650 142.565 67.060 143.185 ;
        RECT 67.230 142.395 67.400 143.365 ;
        RECT 66.705 142.225 67.400 142.395 ;
        RECT 65.020 141.555 65.400 141.935 ;
        RECT 65.640 141.770 66.470 141.940 ;
        RECT 66.705 141.725 66.875 142.225 ;
        RECT 67.045 141.555 67.375 142.055 ;
        RECT 67.590 141.725 67.815 143.845 ;
        RECT 67.985 143.725 68.315 144.105 ;
        RECT 68.485 143.555 68.655 143.845 ;
        RECT 68.920 143.560 74.265 144.105 ;
        RECT 67.990 143.385 68.655 143.555 ;
        RECT 67.990 142.395 68.220 143.385 ;
        RECT 68.390 142.565 68.740 143.215 ;
        RECT 67.990 142.225 68.655 142.395 ;
        RECT 67.985 141.555 68.315 142.055 ;
        RECT 68.485 141.725 68.655 142.225 ;
        RECT 70.510 141.990 70.860 143.240 ;
        RECT 72.340 142.730 72.680 143.560 ;
        RECT 74.435 143.380 74.725 144.105 ;
        RECT 75.815 143.335 79.325 144.105 ;
        RECT 79.585 143.555 79.755 143.935 ;
        RECT 79.935 143.725 80.265 144.105 ;
        RECT 79.585 143.385 80.250 143.555 ;
        RECT 80.445 143.430 80.705 143.935 ;
        RECT 68.920 141.555 74.265 141.990 ;
        RECT 74.435 141.555 74.725 142.720 ;
        RECT 75.815 142.645 77.505 143.165 ;
        RECT 77.675 142.815 79.325 143.335 ;
        RECT 79.515 142.835 79.845 143.205 ;
        RECT 80.080 143.130 80.250 143.385 ;
        RECT 80.080 142.800 80.365 143.130 ;
        RECT 80.080 142.655 80.250 142.800 ;
        RECT 75.815 141.555 79.325 142.645 ;
        RECT 79.585 142.485 80.250 142.655 ;
        RECT 80.535 142.630 80.705 143.430 ;
        RECT 80.875 143.335 83.465 144.105 ;
        RECT 79.585 141.725 79.755 142.485 ;
        RECT 79.935 141.555 80.265 142.315 ;
        RECT 80.435 141.725 80.705 142.630 ;
        RECT 80.875 142.645 82.085 143.165 ;
        RECT 82.255 142.815 83.465 143.335 ;
        RECT 83.910 143.295 84.155 143.900 ;
        RECT 84.375 143.570 84.885 144.105 ;
        RECT 83.635 143.125 84.865 143.295 ;
        RECT 80.875 141.555 83.465 142.645 ;
        RECT 83.635 142.315 83.975 143.125 ;
        RECT 84.145 142.560 84.895 142.750 ;
        RECT 83.635 141.905 84.150 142.315 ;
        RECT 84.385 141.555 84.555 142.315 ;
        RECT 84.725 141.895 84.895 142.560 ;
        RECT 85.065 142.575 85.255 143.935 ;
        RECT 85.425 143.425 85.700 143.935 ;
        RECT 85.890 143.570 86.420 143.935 ;
        RECT 86.845 143.705 87.175 144.105 ;
        RECT 86.245 143.535 86.420 143.570 ;
        RECT 85.425 143.255 85.705 143.425 ;
        RECT 85.425 142.775 85.700 143.255 ;
        RECT 85.905 142.575 86.075 143.375 ;
        RECT 85.065 142.405 86.075 142.575 ;
        RECT 86.245 143.365 87.175 143.535 ;
        RECT 87.345 143.365 87.600 143.935 ;
        RECT 86.245 142.235 86.415 143.365 ;
        RECT 87.005 143.195 87.175 143.365 ;
        RECT 85.290 142.065 86.415 142.235 ;
        RECT 86.585 142.865 86.780 143.195 ;
        RECT 87.005 142.865 87.260 143.195 ;
        RECT 86.585 141.895 86.755 142.865 ;
        RECT 87.430 142.695 87.600 143.365 ;
        RECT 88.440 143.325 88.940 143.935 ;
        RECT 88.235 142.865 88.585 143.115 ;
        RECT 88.770 142.695 88.940 143.325 ;
        RECT 89.570 143.455 89.900 143.935 ;
        RECT 90.070 143.645 90.295 144.105 ;
        RECT 90.465 143.455 90.795 143.935 ;
        RECT 89.570 143.285 90.795 143.455 ;
        RECT 90.985 143.305 91.235 144.105 ;
        RECT 91.405 143.305 91.745 143.935 ;
        RECT 89.110 142.915 89.440 143.115 ;
        RECT 89.610 142.915 89.940 143.115 ;
        RECT 90.110 142.915 90.530 143.115 ;
        RECT 90.705 142.945 91.400 143.115 ;
        RECT 90.705 142.695 90.875 142.945 ;
        RECT 91.570 142.695 91.745 143.305 ;
        RECT 92.190 143.295 92.435 143.900 ;
        RECT 92.655 143.570 93.165 144.105 ;
        RECT 84.725 141.725 86.755 141.895 ;
        RECT 86.925 141.555 87.095 142.695 ;
        RECT 87.265 141.725 87.600 142.695 ;
        RECT 88.440 142.525 90.875 142.695 ;
        RECT 88.440 141.725 88.770 142.525 ;
        RECT 88.940 141.555 89.270 142.355 ;
        RECT 89.570 141.725 89.900 142.525 ;
        RECT 90.545 141.555 90.795 142.355 ;
        RECT 91.065 141.555 91.235 142.695 ;
        RECT 91.405 141.725 91.745 142.695 ;
        RECT 91.915 143.125 93.145 143.295 ;
        RECT 91.915 142.315 92.255 143.125 ;
        RECT 92.425 142.560 93.175 142.750 ;
        RECT 91.915 141.905 92.430 142.315 ;
        RECT 92.665 141.555 92.835 142.315 ;
        RECT 93.005 141.895 93.175 142.560 ;
        RECT 93.345 142.575 93.535 143.935 ;
        RECT 93.705 143.425 93.980 143.935 ;
        RECT 94.170 143.570 94.700 143.935 ;
        RECT 95.125 143.705 95.455 144.105 ;
        RECT 94.525 143.535 94.700 143.570 ;
        RECT 93.705 143.255 93.985 143.425 ;
        RECT 93.705 142.775 93.980 143.255 ;
        RECT 94.185 142.575 94.355 143.375 ;
        RECT 93.345 142.405 94.355 142.575 ;
        RECT 94.525 143.365 95.455 143.535 ;
        RECT 95.625 143.365 95.880 143.935 ;
        RECT 94.525 142.235 94.695 143.365 ;
        RECT 95.285 143.195 95.455 143.365 ;
        RECT 93.570 142.065 94.695 142.235 ;
        RECT 94.865 142.865 95.060 143.195 ;
        RECT 95.285 142.865 95.540 143.195 ;
        RECT 94.865 141.895 95.035 142.865 ;
        RECT 95.710 142.695 95.880 143.365 ;
        RECT 93.005 141.725 95.035 141.895 ;
        RECT 95.205 141.555 95.375 142.695 ;
        RECT 95.545 141.725 95.880 142.695 ;
        RECT 96.055 143.305 96.395 143.935 ;
        RECT 96.565 143.305 96.815 144.105 ;
        RECT 97.005 143.455 97.335 143.935 ;
        RECT 97.505 143.645 97.730 144.105 ;
        RECT 97.900 143.455 98.230 143.935 ;
        RECT 96.055 142.695 96.230 143.305 ;
        RECT 97.005 143.285 98.230 143.455 ;
        RECT 98.860 143.325 99.360 143.935 ;
        RECT 100.195 143.380 100.485 144.105 ;
        RECT 96.400 142.945 97.095 143.115 ;
        RECT 96.925 142.695 97.095 142.945 ;
        RECT 97.270 142.915 97.690 143.115 ;
        RECT 97.860 142.915 98.190 143.115 ;
        RECT 98.360 142.915 98.690 143.115 ;
        RECT 98.860 142.695 99.030 143.325 ;
        RECT 101.155 143.285 101.385 144.105 ;
        RECT 101.555 143.305 101.885 143.935 ;
        RECT 99.215 142.865 99.565 143.115 ;
        RECT 101.135 142.865 101.465 143.115 ;
        RECT 96.055 141.725 96.395 142.695 ;
        RECT 96.565 141.555 96.735 142.695 ;
        RECT 96.925 142.525 99.360 142.695 ;
        RECT 97.005 141.555 97.255 142.355 ;
        RECT 97.900 141.725 98.230 142.525 ;
        RECT 98.530 141.555 98.860 142.355 ;
        RECT 99.030 141.725 99.360 142.525 ;
        RECT 100.195 141.555 100.485 142.720 ;
        RECT 101.635 142.705 101.885 143.305 ;
        RECT 102.055 143.285 102.265 144.105 ;
        RECT 102.870 143.425 103.125 143.925 ;
        RECT 103.305 143.645 103.590 144.105 ;
        RECT 102.785 143.395 103.125 143.425 ;
        RECT 102.785 143.255 103.050 143.395 ;
        RECT 101.155 141.555 101.385 142.695 ;
        RECT 101.555 141.725 101.885 142.705 ;
        RECT 102.055 141.555 102.265 142.695 ;
        RECT 102.870 142.535 103.050 143.255 ;
        RECT 103.770 143.195 104.020 143.845 ;
        RECT 103.220 142.865 104.020 143.195 ;
        RECT 102.870 141.865 103.125 142.535 ;
        RECT 103.305 141.555 103.590 142.355 ;
        RECT 103.770 142.275 104.020 142.865 ;
        RECT 104.220 143.510 104.540 143.840 ;
        RECT 104.720 143.625 105.380 144.105 ;
        RECT 105.580 143.715 106.430 143.885 ;
        RECT 104.220 142.615 104.410 143.510 ;
        RECT 104.730 143.185 105.390 143.455 ;
        RECT 105.060 143.125 105.390 143.185 ;
        RECT 104.580 142.955 104.910 143.015 ;
        RECT 105.580 142.955 105.750 143.715 ;
        RECT 106.990 143.645 107.310 144.105 ;
        RECT 107.510 143.465 107.760 143.895 ;
        RECT 108.050 143.665 108.460 144.105 ;
        RECT 108.630 143.725 109.645 143.925 ;
        RECT 105.920 143.295 107.170 143.465 ;
        RECT 105.920 143.175 106.250 143.295 ;
        RECT 104.580 142.785 106.480 142.955 ;
        RECT 104.220 142.445 106.140 142.615 ;
        RECT 104.220 142.425 104.540 142.445 ;
        RECT 103.770 141.765 104.100 142.275 ;
        RECT 104.370 141.815 104.540 142.425 ;
        RECT 106.310 142.275 106.480 142.785 ;
        RECT 106.650 142.715 106.830 143.125 ;
        RECT 107.000 142.535 107.170 143.295 ;
        RECT 104.710 141.555 105.040 142.245 ;
        RECT 105.270 142.105 106.480 142.275 ;
        RECT 106.650 142.225 107.170 142.535 ;
        RECT 107.340 143.125 107.760 143.465 ;
        RECT 108.050 143.125 108.460 143.455 ;
        RECT 107.340 142.355 107.530 143.125 ;
        RECT 108.630 142.995 108.800 143.725 ;
        RECT 109.945 143.555 110.115 143.885 ;
        RECT 110.285 143.725 110.615 144.105 ;
        RECT 108.970 143.175 109.320 143.545 ;
        RECT 108.630 142.955 109.050 142.995 ;
        RECT 107.700 142.785 109.050 142.955 ;
        RECT 107.700 142.625 107.950 142.785 ;
        RECT 108.460 142.355 108.710 142.615 ;
        RECT 107.340 142.105 108.710 142.355 ;
        RECT 105.270 141.815 105.510 142.105 ;
        RECT 106.310 142.025 106.480 142.105 ;
        RECT 105.710 141.555 106.130 141.935 ;
        RECT 106.310 141.775 106.940 142.025 ;
        RECT 107.410 141.555 107.740 141.935 ;
        RECT 107.910 141.815 108.080 142.105 ;
        RECT 108.880 141.940 109.050 142.785 ;
        RECT 109.500 142.615 109.720 143.485 ;
        RECT 109.945 143.365 110.640 143.555 ;
        RECT 109.220 142.235 109.720 142.615 ;
        RECT 109.890 142.565 110.300 143.185 ;
        RECT 110.470 142.395 110.640 143.365 ;
        RECT 109.945 142.225 110.640 142.395 ;
        RECT 108.260 141.555 108.640 141.935 ;
        RECT 108.880 141.770 109.710 141.940 ;
        RECT 109.945 141.725 110.115 142.225 ;
        RECT 110.285 141.555 110.615 142.055 ;
        RECT 110.830 141.725 111.055 143.845 ;
        RECT 111.225 143.725 111.555 144.105 ;
        RECT 111.725 143.555 111.895 143.845 ;
        RECT 111.230 143.385 111.895 143.555 ;
        RECT 111.230 142.395 111.460 143.385 ;
        RECT 112.155 143.355 113.365 144.105 ;
        RECT 111.630 142.565 111.980 143.215 ;
        RECT 112.155 142.645 112.675 143.185 ;
        RECT 112.845 142.815 113.365 143.355 ;
        RECT 111.230 142.225 111.895 142.395 ;
        RECT 111.225 141.555 111.555 142.055 ;
        RECT 111.725 141.725 111.895 142.225 ;
        RECT 112.155 141.555 113.365 142.645 ;
        RECT 15.010 141.385 113.450 141.555 ;
        RECT 15.095 140.295 16.305 141.385 ;
        RECT 15.095 139.585 15.615 140.125 ;
        RECT 15.785 139.755 16.305 140.295 ;
        RECT 17.485 140.455 17.655 141.215 ;
        RECT 17.835 140.625 18.165 141.385 ;
        RECT 17.485 140.285 18.150 140.455 ;
        RECT 18.335 140.310 18.605 141.215 ;
        RECT 17.980 140.140 18.150 140.285 ;
        RECT 17.415 139.735 17.745 140.105 ;
        RECT 17.980 139.810 18.265 140.140 ;
        RECT 15.095 138.835 16.305 139.585 ;
        RECT 17.980 139.555 18.150 139.810 ;
        RECT 17.485 139.385 18.150 139.555 ;
        RECT 18.435 139.510 18.605 140.310 ;
        RECT 18.835 140.245 19.045 141.385 ;
        RECT 19.215 140.235 19.545 141.215 ;
        RECT 19.715 140.245 19.945 141.385 ;
        RECT 20.245 140.715 20.415 141.215 ;
        RECT 20.585 140.885 20.915 141.385 ;
        RECT 20.245 140.545 20.910 140.715 ;
        RECT 17.485 139.005 17.655 139.385 ;
        RECT 17.835 138.835 18.165 139.215 ;
        RECT 18.345 139.005 18.605 139.510 ;
        RECT 18.835 138.835 19.045 139.655 ;
        RECT 19.215 139.635 19.465 140.235 ;
        RECT 19.635 139.825 19.965 140.075 ;
        RECT 20.160 139.725 20.510 140.375 ;
        RECT 19.215 139.005 19.545 139.635 ;
        RECT 19.715 138.835 19.945 139.655 ;
        RECT 20.680 139.555 20.910 140.545 ;
        RECT 20.245 139.385 20.910 139.555 ;
        RECT 20.245 139.095 20.415 139.385 ;
        RECT 20.585 138.835 20.915 139.215 ;
        RECT 21.085 139.095 21.310 141.215 ;
        RECT 21.525 140.885 21.855 141.385 ;
        RECT 22.025 140.715 22.195 141.215 ;
        RECT 22.430 141.000 23.260 141.170 ;
        RECT 23.500 141.005 23.880 141.385 ;
        RECT 21.500 140.545 22.195 140.715 ;
        RECT 21.500 139.575 21.670 140.545 ;
        RECT 21.840 139.755 22.250 140.375 ;
        RECT 22.420 140.325 22.920 140.705 ;
        RECT 21.500 139.385 22.195 139.575 ;
        RECT 22.420 139.455 22.640 140.325 ;
        RECT 23.090 140.155 23.260 141.000 ;
        RECT 24.060 140.835 24.230 141.125 ;
        RECT 24.400 141.005 24.730 141.385 ;
        RECT 25.200 140.915 25.830 141.165 ;
        RECT 26.010 141.005 26.430 141.385 ;
        RECT 25.660 140.835 25.830 140.915 ;
        RECT 26.630 140.835 26.870 141.125 ;
        RECT 23.430 140.585 24.800 140.835 ;
        RECT 23.430 140.325 23.680 140.585 ;
        RECT 24.190 140.155 24.440 140.315 ;
        RECT 23.090 139.985 24.440 140.155 ;
        RECT 23.090 139.945 23.510 139.985 ;
        RECT 22.820 139.395 23.170 139.765 ;
        RECT 21.525 138.835 21.855 139.215 ;
        RECT 22.025 139.055 22.195 139.385 ;
        RECT 23.340 139.215 23.510 139.945 ;
        RECT 24.610 139.815 24.800 140.585 ;
        RECT 23.680 139.485 24.090 139.815 ;
        RECT 24.380 139.475 24.800 139.815 ;
        RECT 24.970 140.405 25.490 140.715 ;
        RECT 25.660 140.665 26.870 140.835 ;
        RECT 27.100 140.695 27.430 141.385 ;
        RECT 24.970 139.645 25.140 140.405 ;
        RECT 25.310 139.815 25.490 140.225 ;
        RECT 25.660 140.155 25.830 140.665 ;
        RECT 27.600 140.515 27.770 141.125 ;
        RECT 28.040 140.665 28.370 141.175 ;
        RECT 27.600 140.495 27.920 140.515 ;
        RECT 26.000 140.325 27.920 140.495 ;
        RECT 25.660 139.985 27.560 140.155 ;
        RECT 25.890 139.645 26.220 139.765 ;
        RECT 24.970 139.475 26.220 139.645 ;
        RECT 22.495 139.015 23.510 139.215 ;
        RECT 23.680 138.835 24.090 139.275 ;
        RECT 24.380 139.045 24.630 139.475 ;
        RECT 24.830 138.835 25.150 139.295 ;
        RECT 26.390 139.225 26.560 139.985 ;
        RECT 27.230 139.925 27.560 139.985 ;
        RECT 26.750 139.755 27.080 139.815 ;
        RECT 26.750 139.485 27.410 139.755 ;
        RECT 27.730 139.430 27.920 140.325 ;
        RECT 25.710 139.055 26.560 139.225 ;
        RECT 26.760 138.835 27.420 139.315 ;
        RECT 27.600 139.100 27.920 139.430 ;
        RECT 28.120 140.075 28.370 140.665 ;
        RECT 28.550 140.585 28.835 141.385 ;
        RECT 29.015 140.405 29.270 141.075 ;
        RECT 30.935 140.715 31.215 141.385 ;
        RECT 31.385 140.495 31.685 141.045 ;
        RECT 31.885 140.665 32.215 141.385 ;
        RECT 32.405 140.665 32.865 141.215 ;
        RECT 33.695 140.715 33.975 141.385 ;
        RECT 28.120 139.745 28.920 140.075 ;
        RECT 29.090 140.025 29.270 140.405 ;
        RECT 30.750 140.075 31.015 140.435 ;
        RECT 31.385 140.325 32.325 140.495 ;
        RECT 32.155 140.075 32.325 140.325 ;
        RECT 29.090 139.855 29.355 140.025 ;
        RECT 28.120 139.095 28.370 139.745 ;
        RECT 29.090 139.545 29.270 139.855 ;
        RECT 30.750 139.825 31.425 140.075 ;
        RECT 31.645 139.825 31.985 140.075 ;
        RECT 32.155 139.745 32.445 140.075 ;
        RECT 32.155 139.655 32.325 139.745 ;
        RECT 28.550 138.835 28.835 139.295 ;
        RECT 29.015 139.015 29.270 139.545 ;
        RECT 30.935 139.465 32.325 139.655 ;
        RECT 30.935 139.105 31.265 139.465 ;
        RECT 32.615 139.295 32.865 140.665 ;
        RECT 34.145 140.495 34.445 141.045 ;
        RECT 34.645 140.665 34.975 141.385 ;
        RECT 35.165 140.665 35.625 141.215 ;
        RECT 33.510 140.075 33.775 140.435 ;
        RECT 34.145 140.325 35.085 140.495 ;
        RECT 34.915 140.075 35.085 140.325 ;
        RECT 33.510 139.825 34.185 140.075 ;
        RECT 34.405 139.825 34.745 140.075 ;
        RECT 34.915 139.745 35.205 140.075 ;
        RECT 34.915 139.655 35.085 139.745 ;
        RECT 31.885 138.835 32.135 139.295 ;
        RECT 32.305 139.005 32.865 139.295 ;
        RECT 33.695 139.465 35.085 139.655 ;
        RECT 33.695 139.105 34.025 139.465 ;
        RECT 35.375 139.295 35.625 140.665 ;
        RECT 35.795 140.220 36.085 141.385 ;
        RECT 36.345 140.715 36.515 141.215 ;
        RECT 36.685 140.885 37.015 141.385 ;
        RECT 36.345 140.545 37.010 140.715 ;
        RECT 36.260 139.725 36.610 140.375 ;
        RECT 34.645 138.835 34.895 139.295 ;
        RECT 35.065 139.005 35.625 139.295 ;
        RECT 35.795 138.835 36.085 139.560 ;
        RECT 36.780 139.555 37.010 140.545 ;
        RECT 36.345 139.385 37.010 139.555 ;
        RECT 36.345 139.095 36.515 139.385 ;
        RECT 36.685 138.835 37.015 139.215 ;
        RECT 37.185 139.095 37.410 141.215 ;
        RECT 37.625 140.885 37.955 141.385 ;
        RECT 38.125 140.715 38.295 141.215 ;
        RECT 38.530 141.000 39.360 141.170 ;
        RECT 39.600 141.005 39.980 141.385 ;
        RECT 37.600 140.545 38.295 140.715 ;
        RECT 37.600 139.575 37.770 140.545 ;
        RECT 37.940 139.755 38.350 140.375 ;
        RECT 38.520 140.325 39.020 140.705 ;
        RECT 37.600 139.385 38.295 139.575 ;
        RECT 38.520 139.455 38.740 140.325 ;
        RECT 39.190 140.155 39.360 141.000 ;
        RECT 40.160 140.835 40.330 141.125 ;
        RECT 40.500 141.005 40.830 141.385 ;
        RECT 41.300 140.915 41.930 141.165 ;
        RECT 42.110 141.005 42.530 141.385 ;
        RECT 41.760 140.835 41.930 140.915 ;
        RECT 42.730 140.835 42.970 141.125 ;
        RECT 39.530 140.585 40.900 140.835 ;
        RECT 39.530 140.325 39.780 140.585 ;
        RECT 40.290 140.155 40.540 140.315 ;
        RECT 39.190 139.985 40.540 140.155 ;
        RECT 39.190 139.945 39.610 139.985 ;
        RECT 38.920 139.395 39.270 139.765 ;
        RECT 37.625 138.835 37.955 139.215 ;
        RECT 38.125 139.055 38.295 139.385 ;
        RECT 39.440 139.215 39.610 139.945 ;
        RECT 40.710 139.815 40.900 140.585 ;
        RECT 39.780 139.485 40.190 139.815 ;
        RECT 40.480 139.475 40.900 139.815 ;
        RECT 41.070 140.405 41.590 140.715 ;
        RECT 41.760 140.665 42.970 140.835 ;
        RECT 43.200 140.695 43.530 141.385 ;
        RECT 41.070 139.645 41.240 140.405 ;
        RECT 41.410 139.815 41.590 140.225 ;
        RECT 41.760 140.155 41.930 140.665 ;
        RECT 43.700 140.515 43.870 141.125 ;
        RECT 44.140 140.665 44.470 141.175 ;
        RECT 43.700 140.495 44.020 140.515 ;
        RECT 42.100 140.325 44.020 140.495 ;
        RECT 41.760 139.985 43.660 140.155 ;
        RECT 41.990 139.645 42.320 139.765 ;
        RECT 41.070 139.475 42.320 139.645 ;
        RECT 38.595 139.015 39.610 139.215 ;
        RECT 39.780 138.835 40.190 139.275 ;
        RECT 40.480 139.045 40.730 139.475 ;
        RECT 40.930 138.835 41.250 139.295 ;
        RECT 42.490 139.225 42.660 139.985 ;
        RECT 43.330 139.925 43.660 139.985 ;
        RECT 42.850 139.755 43.180 139.815 ;
        RECT 42.850 139.485 43.510 139.755 ;
        RECT 43.830 139.430 44.020 140.325 ;
        RECT 41.810 139.055 42.660 139.225 ;
        RECT 42.860 138.835 43.520 139.315 ;
        RECT 43.700 139.100 44.020 139.430 ;
        RECT 44.220 140.075 44.470 140.665 ;
        RECT 44.650 140.585 44.935 141.385 ;
        RECT 45.115 140.405 45.370 141.075 ;
        RECT 44.220 139.745 45.020 140.075 ;
        RECT 44.220 139.095 44.470 139.745 ;
        RECT 45.190 139.685 45.370 140.405 ;
        RECT 45.915 140.310 46.185 141.215 ;
        RECT 46.355 140.625 46.685 141.385 ;
        RECT 46.865 140.455 47.035 141.215 ;
        RECT 45.190 139.545 45.455 139.685 ;
        RECT 45.115 139.515 45.455 139.545 ;
        RECT 44.650 138.835 44.935 139.295 ;
        RECT 45.115 139.015 45.370 139.515 ;
        RECT 45.915 139.510 46.085 140.310 ;
        RECT 46.370 140.285 47.035 140.455 ;
        RECT 47.500 140.415 47.830 141.215 ;
        RECT 48.000 140.585 48.330 141.385 ;
        RECT 48.630 140.415 48.960 141.215 ;
        RECT 49.605 140.585 49.855 141.385 ;
        RECT 46.370 140.140 46.540 140.285 ;
        RECT 47.500 140.245 49.935 140.415 ;
        RECT 50.125 140.245 50.295 141.385 ;
        RECT 50.465 140.245 50.805 141.215 ;
        RECT 46.255 139.810 46.540 140.140 ;
        RECT 46.370 139.555 46.540 139.810 ;
        RECT 46.775 139.735 47.105 140.105 ;
        RECT 47.295 139.825 47.645 140.075 ;
        RECT 47.830 139.615 48.000 140.245 ;
        RECT 48.170 139.825 48.500 140.025 ;
        RECT 48.670 139.825 49.000 140.025 ;
        RECT 49.170 139.825 49.590 140.025 ;
        RECT 49.765 139.995 49.935 140.245 ;
        RECT 49.765 139.825 50.460 139.995 ;
        RECT 45.915 139.005 46.175 139.510 ;
        RECT 46.370 139.385 47.035 139.555 ;
        RECT 46.355 138.835 46.685 139.215 ;
        RECT 46.865 139.005 47.035 139.385 ;
        RECT 47.500 139.005 48.000 139.615 ;
        RECT 48.630 139.485 49.855 139.655 ;
        RECT 50.630 139.635 50.805 140.245 ;
        RECT 50.975 140.625 51.490 141.035 ;
        RECT 51.725 140.625 51.895 141.385 ;
        RECT 52.065 141.045 54.095 141.215 ;
        RECT 50.975 139.815 51.315 140.625 ;
        RECT 52.065 140.380 52.235 141.045 ;
        RECT 52.630 140.705 53.755 140.875 ;
        RECT 51.485 140.190 52.235 140.380 ;
        RECT 52.405 140.365 53.415 140.535 ;
        RECT 50.975 139.645 52.205 139.815 ;
        RECT 48.630 139.005 48.960 139.485 ;
        RECT 49.130 138.835 49.355 139.295 ;
        RECT 49.525 139.005 49.855 139.485 ;
        RECT 50.045 138.835 50.295 139.635 ;
        RECT 50.465 139.005 50.805 139.635 ;
        RECT 51.250 139.040 51.495 139.645 ;
        RECT 51.715 138.835 52.225 139.370 ;
        RECT 52.405 139.005 52.595 140.365 ;
        RECT 52.765 139.685 53.040 140.165 ;
        RECT 52.765 139.515 53.045 139.685 ;
        RECT 53.245 139.565 53.415 140.365 ;
        RECT 53.585 139.575 53.755 140.705 ;
        RECT 53.925 140.075 54.095 141.045 ;
        RECT 54.265 140.245 54.435 141.385 ;
        RECT 54.605 140.245 54.940 141.215 ;
        RECT 55.665 140.455 55.835 141.215 ;
        RECT 56.015 140.625 56.345 141.385 ;
        RECT 55.665 140.285 56.330 140.455 ;
        RECT 56.515 140.310 56.785 141.215 ;
        RECT 53.925 139.745 54.120 140.075 ;
        RECT 54.345 139.745 54.600 140.075 ;
        RECT 54.345 139.575 54.515 139.745 ;
        RECT 54.770 139.575 54.940 140.245 ;
        RECT 56.160 140.140 56.330 140.285 ;
        RECT 55.595 139.735 55.925 140.105 ;
        RECT 56.160 139.810 56.445 140.140 ;
        RECT 52.765 139.005 53.040 139.515 ;
        RECT 53.585 139.405 54.515 139.575 ;
        RECT 53.585 139.370 53.760 139.405 ;
        RECT 53.230 139.005 53.760 139.370 ;
        RECT 54.185 138.835 54.515 139.235 ;
        RECT 54.685 139.005 54.940 139.575 ;
        RECT 56.160 139.555 56.330 139.810 ;
        RECT 55.665 139.385 56.330 139.555 ;
        RECT 56.615 139.510 56.785 140.310 ;
        RECT 57.415 140.625 57.930 141.035 ;
        RECT 58.165 140.625 58.335 141.385 ;
        RECT 58.505 141.045 60.535 141.215 ;
        RECT 57.415 139.815 57.755 140.625 ;
        RECT 58.505 140.380 58.675 141.045 ;
        RECT 59.070 140.705 60.195 140.875 ;
        RECT 57.925 140.190 58.675 140.380 ;
        RECT 58.845 140.365 59.855 140.535 ;
        RECT 57.415 139.645 58.645 139.815 ;
        RECT 55.665 139.005 55.835 139.385 ;
        RECT 56.015 138.835 56.345 139.215 ;
        RECT 56.525 139.005 56.785 139.510 ;
        RECT 57.690 139.040 57.935 139.645 ;
        RECT 58.155 138.835 58.665 139.370 ;
        RECT 58.845 139.005 59.035 140.365 ;
        RECT 59.205 139.345 59.480 140.165 ;
        RECT 59.685 139.565 59.855 140.365 ;
        RECT 60.025 139.575 60.195 140.705 ;
        RECT 60.365 140.075 60.535 141.045 ;
        RECT 60.705 140.245 60.875 141.385 ;
        RECT 61.045 140.245 61.380 141.215 ;
        RECT 60.365 139.745 60.560 140.075 ;
        RECT 60.785 139.745 61.040 140.075 ;
        RECT 60.785 139.575 60.955 139.745 ;
        RECT 61.210 139.575 61.380 140.245 ;
        RECT 61.555 140.220 61.845 141.385 ;
        RECT 62.995 140.245 63.205 141.385 ;
        RECT 63.375 140.235 63.705 141.215 ;
        RECT 63.875 140.245 64.105 141.385 ;
        RECT 64.865 140.455 65.035 141.215 ;
        RECT 65.215 140.625 65.545 141.385 ;
        RECT 64.865 140.285 65.530 140.455 ;
        RECT 65.715 140.310 65.985 141.215 ;
        RECT 60.025 139.405 60.955 139.575 ;
        RECT 60.025 139.370 60.200 139.405 ;
        RECT 59.205 139.175 59.485 139.345 ;
        RECT 59.205 139.005 59.480 139.175 ;
        RECT 59.670 139.005 60.200 139.370 ;
        RECT 60.625 138.835 60.955 139.235 ;
        RECT 61.125 139.005 61.380 139.575 ;
        RECT 61.555 138.835 61.845 139.560 ;
        RECT 62.995 138.835 63.205 139.655 ;
        RECT 63.375 139.635 63.625 140.235 ;
        RECT 65.360 140.140 65.530 140.285 ;
        RECT 63.795 139.825 64.125 140.075 ;
        RECT 64.795 139.735 65.125 140.105 ;
        RECT 65.360 139.810 65.645 140.140 ;
        RECT 63.375 139.005 63.705 139.635 ;
        RECT 63.875 138.835 64.105 139.655 ;
        RECT 65.360 139.555 65.530 139.810 ;
        RECT 64.865 139.385 65.530 139.555 ;
        RECT 65.815 139.510 65.985 140.310 ;
        RECT 67.075 140.295 70.585 141.385 ;
        RECT 70.760 140.875 72.415 141.165 ;
        RECT 70.760 140.535 72.350 140.705 ;
        RECT 72.585 140.585 72.865 141.385 ;
        RECT 67.075 139.775 68.765 140.295 ;
        RECT 70.760 140.245 71.080 140.535 ;
        RECT 72.180 140.415 72.350 140.535 ;
        RECT 68.935 139.605 70.585 140.125 ;
        RECT 64.865 139.005 65.035 139.385 ;
        RECT 65.215 138.835 65.545 139.215 ;
        RECT 65.725 139.005 65.985 139.510 ;
        RECT 67.075 138.835 70.585 139.605 ;
        RECT 70.760 139.505 71.110 140.075 ;
        RECT 71.280 139.745 71.990 140.365 ;
        RECT 72.180 140.245 72.905 140.415 ;
        RECT 73.075 140.245 73.345 141.215 ;
        RECT 72.735 140.075 72.905 140.245 ;
        RECT 72.160 139.745 72.565 140.075 ;
        RECT 72.735 139.745 73.005 140.075 ;
        RECT 72.735 139.575 72.905 139.745 ;
        RECT 71.295 139.405 72.905 139.575 ;
        RECT 73.175 139.510 73.345 140.245 ;
        RECT 73.515 140.625 74.030 141.035 ;
        RECT 74.265 140.625 74.435 141.385 ;
        RECT 74.605 141.045 76.635 141.215 ;
        RECT 73.515 139.815 73.855 140.625 ;
        RECT 74.605 140.380 74.775 141.045 ;
        RECT 75.170 140.705 76.295 140.875 ;
        RECT 74.025 140.190 74.775 140.380 ;
        RECT 74.945 140.365 75.955 140.535 ;
        RECT 73.515 139.645 74.745 139.815 ;
        RECT 70.765 138.835 71.095 139.335 ;
        RECT 71.295 139.055 71.465 139.405 ;
        RECT 71.665 138.835 71.995 139.235 ;
        RECT 72.165 139.055 72.335 139.405 ;
        RECT 72.505 138.835 72.885 139.235 ;
        RECT 73.075 139.165 73.345 139.510 ;
        RECT 73.790 139.040 74.035 139.645 ;
        RECT 74.255 138.835 74.765 139.370 ;
        RECT 74.945 139.005 75.135 140.365 ;
        RECT 75.305 139.345 75.580 140.165 ;
        RECT 75.785 139.565 75.955 140.365 ;
        RECT 76.125 139.575 76.295 140.705 ;
        RECT 76.465 140.075 76.635 141.045 ;
        RECT 76.805 140.245 76.975 141.385 ;
        RECT 77.145 140.245 77.480 141.215 ;
        RECT 76.465 139.745 76.660 140.075 ;
        RECT 76.885 139.745 77.140 140.075 ;
        RECT 76.885 139.575 77.055 139.745 ;
        RECT 77.310 139.575 77.480 140.245 ;
        RECT 78.030 140.405 78.285 141.075 ;
        RECT 78.465 140.585 78.750 141.385 ;
        RECT 78.930 140.665 79.260 141.175 ;
        RECT 78.030 139.685 78.210 140.405 ;
        RECT 78.930 140.075 79.180 140.665 ;
        RECT 79.530 140.515 79.700 141.125 ;
        RECT 79.870 140.695 80.200 141.385 ;
        RECT 80.430 140.835 80.670 141.125 ;
        RECT 80.870 141.005 81.290 141.385 ;
        RECT 81.470 140.915 82.100 141.165 ;
        RECT 82.570 141.005 82.900 141.385 ;
        RECT 81.470 140.835 81.640 140.915 ;
        RECT 83.070 140.835 83.240 141.125 ;
        RECT 83.420 141.005 83.800 141.385 ;
        RECT 84.040 141.000 84.870 141.170 ;
        RECT 80.430 140.665 81.640 140.835 ;
        RECT 78.380 139.745 79.180 140.075 ;
        RECT 76.125 139.405 77.055 139.575 ;
        RECT 76.125 139.370 76.300 139.405 ;
        RECT 75.305 139.175 75.585 139.345 ;
        RECT 75.305 139.005 75.580 139.175 ;
        RECT 75.770 139.005 76.300 139.370 ;
        RECT 76.725 138.835 77.055 139.235 ;
        RECT 77.225 139.005 77.480 139.575 ;
        RECT 77.945 139.545 78.210 139.685 ;
        RECT 77.945 139.515 78.285 139.545 ;
        RECT 78.030 139.015 78.285 139.515 ;
        RECT 78.465 138.835 78.750 139.295 ;
        RECT 78.930 139.095 79.180 139.745 ;
        RECT 79.380 140.495 79.700 140.515 ;
        RECT 79.380 140.325 81.300 140.495 ;
        RECT 79.380 139.430 79.570 140.325 ;
        RECT 81.470 140.155 81.640 140.665 ;
        RECT 81.810 140.405 82.330 140.715 ;
        RECT 79.740 139.985 81.640 140.155 ;
        RECT 79.740 139.925 80.070 139.985 ;
        RECT 80.220 139.755 80.550 139.815 ;
        RECT 79.890 139.485 80.550 139.755 ;
        RECT 79.380 139.100 79.700 139.430 ;
        RECT 79.880 138.835 80.540 139.315 ;
        RECT 80.740 139.225 80.910 139.985 ;
        RECT 81.810 139.815 81.990 140.225 ;
        RECT 81.080 139.645 81.410 139.765 ;
        RECT 82.160 139.645 82.330 140.405 ;
        RECT 81.080 139.475 82.330 139.645 ;
        RECT 82.500 140.585 83.870 140.835 ;
        RECT 82.500 139.815 82.690 140.585 ;
        RECT 83.620 140.325 83.870 140.585 ;
        RECT 82.860 140.155 83.110 140.315 ;
        RECT 84.040 140.155 84.210 141.000 ;
        RECT 85.105 140.715 85.275 141.215 ;
        RECT 85.445 140.885 85.775 141.385 ;
        RECT 84.380 140.325 84.880 140.705 ;
        RECT 85.105 140.545 85.800 140.715 ;
        RECT 82.860 139.985 84.210 140.155 ;
        RECT 83.790 139.945 84.210 139.985 ;
        RECT 82.500 139.475 82.920 139.815 ;
        RECT 83.210 139.485 83.620 139.815 ;
        RECT 80.740 139.055 81.590 139.225 ;
        RECT 82.150 138.835 82.470 139.295 ;
        RECT 82.670 139.045 82.920 139.475 ;
        RECT 83.210 138.835 83.620 139.275 ;
        RECT 83.790 139.215 83.960 139.945 ;
        RECT 84.130 139.395 84.480 139.765 ;
        RECT 84.660 139.455 84.880 140.325 ;
        RECT 85.050 139.755 85.460 140.375 ;
        RECT 85.630 139.575 85.800 140.545 ;
        RECT 85.105 139.385 85.800 139.575 ;
        RECT 83.790 139.015 84.805 139.215 ;
        RECT 85.105 139.055 85.275 139.385 ;
        RECT 85.445 138.835 85.775 139.215 ;
        RECT 85.990 139.095 86.215 141.215 ;
        RECT 86.385 140.885 86.715 141.385 ;
        RECT 86.885 140.715 87.055 141.215 ;
        RECT 86.390 140.545 87.055 140.715 ;
        RECT 86.390 139.555 86.620 140.545 ;
        RECT 86.790 139.725 87.140 140.375 ;
        RECT 87.315 140.220 87.605 141.385 ;
        RECT 88.150 141.045 88.405 141.075 ;
        RECT 88.065 140.875 88.405 141.045 ;
        RECT 88.150 140.405 88.405 140.875 ;
        RECT 88.585 140.585 88.870 141.385 ;
        RECT 89.050 140.665 89.380 141.175 ;
        RECT 86.390 139.385 87.055 139.555 ;
        RECT 86.385 138.835 86.715 139.215 ;
        RECT 86.885 139.095 87.055 139.385 ;
        RECT 87.315 138.835 87.605 139.560 ;
        RECT 88.150 139.545 88.330 140.405 ;
        RECT 89.050 140.075 89.300 140.665 ;
        RECT 89.650 140.515 89.820 141.125 ;
        RECT 89.990 140.695 90.320 141.385 ;
        RECT 90.550 140.835 90.790 141.125 ;
        RECT 90.990 141.005 91.410 141.385 ;
        RECT 91.590 140.915 92.220 141.165 ;
        RECT 92.690 141.005 93.020 141.385 ;
        RECT 91.590 140.835 91.760 140.915 ;
        RECT 93.190 140.835 93.360 141.125 ;
        RECT 93.540 141.005 93.920 141.385 ;
        RECT 94.160 141.000 94.990 141.170 ;
        RECT 90.550 140.665 91.760 140.835 ;
        RECT 88.500 139.745 89.300 140.075 ;
        RECT 88.150 139.015 88.405 139.545 ;
        RECT 88.585 138.835 88.870 139.295 ;
        RECT 89.050 139.095 89.300 139.745 ;
        RECT 89.500 140.495 89.820 140.515 ;
        RECT 89.500 140.325 91.420 140.495 ;
        RECT 89.500 139.430 89.690 140.325 ;
        RECT 91.590 140.155 91.760 140.665 ;
        RECT 91.930 140.405 92.450 140.715 ;
        RECT 89.860 139.985 91.760 140.155 ;
        RECT 89.860 139.925 90.190 139.985 ;
        RECT 90.340 139.755 90.670 139.815 ;
        RECT 90.010 139.485 90.670 139.755 ;
        RECT 89.500 139.100 89.820 139.430 ;
        RECT 90.000 138.835 90.660 139.315 ;
        RECT 90.860 139.225 91.030 139.985 ;
        RECT 91.930 139.815 92.110 140.225 ;
        RECT 91.200 139.645 91.530 139.765 ;
        RECT 92.280 139.645 92.450 140.405 ;
        RECT 91.200 139.475 92.450 139.645 ;
        RECT 92.620 140.585 93.990 140.835 ;
        RECT 92.620 139.815 92.810 140.585 ;
        RECT 93.740 140.325 93.990 140.585 ;
        RECT 92.980 140.155 93.230 140.315 ;
        RECT 94.160 140.155 94.330 141.000 ;
        RECT 95.225 140.715 95.395 141.215 ;
        RECT 95.565 140.885 95.895 141.385 ;
        RECT 94.500 140.325 95.000 140.705 ;
        RECT 95.225 140.545 95.920 140.715 ;
        RECT 92.980 139.985 94.330 140.155 ;
        RECT 93.910 139.945 94.330 139.985 ;
        RECT 92.620 139.475 93.040 139.815 ;
        RECT 93.330 139.485 93.740 139.815 ;
        RECT 90.860 139.055 91.710 139.225 ;
        RECT 92.270 138.835 92.590 139.295 ;
        RECT 92.790 139.045 93.040 139.475 ;
        RECT 93.330 138.835 93.740 139.275 ;
        RECT 93.910 139.215 94.080 139.945 ;
        RECT 94.250 139.395 94.600 139.765 ;
        RECT 94.780 139.455 95.000 140.325 ;
        RECT 95.170 139.755 95.580 140.375 ;
        RECT 95.750 139.575 95.920 140.545 ;
        RECT 95.225 139.385 95.920 139.575 ;
        RECT 93.910 139.015 94.925 139.215 ;
        RECT 95.225 139.055 95.395 139.385 ;
        RECT 95.565 138.835 95.895 139.215 ;
        RECT 96.110 139.095 96.335 141.215 ;
        RECT 96.505 140.885 96.835 141.385 ;
        RECT 97.005 140.715 97.175 141.215 ;
        RECT 96.510 140.545 97.175 140.715 ;
        RECT 96.510 139.555 96.740 140.545 ;
        RECT 96.910 139.725 97.260 140.375 ;
        RECT 97.435 140.310 97.705 141.215 ;
        RECT 97.875 140.625 98.205 141.385 ;
        RECT 98.385 140.455 98.555 141.215 ;
        RECT 96.510 139.385 97.175 139.555 ;
        RECT 96.505 138.835 96.835 139.215 ;
        RECT 97.005 139.095 97.175 139.385 ;
        RECT 97.435 139.510 97.605 140.310 ;
        RECT 97.890 140.285 98.555 140.455 ;
        RECT 99.650 140.405 99.905 141.075 ;
        RECT 100.085 140.585 100.370 141.385 ;
        RECT 100.550 140.665 100.880 141.175 ;
        RECT 97.890 140.140 98.060 140.285 ;
        RECT 97.775 139.810 98.060 140.140 ;
        RECT 97.890 139.555 98.060 139.810 ;
        RECT 98.295 139.735 98.625 140.105 ;
        RECT 97.435 139.005 97.695 139.510 ;
        RECT 97.890 139.385 98.555 139.555 ;
        RECT 97.875 138.835 98.205 139.215 ;
        RECT 98.385 139.005 98.555 139.385 ;
        RECT 99.650 139.545 99.830 140.405 ;
        RECT 100.550 140.075 100.800 140.665 ;
        RECT 101.150 140.515 101.320 141.125 ;
        RECT 101.490 140.695 101.820 141.385 ;
        RECT 102.050 140.835 102.290 141.125 ;
        RECT 102.490 141.005 102.910 141.385 ;
        RECT 103.090 140.915 103.720 141.165 ;
        RECT 104.190 141.005 104.520 141.385 ;
        RECT 103.090 140.835 103.260 140.915 ;
        RECT 104.690 140.835 104.860 141.125 ;
        RECT 105.040 141.005 105.420 141.385 ;
        RECT 105.660 141.000 106.490 141.170 ;
        RECT 102.050 140.665 103.260 140.835 ;
        RECT 100.000 139.745 100.800 140.075 ;
        RECT 99.650 139.345 99.905 139.545 ;
        RECT 99.565 139.175 99.905 139.345 ;
        RECT 99.650 139.015 99.905 139.175 ;
        RECT 100.085 138.835 100.370 139.295 ;
        RECT 100.550 139.095 100.800 139.745 ;
        RECT 101.000 140.495 101.320 140.515 ;
        RECT 101.000 140.325 102.920 140.495 ;
        RECT 101.000 139.430 101.190 140.325 ;
        RECT 103.090 140.155 103.260 140.665 ;
        RECT 103.430 140.405 103.950 140.715 ;
        RECT 101.360 139.985 103.260 140.155 ;
        RECT 101.360 139.925 101.690 139.985 ;
        RECT 101.840 139.755 102.170 139.815 ;
        RECT 101.510 139.485 102.170 139.755 ;
        RECT 101.000 139.100 101.320 139.430 ;
        RECT 101.500 138.835 102.160 139.315 ;
        RECT 102.360 139.225 102.530 139.985 ;
        RECT 103.430 139.815 103.610 140.225 ;
        RECT 102.700 139.645 103.030 139.765 ;
        RECT 103.780 139.645 103.950 140.405 ;
        RECT 102.700 139.475 103.950 139.645 ;
        RECT 104.120 140.585 105.490 140.835 ;
        RECT 104.120 139.815 104.310 140.585 ;
        RECT 105.240 140.325 105.490 140.585 ;
        RECT 104.480 140.155 104.730 140.315 ;
        RECT 105.660 140.155 105.830 141.000 ;
        RECT 106.725 140.715 106.895 141.215 ;
        RECT 107.065 140.885 107.395 141.385 ;
        RECT 106.000 140.325 106.500 140.705 ;
        RECT 106.725 140.545 107.420 140.715 ;
        RECT 104.480 139.985 105.830 140.155 ;
        RECT 105.410 139.945 105.830 139.985 ;
        RECT 104.120 139.475 104.540 139.815 ;
        RECT 104.830 139.485 105.240 139.815 ;
        RECT 102.360 139.055 103.210 139.225 ;
        RECT 103.770 138.835 104.090 139.295 ;
        RECT 104.290 139.045 104.540 139.475 ;
        RECT 104.830 138.835 105.240 139.275 ;
        RECT 105.410 139.215 105.580 139.945 ;
        RECT 105.750 139.395 106.100 139.765 ;
        RECT 106.280 139.455 106.500 140.325 ;
        RECT 106.670 139.755 107.080 140.375 ;
        RECT 107.250 139.575 107.420 140.545 ;
        RECT 106.725 139.385 107.420 139.575 ;
        RECT 105.410 139.015 106.425 139.215 ;
        RECT 106.725 139.055 106.895 139.385 ;
        RECT 107.065 138.835 107.395 139.215 ;
        RECT 107.610 139.095 107.835 141.215 ;
        RECT 108.005 140.885 108.335 141.385 ;
        RECT 108.505 140.715 108.675 141.215 ;
        RECT 108.010 140.545 108.675 140.715 ;
        RECT 108.010 139.555 108.240 140.545 ;
        RECT 109.025 140.455 109.195 141.215 ;
        RECT 109.375 140.625 109.705 141.385 ;
        RECT 108.410 139.725 108.760 140.375 ;
        RECT 109.025 140.285 109.690 140.455 ;
        RECT 109.875 140.310 110.145 141.215 ;
        RECT 109.520 140.140 109.690 140.285 ;
        RECT 108.955 139.735 109.285 140.105 ;
        RECT 109.520 139.810 109.805 140.140 ;
        RECT 109.520 139.555 109.690 139.810 ;
        RECT 108.010 139.385 108.675 139.555 ;
        RECT 108.005 138.835 108.335 139.215 ;
        RECT 108.505 139.095 108.675 139.385 ;
        RECT 109.025 139.385 109.690 139.555 ;
        RECT 109.975 139.510 110.145 140.310 ;
        RECT 110.315 140.295 111.985 141.385 ;
        RECT 112.155 140.295 113.365 141.385 ;
        RECT 110.315 139.775 111.065 140.295 ;
        RECT 111.235 139.605 111.985 140.125 ;
        RECT 112.155 139.755 112.675 140.295 ;
        RECT 109.025 139.005 109.195 139.385 ;
        RECT 109.375 138.835 109.705 139.215 ;
        RECT 109.885 139.005 110.145 139.510 ;
        RECT 110.315 138.835 111.985 139.605 ;
        RECT 112.845 139.585 113.365 140.125 ;
        RECT 112.155 138.835 113.365 139.585 ;
        RECT 15.010 138.665 113.450 138.835 ;
        RECT 15.095 137.915 16.305 138.665 ;
        RECT 17.485 138.115 17.655 138.495 ;
        RECT 17.835 138.285 18.165 138.665 ;
        RECT 17.485 137.945 18.150 138.115 ;
        RECT 18.345 137.990 18.605 138.495 ;
        RECT 15.095 137.375 15.615 137.915 ;
        RECT 15.785 137.205 16.305 137.745 ;
        RECT 17.415 137.395 17.745 137.765 ;
        RECT 17.980 137.690 18.150 137.945 ;
        RECT 17.980 137.360 18.265 137.690 ;
        RECT 17.980 137.215 18.150 137.360 ;
        RECT 15.095 136.115 16.305 137.205 ;
        RECT 17.485 137.045 18.150 137.215 ;
        RECT 18.435 137.190 18.605 137.990 ;
        RECT 17.485 136.285 17.655 137.045 ;
        RECT 17.835 136.115 18.165 136.875 ;
        RECT 18.335 136.285 18.605 137.190 ;
        RECT 18.780 137.925 19.035 138.495 ;
        RECT 19.205 138.265 19.535 138.665 ;
        RECT 19.960 138.130 20.490 138.495 ;
        RECT 20.680 138.325 20.955 138.495 ;
        RECT 20.675 138.155 20.955 138.325 ;
        RECT 19.960 138.095 20.135 138.130 ;
        RECT 19.205 137.925 20.135 138.095 ;
        RECT 18.780 137.255 18.950 137.925 ;
        RECT 19.205 137.755 19.375 137.925 ;
        RECT 19.120 137.425 19.375 137.755 ;
        RECT 19.600 137.425 19.795 137.755 ;
        RECT 18.780 136.285 19.115 137.255 ;
        RECT 19.285 136.115 19.455 137.255 ;
        RECT 19.625 136.455 19.795 137.425 ;
        RECT 19.965 136.795 20.135 137.925 ;
        RECT 20.305 137.135 20.475 137.935 ;
        RECT 20.680 137.335 20.955 138.155 ;
        RECT 21.125 137.135 21.315 138.495 ;
        RECT 21.495 138.130 22.005 138.665 ;
        RECT 22.225 137.855 22.470 138.460 ;
        RECT 22.915 137.940 23.205 138.665 ;
        RECT 21.515 137.685 22.745 137.855 ;
        RECT 23.415 137.845 23.645 138.665 ;
        RECT 23.815 137.865 24.145 138.495 ;
        RECT 20.305 136.965 21.315 137.135 ;
        RECT 21.485 137.120 22.235 137.310 ;
        RECT 19.965 136.625 21.090 136.795 ;
        RECT 21.485 136.455 21.655 137.120 ;
        RECT 22.405 136.875 22.745 137.685 ;
        RECT 23.395 137.425 23.725 137.675 ;
        RECT 19.625 136.285 21.655 136.455 ;
        RECT 21.825 136.115 21.995 136.875 ;
        RECT 22.230 136.465 22.745 136.875 ;
        RECT 22.915 136.115 23.205 137.280 ;
        RECT 23.895 137.265 24.145 137.865 ;
        RECT 24.315 137.845 24.525 138.665 ;
        RECT 24.955 138.035 25.285 138.395 ;
        RECT 25.905 138.205 26.155 138.665 ;
        RECT 26.325 138.205 26.885 138.495 ;
        RECT 24.955 137.845 26.345 138.035 ;
        RECT 26.175 137.755 26.345 137.845 ;
        RECT 23.415 136.115 23.645 137.255 ;
        RECT 23.815 136.285 24.145 137.265 ;
        RECT 24.770 137.425 25.445 137.675 ;
        RECT 25.665 137.425 26.005 137.675 ;
        RECT 26.175 137.425 26.465 137.755 ;
        RECT 24.315 136.115 24.525 137.255 ;
        RECT 24.770 137.065 25.035 137.425 ;
        RECT 26.175 137.175 26.345 137.425 ;
        RECT 25.405 137.005 26.345 137.175 ;
        RECT 24.955 136.115 25.235 136.785 ;
        RECT 25.405 136.455 25.705 137.005 ;
        RECT 26.635 136.835 26.885 138.205 ;
        RECT 25.905 136.115 26.235 136.835 ;
        RECT 26.425 136.285 26.885 136.835 ;
        RECT 27.060 137.925 27.315 138.495 ;
        RECT 27.485 138.265 27.815 138.665 ;
        RECT 28.240 138.130 28.770 138.495 ;
        RECT 28.240 138.095 28.415 138.130 ;
        RECT 27.485 137.925 28.415 138.095 ;
        RECT 28.960 137.985 29.235 138.495 ;
        RECT 27.060 137.255 27.230 137.925 ;
        RECT 27.485 137.755 27.655 137.925 ;
        RECT 27.400 137.425 27.655 137.755 ;
        RECT 27.880 137.425 28.075 137.755 ;
        RECT 27.060 136.285 27.395 137.255 ;
        RECT 27.565 136.115 27.735 137.255 ;
        RECT 27.905 136.455 28.075 137.425 ;
        RECT 28.245 136.795 28.415 137.925 ;
        RECT 28.585 137.135 28.755 137.935 ;
        RECT 28.955 137.815 29.235 137.985 ;
        RECT 28.960 137.335 29.235 137.815 ;
        RECT 29.405 137.135 29.595 138.495 ;
        RECT 29.775 138.130 30.285 138.665 ;
        RECT 30.505 137.855 30.750 138.460 ;
        RECT 31.305 138.185 31.475 138.665 ;
        RECT 31.645 138.015 31.975 138.490 ;
        RECT 32.145 138.185 32.315 138.665 ;
        RECT 32.485 138.015 32.815 138.490 ;
        RECT 32.985 138.185 33.155 138.665 ;
        RECT 33.325 138.015 33.655 138.490 ;
        RECT 33.825 138.185 33.995 138.665 ;
        RECT 34.165 138.015 34.495 138.490 ;
        RECT 34.665 138.185 34.835 138.665 ;
        RECT 35.005 138.015 35.335 138.490 ;
        RECT 35.505 138.185 35.675 138.665 ;
        RECT 35.925 138.490 36.095 138.495 ;
        RECT 35.845 138.015 36.175 138.490 ;
        RECT 36.345 138.185 36.515 138.665 ;
        RECT 36.765 138.490 36.935 138.495 ;
        RECT 36.685 138.015 37.015 138.490 ;
        RECT 37.185 138.185 37.355 138.665 ;
        RECT 37.605 138.490 37.855 138.495 ;
        RECT 37.525 138.015 37.855 138.490 ;
        RECT 38.025 138.185 38.195 138.665 ;
        RECT 38.365 138.015 38.695 138.490 ;
        RECT 38.865 138.185 39.035 138.665 ;
        RECT 39.205 138.015 39.535 138.490 ;
        RECT 39.705 138.185 39.875 138.665 ;
        RECT 40.045 138.015 40.375 138.490 ;
        RECT 40.545 138.185 40.715 138.665 ;
        RECT 40.885 138.015 41.215 138.490 ;
        RECT 41.385 138.185 41.555 138.665 ;
        RECT 41.725 138.015 42.055 138.490 ;
        RECT 29.795 137.685 31.025 137.855 ;
        RECT 28.585 136.965 29.595 137.135 ;
        RECT 29.765 137.120 30.515 137.310 ;
        RECT 28.245 136.625 29.370 136.795 ;
        RECT 29.765 136.455 29.935 137.120 ;
        RECT 30.685 136.875 31.025 137.685 ;
        RECT 31.195 137.845 37.855 138.015 ;
        RECT 38.025 137.845 40.375 138.015 ;
        RECT 40.545 137.845 42.055 138.015 ;
        RECT 42.235 137.990 42.505 138.335 ;
        RECT 42.695 138.265 43.075 138.665 ;
        RECT 43.245 138.095 43.415 138.445 ;
        RECT 43.585 138.265 43.915 138.665 ;
        RECT 44.115 138.095 44.285 138.445 ;
        RECT 44.485 138.165 44.815 138.665 ;
        RECT 31.195 137.305 31.470 137.845 ;
        RECT 38.025 137.675 38.200 137.845 ;
        RECT 40.545 137.675 40.715 137.845 ;
        RECT 31.640 137.475 38.200 137.675 ;
        RECT 38.405 137.475 40.715 137.675 ;
        RECT 40.885 137.475 42.060 137.675 ;
        RECT 38.025 137.305 38.200 137.475 ;
        RECT 40.545 137.305 40.715 137.475 ;
        RECT 31.195 137.135 37.855 137.305 ;
        RECT 38.025 137.135 40.375 137.305 ;
        RECT 40.545 137.135 42.055 137.305 ;
        RECT 27.905 136.285 29.935 136.455 ;
        RECT 30.105 136.115 30.275 136.875 ;
        RECT 30.510 136.465 31.025 136.875 ;
        RECT 31.305 136.115 31.475 136.915 ;
        RECT 31.645 136.285 31.975 137.135 ;
        RECT 32.145 136.115 32.315 136.915 ;
        RECT 32.485 136.285 32.815 137.135 ;
        RECT 32.985 136.115 33.155 136.915 ;
        RECT 33.325 136.285 33.655 137.135 ;
        RECT 33.825 136.115 33.995 136.915 ;
        RECT 34.165 136.285 34.495 137.135 ;
        RECT 34.665 136.115 34.835 136.915 ;
        RECT 35.005 136.285 35.335 137.135 ;
        RECT 35.505 136.115 35.675 136.915 ;
        RECT 35.845 136.285 36.175 137.135 ;
        RECT 36.345 136.115 36.515 136.915 ;
        RECT 36.685 136.285 37.015 137.135 ;
        RECT 37.185 136.115 37.355 136.915 ;
        RECT 37.525 136.285 37.855 137.135 ;
        RECT 38.025 136.115 38.195 136.915 ;
        RECT 38.365 136.285 38.695 137.135 ;
        RECT 38.865 136.115 39.035 136.915 ;
        RECT 39.205 136.285 39.535 137.135 ;
        RECT 39.705 136.115 39.875 136.915 ;
        RECT 40.045 136.285 40.375 137.135 ;
        RECT 40.545 136.115 40.715 136.965 ;
        RECT 40.885 136.285 41.215 137.135 ;
        RECT 41.385 136.115 41.555 136.965 ;
        RECT 41.725 136.285 42.055 137.135 ;
        RECT 42.235 137.255 42.405 137.990 ;
        RECT 42.675 137.925 44.285 138.095 ;
        RECT 42.675 137.755 42.845 137.925 ;
        RECT 42.575 137.425 42.845 137.755 ;
        RECT 43.015 137.425 43.420 137.755 ;
        RECT 42.675 137.255 42.845 137.425 ;
        RECT 43.590 137.305 44.300 137.755 ;
        RECT 44.470 137.425 44.820 137.995 ;
        RECT 44.995 137.865 45.335 138.495 ;
        RECT 45.505 137.865 45.755 138.665 ;
        RECT 45.945 138.015 46.275 138.495 ;
        RECT 46.445 138.205 46.670 138.665 ;
        RECT 46.840 138.015 47.170 138.495 ;
        RECT 44.995 137.815 45.225 137.865 ;
        RECT 45.945 137.845 47.170 138.015 ;
        RECT 47.800 137.885 48.300 138.495 ;
        RECT 48.675 137.940 48.965 138.665 ;
        RECT 50.430 137.955 50.685 138.485 ;
        RECT 50.865 138.205 51.150 138.665 ;
        RECT 42.235 136.285 42.505 137.255 ;
        RECT 42.675 137.085 43.400 137.255 ;
        RECT 43.590 137.135 44.305 137.305 ;
        RECT 44.995 137.255 45.170 137.815 ;
        RECT 45.340 137.505 46.035 137.675 ;
        RECT 45.865 137.255 46.035 137.505 ;
        RECT 46.210 137.475 46.630 137.675 ;
        RECT 46.800 137.475 47.130 137.675 ;
        RECT 47.300 137.475 47.630 137.675 ;
        RECT 47.800 137.255 47.970 137.885 ;
        RECT 48.155 137.425 48.505 137.675 ;
        RECT 43.230 136.965 43.400 137.085 ;
        RECT 44.500 136.965 44.820 137.255 ;
        RECT 42.715 136.115 42.995 136.915 ;
        RECT 43.230 136.795 44.820 136.965 ;
        RECT 43.165 136.335 44.820 136.625 ;
        RECT 44.995 136.285 45.335 137.255 ;
        RECT 45.505 136.115 45.675 137.255 ;
        RECT 45.865 137.085 48.300 137.255 ;
        RECT 45.945 136.115 46.195 136.915 ;
        RECT 46.840 136.285 47.170 137.085 ;
        RECT 47.470 136.115 47.800 136.915 ;
        RECT 47.970 136.285 48.300 137.085 ;
        RECT 48.675 136.115 48.965 137.280 ;
        RECT 50.430 137.095 50.610 137.955 ;
        RECT 51.330 137.755 51.580 138.405 ;
        RECT 50.780 137.425 51.580 137.755 ;
        RECT 50.430 136.625 50.685 137.095 ;
        RECT 50.345 136.455 50.685 136.625 ;
        RECT 50.430 136.425 50.685 136.455 ;
        RECT 50.865 136.115 51.150 136.915 ;
        RECT 51.330 136.835 51.580 137.425 ;
        RECT 51.780 138.070 52.100 138.400 ;
        RECT 52.280 138.185 52.940 138.665 ;
        RECT 53.140 138.275 53.990 138.445 ;
        RECT 51.780 137.175 51.970 138.070 ;
        RECT 52.290 137.745 52.950 138.015 ;
        RECT 52.620 137.685 52.950 137.745 ;
        RECT 52.140 137.515 52.470 137.575 ;
        RECT 53.140 137.515 53.310 138.275 ;
        RECT 54.550 138.205 54.870 138.665 ;
        RECT 55.070 138.025 55.320 138.455 ;
        RECT 55.610 138.225 56.020 138.665 ;
        RECT 56.190 138.285 57.205 138.485 ;
        RECT 53.480 137.855 54.730 138.025 ;
        RECT 53.480 137.735 53.810 137.855 ;
        RECT 52.140 137.345 54.040 137.515 ;
        RECT 51.780 137.005 53.700 137.175 ;
        RECT 51.780 136.985 52.100 137.005 ;
        RECT 51.330 136.325 51.660 136.835 ;
        RECT 51.930 136.375 52.100 136.985 ;
        RECT 53.870 136.835 54.040 137.345 ;
        RECT 54.210 137.275 54.390 137.685 ;
        RECT 54.560 137.095 54.730 137.855 ;
        RECT 52.270 136.115 52.600 136.805 ;
        RECT 52.830 136.665 54.040 136.835 ;
        RECT 54.210 136.785 54.730 137.095 ;
        RECT 54.900 137.685 55.320 138.025 ;
        RECT 55.610 137.685 56.020 138.015 ;
        RECT 54.900 136.915 55.090 137.685 ;
        RECT 56.190 137.555 56.360 138.285 ;
        RECT 57.505 138.115 57.675 138.445 ;
        RECT 57.845 138.285 58.175 138.665 ;
        RECT 56.530 137.735 56.880 138.105 ;
        RECT 56.190 137.515 56.610 137.555 ;
        RECT 55.260 137.345 56.610 137.515 ;
        RECT 55.260 137.185 55.510 137.345 ;
        RECT 56.020 136.915 56.270 137.175 ;
        RECT 54.900 136.665 56.270 136.915 ;
        RECT 52.830 136.375 53.070 136.665 ;
        RECT 53.870 136.585 54.040 136.665 ;
        RECT 53.270 136.115 53.690 136.495 ;
        RECT 53.870 136.335 54.500 136.585 ;
        RECT 54.970 136.115 55.300 136.495 ;
        RECT 55.470 136.375 55.640 136.665 ;
        RECT 56.440 136.500 56.610 137.345 ;
        RECT 57.060 137.175 57.280 138.045 ;
        RECT 57.505 137.925 58.200 138.115 ;
        RECT 56.780 136.795 57.280 137.175 ;
        RECT 57.450 137.125 57.860 137.745 ;
        RECT 58.030 136.955 58.200 137.925 ;
        RECT 57.505 136.785 58.200 136.955 ;
        RECT 55.820 136.115 56.200 136.495 ;
        RECT 56.440 136.330 57.270 136.500 ;
        RECT 57.505 136.285 57.675 136.785 ;
        RECT 57.845 136.115 58.175 136.615 ;
        RECT 58.390 136.285 58.615 138.405 ;
        RECT 58.785 138.285 59.115 138.665 ;
        RECT 59.285 138.115 59.455 138.405 ;
        RECT 58.790 137.945 59.455 138.115 ;
        RECT 58.790 136.955 59.020 137.945 ;
        RECT 59.715 137.895 62.305 138.665 ;
        RECT 62.480 138.120 67.825 138.665 ;
        RECT 68.005 138.165 68.335 138.665 ;
        RECT 59.190 137.125 59.540 137.775 ;
        RECT 59.715 137.205 60.925 137.725 ;
        RECT 61.095 137.375 62.305 137.895 ;
        RECT 58.790 136.785 59.455 136.955 ;
        RECT 58.785 136.115 59.115 136.615 ;
        RECT 59.285 136.285 59.455 136.785 ;
        RECT 59.715 136.115 62.305 137.205 ;
        RECT 64.070 136.550 64.420 137.800 ;
        RECT 65.900 137.290 66.240 138.120 ;
        RECT 68.535 138.095 68.705 138.445 ;
        RECT 68.905 138.265 69.235 138.665 ;
        RECT 69.405 138.095 69.575 138.445 ;
        RECT 69.745 138.265 70.125 138.665 ;
        RECT 68.000 137.425 68.350 137.995 ;
        RECT 68.535 137.925 70.145 138.095 ;
        RECT 70.315 137.990 70.585 138.335 ;
        RECT 69.975 137.755 70.145 137.925 ;
        RECT 68.520 137.305 69.230 137.755 ;
        RECT 69.400 137.425 69.805 137.755 ;
        RECT 69.975 137.425 70.245 137.755 ;
        RECT 68.000 136.965 68.320 137.255 ;
        RECT 68.515 137.135 69.230 137.305 ;
        RECT 69.975 137.255 70.145 137.425 ;
        RECT 70.415 137.255 70.585 137.990 ;
        RECT 69.420 137.085 70.145 137.255 ;
        RECT 69.420 136.965 69.590 137.085 ;
        RECT 68.000 136.795 69.590 136.965 ;
        RECT 62.480 136.115 67.825 136.550 ;
        RECT 68.000 136.335 69.655 136.625 ;
        RECT 69.825 136.115 70.105 136.915 ;
        RECT 70.315 136.285 70.585 137.255 ;
        RECT 70.755 137.865 71.095 138.495 ;
        RECT 71.265 137.865 71.515 138.665 ;
        RECT 71.705 138.015 72.035 138.495 ;
        RECT 72.205 138.205 72.430 138.665 ;
        RECT 72.600 138.015 72.930 138.495 ;
        RECT 70.755 137.815 70.985 137.865 ;
        RECT 71.705 137.845 72.930 138.015 ;
        RECT 73.560 137.885 74.060 138.495 ;
        RECT 74.435 137.940 74.725 138.665 ;
        RECT 75.270 137.985 75.525 138.485 ;
        RECT 75.705 138.205 75.990 138.665 ;
        RECT 75.185 137.955 75.525 137.985 ;
        RECT 70.755 137.255 70.930 137.815 ;
        RECT 71.100 137.505 71.795 137.675 ;
        RECT 71.625 137.255 71.795 137.505 ;
        RECT 71.970 137.475 72.390 137.675 ;
        RECT 72.560 137.475 72.890 137.675 ;
        RECT 73.060 137.475 73.390 137.675 ;
        RECT 73.560 137.255 73.730 137.885 ;
        RECT 75.185 137.815 75.450 137.955 ;
        RECT 73.915 137.425 74.265 137.675 ;
        RECT 70.755 136.285 71.095 137.255 ;
        RECT 71.265 136.115 71.435 137.255 ;
        RECT 71.625 137.085 74.060 137.255 ;
        RECT 71.705 136.115 71.955 136.915 ;
        RECT 72.600 136.285 72.930 137.085 ;
        RECT 73.230 136.115 73.560 136.915 ;
        RECT 73.730 136.285 74.060 137.085 ;
        RECT 74.435 136.115 74.725 137.280 ;
        RECT 75.270 137.095 75.450 137.815 ;
        RECT 76.170 137.755 76.420 138.405 ;
        RECT 75.620 137.425 76.420 137.755 ;
        RECT 75.270 136.425 75.525 137.095 ;
        RECT 75.705 136.115 75.990 136.915 ;
        RECT 76.170 136.835 76.420 137.425 ;
        RECT 76.620 138.070 76.940 138.400 ;
        RECT 77.120 138.185 77.780 138.665 ;
        RECT 77.980 138.275 78.830 138.445 ;
        RECT 76.620 137.175 76.810 138.070 ;
        RECT 77.130 137.745 77.790 138.015 ;
        RECT 77.460 137.685 77.790 137.745 ;
        RECT 76.980 137.515 77.310 137.575 ;
        RECT 77.980 137.515 78.150 138.275 ;
        RECT 79.390 138.205 79.710 138.665 ;
        RECT 79.910 138.025 80.160 138.455 ;
        RECT 80.450 138.225 80.860 138.665 ;
        RECT 81.030 138.285 82.045 138.485 ;
        RECT 78.320 137.855 79.570 138.025 ;
        RECT 78.320 137.735 78.650 137.855 ;
        RECT 76.980 137.345 78.880 137.515 ;
        RECT 76.620 137.005 78.540 137.175 ;
        RECT 76.620 136.985 76.940 137.005 ;
        RECT 76.170 136.325 76.500 136.835 ;
        RECT 76.770 136.375 76.940 136.985 ;
        RECT 78.710 136.835 78.880 137.345 ;
        RECT 79.050 137.275 79.230 137.685 ;
        RECT 79.400 137.095 79.570 137.855 ;
        RECT 77.110 136.115 77.440 136.805 ;
        RECT 77.670 136.665 78.880 136.835 ;
        RECT 79.050 136.785 79.570 137.095 ;
        RECT 79.740 137.685 80.160 138.025 ;
        RECT 80.450 137.685 80.860 138.015 ;
        RECT 79.740 136.915 79.930 137.685 ;
        RECT 81.030 137.555 81.200 138.285 ;
        RECT 82.345 138.115 82.515 138.445 ;
        RECT 82.685 138.285 83.015 138.665 ;
        RECT 81.370 137.735 81.720 138.105 ;
        RECT 81.030 137.515 81.450 137.555 ;
        RECT 80.100 137.345 81.450 137.515 ;
        RECT 80.100 137.185 80.350 137.345 ;
        RECT 80.860 136.915 81.110 137.175 ;
        RECT 79.740 136.665 81.110 136.915 ;
        RECT 77.670 136.375 77.910 136.665 ;
        RECT 78.710 136.585 78.880 136.665 ;
        RECT 78.110 136.115 78.530 136.495 ;
        RECT 78.710 136.335 79.340 136.585 ;
        RECT 79.810 136.115 80.140 136.495 ;
        RECT 80.310 136.375 80.480 136.665 ;
        RECT 81.280 136.500 81.450 137.345 ;
        RECT 81.900 137.175 82.120 138.045 ;
        RECT 82.345 137.925 83.040 138.115 ;
        RECT 81.620 136.795 82.120 137.175 ;
        RECT 82.290 137.125 82.700 137.745 ;
        RECT 82.870 136.955 83.040 137.925 ;
        RECT 82.345 136.785 83.040 136.955 ;
        RECT 80.660 136.115 81.040 136.495 ;
        RECT 81.280 136.330 82.110 136.500 ;
        RECT 82.345 136.285 82.515 136.785 ;
        RECT 82.685 136.115 83.015 136.615 ;
        RECT 83.230 136.285 83.455 138.405 ;
        RECT 83.625 138.285 83.955 138.665 ;
        RECT 84.125 138.115 84.295 138.405 ;
        RECT 83.630 137.945 84.295 138.115 ;
        RECT 83.630 136.955 83.860 137.945 ;
        RECT 84.615 137.845 84.825 138.665 ;
        RECT 84.995 137.865 85.325 138.495 ;
        RECT 84.030 137.125 84.380 137.775 ;
        RECT 84.995 137.265 85.245 137.865 ;
        RECT 85.495 137.845 85.725 138.665 ;
        RECT 86.395 137.990 86.655 138.495 ;
        RECT 86.835 138.285 87.165 138.665 ;
        RECT 87.345 138.115 87.515 138.495 ;
        RECT 85.415 137.425 85.745 137.675 ;
        RECT 83.630 136.785 84.295 136.955 ;
        RECT 83.625 136.115 83.955 136.615 ;
        RECT 84.125 136.285 84.295 136.785 ;
        RECT 84.615 136.115 84.825 137.255 ;
        RECT 84.995 136.285 85.325 137.265 ;
        RECT 85.495 136.115 85.725 137.255 ;
        RECT 86.395 137.190 86.565 137.990 ;
        RECT 86.850 137.945 87.515 138.115 ;
        RECT 86.850 137.690 87.020 137.945 ;
        RECT 87.775 137.895 90.365 138.665 ;
        RECT 86.735 137.360 87.020 137.690 ;
        RECT 87.255 137.395 87.585 137.765 ;
        RECT 86.850 137.215 87.020 137.360 ;
        RECT 86.395 136.285 86.665 137.190 ;
        RECT 86.850 137.045 87.515 137.215 ;
        RECT 86.835 136.115 87.165 136.875 ;
        RECT 87.345 136.285 87.515 137.045 ;
        RECT 87.775 137.205 88.985 137.725 ;
        RECT 89.155 137.375 90.365 137.895 ;
        RECT 90.575 137.845 90.805 138.665 ;
        RECT 90.975 137.865 91.305 138.495 ;
        RECT 90.555 137.425 90.885 137.675 ;
        RECT 91.055 137.265 91.305 137.865 ;
        RECT 91.475 137.845 91.685 138.665 ;
        RECT 92.835 137.990 93.105 138.335 ;
        RECT 93.295 138.265 93.675 138.665 ;
        RECT 93.845 138.095 94.015 138.445 ;
        RECT 94.185 138.265 94.515 138.665 ;
        RECT 94.715 138.095 94.885 138.445 ;
        RECT 95.085 138.165 95.415 138.665 ;
        RECT 95.605 138.165 95.935 138.665 ;
        RECT 87.775 136.115 90.365 137.205 ;
        RECT 90.575 136.115 90.805 137.255 ;
        RECT 90.975 136.285 91.305 137.265 ;
        RECT 92.835 137.255 93.005 137.990 ;
        RECT 93.275 137.925 94.885 138.095 ;
        RECT 96.135 138.095 96.305 138.445 ;
        RECT 96.505 138.265 96.835 138.665 ;
        RECT 97.005 138.095 97.175 138.445 ;
        RECT 97.345 138.265 97.725 138.665 ;
        RECT 93.275 137.755 93.445 137.925 ;
        RECT 93.175 137.425 93.445 137.755 ;
        RECT 93.615 137.425 94.020 137.755 ;
        RECT 93.275 137.255 93.445 137.425 ;
        RECT 91.475 136.115 91.685 137.255 ;
        RECT 92.835 136.285 93.105 137.255 ;
        RECT 93.275 137.085 94.000 137.255 ;
        RECT 94.190 137.135 94.900 137.755 ;
        RECT 95.070 137.425 95.420 137.995 ;
        RECT 95.600 137.425 95.950 137.995 ;
        RECT 96.135 137.925 97.745 138.095 ;
        RECT 97.915 137.990 98.185 138.335 ;
        RECT 97.575 137.755 97.745 137.925 ;
        RECT 93.830 136.965 94.000 137.085 ;
        RECT 95.100 136.965 95.420 137.255 ;
        RECT 93.315 136.115 93.595 136.915 ;
        RECT 93.830 136.795 95.420 136.965 ;
        RECT 95.600 136.965 95.920 137.255 ;
        RECT 96.120 137.135 96.830 137.755 ;
        RECT 97.000 137.425 97.405 137.755 ;
        RECT 97.575 137.425 97.845 137.755 ;
        RECT 97.575 137.255 97.745 137.425 ;
        RECT 98.015 137.255 98.185 137.990 ;
        RECT 98.355 137.895 100.025 138.665 ;
        RECT 100.195 137.940 100.485 138.665 ;
        RECT 97.020 137.085 97.745 137.255 ;
        RECT 97.020 136.965 97.190 137.085 ;
        RECT 95.600 136.795 97.190 136.965 ;
        RECT 93.765 136.335 95.420 136.625 ;
        RECT 95.600 136.335 97.255 136.625 ;
        RECT 97.425 136.115 97.705 136.915 ;
        RECT 97.915 136.285 98.185 137.255 ;
        RECT 98.355 137.205 99.105 137.725 ;
        RECT 99.275 137.375 100.025 137.895 ;
        RECT 100.930 137.855 101.175 138.460 ;
        RECT 101.395 138.130 101.905 138.665 ;
        RECT 100.655 137.685 101.885 137.855 ;
        RECT 98.355 136.115 100.025 137.205 ;
        RECT 100.195 136.115 100.485 137.280 ;
        RECT 100.655 136.875 100.995 137.685 ;
        RECT 101.165 137.120 101.915 137.310 ;
        RECT 100.655 136.465 101.170 136.875 ;
        RECT 101.405 136.115 101.575 136.875 ;
        RECT 101.745 136.455 101.915 137.120 ;
        RECT 102.085 137.135 102.275 138.495 ;
        RECT 102.445 138.325 102.720 138.495 ;
        RECT 102.445 138.155 102.725 138.325 ;
        RECT 102.445 137.335 102.720 138.155 ;
        RECT 102.910 138.130 103.440 138.495 ;
        RECT 103.865 138.265 104.195 138.665 ;
        RECT 103.265 138.095 103.440 138.130 ;
        RECT 102.925 137.135 103.095 137.935 ;
        RECT 102.085 136.965 103.095 137.135 ;
        RECT 103.265 137.925 104.195 138.095 ;
        RECT 104.365 137.925 104.620 138.495 ;
        RECT 105.345 138.115 105.515 138.495 ;
        RECT 105.695 138.285 106.025 138.665 ;
        RECT 105.345 137.945 106.010 138.115 ;
        RECT 106.205 137.990 106.465 138.495 ;
        RECT 106.640 138.120 111.985 138.665 ;
        RECT 103.265 136.795 103.435 137.925 ;
        RECT 104.025 137.755 104.195 137.925 ;
        RECT 102.310 136.625 103.435 136.795 ;
        RECT 103.605 137.425 103.800 137.755 ;
        RECT 104.025 137.425 104.280 137.755 ;
        RECT 103.605 136.455 103.775 137.425 ;
        RECT 104.450 137.255 104.620 137.925 ;
        RECT 105.275 137.395 105.605 137.765 ;
        RECT 105.840 137.690 106.010 137.945 ;
        RECT 101.745 136.285 103.775 136.455 ;
        RECT 103.945 136.115 104.115 137.255 ;
        RECT 104.285 136.285 104.620 137.255 ;
        RECT 105.840 137.360 106.125 137.690 ;
        RECT 105.840 137.215 106.010 137.360 ;
        RECT 105.345 137.045 106.010 137.215 ;
        RECT 106.295 137.190 106.465 137.990 ;
        RECT 105.345 136.285 105.515 137.045 ;
        RECT 105.695 136.115 106.025 136.875 ;
        RECT 106.195 136.285 106.465 137.190 ;
        RECT 108.230 136.550 108.580 137.800 ;
        RECT 110.060 137.290 110.400 138.120 ;
        RECT 112.155 137.915 113.365 138.665 ;
        RECT 112.155 137.205 112.675 137.745 ;
        RECT 112.845 137.375 113.365 137.915 ;
        RECT 106.640 136.115 111.985 136.550 ;
        RECT 112.155 136.115 113.365 137.205 ;
        RECT 15.010 135.945 113.450 136.115 ;
        RECT 15.095 134.855 16.305 135.945 ;
        RECT 15.095 134.145 15.615 134.685 ;
        RECT 15.785 134.315 16.305 134.855 ;
        RECT 16.850 134.965 17.105 135.635 ;
        RECT 17.285 135.145 17.570 135.945 ;
        RECT 17.750 135.225 18.080 135.735 ;
        RECT 15.095 133.395 16.305 134.145 ;
        RECT 16.850 134.105 17.030 134.965 ;
        RECT 17.750 134.635 18.000 135.225 ;
        RECT 18.350 135.075 18.520 135.685 ;
        RECT 18.690 135.255 19.020 135.945 ;
        RECT 19.250 135.395 19.490 135.685 ;
        RECT 19.690 135.565 20.110 135.945 ;
        RECT 20.290 135.475 20.920 135.725 ;
        RECT 21.390 135.565 21.720 135.945 ;
        RECT 20.290 135.395 20.460 135.475 ;
        RECT 21.890 135.395 22.060 135.685 ;
        RECT 22.240 135.565 22.620 135.945 ;
        RECT 22.860 135.560 23.690 135.730 ;
        RECT 19.250 135.225 20.460 135.395 ;
        RECT 17.200 134.305 18.000 134.635 ;
        RECT 16.850 133.905 17.105 134.105 ;
        RECT 16.765 133.735 17.105 133.905 ;
        RECT 16.850 133.575 17.105 133.735 ;
        RECT 17.285 133.395 17.570 133.855 ;
        RECT 17.750 133.655 18.000 134.305 ;
        RECT 18.200 135.055 18.520 135.075 ;
        RECT 18.200 134.885 20.120 135.055 ;
        RECT 18.200 133.990 18.390 134.885 ;
        RECT 20.290 134.715 20.460 135.225 ;
        RECT 20.630 134.965 21.150 135.275 ;
        RECT 18.560 134.545 20.460 134.715 ;
        RECT 18.560 134.485 18.890 134.545 ;
        RECT 19.040 134.315 19.370 134.375 ;
        RECT 18.710 134.045 19.370 134.315 ;
        RECT 18.200 133.660 18.520 133.990 ;
        RECT 18.700 133.395 19.360 133.875 ;
        RECT 19.560 133.785 19.730 134.545 ;
        RECT 20.630 134.375 20.810 134.785 ;
        RECT 19.900 134.205 20.230 134.325 ;
        RECT 20.980 134.205 21.150 134.965 ;
        RECT 19.900 134.035 21.150 134.205 ;
        RECT 21.320 135.145 22.690 135.395 ;
        RECT 21.320 134.375 21.510 135.145 ;
        RECT 22.440 134.885 22.690 135.145 ;
        RECT 21.680 134.715 21.930 134.875 ;
        RECT 22.860 134.715 23.030 135.560 ;
        RECT 23.925 135.275 24.095 135.775 ;
        RECT 24.265 135.445 24.595 135.945 ;
        RECT 23.200 134.885 23.700 135.265 ;
        RECT 23.925 135.105 24.620 135.275 ;
        RECT 21.680 134.545 23.030 134.715 ;
        RECT 22.610 134.505 23.030 134.545 ;
        RECT 21.320 134.035 21.740 134.375 ;
        RECT 22.030 134.045 22.440 134.375 ;
        RECT 19.560 133.615 20.410 133.785 ;
        RECT 20.970 133.395 21.290 133.855 ;
        RECT 21.490 133.605 21.740 134.035 ;
        RECT 22.030 133.395 22.440 133.835 ;
        RECT 22.610 133.775 22.780 134.505 ;
        RECT 22.950 133.955 23.300 134.325 ;
        RECT 23.480 134.015 23.700 134.885 ;
        RECT 23.870 134.315 24.280 134.935 ;
        RECT 24.450 134.135 24.620 135.105 ;
        RECT 23.925 133.945 24.620 134.135 ;
        RECT 22.610 133.575 23.625 133.775 ;
        RECT 23.925 133.615 24.095 133.945 ;
        RECT 24.265 133.395 24.595 133.775 ;
        RECT 24.810 133.655 25.035 135.775 ;
        RECT 25.205 135.445 25.535 135.945 ;
        RECT 25.705 135.275 25.875 135.775 ;
        RECT 25.210 135.105 25.875 135.275 ;
        RECT 25.210 134.115 25.440 135.105 ;
        RECT 26.510 134.965 26.765 135.635 ;
        RECT 26.945 135.145 27.230 135.945 ;
        RECT 27.410 135.225 27.740 135.735 ;
        RECT 25.610 134.285 25.960 134.935 ;
        RECT 25.210 133.945 25.875 134.115 ;
        RECT 25.205 133.395 25.535 133.775 ;
        RECT 25.705 133.655 25.875 133.945 ;
        RECT 26.510 134.105 26.690 134.965 ;
        RECT 27.410 134.635 27.660 135.225 ;
        RECT 28.010 135.075 28.180 135.685 ;
        RECT 28.350 135.255 28.680 135.945 ;
        RECT 28.910 135.395 29.150 135.685 ;
        RECT 29.350 135.565 29.770 135.945 ;
        RECT 29.950 135.475 30.580 135.725 ;
        RECT 31.050 135.565 31.380 135.945 ;
        RECT 29.950 135.395 30.120 135.475 ;
        RECT 31.550 135.395 31.720 135.685 ;
        RECT 31.900 135.565 32.280 135.945 ;
        RECT 32.520 135.560 33.350 135.730 ;
        RECT 28.910 135.225 30.120 135.395 ;
        RECT 26.860 134.305 27.660 134.635 ;
        RECT 26.510 133.905 26.765 134.105 ;
        RECT 26.425 133.735 26.765 133.905 ;
        RECT 26.510 133.575 26.765 133.735 ;
        RECT 26.945 133.395 27.230 133.855 ;
        RECT 27.410 133.655 27.660 134.305 ;
        RECT 27.860 135.055 28.180 135.075 ;
        RECT 27.860 134.885 29.780 135.055 ;
        RECT 27.860 133.990 28.050 134.885 ;
        RECT 29.950 134.715 30.120 135.225 ;
        RECT 30.290 134.965 30.810 135.275 ;
        RECT 28.220 134.545 30.120 134.715 ;
        RECT 28.220 134.485 28.550 134.545 ;
        RECT 28.700 134.315 29.030 134.375 ;
        RECT 28.370 134.045 29.030 134.315 ;
        RECT 27.860 133.660 28.180 133.990 ;
        RECT 28.360 133.395 29.020 133.875 ;
        RECT 29.220 133.785 29.390 134.545 ;
        RECT 30.290 134.375 30.470 134.785 ;
        RECT 29.560 134.205 29.890 134.325 ;
        RECT 30.640 134.205 30.810 134.965 ;
        RECT 29.560 134.035 30.810 134.205 ;
        RECT 30.980 135.145 32.350 135.395 ;
        RECT 30.980 134.375 31.170 135.145 ;
        RECT 32.100 134.885 32.350 135.145 ;
        RECT 31.340 134.715 31.590 134.875 ;
        RECT 32.520 134.715 32.690 135.560 ;
        RECT 33.585 135.275 33.755 135.775 ;
        RECT 33.925 135.445 34.255 135.945 ;
        RECT 32.860 134.885 33.360 135.265 ;
        RECT 33.585 135.105 34.280 135.275 ;
        RECT 31.340 134.545 32.690 134.715 ;
        RECT 32.270 134.505 32.690 134.545 ;
        RECT 30.980 134.035 31.400 134.375 ;
        RECT 31.690 134.045 32.100 134.375 ;
        RECT 29.220 133.615 30.070 133.785 ;
        RECT 30.630 133.395 30.950 133.855 ;
        RECT 31.150 133.605 31.400 134.035 ;
        RECT 31.690 133.395 32.100 133.835 ;
        RECT 32.270 133.775 32.440 134.505 ;
        RECT 32.610 133.955 32.960 134.325 ;
        RECT 33.140 134.015 33.360 134.885 ;
        RECT 33.530 134.315 33.940 134.935 ;
        RECT 34.110 134.135 34.280 135.105 ;
        RECT 33.585 133.945 34.280 134.135 ;
        RECT 32.270 133.575 33.285 133.775 ;
        RECT 33.585 133.615 33.755 133.945 ;
        RECT 33.925 133.395 34.255 133.775 ;
        RECT 34.470 133.655 34.695 135.775 ;
        RECT 34.865 135.445 35.195 135.945 ;
        RECT 35.365 135.275 35.535 135.775 ;
        RECT 34.870 135.105 35.535 135.275 ;
        RECT 34.870 134.115 35.100 135.105 ;
        RECT 35.270 134.285 35.620 134.935 ;
        RECT 35.795 134.780 36.085 135.945 ;
        RECT 36.715 134.805 36.985 135.775 ;
        RECT 37.195 135.145 37.475 135.945 ;
        RECT 37.645 135.435 39.300 135.725 ;
        RECT 37.710 135.095 39.300 135.265 ;
        RECT 37.710 134.975 37.880 135.095 ;
        RECT 37.155 134.805 37.880 134.975 ;
        RECT 34.870 133.945 35.535 134.115 ;
        RECT 34.865 133.395 35.195 133.775 ;
        RECT 35.365 133.655 35.535 133.945 ;
        RECT 35.795 133.395 36.085 134.120 ;
        RECT 36.715 134.070 36.885 134.805 ;
        RECT 37.155 134.635 37.325 134.805 ;
        RECT 37.055 134.305 37.325 134.635 ;
        RECT 37.495 134.305 37.900 134.635 ;
        RECT 38.070 134.305 38.780 134.925 ;
        RECT 38.980 134.805 39.300 135.095 ;
        RECT 39.475 134.805 39.745 135.775 ;
        RECT 39.955 135.145 40.235 135.945 ;
        RECT 40.405 135.435 42.060 135.725 ;
        RECT 40.470 135.095 42.060 135.265 ;
        RECT 40.470 134.975 40.640 135.095 ;
        RECT 39.915 134.805 40.640 134.975 ;
        RECT 37.155 134.135 37.325 134.305 ;
        RECT 36.715 133.725 36.985 134.070 ;
        RECT 37.155 133.965 38.765 134.135 ;
        RECT 38.950 134.065 39.300 134.635 ;
        RECT 39.475 134.070 39.645 134.805 ;
        RECT 39.915 134.635 40.085 134.805 ;
        RECT 39.815 134.305 40.085 134.635 ;
        RECT 40.255 134.305 40.660 134.635 ;
        RECT 40.830 134.305 41.540 134.925 ;
        RECT 41.740 134.805 42.060 135.095 ;
        RECT 42.235 134.855 43.905 135.945 ;
        RECT 39.915 134.135 40.085 134.305 ;
        RECT 37.175 133.395 37.555 133.795 ;
        RECT 37.725 133.615 37.895 133.965 ;
        RECT 38.065 133.395 38.395 133.795 ;
        RECT 38.595 133.615 38.765 133.965 ;
        RECT 38.965 133.395 39.295 133.895 ;
        RECT 39.475 133.725 39.745 134.070 ;
        RECT 39.915 133.965 41.525 134.135 ;
        RECT 41.710 134.065 42.060 134.635 ;
        RECT 42.235 134.335 42.985 134.855 ;
        RECT 44.075 134.805 44.415 135.775 ;
        RECT 44.585 134.805 44.755 135.945 ;
        RECT 45.025 135.145 45.275 135.945 ;
        RECT 45.920 134.975 46.250 135.775 ;
        RECT 46.550 135.145 46.880 135.945 ;
        RECT 47.050 134.975 47.380 135.775 ;
        RECT 44.945 134.805 47.380 134.975 ;
        RECT 47.755 134.805 48.095 135.775 ;
        RECT 48.265 134.805 48.435 135.945 ;
        RECT 48.705 135.145 48.955 135.945 ;
        RECT 49.600 134.975 49.930 135.775 ;
        RECT 50.230 135.145 50.560 135.945 ;
        RECT 50.730 134.975 51.060 135.775 ;
        RECT 48.625 134.805 51.060 134.975 ;
        RECT 51.900 134.805 52.235 135.775 ;
        RECT 52.405 134.805 52.575 135.945 ;
        RECT 52.745 135.605 54.775 135.775 ;
        RECT 43.155 134.165 43.905 134.685 ;
        RECT 39.935 133.395 40.315 133.795 ;
        RECT 40.485 133.615 40.655 133.965 ;
        RECT 40.825 133.395 41.155 133.795 ;
        RECT 41.355 133.615 41.525 133.965 ;
        RECT 41.725 133.395 42.055 133.895 ;
        RECT 42.235 133.395 43.905 134.165 ;
        RECT 44.075 134.245 44.250 134.805 ;
        RECT 44.945 134.555 45.115 134.805 ;
        RECT 44.420 134.385 45.115 134.555 ;
        RECT 45.290 134.385 45.710 134.585 ;
        RECT 45.880 134.385 46.210 134.585 ;
        RECT 46.380 134.385 46.710 134.585 ;
        RECT 44.075 134.195 44.305 134.245 ;
        RECT 44.075 133.565 44.415 134.195 ;
        RECT 44.585 133.395 44.835 134.195 ;
        RECT 45.025 134.045 46.250 134.215 ;
        RECT 45.025 133.565 45.355 134.045 ;
        RECT 45.525 133.395 45.750 133.855 ;
        RECT 45.920 133.565 46.250 134.045 ;
        RECT 46.880 134.175 47.050 134.805 ;
        RECT 47.235 134.385 47.585 134.635 ;
        RECT 47.755 134.195 47.930 134.805 ;
        RECT 48.625 134.555 48.795 134.805 ;
        RECT 48.100 134.385 48.795 134.555 ;
        RECT 48.965 134.415 49.390 134.585 ;
        RECT 48.970 134.385 49.390 134.415 ;
        RECT 49.560 134.385 49.890 134.585 ;
        RECT 50.060 134.385 50.390 134.585 ;
        RECT 46.880 133.565 47.380 134.175 ;
        RECT 47.755 133.565 48.095 134.195 ;
        RECT 48.265 133.395 48.515 134.195 ;
        RECT 48.705 134.045 49.930 134.215 ;
        RECT 48.705 133.565 49.035 134.045 ;
        RECT 49.205 133.395 49.430 133.855 ;
        RECT 49.600 133.565 49.930 134.045 ;
        RECT 50.560 134.175 50.730 134.805 ;
        RECT 50.915 134.385 51.265 134.635 ;
        RECT 50.560 133.565 51.060 134.175 ;
        RECT 51.900 134.135 52.070 134.805 ;
        RECT 52.745 134.635 52.915 135.605 ;
        RECT 52.240 134.305 52.495 134.635 ;
        RECT 52.720 134.305 52.915 134.635 ;
        RECT 53.085 135.265 54.210 135.435 ;
        RECT 52.325 134.135 52.495 134.305 ;
        RECT 53.085 134.135 53.255 135.265 ;
        RECT 51.900 133.565 52.155 134.135 ;
        RECT 52.325 133.965 53.255 134.135 ;
        RECT 53.425 134.925 54.435 135.095 ;
        RECT 53.425 134.125 53.595 134.925 ;
        RECT 53.800 134.245 54.075 134.725 ;
        RECT 53.795 134.075 54.075 134.245 ;
        RECT 53.080 133.930 53.255 133.965 ;
        RECT 52.325 133.395 52.655 133.795 ;
        RECT 53.080 133.565 53.610 133.930 ;
        RECT 53.800 133.565 54.075 134.075 ;
        RECT 54.245 133.565 54.435 134.925 ;
        RECT 54.605 134.940 54.775 135.605 ;
        RECT 54.945 135.185 55.115 135.945 ;
        RECT 55.350 135.185 55.865 135.595 ;
        RECT 54.605 134.750 55.355 134.940 ;
        RECT 55.525 134.375 55.865 135.185 ;
        RECT 56.095 134.805 56.305 135.945 ;
        RECT 54.635 134.205 55.865 134.375 ;
        RECT 56.475 134.795 56.805 135.775 ;
        RECT 56.975 134.805 57.205 135.945 ;
        RECT 57.455 134.805 57.685 135.945 ;
        RECT 57.855 134.795 58.185 135.775 ;
        RECT 58.355 134.805 58.565 135.945 ;
        RECT 58.795 134.855 61.385 135.945 ;
        RECT 54.615 133.395 55.125 133.930 ;
        RECT 55.345 133.600 55.590 134.205 ;
        RECT 56.095 133.395 56.305 134.215 ;
        RECT 56.475 134.195 56.725 134.795 ;
        RECT 56.895 134.385 57.225 134.635 ;
        RECT 57.435 134.385 57.765 134.635 ;
        RECT 56.475 133.565 56.805 134.195 ;
        RECT 56.975 133.395 57.205 134.215 ;
        RECT 57.455 133.395 57.685 134.215 ;
        RECT 57.935 134.195 58.185 134.795 ;
        RECT 58.795 134.335 60.005 134.855 ;
        RECT 61.555 134.780 61.845 135.945 ;
        RECT 62.015 134.855 63.225 135.945 ;
        RECT 63.400 135.520 63.735 135.945 ;
        RECT 63.905 135.340 64.090 135.745 ;
        RECT 63.425 135.165 64.090 135.340 ;
        RECT 64.295 135.165 64.625 135.945 ;
        RECT 57.855 133.565 58.185 134.195 ;
        RECT 58.355 133.395 58.565 134.215 ;
        RECT 60.175 134.165 61.385 134.685 ;
        RECT 62.015 134.315 62.535 134.855 ;
        RECT 58.795 133.395 61.385 134.165 ;
        RECT 62.705 134.145 63.225 134.685 ;
        RECT 61.555 133.395 61.845 134.120 ;
        RECT 62.015 133.395 63.225 134.145 ;
        RECT 63.425 134.135 63.765 135.165 ;
        RECT 64.795 134.975 65.065 135.745 ;
        RECT 63.935 134.805 65.065 134.975 ;
        RECT 63.935 134.305 64.185 134.805 ;
        RECT 63.425 133.965 64.110 134.135 ;
        RECT 64.365 134.055 64.725 134.635 ;
        RECT 63.400 133.395 63.735 133.795 ;
        RECT 63.905 133.565 64.110 133.965 ;
        RECT 64.895 133.895 65.065 134.805 ;
        RECT 65.235 134.855 67.825 135.945 ;
        RECT 68.195 135.275 68.475 135.945 ;
        RECT 68.645 135.055 68.945 135.605 ;
        RECT 69.145 135.225 69.475 135.945 ;
        RECT 69.665 135.225 70.125 135.775 ;
        RECT 65.235 134.335 66.445 134.855 ;
        RECT 66.615 134.165 67.825 134.685 ;
        RECT 68.010 134.635 68.275 134.995 ;
        RECT 68.645 134.885 69.585 135.055 ;
        RECT 69.415 134.635 69.585 134.885 ;
        RECT 68.010 134.385 68.685 134.635 ;
        RECT 68.905 134.385 69.245 134.635 ;
        RECT 69.415 134.305 69.705 134.635 ;
        RECT 69.415 134.215 69.585 134.305 ;
        RECT 64.320 133.395 64.595 133.875 ;
        RECT 64.805 133.565 65.065 133.895 ;
        RECT 65.235 133.395 67.825 134.165 ;
        RECT 68.195 134.025 69.585 134.215 ;
        RECT 68.195 133.665 68.525 134.025 ;
        RECT 69.875 133.855 70.125 135.225 ;
        RECT 70.385 135.200 70.655 135.945 ;
        RECT 71.285 135.940 77.560 135.945 ;
        RECT 70.825 135.030 71.115 135.770 ;
        RECT 71.285 135.215 71.540 135.940 ;
        RECT 71.725 135.045 71.985 135.770 ;
        RECT 72.155 135.215 72.400 135.940 ;
        RECT 72.585 135.045 72.845 135.770 ;
        RECT 73.015 135.215 73.260 135.940 ;
        RECT 73.445 135.045 73.705 135.770 ;
        RECT 73.875 135.215 74.120 135.940 ;
        RECT 74.290 135.045 74.550 135.770 ;
        RECT 74.720 135.215 74.980 135.940 ;
        RECT 75.150 135.045 75.410 135.770 ;
        RECT 75.580 135.215 75.840 135.940 ;
        RECT 76.010 135.045 76.270 135.770 ;
        RECT 76.440 135.215 76.700 135.940 ;
        RECT 76.870 135.045 77.130 135.770 ;
        RECT 77.300 135.145 77.560 135.940 ;
        RECT 71.725 135.030 77.130 135.045 ;
        RECT 70.385 134.805 77.130 135.030 ;
        RECT 70.385 134.215 71.550 134.805 ;
        RECT 77.730 134.635 77.980 135.770 ;
        RECT 78.160 135.135 78.420 135.945 ;
        RECT 78.595 134.635 78.840 135.775 ;
        RECT 79.020 135.135 79.315 135.945 ;
        RECT 79.555 134.805 79.765 135.945 ;
        RECT 79.935 134.795 80.265 135.775 ;
        RECT 80.435 134.805 80.665 135.945 ;
        RECT 80.965 135.015 81.135 135.775 ;
        RECT 81.315 135.185 81.645 135.945 ;
        RECT 80.965 134.845 81.630 135.015 ;
        RECT 81.815 134.870 82.085 135.775 ;
        RECT 71.720 134.385 78.840 134.635 ;
        RECT 70.385 134.045 77.130 134.215 ;
        RECT 69.145 133.395 69.395 133.855 ;
        RECT 69.565 133.565 70.125 133.855 ;
        RECT 70.385 133.395 70.685 133.875 ;
        RECT 70.855 133.590 71.115 134.045 ;
        RECT 71.285 133.395 71.545 133.875 ;
        RECT 71.725 133.590 71.985 134.045 ;
        RECT 72.155 133.395 72.405 133.875 ;
        RECT 72.585 133.590 72.845 134.045 ;
        RECT 73.015 133.395 73.265 133.875 ;
        RECT 73.445 133.590 73.705 134.045 ;
        RECT 73.875 133.395 74.120 133.875 ;
        RECT 74.290 133.590 74.565 134.045 ;
        RECT 74.735 133.395 74.980 133.875 ;
        RECT 75.150 133.590 75.410 134.045 ;
        RECT 75.580 133.395 75.840 133.875 ;
        RECT 76.010 133.590 76.270 134.045 ;
        RECT 76.440 133.395 76.700 133.875 ;
        RECT 76.870 133.590 77.130 134.045 ;
        RECT 77.300 133.395 77.560 133.955 ;
        RECT 77.730 133.575 77.980 134.385 ;
        RECT 78.160 133.395 78.420 133.920 ;
        RECT 78.590 133.575 78.840 134.385 ;
        RECT 79.010 134.075 79.325 134.635 ;
        RECT 79.020 133.395 79.325 133.905 ;
        RECT 79.555 133.395 79.765 134.215 ;
        RECT 79.935 134.195 80.185 134.795 ;
        RECT 81.460 134.700 81.630 134.845 ;
        RECT 80.355 134.385 80.685 134.635 ;
        RECT 80.895 134.295 81.225 134.665 ;
        RECT 81.460 134.370 81.745 134.700 ;
        RECT 79.935 133.565 80.265 134.195 ;
        RECT 80.435 133.395 80.665 134.215 ;
        RECT 81.460 134.115 81.630 134.370 ;
        RECT 80.965 133.945 81.630 134.115 ;
        RECT 81.915 134.070 82.085 134.870 ;
        RECT 82.255 134.855 83.465 135.945 ;
        RECT 83.635 134.855 87.145 135.945 ;
        RECT 82.255 134.315 82.775 134.855 ;
        RECT 82.945 134.145 83.465 134.685 ;
        RECT 83.635 134.335 85.325 134.855 ;
        RECT 87.315 134.780 87.605 135.945 ;
        RECT 87.785 135.135 88.080 135.945 ;
        RECT 85.495 134.165 87.145 134.685 ;
        RECT 88.260 134.635 88.505 135.775 ;
        RECT 88.680 135.135 88.940 135.945 ;
        RECT 89.540 135.940 95.815 135.945 ;
        RECT 89.120 134.635 89.370 135.770 ;
        RECT 89.540 135.145 89.800 135.940 ;
        RECT 89.970 135.045 90.230 135.770 ;
        RECT 90.400 135.215 90.660 135.940 ;
        RECT 90.830 135.045 91.090 135.770 ;
        RECT 91.260 135.215 91.520 135.940 ;
        RECT 91.690 135.045 91.950 135.770 ;
        RECT 92.120 135.215 92.380 135.940 ;
        RECT 92.550 135.045 92.810 135.770 ;
        RECT 92.980 135.215 93.225 135.940 ;
        RECT 93.395 135.045 93.655 135.770 ;
        RECT 93.840 135.215 94.085 135.940 ;
        RECT 94.255 135.045 94.515 135.770 ;
        RECT 94.700 135.215 94.945 135.940 ;
        RECT 95.115 135.045 95.375 135.770 ;
        RECT 95.560 135.215 95.815 135.940 ;
        RECT 89.970 135.030 95.375 135.045 ;
        RECT 95.985 135.030 96.275 135.770 ;
        RECT 96.445 135.200 96.715 135.945 ;
        RECT 97.895 135.225 98.355 135.775 ;
        RECT 98.545 135.225 98.875 135.945 ;
        RECT 89.970 134.805 96.715 135.030 ;
        RECT 80.965 133.565 81.135 133.945 ;
        RECT 81.315 133.395 81.645 133.775 ;
        RECT 81.825 133.565 82.085 134.070 ;
        RECT 82.255 133.395 83.465 134.145 ;
        RECT 83.635 133.395 87.145 134.165 ;
        RECT 87.315 133.395 87.605 134.120 ;
        RECT 87.775 134.075 88.090 134.635 ;
        RECT 88.260 134.385 95.380 134.635 ;
        RECT 87.775 133.395 88.080 133.905 ;
        RECT 88.260 133.575 88.510 134.385 ;
        RECT 88.680 133.395 88.940 133.920 ;
        RECT 89.120 133.575 89.370 134.385 ;
        RECT 95.550 134.215 96.715 134.805 ;
        RECT 89.970 134.045 96.715 134.215 ;
        RECT 89.540 133.395 89.800 133.955 ;
        RECT 89.970 133.590 90.230 134.045 ;
        RECT 90.400 133.395 90.660 133.875 ;
        RECT 90.830 133.590 91.090 134.045 ;
        RECT 91.260 133.395 91.520 133.875 ;
        RECT 91.690 133.590 91.950 134.045 ;
        RECT 92.120 133.395 92.365 133.875 ;
        RECT 92.535 133.590 92.810 134.045 ;
        RECT 92.980 133.395 93.225 133.875 ;
        RECT 93.395 133.590 93.655 134.045 ;
        RECT 93.835 133.395 94.085 133.875 ;
        RECT 94.255 133.590 94.515 134.045 ;
        RECT 94.695 133.395 94.945 133.875 ;
        RECT 95.115 133.590 95.375 134.045 ;
        RECT 95.555 133.395 95.815 133.875 ;
        RECT 95.985 133.590 96.245 134.045 ;
        RECT 96.415 133.395 96.715 133.875 ;
        RECT 97.895 133.855 98.145 135.225 ;
        RECT 99.075 135.055 99.375 135.605 ;
        RECT 99.545 135.275 99.825 135.945 ;
        RECT 101.120 135.510 106.465 135.945 ;
        RECT 106.640 135.510 111.985 135.945 ;
        RECT 98.435 134.885 99.375 135.055 ;
        RECT 98.435 134.635 98.605 134.885 ;
        RECT 99.745 134.635 100.010 134.995 ;
        RECT 98.315 134.305 98.605 134.635 ;
        RECT 98.775 134.385 99.115 134.635 ;
        RECT 99.335 134.385 100.010 134.635 ;
        RECT 98.435 134.215 98.605 134.305 ;
        RECT 102.710 134.260 103.060 135.510 ;
        RECT 98.435 134.025 99.825 134.215 ;
        RECT 97.895 133.565 98.455 133.855 ;
        RECT 98.625 133.395 98.875 133.855 ;
        RECT 99.495 133.665 99.825 134.025 ;
        RECT 104.540 133.940 104.880 134.770 ;
        RECT 108.230 134.260 108.580 135.510 ;
        RECT 112.155 134.855 113.365 135.945 ;
        RECT 110.060 133.940 110.400 134.770 ;
        RECT 112.155 134.315 112.675 134.855 ;
        RECT 112.845 134.145 113.365 134.685 ;
        RECT 101.120 133.395 106.465 133.940 ;
        RECT 106.640 133.395 111.985 133.940 ;
        RECT 112.155 133.395 113.365 134.145 ;
        RECT 15.010 133.225 113.450 133.395 ;
        RECT 15.095 132.475 16.305 133.225 ;
        RECT 15.095 131.935 15.615 132.475 ;
        RECT 16.935 132.455 18.605 133.225 ;
        RECT 15.785 131.765 16.305 132.305 ;
        RECT 15.095 130.675 16.305 131.765 ;
        RECT 16.935 131.765 17.685 132.285 ;
        RECT 17.855 131.935 18.605 132.455 ;
        RECT 19.050 132.415 19.295 133.020 ;
        RECT 19.515 132.690 20.025 133.225 ;
        RECT 18.775 132.245 20.005 132.415 ;
        RECT 16.935 130.675 18.605 131.765 ;
        RECT 18.775 131.435 19.115 132.245 ;
        RECT 19.285 131.680 20.035 131.870 ;
        RECT 18.775 131.025 19.290 131.435 ;
        RECT 19.525 130.675 19.695 131.435 ;
        RECT 19.865 131.015 20.035 131.680 ;
        RECT 20.205 131.695 20.395 133.055 ;
        RECT 20.565 132.205 20.840 133.055 ;
        RECT 21.030 132.690 21.560 133.055 ;
        RECT 21.985 132.825 22.315 133.225 ;
        RECT 21.385 132.655 21.560 132.690 ;
        RECT 20.565 132.035 20.845 132.205 ;
        RECT 20.565 131.895 20.840 132.035 ;
        RECT 21.045 131.695 21.215 132.495 ;
        RECT 20.205 131.525 21.215 131.695 ;
        RECT 21.385 132.485 22.315 132.655 ;
        RECT 22.485 132.485 22.740 133.055 ;
        RECT 22.915 132.500 23.205 133.225 ;
        RECT 23.465 132.675 23.635 132.965 ;
        RECT 23.805 132.845 24.135 133.225 ;
        RECT 23.465 132.505 24.130 132.675 ;
        RECT 21.385 131.355 21.555 132.485 ;
        RECT 22.145 132.315 22.315 132.485 ;
        RECT 20.430 131.185 21.555 131.355 ;
        RECT 21.725 131.985 21.920 132.315 ;
        RECT 22.145 131.985 22.400 132.315 ;
        RECT 21.725 131.015 21.895 131.985 ;
        RECT 22.570 131.815 22.740 132.485 ;
        RECT 19.865 130.845 21.895 131.015 ;
        RECT 22.065 130.675 22.235 131.815 ;
        RECT 22.405 130.845 22.740 131.815 ;
        RECT 22.915 130.675 23.205 131.840 ;
        RECT 23.380 131.685 23.730 132.335 ;
        RECT 23.900 131.515 24.130 132.505 ;
        RECT 23.465 131.345 24.130 131.515 ;
        RECT 23.465 130.845 23.635 131.345 ;
        RECT 23.805 130.675 24.135 131.175 ;
        RECT 24.305 130.845 24.530 132.965 ;
        RECT 24.745 132.845 25.075 133.225 ;
        RECT 25.245 132.675 25.415 133.005 ;
        RECT 25.715 132.845 26.730 133.045 ;
        RECT 24.720 132.485 25.415 132.675 ;
        RECT 24.720 131.515 24.890 132.485 ;
        RECT 25.060 131.685 25.470 132.305 ;
        RECT 25.640 131.735 25.860 132.605 ;
        RECT 26.040 132.295 26.390 132.665 ;
        RECT 26.560 132.115 26.730 132.845 ;
        RECT 26.900 132.785 27.310 133.225 ;
        RECT 27.600 132.585 27.850 133.015 ;
        RECT 28.050 132.765 28.370 133.225 ;
        RECT 28.930 132.835 29.780 133.005 ;
        RECT 26.900 132.245 27.310 132.575 ;
        RECT 27.600 132.245 28.020 132.585 ;
        RECT 26.310 132.075 26.730 132.115 ;
        RECT 26.310 131.905 27.660 132.075 ;
        RECT 24.720 131.345 25.415 131.515 ;
        RECT 25.640 131.355 26.140 131.735 ;
        RECT 24.745 130.675 25.075 131.175 ;
        RECT 25.245 130.845 25.415 131.345 ;
        RECT 26.310 131.060 26.480 131.905 ;
        RECT 27.410 131.745 27.660 131.905 ;
        RECT 26.650 131.475 26.900 131.735 ;
        RECT 27.830 131.475 28.020 132.245 ;
        RECT 26.650 131.225 28.020 131.475 ;
        RECT 28.190 132.415 29.440 132.585 ;
        RECT 28.190 131.655 28.360 132.415 ;
        RECT 29.110 132.295 29.440 132.415 ;
        RECT 28.530 131.835 28.710 132.245 ;
        RECT 29.610 132.075 29.780 132.835 ;
        RECT 29.980 132.745 30.640 133.225 ;
        RECT 30.820 132.630 31.140 132.960 ;
        RECT 29.970 132.305 30.630 132.575 ;
        RECT 29.970 132.245 30.300 132.305 ;
        RECT 30.450 132.075 30.780 132.135 ;
        RECT 28.880 131.905 30.780 132.075 ;
        RECT 28.190 131.345 28.710 131.655 ;
        RECT 28.880 131.395 29.050 131.905 ;
        RECT 30.950 131.735 31.140 132.630 ;
        RECT 29.220 131.565 31.140 131.735 ;
        RECT 30.820 131.545 31.140 131.565 ;
        RECT 31.340 132.315 31.590 132.965 ;
        RECT 31.770 132.765 32.055 133.225 ;
        RECT 32.235 132.515 32.490 133.045 ;
        RECT 33.125 132.745 33.425 133.225 ;
        RECT 33.595 132.575 33.855 133.030 ;
        RECT 34.025 132.745 34.285 133.225 ;
        RECT 34.465 132.575 34.725 133.030 ;
        RECT 34.895 132.745 35.145 133.225 ;
        RECT 35.325 132.575 35.585 133.030 ;
        RECT 35.755 132.745 36.005 133.225 ;
        RECT 36.185 132.575 36.445 133.030 ;
        RECT 36.615 132.745 36.860 133.225 ;
        RECT 37.030 132.575 37.305 133.030 ;
        RECT 37.475 132.745 37.720 133.225 ;
        RECT 37.890 132.575 38.150 133.030 ;
        RECT 38.320 132.745 38.580 133.225 ;
        RECT 38.750 132.575 39.010 133.030 ;
        RECT 39.180 132.745 39.440 133.225 ;
        RECT 39.610 132.575 39.870 133.030 ;
        RECT 40.040 132.665 40.300 133.225 ;
        RECT 31.340 131.985 32.140 132.315 ;
        RECT 28.880 131.225 30.090 131.395 ;
        RECT 25.650 130.890 26.480 131.060 ;
        RECT 26.720 130.675 27.100 131.055 ;
        RECT 27.280 130.935 27.450 131.225 ;
        RECT 28.880 131.145 29.050 131.225 ;
        RECT 27.620 130.675 27.950 131.055 ;
        RECT 28.420 130.895 29.050 131.145 ;
        RECT 29.230 130.675 29.650 131.055 ;
        RECT 29.850 130.935 30.090 131.225 ;
        RECT 30.320 130.675 30.650 131.365 ;
        RECT 30.820 130.935 30.990 131.545 ;
        RECT 31.340 131.395 31.590 131.985 ;
        RECT 32.310 131.655 32.490 132.515 ;
        RECT 33.125 132.405 39.870 132.575 ;
        RECT 33.125 132.205 34.290 132.405 ;
        RECT 40.470 132.235 40.720 133.045 ;
        RECT 40.900 132.700 41.160 133.225 ;
        RECT 41.330 132.235 41.580 133.045 ;
        RECT 41.760 132.715 42.065 133.225 ;
        RECT 42.435 132.595 42.765 132.955 ;
        RECT 43.385 132.765 43.635 133.225 ;
        RECT 43.805 132.765 44.365 133.055 ;
        RECT 33.095 132.035 34.290 132.205 ;
        RECT 31.260 130.885 31.590 131.395 ;
        RECT 31.770 130.675 32.055 131.475 ;
        RECT 32.235 131.185 32.490 131.655 ;
        RECT 33.125 131.815 34.290 132.035 ;
        RECT 34.460 131.985 41.580 132.235 ;
        RECT 41.750 131.985 42.065 132.545 ;
        RECT 42.435 132.405 43.825 132.595 ;
        RECT 43.655 132.315 43.825 132.405 ;
        RECT 42.250 131.985 42.925 132.235 ;
        RECT 43.145 131.985 43.485 132.235 ;
        RECT 43.655 131.985 43.945 132.315 ;
        RECT 33.125 131.590 39.870 131.815 ;
        RECT 32.235 131.015 32.575 131.185 ;
        RECT 32.235 130.985 32.490 131.015 ;
        RECT 33.125 130.675 33.395 131.420 ;
        RECT 33.565 130.850 33.855 131.590 ;
        RECT 34.465 131.575 39.870 131.590 ;
        RECT 34.025 130.680 34.280 131.405 ;
        RECT 34.465 130.850 34.725 131.575 ;
        RECT 34.895 130.680 35.140 131.405 ;
        RECT 35.325 130.850 35.585 131.575 ;
        RECT 35.755 130.680 36.000 131.405 ;
        RECT 36.185 130.850 36.445 131.575 ;
        RECT 36.615 130.680 36.860 131.405 ;
        RECT 37.030 130.850 37.290 131.575 ;
        RECT 37.460 130.680 37.720 131.405 ;
        RECT 37.890 130.850 38.150 131.575 ;
        RECT 38.320 130.680 38.580 131.405 ;
        RECT 38.750 130.850 39.010 131.575 ;
        RECT 39.180 130.680 39.440 131.405 ;
        RECT 39.610 130.850 39.870 131.575 ;
        RECT 40.040 130.680 40.300 131.475 ;
        RECT 40.470 130.850 40.720 131.985 ;
        RECT 34.025 130.675 40.300 130.680 ;
        RECT 40.900 130.675 41.160 131.485 ;
        RECT 41.335 130.845 41.580 131.985 ;
        RECT 42.250 131.625 42.515 131.985 ;
        RECT 43.655 131.735 43.825 131.985 ;
        RECT 42.885 131.565 43.825 131.735 ;
        RECT 41.760 130.675 42.055 131.485 ;
        RECT 42.435 130.675 42.715 131.345 ;
        RECT 42.885 131.015 43.185 131.565 ;
        RECT 44.115 131.395 44.365 132.765 ;
        RECT 43.385 130.675 43.715 131.395 ;
        RECT 43.905 130.845 44.365 131.395 ;
        RECT 44.535 132.765 45.095 133.055 ;
        RECT 45.265 132.765 45.515 133.225 ;
        RECT 44.535 131.395 44.785 132.765 ;
        RECT 46.135 132.595 46.465 132.955 ;
        RECT 45.075 132.405 46.465 132.595 ;
        RECT 46.835 132.455 48.505 133.225 ;
        RECT 48.675 132.500 48.965 133.225 ;
        RECT 49.225 132.675 49.395 133.055 ;
        RECT 49.575 132.845 49.905 133.225 ;
        RECT 49.225 132.505 49.890 132.675 ;
        RECT 50.085 132.550 50.345 133.055 ;
        RECT 45.075 132.315 45.245 132.405 ;
        RECT 44.955 131.985 45.245 132.315 ;
        RECT 45.415 131.985 45.755 132.235 ;
        RECT 45.975 131.985 46.650 132.235 ;
        RECT 45.075 131.735 45.245 131.985 ;
        RECT 45.075 131.565 46.015 131.735 ;
        RECT 46.385 131.625 46.650 131.985 ;
        RECT 46.835 131.765 47.585 132.285 ;
        RECT 47.755 131.935 48.505 132.455 ;
        RECT 49.155 131.955 49.485 132.325 ;
        RECT 49.720 132.250 49.890 132.505 ;
        RECT 49.720 131.920 50.005 132.250 ;
        RECT 44.535 130.845 44.995 131.395 ;
        RECT 45.185 130.675 45.515 131.395 ;
        RECT 45.715 131.015 46.015 131.565 ;
        RECT 46.185 130.675 46.465 131.345 ;
        RECT 46.835 130.675 48.505 131.765 ;
        RECT 48.675 130.675 48.965 131.840 ;
        RECT 49.720 131.775 49.890 131.920 ;
        RECT 49.225 131.605 49.890 131.775 ;
        RECT 50.175 131.750 50.345 132.550 ;
        RECT 50.605 132.675 50.775 132.965 ;
        RECT 50.945 132.845 51.275 133.225 ;
        RECT 50.605 132.505 51.270 132.675 ;
        RECT 49.225 130.845 49.395 131.605 ;
        RECT 49.575 130.675 49.905 131.435 ;
        RECT 50.075 130.845 50.345 131.750 ;
        RECT 50.520 131.685 50.870 132.335 ;
        RECT 51.040 131.515 51.270 132.505 ;
        RECT 50.605 131.345 51.270 131.515 ;
        RECT 50.605 130.845 50.775 131.345 ;
        RECT 50.945 130.675 51.275 131.175 ;
        RECT 51.445 130.845 51.670 132.965 ;
        RECT 51.885 132.845 52.215 133.225 ;
        RECT 52.385 132.675 52.555 133.005 ;
        RECT 52.855 132.845 53.870 133.045 ;
        RECT 51.860 132.485 52.555 132.675 ;
        RECT 51.860 131.515 52.030 132.485 ;
        RECT 52.200 131.685 52.610 132.305 ;
        RECT 52.780 131.735 53.000 132.605 ;
        RECT 53.180 132.295 53.530 132.665 ;
        RECT 53.700 132.115 53.870 132.845 ;
        RECT 54.040 132.785 54.450 133.225 ;
        RECT 54.740 132.585 54.990 133.015 ;
        RECT 55.190 132.765 55.510 133.225 ;
        RECT 56.070 132.835 56.920 133.005 ;
        RECT 54.040 132.245 54.450 132.575 ;
        RECT 54.740 132.245 55.160 132.585 ;
        RECT 53.450 132.075 53.870 132.115 ;
        RECT 53.450 131.905 54.800 132.075 ;
        RECT 51.860 131.345 52.555 131.515 ;
        RECT 52.780 131.355 53.280 131.735 ;
        RECT 51.885 130.675 52.215 131.175 ;
        RECT 52.385 130.845 52.555 131.345 ;
        RECT 53.450 131.060 53.620 131.905 ;
        RECT 54.550 131.745 54.800 131.905 ;
        RECT 53.790 131.475 54.040 131.735 ;
        RECT 54.970 131.475 55.160 132.245 ;
        RECT 53.790 131.225 55.160 131.475 ;
        RECT 55.330 132.415 56.580 132.585 ;
        RECT 55.330 131.655 55.500 132.415 ;
        RECT 56.250 132.295 56.580 132.415 ;
        RECT 55.670 131.835 55.850 132.245 ;
        RECT 56.750 132.075 56.920 132.835 ;
        RECT 57.120 132.745 57.780 133.225 ;
        RECT 57.960 132.630 58.280 132.960 ;
        RECT 57.110 132.305 57.770 132.575 ;
        RECT 57.110 132.245 57.440 132.305 ;
        RECT 57.590 132.075 57.920 132.135 ;
        RECT 56.020 131.905 57.920 132.075 ;
        RECT 55.330 131.345 55.850 131.655 ;
        RECT 56.020 131.395 56.190 131.905 ;
        RECT 58.090 131.735 58.280 132.630 ;
        RECT 56.360 131.565 58.280 131.735 ;
        RECT 57.960 131.545 58.280 131.565 ;
        RECT 58.480 132.315 58.730 132.965 ;
        RECT 58.910 132.765 59.195 133.225 ;
        RECT 59.375 132.515 59.630 133.045 ;
        RECT 60.235 132.745 60.515 133.225 ;
        RECT 60.685 132.575 60.945 132.965 ;
        RECT 61.120 132.745 61.375 133.225 ;
        RECT 61.545 132.575 61.840 132.965 ;
        RECT 62.020 132.745 62.295 133.225 ;
        RECT 62.465 132.725 62.765 133.055 ;
        RECT 58.480 131.985 59.280 132.315 ;
        RECT 56.020 131.225 57.230 131.395 ;
        RECT 52.790 130.890 53.620 131.060 ;
        RECT 53.860 130.675 54.240 131.055 ;
        RECT 54.420 130.935 54.590 131.225 ;
        RECT 56.020 131.145 56.190 131.225 ;
        RECT 54.760 130.675 55.090 131.055 ;
        RECT 55.560 130.895 56.190 131.145 ;
        RECT 56.370 130.675 56.790 131.055 ;
        RECT 56.990 130.935 57.230 131.225 ;
        RECT 57.460 130.675 57.790 131.365 ;
        RECT 57.960 130.935 58.130 131.545 ;
        RECT 58.480 131.395 58.730 131.985 ;
        RECT 59.450 131.655 59.630 132.515 ;
        RECT 60.190 132.405 61.840 132.575 ;
        RECT 60.190 131.895 60.595 132.405 ;
        RECT 60.765 132.065 61.905 132.235 ;
        RECT 60.190 131.725 60.945 131.895 ;
        RECT 58.400 130.885 58.730 131.395 ;
        RECT 58.910 130.675 59.195 131.475 ;
        RECT 59.375 131.185 59.630 131.655 ;
        RECT 59.375 131.015 59.715 131.185 ;
        RECT 59.375 130.985 59.630 131.015 ;
        RECT 60.230 130.675 60.515 131.545 ;
        RECT 60.685 131.475 60.945 131.725 ;
        RECT 61.735 131.815 61.905 132.065 ;
        RECT 62.075 131.985 62.425 132.555 ;
        RECT 62.595 131.815 62.765 132.725 ;
        RECT 62.935 132.475 64.145 133.225 ;
        RECT 61.735 131.645 62.765 131.815 ;
        RECT 60.685 131.305 61.805 131.475 ;
        RECT 60.685 130.845 60.945 131.305 ;
        RECT 61.120 130.675 61.375 131.135 ;
        RECT 61.545 130.845 61.805 131.305 ;
        RECT 61.975 130.675 62.285 131.475 ;
        RECT 62.455 130.845 62.765 131.645 ;
        RECT 62.935 131.765 63.455 132.305 ;
        RECT 63.625 131.935 64.145 132.475 ;
        RECT 64.315 132.765 64.875 133.055 ;
        RECT 65.045 132.765 65.295 133.225 ;
        RECT 62.935 130.675 64.145 131.765 ;
        RECT 64.315 131.395 64.565 132.765 ;
        RECT 65.915 132.595 66.245 132.955 ;
        RECT 64.855 132.405 66.245 132.595 ;
        RECT 67.535 132.765 68.095 133.055 ;
        RECT 68.265 132.765 68.515 133.225 ;
        RECT 64.855 132.315 65.025 132.405 ;
        RECT 64.735 131.985 65.025 132.315 ;
        RECT 65.195 131.985 65.535 132.235 ;
        RECT 65.755 131.985 66.430 132.235 ;
        RECT 64.855 131.735 65.025 131.985 ;
        RECT 64.855 131.565 65.795 131.735 ;
        RECT 66.165 131.625 66.430 131.985 ;
        RECT 64.315 130.845 64.775 131.395 ;
        RECT 64.965 130.675 65.295 131.395 ;
        RECT 65.495 131.015 65.795 131.565 ;
        RECT 67.535 131.395 67.785 132.765 ;
        RECT 69.135 132.595 69.465 132.955 ;
        RECT 68.075 132.405 69.465 132.595 ;
        RECT 70.755 132.425 71.095 133.055 ;
        RECT 71.265 132.425 71.515 133.225 ;
        RECT 71.705 132.575 72.035 133.055 ;
        RECT 72.205 132.765 72.430 133.225 ;
        RECT 72.600 132.575 72.930 133.055 ;
        RECT 68.075 132.315 68.245 132.405 ;
        RECT 67.955 131.985 68.245 132.315 ;
        RECT 68.415 131.985 68.755 132.235 ;
        RECT 68.975 131.985 69.650 132.235 ;
        RECT 68.075 131.735 68.245 131.985 ;
        RECT 68.075 131.565 69.015 131.735 ;
        RECT 69.385 131.625 69.650 131.985 ;
        RECT 70.755 131.815 70.930 132.425 ;
        RECT 71.705 132.405 72.930 132.575 ;
        RECT 73.560 132.445 74.060 133.055 ;
        RECT 74.435 132.500 74.725 133.225 ;
        RECT 74.895 132.550 75.155 133.055 ;
        RECT 75.335 132.845 75.665 133.225 ;
        RECT 75.845 132.675 76.015 133.055 ;
        RECT 76.375 132.760 76.625 133.225 ;
        RECT 71.100 132.065 71.795 132.235 ;
        RECT 71.625 131.815 71.795 132.065 ;
        RECT 71.970 132.035 72.390 132.235 ;
        RECT 72.560 132.035 72.890 132.235 ;
        RECT 73.060 132.035 73.390 132.235 ;
        RECT 73.560 131.815 73.730 132.445 ;
        RECT 73.915 131.985 74.265 132.235 ;
        RECT 65.965 130.675 66.245 131.345 ;
        RECT 67.535 130.845 67.995 131.395 ;
        RECT 68.185 130.675 68.515 131.395 ;
        RECT 68.715 131.015 69.015 131.565 ;
        RECT 69.185 130.675 69.465 131.345 ;
        RECT 70.755 130.845 71.095 131.815 ;
        RECT 71.265 130.675 71.435 131.815 ;
        RECT 71.625 131.645 74.060 131.815 ;
        RECT 71.705 130.675 71.955 131.475 ;
        RECT 72.600 130.845 72.930 131.645 ;
        RECT 73.230 130.675 73.560 131.475 ;
        RECT 73.730 130.845 74.060 131.645 ;
        RECT 74.435 130.675 74.725 131.840 ;
        RECT 74.895 131.750 75.065 132.550 ;
        RECT 75.350 132.505 76.015 132.675 ;
        RECT 76.795 132.585 76.965 133.055 ;
        RECT 77.215 132.765 77.385 133.225 ;
        RECT 77.635 132.585 77.805 133.055 ;
        RECT 78.055 132.765 78.225 133.225 ;
        RECT 78.475 132.585 78.645 133.055 ;
        RECT 79.015 132.765 79.280 133.225 ;
        RECT 79.495 132.765 80.055 133.055 ;
        RECT 80.225 132.765 80.475 133.225 ;
        RECT 75.350 132.250 75.520 132.505 ;
        RECT 76.275 132.405 78.645 132.585 ;
        RECT 75.235 131.920 75.520 132.250 ;
        RECT 75.755 131.955 76.085 132.325 ;
        RECT 75.350 131.775 75.520 131.920 ;
        RECT 76.275 131.815 76.625 132.405 ;
        RECT 76.795 131.985 79.305 132.235 ;
        RECT 74.895 130.845 75.165 131.750 ;
        RECT 75.350 131.605 76.015 131.775 ;
        RECT 76.275 131.645 78.725 131.815 ;
        RECT 76.275 131.625 77.045 131.645 ;
        RECT 75.335 130.675 75.665 131.435 ;
        RECT 75.845 130.845 76.015 131.605 ;
        RECT 76.375 130.675 76.545 131.135 ;
        RECT 76.715 130.845 77.045 131.625 ;
        RECT 77.215 130.675 77.385 131.475 ;
        RECT 77.555 130.845 77.885 131.645 ;
        RECT 78.055 130.675 78.225 131.475 ;
        RECT 78.395 130.845 78.725 131.645 ;
        RECT 78.985 130.675 79.280 131.815 ;
        RECT 79.495 131.395 79.745 132.765 ;
        RECT 81.095 132.595 81.425 132.955 ;
        RECT 80.035 132.405 81.425 132.595 ;
        RECT 81.795 132.455 83.465 133.225 ;
        RECT 80.035 132.315 80.205 132.405 ;
        RECT 79.915 131.985 80.205 132.315 ;
        RECT 80.375 131.985 80.715 132.235 ;
        RECT 80.935 131.985 81.610 132.235 ;
        RECT 80.035 131.735 80.205 131.985 ;
        RECT 80.035 131.565 80.975 131.735 ;
        RECT 81.345 131.625 81.610 131.985 ;
        RECT 81.795 131.765 82.545 132.285 ;
        RECT 82.715 131.935 83.465 132.455 ;
        RECT 84.010 132.515 84.265 133.045 ;
        RECT 84.445 132.765 84.730 133.225 ;
        RECT 79.495 130.845 79.955 131.395 ;
        RECT 80.145 130.675 80.475 131.395 ;
        RECT 80.675 131.015 80.975 131.565 ;
        RECT 81.145 130.675 81.425 131.345 ;
        RECT 81.795 130.675 83.465 131.765 ;
        RECT 84.010 131.655 84.190 132.515 ;
        RECT 84.910 132.315 85.160 132.965 ;
        RECT 84.360 131.985 85.160 132.315 ;
        RECT 84.010 131.185 84.265 131.655 ;
        RECT 83.925 131.015 84.265 131.185 ;
        RECT 84.010 130.985 84.265 131.015 ;
        RECT 84.445 130.675 84.730 131.475 ;
        RECT 84.910 131.395 85.160 131.985 ;
        RECT 85.360 132.630 85.680 132.960 ;
        RECT 85.860 132.745 86.520 133.225 ;
        RECT 86.720 132.835 87.570 133.005 ;
        RECT 85.360 131.735 85.550 132.630 ;
        RECT 85.870 132.305 86.530 132.575 ;
        RECT 86.200 132.245 86.530 132.305 ;
        RECT 85.720 132.075 86.050 132.135 ;
        RECT 86.720 132.075 86.890 132.835 ;
        RECT 88.130 132.765 88.450 133.225 ;
        RECT 88.650 132.585 88.900 133.015 ;
        RECT 89.190 132.785 89.600 133.225 ;
        RECT 89.770 132.845 90.785 133.045 ;
        RECT 87.060 132.415 88.310 132.585 ;
        RECT 87.060 132.295 87.390 132.415 ;
        RECT 85.720 131.905 87.620 132.075 ;
        RECT 85.360 131.565 87.280 131.735 ;
        RECT 85.360 131.545 85.680 131.565 ;
        RECT 84.910 130.885 85.240 131.395 ;
        RECT 85.510 130.935 85.680 131.545 ;
        RECT 87.450 131.395 87.620 131.905 ;
        RECT 87.790 131.835 87.970 132.245 ;
        RECT 88.140 131.655 88.310 132.415 ;
        RECT 85.850 130.675 86.180 131.365 ;
        RECT 86.410 131.225 87.620 131.395 ;
        RECT 87.790 131.345 88.310 131.655 ;
        RECT 88.480 132.245 88.900 132.585 ;
        RECT 89.190 132.245 89.600 132.575 ;
        RECT 88.480 131.475 88.670 132.245 ;
        RECT 89.770 132.115 89.940 132.845 ;
        RECT 91.085 132.675 91.255 133.005 ;
        RECT 91.425 132.845 91.755 133.225 ;
        RECT 90.110 132.295 90.460 132.665 ;
        RECT 89.770 132.075 90.190 132.115 ;
        RECT 88.840 131.905 90.190 132.075 ;
        RECT 88.840 131.745 89.090 131.905 ;
        RECT 89.600 131.475 89.850 131.735 ;
        RECT 88.480 131.225 89.850 131.475 ;
        RECT 86.410 130.935 86.650 131.225 ;
        RECT 87.450 131.145 87.620 131.225 ;
        RECT 86.850 130.675 87.270 131.055 ;
        RECT 87.450 130.895 88.080 131.145 ;
        RECT 88.550 130.675 88.880 131.055 ;
        RECT 89.050 130.935 89.220 131.225 ;
        RECT 90.020 131.060 90.190 131.905 ;
        RECT 90.640 131.735 90.860 132.605 ;
        RECT 91.085 132.485 91.780 132.675 ;
        RECT 90.360 131.355 90.860 131.735 ;
        RECT 91.030 131.685 91.440 132.305 ;
        RECT 91.610 131.515 91.780 132.485 ;
        RECT 91.085 131.345 91.780 131.515 ;
        RECT 89.400 130.675 89.780 131.055 ;
        RECT 90.020 130.890 90.850 131.060 ;
        RECT 91.085 130.845 91.255 131.345 ;
        RECT 91.425 130.675 91.755 131.175 ;
        RECT 91.970 130.845 92.195 132.965 ;
        RECT 92.365 132.845 92.695 133.225 ;
        RECT 92.865 132.675 93.035 132.965 ;
        RECT 92.370 132.505 93.035 132.675 ;
        RECT 92.370 131.515 92.600 132.505 ;
        RECT 93.295 132.455 94.965 133.225 ;
        RECT 92.770 131.685 93.120 132.335 ;
        RECT 93.295 131.765 94.045 132.285 ;
        RECT 94.215 131.935 94.965 132.455 ;
        RECT 95.135 132.765 95.695 133.055 ;
        RECT 95.865 132.765 96.115 133.225 ;
        RECT 92.370 131.345 93.035 131.515 ;
        RECT 92.365 130.675 92.695 131.175 ;
        RECT 92.865 130.845 93.035 131.345 ;
        RECT 93.295 130.675 94.965 131.765 ;
        RECT 95.135 131.395 95.385 132.765 ;
        RECT 96.735 132.595 97.065 132.955 ;
        RECT 95.675 132.405 97.065 132.595 ;
        RECT 97.895 132.765 98.455 133.055 ;
        RECT 98.625 132.765 98.875 133.225 ;
        RECT 95.675 132.315 95.845 132.405 ;
        RECT 95.555 131.985 95.845 132.315 ;
        RECT 96.015 131.985 96.355 132.235 ;
        RECT 96.575 131.985 97.250 132.235 ;
        RECT 95.675 131.735 95.845 131.985 ;
        RECT 95.675 131.565 96.615 131.735 ;
        RECT 96.985 131.625 97.250 131.985 ;
        RECT 95.135 130.845 95.595 131.395 ;
        RECT 95.785 130.675 96.115 131.395 ;
        RECT 96.315 131.015 96.615 131.565 ;
        RECT 97.895 131.395 98.145 132.765 ;
        RECT 99.495 132.595 99.825 132.955 ;
        RECT 98.435 132.405 99.825 132.595 ;
        RECT 100.195 132.500 100.485 133.225 ;
        RECT 100.695 132.405 100.925 133.225 ;
        RECT 101.095 132.425 101.425 133.055 ;
        RECT 98.435 132.315 98.605 132.405 ;
        RECT 98.315 131.985 98.605 132.315 ;
        RECT 98.775 131.985 99.115 132.235 ;
        RECT 99.335 131.985 100.010 132.235 ;
        RECT 100.675 131.985 101.005 132.235 ;
        RECT 98.435 131.735 98.605 131.985 ;
        RECT 98.435 131.565 99.375 131.735 ;
        RECT 99.745 131.625 100.010 131.985 ;
        RECT 96.785 130.675 97.065 131.345 ;
        RECT 97.895 130.845 98.355 131.395 ;
        RECT 98.545 130.675 98.875 131.395 ;
        RECT 99.075 131.015 99.375 131.565 ;
        RECT 99.545 130.675 99.825 131.345 ;
        RECT 100.195 130.675 100.485 131.840 ;
        RECT 101.175 131.825 101.425 132.425 ;
        RECT 101.595 132.405 101.805 133.225 ;
        RECT 102.410 132.515 102.665 133.045 ;
        RECT 102.845 132.765 103.130 133.225 ;
        RECT 102.410 131.865 102.590 132.515 ;
        RECT 103.310 132.315 103.560 132.965 ;
        RECT 102.760 131.985 103.560 132.315 ;
        RECT 100.695 130.675 100.925 131.815 ;
        RECT 101.095 130.845 101.425 131.825 ;
        RECT 101.595 130.675 101.805 131.815 ;
        RECT 102.325 131.695 102.590 131.865 ;
        RECT 102.410 131.655 102.590 131.695 ;
        RECT 102.410 130.985 102.665 131.655 ;
        RECT 102.845 130.675 103.130 131.475 ;
        RECT 103.310 131.395 103.560 131.985 ;
        RECT 103.760 132.630 104.080 132.960 ;
        RECT 104.260 132.745 104.920 133.225 ;
        RECT 105.120 132.835 105.970 133.005 ;
        RECT 103.760 131.735 103.950 132.630 ;
        RECT 104.270 132.305 104.930 132.575 ;
        RECT 104.600 132.245 104.930 132.305 ;
        RECT 104.120 132.075 104.450 132.135 ;
        RECT 105.120 132.075 105.290 132.835 ;
        RECT 106.530 132.765 106.850 133.225 ;
        RECT 107.050 132.585 107.300 133.015 ;
        RECT 107.590 132.785 108.000 133.225 ;
        RECT 108.170 132.845 109.185 133.045 ;
        RECT 105.460 132.415 106.710 132.585 ;
        RECT 105.460 132.295 105.790 132.415 ;
        RECT 104.120 131.905 106.020 132.075 ;
        RECT 103.760 131.565 105.680 131.735 ;
        RECT 103.760 131.545 104.080 131.565 ;
        RECT 103.310 130.885 103.640 131.395 ;
        RECT 103.910 130.935 104.080 131.545 ;
        RECT 105.850 131.395 106.020 131.905 ;
        RECT 106.190 131.835 106.370 132.245 ;
        RECT 106.540 131.655 106.710 132.415 ;
        RECT 104.250 130.675 104.580 131.365 ;
        RECT 104.810 131.225 106.020 131.395 ;
        RECT 106.190 131.345 106.710 131.655 ;
        RECT 106.880 132.245 107.300 132.585 ;
        RECT 107.590 132.245 108.000 132.575 ;
        RECT 106.880 131.475 107.070 132.245 ;
        RECT 108.170 132.115 108.340 132.845 ;
        RECT 109.485 132.675 109.655 133.005 ;
        RECT 109.825 132.845 110.155 133.225 ;
        RECT 108.510 132.295 108.860 132.665 ;
        RECT 108.170 132.075 108.590 132.115 ;
        RECT 107.240 131.905 108.590 132.075 ;
        RECT 107.240 131.745 107.490 131.905 ;
        RECT 108.000 131.475 108.250 131.735 ;
        RECT 106.880 131.225 108.250 131.475 ;
        RECT 104.810 130.935 105.050 131.225 ;
        RECT 105.850 131.145 106.020 131.225 ;
        RECT 105.250 130.675 105.670 131.055 ;
        RECT 105.850 130.895 106.480 131.145 ;
        RECT 106.950 130.675 107.280 131.055 ;
        RECT 107.450 130.935 107.620 131.225 ;
        RECT 108.420 131.060 108.590 131.905 ;
        RECT 109.040 131.735 109.260 132.605 ;
        RECT 109.485 132.485 110.180 132.675 ;
        RECT 108.760 131.355 109.260 131.735 ;
        RECT 109.430 131.685 109.840 132.305 ;
        RECT 110.010 131.515 110.180 132.485 ;
        RECT 109.485 131.345 110.180 131.515 ;
        RECT 107.800 130.675 108.180 131.055 ;
        RECT 108.420 130.890 109.250 131.060 ;
        RECT 109.485 130.845 109.655 131.345 ;
        RECT 109.825 130.675 110.155 131.175 ;
        RECT 110.370 130.845 110.595 132.965 ;
        RECT 110.765 132.845 111.095 133.225 ;
        RECT 111.265 132.675 111.435 132.965 ;
        RECT 110.770 132.505 111.435 132.675 ;
        RECT 110.770 131.515 111.000 132.505 ;
        RECT 112.155 132.475 113.365 133.225 ;
        RECT 111.170 131.685 111.520 132.335 ;
        RECT 112.155 131.765 112.675 132.305 ;
        RECT 112.845 131.935 113.365 132.475 ;
        RECT 110.770 131.345 111.435 131.515 ;
        RECT 110.765 130.675 111.095 131.175 ;
        RECT 111.265 130.845 111.435 131.345 ;
        RECT 112.155 130.675 113.365 131.765 ;
        RECT 15.010 130.505 113.450 130.675 ;
        RECT 15.095 129.415 16.305 130.505 ;
        RECT 16.850 130.165 17.105 130.195 ;
        RECT 16.765 129.995 17.105 130.165 ;
        RECT 15.095 128.705 15.615 129.245 ;
        RECT 15.785 128.875 16.305 129.415 ;
        RECT 16.850 129.525 17.105 129.995 ;
        RECT 17.285 129.705 17.570 130.505 ;
        RECT 17.750 129.785 18.080 130.295 ;
        RECT 15.095 127.955 16.305 128.705 ;
        RECT 16.850 128.665 17.030 129.525 ;
        RECT 17.750 129.195 18.000 129.785 ;
        RECT 18.350 129.635 18.520 130.245 ;
        RECT 18.690 129.815 19.020 130.505 ;
        RECT 19.250 129.955 19.490 130.245 ;
        RECT 19.690 130.125 20.110 130.505 ;
        RECT 20.290 130.035 20.920 130.285 ;
        RECT 21.390 130.125 21.720 130.505 ;
        RECT 20.290 129.955 20.460 130.035 ;
        RECT 21.890 129.955 22.060 130.245 ;
        RECT 22.240 130.125 22.620 130.505 ;
        RECT 22.860 130.120 23.690 130.290 ;
        RECT 19.250 129.785 20.460 129.955 ;
        RECT 17.200 128.865 18.000 129.195 ;
        RECT 16.850 128.135 17.105 128.665 ;
        RECT 17.285 127.955 17.570 128.415 ;
        RECT 17.750 128.215 18.000 128.865 ;
        RECT 18.200 129.615 18.520 129.635 ;
        RECT 18.200 129.445 20.120 129.615 ;
        RECT 18.200 128.550 18.390 129.445 ;
        RECT 20.290 129.275 20.460 129.785 ;
        RECT 20.630 129.525 21.150 129.835 ;
        RECT 18.560 129.105 20.460 129.275 ;
        RECT 18.560 129.045 18.890 129.105 ;
        RECT 19.040 128.875 19.370 128.935 ;
        RECT 18.710 128.605 19.370 128.875 ;
        RECT 18.200 128.220 18.520 128.550 ;
        RECT 18.700 127.955 19.360 128.435 ;
        RECT 19.560 128.345 19.730 129.105 ;
        RECT 20.630 128.935 20.810 129.345 ;
        RECT 19.900 128.765 20.230 128.885 ;
        RECT 20.980 128.765 21.150 129.525 ;
        RECT 19.900 128.595 21.150 128.765 ;
        RECT 21.320 129.705 22.690 129.955 ;
        RECT 21.320 128.935 21.510 129.705 ;
        RECT 22.440 129.445 22.690 129.705 ;
        RECT 21.680 129.275 21.930 129.435 ;
        RECT 22.860 129.275 23.030 130.120 ;
        RECT 23.925 129.835 24.095 130.335 ;
        RECT 24.265 130.005 24.595 130.505 ;
        RECT 23.200 129.445 23.700 129.825 ;
        RECT 23.925 129.665 24.620 129.835 ;
        RECT 21.680 129.105 23.030 129.275 ;
        RECT 22.610 129.065 23.030 129.105 ;
        RECT 21.320 128.595 21.740 128.935 ;
        RECT 22.030 128.605 22.440 128.935 ;
        RECT 19.560 128.175 20.410 128.345 ;
        RECT 20.970 127.955 21.290 128.415 ;
        RECT 21.490 128.165 21.740 128.595 ;
        RECT 22.030 127.955 22.440 128.395 ;
        RECT 22.610 128.335 22.780 129.065 ;
        RECT 22.950 128.515 23.300 128.885 ;
        RECT 23.480 128.575 23.700 129.445 ;
        RECT 23.870 128.875 24.280 129.495 ;
        RECT 24.450 128.695 24.620 129.665 ;
        RECT 23.925 128.505 24.620 128.695 ;
        RECT 22.610 128.135 23.625 128.335 ;
        RECT 23.925 128.175 24.095 128.505 ;
        RECT 24.265 127.955 24.595 128.335 ;
        RECT 24.810 128.215 25.035 130.335 ;
        RECT 25.205 130.005 25.535 130.505 ;
        RECT 25.705 129.835 25.875 130.335 ;
        RECT 25.210 129.665 25.875 129.835 ;
        RECT 25.210 128.675 25.440 129.665 ;
        RECT 25.610 128.845 25.960 129.495 ;
        RECT 26.135 129.430 26.405 130.335 ;
        RECT 26.575 129.745 26.905 130.505 ;
        RECT 27.085 129.575 27.255 130.335 ;
        RECT 25.210 128.505 25.875 128.675 ;
        RECT 25.205 127.955 25.535 128.335 ;
        RECT 25.705 128.215 25.875 128.505 ;
        RECT 26.135 128.630 26.305 129.430 ;
        RECT 26.590 129.405 27.255 129.575 ;
        RECT 26.590 129.260 26.760 129.405 ;
        RECT 28.015 129.365 28.245 130.505 ;
        RECT 28.415 129.355 28.745 130.335 ;
        RECT 28.915 129.365 29.125 130.505 ;
        RECT 29.355 129.785 29.815 130.335 ;
        RECT 30.005 129.785 30.335 130.505 ;
        RECT 26.475 128.930 26.760 129.260 ;
        RECT 26.590 128.675 26.760 128.930 ;
        RECT 26.995 128.855 27.325 129.225 ;
        RECT 27.995 128.945 28.325 129.195 ;
        RECT 26.135 128.125 26.395 128.630 ;
        RECT 26.590 128.505 27.255 128.675 ;
        RECT 26.575 127.955 26.905 128.335 ;
        RECT 27.085 128.125 27.255 128.505 ;
        RECT 28.015 127.955 28.245 128.775 ;
        RECT 28.495 128.755 28.745 129.355 ;
        RECT 28.415 128.125 28.745 128.755 ;
        RECT 28.915 127.955 29.125 128.775 ;
        RECT 29.355 128.415 29.605 129.785 ;
        RECT 30.535 129.615 30.835 130.165 ;
        RECT 31.005 129.835 31.285 130.505 ;
        RECT 29.895 129.445 30.835 129.615 ;
        RECT 31.655 129.745 32.170 130.155 ;
        RECT 32.405 129.745 32.575 130.505 ;
        RECT 32.745 130.165 34.775 130.335 ;
        RECT 29.895 129.195 30.065 129.445 ;
        RECT 31.205 129.195 31.470 129.555 ;
        RECT 29.775 128.865 30.065 129.195 ;
        RECT 30.235 128.945 30.575 129.195 ;
        RECT 30.795 128.945 31.470 129.195 ;
        RECT 29.895 128.775 30.065 128.865 ;
        RECT 31.655 128.935 31.995 129.745 ;
        RECT 32.745 129.500 32.915 130.165 ;
        RECT 33.310 129.825 34.435 129.995 ;
        RECT 32.165 129.310 32.915 129.500 ;
        RECT 33.085 129.485 34.095 129.655 ;
        RECT 29.895 128.585 31.285 128.775 ;
        RECT 31.655 128.765 32.885 128.935 ;
        RECT 29.355 128.125 29.915 128.415 ;
        RECT 30.085 127.955 30.335 128.415 ;
        RECT 30.955 128.225 31.285 128.585 ;
        RECT 31.930 128.160 32.175 128.765 ;
        RECT 32.395 127.955 32.905 128.490 ;
        RECT 33.085 128.125 33.275 129.485 ;
        RECT 33.445 128.465 33.720 129.285 ;
        RECT 33.925 128.685 34.095 129.485 ;
        RECT 34.265 128.695 34.435 129.825 ;
        RECT 34.605 129.195 34.775 130.165 ;
        RECT 34.945 129.365 35.115 130.505 ;
        RECT 35.285 129.365 35.620 130.335 ;
        RECT 34.605 128.865 34.800 129.195 ;
        RECT 35.025 128.865 35.280 129.195 ;
        RECT 35.025 128.695 35.195 128.865 ;
        RECT 35.450 128.695 35.620 129.365 ;
        RECT 35.795 129.340 36.085 130.505 ;
        RECT 36.255 129.430 36.525 130.335 ;
        RECT 36.695 129.745 37.025 130.505 ;
        RECT 37.205 129.575 37.375 130.335 ;
        RECT 34.265 128.525 35.195 128.695 ;
        RECT 34.265 128.490 34.440 128.525 ;
        RECT 33.445 128.295 33.725 128.465 ;
        RECT 33.445 128.125 33.720 128.295 ;
        RECT 33.910 128.125 34.440 128.490 ;
        RECT 34.865 127.955 35.195 128.355 ;
        RECT 35.365 128.125 35.620 128.695 ;
        RECT 35.795 127.955 36.085 128.680 ;
        RECT 36.255 128.630 36.425 129.430 ;
        RECT 36.710 129.405 37.375 129.575 ;
        RECT 36.710 129.260 36.880 129.405 ;
        RECT 36.595 128.930 36.880 129.260 ;
        RECT 37.640 129.365 37.975 130.335 ;
        RECT 38.145 129.365 38.315 130.505 ;
        RECT 38.485 130.165 40.515 130.335 ;
        RECT 36.710 128.675 36.880 128.930 ;
        RECT 37.115 128.855 37.445 129.225 ;
        RECT 37.640 128.695 37.810 129.365 ;
        RECT 38.485 129.195 38.655 130.165 ;
        RECT 37.980 128.865 38.235 129.195 ;
        RECT 38.460 128.865 38.655 129.195 ;
        RECT 38.825 129.825 39.950 129.995 ;
        RECT 38.065 128.695 38.235 128.865 ;
        RECT 38.825 128.695 38.995 129.825 ;
        RECT 36.255 128.125 36.515 128.630 ;
        RECT 36.710 128.505 37.375 128.675 ;
        RECT 36.695 127.955 37.025 128.335 ;
        RECT 37.205 128.125 37.375 128.505 ;
        RECT 37.640 128.125 37.895 128.695 ;
        RECT 38.065 128.525 38.995 128.695 ;
        RECT 39.165 129.485 40.175 129.655 ;
        RECT 39.165 128.685 39.335 129.485 ;
        RECT 38.820 128.490 38.995 128.525 ;
        RECT 38.065 127.955 38.395 128.355 ;
        RECT 38.820 128.125 39.350 128.490 ;
        RECT 39.540 128.465 39.815 129.285 ;
        RECT 39.535 128.295 39.815 128.465 ;
        RECT 39.540 128.125 39.815 128.295 ;
        RECT 39.985 128.125 40.175 129.485 ;
        RECT 40.345 129.500 40.515 130.165 ;
        RECT 40.685 129.745 40.855 130.505 ;
        RECT 41.090 129.745 41.605 130.155 ;
        RECT 40.345 129.310 41.095 129.500 ;
        RECT 41.265 128.935 41.605 129.745 ;
        RECT 40.375 128.765 41.605 128.935 ;
        RECT 41.775 129.415 43.445 130.505 ;
        RECT 43.625 129.695 43.920 130.505 ;
        RECT 41.775 128.895 42.525 129.415 ;
        RECT 40.355 127.955 40.865 128.490 ;
        RECT 41.085 128.160 41.330 128.765 ;
        RECT 42.695 128.725 43.445 129.245 ;
        RECT 44.100 129.195 44.345 130.335 ;
        RECT 44.520 129.695 44.780 130.505 ;
        RECT 45.380 130.500 51.655 130.505 ;
        RECT 44.960 129.195 45.210 130.330 ;
        RECT 45.380 129.705 45.640 130.500 ;
        RECT 45.810 129.605 46.070 130.330 ;
        RECT 46.240 129.775 46.500 130.500 ;
        RECT 46.670 129.605 46.930 130.330 ;
        RECT 47.100 129.775 47.360 130.500 ;
        RECT 47.530 129.605 47.790 130.330 ;
        RECT 47.960 129.775 48.220 130.500 ;
        RECT 48.390 129.605 48.650 130.330 ;
        RECT 48.820 129.775 49.065 130.500 ;
        RECT 49.235 129.605 49.495 130.330 ;
        RECT 49.680 129.775 49.925 130.500 ;
        RECT 50.095 129.605 50.355 130.330 ;
        RECT 50.540 129.775 50.785 130.500 ;
        RECT 50.955 129.605 51.215 130.330 ;
        RECT 51.400 129.775 51.655 130.500 ;
        RECT 45.810 129.590 51.215 129.605 ;
        RECT 51.825 129.590 52.115 130.330 ;
        RECT 52.285 129.760 52.555 130.505 ;
        RECT 53.275 129.745 53.790 130.155 ;
        RECT 54.025 129.745 54.195 130.505 ;
        RECT 54.365 130.165 56.395 130.335 ;
        RECT 45.810 129.365 52.555 129.590 ;
        RECT 41.775 127.955 43.445 128.725 ;
        RECT 43.615 128.635 43.930 129.195 ;
        RECT 44.100 128.945 51.220 129.195 ;
        RECT 43.615 127.955 43.920 128.465 ;
        RECT 44.100 128.135 44.350 128.945 ;
        RECT 44.520 127.955 44.780 128.480 ;
        RECT 44.960 128.135 45.210 128.945 ;
        RECT 51.390 128.775 52.555 129.365 ;
        RECT 45.810 128.605 52.555 128.775 ;
        RECT 53.275 128.935 53.615 129.745 ;
        RECT 54.365 129.500 54.535 130.165 ;
        RECT 54.930 129.825 56.055 129.995 ;
        RECT 53.785 129.310 54.535 129.500 ;
        RECT 54.705 129.485 55.715 129.655 ;
        RECT 53.275 128.765 54.505 128.935 ;
        RECT 45.380 127.955 45.640 128.515 ;
        RECT 45.810 128.150 46.070 128.605 ;
        RECT 46.240 127.955 46.500 128.435 ;
        RECT 46.670 128.150 46.930 128.605 ;
        RECT 47.100 127.955 47.360 128.435 ;
        RECT 47.530 128.150 47.790 128.605 ;
        RECT 47.960 127.955 48.205 128.435 ;
        RECT 48.375 128.150 48.650 128.605 ;
        RECT 48.820 127.955 49.065 128.435 ;
        RECT 49.235 128.150 49.495 128.605 ;
        RECT 49.675 127.955 49.925 128.435 ;
        RECT 50.095 128.150 50.355 128.605 ;
        RECT 50.535 127.955 50.785 128.435 ;
        RECT 50.955 128.150 51.215 128.605 ;
        RECT 51.395 127.955 51.655 128.435 ;
        RECT 51.825 128.150 52.085 128.605 ;
        RECT 52.255 127.955 52.555 128.435 ;
        RECT 53.550 128.160 53.795 128.765 ;
        RECT 54.015 127.955 54.525 128.490 ;
        RECT 54.705 128.125 54.895 129.485 ;
        RECT 55.065 129.145 55.340 129.285 ;
        RECT 55.065 128.975 55.345 129.145 ;
        RECT 55.065 128.125 55.340 128.975 ;
        RECT 55.545 128.685 55.715 129.485 ;
        RECT 55.885 128.695 56.055 129.825 ;
        RECT 56.225 129.195 56.395 130.165 ;
        RECT 56.565 129.365 56.735 130.505 ;
        RECT 56.905 129.365 57.240 130.335 ;
        RECT 56.225 128.865 56.420 129.195 ;
        RECT 56.645 128.865 56.900 129.195 ;
        RECT 56.645 128.695 56.815 128.865 ;
        RECT 57.070 128.695 57.240 129.365 ;
        RECT 57.415 129.745 57.930 130.155 ;
        RECT 58.165 129.745 58.335 130.505 ;
        RECT 58.505 130.165 60.535 130.335 ;
        RECT 57.415 128.935 57.755 129.745 ;
        RECT 58.505 129.500 58.675 130.165 ;
        RECT 59.070 129.825 60.195 129.995 ;
        RECT 57.925 129.310 58.675 129.500 ;
        RECT 58.845 129.485 59.855 129.655 ;
        RECT 57.415 128.765 58.645 128.935 ;
        RECT 55.885 128.525 56.815 128.695 ;
        RECT 55.885 128.490 56.060 128.525 ;
        RECT 55.530 128.125 56.060 128.490 ;
        RECT 56.485 127.955 56.815 128.355 ;
        RECT 56.985 128.125 57.240 128.695 ;
        RECT 57.690 128.160 57.935 128.765 ;
        RECT 58.155 127.955 58.665 128.490 ;
        RECT 58.845 128.125 59.035 129.485 ;
        RECT 59.205 128.805 59.480 129.285 ;
        RECT 59.205 128.635 59.485 128.805 ;
        RECT 59.685 128.685 59.855 129.485 ;
        RECT 60.025 128.695 60.195 129.825 ;
        RECT 60.365 129.195 60.535 130.165 ;
        RECT 60.705 129.365 60.875 130.505 ;
        RECT 61.045 129.365 61.380 130.335 ;
        RECT 60.365 128.865 60.560 129.195 ;
        RECT 60.785 128.865 61.040 129.195 ;
        RECT 60.785 128.695 60.955 128.865 ;
        RECT 61.210 128.695 61.380 129.365 ;
        RECT 61.555 129.340 61.845 130.505 ;
        RECT 62.940 130.080 63.275 130.505 ;
        RECT 63.445 129.900 63.630 130.305 ;
        RECT 62.965 129.725 63.630 129.900 ;
        RECT 63.835 129.725 64.165 130.505 ;
        RECT 59.205 128.125 59.480 128.635 ;
        RECT 60.025 128.525 60.955 128.695 ;
        RECT 60.025 128.490 60.200 128.525 ;
        RECT 59.670 128.125 60.200 128.490 ;
        RECT 60.625 127.955 60.955 128.355 ;
        RECT 61.125 128.125 61.380 128.695 ;
        RECT 62.965 128.695 63.305 129.725 ;
        RECT 64.335 129.535 64.605 130.305 ;
        RECT 63.475 129.365 64.605 129.535 ;
        RECT 63.475 128.865 63.725 129.365 ;
        RECT 61.555 127.955 61.845 128.680 ;
        RECT 62.965 128.525 63.650 128.695 ;
        RECT 63.905 128.615 64.265 129.195 ;
        RECT 62.940 127.955 63.275 128.355 ;
        RECT 63.445 128.125 63.650 128.525 ;
        RECT 64.435 128.455 64.605 129.365 ;
        RECT 63.860 127.955 64.135 128.435 ;
        RECT 64.345 128.125 64.605 128.455 ;
        RECT 64.775 129.535 65.085 130.335 ;
        RECT 65.255 129.705 65.565 130.505 ;
        RECT 65.735 129.875 65.995 130.335 ;
        RECT 66.165 130.045 66.420 130.505 ;
        RECT 66.595 129.875 66.855 130.335 ;
        RECT 65.735 129.705 66.855 129.875 ;
        RECT 64.775 129.365 65.805 129.535 ;
        RECT 64.775 128.455 64.945 129.365 ;
        RECT 65.115 128.625 65.465 129.195 ;
        RECT 65.635 129.115 65.805 129.365 ;
        RECT 66.595 129.455 66.855 129.705 ;
        RECT 67.025 129.635 67.310 130.505 ;
        RECT 66.595 129.285 67.350 129.455 ;
        RECT 65.635 128.945 66.775 129.115 ;
        RECT 66.945 128.775 67.350 129.285 ;
        RECT 67.535 129.415 68.745 130.505 ;
        RECT 68.915 129.745 69.430 130.155 ;
        RECT 69.665 129.745 69.835 130.505 ;
        RECT 70.005 130.165 72.035 130.335 ;
        RECT 67.535 128.875 68.055 129.415 ;
        RECT 65.700 128.605 67.350 128.775 ;
        RECT 68.225 128.705 68.745 129.245 ;
        RECT 68.915 128.935 69.255 129.745 ;
        RECT 70.005 129.500 70.175 130.165 ;
        RECT 70.570 129.825 71.695 129.995 ;
        RECT 69.425 129.310 70.175 129.500 ;
        RECT 70.345 129.485 71.355 129.655 ;
        RECT 68.915 128.765 70.145 128.935 ;
        RECT 64.775 128.125 65.075 128.455 ;
        RECT 65.245 127.955 65.520 128.435 ;
        RECT 65.700 128.215 65.995 128.605 ;
        RECT 66.165 127.955 66.420 128.435 ;
        RECT 66.595 128.215 66.855 128.605 ;
        RECT 67.025 127.955 67.305 128.435 ;
        RECT 67.535 127.955 68.745 128.705 ;
        RECT 69.190 128.160 69.435 128.765 ;
        RECT 69.655 127.955 70.165 128.490 ;
        RECT 70.345 128.125 70.535 129.485 ;
        RECT 70.705 128.465 70.980 129.285 ;
        RECT 71.185 128.685 71.355 129.485 ;
        RECT 71.525 128.695 71.695 129.825 ;
        RECT 71.865 129.195 72.035 130.165 ;
        RECT 72.205 129.365 72.375 130.505 ;
        RECT 72.545 129.365 72.880 130.335 ;
        RECT 73.145 129.835 73.315 130.335 ;
        RECT 73.485 130.005 73.815 130.505 ;
        RECT 73.145 129.665 73.810 129.835 ;
        RECT 71.865 128.865 72.060 129.195 ;
        RECT 72.285 128.865 72.540 129.195 ;
        RECT 72.285 128.695 72.455 128.865 ;
        RECT 72.710 128.695 72.880 129.365 ;
        RECT 73.060 128.845 73.410 129.495 ;
        RECT 71.525 128.525 72.455 128.695 ;
        RECT 71.525 128.490 71.700 128.525 ;
        RECT 70.705 128.295 70.985 128.465 ;
        RECT 70.705 128.125 70.980 128.295 ;
        RECT 71.170 128.125 71.700 128.490 ;
        RECT 72.125 127.955 72.455 128.355 ;
        RECT 72.625 128.125 72.880 128.695 ;
        RECT 73.580 128.675 73.810 129.665 ;
        RECT 73.145 128.505 73.810 128.675 ;
        RECT 73.145 128.215 73.315 128.505 ;
        RECT 73.485 127.955 73.815 128.335 ;
        RECT 73.985 128.215 74.210 130.335 ;
        RECT 74.425 130.005 74.755 130.505 ;
        RECT 74.925 129.835 75.095 130.335 ;
        RECT 75.330 130.120 76.160 130.290 ;
        RECT 76.400 130.125 76.780 130.505 ;
        RECT 74.400 129.665 75.095 129.835 ;
        RECT 74.400 128.695 74.570 129.665 ;
        RECT 74.740 128.875 75.150 129.495 ;
        RECT 75.320 129.445 75.820 129.825 ;
        RECT 74.400 128.505 75.095 128.695 ;
        RECT 75.320 128.575 75.540 129.445 ;
        RECT 75.990 129.275 76.160 130.120 ;
        RECT 76.960 129.955 77.130 130.245 ;
        RECT 77.300 130.125 77.630 130.505 ;
        RECT 78.100 130.035 78.730 130.285 ;
        RECT 78.910 130.125 79.330 130.505 ;
        RECT 78.560 129.955 78.730 130.035 ;
        RECT 79.530 129.955 79.770 130.245 ;
        RECT 76.330 129.705 77.700 129.955 ;
        RECT 76.330 129.445 76.580 129.705 ;
        RECT 77.090 129.275 77.340 129.435 ;
        RECT 75.990 129.105 77.340 129.275 ;
        RECT 75.990 129.065 76.410 129.105 ;
        RECT 75.720 128.515 76.070 128.885 ;
        RECT 74.425 127.955 74.755 128.335 ;
        RECT 74.925 128.175 75.095 128.505 ;
        RECT 76.240 128.335 76.410 129.065 ;
        RECT 77.510 128.935 77.700 129.705 ;
        RECT 76.580 128.605 76.990 128.935 ;
        RECT 77.280 128.595 77.700 128.935 ;
        RECT 77.870 129.525 78.390 129.835 ;
        RECT 78.560 129.785 79.770 129.955 ;
        RECT 80.000 129.815 80.330 130.505 ;
        RECT 77.870 128.765 78.040 129.525 ;
        RECT 78.210 128.935 78.390 129.345 ;
        RECT 78.560 129.275 78.730 129.785 ;
        RECT 80.500 129.635 80.670 130.245 ;
        RECT 80.940 129.785 81.270 130.295 ;
        RECT 80.500 129.615 80.820 129.635 ;
        RECT 78.900 129.445 80.820 129.615 ;
        RECT 78.560 129.105 80.460 129.275 ;
        RECT 78.790 128.765 79.120 128.885 ;
        RECT 77.870 128.595 79.120 128.765 ;
        RECT 75.395 128.135 76.410 128.335 ;
        RECT 76.580 127.955 76.990 128.395 ;
        RECT 77.280 128.165 77.530 128.595 ;
        RECT 77.730 127.955 78.050 128.415 ;
        RECT 79.290 128.345 79.460 129.105 ;
        RECT 80.130 129.045 80.460 129.105 ;
        RECT 79.650 128.875 79.980 128.935 ;
        RECT 79.650 128.605 80.310 128.875 ;
        RECT 80.630 128.550 80.820 129.445 ;
        RECT 78.610 128.175 79.460 128.345 ;
        RECT 79.660 127.955 80.320 128.435 ;
        RECT 80.500 128.220 80.820 128.550 ;
        RECT 81.020 129.195 81.270 129.785 ;
        RECT 81.450 129.705 81.735 130.505 ;
        RECT 81.915 129.525 82.170 130.195 ;
        RECT 81.020 128.865 81.820 129.195 ;
        RECT 81.020 128.215 81.270 128.865 ;
        RECT 81.990 128.665 82.170 129.525 ;
        RECT 83.175 129.745 83.690 130.155 ;
        RECT 83.925 129.745 84.095 130.505 ;
        RECT 84.265 130.165 86.295 130.335 ;
        RECT 83.175 128.935 83.515 129.745 ;
        RECT 84.265 129.500 84.435 130.165 ;
        RECT 84.830 129.825 85.955 129.995 ;
        RECT 83.685 129.310 84.435 129.500 ;
        RECT 84.605 129.485 85.615 129.655 ;
        RECT 83.175 128.765 84.405 128.935 ;
        RECT 81.915 128.465 82.170 128.665 ;
        RECT 81.450 127.955 81.735 128.415 ;
        RECT 81.915 128.295 82.255 128.465 ;
        RECT 81.915 128.135 82.170 128.295 ;
        RECT 83.450 128.160 83.695 128.765 ;
        RECT 83.915 127.955 84.425 128.490 ;
        RECT 84.605 128.125 84.795 129.485 ;
        RECT 84.965 128.805 85.240 129.285 ;
        RECT 84.965 128.635 85.245 128.805 ;
        RECT 85.445 128.685 85.615 129.485 ;
        RECT 85.785 128.695 85.955 129.825 ;
        RECT 86.125 129.195 86.295 130.165 ;
        RECT 86.465 129.365 86.635 130.505 ;
        RECT 86.805 129.365 87.140 130.335 ;
        RECT 86.125 128.865 86.320 129.195 ;
        RECT 86.545 128.865 86.800 129.195 ;
        RECT 86.545 128.695 86.715 128.865 ;
        RECT 86.970 128.695 87.140 129.365 ;
        RECT 87.315 129.340 87.605 130.505 ;
        RECT 88.435 129.835 88.715 130.505 ;
        RECT 88.885 129.615 89.185 130.165 ;
        RECT 89.385 129.785 89.715 130.505 ;
        RECT 89.905 129.785 90.365 130.335 ;
        RECT 88.250 129.195 88.515 129.555 ;
        RECT 88.885 129.445 89.825 129.615 ;
        RECT 89.655 129.195 89.825 129.445 ;
        RECT 88.250 128.945 88.925 129.195 ;
        RECT 89.145 128.945 89.485 129.195 ;
        RECT 89.655 128.865 89.945 129.195 ;
        RECT 89.655 128.775 89.825 128.865 ;
        RECT 84.965 128.125 85.240 128.635 ;
        RECT 85.785 128.525 86.715 128.695 ;
        RECT 85.785 128.490 85.960 128.525 ;
        RECT 85.430 128.125 85.960 128.490 ;
        RECT 86.385 127.955 86.715 128.355 ;
        RECT 86.885 128.125 87.140 128.695 ;
        RECT 87.315 127.955 87.605 128.680 ;
        RECT 88.435 128.585 89.825 128.775 ;
        RECT 88.435 128.225 88.765 128.585 ;
        RECT 90.115 128.415 90.365 129.785 ;
        RECT 90.625 129.575 90.795 130.335 ;
        RECT 90.975 129.745 91.305 130.505 ;
        RECT 90.625 129.405 91.290 129.575 ;
        RECT 91.475 129.430 91.745 130.335 ;
        RECT 91.120 129.260 91.290 129.405 ;
        RECT 90.555 128.855 90.885 129.225 ;
        RECT 91.120 128.930 91.405 129.260 ;
        RECT 91.120 128.675 91.290 128.930 ;
        RECT 89.385 127.955 89.635 128.415 ;
        RECT 89.805 128.125 90.365 128.415 ;
        RECT 90.625 128.505 91.290 128.675 ;
        RECT 91.575 128.630 91.745 129.430 ;
        RECT 91.915 129.415 93.125 130.505 ;
        RECT 93.495 129.835 93.775 130.505 ;
        RECT 93.945 129.615 94.245 130.165 ;
        RECT 94.445 129.785 94.775 130.505 ;
        RECT 94.965 129.785 95.425 130.335 ;
        RECT 91.915 128.875 92.435 129.415 ;
        RECT 92.605 128.705 93.125 129.245 ;
        RECT 93.310 129.195 93.575 129.555 ;
        RECT 93.945 129.445 94.885 129.615 ;
        RECT 94.715 129.195 94.885 129.445 ;
        RECT 93.310 128.945 93.985 129.195 ;
        RECT 94.205 128.945 94.545 129.195 ;
        RECT 94.715 128.865 95.005 129.195 ;
        RECT 94.715 128.775 94.885 128.865 ;
        RECT 90.625 128.125 90.795 128.505 ;
        RECT 90.975 127.955 91.305 128.335 ;
        RECT 91.485 128.125 91.745 128.630 ;
        RECT 91.915 127.955 93.125 128.705 ;
        RECT 93.495 128.585 94.885 128.775 ;
        RECT 93.495 128.225 93.825 128.585 ;
        RECT 95.175 128.415 95.425 129.785 ;
        RECT 94.445 127.955 94.695 128.415 ;
        RECT 94.865 128.125 95.425 128.415 ;
        RECT 96.515 129.785 96.975 130.335 ;
        RECT 97.165 129.785 97.495 130.505 ;
        RECT 96.515 128.415 96.765 129.785 ;
        RECT 97.695 129.615 97.995 130.165 ;
        RECT 98.165 129.835 98.445 130.505 ;
        RECT 97.055 129.445 97.995 129.615 ;
        RECT 99.735 129.745 100.250 130.155 ;
        RECT 100.485 129.745 100.655 130.505 ;
        RECT 100.825 130.165 102.855 130.335 ;
        RECT 97.055 129.195 97.225 129.445 ;
        RECT 98.365 129.195 98.630 129.555 ;
        RECT 96.935 128.865 97.225 129.195 ;
        RECT 97.395 128.945 97.735 129.195 ;
        RECT 97.955 128.945 98.630 129.195 ;
        RECT 97.055 128.775 97.225 128.865 ;
        RECT 99.735 128.935 100.075 129.745 ;
        RECT 100.825 129.500 100.995 130.165 ;
        RECT 101.390 129.825 102.515 129.995 ;
        RECT 100.245 129.310 100.995 129.500 ;
        RECT 101.165 129.485 102.175 129.655 ;
        RECT 97.055 128.585 98.445 128.775 ;
        RECT 99.735 128.765 100.965 128.935 ;
        RECT 96.515 128.125 97.075 128.415 ;
        RECT 97.245 127.955 97.495 128.415 ;
        RECT 98.115 128.225 98.445 128.585 ;
        RECT 100.010 128.160 100.255 128.765 ;
        RECT 100.475 127.955 100.985 128.490 ;
        RECT 101.165 128.125 101.355 129.485 ;
        RECT 101.525 129.145 101.800 129.285 ;
        RECT 101.525 128.975 101.805 129.145 ;
        RECT 101.525 128.125 101.800 128.975 ;
        RECT 102.005 128.685 102.175 129.485 ;
        RECT 102.345 128.695 102.515 129.825 ;
        RECT 102.685 129.195 102.855 130.165 ;
        RECT 103.025 129.365 103.195 130.505 ;
        RECT 103.365 129.365 103.700 130.335 ;
        RECT 102.685 128.865 102.880 129.195 ;
        RECT 103.105 128.865 103.360 129.195 ;
        RECT 103.105 128.695 103.275 128.865 ;
        RECT 103.530 128.695 103.700 129.365 ;
        RECT 103.875 129.745 104.390 130.155 ;
        RECT 104.625 129.745 104.795 130.505 ;
        RECT 104.965 130.165 106.995 130.335 ;
        RECT 103.875 128.935 104.215 129.745 ;
        RECT 104.965 129.500 105.135 130.165 ;
        RECT 105.530 129.825 106.655 129.995 ;
        RECT 104.385 129.310 105.135 129.500 ;
        RECT 105.305 129.485 106.315 129.655 ;
        RECT 103.875 128.765 105.105 128.935 ;
        RECT 102.345 128.525 103.275 128.695 ;
        RECT 102.345 128.490 102.520 128.525 ;
        RECT 101.990 128.125 102.520 128.490 ;
        RECT 102.945 127.955 103.275 128.355 ;
        RECT 103.445 128.125 103.700 128.695 ;
        RECT 104.150 128.160 104.395 128.765 ;
        RECT 104.615 127.955 105.125 128.490 ;
        RECT 105.305 128.125 105.495 129.485 ;
        RECT 105.665 128.465 105.940 129.285 ;
        RECT 106.145 128.685 106.315 129.485 ;
        RECT 106.485 128.695 106.655 129.825 ;
        RECT 106.825 129.195 106.995 130.165 ;
        RECT 107.165 129.365 107.335 130.505 ;
        RECT 107.505 129.365 107.840 130.335 ;
        RECT 108.105 129.575 108.275 130.335 ;
        RECT 108.455 129.745 108.785 130.505 ;
        RECT 108.105 129.405 108.770 129.575 ;
        RECT 108.955 129.430 109.225 130.335 ;
        RECT 106.825 128.865 107.020 129.195 ;
        RECT 107.245 128.865 107.500 129.195 ;
        RECT 107.245 128.695 107.415 128.865 ;
        RECT 107.670 128.695 107.840 129.365 ;
        RECT 108.600 129.260 108.770 129.405 ;
        RECT 108.035 128.855 108.365 129.225 ;
        RECT 108.600 128.930 108.885 129.260 ;
        RECT 106.485 128.525 107.415 128.695 ;
        RECT 106.485 128.490 106.660 128.525 ;
        RECT 105.665 128.295 105.945 128.465 ;
        RECT 105.665 128.125 105.940 128.295 ;
        RECT 106.130 128.125 106.660 128.490 ;
        RECT 107.085 127.955 107.415 128.355 ;
        RECT 107.585 128.125 107.840 128.695 ;
        RECT 108.600 128.675 108.770 128.930 ;
        RECT 108.105 128.505 108.770 128.675 ;
        RECT 109.055 128.630 109.225 129.430 ;
        RECT 109.395 129.415 111.985 130.505 ;
        RECT 112.155 129.415 113.365 130.505 ;
        RECT 109.395 128.895 110.605 129.415 ;
        RECT 110.775 128.725 111.985 129.245 ;
        RECT 112.155 128.875 112.675 129.415 ;
        RECT 108.105 128.125 108.275 128.505 ;
        RECT 108.455 127.955 108.785 128.335 ;
        RECT 108.965 128.125 109.225 128.630 ;
        RECT 109.395 127.955 111.985 128.725 ;
        RECT 112.845 128.705 113.365 129.245 ;
        RECT 112.155 127.955 113.365 128.705 ;
        RECT 15.010 127.785 113.450 127.955 ;
        RECT 15.095 127.035 16.305 127.785 ;
        RECT 15.095 126.495 15.615 127.035 ;
        RECT 16.475 127.015 19.985 127.785 ;
        RECT 15.785 126.325 16.305 126.865 ;
        RECT 15.095 125.235 16.305 126.325 ;
        RECT 16.475 126.325 18.165 126.845 ;
        RECT 18.335 126.495 19.985 127.015 ;
        RECT 20.215 126.965 20.425 127.785 ;
        RECT 20.595 126.985 20.925 127.615 ;
        RECT 20.595 126.385 20.845 126.985 ;
        RECT 21.095 126.965 21.325 127.785 ;
        RECT 21.535 127.035 22.745 127.785 ;
        RECT 22.915 127.060 23.205 127.785 ;
        RECT 21.015 126.545 21.345 126.795 ;
        RECT 16.475 125.235 19.985 126.325 ;
        RECT 20.215 125.235 20.425 126.375 ;
        RECT 20.595 125.405 20.925 126.385 ;
        RECT 21.095 125.235 21.325 126.375 ;
        RECT 21.535 126.325 22.055 126.865 ;
        RECT 22.225 126.495 22.745 127.035 ;
        RECT 24.300 127.045 24.555 127.615 ;
        RECT 24.725 127.385 25.055 127.785 ;
        RECT 25.480 127.250 26.010 127.615 ;
        RECT 26.200 127.445 26.475 127.615 ;
        RECT 26.195 127.275 26.475 127.445 ;
        RECT 25.480 127.215 25.655 127.250 ;
        RECT 24.725 127.045 25.655 127.215 ;
        RECT 21.535 125.235 22.745 126.325 ;
        RECT 22.915 125.235 23.205 126.400 ;
        RECT 24.300 126.375 24.470 127.045 ;
        RECT 24.725 126.875 24.895 127.045 ;
        RECT 24.640 126.545 24.895 126.875 ;
        RECT 25.120 126.545 25.315 126.875 ;
        RECT 24.300 125.405 24.635 126.375 ;
        RECT 24.805 125.235 24.975 126.375 ;
        RECT 25.145 125.575 25.315 126.545 ;
        RECT 25.485 125.915 25.655 127.045 ;
        RECT 25.825 126.255 25.995 127.055 ;
        RECT 26.200 126.455 26.475 127.275 ;
        RECT 26.645 126.255 26.835 127.615 ;
        RECT 27.015 127.250 27.525 127.785 ;
        RECT 27.745 126.975 27.990 127.580 ;
        RECT 28.895 127.015 31.485 127.785 ;
        RECT 32.030 127.445 32.285 127.605 ;
        RECT 31.945 127.275 32.285 127.445 ;
        RECT 32.465 127.325 32.750 127.785 ;
        RECT 27.035 126.805 28.265 126.975 ;
        RECT 25.825 126.085 26.835 126.255 ;
        RECT 27.005 126.240 27.755 126.430 ;
        RECT 25.485 125.745 26.610 125.915 ;
        RECT 27.005 125.575 27.175 126.240 ;
        RECT 27.925 125.995 28.265 126.805 ;
        RECT 25.145 125.405 27.175 125.575 ;
        RECT 27.345 125.235 27.515 125.995 ;
        RECT 27.750 125.585 28.265 125.995 ;
        RECT 28.895 126.325 30.105 126.845 ;
        RECT 30.275 126.495 31.485 127.015 ;
        RECT 32.030 127.075 32.285 127.275 ;
        RECT 28.895 125.235 31.485 126.325 ;
        RECT 32.030 126.215 32.210 127.075 ;
        RECT 32.930 126.875 33.180 127.525 ;
        RECT 32.380 126.545 33.180 126.875 ;
        RECT 32.030 125.545 32.285 126.215 ;
        RECT 32.465 125.235 32.750 126.035 ;
        RECT 32.930 125.955 33.180 126.545 ;
        RECT 33.380 127.190 33.700 127.520 ;
        RECT 33.880 127.305 34.540 127.785 ;
        RECT 34.740 127.395 35.590 127.565 ;
        RECT 33.380 126.295 33.570 127.190 ;
        RECT 33.890 126.865 34.550 127.135 ;
        RECT 34.220 126.805 34.550 126.865 ;
        RECT 33.740 126.635 34.070 126.695 ;
        RECT 34.740 126.635 34.910 127.395 ;
        RECT 36.150 127.325 36.470 127.785 ;
        RECT 36.670 127.145 36.920 127.575 ;
        RECT 37.210 127.345 37.620 127.785 ;
        RECT 37.790 127.405 38.805 127.605 ;
        RECT 35.080 126.975 36.330 127.145 ;
        RECT 35.080 126.855 35.410 126.975 ;
        RECT 33.740 126.465 35.640 126.635 ;
        RECT 33.380 126.125 35.300 126.295 ;
        RECT 33.380 126.105 33.700 126.125 ;
        RECT 32.930 125.445 33.260 125.955 ;
        RECT 33.530 125.495 33.700 126.105 ;
        RECT 35.470 125.955 35.640 126.465 ;
        RECT 35.810 126.395 35.990 126.805 ;
        RECT 36.160 126.215 36.330 126.975 ;
        RECT 33.870 125.235 34.200 125.925 ;
        RECT 34.430 125.785 35.640 125.955 ;
        RECT 35.810 125.905 36.330 126.215 ;
        RECT 36.500 126.805 36.920 127.145 ;
        RECT 37.210 126.805 37.620 127.135 ;
        RECT 36.500 126.035 36.690 126.805 ;
        RECT 37.790 126.675 37.960 127.405 ;
        RECT 39.105 127.235 39.275 127.565 ;
        RECT 39.445 127.405 39.775 127.785 ;
        RECT 38.130 126.855 38.480 127.225 ;
        RECT 37.790 126.635 38.210 126.675 ;
        RECT 36.860 126.465 38.210 126.635 ;
        RECT 36.860 126.305 37.110 126.465 ;
        RECT 37.620 126.035 37.870 126.295 ;
        RECT 36.500 125.785 37.870 126.035 ;
        RECT 34.430 125.495 34.670 125.785 ;
        RECT 35.470 125.705 35.640 125.785 ;
        RECT 34.870 125.235 35.290 125.615 ;
        RECT 35.470 125.455 36.100 125.705 ;
        RECT 36.570 125.235 36.900 125.615 ;
        RECT 37.070 125.495 37.240 125.785 ;
        RECT 38.040 125.620 38.210 126.465 ;
        RECT 38.660 126.295 38.880 127.165 ;
        RECT 39.105 127.045 39.800 127.235 ;
        RECT 38.380 125.915 38.880 126.295 ;
        RECT 39.050 126.245 39.460 126.865 ;
        RECT 39.630 126.075 39.800 127.045 ;
        RECT 39.105 125.905 39.800 126.075 ;
        RECT 37.420 125.235 37.800 125.615 ;
        RECT 38.040 125.450 38.870 125.620 ;
        RECT 39.105 125.405 39.275 125.905 ;
        RECT 39.445 125.235 39.775 125.735 ;
        RECT 39.990 125.405 40.215 127.525 ;
        RECT 40.385 127.405 40.715 127.785 ;
        RECT 40.885 127.235 41.055 127.525 ;
        RECT 40.390 127.065 41.055 127.235 ;
        RECT 41.315 127.325 41.875 127.615 ;
        RECT 42.045 127.325 42.295 127.785 ;
        RECT 40.390 126.075 40.620 127.065 ;
        RECT 40.790 126.245 41.140 126.895 ;
        RECT 40.390 125.905 41.055 126.075 ;
        RECT 40.385 125.235 40.715 125.735 ;
        RECT 40.885 125.405 41.055 125.905 ;
        RECT 41.315 125.955 41.565 127.325 ;
        RECT 42.915 127.155 43.245 127.515 ;
        RECT 41.855 126.965 43.245 127.155 ;
        RECT 44.075 127.325 44.635 127.615 ;
        RECT 44.805 127.325 45.055 127.785 ;
        RECT 41.855 126.875 42.025 126.965 ;
        RECT 41.735 126.545 42.025 126.875 ;
        RECT 42.195 126.545 42.535 126.795 ;
        RECT 42.755 126.545 43.430 126.795 ;
        RECT 41.855 126.295 42.025 126.545 ;
        RECT 41.855 126.125 42.795 126.295 ;
        RECT 43.165 126.185 43.430 126.545 ;
        RECT 41.315 125.405 41.775 125.955 ;
        RECT 41.965 125.235 42.295 125.955 ;
        RECT 42.495 125.575 42.795 126.125 ;
        RECT 44.075 125.955 44.325 127.325 ;
        RECT 45.675 127.155 46.005 127.515 ;
        RECT 44.615 126.965 46.005 127.155 ;
        RECT 46.575 127.155 46.905 127.515 ;
        RECT 47.525 127.325 47.775 127.785 ;
        RECT 47.945 127.325 48.505 127.615 ;
        RECT 46.575 126.965 47.965 127.155 ;
        RECT 44.615 126.875 44.785 126.965 ;
        RECT 44.495 126.545 44.785 126.875 ;
        RECT 47.795 126.875 47.965 126.965 ;
        RECT 44.955 126.545 45.295 126.795 ;
        RECT 45.515 126.545 46.190 126.795 ;
        RECT 44.615 126.295 44.785 126.545 ;
        RECT 44.615 126.125 45.555 126.295 ;
        RECT 45.925 126.185 46.190 126.545 ;
        RECT 46.390 126.545 47.065 126.795 ;
        RECT 47.285 126.545 47.625 126.795 ;
        RECT 47.795 126.545 48.085 126.875 ;
        RECT 46.390 126.185 46.655 126.545 ;
        RECT 47.795 126.295 47.965 126.545 ;
        RECT 42.965 125.235 43.245 125.905 ;
        RECT 44.075 125.405 44.535 125.955 ;
        RECT 44.725 125.235 45.055 125.955 ;
        RECT 45.255 125.575 45.555 126.125 ;
        RECT 47.025 126.125 47.965 126.295 ;
        RECT 45.725 125.235 46.005 125.905 ;
        RECT 46.575 125.235 46.855 125.905 ;
        RECT 47.025 125.575 47.325 126.125 ;
        RECT 48.255 125.955 48.505 127.325 ;
        RECT 48.675 127.060 48.965 127.785 ;
        RECT 49.695 127.320 49.945 127.785 ;
        RECT 50.115 127.145 50.285 127.615 ;
        RECT 50.535 127.325 50.705 127.785 ;
        RECT 50.955 127.145 51.125 127.615 ;
        RECT 51.375 127.325 51.545 127.785 ;
        RECT 51.795 127.145 51.965 127.615 ;
        RECT 52.335 127.325 52.600 127.785 ;
        RECT 49.595 126.965 51.965 127.145 ;
        RECT 52.815 127.015 55.405 127.785 ;
        RECT 55.665 127.235 55.835 127.615 ;
        RECT 56.015 127.405 56.345 127.785 ;
        RECT 55.665 127.065 56.330 127.235 ;
        RECT 56.525 127.110 56.785 127.615 ;
        RECT 57.330 127.445 57.585 127.605 ;
        RECT 57.245 127.275 57.585 127.445 ;
        RECT 57.765 127.325 58.050 127.785 ;
        RECT 47.525 125.235 47.855 125.955 ;
        RECT 48.045 125.405 48.505 125.955 ;
        RECT 48.675 125.235 48.965 126.400 ;
        RECT 49.595 126.375 49.945 126.965 ;
        RECT 50.115 126.545 52.625 126.795 ;
        RECT 49.595 126.205 52.045 126.375 ;
        RECT 49.595 126.185 50.365 126.205 ;
        RECT 49.695 125.235 49.865 125.695 ;
        RECT 50.035 125.405 50.365 126.185 ;
        RECT 50.535 125.235 50.705 126.035 ;
        RECT 50.875 125.405 51.205 126.205 ;
        RECT 51.375 125.235 51.545 126.035 ;
        RECT 51.715 125.405 52.045 126.205 ;
        RECT 52.305 125.235 52.600 126.375 ;
        RECT 52.815 126.325 54.025 126.845 ;
        RECT 54.195 126.495 55.405 127.015 ;
        RECT 55.595 126.515 55.925 126.885 ;
        RECT 56.160 126.810 56.330 127.065 ;
        RECT 56.160 126.480 56.445 126.810 ;
        RECT 56.160 126.335 56.330 126.480 ;
        RECT 52.815 125.235 55.405 126.325 ;
        RECT 55.665 126.165 56.330 126.335 ;
        RECT 56.615 126.310 56.785 127.110 ;
        RECT 55.665 125.405 55.835 126.165 ;
        RECT 56.015 125.235 56.345 125.995 ;
        RECT 56.515 125.405 56.785 126.310 ;
        RECT 57.330 127.075 57.585 127.275 ;
        RECT 57.330 126.215 57.510 127.075 ;
        RECT 58.230 126.875 58.480 127.525 ;
        RECT 57.680 126.545 58.480 126.875 ;
        RECT 57.330 125.545 57.585 126.215 ;
        RECT 57.765 125.235 58.050 126.035 ;
        RECT 58.230 125.955 58.480 126.545 ;
        RECT 58.680 127.190 59.000 127.520 ;
        RECT 59.180 127.305 59.840 127.785 ;
        RECT 60.040 127.395 60.890 127.565 ;
        RECT 58.680 126.295 58.870 127.190 ;
        RECT 59.190 126.865 59.850 127.135 ;
        RECT 59.520 126.805 59.850 126.865 ;
        RECT 59.040 126.635 59.370 126.695 ;
        RECT 60.040 126.635 60.210 127.395 ;
        RECT 61.450 127.325 61.770 127.785 ;
        RECT 61.970 127.145 62.220 127.575 ;
        RECT 62.510 127.345 62.920 127.785 ;
        RECT 63.090 127.405 64.105 127.605 ;
        RECT 60.380 126.975 61.630 127.145 ;
        RECT 60.380 126.855 60.710 126.975 ;
        RECT 59.040 126.465 60.940 126.635 ;
        RECT 58.680 126.125 60.600 126.295 ;
        RECT 58.680 126.105 59.000 126.125 ;
        RECT 58.230 125.445 58.560 125.955 ;
        RECT 58.830 125.495 59.000 126.105 ;
        RECT 60.770 125.955 60.940 126.465 ;
        RECT 61.110 126.395 61.290 126.805 ;
        RECT 61.460 126.215 61.630 126.975 ;
        RECT 59.170 125.235 59.500 125.925 ;
        RECT 59.730 125.785 60.940 125.955 ;
        RECT 61.110 125.905 61.630 126.215 ;
        RECT 61.800 126.805 62.220 127.145 ;
        RECT 62.510 126.805 62.920 127.135 ;
        RECT 61.800 126.035 61.990 126.805 ;
        RECT 63.090 126.675 63.260 127.405 ;
        RECT 64.405 127.235 64.575 127.565 ;
        RECT 64.745 127.405 65.075 127.785 ;
        RECT 63.430 126.855 63.780 127.225 ;
        RECT 63.090 126.635 63.510 126.675 ;
        RECT 62.160 126.465 63.510 126.635 ;
        RECT 62.160 126.305 62.410 126.465 ;
        RECT 62.920 126.035 63.170 126.295 ;
        RECT 61.800 125.785 63.170 126.035 ;
        RECT 59.730 125.495 59.970 125.785 ;
        RECT 60.770 125.705 60.940 125.785 ;
        RECT 60.170 125.235 60.590 125.615 ;
        RECT 60.770 125.455 61.400 125.705 ;
        RECT 61.870 125.235 62.200 125.615 ;
        RECT 62.370 125.495 62.540 125.785 ;
        RECT 63.340 125.620 63.510 126.465 ;
        RECT 63.960 126.295 64.180 127.165 ;
        RECT 64.405 127.045 65.100 127.235 ;
        RECT 63.680 125.915 64.180 126.295 ;
        RECT 64.350 126.245 64.760 126.865 ;
        RECT 64.930 126.075 65.100 127.045 ;
        RECT 64.405 125.905 65.100 126.075 ;
        RECT 62.720 125.235 63.100 125.615 ;
        RECT 63.340 125.450 64.170 125.620 ;
        RECT 64.405 125.405 64.575 125.905 ;
        RECT 64.745 125.235 65.075 125.735 ;
        RECT 65.290 125.405 65.515 127.525 ;
        RECT 65.685 127.405 66.015 127.785 ;
        RECT 66.185 127.235 66.355 127.525 ;
        RECT 65.690 127.065 66.355 127.235 ;
        RECT 65.690 126.075 65.920 127.065 ;
        RECT 66.615 127.035 67.825 127.785 ;
        RECT 66.090 126.245 66.440 126.895 ;
        RECT 66.615 126.325 67.135 126.865 ;
        RECT 67.305 126.495 67.825 127.035 ;
        RECT 67.995 127.110 68.255 127.615 ;
        RECT 68.435 127.405 68.765 127.785 ;
        RECT 68.945 127.235 69.115 127.615 ;
        RECT 65.690 125.905 66.355 126.075 ;
        RECT 65.685 125.235 66.015 125.735 ;
        RECT 66.185 125.405 66.355 125.905 ;
        RECT 66.615 125.235 67.825 126.325 ;
        RECT 67.995 126.310 68.165 127.110 ;
        RECT 68.450 127.065 69.115 127.235 ;
        RECT 68.450 126.810 68.620 127.065 ;
        RECT 69.380 127.045 69.635 127.615 ;
        RECT 69.805 127.385 70.135 127.785 ;
        RECT 70.560 127.250 71.090 127.615 ;
        RECT 70.560 127.215 70.735 127.250 ;
        RECT 69.805 127.045 70.735 127.215 ;
        RECT 68.335 126.480 68.620 126.810 ;
        RECT 68.855 126.515 69.185 126.885 ;
        RECT 68.450 126.335 68.620 126.480 ;
        RECT 69.380 126.375 69.550 127.045 ;
        RECT 69.805 126.875 69.975 127.045 ;
        RECT 69.720 126.545 69.975 126.875 ;
        RECT 70.200 126.545 70.395 126.875 ;
        RECT 67.995 125.405 68.265 126.310 ;
        RECT 68.450 126.165 69.115 126.335 ;
        RECT 68.435 125.235 68.765 125.995 ;
        RECT 68.945 125.405 69.115 126.165 ;
        RECT 69.380 125.405 69.715 126.375 ;
        RECT 69.885 125.235 70.055 126.375 ;
        RECT 70.225 125.575 70.395 126.545 ;
        RECT 70.565 125.915 70.735 127.045 ;
        RECT 70.905 126.255 71.075 127.055 ;
        RECT 71.280 126.765 71.555 127.615 ;
        RECT 71.275 126.595 71.555 126.765 ;
        RECT 71.280 126.455 71.555 126.595 ;
        RECT 71.725 126.255 71.915 127.615 ;
        RECT 72.095 127.250 72.605 127.785 ;
        RECT 72.825 126.975 73.070 127.580 ;
        RECT 74.435 127.060 74.725 127.785 ;
        RECT 74.895 127.325 75.455 127.615 ;
        RECT 75.625 127.325 75.875 127.785 ;
        RECT 72.115 126.805 73.345 126.975 ;
        RECT 70.905 126.085 71.915 126.255 ;
        RECT 72.085 126.240 72.835 126.430 ;
        RECT 70.565 125.745 71.690 125.915 ;
        RECT 72.085 125.575 72.255 126.240 ;
        RECT 73.005 125.995 73.345 126.805 ;
        RECT 70.225 125.405 72.255 125.575 ;
        RECT 72.425 125.235 72.595 125.995 ;
        RECT 72.830 125.585 73.345 125.995 ;
        RECT 74.435 125.235 74.725 126.400 ;
        RECT 74.895 125.955 75.145 127.325 ;
        RECT 76.495 127.155 76.825 127.515 ;
        RECT 75.435 126.965 76.825 127.155 ;
        RECT 77.235 126.965 77.465 127.785 ;
        RECT 77.635 126.985 77.965 127.615 ;
        RECT 75.435 126.875 75.605 126.965 ;
        RECT 75.315 126.545 75.605 126.875 ;
        RECT 75.775 126.545 76.115 126.795 ;
        RECT 76.335 126.545 77.010 126.795 ;
        RECT 77.215 126.545 77.545 126.795 ;
        RECT 75.435 126.295 75.605 126.545 ;
        RECT 75.435 126.125 76.375 126.295 ;
        RECT 76.745 126.185 77.010 126.545 ;
        RECT 77.715 126.385 77.965 126.985 ;
        RECT 78.135 126.965 78.345 127.785 ;
        RECT 78.575 127.015 81.165 127.785 ;
        RECT 81.340 127.240 86.685 127.785 ;
        RECT 74.895 125.405 75.355 125.955 ;
        RECT 75.545 125.235 75.875 125.955 ;
        RECT 76.075 125.575 76.375 126.125 ;
        RECT 76.545 125.235 76.825 125.905 ;
        RECT 77.235 125.235 77.465 126.375 ;
        RECT 77.635 125.405 77.965 126.385 ;
        RECT 78.135 125.235 78.345 126.375 ;
        RECT 78.575 126.325 79.785 126.845 ;
        RECT 79.955 126.495 81.165 127.015 ;
        RECT 78.575 125.235 81.165 126.325 ;
        RECT 82.930 125.670 83.280 126.920 ;
        RECT 84.760 126.410 85.100 127.240 ;
        RECT 86.895 126.965 87.125 127.785 ;
        RECT 87.295 126.985 87.625 127.615 ;
        RECT 86.875 126.545 87.205 126.795 ;
        RECT 87.375 126.385 87.625 126.985 ;
        RECT 87.795 126.965 88.005 127.785 ;
        RECT 89.430 126.975 89.675 127.580 ;
        RECT 89.895 127.250 90.405 127.785 ;
        RECT 81.340 125.235 86.685 125.670 ;
        RECT 86.895 125.235 87.125 126.375 ;
        RECT 87.295 125.405 87.625 126.385 ;
        RECT 89.155 126.805 90.385 126.975 ;
        RECT 87.795 125.235 88.005 126.375 ;
        RECT 89.155 125.995 89.495 126.805 ;
        RECT 89.665 126.240 90.415 126.430 ;
        RECT 89.155 125.585 89.670 125.995 ;
        RECT 89.905 125.235 90.075 125.995 ;
        RECT 90.245 125.575 90.415 126.240 ;
        RECT 90.585 126.255 90.775 127.615 ;
        RECT 90.945 126.765 91.220 127.615 ;
        RECT 91.410 127.250 91.940 127.615 ;
        RECT 92.365 127.385 92.695 127.785 ;
        RECT 91.765 127.215 91.940 127.250 ;
        RECT 90.945 126.595 91.225 126.765 ;
        RECT 90.945 126.455 91.220 126.595 ;
        RECT 91.425 126.255 91.595 127.055 ;
        RECT 90.585 126.085 91.595 126.255 ;
        RECT 91.765 127.045 92.695 127.215 ;
        RECT 92.865 127.045 93.120 127.615 ;
        RECT 91.765 125.915 91.935 127.045 ;
        RECT 92.525 126.875 92.695 127.045 ;
        RECT 90.810 125.745 91.935 125.915 ;
        RECT 92.105 126.545 92.300 126.875 ;
        RECT 92.525 126.545 92.780 126.875 ;
        RECT 92.105 125.575 92.275 126.545 ;
        RECT 92.950 126.375 93.120 127.045 ;
        RECT 93.335 126.965 93.565 127.785 ;
        RECT 93.735 126.985 94.065 127.615 ;
        RECT 93.315 126.545 93.645 126.795 ;
        RECT 93.815 126.385 94.065 126.985 ;
        RECT 94.235 126.965 94.445 127.785 ;
        RECT 94.950 126.975 95.195 127.580 ;
        RECT 95.415 127.250 95.925 127.785 ;
        RECT 90.245 125.405 92.275 125.575 ;
        RECT 92.445 125.235 92.615 126.375 ;
        RECT 92.785 125.405 93.120 126.375 ;
        RECT 93.335 125.235 93.565 126.375 ;
        RECT 93.735 125.405 94.065 126.385 ;
        RECT 94.675 126.805 95.905 126.975 ;
        RECT 94.235 125.235 94.445 126.375 ;
        RECT 94.675 125.995 95.015 126.805 ;
        RECT 95.185 126.240 95.935 126.430 ;
        RECT 94.675 125.585 95.190 125.995 ;
        RECT 95.425 125.235 95.595 125.995 ;
        RECT 95.765 125.575 95.935 126.240 ;
        RECT 96.105 126.255 96.295 127.615 ;
        RECT 96.465 126.765 96.740 127.615 ;
        RECT 96.930 127.250 97.460 127.615 ;
        RECT 97.885 127.385 98.215 127.785 ;
        RECT 97.285 127.215 97.460 127.250 ;
        RECT 96.465 126.595 96.745 126.765 ;
        RECT 96.465 126.455 96.740 126.595 ;
        RECT 96.945 126.255 97.115 127.055 ;
        RECT 96.105 126.085 97.115 126.255 ;
        RECT 97.285 127.045 98.215 127.215 ;
        RECT 98.385 127.045 98.640 127.615 ;
        RECT 97.285 125.915 97.455 127.045 ;
        RECT 98.045 126.875 98.215 127.045 ;
        RECT 96.330 125.745 97.455 125.915 ;
        RECT 97.625 126.545 97.820 126.875 ;
        RECT 98.045 126.545 98.300 126.875 ;
        RECT 97.625 125.575 97.795 126.545 ;
        RECT 98.470 126.375 98.640 127.045 ;
        RECT 98.855 126.965 99.085 127.785 ;
        RECT 99.255 126.985 99.585 127.615 ;
        RECT 98.835 126.545 99.165 126.795 ;
        RECT 99.335 126.385 99.585 126.985 ;
        RECT 99.755 126.965 99.965 127.785 ;
        RECT 100.195 127.060 100.485 127.785 ;
        RECT 100.695 126.965 100.925 127.785 ;
        RECT 101.095 126.985 101.425 127.615 ;
        RECT 100.675 126.545 101.005 126.795 ;
        RECT 95.765 125.405 97.795 125.575 ;
        RECT 97.965 125.235 98.135 126.375 ;
        RECT 98.305 125.405 98.640 126.375 ;
        RECT 98.855 125.235 99.085 126.375 ;
        RECT 99.255 125.405 99.585 126.385 ;
        RECT 99.755 125.235 99.965 126.375 ;
        RECT 100.195 125.235 100.485 126.400 ;
        RECT 101.175 126.385 101.425 126.985 ;
        RECT 101.595 126.965 101.805 127.785 ;
        RECT 102.410 127.445 102.665 127.605 ;
        RECT 102.325 127.275 102.665 127.445 ;
        RECT 102.845 127.325 103.130 127.785 ;
        RECT 102.410 127.075 102.665 127.275 ;
        RECT 100.695 125.235 100.925 126.375 ;
        RECT 101.095 125.405 101.425 126.385 ;
        RECT 101.595 125.235 101.805 126.375 ;
        RECT 102.410 126.215 102.590 127.075 ;
        RECT 103.310 126.875 103.560 127.525 ;
        RECT 102.760 126.545 103.560 126.875 ;
        RECT 102.410 125.545 102.665 126.215 ;
        RECT 102.845 125.235 103.130 126.035 ;
        RECT 103.310 125.955 103.560 126.545 ;
        RECT 103.760 127.190 104.080 127.520 ;
        RECT 104.260 127.305 104.920 127.785 ;
        RECT 105.120 127.395 105.970 127.565 ;
        RECT 103.760 126.295 103.950 127.190 ;
        RECT 104.270 126.865 104.930 127.135 ;
        RECT 104.600 126.805 104.930 126.865 ;
        RECT 104.120 126.635 104.450 126.695 ;
        RECT 105.120 126.635 105.290 127.395 ;
        RECT 106.530 127.325 106.850 127.785 ;
        RECT 107.050 127.145 107.300 127.575 ;
        RECT 107.590 127.345 108.000 127.785 ;
        RECT 108.170 127.405 109.185 127.605 ;
        RECT 105.460 126.975 106.710 127.145 ;
        RECT 105.460 126.855 105.790 126.975 ;
        RECT 104.120 126.465 106.020 126.635 ;
        RECT 103.760 126.125 105.680 126.295 ;
        RECT 103.760 126.105 104.080 126.125 ;
        RECT 103.310 125.445 103.640 125.955 ;
        RECT 103.910 125.495 104.080 126.105 ;
        RECT 105.850 125.955 106.020 126.465 ;
        RECT 106.190 126.395 106.370 126.805 ;
        RECT 106.540 126.215 106.710 126.975 ;
        RECT 104.250 125.235 104.580 125.925 ;
        RECT 104.810 125.785 106.020 125.955 ;
        RECT 106.190 125.905 106.710 126.215 ;
        RECT 106.880 126.805 107.300 127.145 ;
        RECT 107.590 126.805 108.000 127.135 ;
        RECT 106.880 126.035 107.070 126.805 ;
        RECT 108.170 126.675 108.340 127.405 ;
        RECT 109.485 127.235 109.655 127.565 ;
        RECT 109.825 127.405 110.155 127.785 ;
        RECT 108.510 126.855 108.860 127.225 ;
        RECT 108.170 126.635 108.590 126.675 ;
        RECT 107.240 126.465 108.590 126.635 ;
        RECT 107.240 126.305 107.490 126.465 ;
        RECT 108.000 126.035 108.250 126.295 ;
        RECT 106.880 125.785 108.250 126.035 ;
        RECT 104.810 125.495 105.050 125.785 ;
        RECT 105.850 125.705 106.020 125.785 ;
        RECT 105.250 125.235 105.670 125.615 ;
        RECT 105.850 125.455 106.480 125.705 ;
        RECT 106.950 125.235 107.280 125.615 ;
        RECT 107.450 125.495 107.620 125.785 ;
        RECT 108.420 125.620 108.590 126.465 ;
        RECT 109.040 126.295 109.260 127.165 ;
        RECT 109.485 127.045 110.180 127.235 ;
        RECT 108.760 125.915 109.260 126.295 ;
        RECT 109.430 126.245 109.840 126.865 ;
        RECT 110.010 126.075 110.180 127.045 ;
        RECT 109.485 125.905 110.180 126.075 ;
        RECT 107.800 125.235 108.180 125.615 ;
        RECT 108.420 125.450 109.250 125.620 ;
        RECT 109.485 125.405 109.655 125.905 ;
        RECT 109.825 125.235 110.155 125.735 ;
        RECT 110.370 125.405 110.595 127.525 ;
        RECT 110.765 127.405 111.095 127.785 ;
        RECT 111.265 127.235 111.435 127.525 ;
        RECT 110.770 127.065 111.435 127.235 ;
        RECT 110.770 126.075 111.000 127.065 ;
        RECT 112.155 127.035 113.365 127.785 ;
        RECT 111.170 126.245 111.520 126.895 ;
        RECT 112.155 126.325 112.675 126.865 ;
        RECT 112.845 126.495 113.365 127.035 ;
        RECT 110.770 125.905 111.435 126.075 ;
        RECT 110.765 125.235 111.095 125.735 ;
        RECT 111.265 125.405 111.435 125.905 ;
        RECT 112.155 125.235 113.365 126.325 ;
        RECT 15.010 125.065 113.450 125.235 ;
        RECT 15.095 123.975 16.305 125.065 ;
        RECT 15.095 123.265 15.615 123.805 ;
        RECT 15.785 123.435 16.305 123.975 ;
        RECT 16.935 123.975 18.605 125.065 ;
        RECT 16.935 123.455 17.685 123.975 ;
        RECT 18.835 123.925 19.045 125.065 ;
        RECT 19.215 123.915 19.545 124.895 ;
        RECT 19.715 123.925 19.945 125.065 ;
        RECT 20.530 124.725 20.785 124.755 ;
        RECT 20.445 124.555 20.785 124.725 ;
        RECT 20.530 124.085 20.785 124.555 ;
        RECT 20.965 124.265 21.250 125.065 ;
        RECT 21.430 124.345 21.760 124.855 ;
        RECT 17.855 123.285 18.605 123.805 ;
        RECT 15.095 122.515 16.305 123.265 ;
        RECT 16.935 122.515 18.605 123.285 ;
        RECT 18.835 122.515 19.045 123.335 ;
        RECT 19.215 123.315 19.465 123.915 ;
        RECT 19.635 123.505 19.965 123.755 ;
        RECT 19.215 122.685 19.545 123.315 ;
        RECT 19.715 122.515 19.945 123.335 ;
        RECT 20.530 123.225 20.710 124.085 ;
        RECT 21.430 123.755 21.680 124.345 ;
        RECT 22.030 124.195 22.200 124.805 ;
        RECT 22.370 124.375 22.700 125.065 ;
        RECT 22.930 124.515 23.170 124.805 ;
        RECT 23.370 124.685 23.790 125.065 ;
        RECT 23.970 124.595 24.600 124.845 ;
        RECT 25.070 124.685 25.400 125.065 ;
        RECT 23.970 124.515 24.140 124.595 ;
        RECT 25.570 124.515 25.740 124.805 ;
        RECT 25.920 124.685 26.300 125.065 ;
        RECT 26.540 124.680 27.370 124.850 ;
        RECT 22.930 124.345 24.140 124.515 ;
        RECT 20.880 123.425 21.680 123.755 ;
        RECT 20.530 122.695 20.785 123.225 ;
        RECT 20.965 122.515 21.250 122.975 ;
        RECT 21.430 122.775 21.680 123.425 ;
        RECT 21.880 124.175 22.200 124.195 ;
        RECT 21.880 124.005 23.800 124.175 ;
        RECT 21.880 123.110 22.070 124.005 ;
        RECT 23.970 123.835 24.140 124.345 ;
        RECT 24.310 124.085 24.830 124.395 ;
        RECT 22.240 123.665 24.140 123.835 ;
        RECT 22.240 123.605 22.570 123.665 ;
        RECT 22.720 123.435 23.050 123.495 ;
        RECT 22.390 123.165 23.050 123.435 ;
        RECT 21.880 122.780 22.200 123.110 ;
        RECT 22.380 122.515 23.040 122.995 ;
        RECT 23.240 122.905 23.410 123.665 ;
        RECT 24.310 123.495 24.490 123.905 ;
        RECT 23.580 123.325 23.910 123.445 ;
        RECT 24.660 123.325 24.830 124.085 ;
        RECT 23.580 123.155 24.830 123.325 ;
        RECT 25.000 124.265 26.370 124.515 ;
        RECT 25.000 123.495 25.190 124.265 ;
        RECT 26.120 124.005 26.370 124.265 ;
        RECT 25.360 123.835 25.610 123.995 ;
        RECT 26.540 123.835 26.710 124.680 ;
        RECT 27.605 124.395 27.775 124.895 ;
        RECT 27.945 124.565 28.275 125.065 ;
        RECT 26.880 124.005 27.380 124.385 ;
        RECT 27.605 124.225 28.300 124.395 ;
        RECT 25.360 123.665 26.710 123.835 ;
        RECT 26.290 123.625 26.710 123.665 ;
        RECT 25.000 123.155 25.420 123.495 ;
        RECT 25.710 123.165 26.120 123.495 ;
        RECT 23.240 122.735 24.090 122.905 ;
        RECT 24.650 122.515 24.970 122.975 ;
        RECT 25.170 122.725 25.420 123.155 ;
        RECT 25.710 122.515 26.120 122.955 ;
        RECT 26.290 122.895 26.460 123.625 ;
        RECT 26.630 123.075 26.980 123.445 ;
        RECT 27.160 123.135 27.380 124.005 ;
        RECT 27.550 123.435 27.960 124.055 ;
        RECT 28.130 123.255 28.300 124.225 ;
        RECT 27.605 123.065 28.300 123.255 ;
        RECT 26.290 122.695 27.305 122.895 ;
        RECT 27.605 122.735 27.775 123.065 ;
        RECT 27.945 122.515 28.275 122.895 ;
        RECT 28.490 122.775 28.715 124.895 ;
        RECT 28.885 124.565 29.215 125.065 ;
        RECT 29.385 124.395 29.555 124.895 ;
        RECT 28.890 124.225 29.555 124.395 ;
        RECT 30.275 124.305 30.790 124.715 ;
        RECT 31.025 124.305 31.195 125.065 ;
        RECT 31.365 124.725 33.395 124.895 ;
        RECT 28.890 123.235 29.120 124.225 ;
        RECT 29.290 123.405 29.640 124.055 ;
        RECT 30.275 123.495 30.615 124.305 ;
        RECT 31.365 124.060 31.535 124.725 ;
        RECT 31.930 124.385 33.055 124.555 ;
        RECT 30.785 123.870 31.535 124.060 ;
        RECT 31.705 124.045 32.715 124.215 ;
        RECT 30.275 123.325 31.505 123.495 ;
        RECT 28.890 123.065 29.555 123.235 ;
        RECT 28.885 122.515 29.215 122.895 ;
        RECT 29.385 122.775 29.555 123.065 ;
        RECT 30.550 122.720 30.795 123.325 ;
        RECT 31.015 122.515 31.525 123.050 ;
        RECT 31.705 122.685 31.895 124.045 ;
        RECT 32.065 123.025 32.340 123.845 ;
        RECT 32.545 123.245 32.715 124.045 ;
        RECT 32.885 123.255 33.055 124.385 ;
        RECT 33.225 123.755 33.395 124.725 ;
        RECT 33.565 123.925 33.735 125.065 ;
        RECT 33.905 123.925 34.240 124.895 ;
        RECT 33.225 123.425 33.420 123.755 ;
        RECT 33.645 123.425 33.900 123.755 ;
        RECT 33.645 123.255 33.815 123.425 ;
        RECT 34.070 123.255 34.240 123.925 ;
        RECT 34.415 123.975 35.625 125.065 ;
        RECT 34.415 123.435 34.935 123.975 ;
        RECT 35.795 123.900 36.085 125.065 ;
        RECT 36.255 123.975 37.925 125.065 ;
        RECT 38.185 124.135 38.355 124.895 ;
        RECT 38.535 124.305 38.865 125.065 ;
        RECT 35.105 123.265 35.625 123.805 ;
        RECT 36.255 123.455 37.005 123.975 ;
        RECT 38.185 123.965 38.850 124.135 ;
        RECT 39.035 123.990 39.305 124.895 ;
        RECT 39.675 124.395 39.955 125.065 ;
        RECT 40.125 124.175 40.425 124.725 ;
        RECT 40.625 124.345 40.955 125.065 ;
        RECT 41.145 124.345 41.605 124.895 ;
        RECT 38.680 123.820 38.850 123.965 ;
        RECT 37.175 123.285 37.925 123.805 ;
        RECT 38.115 123.415 38.445 123.785 ;
        RECT 38.680 123.490 38.965 123.820 ;
        RECT 32.885 123.085 33.815 123.255 ;
        RECT 32.885 123.050 33.060 123.085 ;
        RECT 32.065 122.855 32.345 123.025 ;
        RECT 32.065 122.685 32.340 122.855 ;
        RECT 32.530 122.685 33.060 123.050 ;
        RECT 33.485 122.515 33.815 122.915 ;
        RECT 33.985 122.685 34.240 123.255 ;
        RECT 34.415 122.515 35.625 123.265 ;
        RECT 35.795 122.515 36.085 123.240 ;
        RECT 36.255 122.515 37.925 123.285 ;
        RECT 38.680 123.235 38.850 123.490 ;
        RECT 38.185 123.065 38.850 123.235 ;
        RECT 39.135 123.190 39.305 123.990 ;
        RECT 39.490 123.755 39.755 124.115 ;
        RECT 40.125 124.005 41.065 124.175 ;
        RECT 40.895 123.755 41.065 124.005 ;
        RECT 39.490 123.505 40.165 123.755 ;
        RECT 40.385 123.505 40.725 123.755 ;
        RECT 40.895 123.425 41.185 123.755 ;
        RECT 40.895 123.335 41.065 123.425 ;
        RECT 38.185 122.685 38.355 123.065 ;
        RECT 38.535 122.515 38.865 122.895 ;
        RECT 39.045 122.685 39.305 123.190 ;
        RECT 39.675 123.145 41.065 123.335 ;
        RECT 39.675 122.785 40.005 123.145 ;
        RECT 41.355 122.975 41.605 124.345 ;
        RECT 40.625 122.515 40.875 122.975 ;
        RECT 41.045 122.685 41.605 122.975 ;
        RECT 41.780 123.925 42.115 124.895 ;
        RECT 42.285 123.925 42.455 125.065 ;
        RECT 42.625 124.725 44.655 124.895 ;
        RECT 41.780 123.255 41.950 123.925 ;
        RECT 42.625 123.755 42.795 124.725 ;
        RECT 42.120 123.425 42.375 123.755 ;
        RECT 42.600 123.425 42.795 123.755 ;
        RECT 42.965 124.385 44.090 124.555 ;
        RECT 42.205 123.255 42.375 123.425 ;
        RECT 42.965 123.255 43.135 124.385 ;
        RECT 41.780 122.685 42.035 123.255 ;
        RECT 42.205 123.085 43.135 123.255 ;
        RECT 43.305 124.045 44.315 124.215 ;
        RECT 43.305 123.245 43.475 124.045 ;
        RECT 43.680 123.365 43.955 123.845 ;
        RECT 43.675 123.195 43.955 123.365 ;
        RECT 42.960 123.050 43.135 123.085 ;
        RECT 42.205 122.515 42.535 122.915 ;
        RECT 42.960 122.685 43.490 123.050 ;
        RECT 43.680 122.685 43.955 123.195 ;
        RECT 44.125 122.685 44.315 124.045 ;
        RECT 44.485 124.060 44.655 124.725 ;
        RECT 44.825 124.305 44.995 125.065 ;
        RECT 45.230 124.305 45.745 124.715 ;
        RECT 44.485 123.870 45.235 124.060 ;
        RECT 45.405 123.495 45.745 124.305 ;
        RECT 44.515 123.325 45.745 123.495 ;
        RECT 45.915 124.305 46.430 124.715 ;
        RECT 46.665 124.305 46.835 125.065 ;
        RECT 47.005 124.725 49.035 124.895 ;
        RECT 45.915 123.495 46.255 124.305 ;
        RECT 47.005 124.060 47.175 124.725 ;
        RECT 47.570 124.385 48.695 124.555 ;
        RECT 46.425 123.870 47.175 124.060 ;
        RECT 47.345 124.045 48.355 124.215 ;
        RECT 45.915 123.325 47.145 123.495 ;
        RECT 44.495 122.515 45.005 123.050 ;
        RECT 45.225 122.720 45.470 123.325 ;
        RECT 46.190 122.720 46.435 123.325 ;
        RECT 46.655 122.515 47.165 123.050 ;
        RECT 47.345 122.685 47.535 124.045 ;
        RECT 47.705 123.365 47.980 123.845 ;
        RECT 47.705 123.195 47.985 123.365 ;
        RECT 48.185 123.245 48.355 124.045 ;
        RECT 48.525 123.255 48.695 124.385 ;
        RECT 48.865 123.755 49.035 124.725 ;
        RECT 49.205 123.925 49.375 125.065 ;
        RECT 49.545 123.925 49.880 124.895 ;
        RECT 48.865 123.425 49.060 123.755 ;
        RECT 49.285 123.425 49.540 123.755 ;
        RECT 49.285 123.255 49.455 123.425 ;
        RECT 49.710 123.255 49.880 123.925 ;
        RECT 50.055 123.975 51.725 125.065 ;
        RECT 52.270 124.725 52.525 124.755 ;
        RECT 52.185 124.555 52.525 124.725 ;
        RECT 52.270 124.085 52.525 124.555 ;
        RECT 52.705 124.265 52.990 125.065 ;
        RECT 53.170 124.345 53.500 124.855 ;
        RECT 50.055 123.455 50.805 123.975 ;
        RECT 50.975 123.285 51.725 123.805 ;
        RECT 47.705 122.685 47.980 123.195 ;
        RECT 48.525 123.085 49.455 123.255 ;
        RECT 48.525 123.050 48.700 123.085 ;
        RECT 48.170 122.685 48.700 123.050 ;
        RECT 49.125 122.515 49.455 122.915 ;
        RECT 49.625 122.685 49.880 123.255 ;
        RECT 50.055 122.515 51.725 123.285 ;
        RECT 52.270 123.225 52.450 124.085 ;
        RECT 53.170 123.755 53.420 124.345 ;
        RECT 53.770 124.195 53.940 124.805 ;
        RECT 54.110 124.375 54.440 125.065 ;
        RECT 54.670 124.515 54.910 124.805 ;
        RECT 55.110 124.685 55.530 125.065 ;
        RECT 55.710 124.595 56.340 124.845 ;
        RECT 56.810 124.685 57.140 125.065 ;
        RECT 55.710 124.515 55.880 124.595 ;
        RECT 57.310 124.515 57.480 124.805 ;
        RECT 57.660 124.685 58.040 125.065 ;
        RECT 58.280 124.680 59.110 124.850 ;
        RECT 54.670 124.345 55.880 124.515 ;
        RECT 52.620 123.425 53.420 123.755 ;
        RECT 52.270 122.695 52.525 123.225 ;
        RECT 52.705 122.515 52.990 122.975 ;
        RECT 53.170 122.775 53.420 123.425 ;
        RECT 53.620 124.175 53.940 124.195 ;
        RECT 53.620 124.005 55.540 124.175 ;
        RECT 53.620 123.110 53.810 124.005 ;
        RECT 55.710 123.835 55.880 124.345 ;
        RECT 56.050 124.085 56.570 124.395 ;
        RECT 53.980 123.665 55.880 123.835 ;
        RECT 53.980 123.605 54.310 123.665 ;
        RECT 54.460 123.435 54.790 123.495 ;
        RECT 54.130 123.165 54.790 123.435 ;
        RECT 53.620 122.780 53.940 123.110 ;
        RECT 54.120 122.515 54.780 122.995 ;
        RECT 54.980 122.905 55.150 123.665 ;
        RECT 56.050 123.495 56.230 123.905 ;
        RECT 55.320 123.325 55.650 123.445 ;
        RECT 56.400 123.325 56.570 124.085 ;
        RECT 55.320 123.155 56.570 123.325 ;
        RECT 56.740 124.265 58.110 124.515 ;
        RECT 56.740 123.495 56.930 124.265 ;
        RECT 57.860 124.005 58.110 124.265 ;
        RECT 57.100 123.835 57.350 123.995 ;
        RECT 58.280 123.835 58.450 124.680 ;
        RECT 59.345 124.395 59.515 124.895 ;
        RECT 59.685 124.565 60.015 125.065 ;
        RECT 58.620 124.005 59.120 124.385 ;
        RECT 59.345 124.225 60.040 124.395 ;
        RECT 57.100 123.665 58.450 123.835 ;
        RECT 58.030 123.625 58.450 123.665 ;
        RECT 56.740 123.155 57.160 123.495 ;
        RECT 57.450 123.165 57.860 123.495 ;
        RECT 54.980 122.735 55.830 122.905 ;
        RECT 56.390 122.515 56.710 122.975 ;
        RECT 56.910 122.725 57.160 123.155 ;
        RECT 57.450 122.515 57.860 122.955 ;
        RECT 58.030 122.895 58.200 123.625 ;
        RECT 58.370 123.075 58.720 123.445 ;
        RECT 58.900 123.135 59.120 124.005 ;
        RECT 59.290 123.435 59.700 124.055 ;
        RECT 59.870 123.255 60.040 124.225 ;
        RECT 59.345 123.065 60.040 123.255 ;
        RECT 58.030 122.695 59.045 122.895 ;
        RECT 59.345 122.735 59.515 123.065 ;
        RECT 59.685 122.515 60.015 122.895 ;
        RECT 60.230 122.775 60.455 124.895 ;
        RECT 60.625 124.565 60.955 125.065 ;
        RECT 61.125 124.395 61.295 124.895 ;
        RECT 60.630 124.225 61.295 124.395 ;
        RECT 60.630 123.235 60.860 124.225 ;
        RECT 61.030 123.405 61.380 124.055 ;
        RECT 61.555 123.900 61.845 125.065 ;
        RECT 62.075 123.925 62.285 125.065 ;
        RECT 62.455 123.915 62.785 124.895 ;
        RECT 62.955 123.925 63.185 125.065 ;
        RECT 63.485 124.135 63.655 124.895 ;
        RECT 63.835 124.305 64.165 125.065 ;
        RECT 63.485 123.965 64.150 124.135 ;
        RECT 64.335 123.990 64.605 124.895 ;
        RECT 60.630 123.065 61.295 123.235 ;
        RECT 60.625 122.515 60.955 122.895 ;
        RECT 61.125 122.775 61.295 123.065 ;
        RECT 61.555 122.515 61.845 123.240 ;
        RECT 62.075 122.515 62.285 123.335 ;
        RECT 62.455 123.315 62.705 123.915 ;
        RECT 63.980 123.820 64.150 123.965 ;
        RECT 62.875 123.505 63.205 123.755 ;
        RECT 63.415 123.415 63.745 123.785 ;
        RECT 63.980 123.490 64.265 123.820 ;
        RECT 62.455 122.685 62.785 123.315 ;
        RECT 62.955 122.515 63.185 123.335 ;
        RECT 63.980 123.235 64.150 123.490 ;
        RECT 63.485 123.065 64.150 123.235 ;
        RECT 64.435 123.190 64.605 123.990 ;
        RECT 64.775 123.975 66.445 125.065 ;
        RECT 64.775 123.455 65.525 123.975 ;
        RECT 66.655 123.925 66.885 125.065 ;
        RECT 67.055 123.915 67.385 124.895 ;
        RECT 67.555 123.925 67.765 125.065 ;
        RECT 68.370 124.725 68.625 124.755 ;
        RECT 68.285 124.555 68.625 124.725 ;
        RECT 68.370 124.085 68.625 124.555 ;
        RECT 68.805 124.265 69.090 125.065 ;
        RECT 69.270 124.345 69.600 124.855 ;
        RECT 65.695 123.285 66.445 123.805 ;
        RECT 66.635 123.505 66.965 123.755 ;
        RECT 63.485 122.685 63.655 123.065 ;
        RECT 63.835 122.515 64.165 122.895 ;
        RECT 64.345 122.685 64.605 123.190 ;
        RECT 64.775 122.515 66.445 123.285 ;
        RECT 66.655 122.515 66.885 123.335 ;
        RECT 67.135 123.315 67.385 123.915 ;
        RECT 67.055 122.685 67.385 123.315 ;
        RECT 67.555 122.515 67.765 123.335 ;
        RECT 68.370 123.225 68.550 124.085 ;
        RECT 69.270 123.755 69.520 124.345 ;
        RECT 69.870 124.195 70.040 124.805 ;
        RECT 70.210 124.375 70.540 125.065 ;
        RECT 70.770 124.515 71.010 124.805 ;
        RECT 71.210 124.685 71.630 125.065 ;
        RECT 71.810 124.595 72.440 124.845 ;
        RECT 72.910 124.685 73.240 125.065 ;
        RECT 71.810 124.515 71.980 124.595 ;
        RECT 73.410 124.515 73.580 124.805 ;
        RECT 73.760 124.685 74.140 125.065 ;
        RECT 74.380 124.680 75.210 124.850 ;
        RECT 70.770 124.345 71.980 124.515 ;
        RECT 68.720 123.425 69.520 123.755 ;
        RECT 68.370 122.695 68.625 123.225 ;
        RECT 68.805 122.515 69.090 122.975 ;
        RECT 69.270 122.775 69.520 123.425 ;
        RECT 69.720 124.175 70.040 124.195 ;
        RECT 69.720 124.005 71.640 124.175 ;
        RECT 69.720 123.110 69.910 124.005 ;
        RECT 71.810 123.835 71.980 124.345 ;
        RECT 72.150 124.085 72.670 124.395 ;
        RECT 70.080 123.665 71.980 123.835 ;
        RECT 70.080 123.605 70.410 123.665 ;
        RECT 70.560 123.435 70.890 123.495 ;
        RECT 70.230 123.165 70.890 123.435 ;
        RECT 69.720 122.780 70.040 123.110 ;
        RECT 70.220 122.515 70.880 122.995 ;
        RECT 71.080 122.905 71.250 123.665 ;
        RECT 72.150 123.495 72.330 123.905 ;
        RECT 71.420 123.325 71.750 123.445 ;
        RECT 72.500 123.325 72.670 124.085 ;
        RECT 71.420 123.155 72.670 123.325 ;
        RECT 72.840 124.265 74.210 124.515 ;
        RECT 72.840 123.495 73.030 124.265 ;
        RECT 73.960 124.005 74.210 124.265 ;
        RECT 73.200 123.835 73.450 123.995 ;
        RECT 74.380 123.835 74.550 124.680 ;
        RECT 75.445 124.395 75.615 124.895 ;
        RECT 75.785 124.565 76.115 125.065 ;
        RECT 74.720 124.005 75.220 124.385 ;
        RECT 75.445 124.225 76.140 124.395 ;
        RECT 73.200 123.665 74.550 123.835 ;
        RECT 74.130 123.625 74.550 123.665 ;
        RECT 72.840 123.155 73.260 123.495 ;
        RECT 73.550 123.165 73.960 123.495 ;
        RECT 71.080 122.735 71.930 122.905 ;
        RECT 72.490 122.515 72.810 122.975 ;
        RECT 73.010 122.725 73.260 123.155 ;
        RECT 73.550 122.515 73.960 122.955 ;
        RECT 74.130 122.895 74.300 123.625 ;
        RECT 74.470 123.075 74.820 123.445 ;
        RECT 75.000 123.135 75.220 124.005 ;
        RECT 75.390 123.435 75.800 124.055 ;
        RECT 75.970 123.255 76.140 124.225 ;
        RECT 75.445 123.065 76.140 123.255 ;
        RECT 74.130 122.695 75.145 122.895 ;
        RECT 75.445 122.735 75.615 123.065 ;
        RECT 75.785 122.515 76.115 122.895 ;
        RECT 76.330 122.775 76.555 124.895 ;
        RECT 76.725 124.565 77.055 125.065 ;
        RECT 77.225 124.395 77.395 124.895 ;
        RECT 76.730 124.225 77.395 124.395 ;
        RECT 76.730 123.235 76.960 124.225 ;
        RECT 77.130 123.405 77.480 124.055 ;
        RECT 77.655 123.975 81.165 125.065 ;
        RECT 81.335 124.305 81.850 124.715 ;
        RECT 82.085 124.305 82.255 125.065 ;
        RECT 82.425 124.725 84.455 124.895 ;
        RECT 77.655 123.455 79.345 123.975 ;
        RECT 79.515 123.285 81.165 123.805 ;
        RECT 81.335 123.495 81.675 124.305 ;
        RECT 82.425 124.060 82.595 124.725 ;
        RECT 82.990 124.385 84.115 124.555 ;
        RECT 81.845 123.870 82.595 124.060 ;
        RECT 82.765 124.045 83.775 124.215 ;
        RECT 81.335 123.325 82.565 123.495 ;
        RECT 76.730 123.065 77.395 123.235 ;
        RECT 76.725 122.515 77.055 122.895 ;
        RECT 77.225 122.775 77.395 123.065 ;
        RECT 77.655 122.515 81.165 123.285 ;
        RECT 81.610 122.720 81.855 123.325 ;
        RECT 82.075 122.515 82.585 123.050 ;
        RECT 82.765 122.685 82.955 124.045 ;
        RECT 83.125 123.025 83.400 123.845 ;
        RECT 83.605 123.245 83.775 124.045 ;
        RECT 83.945 123.255 84.115 124.385 ;
        RECT 84.285 123.755 84.455 124.725 ;
        RECT 84.625 123.925 84.795 125.065 ;
        RECT 84.965 123.925 85.300 124.895 ;
        RECT 84.285 123.425 84.480 123.755 ;
        RECT 84.705 123.425 84.960 123.755 ;
        RECT 84.705 123.255 84.875 123.425 ;
        RECT 85.130 123.255 85.300 123.925 ;
        RECT 85.475 123.975 87.145 125.065 ;
        RECT 85.475 123.455 86.225 123.975 ;
        RECT 87.315 123.900 87.605 125.065 ;
        RECT 87.775 123.975 90.365 125.065 ;
        RECT 90.910 124.725 91.165 124.755 ;
        RECT 90.825 124.555 91.165 124.725 ;
        RECT 90.910 124.085 91.165 124.555 ;
        RECT 91.345 124.265 91.630 125.065 ;
        RECT 91.810 124.345 92.140 124.855 ;
        RECT 86.395 123.285 87.145 123.805 ;
        RECT 87.775 123.455 88.985 123.975 ;
        RECT 89.155 123.285 90.365 123.805 ;
        RECT 83.945 123.085 84.875 123.255 ;
        RECT 83.945 123.050 84.120 123.085 ;
        RECT 83.125 122.855 83.405 123.025 ;
        RECT 83.125 122.685 83.400 122.855 ;
        RECT 83.590 122.685 84.120 123.050 ;
        RECT 84.545 122.515 84.875 122.915 ;
        RECT 85.045 122.685 85.300 123.255 ;
        RECT 85.475 122.515 87.145 123.285 ;
        RECT 87.315 122.515 87.605 123.240 ;
        RECT 87.775 122.515 90.365 123.285 ;
        RECT 90.910 123.225 91.090 124.085 ;
        RECT 91.810 123.755 92.060 124.345 ;
        RECT 92.410 124.195 92.580 124.805 ;
        RECT 92.750 124.375 93.080 125.065 ;
        RECT 93.310 124.515 93.550 124.805 ;
        RECT 93.750 124.685 94.170 125.065 ;
        RECT 94.350 124.595 94.980 124.845 ;
        RECT 95.450 124.685 95.780 125.065 ;
        RECT 94.350 124.515 94.520 124.595 ;
        RECT 95.950 124.515 96.120 124.805 ;
        RECT 96.300 124.685 96.680 125.065 ;
        RECT 96.920 124.680 97.750 124.850 ;
        RECT 93.310 124.345 94.520 124.515 ;
        RECT 91.260 123.425 92.060 123.755 ;
        RECT 90.910 122.695 91.165 123.225 ;
        RECT 91.345 122.515 91.630 122.975 ;
        RECT 91.810 122.775 92.060 123.425 ;
        RECT 92.260 124.175 92.580 124.195 ;
        RECT 92.260 124.005 94.180 124.175 ;
        RECT 92.260 123.110 92.450 124.005 ;
        RECT 94.350 123.835 94.520 124.345 ;
        RECT 94.690 124.085 95.210 124.395 ;
        RECT 92.620 123.665 94.520 123.835 ;
        RECT 92.620 123.605 92.950 123.665 ;
        RECT 93.100 123.435 93.430 123.495 ;
        RECT 92.770 123.165 93.430 123.435 ;
        RECT 92.260 122.780 92.580 123.110 ;
        RECT 92.760 122.515 93.420 122.995 ;
        RECT 93.620 122.905 93.790 123.665 ;
        RECT 94.690 123.495 94.870 123.905 ;
        RECT 93.960 123.325 94.290 123.445 ;
        RECT 95.040 123.325 95.210 124.085 ;
        RECT 93.960 123.155 95.210 123.325 ;
        RECT 95.380 124.265 96.750 124.515 ;
        RECT 95.380 123.495 95.570 124.265 ;
        RECT 96.500 124.005 96.750 124.265 ;
        RECT 95.740 123.835 95.990 123.995 ;
        RECT 96.920 123.835 97.090 124.680 ;
        RECT 97.985 124.395 98.155 124.895 ;
        RECT 98.325 124.565 98.655 125.065 ;
        RECT 97.260 124.005 97.760 124.385 ;
        RECT 97.985 124.225 98.680 124.395 ;
        RECT 95.740 123.665 97.090 123.835 ;
        RECT 96.670 123.625 97.090 123.665 ;
        RECT 95.380 123.155 95.800 123.495 ;
        RECT 96.090 123.165 96.500 123.495 ;
        RECT 93.620 122.735 94.470 122.905 ;
        RECT 95.030 122.515 95.350 122.975 ;
        RECT 95.550 122.725 95.800 123.155 ;
        RECT 96.090 122.515 96.500 122.955 ;
        RECT 96.670 122.895 96.840 123.625 ;
        RECT 97.010 123.075 97.360 123.445 ;
        RECT 97.540 123.135 97.760 124.005 ;
        RECT 97.930 123.435 98.340 124.055 ;
        RECT 98.510 123.255 98.680 124.225 ;
        RECT 97.985 123.065 98.680 123.255 ;
        RECT 96.670 122.695 97.685 122.895 ;
        RECT 97.985 122.735 98.155 123.065 ;
        RECT 98.325 122.515 98.655 122.895 ;
        RECT 98.870 122.775 99.095 124.895 ;
        RECT 99.265 124.565 99.595 125.065 ;
        RECT 99.765 124.395 99.935 124.895 ;
        RECT 99.270 124.225 99.935 124.395 ;
        RECT 100.570 124.385 100.825 124.755 ;
        RECT 99.270 123.235 99.500 124.225 ;
        RECT 100.485 124.215 100.825 124.385 ;
        RECT 101.005 124.265 101.290 125.065 ;
        RECT 101.470 124.345 101.800 124.855 ;
        RECT 100.570 124.085 100.825 124.215 ;
        RECT 99.670 123.405 100.020 124.055 ;
        RECT 99.270 123.065 99.935 123.235 ;
        RECT 99.265 122.515 99.595 122.895 ;
        RECT 99.765 122.775 99.935 123.065 ;
        RECT 100.570 123.225 100.750 124.085 ;
        RECT 101.470 123.755 101.720 124.345 ;
        RECT 102.070 124.195 102.240 124.805 ;
        RECT 102.410 124.375 102.740 125.065 ;
        RECT 102.970 124.515 103.210 124.805 ;
        RECT 103.410 124.685 103.830 125.065 ;
        RECT 104.010 124.595 104.640 124.845 ;
        RECT 105.110 124.685 105.440 125.065 ;
        RECT 104.010 124.515 104.180 124.595 ;
        RECT 105.610 124.515 105.780 124.805 ;
        RECT 105.960 124.685 106.340 125.065 ;
        RECT 106.580 124.680 107.410 124.850 ;
        RECT 102.970 124.345 104.180 124.515 ;
        RECT 100.920 123.425 101.720 123.755 ;
        RECT 100.570 122.695 100.825 123.225 ;
        RECT 101.005 122.515 101.290 122.975 ;
        RECT 101.470 122.775 101.720 123.425 ;
        RECT 101.920 124.175 102.240 124.195 ;
        RECT 101.920 124.005 103.840 124.175 ;
        RECT 101.920 123.110 102.110 124.005 ;
        RECT 104.010 123.835 104.180 124.345 ;
        RECT 104.350 124.085 104.870 124.395 ;
        RECT 102.280 123.665 104.180 123.835 ;
        RECT 102.280 123.605 102.610 123.665 ;
        RECT 102.760 123.435 103.090 123.495 ;
        RECT 102.430 123.165 103.090 123.435 ;
        RECT 101.920 122.780 102.240 123.110 ;
        RECT 102.420 122.515 103.080 122.995 ;
        RECT 103.280 122.905 103.450 123.665 ;
        RECT 104.350 123.495 104.530 123.905 ;
        RECT 103.620 123.325 103.950 123.445 ;
        RECT 104.700 123.325 104.870 124.085 ;
        RECT 103.620 123.155 104.870 123.325 ;
        RECT 105.040 124.265 106.410 124.515 ;
        RECT 105.040 123.495 105.230 124.265 ;
        RECT 106.160 124.005 106.410 124.265 ;
        RECT 105.400 123.835 105.650 123.995 ;
        RECT 106.580 123.835 106.750 124.680 ;
        RECT 107.645 124.395 107.815 124.895 ;
        RECT 107.985 124.565 108.315 125.065 ;
        RECT 106.920 124.005 107.420 124.385 ;
        RECT 107.645 124.225 108.340 124.395 ;
        RECT 105.400 123.665 106.750 123.835 ;
        RECT 106.330 123.625 106.750 123.665 ;
        RECT 105.040 123.155 105.460 123.495 ;
        RECT 105.750 123.165 106.160 123.495 ;
        RECT 103.280 122.735 104.130 122.905 ;
        RECT 104.690 122.515 105.010 122.975 ;
        RECT 105.210 122.725 105.460 123.155 ;
        RECT 105.750 122.515 106.160 122.955 ;
        RECT 106.330 122.895 106.500 123.625 ;
        RECT 106.670 123.075 107.020 123.445 ;
        RECT 107.200 123.135 107.420 124.005 ;
        RECT 107.590 123.435 108.000 124.055 ;
        RECT 108.170 123.255 108.340 124.225 ;
        RECT 107.645 123.065 108.340 123.255 ;
        RECT 106.330 122.695 107.345 122.895 ;
        RECT 107.645 122.735 107.815 123.065 ;
        RECT 107.985 122.515 108.315 122.895 ;
        RECT 108.530 122.775 108.755 124.895 ;
        RECT 108.925 124.565 109.255 125.065 ;
        RECT 109.425 124.395 109.595 124.895 ;
        RECT 108.930 124.225 109.595 124.395 ;
        RECT 108.930 123.235 109.160 124.225 ;
        RECT 109.330 123.405 109.680 124.055 ;
        RECT 110.315 123.975 111.985 125.065 ;
        RECT 112.155 123.975 113.365 125.065 ;
        RECT 110.315 123.455 111.065 123.975 ;
        RECT 111.235 123.285 111.985 123.805 ;
        RECT 112.155 123.435 112.675 123.975 ;
        RECT 108.930 123.065 109.595 123.235 ;
        RECT 108.925 122.515 109.255 122.895 ;
        RECT 109.425 122.775 109.595 123.065 ;
        RECT 110.315 122.515 111.985 123.285 ;
        RECT 112.845 123.265 113.365 123.805 ;
        RECT 112.155 122.515 113.365 123.265 ;
        RECT 15.010 122.345 113.450 122.515 ;
        RECT 15.095 121.595 16.305 122.345 ;
        RECT 17.485 121.795 17.655 122.175 ;
        RECT 17.835 121.965 18.165 122.345 ;
        RECT 17.485 121.625 18.150 121.795 ;
        RECT 18.345 121.670 18.605 122.175 ;
        RECT 15.095 121.055 15.615 121.595 ;
        RECT 15.785 120.885 16.305 121.425 ;
        RECT 17.415 121.075 17.745 121.445 ;
        RECT 17.980 121.370 18.150 121.625 ;
        RECT 17.980 121.040 18.265 121.370 ;
        RECT 17.980 120.895 18.150 121.040 ;
        RECT 15.095 119.795 16.305 120.885 ;
        RECT 17.485 120.725 18.150 120.895 ;
        RECT 18.435 120.870 18.605 121.670 ;
        RECT 17.485 119.965 17.655 120.725 ;
        RECT 17.835 119.795 18.165 120.555 ;
        RECT 18.335 119.965 18.605 120.870 ;
        RECT 18.780 121.605 19.035 122.175 ;
        RECT 19.205 121.945 19.535 122.345 ;
        RECT 19.960 121.810 20.490 122.175 ;
        RECT 19.960 121.775 20.135 121.810 ;
        RECT 19.205 121.605 20.135 121.775 ;
        RECT 20.680 121.665 20.955 122.175 ;
        RECT 18.780 120.935 18.950 121.605 ;
        RECT 19.205 121.435 19.375 121.605 ;
        RECT 19.120 121.105 19.375 121.435 ;
        RECT 19.600 121.105 19.795 121.435 ;
        RECT 18.780 119.965 19.115 120.935 ;
        RECT 19.285 119.795 19.455 120.935 ;
        RECT 19.625 120.135 19.795 121.105 ;
        RECT 19.965 120.475 20.135 121.605 ;
        RECT 20.305 120.815 20.475 121.615 ;
        RECT 20.675 121.495 20.955 121.665 ;
        RECT 20.680 121.015 20.955 121.495 ;
        RECT 21.125 120.815 21.315 122.175 ;
        RECT 21.495 121.810 22.005 122.345 ;
        RECT 22.225 121.535 22.470 122.140 ;
        RECT 22.915 121.620 23.205 122.345 ;
        RECT 21.515 121.365 22.745 121.535 ;
        RECT 23.415 121.525 23.645 122.345 ;
        RECT 23.815 121.545 24.145 122.175 ;
        RECT 20.305 120.645 21.315 120.815 ;
        RECT 21.485 120.800 22.235 120.990 ;
        RECT 19.965 120.305 21.090 120.475 ;
        RECT 21.485 120.135 21.655 120.800 ;
        RECT 22.405 120.555 22.745 121.365 ;
        RECT 23.395 121.105 23.725 121.355 ;
        RECT 19.625 119.965 21.655 120.135 ;
        RECT 21.825 119.795 21.995 120.555 ;
        RECT 22.230 120.145 22.745 120.555 ;
        RECT 22.915 119.795 23.205 120.960 ;
        RECT 23.895 120.945 24.145 121.545 ;
        RECT 24.315 121.525 24.525 122.345 ;
        RECT 25.765 121.795 25.935 122.175 ;
        RECT 26.115 121.965 26.445 122.345 ;
        RECT 25.765 121.625 26.430 121.795 ;
        RECT 26.625 121.670 26.885 122.175 ;
        RECT 27.430 122.005 27.685 122.165 ;
        RECT 27.345 121.835 27.685 122.005 ;
        RECT 27.865 121.885 28.150 122.345 ;
        RECT 25.695 121.075 26.025 121.445 ;
        RECT 26.260 121.370 26.430 121.625 ;
        RECT 23.415 119.795 23.645 120.935 ;
        RECT 23.815 119.965 24.145 120.945 ;
        RECT 26.260 121.040 26.545 121.370 ;
        RECT 24.315 119.795 24.525 120.935 ;
        RECT 26.260 120.895 26.430 121.040 ;
        RECT 25.765 120.725 26.430 120.895 ;
        RECT 26.715 120.870 26.885 121.670 ;
        RECT 25.765 119.965 25.935 120.725 ;
        RECT 26.115 119.795 26.445 120.555 ;
        RECT 26.615 119.965 26.885 120.870 ;
        RECT 27.430 121.635 27.685 121.835 ;
        RECT 27.430 120.775 27.610 121.635 ;
        RECT 28.330 121.435 28.580 122.085 ;
        RECT 27.780 121.105 28.580 121.435 ;
        RECT 27.430 120.105 27.685 120.775 ;
        RECT 27.865 119.795 28.150 120.595 ;
        RECT 28.330 120.515 28.580 121.105 ;
        RECT 28.780 121.750 29.100 122.080 ;
        RECT 29.280 121.865 29.940 122.345 ;
        RECT 30.140 121.955 30.990 122.125 ;
        RECT 28.780 120.855 28.970 121.750 ;
        RECT 29.290 121.425 29.950 121.695 ;
        RECT 29.620 121.365 29.950 121.425 ;
        RECT 29.140 121.195 29.470 121.255 ;
        RECT 30.140 121.195 30.310 121.955 ;
        RECT 31.550 121.885 31.870 122.345 ;
        RECT 32.070 121.705 32.320 122.135 ;
        RECT 32.610 121.905 33.020 122.345 ;
        RECT 33.190 121.965 34.205 122.165 ;
        RECT 30.480 121.535 31.730 121.705 ;
        RECT 30.480 121.415 30.810 121.535 ;
        RECT 29.140 121.025 31.040 121.195 ;
        RECT 28.780 120.685 30.700 120.855 ;
        RECT 28.780 120.665 29.100 120.685 ;
        RECT 28.330 120.005 28.660 120.515 ;
        RECT 28.930 120.055 29.100 120.665 ;
        RECT 30.870 120.515 31.040 121.025 ;
        RECT 31.210 120.955 31.390 121.365 ;
        RECT 31.560 120.775 31.730 121.535 ;
        RECT 29.270 119.795 29.600 120.485 ;
        RECT 29.830 120.345 31.040 120.515 ;
        RECT 31.210 120.465 31.730 120.775 ;
        RECT 31.900 121.365 32.320 121.705 ;
        RECT 32.610 121.365 33.020 121.695 ;
        RECT 31.900 120.595 32.090 121.365 ;
        RECT 33.190 121.235 33.360 121.965 ;
        RECT 34.505 121.795 34.675 122.125 ;
        RECT 34.845 121.965 35.175 122.345 ;
        RECT 33.530 121.415 33.880 121.785 ;
        RECT 33.190 121.195 33.610 121.235 ;
        RECT 32.260 121.025 33.610 121.195 ;
        RECT 32.260 120.865 32.510 121.025 ;
        RECT 33.020 120.595 33.270 120.855 ;
        RECT 31.900 120.345 33.270 120.595 ;
        RECT 29.830 120.055 30.070 120.345 ;
        RECT 30.870 120.265 31.040 120.345 ;
        RECT 30.270 119.795 30.690 120.175 ;
        RECT 30.870 120.015 31.500 120.265 ;
        RECT 31.970 119.795 32.300 120.175 ;
        RECT 32.470 120.055 32.640 120.345 ;
        RECT 33.440 120.180 33.610 121.025 ;
        RECT 34.060 120.855 34.280 121.725 ;
        RECT 34.505 121.605 35.200 121.795 ;
        RECT 33.780 120.475 34.280 120.855 ;
        RECT 34.450 120.805 34.860 121.425 ;
        RECT 35.030 120.635 35.200 121.605 ;
        RECT 34.505 120.465 35.200 120.635 ;
        RECT 32.820 119.795 33.200 120.175 ;
        RECT 33.440 120.010 34.270 120.180 ;
        RECT 34.505 119.965 34.675 120.465 ;
        RECT 34.845 119.795 35.175 120.295 ;
        RECT 35.390 119.965 35.615 122.085 ;
        RECT 35.785 121.965 36.115 122.345 ;
        RECT 36.285 121.795 36.455 122.085 ;
        RECT 35.790 121.625 36.455 121.795 ;
        RECT 35.790 120.635 36.020 121.625 ;
        RECT 36.715 121.595 37.925 122.345 ;
        RECT 38.470 122.005 38.725 122.165 ;
        RECT 38.385 121.835 38.725 122.005 ;
        RECT 38.905 121.885 39.190 122.345 ;
        RECT 36.190 120.805 36.540 121.455 ;
        RECT 36.715 120.885 37.235 121.425 ;
        RECT 37.405 121.055 37.925 121.595 ;
        RECT 38.470 121.635 38.725 121.835 ;
        RECT 35.790 120.465 36.455 120.635 ;
        RECT 35.785 119.795 36.115 120.295 ;
        RECT 36.285 119.965 36.455 120.465 ;
        RECT 36.715 119.795 37.925 120.885 ;
        RECT 38.470 120.775 38.650 121.635 ;
        RECT 39.370 121.435 39.620 122.085 ;
        RECT 38.820 121.105 39.620 121.435 ;
        RECT 38.470 120.105 38.725 120.775 ;
        RECT 38.905 119.795 39.190 120.595 ;
        RECT 39.370 120.515 39.620 121.105 ;
        RECT 39.820 121.750 40.140 122.080 ;
        RECT 40.320 121.865 40.980 122.345 ;
        RECT 41.180 121.955 42.030 122.125 ;
        RECT 39.820 120.855 40.010 121.750 ;
        RECT 40.330 121.425 40.990 121.695 ;
        RECT 40.660 121.365 40.990 121.425 ;
        RECT 40.180 121.195 40.510 121.255 ;
        RECT 41.180 121.195 41.350 121.955 ;
        RECT 42.590 121.885 42.910 122.345 ;
        RECT 43.110 121.705 43.360 122.135 ;
        RECT 43.650 121.905 44.060 122.345 ;
        RECT 44.230 121.965 45.245 122.165 ;
        RECT 41.520 121.535 42.770 121.705 ;
        RECT 41.520 121.415 41.850 121.535 ;
        RECT 40.180 121.025 42.080 121.195 ;
        RECT 39.820 120.685 41.740 120.855 ;
        RECT 39.820 120.665 40.140 120.685 ;
        RECT 39.370 120.005 39.700 120.515 ;
        RECT 39.970 120.055 40.140 120.665 ;
        RECT 41.910 120.515 42.080 121.025 ;
        RECT 42.250 120.955 42.430 121.365 ;
        RECT 42.600 120.775 42.770 121.535 ;
        RECT 40.310 119.795 40.640 120.485 ;
        RECT 40.870 120.345 42.080 120.515 ;
        RECT 42.250 120.465 42.770 120.775 ;
        RECT 42.940 121.365 43.360 121.705 ;
        RECT 43.650 121.365 44.060 121.695 ;
        RECT 42.940 120.595 43.130 121.365 ;
        RECT 44.230 121.235 44.400 121.965 ;
        RECT 45.545 121.795 45.715 122.125 ;
        RECT 45.885 121.965 46.215 122.345 ;
        RECT 44.570 121.415 44.920 121.785 ;
        RECT 44.230 121.195 44.650 121.235 ;
        RECT 43.300 121.025 44.650 121.195 ;
        RECT 43.300 120.865 43.550 121.025 ;
        RECT 44.060 120.595 44.310 120.855 ;
        RECT 42.940 120.345 44.310 120.595 ;
        RECT 40.870 120.055 41.110 120.345 ;
        RECT 41.910 120.265 42.080 120.345 ;
        RECT 41.310 119.795 41.730 120.175 ;
        RECT 41.910 120.015 42.540 120.265 ;
        RECT 43.010 119.795 43.340 120.175 ;
        RECT 43.510 120.055 43.680 120.345 ;
        RECT 44.480 120.180 44.650 121.025 ;
        RECT 45.100 120.855 45.320 121.725 ;
        RECT 45.545 121.605 46.240 121.795 ;
        RECT 44.820 120.475 45.320 120.855 ;
        RECT 45.490 120.805 45.900 121.425 ;
        RECT 46.070 120.635 46.240 121.605 ;
        RECT 45.545 120.465 46.240 120.635 ;
        RECT 43.860 119.795 44.240 120.175 ;
        RECT 44.480 120.010 45.310 120.180 ;
        RECT 45.545 119.965 45.715 120.465 ;
        RECT 45.885 119.795 46.215 120.295 ;
        RECT 46.430 119.965 46.655 122.085 ;
        RECT 46.825 121.965 47.155 122.345 ;
        RECT 47.325 121.795 47.495 122.085 ;
        RECT 46.830 121.625 47.495 121.795 ;
        RECT 46.830 120.635 47.060 121.625 ;
        RECT 48.675 121.620 48.965 122.345 ;
        RECT 49.195 121.525 49.405 122.345 ;
        RECT 49.575 121.545 49.905 122.175 ;
        RECT 47.230 120.805 47.580 121.455 ;
        RECT 46.830 120.465 47.495 120.635 ;
        RECT 46.825 119.795 47.155 120.295 ;
        RECT 47.325 119.965 47.495 120.465 ;
        RECT 48.675 119.795 48.965 120.960 ;
        RECT 49.575 120.945 49.825 121.545 ;
        RECT 50.075 121.525 50.305 122.345 ;
        RECT 50.605 121.795 50.775 122.175 ;
        RECT 50.955 121.965 51.285 122.345 ;
        RECT 50.605 121.625 51.270 121.795 ;
        RECT 51.465 121.670 51.725 122.175 ;
        RECT 49.995 121.105 50.325 121.355 ;
        RECT 50.535 121.075 50.865 121.445 ;
        RECT 51.100 121.370 51.270 121.625 ;
        RECT 51.100 121.040 51.385 121.370 ;
        RECT 49.195 119.795 49.405 120.935 ;
        RECT 49.575 119.965 49.905 120.945 ;
        RECT 50.075 119.795 50.305 120.935 ;
        RECT 51.100 120.895 51.270 121.040 ;
        RECT 50.605 120.725 51.270 120.895 ;
        RECT 51.555 120.870 51.725 121.670 ;
        RECT 52.045 121.545 52.375 122.345 ;
        RECT 52.545 121.695 52.715 122.175 ;
        RECT 52.885 121.865 53.215 122.345 ;
        RECT 53.385 121.695 53.555 122.175 ;
        RECT 53.805 121.865 54.045 122.345 ;
        RECT 54.225 121.695 54.395 122.175 ;
        RECT 52.545 121.525 53.555 121.695 ;
        RECT 53.760 121.525 54.395 121.695 ;
        RECT 54.655 121.595 55.865 122.345 ;
        RECT 52.545 120.985 53.040 121.525 ;
        RECT 53.760 121.355 53.930 121.525 ;
        RECT 53.430 121.185 53.930 121.355 ;
        RECT 50.605 119.965 50.775 120.725 ;
        RECT 50.955 119.795 51.285 120.555 ;
        RECT 51.455 119.965 51.725 120.870 ;
        RECT 52.045 119.795 52.375 120.945 ;
        RECT 52.545 120.815 53.555 120.985 ;
        RECT 52.545 119.965 52.715 120.815 ;
        RECT 52.885 119.795 53.215 120.595 ;
        RECT 53.385 119.965 53.555 120.815 ;
        RECT 53.760 120.945 53.930 121.185 ;
        RECT 54.100 121.115 54.480 121.355 ;
        RECT 53.760 120.775 54.475 120.945 ;
        RECT 53.735 119.795 53.975 120.595 ;
        RECT 54.145 119.965 54.475 120.775 ;
        RECT 54.655 120.885 55.175 121.425 ;
        RECT 55.345 121.055 55.865 121.595 ;
        RECT 56.095 121.525 56.305 122.345 ;
        RECT 56.475 121.545 56.805 122.175 ;
        RECT 56.475 120.945 56.725 121.545 ;
        RECT 56.975 121.525 57.205 122.345 ;
        RECT 57.415 121.575 59.085 122.345 ;
        RECT 59.260 121.800 64.605 122.345 ;
        RECT 56.895 121.105 57.225 121.355 ;
        RECT 54.655 119.795 55.865 120.885 ;
        RECT 56.095 119.795 56.305 120.935 ;
        RECT 56.475 119.965 56.805 120.945 ;
        RECT 56.975 119.795 57.205 120.935 ;
        RECT 57.415 120.885 58.165 121.405 ;
        RECT 58.335 121.055 59.085 121.575 ;
        RECT 57.415 119.795 59.085 120.885 ;
        RECT 60.850 120.230 61.200 121.480 ;
        RECT 62.680 120.970 63.020 121.800 ;
        RECT 64.865 121.795 65.035 122.085 ;
        RECT 65.205 121.965 65.535 122.345 ;
        RECT 64.865 121.625 65.530 121.795 ;
        RECT 64.780 120.805 65.130 121.455 ;
        RECT 65.300 120.635 65.530 121.625 ;
        RECT 64.865 120.465 65.530 120.635 ;
        RECT 59.260 119.795 64.605 120.230 ;
        RECT 64.865 119.965 65.035 120.465 ;
        RECT 65.205 119.795 65.535 120.295 ;
        RECT 65.705 119.965 65.930 122.085 ;
        RECT 66.145 121.965 66.475 122.345 ;
        RECT 66.645 121.795 66.815 122.125 ;
        RECT 67.115 121.965 68.130 122.165 ;
        RECT 66.120 121.605 66.815 121.795 ;
        RECT 66.120 120.635 66.290 121.605 ;
        RECT 66.460 120.805 66.870 121.425 ;
        RECT 67.040 120.855 67.260 121.725 ;
        RECT 67.440 121.415 67.790 121.785 ;
        RECT 67.960 121.235 68.130 121.965 ;
        RECT 68.300 121.905 68.710 122.345 ;
        RECT 69.000 121.705 69.250 122.135 ;
        RECT 69.450 121.885 69.770 122.345 ;
        RECT 70.330 121.955 71.180 122.125 ;
        RECT 68.300 121.365 68.710 121.695 ;
        RECT 69.000 121.365 69.420 121.705 ;
        RECT 67.710 121.195 68.130 121.235 ;
        RECT 67.710 121.025 69.060 121.195 ;
        RECT 66.120 120.465 66.815 120.635 ;
        RECT 67.040 120.475 67.540 120.855 ;
        RECT 66.145 119.795 66.475 120.295 ;
        RECT 66.645 119.965 66.815 120.465 ;
        RECT 67.710 120.180 67.880 121.025 ;
        RECT 68.810 120.865 69.060 121.025 ;
        RECT 68.050 120.595 68.300 120.855 ;
        RECT 69.230 120.595 69.420 121.365 ;
        RECT 68.050 120.345 69.420 120.595 ;
        RECT 69.590 121.535 70.840 121.705 ;
        RECT 69.590 120.775 69.760 121.535 ;
        RECT 70.510 121.415 70.840 121.535 ;
        RECT 69.930 120.955 70.110 121.365 ;
        RECT 71.010 121.195 71.180 121.955 ;
        RECT 71.380 121.865 72.040 122.345 ;
        RECT 72.220 121.750 72.540 122.080 ;
        RECT 71.370 121.425 72.030 121.695 ;
        RECT 71.370 121.365 71.700 121.425 ;
        RECT 71.850 121.195 72.180 121.255 ;
        RECT 70.280 121.025 72.180 121.195 ;
        RECT 69.590 120.465 70.110 120.775 ;
        RECT 70.280 120.515 70.450 121.025 ;
        RECT 72.350 120.855 72.540 121.750 ;
        RECT 70.620 120.685 72.540 120.855 ;
        RECT 72.220 120.665 72.540 120.685 ;
        RECT 72.740 121.435 72.990 122.085 ;
        RECT 73.170 121.885 73.455 122.345 ;
        RECT 73.635 122.005 73.890 122.165 ;
        RECT 73.635 121.835 73.975 122.005 ;
        RECT 73.635 121.635 73.890 121.835 ;
        RECT 72.740 121.105 73.540 121.435 ;
        RECT 70.280 120.345 71.490 120.515 ;
        RECT 67.050 120.010 67.880 120.180 ;
        RECT 68.120 119.795 68.500 120.175 ;
        RECT 68.680 120.055 68.850 120.345 ;
        RECT 70.280 120.265 70.450 120.345 ;
        RECT 69.020 119.795 69.350 120.175 ;
        RECT 69.820 120.015 70.450 120.265 ;
        RECT 70.630 119.795 71.050 120.175 ;
        RECT 71.250 120.055 71.490 120.345 ;
        RECT 71.720 119.795 72.050 120.485 ;
        RECT 72.220 120.055 72.390 120.665 ;
        RECT 72.740 120.515 72.990 121.105 ;
        RECT 73.710 120.775 73.890 121.635 ;
        RECT 74.435 121.620 74.725 122.345 ;
        RECT 74.985 121.795 75.155 122.175 ;
        RECT 75.335 121.965 75.665 122.345 ;
        RECT 74.985 121.625 75.650 121.795 ;
        RECT 75.845 121.670 76.105 122.175 ;
        RECT 74.915 121.075 75.245 121.445 ;
        RECT 75.480 121.370 75.650 121.625 ;
        RECT 75.480 121.040 75.765 121.370 ;
        RECT 72.660 120.005 72.990 120.515 ;
        RECT 73.170 119.795 73.455 120.595 ;
        RECT 73.635 120.105 73.890 120.775 ;
        RECT 74.435 119.795 74.725 120.960 ;
        RECT 75.480 120.895 75.650 121.040 ;
        RECT 74.985 120.725 75.650 120.895 ;
        RECT 75.935 120.870 76.105 121.670 ;
        RECT 76.275 121.595 77.485 122.345 ;
        RECT 74.985 119.965 75.155 120.725 ;
        RECT 75.335 119.795 75.665 120.555 ;
        RECT 75.835 119.965 76.105 120.870 ;
        RECT 76.275 120.885 76.795 121.425 ;
        RECT 76.965 121.055 77.485 121.595 ;
        RECT 78.030 121.635 78.285 122.165 ;
        RECT 78.465 121.885 78.750 122.345 ;
        RECT 76.275 119.795 77.485 120.885 ;
        RECT 78.030 120.775 78.210 121.635 ;
        RECT 78.930 121.435 79.180 122.085 ;
        RECT 78.380 121.105 79.180 121.435 ;
        RECT 78.030 120.305 78.285 120.775 ;
        RECT 77.945 120.135 78.285 120.305 ;
        RECT 78.030 120.105 78.285 120.135 ;
        RECT 78.465 119.795 78.750 120.595 ;
        RECT 78.930 120.515 79.180 121.105 ;
        RECT 79.380 121.750 79.700 122.080 ;
        RECT 79.880 121.865 80.540 122.345 ;
        RECT 80.740 121.955 81.590 122.125 ;
        RECT 79.380 120.855 79.570 121.750 ;
        RECT 79.890 121.425 80.550 121.695 ;
        RECT 80.220 121.365 80.550 121.425 ;
        RECT 79.740 121.195 80.070 121.255 ;
        RECT 80.740 121.195 80.910 121.955 ;
        RECT 82.150 121.885 82.470 122.345 ;
        RECT 82.670 121.705 82.920 122.135 ;
        RECT 83.210 121.905 83.620 122.345 ;
        RECT 83.790 121.965 84.805 122.165 ;
        RECT 81.080 121.535 82.330 121.705 ;
        RECT 81.080 121.415 81.410 121.535 ;
        RECT 79.740 121.025 81.640 121.195 ;
        RECT 79.380 120.685 81.300 120.855 ;
        RECT 79.380 120.665 79.700 120.685 ;
        RECT 78.930 120.005 79.260 120.515 ;
        RECT 79.530 120.055 79.700 120.665 ;
        RECT 81.470 120.515 81.640 121.025 ;
        RECT 81.810 120.955 81.990 121.365 ;
        RECT 82.160 120.775 82.330 121.535 ;
        RECT 79.870 119.795 80.200 120.485 ;
        RECT 80.430 120.345 81.640 120.515 ;
        RECT 81.810 120.465 82.330 120.775 ;
        RECT 82.500 121.365 82.920 121.705 ;
        RECT 83.210 121.365 83.620 121.695 ;
        RECT 82.500 120.595 82.690 121.365 ;
        RECT 83.790 121.235 83.960 121.965 ;
        RECT 85.105 121.795 85.275 122.125 ;
        RECT 85.445 121.965 85.775 122.345 ;
        RECT 84.130 121.415 84.480 121.785 ;
        RECT 83.790 121.195 84.210 121.235 ;
        RECT 82.860 121.025 84.210 121.195 ;
        RECT 82.860 120.865 83.110 121.025 ;
        RECT 83.620 120.595 83.870 120.855 ;
        RECT 82.500 120.345 83.870 120.595 ;
        RECT 80.430 120.055 80.670 120.345 ;
        RECT 81.470 120.265 81.640 120.345 ;
        RECT 80.870 119.795 81.290 120.175 ;
        RECT 81.470 120.015 82.100 120.265 ;
        RECT 82.570 119.795 82.900 120.175 ;
        RECT 83.070 120.055 83.240 120.345 ;
        RECT 84.040 120.180 84.210 121.025 ;
        RECT 84.660 120.855 84.880 121.725 ;
        RECT 85.105 121.605 85.800 121.795 ;
        RECT 84.380 120.475 84.880 120.855 ;
        RECT 85.050 120.805 85.460 121.425 ;
        RECT 85.630 120.635 85.800 121.605 ;
        RECT 85.105 120.465 85.800 120.635 ;
        RECT 83.420 119.795 83.800 120.175 ;
        RECT 84.040 120.010 84.870 120.180 ;
        RECT 85.105 119.965 85.275 120.465 ;
        RECT 85.445 119.795 85.775 120.295 ;
        RECT 85.990 119.965 86.215 122.085 ;
        RECT 86.385 121.965 86.715 122.345 ;
        RECT 86.885 121.795 87.055 122.085 ;
        RECT 87.690 122.005 87.945 122.165 ;
        RECT 87.605 121.835 87.945 122.005 ;
        RECT 88.125 121.885 88.410 122.345 ;
        RECT 86.390 121.625 87.055 121.795 ;
        RECT 87.690 121.635 87.945 121.835 ;
        RECT 86.390 120.635 86.620 121.625 ;
        RECT 86.790 120.805 87.140 121.455 ;
        RECT 87.690 120.775 87.870 121.635 ;
        RECT 88.590 121.435 88.840 122.085 ;
        RECT 88.040 121.105 88.840 121.435 ;
        RECT 86.390 120.465 87.055 120.635 ;
        RECT 86.385 119.795 86.715 120.295 ;
        RECT 86.885 119.965 87.055 120.465 ;
        RECT 87.690 120.105 87.945 120.775 ;
        RECT 88.125 119.795 88.410 120.595 ;
        RECT 88.590 120.515 88.840 121.105 ;
        RECT 89.040 121.750 89.360 122.080 ;
        RECT 89.540 121.865 90.200 122.345 ;
        RECT 90.400 121.955 91.250 122.125 ;
        RECT 89.040 120.855 89.230 121.750 ;
        RECT 89.550 121.425 90.210 121.695 ;
        RECT 89.880 121.365 90.210 121.425 ;
        RECT 89.400 121.195 89.730 121.255 ;
        RECT 90.400 121.195 90.570 121.955 ;
        RECT 91.810 121.885 92.130 122.345 ;
        RECT 92.330 121.705 92.580 122.135 ;
        RECT 92.870 121.905 93.280 122.345 ;
        RECT 93.450 121.965 94.465 122.165 ;
        RECT 90.740 121.535 91.990 121.705 ;
        RECT 90.740 121.415 91.070 121.535 ;
        RECT 89.400 121.025 91.300 121.195 ;
        RECT 89.040 120.685 90.960 120.855 ;
        RECT 89.040 120.665 89.360 120.685 ;
        RECT 88.590 120.005 88.920 120.515 ;
        RECT 89.190 120.055 89.360 120.665 ;
        RECT 91.130 120.515 91.300 121.025 ;
        RECT 91.470 120.955 91.650 121.365 ;
        RECT 91.820 120.775 91.990 121.535 ;
        RECT 89.530 119.795 89.860 120.485 ;
        RECT 90.090 120.345 91.300 120.515 ;
        RECT 91.470 120.465 91.990 120.775 ;
        RECT 92.160 121.365 92.580 121.705 ;
        RECT 92.870 121.365 93.280 121.695 ;
        RECT 92.160 120.595 92.350 121.365 ;
        RECT 93.450 121.235 93.620 121.965 ;
        RECT 94.765 121.795 94.935 122.125 ;
        RECT 95.105 121.965 95.435 122.345 ;
        RECT 93.790 121.415 94.140 121.785 ;
        RECT 93.450 121.195 93.870 121.235 ;
        RECT 92.520 121.025 93.870 121.195 ;
        RECT 92.520 120.865 92.770 121.025 ;
        RECT 93.280 120.595 93.530 120.855 ;
        RECT 92.160 120.345 93.530 120.595 ;
        RECT 90.090 120.055 90.330 120.345 ;
        RECT 91.130 120.265 91.300 120.345 ;
        RECT 90.530 119.795 90.950 120.175 ;
        RECT 91.130 120.015 91.760 120.265 ;
        RECT 92.230 119.795 92.560 120.175 ;
        RECT 92.730 120.055 92.900 120.345 ;
        RECT 93.700 120.180 93.870 121.025 ;
        RECT 94.320 120.855 94.540 121.725 ;
        RECT 94.765 121.605 95.460 121.795 ;
        RECT 94.040 120.475 94.540 120.855 ;
        RECT 94.710 120.805 95.120 121.425 ;
        RECT 95.290 120.635 95.460 121.605 ;
        RECT 94.765 120.465 95.460 120.635 ;
        RECT 93.080 119.795 93.460 120.175 ;
        RECT 93.700 120.010 94.530 120.180 ;
        RECT 94.765 119.965 94.935 120.465 ;
        RECT 95.105 119.795 95.435 120.295 ;
        RECT 95.650 119.965 95.875 122.085 ;
        RECT 96.045 121.965 96.375 122.345 ;
        RECT 96.545 121.795 96.715 122.085 ;
        RECT 96.050 121.625 96.715 121.795 ;
        RECT 97.435 121.670 97.695 122.175 ;
        RECT 97.875 121.965 98.205 122.345 ;
        RECT 98.385 121.795 98.555 122.175 ;
        RECT 96.050 120.635 96.280 121.625 ;
        RECT 96.450 120.805 96.800 121.455 ;
        RECT 97.435 120.870 97.605 121.670 ;
        RECT 97.890 121.625 98.555 121.795 ;
        RECT 97.890 121.370 98.060 121.625 ;
        RECT 98.815 121.595 100.025 122.345 ;
        RECT 100.195 121.620 100.485 122.345 ;
        RECT 97.775 121.040 98.060 121.370 ;
        RECT 98.295 121.075 98.625 121.445 ;
        RECT 97.890 120.895 98.060 121.040 ;
        RECT 96.050 120.465 96.715 120.635 ;
        RECT 96.045 119.795 96.375 120.295 ;
        RECT 96.545 119.965 96.715 120.465 ;
        RECT 97.435 119.965 97.705 120.870 ;
        RECT 97.890 120.725 98.555 120.895 ;
        RECT 97.875 119.795 98.205 120.555 ;
        RECT 98.385 119.965 98.555 120.725 ;
        RECT 98.815 120.885 99.335 121.425 ;
        RECT 99.505 121.055 100.025 121.595 ;
        RECT 100.930 121.535 101.175 122.140 ;
        RECT 101.395 121.810 101.905 122.345 ;
        RECT 100.655 121.365 101.885 121.535 ;
        RECT 98.815 119.795 100.025 120.885 ;
        RECT 100.195 119.795 100.485 120.960 ;
        RECT 100.655 120.555 100.995 121.365 ;
        RECT 101.165 120.800 101.915 120.990 ;
        RECT 100.655 120.145 101.170 120.555 ;
        RECT 101.405 119.795 101.575 120.555 ;
        RECT 101.745 120.135 101.915 120.800 ;
        RECT 102.085 120.815 102.275 122.175 ;
        RECT 102.445 122.005 102.720 122.175 ;
        RECT 102.445 121.835 102.725 122.005 ;
        RECT 102.445 121.015 102.720 121.835 ;
        RECT 102.910 121.810 103.440 122.175 ;
        RECT 103.865 121.945 104.195 122.345 ;
        RECT 103.265 121.775 103.440 121.810 ;
        RECT 102.925 120.815 103.095 121.615 ;
        RECT 102.085 120.645 103.095 120.815 ;
        RECT 103.265 121.605 104.195 121.775 ;
        RECT 104.365 121.605 104.620 122.175 ;
        RECT 104.885 121.795 105.055 122.175 ;
        RECT 105.235 121.965 105.565 122.345 ;
        RECT 104.885 121.625 105.550 121.795 ;
        RECT 105.745 121.670 106.005 122.175 ;
        RECT 103.265 120.475 103.435 121.605 ;
        RECT 104.025 121.435 104.195 121.605 ;
        RECT 102.310 120.305 103.435 120.475 ;
        RECT 103.605 121.105 103.800 121.435 ;
        RECT 104.025 121.105 104.280 121.435 ;
        RECT 103.605 120.135 103.775 121.105 ;
        RECT 104.450 120.935 104.620 121.605 ;
        RECT 104.815 121.075 105.145 121.445 ;
        RECT 105.380 121.370 105.550 121.625 ;
        RECT 101.745 119.965 103.775 120.135 ;
        RECT 103.945 119.795 104.115 120.935 ;
        RECT 104.285 119.965 104.620 120.935 ;
        RECT 105.380 121.040 105.665 121.370 ;
        RECT 105.380 120.895 105.550 121.040 ;
        RECT 104.885 120.725 105.550 120.895 ;
        RECT 105.835 120.870 106.005 121.670 ;
        RECT 106.725 121.795 106.895 122.175 ;
        RECT 107.075 121.965 107.405 122.345 ;
        RECT 106.725 121.625 107.390 121.795 ;
        RECT 107.585 121.670 107.845 122.175 ;
        RECT 106.655 121.075 106.985 121.445 ;
        RECT 107.220 121.370 107.390 121.625 ;
        RECT 107.220 121.040 107.505 121.370 ;
        RECT 107.220 120.895 107.390 121.040 ;
        RECT 104.885 119.965 105.055 120.725 ;
        RECT 105.235 119.795 105.565 120.555 ;
        RECT 105.735 119.965 106.005 120.870 ;
        RECT 106.725 120.725 107.390 120.895 ;
        RECT 107.675 120.870 107.845 121.670 ;
        RECT 108.475 121.575 111.985 122.345 ;
        RECT 112.155 121.595 113.365 122.345 ;
        RECT 106.725 119.965 106.895 120.725 ;
        RECT 107.075 119.795 107.405 120.555 ;
        RECT 107.575 119.965 107.845 120.870 ;
        RECT 108.475 120.885 110.165 121.405 ;
        RECT 110.335 121.055 111.985 121.575 ;
        RECT 112.155 120.885 112.675 121.425 ;
        RECT 112.845 121.055 113.365 121.595 ;
        RECT 108.475 119.795 111.985 120.885 ;
        RECT 112.155 119.795 113.365 120.885 ;
        RECT 15.010 119.625 113.450 119.795 ;
        RECT 15.095 118.535 16.305 119.625 ;
        RECT 15.095 117.825 15.615 118.365 ;
        RECT 15.785 117.995 16.305 118.535 ;
        RECT 16.475 118.535 19.065 119.625 ;
        RECT 19.545 118.785 19.715 119.625 ;
        RECT 19.925 118.615 20.175 119.455 ;
        RECT 20.385 118.785 20.555 119.625 ;
        RECT 20.725 118.615 21.015 119.455 ;
        RECT 16.475 118.015 17.685 118.535 ;
        RECT 19.290 118.445 21.015 118.615 ;
        RECT 21.225 118.565 21.395 119.625 ;
        RECT 21.690 119.245 22.020 119.625 ;
        RECT 22.200 119.075 22.370 119.365 ;
        RECT 22.540 119.165 22.790 119.625 ;
        RECT 21.570 118.905 22.370 119.075 ;
        RECT 22.960 119.115 23.830 119.455 ;
        RECT 17.855 117.845 19.065 118.365 ;
        RECT 15.095 117.075 16.305 117.825 ;
        RECT 16.475 117.075 19.065 117.845 ;
        RECT 19.290 117.895 19.700 118.445 ;
        RECT 21.570 118.285 21.740 118.905 ;
        RECT 22.960 118.735 23.130 119.115 ;
        RECT 24.065 118.995 24.235 119.455 ;
        RECT 24.405 119.165 24.775 119.625 ;
        RECT 25.070 119.025 25.240 119.365 ;
        RECT 25.410 119.195 25.740 119.625 ;
        RECT 25.975 119.025 26.145 119.365 ;
        RECT 21.910 118.565 23.130 118.735 ;
        RECT 23.300 118.655 23.760 118.945 ;
        RECT 24.065 118.825 24.625 118.995 ;
        RECT 25.070 118.855 26.145 119.025 ;
        RECT 26.315 119.125 26.995 119.455 ;
        RECT 27.210 119.125 27.460 119.455 ;
        RECT 27.630 119.165 27.880 119.625 ;
        RECT 24.455 118.685 24.625 118.825 ;
        RECT 23.300 118.645 24.265 118.655 ;
        RECT 22.960 118.475 23.130 118.565 ;
        RECT 23.590 118.485 24.265 118.645 ;
        RECT 21.570 118.275 21.915 118.285 ;
        RECT 19.885 118.065 21.915 118.275 ;
        RECT 19.290 117.725 21.055 117.895 ;
        RECT 19.545 117.075 19.715 117.545 ;
        RECT 19.885 117.245 20.215 117.725 ;
        RECT 20.385 117.075 20.555 117.545 ;
        RECT 20.725 117.245 21.055 117.725 ;
        RECT 21.225 117.075 21.395 117.885 ;
        RECT 21.590 117.810 21.915 118.065 ;
        RECT 21.595 117.455 21.915 117.810 ;
        RECT 22.085 118.025 22.625 118.395 ;
        RECT 22.960 118.305 23.365 118.475 ;
        RECT 22.085 117.625 22.325 118.025 ;
        RECT 22.805 117.855 23.025 118.135 ;
        RECT 22.495 117.685 23.025 117.855 ;
        RECT 22.495 117.455 22.665 117.685 ;
        RECT 23.195 117.525 23.365 118.305 ;
        RECT 23.535 117.695 23.885 118.315 ;
        RECT 24.055 117.695 24.265 118.485 ;
        RECT 24.455 118.515 25.955 118.685 ;
        RECT 24.455 117.825 24.625 118.515 ;
        RECT 26.315 118.345 26.485 119.125 ;
        RECT 27.290 118.995 27.460 119.125 ;
        RECT 24.795 118.175 26.485 118.345 ;
        RECT 26.655 118.565 27.120 118.955 ;
        RECT 27.290 118.825 27.685 118.995 ;
        RECT 24.795 117.995 24.965 118.175 ;
        RECT 21.595 117.285 22.665 117.455 ;
        RECT 22.835 117.075 23.025 117.515 ;
        RECT 23.195 117.245 24.145 117.525 ;
        RECT 24.455 117.435 24.715 117.825 ;
        RECT 25.135 117.755 25.925 118.005 ;
        RECT 24.365 117.265 24.715 117.435 ;
        RECT 24.925 117.075 25.255 117.535 ;
        RECT 26.130 117.465 26.300 118.175 ;
        RECT 26.655 117.975 26.825 118.565 ;
        RECT 26.470 117.755 26.825 117.975 ;
        RECT 26.995 117.755 27.345 118.375 ;
        RECT 27.515 117.465 27.685 118.825 ;
        RECT 28.050 118.655 28.375 119.440 ;
        RECT 27.855 117.605 28.315 118.655 ;
        RECT 26.130 117.295 26.985 117.465 ;
        RECT 27.190 117.295 27.685 117.465 ;
        RECT 27.855 117.075 28.185 117.435 ;
        RECT 28.545 117.335 28.715 119.455 ;
        RECT 28.885 119.125 29.215 119.625 ;
        RECT 29.385 118.955 29.640 119.455 ;
        RECT 28.890 118.785 29.640 118.955 ;
        RECT 28.890 117.795 29.120 118.785 ;
        RECT 29.290 117.965 29.640 118.615 ;
        RECT 30.315 118.485 30.545 119.625 ;
        RECT 30.715 118.475 31.045 119.455 ;
        RECT 31.215 118.485 31.425 119.625 ;
        RECT 31.655 118.535 33.325 119.625 ;
        RECT 33.585 118.695 33.755 119.455 ;
        RECT 33.935 118.865 34.265 119.625 ;
        RECT 30.295 118.065 30.625 118.315 ;
        RECT 28.890 117.625 29.640 117.795 ;
        RECT 28.885 117.075 29.215 117.455 ;
        RECT 29.385 117.335 29.640 117.625 ;
        RECT 30.315 117.075 30.545 117.895 ;
        RECT 30.795 117.875 31.045 118.475 ;
        RECT 31.655 118.015 32.405 118.535 ;
        RECT 33.585 118.525 34.250 118.695 ;
        RECT 34.435 118.550 34.705 119.455 ;
        RECT 34.080 118.380 34.250 118.525 ;
        RECT 30.715 117.245 31.045 117.875 ;
        RECT 31.215 117.075 31.425 117.895 ;
        RECT 32.575 117.845 33.325 118.365 ;
        RECT 33.515 117.975 33.845 118.345 ;
        RECT 34.080 118.050 34.365 118.380 ;
        RECT 31.655 117.075 33.325 117.845 ;
        RECT 34.080 117.795 34.250 118.050 ;
        RECT 33.585 117.625 34.250 117.795 ;
        RECT 34.535 117.750 34.705 118.550 ;
        RECT 35.795 118.460 36.085 119.625 ;
        RECT 36.255 118.535 37.465 119.625 ;
        RECT 37.635 118.535 41.145 119.625 ;
        RECT 36.255 117.995 36.775 118.535 ;
        RECT 36.945 117.825 37.465 118.365 ;
        RECT 37.635 118.015 39.325 118.535 ;
        RECT 41.355 118.485 41.585 119.625 ;
        RECT 41.755 118.475 42.085 119.455 ;
        RECT 42.255 118.485 42.465 119.625 ;
        RECT 43.245 118.695 43.415 119.455 ;
        RECT 43.595 118.865 43.925 119.625 ;
        RECT 43.245 118.525 43.910 118.695 ;
        RECT 44.095 118.550 44.365 119.455 ;
        RECT 44.910 119.285 45.165 119.315 ;
        RECT 44.825 119.115 45.165 119.285 ;
        RECT 39.495 117.845 41.145 118.365 ;
        RECT 41.335 118.065 41.665 118.315 ;
        RECT 33.585 117.245 33.755 117.625 ;
        RECT 33.935 117.075 34.265 117.455 ;
        RECT 34.445 117.245 34.705 117.750 ;
        RECT 35.795 117.075 36.085 117.800 ;
        RECT 36.255 117.075 37.465 117.825 ;
        RECT 37.635 117.075 41.145 117.845 ;
        RECT 41.355 117.075 41.585 117.895 ;
        RECT 41.835 117.875 42.085 118.475 ;
        RECT 43.740 118.380 43.910 118.525 ;
        RECT 43.175 117.975 43.505 118.345 ;
        RECT 43.740 118.050 44.025 118.380 ;
        RECT 41.755 117.245 42.085 117.875 ;
        RECT 42.255 117.075 42.465 117.895 ;
        RECT 43.740 117.795 43.910 118.050 ;
        RECT 43.245 117.625 43.910 117.795 ;
        RECT 44.195 117.750 44.365 118.550 ;
        RECT 43.245 117.245 43.415 117.625 ;
        RECT 43.595 117.075 43.925 117.455 ;
        RECT 44.105 117.245 44.365 117.750 ;
        RECT 44.910 118.645 45.165 119.115 ;
        RECT 45.345 118.825 45.630 119.625 ;
        RECT 45.810 118.905 46.140 119.415 ;
        RECT 44.910 117.785 45.090 118.645 ;
        RECT 45.810 118.315 46.060 118.905 ;
        RECT 46.410 118.755 46.580 119.365 ;
        RECT 46.750 118.935 47.080 119.625 ;
        RECT 47.310 119.075 47.550 119.365 ;
        RECT 47.750 119.245 48.170 119.625 ;
        RECT 48.350 119.155 48.980 119.405 ;
        RECT 49.450 119.245 49.780 119.625 ;
        RECT 48.350 119.075 48.520 119.155 ;
        RECT 49.950 119.075 50.120 119.365 ;
        RECT 50.300 119.245 50.680 119.625 ;
        RECT 50.920 119.240 51.750 119.410 ;
        RECT 47.310 118.905 48.520 119.075 ;
        RECT 45.260 117.985 46.060 118.315 ;
        RECT 44.910 117.255 45.165 117.785 ;
        RECT 45.345 117.075 45.630 117.535 ;
        RECT 45.810 117.335 46.060 117.985 ;
        RECT 46.260 118.735 46.580 118.755 ;
        RECT 46.260 118.565 48.180 118.735 ;
        RECT 46.260 117.670 46.450 118.565 ;
        RECT 48.350 118.395 48.520 118.905 ;
        RECT 48.690 118.645 49.210 118.955 ;
        RECT 46.620 118.225 48.520 118.395 ;
        RECT 46.620 118.165 46.950 118.225 ;
        RECT 47.100 117.995 47.430 118.055 ;
        RECT 46.770 117.725 47.430 117.995 ;
        RECT 46.260 117.340 46.580 117.670 ;
        RECT 46.760 117.075 47.420 117.555 ;
        RECT 47.620 117.465 47.790 118.225 ;
        RECT 48.690 118.055 48.870 118.465 ;
        RECT 47.960 117.885 48.290 118.005 ;
        RECT 49.040 117.885 49.210 118.645 ;
        RECT 47.960 117.715 49.210 117.885 ;
        RECT 49.380 118.825 50.750 119.075 ;
        RECT 49.380 118.055 49.570 118.825 ;
        RECT 50.500 118.565 50.750 118.825 ;
        RECT 49.740 118.395 49.990 118.555 ;
        RECT 50.920 118.395 51.090 119.240 ;
        RECT 51.985 118.955 52.155 119.455 ;
        RECT 52.325 119.125 52.655 119.625 ;
        RECT 51.260 118.565 51.760 118.945 ;
        RECT 51.985 118.785 52.680 118.955 ;
        RECT 49.740 118.225 51.090 118.395 ;
        RECT 50.670 118.185 51.090 118.225 ;
        RECT 49.380 117.715 49.800 118.055 ;
        RECT 50.090 117.725 50.500 118.055 ;
        RECT 47.620 117.295 48.470 117.465 ;
        RECT 49.030 117.075 49.350 117.535 ;
        RECT 49.550 117.285 49.800 117.715 ;
        RECT 50.090 117.075 50.500 117.515 ;
        RECT 50.670 117.455 50.840 118.185 ;
        RECT 51.010 117.635 51.360 118.005 ;
        RECT 51.540 117.695 51.760 118.565 ;
        RECT 51.930 117.995 52.340 118.615 ;
        RECT 52.510 117.815 52.680 118.785 ;
        RECT 51.985 117.625 52.680 117.815 ;
        RECT 50.670 117.255 51.685 117.455 ;
        RECT 51.985 117.295 52.155 117.625 ;
        RECT 52.325 117.075 52.655 117.455 ;
        RECT 52.870 117.335 53.095 119.455 ;
        RECT 53.265 119.125 53.595 119.625 ;
        RECT 53.765 118.955 53.935 119.455 ;
        RECT 53.270 118.785 53.935 118.955 ;
        RECT 53.270 117.795 53.500 118.785 ;
        RECT 53.670 117.965 54.020 118.615 ;
        RECT 54.195 118.535 55.865 119.625 ;
        RECT 56.040 119.190 61.385 119.625 ;
        RECT 54.195 118.015 54.945 118.535 ;
        RECT 55.115 117.845 55.865 118.365 ;
        RECT 57.630 117.940 57.980 119.190 ;
        RECT 61.555 118.460 61.845 119.625 ;
        RECT 62.015 118.535 64.605 119.625 ;
        RECT 64.780 119.190 70.125 119.625 ;
        RECT 53.270 117.625 53.935 117.795 ;
        RECT 53.265 117.075 53.595 117.455 ;
        RECT 53.765 117.335 53.935 117.625 ;
        RECT 54.195 117.075 55.865 117.845 ;
        RECT 59.460 117.620 59.800 118.450 ;
        RECT 62.015 118.015 63.225 118.535 ;
        RECT 63.395 117.845 64.605 118.365 ;
        RECT 66.370 117.940 66.720 119.190 ;
        RECT 70.335 118.485 70.565 119.625 ;
        RECT 70.735 118.475 71.065 119.455 ;
        RECT 71.235 118.485 71.445 119.625 ;
        RECT 71.675 118.865 72.190 119.275 ;
        RECT 72.425 118.865 72.595 119.625 ;
        RECT 72.765 119.285 74.795 119.455 ;
        RECT 56.040 117.075 61.385 117.620 ;
        RECT 61.555 117.075 61.845 117.800 ;
        RECT 62.015 117.075 64.605 117.845 ;
        RECT 68.200 117.620 68.540 118.450 ;
        RECT 70.315 118.065 70.645 118.315 ;
        RECT 64.780 117.075 70.125 117.620 ;
        RECT 70.335 117.075 70.565 117.895 ;
        RECT 70.815 117.875 71.065 118.475 ;
        RECT 71.675 118.055 72.015 118.865 ;
        RECT 72.765 118.620 72.935 119.285 ;
        RECT 73.330 118.945 74.455 119.115 ;
        RECT 72.185 118.430 72.935 118.620 ;
        RECT 73.105 118.605 74.115 118.775 ;
        RECT 70.735 117.245 71.065 117.875 ;
        RECT 71.235 117.075 71.445 117.895 ;
        RECT 71.675 117.885 72.905 118.055 ;
        RECT 71.950 117.280 72.195 117.885 ;
        RECT 72.415 117.075 72.925 117.610 ;
        RECT 73.105 117.245 73.295 118.605 ;
        RECT 73.465 117.585 73.740 118.405 ;
        RECT 73.945 117.805 74.115 118.605 ;
        RECT 74.285 117.815 74.455 118.945 ;
        RECT 74.625 118.315 74.795 119.285 ;
        RECT 74.965 118.485 75.135 119.625 ;
        RECT 75.305 118.485 75.640 119.455 ;
        RECT 75.820 119.190 81.165 119.625 ;
        RECT 74.625 117.985 74.820 118.315 ;
        RECT 75.045 117.985 75.300 118.315 ;
        RECT 75.045 117.815 75.215 117.985 ;
        RECT 75.470 117.815 75.640 118.485 ;
        RECT 77.410 117.940 77.760 119.190 ;
        RECT 81.395 118.485 81.605 119.625 ;
        RECT 81.775 118.475 82.105 119.455 ;
        RECT 82.275 118.485 82.505 119.625 ;
        RECT 83.215 118.485 83.445 119.625 ;
        RECT 83.615 118.475 83.945 119.455 ;
        RECT 84.115 118.485 84.325 119.625 ;
        RECT 84.645 118.695 84.815 119.455 ;
        RECT 84.995 118.865 85.325 119.625 ;
        RECT 84.645 118.525 85.310 118.695 ;
        RECT 85.495 118.550 85.765 119.455 ;
        RECT 74.285 117.645 75.215 117.815 ;
        RECT 74.285 117.610 74.460 117.645 ;
        RECT 73.465 117.415 73.745 117.585 ;
        RECT 73.465 117.245 73.740 117.415 ;
        RECT 73.930 117.245 74.460 117.610 ;
        RECT 74.885 117.075 75.215 117.475 ;
        RECT 75.385 117.245 75.640 117.815 ;
        RECT 79.240 117.620 79.580 118.450 ;
        RECT 75.820 117.075 81.165 117.620 ;
        RECT 81.395 117.075 81.605 117.895 ;
        RECT 81.775 117.875 82.025 118.475 ;
        RECT 82.195 118.065 82.525 118.315 ;
        RECT 83.195 118.065 83.525 118.315 ;
        RECT 81.775 117.245 82.105 117.875 ;
        RECT 82.275 117.075 82.505 117.895 ;
        RECT 83.215 117.075 83.445 117.895 ;
        RECT 83.695 117.875 83.945 118.475 ;
        RECT 85.140 118.380 85.310 118.525 ;
        RECT 84.575 117.975 84.905 118.345 ;
        RECT 85.140 118.050 85.425 118.380 ;
        RECT 83.615 117.245 83.945 117.875 ;
        RECT 84.115 117.075 84.325 117.895 ;
        RECT 85.140 117.795 85.310 118.050 ;
        RECT 84.645 117.625 85.310 117.795 ;
        RECT 85.595 117.750 85.765 118.550 ;
        RECT 85.935 118.535 87.145 119.625 ;
        RECT 85.935 117.995 86.455 118.535 ;
        RECT 87.315 118.460 87.605 119.625 ;
        RECT 88.235 118.535 90.825 119.625 ;
        RECT 91.085 118.695 91.255 119.455 ;
        RECT 91.435 118.865 91.765 119.625 ;
        RECT 86.625 117.825 87.145 118.365 ;
        RECT 88.235 118.015 89.445 118.535 ;
        RECT 91.085 118.525 91.750 118.695 ;
        RECT 91.935 118.550 92.205 119.455 ;
        RECT 91.580 118.380 91.750 118.525 ;
        RECT 89.615 117.845 90.825 118.365 ;
        RECT 91.015 117.975 91.345 118.345 ;
        RECT 91.580 118.050 91.865 118.380 ;
        RECT 84.645 117.245 84.815 117.625 ;
        RECT 84.995 117.075 85.325 117.455 ;
        RECT 85.505 117.245 85.765 117.750 ;
        RECT 85.935 117.075 87.145 117.825 ;
        RECT 87.315 117.075 87.605 117.800 ;
        RECT 88.235 117.075 90.825 117.845 ;
        RECT 91.580 117.795 91.750 118.050 ;
        RECT 91.085 117.625 91.750 117.795 ;
        RECT 92.035 117.750 92.205 118.550 ;
        RECT 92.835 118.535 94.505 119.625 ;
        RECT 94.680 119.190 100.025 119.625 ;
        RECT 100.200 119.190 105.545 119.625 ;
        RECT 92.835 118.015 93.585 118.535 ;
        RECT 93.755 117.845 94.505 118.365 ;
        RECT 96.270 117.940 96.620 119.190 ;
        RECT 91.085 117.245 91.255 117.625 ;
        RECT 91.435 117.075 91.765 117.455 ;
        RECT 91.945 117.245 92.205 117.750 ;
        RECT 92.835 117.075 94.505 117.845 ;
        RECT 98.100 117.620 98.440 118.450 ;
        RECT 101.790 117.940 102.140 119.190 ;
        RECT 105.755 118.485 105.985 119.625 ;
        RECT 106.155 118.475 106.485 119.455 ;
        RECT 106.655 118.485 106.865 119.625 ;
        RECT 107.185 118.695 107.355 119.455 ;
        RECT 107.535 118.865 107.865 119.625 ;
        RECT 107.185 118.525 107.850 118.695 ;
        RECT 108.035 118.550 108.305 119.455 ;
        RECT 103.620 117.620 103.960 118.450 ;
        RECT 105.735 118.065 106.065 118.315 ;
        RECT 94.680 117.075 100.025 117.620 ;
        RECT 100.200 117.075 105.545 117.620 ;
        RECT 105.755 117.075 105.985 117.895 ;
        RECT 106.235 117.875 106.485 118.475 ;
        RECT 107.680 118.380 107.850 118.525 ;
        RECT 107.115 117.975 107.445 118.345 ;
        RECT 107.680 118.050 107.965 118.380 ;
        RECT 106.155 117.245 106.485 117.875 ;
        RECT 106.655 117.075 106.865 117.895 ;
        RECT 107.680 117.795 107.850 118.050 ;
        RECT 107.185 117.625 107.850 117.795 ;
        RECT 108.135 117.750 108.305 118.550 ;
        RECT 107.185 117.245 107.355 117.625 ;
        RECT 107.535 117.075 107.865 117.455 ;
        RECT 108.045 117.245 108.305 117.750 ;
        RECT 108.475 118.550 108.745 119.455 ;
        RECT 108.915 118.865 109.245 119.625 ;
        RECT 109.425 118.695 109.595 119.455 ;
        RECT 108.475 117.750 108.645 118.550 ;
        RECT 108.930 118.525 109.595 118.695 ;
        RECT 110.315 118.535 111.985 119.625 ;
        RECT 112.155 118.535 113.365 119.625 ;
        RECT 108.930 118.380 109.100 118.525 ;
        RECT 108.815 118.050 109.100 118.380 ;
        RECT 108.930 117.795 109.100 118.050 ;
        RECT 109.335 117.975 109.665 118.345 ;
        RECT 110.315 118.015 111.065 118.535 ;
        RECT 111.235 117.845 111.985 118.365 ;
        RECT 112.155 117.995 112.675 118.535 ;
        RECT 108.475 117.245 108.735 117.750 ;
        RECT 108.930 117.625 109.595 117.795 ;
        RECT 108.915 117.075 109.245 117.455 ;
        RECT 109.425 117.245 109.595 117.625 ;
        RECT 110.315 117.075 111.985 117.845 ;
        RECT 112.845 117.825 113.365 118.365 ;
        RECT 112.155 117.075 113.365 117.825 ;
        RECT 15.010 116.905 113.450 117.075 ;
        RECT 15.095 116.155 16.305 116.905 ;
        RECT 17.400 116.360 22.745 116.905 ;
        RECT 15.095 115.615 15.615 116.155 ;
        RECT 15.785 115.445 16.305 115.985 ;
        RECT 15.095 114.355 16.305 115.445 ;
        RECT 18.990 114.790 19.340 116.040 ;
        RECT 20.820 115.530 21.160 116.360 ;
        RECT 22.915 116.180 23.205 116.905 ;
        RECT 23.685 116.435 23.855 116.905 ;
        RECT 24.025 116.255 24.355 116.735 ;
        RECT 24.525 116.435 24.695 116.905 ;
        RECT 24.865 116.255 25.195 116.735 ;
        RECT 23.430 116.085 25.195 116.255 ;
        RECT 25.365 116.095 25.535 116.905 ;
        RECT 25.735 116.525 26.805 116.695 ;
        RECT 25.735 116.170 26.055 116.525 ;
        RECT 23.430 115.535 23.840 116.085 ;
        RECT 25.730 115.915 26.055 116.170 ;
        RECT 24.025 115.705 26.055 115.915 ;
        RECT 25.710 115.695 26.055 115.705 ;
        RECT 26.225 115.955 26.465 116.355 ;
        RECT 26.635 116.295 26.805 116.525 ;
        RECT 26.975 116.465 27.165 116.905 ;
        RECT 27.335 116.455 28.285 116.735 ;
        RECT 28.505 116.545 28.855 116.715 ;
        RECT 26.635 116.125 27.165 116.295 ;
        RECT 17.400 114.355 22.745 114.790 ;
        RECT 22.915 114.355 23.205 115.520 ;
        RECT 23.430 115.365 25.155 115.535 ;
        RECT 23.685 114.355 23.855 115.195 ;
        RECT 24.065 114.525 24.315 115.365 ;
        RECT 24.525 114.355 24.695 115.195 ;
        RECT 24.865 114.525 25.155 115.365 ;
        RECT 25.365 114.355 25.535 115.415 ;
        RECT 25.710 115.075 25.880 115.695 ;
        RECT 26.225 115.585 26.765 115.955 ;
        RECT 26.945 115.845 27.165 116.125 ;
        RECT 27.335 115.675 27.505 116.455 ;
        RECT 27.100 115.505 27.505 115.675 ;
        RECT 27.675 115.665 28.025 116.285 ;
        RECT 27.100 115.415 27.270 115.505 ;
        RECT 28.195 115.495 28.405 116.285 ;
        RECT 26.050 115.245 27.270 115.415 ;
        RECT 27.730 115.335 28.405 115.495 ;
        RECT 25.710 114.905 26.510 115.075 ;
        RECT 25.830 114.355 26.160 114.735 ;
        RECT 26.340 114.615 26.510 114.905 ;
        RECT 27.100 114.865 27.270 115.245 ;
        RECT 27.440 115.325 28.405 115.335 ;
        RECT 28.595 116.155 28.855 116.545 ;
        RECT 29.065 116.445 29.395 116.905 ;
        RECT 30.270 116.515 31.125 116.685 ;
        RECT 31.330 116.515 31.825 116.685 ;
        RECT 31.995 116.545 32.325 116.905 ;
        RECT 28.595 115.465 28.765 116.155 ;
        RECT 28.935 115.805 29.105 115.985 ;
        RECT 29.275 115.975 30.065 116.225 ;
        RECT 30.270 115.805 30.440 116.515 ;
        RECT 30.610 116.005 30.965 116.225 ;
        RECT 28.935 115.635 30.625 115.805 ;
        RECT 27.440 115.035 27.900 115.325 ;
        RECT 28.595 115.295 30.095 115.465 ;
        RECT 28.595 115.155 28.765 115.295 ;
        RECT 28.205 114.985 28.765 115.155 ;
        RECT 26.680 114.355 26.930 114.815 ;
        RECT 27.100 114.525 27.970 114.865 ;
        RECT 28.205 114.525 28.375 114.985 ;
        RECT 29.210 114.955 30.285 115.125 ;
        RECT 28.545 114.355 28.915 114.815 ;
        RECT 29.210 114.615 29.380 114.955 ;
        RECT 29.550 114.355 29.880 114.785 ;
        RECT 30.115 114.615 30.285 114.955 ;
        RECT 30.455 114.855 30.625 115.635 ;
        RECT 30.795 115.415 30.965 116.005 ;
        RECT 31.135 115.605 31.485 116.225 ;
        RECT 30.795 115.025 31.260 115.415 ;
        RECT 31.655 115.155 31.825 116.515 ;
        RECT 31.995 115.325 32.455 116.375 ;
        RECT 31.430 114.985 31.825 115.155 ;
        RECT 31.430 114.855 31.600 114.985 ;
        RECT 30.455 114.525 31.135 114.855 ;
        RECT 31.350 114.525 31.600 114.855 ;
        RECT 31.770 114.355 32.020 114.815 ;
        RECT 32.190 114.540 32.515 115.325 ;
        RECT 32.685 114.525 32.855 116.645 ;
        RECT 33.025 116.525 33.355 116.905 ;
        RECT 33.525 116.355 33.780 116.645 ;
        RECT 33.030 116.185 33.780 116.355 ;
        RECT 34.415 116.230 34.675 116.735 ;
        RECT 34.855 116.525 35.185 116.905 ;
        RECT 35.365 116.355 35.535 116.735 ;
        RECT 36.260 116.360 41.605 116.905 ;
        RECT 41.780 116.360 47.125 116.905 ;
        RECT 33.030 115.195 33.260 116.185 ;
        RECT 33.430 115.365 33.780 116.015 ;
        RECT 34.415 115.430 34.585 116.230 ;
        RECT 34.870 116.185 35.535 116.355 ;
        RECT 34.870 115.930 35.040 116.185 ;
        RECT 34.755 115.600 35.040 115.930 ;
        RECT 35.275 115.635 35.605 116.005 ;
        RECT 34.870 115.455 35.040 115.600 ;
        RECT 33.030 115.025 33.780 115.195 ;
        RECT 33.025 114.355 33.355 114.855 ;
        RECT 33.525 114.525 33.780 115.025 ;
        RECT 34.415 114.525 34.685 115.430 ;
        RECT 34.870 115.285 35.535 115.455 ;
        RECT 34.855 114.355 35.185 115.115 ;
        RECT 35.365 114.525 35.535 115.285 ;
        RECT 37.850 114.790 38.200 116.040 ;
        RECT 39.680 115.530 40.020 116.360 ;
        RECT 43.370 114.790 43.720 116.040 ;
        RECT 45.200 115.530 45.540 116.360 ;
        RECT 47.385 116.355 47.555 116.735 ;
        RECT 47.735 116.525 48.065 116.905 ;
        RECT 47.385 116.185 48.050 116.355 ;
        RECT 48.245 116.230 48.505 116.735 ;
        RECT 47.315 115.635 47.645 116.005 ;
        RECT 47.880 115.930 48.050 116.185 ;
        RECT 47.880 115.600 48.165 115.930 ;
        RECT 47.880 115.455 48.050 115.600 ;
        RECT 47.385 115.285 48.050 115.455 ;
        RECT 48.335 115.430 48.505 116.230 ;
        RECT 48.675 116.180 48.965 116.905 ;
        RECT 49.135 116.155 50.345 116.905 ;
        RECT 50.520 116.360 55.865 116.905 ;
        RECT 36.260 114.355 41.605 114.790 ;
        RECT 41.780 114.355 47.125 114.790 ;
        RECT 47.385 114.525 47.555 115.285 ;
        RECT 47.735 114.355 48.065 115.115 ;
        RECT 48.235 114.525 48.505 115.430 ;
        RECT 48.675 114.355 48.965 115.520 ;
        RECT 49.135 115.445 49.655 115.985 ;
        RECT 49.825 115.615 50.345 116.155 ;
        RECT 49.135 114.355 50.345 115.445 ;
        RECT 52.110 114.790 52.460 116.040 ;
        RECT 53.940 115.530 54.280 116.360 ;
        RECT 56.125 116.255 56.295 116.735 ;
        RECT 56.475 116.425 56.715 116.905 ;
        RECT 56.965 116.255 57.135 116.735 ;
        RECT 57.305 116.425 57.635 116.905 ;
        RECT 57.805 116.255 57.975 116.735 ;
        RECT 56.125 116.085 56.760 116.255 ;
        RECT 56.965 116.085 57.975 116.255 ;
        RECT 58.145 116.105 58.475 116.905 ;
        RECT 58.800 116.360 64.145 116.905 ;
        RECT 64.320 116.360 69.665 116.905 ;
        RECT 56.590 115.915 56.760 116.085 ;
        RECT 56.040 115.675 56.420 115.915 ;
        RECT 56.590 115.745 57.090 115.915 ;
        RECT 56.590 115.505 56.760 115.745 ;
        RECT 57.480 115.545 57.975 116.085 ;
        RECT 56.045 115.335 56.760 115.505 ;
        RECT 56.965 115.375 57.975 115.545 ;
        RECT 50.520 114.355 55.865 114.790 ;
        RECT 56.045 114.525 56.375 115.335 ;
        RECT 56.545 114.355 56.785 115.155 ;
        RECT 56.965 114.525 57.135 115.375 ;
        RECT 57.305 114.355 57.635 115.155 ;
        RECT 57.805 114.525 57.975 115.375 ;
        RECT 58.145 114.355 58.475 115.505 ;
        RECT 60.390 114.790 60.740 116.040 ;
        RECT 62.220 115.530 62.560 116.360 ;
        RECT 65.910 114.790 66.260 116.040 ;
        RECT 67.740 115.530 68.080 116.360 ;
        RECT 69.895 116.085 70.105 116.905 ;
        RECT 70.275 116.105 70.605 116.735 ;
        RECT 70.275 115.505 70.525 116.105 ;
        RECT 70.775 116.085 71.005 116.905 ;
        RECT 71.765 116.255 71.935 116.735 ;
        RECT 72.115 116.425 72.355 116.905 ;
        RECT 72.605 116.255 72.775 116.735 ;
        RECT 72.945 116.425 73.275 116.905 ;
        RECT 73.445 116.255 73.615 116.735 ;
        RECT 71.765 116.085 72.400 116.255 ;
        RECT 72.605 116.085 73.615 116.255 ;
        RECT 73.785 116.105 74.115 116.905 ;
        RECT 74.435 116.180 74.725 116.905 ;
        RECT 74.895 116.135 77.485 116.905 ;
        RECT 77.745 116.355 77.915 116.735 ;
        RECT 78.095 116.525 78.425 116.905 ;
        RECT 77.745 116.185 78.410 116.355 ;
        RECT 78.605 116.230 78.865 116.735 ;
        RECT 72.230 115.915 72.400 116.085 ;
        RECT 73.115 116.055 73.615 116.085 ;
        RECT 70.695 115.665 71.025 115.915 ;
        RECT 71.680 115.675 72.060 115.915 ;
        RECT 72.230 115.745 72.730 115.915 ;
        RECT 72.230 115.505 72.400 115.745 ;
        RECT 73.120 115.545 73.615 116.055 ;
        RECT 58.800 114.355 64.145 114.790 ;
        RECT 64.320 114.355 69.665 114.790 ;
        RECT 69.895 114.355 70.105 115.495 ;
        RECT 70.275 114.525 70.605 115.505 ;
        RECT 70.775 114.355 71.005 115.495 ;
        RECT 71.685 115.335 72.400 115.505 ;
        RECT 72.605 115.375 73.615 115.545 ;
        RECT 71.685 114.525 72.015 115.335 ;
        RECT 72.185 114.355 72.425 115.155 ;
        RECT 72.605 114.525 72.775 115.375 ;
        RECT 72.945 114.355 73.275 115.155 ;
        RECT 73.445 114.525 73.615 115.375 ;
        RECT 73.785 114.355 74.115 115.505 ;
        RECT 74.435 114.355 74.725 115.520 ;
        RECT 74.895 115.445 76.105 115.965 ;
        RECT 76.275 115.615 77.485 116.135 ;
        RECT 77.675 115.635 78.005 116.005 ;
        RECT 78.240 115.930 78.410 116.185 ;
        RECT 78.240 115.600 78.525 115.930 ;
        RECT 78.240 115.455 78.410 115.600 ;
        RECT 74.895 114.355 77.485 115.445 ;
        RECT 77.745 115.285 78.410 115.455 ;
        RECT 78.695 115.430 78.865 116.230 ;
        RECT 79.495 116.135 83.005 116.905 ;
        RECT 77.745 114.525 77.915 115.285 ;
        RECT 78.095 114.355 78.425 115.115 ;
        RECT 78.595 114.525 78.865 115.430 ;
        RECT 79.495 115.445 81.185 115.965 ;
        RECT 81.355 115.615 83.005 116.135 ;
        RECT 83.235 116.085 83.445 116.905 ;
        RECT 83.615 116.105 83.945 116.735 ;
        RECT 83.615 115.505 83.865 116.105 ;
        RECT 84.115 116.085 84.345 116.905 ;
        RECT 84.555 116.155 85.765 116.905 ;
        RECT 84.035 115.665 84.365 115.915 ;
        RECT 79.495 114.355 83.005 115.445 ;
        RECT 83.235 114.355 83.445 115.495 ;
        RECT 83.615 114.525 83.945 115.505 ;
        RECT 84.115 114.355 84.345 115.495 ;
        RECT 84.555 115.445 85.075 115.985 ;
        RECT 85.245 115.615 85.765 116.155 ;
        RECT 85.935 116.135 89.445 116.905 ;
        RECT 89.705 116.355 89.875 116.735 ;
        RECT 90.055 116.525 90.385 116.905 ;
        RECT 89.705 116.185 90.370 116.355 ;
        RECT 90.565 116.230 90.825 116.735 ;
        RECT 85.935 115.445 87.625 115.965 ;
        RECT 87.795 115.615 89.445 116.135 ;
        RECT 89.635 115.635 89.965 116.005 ;
        RECT 90.200 115.930 90.370 116.185 ;
        RECT 90.200 115.600 90.485 115.930 ;
        RECT 90.200 115.455 90.370 115.600 ;
        RECT 84.555 114.355 85.765 115.445 ;
        RECT 85.935 114.355 89.445 115.445 ;
        RECT 89.705 115.285 90.370 115.455 ;
        RECT 90.655 115.430 90.825 116.230 ;
        RECT 90.995 116.135 94.505 116.905 ;
        RECT 94.765 116.355 94.935 116.735 ;
        RECT 95.115 116.525 95.445 116.905 ;
        RECT 94.765 116.185 95.430 116.355 ;
        RECT 95.625 116.230 95.885 116.735 ;
        RECT 89.705 114.525 89.875 115.285 ;
        RECT 90.055 114.355 90.385 115.115 ;
        RECT 90.555 114.525 90.825 115.430 ;
        RECT 90.995 115.445 92.685 115.965 ;
        RECT 92.855 115.615 94.505 116.135 ;
        RECT 94.695 115.635 95.025 116.005 ;
        RECT 95.260 115.930 95.430 116.185 ;
        RECT 95.260 115.600 95.545 115.930 ;
        RECT 95.260 115.455 95.430 115.600 ;
        RECT 90.995 114.355 94.505 115.445 ;
        RECT 94.765 115.285 95.430 115.455 ;
        RECT 95.715 115.430 95.885 116.230 ;
        RECT 96.055 116.135 98.645 116.905 ;
        RECT 98.905 116.355 99.075 116.735 ;
        RECT 99.255 116.525 99.585 116.905 ;
        RECT 98.905 116.185 99.570 116.355 ;
        RECT 99.765 116.230 100.025 116.735 ;
        RECT 94.765 114.525 94.935 115.285 ;
        RECT 95.115 114.355 95.445 115.115 ;
        RECT 95.615 114.525 95.885 115.430 ;
        RECT 96.055 115.445 97.265 115.965 ;
        RECT 97.435 115.615 98.645 116.135 ;
        RECT 98.835 115.635 99.165 116.005 ;
        RECT 99.400 115.930 99.570 116.185 ;
        RECT 99.400 115.600 99.685 115.930 ;
        RECT 99.400 115.455 99.570 115.600 ;
        RECT 96.055 114.355 98.645 115.445 ;
        RECT 98.905 115.285 99.570 115.455 ;
        RECT 99.855 115.430 100.025 116.230 ;
        RECT 100.195 116.180 100.485 116.905 ;
        RECT 101.580 116.355 101.835 116.645 ;
        RECT 102.005 116.525 102.335 116.905 ;
        RECT 101.580 116.185 102.330 116.355 ;
        RECT 98.905 114.525 99.075 115.285 ;
        RECT 99.255 114.355 99.585 115.115 ;
        RECT 99.755 114.525 100.025 115.430 ;
        RECT 100.195 114.355 100.485 115.520 ;
        RECT 101.580 115.365 101.930 116.015 ;
        RECT 102.100 115.195 102.330 116.185 ;
        RECT 101.580 115.025 102.330 115.195 ;
        RECT 101.580 114.525 101.835 115.025 ;
        RECT 102.005 114.355 102.335 114.855 ;
        RECT 102.505 114.525 102.675 116.645 ;
        RECT 103.035 116.545 103.365 116.905 ;
        RECT 103.535 116.515 104.030 116.685 ;
        RECT 104.235 116.515 105.090 116.685 ;
        RECT 102.905 115.325 103.365 116.375 ;
        RECT 102.845 114.540 103.170 115.325 ;
        RECT 103.535 115.155 103.705 116.515 ;
        RECT 103.875 115.605 104.225 116.225 ;
        RECT 104.395 116.005 104.750 116.225 ;
        RECT 104.395 115.415 104.565 116.005 ;
        RECT 104.920 115.805 105.090 116.515 ;
        RECT 105.965 116.445 106.295 116.905 ;
        RECT 106.505 116.545 106.855 116.715 ;
        RECT 105.295 115.975 106.085 116.225 ;
        RECT 106.505 116.155 106.765 116.545 ;
        RECT 107.075 116.455 108.025 116.735 ;
        RECT 108.195 116.465 108.385 116.905 ;
        RECT 108.555 116.525 109.625 116.695 ;
        RECT 106.255 115.805 106.425 115.985 ;
        RECT 103.535 114.985 103.930 115.155 ;
        RECT 104.100 115.025 104.565 115.415 ;
        RECT 104.735 115.635 106.425 115.805 ;
        RECT 103.760 114.855 103.930 114.985 ;
        RECT 104.735 114.855 104.905 115.635 ;
        RECT 106.595 115.465 106.765 116.155 ;
        RECT 105.265 115.295 106.765 115.465 ;
        RECT 106.955 115.495 107.165 116.285 ;
        RECT 107.335 115.665 107.685 116.285 ;
        RECT 107.855 115.675 108.025 116.455 ;
        RECT 108.555 116.295 108.725 116.525 ;
        RECT 108.195 116.125 108.725 116.295 ;
        RECT 108.195 115.845 108.415 116.125 ;
        RECT 108.895 115.955 109.135 116.355 ;
        RECT 107.855 115.505 108.260 115.675 ;
        RECT 108.595 115.585 109.135 115.955 ;
        RECT 109.305 116.170 109.625 116.525 ;
        RECT 109.305 115.915 109.630 116.170 ;
        RECT 109.825 116.095 109.995 116.905 ;
        RECT 110.165 116.255 110.495 116.735 ;
        RECT 110.665 116.435 110.835 116.905 ;
        RECT 111.005 116.255 111.335 116.735 ;
        RECT 111.505 116.435 111.675 116.905 ;
        RECT 110.165 116.085 111.930 116.255 ;
        RECT 112.155 116.155 113.365 116.905 ;
        RECT 109.305 115.705 111.335 115.915 ;
        RECT 109.305 115.695 109.650 115.705 ;
        RECT 106.955 115.335 107.630 115.495 ;
        RECT 108.090 115.415 108.260 115.505 ;
        RECT 106.955 115.325 107.920 115.335 ;
        RECT 106.595 115.155 106.765 115.295 ;
        RECT 103.340 114.355 103.590 114.815 ;
        RECT 103.760 114.525 104.010 114.855 ;
        RECT 104.225 114.525 104.905 114.855 ;
        RECT 105.075 114.955 106.150 115.125 ;
        RECT 106.595 114.985 107.155 115.155 ;
        RECT 107.460 115.035 107.920 115.325 ;
        RECT 108.090 115.245 109.310 115.415 ;
        RECT 105.075 114.615 105.245 114.955 ;
        RECT 105.480 114.355 105.810 114.785 ;
        RECT 105.980 114.615 106.150 114.955 ;
        RECT 106.445 114.355 106.815 114.815 ;
        RECT 106.985 114.525 107.155 114.985 ;
        RECT 108.090 114.865 108.260 115.245 ;
        RECT 109.480 115.075 109.650 115.695 ;
        RECT 111.520 115.535 111.930 116.085 ;
        RECT 107.390 114.525 108.260 114.865 ;
        RECT 108.850 114.905 109.650 115.075 ;
        RECT 108.430 114.355 108.680 114.815 ;
        RECT 108.850 114.615 109.020 114.905 ;
        RECT 109.200 114.355 109.530 114.735 ;
        RECT 109.825 114.355 109.995 115.415 ;
        RECT 110.205 115.365 111.930 115.535 ;
        RECT 112.155 115.445 112.675 115.985 ;
        RECT 112.845 115.615 113.365 116.155 ;
        RECT 110.205 114.525 110.495 115.365 ;
        RECT 110.665 114.355 110.835 115.195 ;
        RECT 111.045 114.525 111.295 115.365 ;
        RECT 111.505 114.355 111.675 115.195 ;
        RECT 112.155 114.355 113.365 115.445 ;
        RECT 15.010 114.185 113.450 114.355 ;
        RECT 15.095 113.095 16.305 114.185 ;
        RECT 16.940 113.750 22.285 114.185 ;
        RECT 15.095 112.385 15.615 112.925 ;
        RECT 15.785 112.555 16.305 113.095 ;
        RECT 18.530 112.500 18.880 113.750 ;
        RECT 22.545 113.255 22.715 114.015 ;
        RECT 22.895 113.425 23.225 114.185 ;
        RECT 22.545 113.085 23.210 113.255 ;
        RECT 23.395 113.110 23.665 114.015 ;
        RECT 15.095 111.635 16.305 112.385 ;
        RECT 20.360 112.180 20.700 113.010 ;
        RECT 23.040 112.940 23.210 113.085 ;
        RECT 22.475 112.535 22.805 112.905 ;
        RECT 23.040 112.610 23.325 112.940 ;
        RECT 23.040 112.355 23.210 112.610 ;
        RECT 22.545 112.185 23.210 112.355 ;
        RECT 23.495 112.310 23.665 113.110 ;
        RECT 23.925 113.255 24.095 114.015 ;
        RECT 24.275 113.425 24.605 114.185 ;
        RECT 23.925 113.085 24.590 113.255 ;
        RECT 24.775 113.110 25.045 114.015 ;
        RECT 25.525 113.345 25.695 114.185 ;
        RECT 25.905 113.175 26.155 114.015 ;
        RECT 26.365 113.345 26.535 114.185 ;
        RECT 26.705 113.175 26.995 114.015 ;
        RECT 24.420 112.940 24.590 113.085 ;
        RECT 23.855 112.535 24.185 112.905 ;
        RECT 24.420 112.610 24.705 112.940 ;
        RECT 24.420 112.355 24.590 112.610 ;
        RECT 16.940 111.635 22.285 112.180 ;
        RECT 22.545 111.805 22.715 112.185 ;
        RECT 22.895 111.635 23.225 112.015 ;
        RECT 23.405 111.805 23.665 112.310 ;
        RECT 23.925 112.185 24.590 112.355 ;
        RECT 24.875 112.310 25.045 113.110 ;
        RECT 23.925 111.805 24.095 112.185 ;
        RECT 24.275 111.635 24.605 112.015 ;
        RECT 24.785 111.805 25.045 112.310 ;
        RECT 25.270 113.005 26.995 113.175 ;
        RECT 27.205 113.125 27.375 114.185 ;
        RECT 27.670 113.805 28.000 114.185 ;
        RECT 28.180 113.635 28.350 113.925 ;
        RECT 28.520 113.725 28.770 114.185 ;
        RECT 27.550 113.465 28.350 113.635 ;
        RECT 28.940 113.675 29.810 114.015 ;
        RECT 25.270 112.455 25.680 113.005 ;
        RECT 27.550 112.845 27.720 113.465 ;
        RECT 28.940 113.295 29.110 113.675 ;
        RECT 30.045 113.555 30.215 114.015 ;
        RECT 30.385 113.725 30.755 114.185 ;
        RECT 31.050 113.585 31.220 113.925 ;
        RECT 31.390 113.755 31.720 114.185 ;
        RECT 31.955 113.585 32.125 113.925 ;
        RECT 27.890 113.125 29.110 113.295 ;
        RECT 29.280 113.215 29.740 113.505 ;
        RECT 30.045 113.385 30.605 113.555 ;
        RECT 31.050 113.415 32.125 113.585 ;
        RECT 32.295 113.685 32.975 114.015 ;
        RECT 33.190 113.685 33.440 114.015 ;
        RECT 33.610 113.725 33.860 114.185 ;
        RECT 30.435 113.245 30.605 113.385 ;
        RECT 29.280 113.205 30.245 113.215 ;
        RECT 28.940 113.035 29.110 113.125 ;
        RECT 29.570 113.045 30.245 113.205 ;
        RECT 27.550 112.835 27.895 112.845 ;
        RECT 25.865 112.625 27.895 112.835 ;
        RECT 25.270 112.285 27.035 112.455 ;
        RECT 25.525 111.635 25.695 112.105 ;
        RECT 25.865 111.805 26.195 112.285 ;
        RECT 26.365 111.635 26.535 112.105 ;
        RECT 26.705 111.805 27.035 112.285 ;
        RECT 27.205 111.635 27.375 112.445 ;
        RECT 27.570 112.370 27.895 112.625 ;
        RECT 27.575 112.015 27.895 112.370 ;
        RECT 28.065 112.585 28.605 112.955 ;
        RECT 28.940 112.865 29.345 113.035 ;
        RECT 28.065 112.185 28.305 112.585 ;
        RECT 28.785 112.415 29.005 112.695 ;
        RECT 28.475 112.245 29.005 112.415 ;
        RECT 28.475 112.015 28.645 112.245 ;
        RECT 29.175 112.085 29.345 112.865 ;
        RECT 29.515 112.255 29.865 112.875 ;
        RECT 30.035 112.255 30.245 113.045 ;
        RECT 30.435 113.075 31.935 113.245 ;
        RECT 30.435 112.385 30.605 113.075 ;
        RECT 32.295 112.905 32.465 113.685 ;
        RECT 33.270 113.555 33.440 113.685 ;
        RECT 30.775 112.735 32.465 112.905 ;
        RECT 32.635 113.125 33.100 113.515 ;
        RECT 33.270 113.385 33.665 113.555 ;
        RECT 30.775 112.555 30.945 112.735 ;
        RECT 27.575 111.845 28.645 112.015 ;
        RECT 28.815 111.635 29.005 112.075 ;
        RECT 29.175 111.805 30.125 112.085 ;
        RECT 30.435 111.995 30.695 112.385 ;
        RECT 31.115 112.315 31.905 112.565 ;
        RECT 30.345 111.825 30.695 111.995 ;
        RECT 30.905 111.635 31.235 112.095 ;
        RECT 32.110 112.025 32.280 112.735 ;
        RECT 32.635 112.535 32.805 113.125 ;
        RECT 32.450 112.315 32.805 112.535 ;
        RECT 32.975 112.315 33.325 112.935 ;
        RECT 33.495 112.025 33.665 113.385 ;
        RECT 34.030 113.215 34.355 114.000 ;
        RECT 33.835 112.165 34.295 113.215 ;
        RECT 32.110 111.855 32.965 112.025 ;
        RECT 33.170 111.855 33.665 112.025 ;
        RECT 33.835 111.635 34.165 111.995 ;
        RECT 34.525 111.895 34.695 114.015 ;
        RECT 34.865 113.685 35.195 114.185 ;
        RECT 35.365 113.515 35.620 114.015 ;
        RECT 34.870 113.345 35.620 113.515 ;
        RECT 34.870 112.355 35.100 113.345 ;
        RECT 35.270 112.525 35.620 113.175 ;
        RECT 35.795 113.020 36.085 114.185 ;
        RECT 37.235 113.045 37.445 114.185 ;
        RECT 37.615 113.035 37.945 114.015 ;
        RECT 38.115 113.045 38.345 114.185 ;
        RECT 38.555 113.095 40.225 114.185 ;
        RECT 40.395 113.110 40.665 114.015 ;
        RECT 40.835 113.425 41.165 114.185 ;
        RECT 41.345 113.255 41.515 114.015 ;
        RECT 34.870 112.185 35.620 112.355 ;
        RECT 34.865 111.635 35.195 112.015 ;
        RECT 35.365 111.895 35.620 112.185 ;
        RECT 35.795 111.635 36.085 112.360 ;
        RECT 37.235 111.635 37.445 112.455 ;
        RECT 37.615 112.435 37.865 113.035 ;
        RECT 38.035 112.625 38.365 112.875 ;
        RECT 38.555 112.575 39.305 113.095 ;
        RECT 37.615 111.805 37.945 112.435 ;
        RECT 38.115 111.635 38.345 112.455 ;
        RECT 39.475 112.405 40.225 112.925 ;
        RECT 38.555 111.635 40.225 112.405 ;
        RECT 40.395 112.310 40.565 113.110 ;
        RECT 40.850 113.085 41.515 113.255 ;
        RECT 42.325 113.255 42.495 114.015 ;
        RECT 42.675 113.425 43.005 114.185 ;
        RECT 42.325 113.085 42.990 113.255 ;
        RECT 43.175 113.110 43.445 114.015 ;
        RECT 43.925 113.345 44.095 114.185 ;
        RECT 44.305 113.175 44.555 114.015 ;
        RECT 44.765 113.345 44.935 114.185 ;
        RECT 45.105 113.175 45.395 114.015 ;
        RECT 40.850 112.940 41.020 113.085 ;
        RECT 40.735 112.610 41.020 112.940 ;
        RECT 42.820 112.940 42.990 113.085 ;
        RECT 40.850 112.355 41.020 112.610 ;
        RECT 41.255 112.535 41.585 112.905 ;
        RECT 42.255 112.535 42.585 112.905 ;
        RECT 42.820 112.610 43.105 112.940 ;
        RECT 42.820 112.355 42.990 112.610 ;
        RECT 40.395 111.805 40.655 112.310 ;
        RECT 40.850 112.185 41.515 112.355 ;
        RECT 40.835 111.635 41.165 112.015 ;
        RECT 41.345 111.805 41.515 112.185 ;
        RECT 42.325 112.185 42.990 112.355 ;
        RECT 43.275 112.310 43.445 113.110 ;
        RECT 42.325 111.805 42.495 112.185 ;
        RECT 42.675 111.635 43.005 112.015 ;
        RECT 43.185 111.805 43.445 112.310 ;
        RECT 43.670 113.005 45.395 113.175 ;
        RECT 45.605 113.125 45.775 114.185 ;
        RECT 46.070 113.805 46.400 114.185 ;
        RECT 46.580 113.635 46.750 113.925 ;
        RECT 46.920 113.725 47.170 114.185 ;
        RECT 45.950 113.465 46.750 113.635 ;
        RECT 47.340 113.675 48.210 114.015 ;
        RECT 43.670 112.455 44.080 113.005 ;
        RECT 45.950 112.845 46.120 113.465 ;
        RECT 47.340 113.295 47.510 113.675 ;
        RECT 48.445 113.555 48.615 114.015 ;
        RECT 48.785 113.725 49.155 114.185 ;
        RECT 49.450 113.585 49.620 113.925 ;
        RECT 49.790 113.755 50.120 114.185 ;
        RECT 50.355 113.585 50.525 113.925 ;
        RECT 46.290 113.125 47.510 113.295 ;
        RECT 47.680 113.215 48.140 113.505 ;
        RECT 48.445 113.385 49.005 113.555 ;
        RECT 49.450 113.415 50.525 113.585 ;
        RECT 50.695 113.685 51.375 114.015 ;
        RECT 51.590 113.685 51.840 114.015 ;
        RECT 52.010 113.725 52.260 114.185 ;
        RECT 48.835 113.245 49.005 113.385 ;
        RECT 47.680 113.205 48.645 113.215 ;
        RECT 47.340 113.035 47.510 113.125 ;
        RECT 47.970 113.045 48.645 113.205 ;
        RECT 45.950 112.835 46.295 112.845 ;
        RECT 44.265 112.625 46.295 112.835 ;
        RECT 43.670 112.285 45.435 112.455 ;
        RECT 43.925 111.635 44.095 112.105 ;
        RECT 44.265 111.805 44.595 112.285 ;
        RECT 44.765 111.635 44.935 112.105 ;
        RECT 45.105 111.805 45.435 112.285 ;
        RECT 45.605 111.635 45.775 112.445 ;
        RECT 45.970 112.370 46.295 112.625 ;
        RECT 45.975 112.015 46.295 112.370 ;
        RECT 46.465 112.585 47.005 112.955 ;
        RECT 47.340 112.865 47.745 113.035 ;
        RECT 46.465 112.185 46.705 112.585 ;
        RECT 47.185 112.415 47.405 112.695 ;
        RECT 46.875 112.245 47.405 112.415 ;
        RECT 46.875 112.015 47.045 112.245 ;
        RECT 47.575 112.085 47.745 112.865 ;
        RECT 47.915 112.255 48.265 112.875 ;
        RECT 48.435 112.255 48.645 113.045 ;
        RECT 48.835 113.075 50.335 113.245 ;
        RECT 48.835 112.385 49.005 113.075 ;
        RECT 50.695 112.905 50.865 113.685 ;
        RECT 51.670 113.555 51.840 113.685 ;
        RECT 49.175 112.735 50.865 112.905 ;
        RECT 51.035 113.125 51.500 113.515 ;
        RECT 51.670 113.385 52.065 113.555 ;
        RECT 49.175 112.555 49.345 112.735 ;
        RECT 45.975 111.845 47.045 112.015 ;
        RECT 47.215 111.635 47.405 112.075 ;
        RECT 47.575 111.805 48.525 112.085 ;
        RECT 48.835 111.995 49.095 112.385 ;
        RECT 49.515 112.315 50.305 112.565 ;
        RECT 48.745 111.825 49.095 111.995 ;
        RECT 49.305 111.635 49.635 112.095 ;
        RECT 50.510 112.025 50.680 112.735 ;
        RECT 51.035 112.535 51.205 113.125 ;
        RECT 50.850 112.315 51.205 112.535 ;
        RECT 51.375 112.315 51.725 112.935 ;
        RECT 51.895 112.025 52.065 113.385 ;
        RECT 52.430 113.215 52.755 114.000 ;
        RECT 52.235 112.165 52.695 113.215 ;
        RECT 50.510 111.855 51.365 112.025 ;
        RECT 51.570 111.855 52.065 112.025 ;
        RECT 52.235 111.635 52.565 111.995 ;
        RECT 52.925 111.895 53.095 114.015 ;
        RECT 53.265 113.685 53.595 114.185 ;
        RECT 53.765 113.515 54.020 114.015 ;
        RECT 53.270 113.345 54.020 113.515 ;
        RECT 53.270 112.355 53.500 113.345 ;
        RECT 54.285 113.255 54.455 114.015 ;
        RECT 54.635 113.425 54.965 114.185 ;
        RECT 53.670 112.525 54.020 113.175 ;
        RECT 54.285 113.085 54.950 113.255 ;
        RECT 55.135 113.110 55.405 114.015 ;
        RECT 54.780 112.940 54.950 113.085 ;
        RECT 54.215 112.535 54.545 112.905 ;
        RECT 54.780 112.610 55.065 112.940 ;
        RECT 54.780 112.355 54.950 112.610 ;
        RECT 53.270 112.185 54.020 112.355 ;
        RECT 53.265 111.635 53.595 112.015 ;
        RECT 53.765 111.895 54.020 112.185 ;
        RECT 54.285 112.185 54.950 112.355 ;
        RECT 55.235 112.310 55.405 113.110 ;
        RECT 56.535 113.045 56.765 114.185 ;
        RECT 56.935 113.035 57.265 114.015 ;
        RECT 57.435 113.045 57.645 114.185 ;
        RECT 57.915 113.045 58.145 114.185 ;
        RECT 58.315 113.035 58.645 114.015 ;
        RECT 58.815 113.045 59.025 114.185 ;
        RECT 59.715 113.110 59.985 114.015 ;
        RECT 60.155 113.425 60.485 114.185 ;
        RECT 60.665 113.255 60.835 114.015 ;
        RECT 56.515 112.625 56.845 112.875 ;
        RECT 54.285 111.805 54.455 112.185 ;
        RECT 54.635 111.635 54.965 112.015 ;
        RECT 55.145 111.805 55.405 112.310 ;
        RECT 56.535 111.635 56.765 112.455 ;
        RECT 57.015 112.435 57.265 113.035 ;
        RECT 57.895 112.625 58.225 112.875 ;
        RECT 56.935 111.805 57.265 112.435 ;
        RECT 57.435 111.635 57.645 112.455 ;
        RECT 57.915 111.635 58.145 112.455 ;
        RECT 58.395 112.435 58.645 113.035 ;
        RECT 58.315 111.805 58.645 112.435 ;
        RECT 58.815 111.635 59.025 112.455 ;
        RECT 59.715 112.310 59.885 113.110 ;
        RECT 60.170 113.085 60.835 113.255 ;
        RECT 60.170 112.940 60.340 113.085 ;
        RECT 61.555 113.020 61.845 114.185 ;
        RECT 63.025 113.255 63.195 114.015 ;
        RECT 63.375 113.425 63.705 114.185 ;
        RECT 63.025 113.085 63.690 113.255 ;
        RECT 63.875 113.110 64.145 114.015 ;
        RECT 64.625 113.345 64.795 114.185 ;
        RECT 65.005 113.175 65.255 114.015 ;
        RECT 65.465 113.345 65.635 114.185 ;
        RECT 65.805 113.175 66.095 114.015 ;
        RECT 60.055 112.610 60.340 112.940 ;
        RECT 63.520 112.940 63.690 113.085 ;
        RECT 60.170 112.355 60.340 112.610 ;
        RECT 60.575 112.535 60.905 112.905 ;
        RECT 62.955 112.535 63.285 112.905 ;
        RECT 63.520 112.610 63.805 112.940 ;
        RECT 59.715 111.805 59.975 112.310 ;
        RECT 60.170 112.185 60.835 112.355 ;
        RECT 60.155 111.635 60.485 112.015 ;
        RECT 60.665 111.805 60.835 112.185 ;
        RECT 61.555 111.635 61.845 112.360 ;
        RECT 63.520 112.355 63.690 112.610 ;
        RECT 63.025 112.185 63.690 112.355 ;
        RECT 63.975 112.310 64.145 113.110 ;
        RECT 63.025 111.805 63.195 112.185 ;
        RECT 63.375 111.635 63.705 112.015 ;
        RECT 63.885 111.805 64.145 112.310 ;
        RECT 64.370 113.005 66.095 113.175 ;
        RECT 66.305 113.125 66.475 114.185 ;
        RECT 66.770 113.805 67.100 114.185 ;
        RECT 67.280 113.635 67.450 113.925 ;
        RECT 67.620 113.725 67.870 114.185 ;
        RECT 66.650 113.465 67.450 113.635 ;
        RECT 68.040 113.675 68.910 114.015 ;
        RECT 64.370 112.455 64.780 113.005 ;
        RECT 66.650 112.845 66.820 113.465 ;
        RECT 68.040 113.295 68.210 113.675 ;
        RECT 69.145 113.555 69.315 114.015 ;
        RECT 69.485 113.725 69.855 114.185 ;
        RECT 70.150 113.585 70.320 113.925 ;
        RECT 70.490 113.755 70.820 114.185 ;
        RECT 71.055 113.585 71.225 113.925 ;
        RECT 66.990 113.125 68.210 113.295 ;
        RECT 68.380 113.215 68.840 113.505 ;
        RECT 69.145 113.385 69.705 113.555 ;
        RECT 70.150 113.415 71.225 113.585 ;
        RECT 71.395 113.685 72.075 114.015 ;
        RECT 72.290 113.685 72.540 114.015 ;
        RECT 72.710 113.725 72.960 114.185 ;
        RECT 69.535 113.245 69.705 113.385 ;
        RECT 68.380 113.205 69.345 113.215 ;
        RECT 68.040 113.035 68.210 113.125 ;
        RECT 68.670 113.045 69.345 113.205 ;
        RECT 66.650 112.835 66.995 112.845 ;
        RECT 64.965 112.625 66.995 112.835 ;
        RECT 64.370 112.285 66.135 112.455 ;
        RECT 64.625 111.635 64.795 112.105 ;
        RECT 64.965 111.805 65.295 112.285 ;
        RECT 65.465 111.635 65.635 112.105 ;
        RECT 65.805 111.805 66.135 112.285 ;
        RECT 66.305 111.635 66.475 112.445 ;
        RECT 66.670 112.370 66.995 112.625 ;
        RECT 66.675 112.015 66.995 112.370 ;
        RECT 67.165 112.585 67.705 112.955 ;
        RECT 68.040 112.865 68.445 113.035 ;
        RECT 67.165 112.185 67.405 112.585 ;
        RECT 67.885 112.415 68.105 112.695 ;
        RECT 67.575 112.245 68.105 112.415 ;
        RECT 67.575 112.015 67.745 112.245 ;
        RECT 68.275 112.085 68.445 112.865 ;
        RECT 68.615 112.255 68.965 112.875 ;
        RECT 69.135 112.255 69.345 113.045 ;
        RECT 69.535 113.075 71.035 113.245 ;
        RECT 69.535 112.385 69.705 113.075 ;
        RECT 71.395 112.905 71.565 113.685 ;
        RECT 72.370 113.555 72.540 113.685 ;
        RECT 69.875 112.735 71.565 112.905 ;
        RECT 71.735 113.125 72.200 113.515 ;
        RECT 72.370 113.385 72.765 113.555 ;
        RECT 69.875 112.555 70.045 112.735 ;
        RECT 66.675 111.845 67.745 112.015 ;
        RECT 67.915 111.635 68.105 112.075 ;
        RECT 68.275 111.805 69.225 112.085 ;
        RECT 69.535 111.995 69.795 112.385 ;
        RECT 70.215 112.315 71.005 112.565 ;
        RECT 69.445 111.825 69.795 111.995 ;
        RECT 70.005 111.635 70.335 112.095 ;
        RECT 71.210 112.025 71.380 112.735 ;
        RECT 71.735 112.535 71.905 113.125 ;
        RECT 71.550 112.315 71.905 112.535 ;
        RECT 72.075 112.315 72.425 112.935 ;
        RECT 72.595 112.025 72.765 113.385 ;
        RECT 73.130 113.215 73.455 114.000 ;
        RECT 72.935 112.165 73.395 113.215 ;
        RECT 71.210 111.855 72.065 112.025 ;
        RECT 72.270 111.855 72.765 112.025 ;
        RECT 72.935 111.635 73.265 111.995 ;
        RECT 73.625 111.895 73.795 114.015 ;
        RECT 73.965 113.685 74.295 114.185 ;
        RECT 74.465 113.515 74.720 114.015 ;
        RECT 73.970 113.345 74.720 113.515 ;
        RECT 75.205 113.345 75.375 114.185 ;
        RECT 73.970 112.355 74.200 113.345 ;
        RECT 75.585 113.175 75.835 114.015 ;
        RECT 76.045 113.345 76.215 114.185 ;
        RECT 76.385 113.175 76.675 114.015 ;
        RECT 74.370 112.525 74.720 113.175 ;
        RECT 74.950 113.005 76.675 113.175 ;
        RECT 76.885 113.125 77.055 114.185 ;
        RECT 77.350 113.805 77.680 114.185 ;
        RECT 77.860 113.635 78.030 113.925 ;
        RECT 78.200 113.725 78.450 114.185 ;
        RECT 77.230 113.465 78.030 113.635 ;
        RECT 78.620 113.675 79.490 114.015 ;
        RECT 74.950 112.455 75.360 113.005 ;
        RECT 77.230 112.845 77.400 113.465 ;
        RECT 78.620 113.295 78.790 113.675 ;
        RECT 79.725 113.555 79.895 114.015 ;
        RECT 80.065 113.725 80.435 114.185 ;
        RECT 80.730 113.585 80.900 113.925 ;
        RECT 81.070 113.755 81.400 114.185 ;
        RECT 81.635 113.585 81.805 113.925 ;
        RECT 77.570 113.125 78.790 113.295 ;
        RECT 78.960 113.215 79.420 113.505 ;
        RECT 79.725 113.385 80.285 113.555 ;
        RECT 80.730 113.415 81.805 113.585 ;
        RECT 81.975 113.685 82.655 114.015 ;
        RECT 82.870 113.685 83.120 114.015 ;
        RECT 83.290 113.725 83.540 114.185 ;
        RECT 80.115 113.245 80.285 113.385 ;
        RECT 78.960 113.205 79.925 113.215 ;
        RECT 78.620 113.035 78.790 113.125 ;
        RECT 79.250 113.045 79.925 113.205 ;
        RECT 77.230 112.835 77.575 112.845 ;
        RECT 75.545 112.625 77.575 112.835 ;
        RECT 73.970 112.185 74.720 112.355 ;
        RECT 74.950 112.285 76.715 112.455 ;
        RECT 73.965 111.635 74.295 112.015 ;
        RECT 74.465 111.895 74.720 112.185 ;
        RECT 75.205 111.635 75.375 112.105 ;
        RECT 75.545 111.805 75.875 112.285 ;
        RECT 76.045 111.635 76.215 112.105 ;
        RECT 76.385 111.805 76.715 112.285 ;
        RECT 76.885 111.635 77.055 112.445 ;
        RECT 77.250 112.370 77.575 112.625 ;
        RECT 77.255 112.015 77.575 112.370 ;
        RECT 77.745 112.585 78.285 112.955 ;
        RECT 78.620 112.865 79.025 113.035 ;
        RECT 77.745 112.185 77.985 112.585 ;
        RECT 78.465 112.415 78.685 112.695 ;
        RECT 78.155 112.245 78.685 112.415 ;
        RECT 78.155 112.015 78.325 112.245 ;
        RECT 78.855 112.085 79.025 112.865 ;
        RECT 79.195 112.255 79.545 112.875 ;
        RECT 79.715 112.255 79.925 113.045 ;
        RECT 80.115 113.075 81.615 113.245 ;
        RECT 80.115 112.385 80.285 113.075 ;
        RECT 81.975 112.905 82.145 113.685 ;
        RECT 82.950 113.555 83.120 113.685 ;
        RECT 80.455 112.735 82.145 112.905 ;
        RECT 82.315 113.125 82.780 113.515 ;
        RECT 82.950 113.385 83.345 113.555 ;
        RECT 80.455 112.555 80.625 112.735 ;
        RECT 77.255 111.845 78.325 112.015 ;
        RECT 78.495 111.635 78.685 112.075 ;
        RECT 78.855 111.805 79.805 112.085 ;
        RECT 80.115 111.995 80.375 112.385 ;
        RECT 80.795 112.315 81.585 112.565 ;
        RECT 80.025 111.825 80.375 111.995 ;
        RECT 80.585 111.635 80.915 112.095 ;
        RECT 81.790 112.025 81.960 112.735 ;
        RECT 82.315 112.535 82.485 113.125 ;
        RECT 82.130 112.315 82.485 112.535 ;
        RECT 82.655 112.315 83.005 112.935 ;
        RECT 83.175 112.025 83.345 113.385 ;
        RECT 83.710 113.215 84.035 114.000 ;
        RECT 83.515 112.165 83.975 113.215 ;
        RECT 81.790 111.855 82.645 112.025 ;
        RECT 82.850 111.855 83.345 112.025 ;
        RECT 83.515 111.635 83.845 111.995 ;
        RECT 84.205 111.895 84.375 114.015 ;
        RECT 84.545 113.685 84.875 114.185 ;
        RECT 85.045 113.515 85.300 114.015 ;
        RECT 84.550 113.345 85.300 113.515 ;
        RECT 84.550 112.355 84.780 113.345 ;
        RECT 84.950 112.525 85.300 113.175 ;
        RECT 85.475 113.110 85.745 114.015 ;
        RECT 85.915 113.425 86.245 114.185 ;
        RECT 86.425 113.255 86.595 114.015 ;
        RECT 84.550 112.185 85.300 112.355 ;
        RECT 84.545 111.635 84.875 112.015 ;
        RECT 85.045 111.895 85.300 112.185 ;
        RECT 85.475 112.310 85.645 113.110 ;
        RECT 85.930 113.085 86.595 113.255 ;
        RECT 85.930 112.940 86.100 113.085 ;
        RECT 87.315 113.020 87.605 114.185 ;
        RECT 89.005 113.345 89.175 114.185 ;
        RECT 89.385 113.175 89.635 114.015 ;
        RECT 89.845 113.345 90.015 114.185 ;
        RECT 90.185 113.175 90.475 114.015 ;
        RECT 85.815 112.610 86.100 112.940 ;
        RECT 88.750 113.005 90.475 113.175 ;
        RECT 90.685 113.125 90.855 114.185 ;
        RECT 91.150 113.805 91.480 114.185 ;
        RECT 91.660 113.635 91.830 113.925 ;
        RECT 92.000 113.725 92.250 114.185 ;
        RECT 91.030 113.465 91.830 113.635 ;
        RECT 92.420 113.675 93.290 114.015 ;
        RECT 85.930 112.355 86.100 112.610 ;
        RECT 86.335 112.535 86.665 112.905 ;
        RECT 88.750 112.455 89.160 113.005 ;
        RECT 91.030 112.845 91.200 113.465 ;
        RECT 92.420 113.295 92.590 113.675 ;
        RECT 93.525 113.555 93.695 114.015 ;
        RECT 93.865 113.725 94.235 114.185 ;
        RECT 94.530 113.585 94.700 113.925 ;
        RECT 94.870 113.755 95.200 114.185 ;
        RECT 95.435 113.585 95.605 113.925 ;
        RECT 91.370 113.125 92.590 113.295 ;
        RECT 92.760 113.215 93.220 113.505 ;
        RECT 93.525 113.385 94.085 113.555 ;
        RECT 94.530 113.415 95.605 113.585 ;
        RECT 95.775 113.685 96.455 114.015 ;
        RECT 96.670 113.685 96.920 114.015 ;
        RECT 97.090 113.725 97.340 114.185 ;
        RECT 93.915 113.245 94.085 113.385 ;
        RECT 92.760 113.205 93.725 113.215 ;
        RECT 92.420 113.035 92.590 113.125 ;
        RECT 93.050 113.045 93.725 113.205 ;
        RECT 91.030 112.835 91.375 112.845 ;
        RECT 89.345 112.625 91.375 112.835 ;
        RECT 85.475 111.805 85.735 112.310 ;
        RECT 85.930 112.185 86.595 112.355 ;
        RECT 85.915 111.635 86.245 112.015 ;
        RECT 86.425 111.805 86.595 112.185 ;
        RECT 87.315 111.635 87.605 112.360 ;
        RECT 88.750 112.285 90.515 112.455 ;
        RECT 89.005 111.635 89.175 112.105 ;
        RECT 89.345 111.805 89.675 112.285 ;
        RECT 89.845 111.635 90.015 112.105 ;
        RECT 90.185 111.805 90.515 112.285 ;
        RECT 90.685 111.635 90.855 112.445 ;
        RECT 91.050 112.370 91.375 112.625 ;
        RECT 91.055 112.015 91.375 112.370 ;
        RECT 91.545 112.585 92.085 112.955 ;
        RECT 92.420 112.865 92.825 113.035 ;
        RECT 91.545 112.185 91.785 112.585 ;
        RECT 92.265 112.415 92.485 112.695 ;
        RECT 91.955 112.245 92.485 112.415 ;
        RECT 91.955 112.015 92.125 112.245 ;
        RECT 92.655 112.085 92.825 112.865 ;
        RECT 92.995 112.255 93.345 112.875 ;
        RECT 93.515 112.255 93.725 113.045 ;
        RECT 93.915 113.075 95.415 113.245 ;
        RECT 93.915 112.385 94.085 113.075 ;
        RECT 95.775 112.905 95.945 113.685 ;
        RECT 96.750 113.555 96.920 113.685 ;
        RECT 94.255 112.735 95.945 112.905 ;
        RECT 96.115 113.125 96.580 113.515 ;
        RECT 96.750 113.385 97.145 113.555 ;
        RECT 94.255 112.555 94.425 112.735 ;
        RECT 91.055 111.845 92.125 112.015 ;
        RECT 92.295 111.635 92.485 112.075 ;
        RECT 92.655 111.805 93.605 112.085 ;
        RECT 93.915 111.995 94.175 112.385 ;
        RECT 94.595 112.315 95.385 112.565 ;
        RECT 93.825 111.825 94.175 111.995 ;
        RECT 94.385 111.635 94.715 112.095 ;
        RECT 95.590 112.025 95.760 112.735 ;
        RECT 96.115 112.535 96.285 113.125 ;
        RECT 95.930 112.315 96.285 112.535 ;
        RECT 96.455 112.315 96.805 112.935 ;
        RECT 96.975 112.025 97.145 113.385 ;
        RECT 97.510 113.215 97.835 114.000 ;
        RECT 97.315 112.165 97.775 113.215 ;
        RECT 95.590 111.855 96.445 112.025 ;
        RECT 96.650 111.855 97.145 112.025 ;
        RECT 97.315 111.635 97.645 111.995 ;
        RECT 98.005 111.895 98.175 114.015 ;
        RECT 98.345 113.685 98.675 114.185 ;
        RECT 98.845 113.515 99.100 114.015 ;
        RECT 98.350 113.345 99.100 113.515 ;
        RECT 98.350 112.355 98.580 113.345 ;
        RECT 98.750 112.525 99.100 113.175 ;
        RECT 99.275 113.110 99.545 114.015 ;
        RECT 99.715 113.425 100.045 114.185 ;
        RECT 100.225 113.255 100.395 114.015 ;
        RECT 101.885 113.345 102.055 114.185 ;
        RECT 98.350 112.185 99.100 112.355 ;
        RECT 98.345 111.635 98.675 112.015 ;
        RECT 98.845 111.895 99.100 112.185 ;
        RECT 99.275 112.310 99.445 113.110 ;
        RECT 99.730 113.085 100.395 113.255 ;
        RECT 102.265 113.175 102.515 114.015 ;
        RECT 102.725 113.345 102.895 114.185 ;
        RECT 103.065 113.175 103.355 114.015 ;
        RECT 99.730 112.940 99.900 113.085 ;
        RECT 99.615 112.610 99.900 112.940 ;
        RECT 101.630 113.005 103.355 113.175 ;
        RECT 103.565 113.125 103.735 114.185 ;
        RECT 104.030 113.805 104.360 114.185 ;
        RECT 104.540 113.635 104.710 113.925 ;
        RECT 104.880 113.725 105.130 114.185 ;
        RECT 103.910 113.465 104.710 113.635 ;
        RECT 105.300 113.675 106.170 114.015 ;
        RECT 99.730 112.355 99.900 112.610 ;
        RECT 100.135 112.535 100.465 112.905 ;
        RECT 101.630 112.455 102.040 113.005 ;
        RECT 103.910 112.845 104.080 113.465 ;
        RECT 105.300 113.295 105.470 113.675 ;
        RECT 106.405 113.555 106.575 114.015 ;
        RECT 106.745 113.725 107.115 114.185 ;
        RECT 107.410 113.585 107.580 113.925 ;
        RECT 107.750 113.755 108.080 114.185 ;
        RECT 108.315 113.585 108.485 113.925 ;
        RECT 104.250 113.125 105.470 113.295 ;
        RECT 105.640 113.215 106.100 113.505 ;
        RECT 106.405 113.385 106.965 113.555 ;
        RECT 107.410 113.415 108.485 113.585 ;
        RECT 108.655 113.685 109.335 114.015 ;
        RECT 109.550 113.685 109.800 114.015 ;
        RECT 109.970 113.725 110.220 114.185 ;
        RECT 106.795 113.245 106.965 113.385 ;
        RECT 105.640 113.205 106.605 113.215 ;
        RECT 105.300 113.035 105.470 113.125 ;
        RECT 105.930 113.045 106.605 113.205 ;
        RECT 103.910 112.835 104.255 112.845 ;
        RECT 102.225 112.625 104.255 112.835 ;
        RECT 99.275 111.805 99.535 112.310 ;
        RECT 99.730 112.185 100.395 112.355 ;
        RECT 101.630 112.285 103.395 112.455 ;
        RECT 99.715 111.635 100.045 112.015 ;
        RECT 100.225 111.805 100.395 112.185 ;
        RECT 101.885 111.635 102.055 112.105 ;
        RECT 102.225 111.805 102.555 112.285 ;
        RECT 102.725 111.635 102.895 112.105 ;
        RECT 103.065 111.805 103.395 112.285 ;
        RECT 103.565 111.635 103.735 112.445 ;
        RECT 103.930 112.370 104.255 112.625 ;
        RECT 103.935 112.015 104.255 112.370 ;
        RECT 104.425 112.585 104.965 112.955 ;
        RECT 105.300 112.865 105.705 113.035 ;
        RECT 104.425 112.185 104.665 112.585 ;
        RECT 105.145 112.415 105.365 112.695 ;
        RECT 104.835 112.245 105.365 112.415 ;
        RECT 104.835 112.015 105.005 112.245 ;
        RECT 105.535 112.085 105.705 112.865 ;
        RECT 105.875 112.255 106.225 112.875 ;
        RECT 106.395 112.255 106.605 113.045 ;
        RECT 106.795 113.075 108.295 113.245 ;
        RECT 106.795 112.385 106.965 113.075 ;
        RECT 108.655 112.905 108.825 113.685 ;
        RECT 109.630 113.555 109.800 113.685 ;
        RECT 107.135 112.735 108.825 112.905 ;
        RECT 108.995 113.125 109.460 113.515 ;
        RECT 109.630 113.385 110.025 113.555 ;
        RECT 107.135 112.555 107.305 112.735 ;
        RECT 103.935 111.845 105.005 112.015 ;
        RECT 105.175 111.635 105.365 112.075 ;
        RECT 105.535 111.805 106.485 112.085 ;
        RECT 106.795 111.995 107.055 112.385 ;
        RECT 107.475 112.315 108.265 112.565 ;
        RECT 106.705 111.825 107.055 111.995 ;
        RECT 107.265 111.635 107.595 112.095 ;
        RECT 108.470 112.025 108.640 112.735 ;
        RECT 108.995 112.535 109.165 113.125 ;
        RECT 108.810 112.315 109.165 112.535 ;
        RECT 109.335 112.315 109.685 112.935 ;
        RECT 109.855 112.025 110.025 113.385 ;
        RECT 110.390 113.215 110.715 114.000 ;
        RECT 110.195 112.165 110.655 113.215 ;
        RECT 108.470 111.855 109.325 112.025 ;
        RECT 109.530 111.855 110.025 112.025 ;
        RECT 110.195 111.635 110.525 111.995 ;
        RECT 110.885 111.895 111.055 114.015 ;
        RECT 111.225 113.685 111.555 114.185 ;
        RECT 111.725 113.515 111.980 114.015 ;
        RECT 111.230 113.345 111.980 113.515 ;
        RECT 111.230 112.355 111.460 113.345 ;
        RECT 111.630 112.525 111.980 113.175 ;
        RECT 112.155 113.095 113.365 114.185 ;
        RECT 112.155 112.555 112.675 113.095 ;
        RECT 112.845 112.385 113.365 112.925 ;
        RECT 111.230 112.185 111.980 112.355 ;
        RECT 111.225 111.635 111.555 112.015 ;
        RECT 111.725 111.895 111.980 112.185 ;
        RECT 112.155 111.635 113.365 112.385 ;
        RECT 15.010 111.465 113.450 111.635 ;
        RECT 15.095 110.715 16.305 111.465 ;
        RECT 15.095 110.175 15.615 110.715 ;
        RECT 16.475 110.695 19.985 111.465 ;
        RECT 15.785 110.005 16.305 110.545 ;
        RECT 15.095 108.915 16.305 110.005 ;
        RECT 16.475 110.005 18.165 110.525 ;
        RECT 18.335 110.175 19.985 110.695 ;
        RECT 20.215 110.645 20.425 111.465 ;
        RECT 20.595 110.665 20.925 111.295 ;
        RECT 20.595 110.065 20.845 110.665 ;
        RECT 21.095 110.645 21.325 111.465 ;
        RECT 21.575 110.645 21.805 111.465 ;
        RECT 21.975 110.665 22.305 111.295 ;
        RECT 21.015 110.225 21.345 110.475 ;
        RECT 21.555 110.225 21.885 110.475 ;
        RECT 22.055 110.065 22.305 110.665 ;
        RECT 22.475 110.645 22.685 111.465 ;
        RECT 22.915 110.740 23.205 111.465 ;
        RECT 23.415 110.645 23.645 111.465 ;
        RECT 23.815 110.665 24.145 111.295 ;
        RECT 23.395 110.225 23.725 110.475 ;
        RECT 16.475 108.915 19.985 110.005 ;
        RECT 20.215 108.915 20.425 110.055 ;
        RECT 20.595 109.085 20.925 110.065 ;
        RECT 21.095 108.915 21.325 110.055 ;
        RECT 21.575 108.915 21.805 110.055 ;
        RECT 21.975 109.085 22.305 110.065 ;
        RECT 22.475 108.915 22.685 110.055 ;
        RECT 22.915 108.915 23.205 110.080 ;
        RECT 23.895 110.065 24.145 110.665 ;
        RECT 24.315 110.645 24.525 111.465 ;
        RECT 24.795 110.645 25.025 111.465 ;
        RECT 25.195 110.665 25.525 111.295 ;
        RECT 24.775 110.225 25.105 110.475 ;
        RECT 25.275 110.065 25.525 110.665 ;
        RECT 25.695 110.645 25.905 111.465 ;
        RECT 26.225 110.915 26.395 111.295 ;
        RECT 26.575 111.085 26.905 111.465 ;
        RECT 26.225 110.745 26.890 110.915 ;
        RECT 27.085 110.790 27.345 111.295 ;
        RECT 26.155 110.195 26.485 110.565 ;
        RECT 26.720 110.490 26.890 110.745 ;
        RECT 23.415 108.915 23.645 110.055 ;
        RECT 23.815 109.085 24.145 110.065 ;
        RECT 24.315 108.915 24.525 110.055 ;
        RECT 24.795 108.915 25.025 110.055 ;
        RECT 25.195 109.085 25.525 110.065 ;
        RECT 26.720 110.160 27.005 110.490 ;
        RECT 25.695 108.915 25.905 110.055 ;
        RECT 26.720 110.015 26.890 110.160 ;
        RECT 26.225 109.845 26.890 110.015 ;
        RECT 27.175 109.990 27.345 110.790 ;
        RECT 27.520 110.915 27.775 111.205 ;
        RECT 27.945 111.085 28.275 111.465 ;
        RECT 27.520 110.745 28.270 110.915 ;
        RECT 26.225 109.085 26.395 109.845 ;
        RECT 26.575 108.915 26.905 109.675 ;
        RECT 27.075 109.085 27.345 109.990 ;
        RECT 27.520 109.925 27.870 110.575 ;
        RECT 28.040 109.755 28.270 110.745 ;
        RECT 27.520 109.585 28.270 109.755 ;
        RECT 27.520 109.085 27.775 109.585 ;
        RECT 27.945 108.915 28.275 109.415 ;
        RECT 28.445 109.085 28.615 111.205 ;
        RECT 28.975 111.105 29.305 111.465 ;
        RECT 29.475 111.075 29.970 111.245 ;
        RECT 30.175 111.075 31.030 111.245 ;
        RECT 28.845 109.885 29.305 110.935 ;
        RECT 28.785 109.100 29.110 109.885 ;
        RECT 29.475 109.715 29.645 111.075 ;
        RECT 29.815 110.165 30.165 110.785 ;
        RECT 30.335 110.565 30.690 110.785 ;
        RECT 30.335 109.975 30.505 110.565 ;
        RECT 30.860 110.365 31.030 111.075 ;
        RECT 31.905 111.005 32.235 111.465 ;
        RECT 32.445 111.105 32.795 111.275 ;
        RECT 31.235 110.535 32.025 110.785 ;
        RECT 32.445 110.715 32.705 111.105 ;
        RECT 33.015 111.015 33.965 111.295 ;
        RECT 34.135 111.025 34.325 111.465 ;
        RECT 34.495 111.085 35.565 111.255 ;
        RECT 32.195 110.365 32.365 110.545 ;
        RECT 29.475 109.545 29.870 109.715 ;
        RECT 30.040 109.585 30.505 109.975 ;
        RECT 30.675 110.195 32.365 110.365 ;
        RECT 29.700 109.415 29.870 109.545 ;
        RECT 30.675 109.415 30.845 110.195 ;
        RECT 32.535 110.025 32.705 110.715 ;
        RECT 31.205 109.855 32.705 110.025 ;
        RECT 32.895 110.055 33.105 110.845 ;
        RECT 33.275 110.225 33.625 110.845 ;
        RECT 33.795 110.235 33.965 111.015 ;
        RECT 34.495 110.855 34.665 111.085 ;
        RECT 34.135 110.685 34.665 110.855 ;
        RECT 34.135 110.405 34.355 110.685 ;
        RECT 34.835 110.515 35.075 110.915 ;
        RECT 33.795 110.065 34.200 110.235 ;
        RECT 34.535 110.145 35.075 110.515 ;
        RECT 35.245 110.730 35.565 111.085 ;
        RECT 35.245 110.475 35.570 110.730 ;
        RECT 35.765 110.655 35.935 111.465 ;
        RECT 36.105 110.815 36.435 111.295 ;
        RECT 36.605 110.995 36.775 111.465 ;
        RECT 36.945 110.815 37.275 111.295 ;
        RECT 37.445 110.995 37.615 111.465 ;
        RECT 38.405 110.995 38.575 111.465 ;
        RECT 38.745 110.815 39.075 111.295 ;
        RECT 39.245 110.995 39.415 111.465 ;
        RECT 39.585 110.815 39.915 111.295 ;
        RECT 36.105 110.645 37.870 110.815 ;
        RECT 35.245 110.265 37.275 110.475 ;
        RECT 35.245 110.255 35.590 110.265 ;
        RECT 32.895 109.895 33.570 110.055 ;
        RECT 34.030 109.975 34.200 110.065 ;
        RECT 32.895 109.885 33.860 109.895 ;
        RECT 32.535 109.715 32.705 109.855 ;
        RECT 29.280 108.915 29.530 109.375 ;
        RECT 29.700 109.085 29.950 109.415 ;
        RECT 30.165 109.085 30.845 109.415 ;
        RECT 31.015 109.515 32.090 109.685 ;
        RECT 32.535 109.545 33.095 109.715 ;
        RECT 33.400 109.595 33.860 109.885 ;
        RECT 34.030 109.805 35.250 109.975 ;
        RECT 31.015 109.175 31.185 109.515 ;
        RECT 31.420 108.915 31.750 109.345 ;
        RECT 31.920 109.175 32.090 109.515 ;
        RECT 32.385 108.915 32.755 109.375 ;
        RECT 32.925 109.085 33.095 109.545 ;
        RECT 34.030 109.425 34.200 109.805 ;
        RECT 35.420 109.635 35.590 110.255 ;
        RECT 37.460 110.095 37.870 110.645 ;
        RECT 33.330 109.085 34.200 109.425 ;
        RECT 34.790 109.465 35.590 109.635 ;
        RECT 34.370 108.915 34.620 109.375 ;
        RECT 34.790 109.175 34.960 109.465 ;
        RECT 35.140 108.915 35.470 109.295 ;
        RECT 35.765 108.915 35.935 109.975 ;
        RECT 36.145 109.925 37.870 110.095 ;
        RECT 38.150 110.645 39.915 110.815 ;
        RECT 40.085 110.655 40.255 111.465 ;
        RECT 40.455 111.085 41.525 111.255 ;
        RECT 40.455 110.730 40.775 111.085 ;
        RECT 38.150 110.095 38.560 110.645 ;
        RECT 40.450 110.475 40.775 110.730 ;
        RECT 38.745 110.265 40.775 110.475 ;
        RECT 40.430 110.255 40.775 110.265 ;
        RECT 40.945 110.515 41.185 110.915 ;
        RECT 41.355 110.855 41.525 111.085 ;
        RECT 41.695 111.025 41.885 111.465 ;
        RECT 42.055 111.015 43.005 111.295 ;
        RECT 43.225 111.105 43.575 111.275 ;
        RECT 41.355 110.685 41.885 110.855 ;
        RECT 38.150 109.925 39.875 110.095 ;
        RECT 36.145 109.085 36.435 109.925 ;
        RECT 36.605 108.915 36.775 109.755 ;
        RECT 36.985 109.085 37.235 109.925 ;
        RECT 37.445 108.915 37.615 109.755 ;
        RECT 38.405 108.915 38.575 109.755 ;
        RECT 38.785 109.085 39.035 109.925 ;
        RECT 39.245 108.915 39.415 109.755 ;
        RECT 39.585 109.085 39.875 109.925 ;
        RECT 40.085 108.915 40.255 109.975 ;
        RECT 40.430 109.635 40.600 110.255 ;
        RECT 40.945 110.145 41.485 110.515 ;
        RECT 41.665 110.405 41.885 110.685 ;
        RECT 42.055 110.235 42.225 111.015 ;
        RECT 41.820 110.065 42.225 110.235 ;
        RECT 42.395 110.225 42.745 110.845 ;
        RECT 41.820 109.975 41.990 110.065 ;
        RECT 42.915 110.055 43.125 110.845 ;
        RECT 40.770 109.805 41.990 109.975 ;
        RECT 42.450 109.895 43.125 110.055 ;
        RECT 40.430 109.465 41.230 109.635 ;
        RECT 40.550 108.915 40.880 109.295 ;
        RECT 41.060 109.175 41.230 109.465 ;
        RECT 41.820 109.425 41.990 109.805 ;
        RECT 42.160 109.885 43.125 109.895 ;
        RECT 43.315 110.715 43.575 111.105 ;
        RECT 43.785 111.005 44.115 111.465 ;
        RECT 44.990 111.075 45.845 111.245 ;
        RECT 46.050 111.075 46.545 111.245 ;
        RECT 46.715 111.105 47.045 111.465 ;
        RECT 43.315 110.025 43.485 110.715 ;
        RECT 43.655 110.365 43.825 110.545 ;
        RECT 43.995 110.535 44.785 110.785 ;
        RECT 44.990 110.365 45.160 111.075 ;
        RECT 45.330 110.565 45.685 110.785 ;
        RECT 43.655 110.195 45.345 110.365 ;
        RECT 42.160 109.595 42.620 109.885 ;
        RECT 43.315 109.855 44.815 110.025 ;
        RECT 43.315 109.715 43.485 109.855 ;
        RECT 42.925 109.545 43.485 109.715 ;
        RECT 41.400 108.915 41.650 109.375 ;
        RECT 41.820 109.085 42.690 109.425 ;
        RECT 42.925 109.085 43.095 109.545 ;
        RECT 43.930 109.515 45.005 109.685 ;
        RECT 43.265 108.915 43.635 109.375 ;
        RECT 43.930 109.175 44.100 109.515 ;
        RECT 44.270 108.915 44.600 109.345 ;
        RECT 44.835 109.175 45.005 109.515 ;
        RECT 45.175 109.415 45.345 110.195 ;
        RECT 45.515 109.975 45.685 110.565 ;
        RECT 45.855 110.165 46.205 110.785 ;
        RECT 45.515 109.585 45.980 109.975 ;
        RECT 46.375 109.715 46.545 111.075 ;
        RECT 46.715 109.885 47.175 110.935 ;
        RECT 46.150 109.545 46.545 109.715 ;
        RECT 46.150 109.415 46.320 109.545 ;
        RECT 45.175 109.085 45.855 109.415 ;
        RECT 46.070 109.085 46.320 109.415 ;
        RECT 46.490 108.915 46.740 109.375 ;
        RECT 46.910 109.100 47.235 109.885 ;
        RECT 47.405 109.085 47.575 111.205 ;
        RECT 47.745 111.085 48.075 111.465 ;
        RECT 48.245 110.915 48.500 111.205 ;
        RECT 47.750 110.745 48.500 110.915 ;
        RECT 47.750 109.755 47.980 110.745 ;
        RECT 48.675 110.740 48.965 111.465 ;
        RECT 49.445 110.995 49.615 111.465 ;
        RECT 49.785 110.815 50.115 111.295 ;
        RECT 50.285 110.995 50.455 111.465 ;
        RECT 50.625 110.815 50.955 111.295 ;
        RECT 49.190 110.645 50.955 110.815 ;
        RECT 51.125 110.655 51.295 111.465 ;
        RECT 51.495 111.085 52.565 111.255 ;
        RECT 51.495 110.730 51.815 111.085 ;
        RECT 48.150 109.925 48.500 110.575 ;
        RECT 49.190 110.095 49.600 110.645 ;
        RECT 51.490 110.475 51.815 110.730 ;
        RECT 49.785 110.265 51.815 110.475 ;
        RECT 51.470 110.255 51.815 110.265 ;
        RECT 51.985 110.515 52.225 110.915 ;
        RECT 52.395 110.855 52.565 111.085 ;
        RECT 52.735 111.025 52.925 111.465 ;
        RECT 53.095 111.015 54.045 111.295 ;
        RECT 54.265 111.105 54.615 111.275 ;
        RECT 52.395 110.685 52.925 110.855 ;
        RECT 47.750 109.585 48.500 109.755 ;
        RECT 47.745 108.915 48.075 109.415 ;
        RECT 48.245 109.085 48.500 109.585 ;
        RECT 48.675 108.915 48.965 110.080 ;
        RECT 49.190 109.925 50.915 110.095 ;
        RECT 49.445 108.915 49.615 109.755 ;
        RECT 49.825 109.085 50.075 109.925 ;
        RECT 50.285 108.915 50.455 109.755 ;
        RECT 50.625 109.085 50.915 109.925 ;
        RECT 51.125 108.915 51.295 109.975 ;
        RECT 51.470 109.635 51.640 110.255 ;
        RECT 51.985 110.145 52.525 110.515 ;
        RECT 52.705 110.405 52.925 110.685 ;
        RECT 53.095 110.235 53.265 111.015 ;
        RECT 52.860 110.065 53.265 110.235 ;
        RECT 53.435 110.225 53.785 110.845 ;
        RECT 52.860 109.975 53.030 110.065 ;
        RECT 53.955 110.055 54.165 110.845 ;
        RECT 51.810 109.805 53.030 109.975 ;
        RECT 53.490 109.895 54.165 110.055 ;
        RECT 51.470 109.465 52.270 109.635 ;
        RECT 51.590 108.915 51.920 109.295 ;
        RECT 52.100 109.175 52.270 109.465 ;
        RECT 52.860 109.425 53.030 109.805 ;
        RECT 53.200 109.885 54.165 109.895 ;
        RECT 54.355 110.715 54.615 111.105 ;
        RECT 54.825 111.005 55.155 111.465 ;
        RECT 56.030 111.075 56.885 111.245 ;
        RECT 57.090 111.075 57.585 111.245 ;
        RECT 57.755 111.105 58.085 111.465 ;
        RECT 54.355 110.025 54.525 110.715 ;
        RECT 54.695 110.365 54.865 110.545 ;
        RECT 55.035 110.535 55.825 110.785 ;
        RECT 56.030 110.365 56.200 111.075 ;
        RECT 56.370 110.565 56.725 110.785 ;
        RECT 54.695 110.195 56.385 110.365 ;
        RECT 53.200 109.595 53.660 109.885 ;
        RECT 54.355 109.855 55.855 110.025 ;
        RECT 54.355 109.715 54.525 109.855 ;
        RECT 53.965 109.545 54.525 109.715 ;
        RECT 52.440 108.915 52.690 109.375 ;
        RECT 52.860 109.085 53.730 109.425 ;
        RECT 53.965 109.085 54.135 109.545 ;
        RECT 54.970 109.515 56.045 109.685 ;
        RECT 54.305 108.915 54.675 109.375 ;
        RECT 54.970 109.175 55.140 109.515 ;
        RECT 55.310 108.915 55.640 109.345 ;
        RECT 55.875 109.175 56.045 109.515 ;
        RECT 56.215 109.415 56.385 110.195 ;
        RECT 56.555 109.975 56.725 110.565 ;
        RECT 56.895 110.165 57.245 110.785 ;
        RECT 56.555 109.585 57.020 109.975 ;
        RECT 57.415 109.715 57.585 111.075 ;
        RECT 57.755 109.885 58.215 110.935 ;
        RECT 57.190 109.545 57.585 109.715 ;
        RECT 57.190 109.415 57.360 109.545 ;
        RECT 56.215 109.085 56.895 109.415 ;
        RECT 57.110 109.085 57.360 109.415 ;
        RECT 57.530 108.915 57.780 109.375 ;
        RECT 57.950 109.100 58.275 109.885 ;
        RECT 58.445 109.085 58.615 111.205 ;
        RECT 58.785 111.085 59.115 111.465 ;
        RECT 59.285 110.915 59.540 111.205 ;
        RECT 60.025 110.995 60.195 111.465 ;
        RECT 58.790 110.745 59.540 110.915 ;
        RECT 60.365 110.815 60.695 111.295 ;
        RECT 60.865 110.995 61.035 111.465 ;
        RECT 61.205 110.815 61.535 111.295 ;
        RECT 58.790 109.755 59.020 110.745 ;
        RECT 59.770 110.645 61.535 110.815 ;
        RECT 61.705 110.655 61.875 111.465 ;
        RECT 62.075 111.085 63.145 111.255 ;
        RECT 62.075 110.730 62.395 111.085 ;
        RECT 59.190 109.925 59.540 110.575 ;
        RECT 59.770 110.095 60.180 110.645 ;
        RECT 62.070 110.475 62.395 110.730 ;
        RECT 60.365 110.265 62.395 110.475 ;
        RECT 62.050 110.255 62.395 110.265 ;
        RECT 62.565 110.515 62.805 110.915 ;
        RECT 62.975 110.855 63.145 111.085 ;
        RECT 63.315 111.025 63.505 111.465 ;
        RECT 63.675 111.015 64.625 111.295 ;
        RECT 64.845 111.105 65.195 111.275 ;
        RECT 62.975 110.685 63.505 110.855 ;
        RECT 59.770 109.925 61.495 110.095 ;
        RECT 58.790 109.585 59.540 109.755 ;
        RECT 58.785 108.915 59.115 109.415 ;
        RECT 59.285 109.085 59.540 109.585 ;
        RECT 60.025 108.915 60.195 109.755 ;
        RECT 60.405 109.085 60.655 109.925 ;
        RECT 60.865 108.915 61.035 109.755 ;
        RECT 61.205 109.085 61.495 109.925 ;
        RECT 61.705 108.915 61.875 109.975 ;
        RECT 62.050 109.635 62.220 110.255 ;
        RECT 62.565 110.145 63.105 110.515 ;
        RECT 63.285 110.405 63.505 110.685 ;
        RECT 63.675 110.235 63.845 111.015 ;
        RECT 63.440 110.065 63.845 110.235 ;
        RECT 64.015 110.225 64.365 110.845 ;
        RECT 63.440 109.975 63.610 110.065 ;
        RECT 64.535 110.055 64.745 110.845 ;
        RECT 62.390 109.805 63.610 109.975 ;
        RECT 64.070 109.895 64.745 110.055 ;
        RECT 62.050 109.465 62.850 109.635 ;
        RECT 62.170 108.915 62.500 109.295 ;
        RECT 62.680 109.175 62.850 109.465 ;
        RECT 63.440 109.425 63.610 109.805 ;
        RECT 63.780 109.885 64.745 109.895 ;
        RECT 64.935 110.715 65.195 111.105 ;
        RECT 65.405 111.005 65.735 111.465 ;
        RECT 66.610 111.075 67.465 111.245 ;
        RECT 67.670 111.075 68.165 111.245 ;
        RECT 68.335 111.105 68.665 111.465 ;
        RECT 64.935 110.025 65.105 110.715 ;
        RECT 65.275 110.365 65.445 110.545 ;
        RECT 65.615 110.535 66.405 110.785 ;
        RECT 66.610 110.365 66.780 111.075 ;
        RECT 66.950 110.565 67.305 110.785 ;
        RECT 65.275 110.195 66.965 110.365 ;
        RECT 63.780 109.595 64.240 109.885 ;
        RECT 64.935 109.855 66.435 110.025 ;
        RECT 64.935 109.715 65.105 109.855 ;
        RECT 64.545 109.545 65.105 109.715 ;
        RECT 63.020 108.915 63.270 109.375 ;
        RECT 63.440 109.085 64.310 109.425 ;
        RECT 64.545 109.085 64.715 109.545 ;
        RECT 65.550 109.515 66.625 109.685 ;
        RECT 64.885 108.915 65.255 109.375 ;
        RECT 65.550 109.175 65.720 109.515 ;
        RECT 65.890 108.915 66.220 109.345 ;
        RECT 66.455 109.175 66.625 109.515 ;
        RECT 66.795 109.415 66.965 110.195 ;
        RECT 67.135 109.975 67.305 110.565 ;
        RECT 67.475 110.165 67.825 110.785 ;
        RECT 67.135 109.585 67.600 109.975 ;
        RECT 67.995 109.715 68.165 111.075 ;
        RECT 68.335 109.885 68.795 110.935 ;
        RECT 67.770 109.545 68.165 109.715 ;
        RECT 67.770 109.415 67.940 109.545 ;
        RECT 66.795 109.085 67.475 109.415 ;
        RECT 67.690 109.085 67.940 109.415 ;
        RECT 68.110 108.915 68.360 109.375 ;
        RECT 68.530 109.100 68.855 109.885 ;
        RECT 69.025 109.085 69.195 111.205 ;
        RECT 69.365 111.085 69.695 111.465 ;
        RECT 69.865 110.915 70.120 111.205 ;
        RECT 69.370 110.745 70.120 110.915 ;
        RECT 70.845 110.915 71.015 111.295 ;
        RECT 71.195 111.085 71.525 111.465 ;
        RECT 70.845 110.745 71.510 110.915 ;
        RECT 71.705 110.790 71.965 111.295 ;
        RECT 69.370 109.755 69.600 110.745 ;
        RECT 69.770 109.925 70.120 110.575 ;
        RECT 70.775 110.195 71.105 110.565 ;
        RECT 71.340 110.490 71.510 110.745 ;
        RECT 71.340 110.160 71.625 110.490 ;
        RECT 71.340 110.015 71.510 110.160 ;
        RECT 70.845 109.845 71.510 110.015 ;
        RECT 71.795 109.990 71.965 110.790 ;
        RECT 72.225 110.915 72.395 111.295 ;
        RECT 72.575 111.085 72.905 111.465 ;
        RECT 72.225 110.745 72.890 110.915 ;
        RECT 73.085 110.790 73.345 111.295 ;
        RECT 72.155 110.195 72.485 110.565 ;
        RECT 72.720 110.490 72.890 110.745 ;
        RECT 72.720 110.160 73.005 110.490 ;
        RECT 72.720 110.015 72.890 110.160 ;
        RECT 69.370 109.585 70.120 109.755 ;
        RECT 69.365 108.915 69.695 109.415 ;
        RECT 69.865 109.085 70.120 109.585 ;
        RECT 70.845 109.085 71.015 109.845 ;
        RECT 71.195 108.915 71.525 109.675 ;
        RECT 71.695 109.085 71.965 109.990 ;
        RECT 72.225 109.845 72.890 110.015 ;
        RECT 73.175 109.990 73.345 110.790 ;
        RECT 74.435 110.740 74.725 111.465 ;
        RECT 75.205 110.995 75.375 111.465 ;
        RECT 75.545 110.815 75.875 111.295 ;
        RECT 76.045 110.995 76.215 111.465 ;
        RECT 76.385 110.815 76.715 111.295 ;
        RECT 74.950 110.645 76.715 110.815 ;
        RECT 76.885 110.655 77.055 111.465 ;
        RECT 77.255 111.085 78.325 111.255 ;
        RECT 77.255 110.730 77.575 111.085 ;
        RECT 74.950 110.095 75.360 110.645 ;
        RECT 77.250 110.475 77.575 110.730 ;
        RECT 75.545 110.265 77.575 110.475 ;
        RECT 77.230 110.255 77.575 110.265 ;
        RECT 77.745 110.515 77.985 110.915 ;
        RECT 78.155 110.855 78.325 111.085 ;
        RECT 78.495 111.025 78.685 111.465 ;
        RECT 78.855 111.015 79.805 111.295 ;
        RECT 80.025 111.105 80.375 111.275 ;
        RECT 78.155 110.685 78.685 110.855 ;
        RECT 72.225 109.085 72.395 109.845 ;
        RECT 72.575 108.915 72.905 109.675 ;
        RECT 73.075 109.085 73.345 109.990 ;
        RECT 74.435 108.915 74.725 110.080 ;
        RECT 74.950 109.925 76.675 110.095 ;
        RECT 75.205 108.915 75.375 109.755 ;
        RECT 75.585 109.085 75.835 109.925 ;
        RECT 76.045 108.915 76.215 109.755 ;
        RECT 76.385 109.085 76.675 109.925 ;
        RECT 76.885 108.915 77.055 109.975 ;
        RECT 77.230 109.635 77.400 110.255 ;
        RECT 77.745 110.145 78.285 110.515 ;
        RECT 78.465 110.405 78.685 110.685 ;
        RECT 78.855 110.235 79.025 111.015 ;
        RECT 78.620 110.065 79.025 110.235 ;
        RECT 79.195 110.225 79.545 110.845 ;
        RECT 78.620 109.975 78.790 110.065 ;
        RECT 79.715 110.055 79.925 110.845 ;
        RECT 77.570 109.805 78.790 109.975 ;
        RECT 79.250 109.895 79.925 110.055 ;
        RECT 77.230 109.465 78.030 109.635 ;
        RECT 77.350 108.915 77.680 109.295 ;
        RECT 77.860 109.175 78.030 109.465 ;
        RECT 78.620 109.425 78.790 109.805 ;
        RECT 78.960 109.885 79.925 109.895 ;
        RECT 80.115 110.715 80.375 111.105 ;
        RECT 80.585 111.005 80.915 111.465 ;
        RECT 81.790 111.075 82.645 111.245 ;
        RECT 82.850 111.075 83.345 111.245 ;
        RECT 83.515 111.105 83.845 111.465 ;
        RECT 80.115 110.025 80.285 110.715 ;
        RECT 80.455 110.365 80.625 110.545 ;
        RECT 80.795 110.535 81.585 110.785 ;
        RECT 81.790 110.365 81.960 111.075 ;
        RECT 82.130 110.565 82.485 110.785 ;
        RECT 80.455 110.195 82.145 110.365 ;
        RECT 78.960 109.595 79.420 109.885 ;
        RECT 80.115 109.855 81.615 110.025 ;
        RECT 80.115 109.715 80.285 109.855 ;
        RECT 79.725 109.545 80.285 109.715 ;
        RECT 78.200 108.915 78.450 109.375 ;
        RECT 78.620 109.085 79.490 109.425 ;
        RECT 79.725 109.085 79.895 109.545 ;
        RECT 80.730 109.515 81.805 109.685 ;
        RECT 80.065 108.915 80.435 109.375 ;
        RECT 80.730 109.175 80.900 109.515 ;
        RECT 81.070 108.915 81.400 109.345 ;
        RECT 81.635 109.175 81.805 109.515 ;
        RECT 81.975 109.415 82.145 110.195 ;
        RECT 82.315 109.975 82.485 110.565 ;
        RECT 82.655 110.165 83.005 110.785 ;
        RECT 82.315 109.585 82.780 109.975 ;
        RECT 83.175 109.715 83.345 111.075 ;
        RECT 83.515 109.885 83.975 110.935 ;
        RECT 82.950 109.545 83.345 109.715 ;
        RECT 82.950 109.415 83.120 109.545 ;
        RECT 81.975 109.085 82.655 109.415 ;
        RECT 82.870 109.085 83.120 109.415 ;
        RECT 83.290 108.915 83.540 109.375 ;
        RECT 83.710 109.100 84.035 109.885 ;
        RECT 84.205 109.085 84.375 111.205 ;
        RECT 84.545 111.085 84.875 111.465 ;
        RECT 85.045 110.915 85.300 111.205 ;
        RECT 85.785 110.995 85.955 111.465 ;
        RECT 84.550 110.745 85.300 110.915 ;
        RECT 86.125 110.815 86.455 111.295 ;
        RECT 86.625 110.995 86.795 111.465 ;
        RECT 86.965 110.815 87.295 111.295 ;
        RECT 84.550 109.755 84.780 110.745 ;
        RECT 85.530 110.645 87.295 110.815 ;
        RECT 87.465 110.655 87.635 111.465 ;
        RECT 87.835 111.085 88.905 111.255 ;
        RECT 87.835 110.730 88.155 111.085 ;
        RECT 84.950 109.925 85.300 110.575 ;
        RECT 85.530 110.095 85.940 110.645 ;
        RECT 87.830 110.475 88.155 110.730 ;
        RECT 86.125 110.265 88.155 110.475 ;
        RECT 87.810 110.255 88.155 110.265 ;
        RECT 88.325 110.515 88.565 110.915 ;
        RECT 88.735 110.855 88.905 111.085 ;
        RECT 89.075 111.025 89.265 111.465 ;
        RECT 89.435 111.015 90.385 111.295 ;
        RECT 90.605 111.105 90.955 111.275 ;
        RECT 88.735 110.685 89.265 110.855 ;
        RECT 85.530 109.925 87.255 110.095 ;
        RECT 84.550 109.585 85.300 109.755 ;
        RECT 84.545 108.915 84.875 109.415 ;
        RECT 85.045 109.085 85.300 109.585 ;
        RECT 85.785 108.915 85.955 109.755 ;
        RECT 86.165 109.085 86.415 109.925 ;
        RECT 86.625 108.915 86.795 109.755 ;
        RECT 86.965 109.085 87.255 109.925 ;
        RECT 87.465 108.915 87.635 109.975 ;
        RECT 87.810 109.635 87.980 110.255 ;
        RECT 88.325 110.145 88.865 110.515 ;
        RECT 89.045 110.405 89.265 110.685 ;
        RECT 89.435 110.235 89.605 111.015 ;
        RECT 89.200 110.065 89.605 110.235 ;
        RECT 89.775 110.225 90.125 110.845 ;
        RECT 89.200 109.975 89.370 110.065 ;
        RECT 90.295 110.055 90.505 110.845 ;
        RECT 88.150 109.805 89.370 109.975 ;
        RECT 89.830 109.895 90.505 110.055 ;
        RECT 87.810 109.465 88.610 109.635 ;
        RECT 87.930 108.915 88.260 109.295 ;
        RECT 88.440 109.175 88.610 109.465 ;
        RECT 89.200 109.425 89.370 109.805 ;
        RECT 89.540 109.885 90.505 109.895 ;
        RECT 90.695 110.715 90.955 111.105 ;
        RECT 91.165 111.005 91.495 111.465 ;
        RECT 92.370 111.075 93.225 111.245 ;
        RECT 93.430 111.075 93.925 111.245 ;
        RECT 94.095 111.105 94.425 111.465 ;
        RECT 90.695 110.025 90.865 110.715 ;
        RECT 91.035 110.365 91.205 110.545 ;
        RECT 91.375 110.535 92.165 110.785 ;
        RECT 92.370 110.365 92.540 111.075 ;
        RECT 92.710 110.565 93.065 110.785 ;
        RECT 91.035 110.195 92.725 110.365 ;
        RECT 89.540 109.595 90.000 109.885 ;
        RECT 90.695 109.855 92.195 110.025 ;
        RECT 90.695 109.715 90.865 109.855 ;
        RECT 90.305 109.545 90.865 109.715 ;
        RECT 88.780 108.915 89.030 109.375 ;
        RECT 89.200 109.085 90.070 109.425 ;
        RECT 90.305 109.085 90.475 109.545 ;
        RECT 91.310 109.515 92.385 109.685 ;
        RECT 90.645 108.915 91.015 109.375 ;
        RECT 91.310 109.175 91.480 109.515 ;
        RECT 91.650 108.915 91.980 109.345 ;
        RECT 92.215 109.175 92.385 109.515 ;
        RECT 92.555 109.415 92.725 110.195 ;
        RECT 92.895 109.975 93.065 110.565 ;
        RECT 93.235 110.165 93.585 110.785 ;
        RECT 92.895 109.585 93.360 109.975 ;
        RECT 93.755 109.715 93.925 111.075 ;
        RECT 94.095 109.885 94.555 110.935 ;
        RECT 93.530 109.545 93.925 109.715 ;
        RECT 93.530 109.415 93.700 109.545 ;
        RECT 92.555 109.085 93.235 109.415 ;
        RECT 93.450 109.085 93.700 109.415 ;
        RECT 93.870 108.915 94.120 109.375 ;
        RECT 94.290 109.100 94.615 109.885 ;
        RECT 94.785 109.085 94.955 111.205 ;
        RECT 95.125 111.085 95.455 111.465 ;
        RECT 95.625 110.915 95.880 111.205 ;
        RECT 95.130 110.745 95.880 110.915 ;
        RECT 95.130 109.755 95.360 110.745 ;
        RECT 96.115 110.645 96.325 111.465 ;
        RECT 96.495 110.665 96.825 111.295 ;
        RECT 95.530 109.925 95.880 110.575 ;
        RECT 96.495 110.065 96.745 110.665 ;
        RECT 96.995 110.645 97.225 111.465 ;
        RECT 97.495 110.645 97.705 111.465 ;
        RECT 97.875 110.665 98.205 111.295 ;
        RECT 96.915 110.225 97.245 110.475 ;
        RECT 97.875 110.065 98.125 110.665 ;
        RECT 98.375 110.645 98.605 111.465 ;
        RECT 98.855 110.645 99.085 111.465 ;
        RECT 99.255 110.665 99.585 111.295 ;
        RECT 98.295 110.225 98.625 110.475 ;
        RECT 98.835 110.225 99.165 110.475 ;
        RECT 99.335 110.065 99.585 110.665 ;
        RECT 99.755 110.645 99.965 111.465 ;
        RECT 100.195 110.740 100.485 111.465 ;
        RECT 100.965 110.995 101.135 111.465 ;
        RECT 101.305 110.815 101.635 111.295 ;
        RECT 101.805 110.995 101.975 111.465 ;
        RECT 102.145 110.815 102.475 111.295 ;
        RECT 100.710 110.645 102.475 110.815 ;
        RECT 102.645 110.655 102.815 111.465 ;
        RECT 103.015 111.085 104.085 111.255 ;
        RECT 103.015 110.730 103.335 111.085 ;
        RECT 100.710 110.095 101.120 110.645 ;
        RECT 103.010 110.475 103.335 110.730 ;
        RECT 101.305 110.265 103.335 110.475 ;
        RECT 102.990 110.255 103.335 110.265 ;
        RECT 103.505 110.515 103.745 110.915 ;
        RECT 103.915 110.855 104.085 111.085 ;
        RECT 104.255 111.025 104.445 111.465 ;
        RECT 104.615 111.015 105.565 111.295 ;
        RECT 105.785 111.105 106.135 111.275 ;
        RECT 103.915 110.685 104.445 110.855 ;
        RECT 95.130 109.585 95.880 109.755 ;
        RECT 95.125 108.915 95.455 109.415 ;
        RECT 95.625 109.085 95.880 109.585 ;
        RECT 96.115 108.915 96.325 110.055 ;
        RECT 96.495 109.085 96.825 110.065 ;
        RECT 96.995 108.915 97.225 110.055 ;
        RECT 97.495 108.915 97.705 110.055 ;
        RECT 97.875 109.085 98.205 110.065 ;
        RECT 98.375 108.915 98.605 110.055 ;
        RECT 98.855 108.915 99.085 110.055 ;
        RECT 99.255 109.085 99.585 110.065 ;
        RECT 99.755 108.915 99.965 110.055 ;
        RECT 100.195 108.915 100.485 110.080 ;
        RECT 100.710 109.925 102.435 110.095 ;
        RECT 100.965 108.915 101.135 109.755 ;
        RECT 101.345 109.085 101.595 109.925 ;
        RECT 101.805 108.915 101.975 109.755 ;
        RECT 102.145 109.085 102.435 109.925 ;
        RECT 102.645 108.915 102.815 109.975 ;
        RECT 102.990 109.635 103.160 110.255 ;
        RECT 103.505 110.145 104.045 110.515 ;
        RECT 104.225 110.405 104.445 110.685 ;
        RECT 104.615 110.235 104.785 111.015 ;
        RECT 104.380 110.065 104.785 110.235 ;
        RECT 104.955 110.225 105.305 110.845 ;
        RECT 104.380 109.975 104.550 110.065 ;
        RECT 105.475 110.055 105.685 110.845 ;
        RECT 103.330 109.805 104.550 109.975 ;
        RECT 105.010 109.895 105.685 110.055 ;
        RECT 102.990 109.465 103.790 109.635 ;
        RECT 103.110 108.915 103.440 109.295 ;
        RECT 103.620 109.175 103.790 109.465 ;
        RECT 104.380 109.425 104.550 109.805 ;
        RECT 104.720 109.885 105.685 109.895 ;
        RECT 105.875 110.715 106.135 111.105 ;
        RECT 106.345 111.005 106.675 111.465 ;
        RECT 107.550 111.075 108.405 111.245 ;
        RECT 108.610 111.075 109.105 111.245 ;
        RECT 109.275 111.105 109.605 111.465 ;
        RECT 105.875 110.025 106.045 110.715 ;
        RECT 106.215 110.365 106.385 110.545 ;
        RECT 106.555 110.535 107.345 110.785 ;
        RECT 107.550 110.365 107.720 111.075 ;
        RECT 107.890 110.565 108.245 110.785 ;
        RECT 106.215 110.195 107.905 110.365 ;
        RECT 104.720 109.595 105.180 109.885 ;
        RECT 105.875 109.855 107.375 110.025 ;
        RECT 105.875 109.715 106.045 109.855 ;
        RECT 105.485 109.545 106.045 109.715 ;
        RECT 103.960 108.915 104.210 109.375 ;
        RECT 104.380 109.085 105.250 109.425 ;
        RECT 105.485 109.085 105.655 109.545 ;
        RECT 106.490 109.515 107.565 109.685 ;
        RECT 105.825 108.915 106.195 109.375 ;
        RECT 106.490 109.175 106.660 109.515 ;
        RECT 106.830 108.915 107.160 109.345 ;
        RECT 107.395 109.175 107.565 109.515 ;
        RECT 107.735 109.415 107.905 110.195 ;
        RECT 108.075 109.975 108.245 110.565 ;
        RECT 108.415 110.165 108.765 110.785 ;
        RECT 108.075 109.585 108.540 109.975 ;
        RECT 108.935 109.715 109.105 111.075 ;
        RECT 109.275 109.885 109.735 110.935 ;
        RECT 108.710 109.545 109.105 109.715 ;
        RECT 108.710 109.415 108.880 109.545 ;
        RECT 107.735 109.085 108.415 109.415 ;
        RECT 108.630 109.085 108.880 109.415 ;
        RECT 109.050 108.915 109.300 109.375 ;
        RECT 109.470 109.100 109.795 109.885 ;
        RECT 109.965 109.085 110.135 111.205 ;
        RECT 110.305 111.085 110.635 111.465 ;
        RECT 110.805 110.915 111.060 111.205 ;
        RECT 110.310 110.745 111.060 110.915 ;
        RECT 110.310 109.755 110.540 110.745 ;
        RECT 112.155 110.715 113.365 111.465 ;
        RECT 110.710 109.925 111.060 110.575 ;
        RECT 112.155 110.005 112.675 110.545 ;
        RECT 112.845 110.175 113.365 110.715 ;
        RECT 110.310 109.585 111.060 109.755 ;
        RECT 110.305 108.915 110.635 109.415 ;
        RECT 110.805 109.085 111.060 109.585 ;
        RECT 112.155 108.915 113.365 110.005 ;
        RECT 15.010 108.745 113.450 108.915 ;
        RECT 15.095 107.655 16.305 108.745 ;
        RECT 17.400 108.310 22.745 108.745 ;
        RECT 15.095 106.945 15.615 107.485 ;
        RECT 15.785 107.115 16.305 107.655 ;
        RECT 18.990 107.060 19.340 108.310 ;
        RECT 22.915 107.580 23.205 108.745 ;
        RECT 23.685 107.905 23.855 108.745 ;
        RECT 24.065 107.735 24.315 108.575 ;
        RECT 24.525 107.905 24.695 108.745 ;
        RECT 24.865 107.735 25.155 108.575 ;
        RECT 15.095 106.195 16.305 106.945 ;
        RECT 20.820 106.740 21.160 107.570 ;
        RECT 23.430 107.565 25.155 107.735 ;
        RECT 25.365 107.685 25.535 108.745 ;
        RECT 25.830 108.365 26.160 108.745 ;
        RECT 26.340 108.195 26.510 108.485 ;
        RECT 26.680 108.285 26.930 108.745 ;
        RECT 25.710 108.025 26.510 108.195 ;
        RECT 27.100 108.235 27.970 108.575 ;
        RECT 23.430 107.015 23.840 107.565 ;
        RECT 25.710 107.405 25.880 108.025 ;
        RECT 27.100 107.855 27.270 108.235 ;
        RECT 28.205 108.115 28.375 108.575 ;
        RECT 28.545 108.285 28.915 108.745 ;
        RECT 29.210 108.145 29.380 108.485 ;
        RECT 29.550 108.315 29.880 108.745 ;
        RECT 30.115 108.145 30.285 108.485 ;
        RECT 26.050 107.685 27.270 107.855 ;
        RECT 27.440 107.775 27.900 108.065 ;
        RECT 28.205 107.945 28.765 108.115 ;
        RECT 29.210 107.975 30.285 108.145 ;
        RECT 30.455 108.245 31.135 108.575 ;
        RECT 31.350 108.245 31.600 108.575 ;
        RECT 31.770 108.285 32.020 108.745 ;
        RECT 28.595 107.805 28.765 107.945 ;
        RECT 27.440 107.765 28.405 107.775 ;
        RECT 27.100 107.595 27.270 107.685 ;
        RECT 27.730 107.605 28.405 107.765 ;
        RECT 25.710 107.395 26.055 107.405 ;
        RECT 24.025 107.185 26.055 107.395 ;
        RECT 17.400 106.195 22.745 106.740 ;
        RECT 22.915 106.195 23.205 106.920 ;
        RECT 23.430 106.845 25.195 107.015 ;
        RECT 23.685 106.195 23.855 106.665 ;
        RECT 24.025 106.365 24.355 106.845 ;
        RECT 24.525 106.195 24.695 106.665 ;
        RECT 24.865 106.365 25.195 106.845 ;
        RECT 25.365 106.195 25.535 107.005 ;
        RECT 25.730 106.930 26.055 107.185 ;
        RECT 25.735 106.575 26.055 106.930 ;
        RECT 26.225 107.145 26.765 107.515 ;
        RECT 27.100 107.425 27.505 107.595 ;
        RECT 26.225 106.745 26.465 107.145 ;
        RECT 26.945 106.975 27.165 107.255 ;
        RECT 26.635 106.805 27.165 106.975 ;
        RECT 26.635 106.575 26.805 106.805 ;
        RECT 27.335 106.645 27.505 107.425 ;
        RECT 27.675 106.815 28.025 107.435 ;
        RECT 28.195 106.815 28.405 107.605 ;
        RECT 28.595 107.635 30.095 107.805 ;
        RECT 28.595 106.945 28.765 107.635 ;
        RECT 30.455 107.465 30.625 108.245 ;
        RECT 31.430 108.115 31.600 108.245 ;
        RECT 28.935 107.295 30.625 107.465 ;
        RECT 30.795 107.685 31.260 108.075 ;
        RECT 31.430 107.945 31.825 108.115 ;
        RECT 28.935 107.115 29.105 107.295 ;
        RECT 25.735 106.405 26.805 106.575 ;
        RECT 26.975 106.195 27.165 106.635 ;
        RECT 27.335 106.365 28.285 106.645 ;
        RECT 28.595 106.555 28.855 106.945 ;
        RECT 29.275 106.875 30.065 107.125 ;
        RECT 28.505 106.385 28.855 106.555 ;
        RECT 29.065 106.195 29.395 106.655 ;
        RECT 30.270 106.585 30.440 107.295 ;
        RECT 30.795 107.095 30.965 107.685 ;
        RECT 30.610 106.875 30.965 107.095 ;
        RECT 31.135 106.875 31.485 107.495 ;
        RECT 31.655 106.585 31.825 107.945 ;
        RECT 32.190 107.775 32.515 108.560 ;
        RECT 31.995 106.725 32.455 107.775 ;
        RECT 30.270 106.415 31.125 106.585 ;
        RECT 31.330 106.415 31.825 106.585 ;
        RECT 31.995 106.195 32.325 106.555 ;
        RECT 32.685 106.455 32.855 108.575 ;
        RECT 33.025 108.245 33.355 108.745 ;
        RECT 33.525 108.075 33.780 108.575 ;
        RECT 33.030 107.905 33.780 108.075 ;
        RECT 33.030 106.915 33.260 107.905 ;
        RECT 33.430 107.085 33.780 107.735 ;
        RECT 33.955 107.655 35.625 108.745 ;
        RECT 33.955 107.135 34.705 107.655 ;
        RECT 35.795 107.580 36.085 108.745 ;
        RECT 36.720 108.310 42.065 108.745 ;
        RECT 34.875 106.965 35.625 107.485 ;
        RECT 38.310 107.060 38.660 108.310 ;
        RECT 42.295 107.605 42.505 108.745 ;
        RECT 42.675 107.595 43.005 108.575 ;
        RECT 43.175 107.605 43.405 108.745 ;
        RECT 43.615 107.655 47.125 108.745 ;
        RECT 33.030 106.745 33.780 106.915 ;
        RECT 33.025 106.195 33.355 106.575 ;
        RECT 33.525 106.455 33.780 106.745 ;
        RECT 33.955 106.195 35.625 106.965 ;
        RECT 35.795 106.195 36.085 106.920 ;
        RECT 40.140 106.740 40.480 107.570 ;
        RECT 36.720 106.195 42.065 106.740 ;
        RECT 42.295 106.195 42.505 107.015 ;
        RECT 42.675 106.995 42.925 107.595 ;
        RECT 43.095 107.185 43.425 107.435 ;
        RECT 43.615 107.135 45.305 107.655 ;
        RECT 47.335 107.605 47.565 108.745 ;
        RECT 47.735 107.595 48.065 108.575 ;
        RECT 48.235 107.605 48.445 108.745 ;
        RECT 42.675 106.365 43.005 106.995 ;
        RECT 43.175 106.195 43.405 107.015 ;
        RECT 45.475 106.965 47.125 107.485 ;
        RECT 47.315 107.185 47.645 107.435 ;
        RECT 43.615 106.195 47.125 106.965 ;
        RECT 47.335 106.195 47.565 107.015 ;
        RECT 47.815 106.995 48.065 107.595 ;
        RECT 48.675 107.580 48.965 108.745 ;
        RECT 49.635 107.605 49.865 108.745 ;
        RECT 50.035 107.595 50.365 108.575 ;
        RECT 50.535 107.605 50.745 108.745 ;
        RECT 51.285 107.905 51.455 108.745 ;
        RECT 51.665 107.735 51.915 108.575 ;
        RECT 52.125 107.905 52.295 108.745 ;
        RECT 52.465 107.735 52.755 108.575 ;
        RECT 49.615 107.185 49.945 107.435 ;
        RECT 47.735 106.365 48.065 106.995 ;
        RECT 48.235 106.195 48.445 107.015 ;
        RECT 48.675 106.195 48.965 106.920 ;
        RECT 49.635 106.195 49.865 107.015 ;
        RECT 50.115 106.995 50.365 107.595 ;
        RECT 51.030 107.565 52.755 107.735 ;
        RECT 52.965 107.685 53.135 108.745 ;
        RECT 53.430 108.365 53.760 108.745 ;
        RECT 53.940 108.195 54.110 108.485 ;
        RECT 54.280 108.285 54.530 108.745 ;
        RECT 53.310 108.025 54.110 108.195 ;
        RECT 54.700 108.235 55.570 108.575 ;
        RECT 51.030 107.015 51.440 107.565 ;
        RECT 53.310 107.405 53.480 108.025 ;
        RECT 54.700 107.855 54.870 108.235 ;
        RECT 55.805 108.115 55.975 108.575 ;
        RECT 56.145 108.285 56.515 108.745 ;
        RECT 56.810 108.145 56.980 108.485 ;
        RECT 57.150 108.315 57.480 108.745 ;
        RECT 57.715 108.145 57.885 108.485 ;
        RECT 53.650 107.685 54.870 107.855 ;
        RECT 55.040 107.775 55.500 108.065 ;
        RECT 55.805 107.945 56.365 108.115 ;
        RECT 56.810 107.975 57.885 108.145 ;
        RECT 58.055 108.245 58.735 108.575 ;
        RECT 58.950 108.245 59.200 108.575 ;
        RECT 59.370 108.285 59.620 108.745 ;
        RECT 56.195 107.805 56.365 107.945 ;
        RECT 55.040 107.765 56.005 107.775 ;
        RECT 54.700 107.595 54.870 107.685 ;
        RECT 55.330 107.605 56.005 107.765 ;
        RECT 53.310 107.395 53.655 107.405 ;
        RECT 51.625 107.185 53.655 107.395 ;
        RECT 50.035 106.365 50.365 106.995 ;
        RECT 50.535 106.195 50.745 107.015 ;
        RECT 51.030 106.845 52.795 107.015 ;
        RECT 51.285 106.195 51.455 106.665 ;
        RECT 51.625 106.365 51.955 106.845 ;
        RECT 52.125 106.195 52.295 106.665 ;
        RECT 52.465 106.365 52.795 106.845 ;
        RECT 52.965 106.195 53.135 107.005 ;
        RECT 53.330 106.930 53.655 107.185 ;
        RECT 53.335 106.575 53.655 106.930 ;
        RECT 53.825 107.145 54.365 107.515 ;
        RECT 54.700 107.425 55.105 107.595 ;
        RECT 53.825 106.745 54.065 107.145 ;
        RECT 54.545 106.975 54.765 107.255 ;
        RECT 54.235 106.805 54.765 106.975 ;
        RECT 54.235 106.575 54.405 106.805 ;
        RECT 54.935 106.645 55.105 107.425 ;
        RECT 55.275 106.815 55.625 107.435 ;
        RECT 55.795 106.815 56.005 107.605 ;
        RECT 56.195 107.635 57.695 107.805 ;
        RECT 56.195 106.945 56.365 107.635 ;
        RECT 58.055 107.465 58.225 108.245 ;
        RECT 59.030 108.115 59.200 108.245 ;
        RECT 56.535 107.295 58.225 107.465 ;
        RECT 58.395 107.685 58.860 108.075 ;
        RECT 59.030 107.945 59.425 108.115 ;
        RECT 56.535 107.115 56.705 107.295 ;
        RECT 53.335 106.405 54.405 106.575 ;
        RECT 54.575 106.195 54.765 106.635 ;
        RECT 54.935 106.365 55.885 106.645 ;
        RECT 56.195 106.555 56.455 106.945 ;
        RECT 56.875 106.875 57.665 107.125 ;
        RECT 56.105 106.385 56.455 106.555 ;
        RECT 56.665 106.195 56.995 106.655 ;
        RECT 57.870 106.585 58.040 107.295 ;
        RECT 58.395 107.095 58.565 107.685 ;
        RECT 58.210 106.875 58.565 107.095 ;
        RECT 58.735 106.875 59.085 107.495 ;
        RECT 59.255 106.585 59.425 107.945 ;
        RECT 59.790 107.775 60.115 108.560 ;
        RECT 59.595 106.725 60.055 107.775 ;
        RECT 57.870 106.415 58.725 106.585 ;
        RECT 58.930 106.415 59.425 106.585 ;
        RECT 59.595 106.195 59.925 106.555 ;
        RECT 60.285 106.455 60.455 108.575 ;
        RECT 60.625 108.245 60.955 108.745 ;
        RECT 61.125 108.075 61.380 108.575 ;
        RECT 60.630 107.905 61.380 108.075 ;
        RECT 60.630 106.915 60.860 107.905 ;
        RECT 61.030 107.085 61.380 107.735 ;
        RECT 61.555 107.580 61.845 108.745 ;
        RECT 62.475 107.655 65.065 108.745 ;
        RECT 65.240 108.310 70.585 108.745 ;
        RECT 62.475 107.135 63.685 107.655 ;
        RECT 63.855 106.965 65.065 107.485 ;
        RECT 66.830 107.060 67.180 108.310 ;
        RECT 70.815 107.605 71.025 108.745 ;
        RECT 71.195 107.595 71.525 108.575 ;
        RECT 71.695 107.605 71.925 108.745 ;
        RECT 72.635 107.605 72.865 108.745 ;
        RECT 73.035 107.595 73.365 108.575 ;
        RECT 73.535 107.605 73.745 108.745 ;
        RECT 60.630 106.745 61.380 106.915 ;
        RECT 60.625 106.195 60.955 106.575 ;
        RECT 61.125 106.455 61.380 106.745 ;
        RECT 61.555 106.195 61.845 106.920 ;
        RECT 62.475 106.195 65.065 106.965 ;
        RECT 68.660 106.740 69.000 107.570 ;
        RECT 65.240 106.195 70.585 106.740 ;
        RECT 70.815 106.195 71.025 107.015 ;
        RECT 71.195 106.995 71.445 107.595 ;
        RECT 71.615 107.185 71.945 107.435 ;
        RECT 72.615 107.185 72.945 107.435 ;
        RECT 71.195 106.365 71.525 106.995 ;
        RECT 71.695 106.195 71.925 107.015 ;
        RECT 72.635 106.195 72.865 107.015 ;
        RECT 73.115 106.995 73.365 107.595 ;
        RECT 74.435 107.580 74.725 108.745 ;
        RECT 75.395 107.605 75.625 108.745 ;
        RECT 75.795 107.595 76.125 108.575 ;
        RECT 76.295 107.605 76.505 108.745 ;
        RECT 77.045 107.905 77.215 108.745 ;
        RECT 77.425 107.735 77.675 108.575 ;
        RECT 77.885 107.905 78.055 108.745 ;
        RECT 78.225 107.735 78.515 108.575 ;
        RECT 75.375 107.185 75.705 107.435 ;
        RECT 73.035 106.365 73.365 106.995 ;
        RECT 73.535 106.195 73.745 107.015 ;
        RECT 74.435 106.195 74.725 106.920 ;
        RECT 75.395 106.195 75.625 107.015 ;
        RECT 75.875 106.995 76.125 107.595 ;
        RECT 76.790 107.565 78.515 107.735 ;
        RECT 78.725 107.685 78.895 108.745 ;
        RECT 79.190 108.365 79.520 108.745 ;
        RECT 79.700 108.195 79.870 108.485 ;
        RECT 80.040 108.285 80.290 108.745 ;
        RECT 79.070 108.025 79.870 108.195 ;
        RECT 80.460 108.235 81.330 108.575 ;
        RECT 76.790 107.015 77.200 107.565 ;
        RECT 79.070 107.405 79.240 108.025 ;
        RECT 80.460 107.855 80.630 108.235 ;
        RECT 81.565 108.115 81.735 108.575 ;
        RECT 81.905 108.285 82.275 108.745 ;
        RECT 82.570 108.145 82.740 108.485 ;
        RECT 82.910 108.315 83.240 108.745 ;
        RECT 83.475 108.145 83.645 108.485 ;
        RECT 79.410 107.685 80.630 107.855 ;
        RECT 80.800 107.775 81.260 108.065 ;
        RECT 81.565 107.945 82.125 108.115 ;
        RECT 82.570 107.975 83.645 108.145 ;
        RECT 83.815 108.245 84.495 108.575 ;
        RECT 84.710 108.245 84.960 108.575 ;
        RECT 85.130 108.285 85.380 108.745 ;
        RECT 81.955 107.805 82.125 107.945 ;
        RECT 80.800 107.765 81.765 107.775 ;
        RECT 80.460 107.595 80.630 107.685 ;
        RECT 81.090 107.605 81.765 107.765 ;
        RECT 79.070 107.395 79.415 107.405 ;
        RECT 77.385 107.185 79.415 107.395 ;
        RECT 75.795 106.365 76.125 106.995 ;
        RECT 76.295 106.195 76.505 107.015 ;
        RECT 76.790 106.845 78.555 107.015 ;
        RECT 77.045 106.195 77.215 106.665 ;
        RECT 77.385 106.365 77.715 106.845 ;
        RECT 77.885 106.195 78.055 106.665 ;
        RECT 78.225 106.365 78.555 106.845 ;
        RECT 78.725 106.195 78.895 107.005 ;
        RECT 79.090 106.930 79.415 107.185 ;
        RECT 79.095 106.575 79.415 106.930 ;
        RECT 79.585 107.145 80.125 107.515 ;
        RECT 80.460 107.425 80.865 107.595 ;
        RECT 79.585 106.745 79.825 107.145 ;
        RECT 80.305 106.975 80.525 107.255 ;
        RECT 79.995 106.805 80.525 106.975 ;
        RECT 79.995 106.575 80.165 106.805 ;
        RECT 80.695 106.645 80.865 107.425 ;
        RECT 81.035 106.815 81.385 107.435 ;
        RECT 81.555 106.815 81.765 107.605 ;
        RECT 81.955 107.635 83.455 107.805 ;
        RECT 81.955 106.945 82.125 107.635 ;
        RECT 83.815 107.465 83.985 108.245 ;
        RECT 84.790 108.115 84.960 108.245 ;
        RECT 82.295 107.295 83.985 107.465 ;
        RECT 84.155 107.685 84.620 108.075 ;
        RECT 84.790 107.945 85.185 108.115 ;
        RECT 82.295 107.115 82.465 107.295 ;
        RECT 79.095 106.405 80.165 106.575 ;
        RECT 80.335 106.195 80.525 106.635 ;
        RECT 80.695 106.365 81.645 106.645 ;
        RECT 81.955 106.555 82.215 106.945 ;
        RECT 82.635 106.875 83.425 107.125 ;
        RECT 81.865 106.385 82.215 106.555 ;
        RECT 82.425 106.195 82.755 106.655 ;
        RECT 83.630 106.585 83.800 107.295 ;
        RECT 84.155 107.095 84.325 107.685 ;
        RECT 83.970 106.875 84.325 107.095 ;
        RECT 84.495 106.875 84.845 107.495 ;
        RECT 85.015 106.585 85.185 107.945 ;
        RECT 85.550 107.775 85.875 108.560 ;
        RECT 85.355 106.725 85.815 107.775 ;
        RECT 83.630 106.415 84.485 106.585 ;
        RECT 84.690 106.415 85.185 106.585 ;
        RECT 85.355 106.195 85.685 106.555 ;
        RECT 86.045 106.455 86.215 108.575 ;
        RECT 86.385 108.245 86.715 108.745 ;
        RECT 86.885 108.075 87.140 108.575 ;
        RECT 86.390 107.905 87.140 108.075 ;
        RECT 86.390 106.915 86.620 107.905 ;
        RECT 86.790 107.085 87.140 107.735 ;
        RECT 87.315 107.580 87.605 108.745 ;
        RECT 88.275 107.605 88.505 108.745 ;
        RECT 88.675 107.595 89.005 108.575 ;
        RECT 89.175 107.605 89.385 108.745 ;
        RECT 89.925 107.905 90.095 108.745 ;
        RECT 90.305 107.735 90.555 108.575 ;
        RECT 90.765 107.905 90.935 108.745 ;
        RECT 91.105 107.735 91.395 108.575 ;
        RECT 88.255 107.185 88.585 107.435 ;
        RECT 86.390 106.745 87.140 106.915 ;
        RECT 86.385 106.195 86.715 106.575 ;
        RECT 86.885 106.455 87.140 106.745 ;
        RECT 87.315 106.195 87.605 106.920 ;
        RECT 88.275 106.195 88.505 107.015 ;
        RECT 88.755 106.995 89.005 107.595 ;
        RECT 89.670 107.565 91.395 107.735 ;
        RECT 91.605 107.685 91.775 108.745 ;
        RECT 92.070 108.365 92.400 108.745 ;
        RECT 92.580 108.195 92.750 108.485 ;
        RECT 92.920 108.285 93.170 108.745 ;
        RECT 91.950 108.025 92.750 108.195 ;
        RECT 93.340 108.235 94.210 108.575 ;
        RECT 89.670 107.015 90.080 107.565 ;
        RECT 91.950 107.405 92.120 108.025 ;
        RECT 93.340 107.855 93.510 108.235 ;
        RECT 94.445 108.115 94.615 108.575 ;
        RECT 94.785 108.285 95.155 108.745 ;
        RECT 95.450 108.145 95.620 108.485 ;
        RECT 95.790 108.315 96.120 108.745 ;
        RECT 96.355 108.145 96.525 108.485 ;
        RECT 92.290 107.685 93.510 107.855 ;
        RECT 93.680 107.775 94.140 108.065 ;
        RECT 94.445 107.945 95.005 108.115 ;
        RECT 95.450 107.975 96.525 108.145 ;
        RECT 96.695 108.245 97.375 108.575 ;
        RECT 97.590 108.245 97.840 108.575 ;
        RECT 98.010 108.285 98.260 108.745 ;
        RECT 94.835 107.805 95.005 107.945 ;
        RECT 93.680 107.765 94.645 107.775 ;
        RECT 93.340 107.595 93.510 107.685 ;
        RECT 93.970 107.605 94.645 107.765 ;
        RECT 91.950 107.395 92.295 107.405 ;
        RECT 90.265 107.185 92.295 107.395 ;
        RECT 88.675 106.365 89.005 106.995 ;
        RECT 89.175 106.195 89.385 107.015 ;
        RECT 89.670 106.845 91.435 107.015 ;
        RECT 89.925 106.195 90.095 106.665 ;
        RECT 90.265 106.365 90.595 106.845 ;
        RECT 90.765 106.195 90.935 106.665 ;
        RECT 91.105 106.365 91.435 106.845 ;
        RECT 91.605 106.195 91.775 107.005 ;
        RECT 91.970 106.930 92.295 107.185 ;
        RECT 91.975 106.575 92.295 106.930 ;
        RECT 92.465 107.145 93.005 107.515 ;
        RECT 93.340 107.425 93.745 107.595 ;
        RECT 92.465 106.745 92.705 107.145 ;
        RECT 93.185 106.975 93.405 107.255 ;
        RECT 92.875 106.805 93.405 106.975 ;
        RECT 92.875 106.575 93.045 106.805 ;
        RECT 93.575 106.645 93.745 107.425 ;
        RECT 93.915 106.815 94.265 107.435 ;
        RECT 94.435 106.815 94.645 107.605 ;
        RECT 94.835 107.635 96.335 107.805 ;
        RECT 94.835 106.945 95.005 107.635 ;
        RECT 96.695 107.465 96.865 108.245 ;
        RECT 97.670 108.115 97.840 108.245 ;
        RECT 95.175 107.295 96.865 107.465 ;
        RECT 97.035 107.685 97.500 108.075 ;
        RECT 97.670 107.945 98.065 108.115 ;
        RECT 95.175 107.115 95.345 107.295 ;
        RECT 91.975 106.405 93.045 106.575 ;
        RECT 93.215 106.195 93.405 106.635 ;
        RECT 93.575 106.365 94.525 106.645 ;
        RECT 94.835 106.555 95.095 106.945 ;
        RECT 95.515 106.875 96.305 107.125 ;
        RECT 94.745 106.385 95.095 106.555 ;
        RECT 95.305 106.195 95.635 106.655 ;
        RECT 96.510 106.585 96.680 107.295 ;
        RECT 97.035 107.095 97.205 107.685 ;
        RECT 96.850 106.875 97.205 107.095 ;
        RECT 97.375 106.875 97.725 107.495 ;
        RECT 97.895 106.585 98.065 107.945 ;
        RECT 98.430 107.775 98.755 108.560 ;
        RECT 98.235 106.725 98.695 107.775 ;
        RECT 96.510 106.415 97.365 106.585 ;
        RECT 97.570 106.415 98.065 106.585 ;
        RECT 98.235 106.195 98.565 106.555 ;
        RECT 98.925 106.455 99.095 108.575 ;
        RECT 99.265 108.245 99.595 108.745 ;
        RECT 99.765 108.075 100.020 108.575 ;
        RECT 99.270 107.905 100.020 108.075 ;
        RECT 99.270 106.915 99.500 107.905 ;
        RECT 99.670 107.085 100.020 107.735 ;
        RECT 100.195 107.580 100.485 108.745 ;
        RECT 100.655 107.655 101.865 108.745 ;
        RECT 102.035 107.655 105.545 108.745 ;
        RECT 100.655 107.115 101.175 107.655 ;
        RECT 101.345 106.945 101.865 107.485 ;
        RECT 102.035 107.135 103.725 107.655 ;
        RECT 105.775 107.605 105.985 108.745 ;
        RECT 106.155 107.595 106.485 108.575 ;
        RECT 106.655 107.605 106.885 108.745 ;
        RECT 107.095 107.655 110.605 108.745 ;
        RECT 110.775 107.670 111.045 108.575 ;
        RECT 111.215 107.985 111.545 108.745 ;
        RECT 111.725 107.815 111.905 108.575 ;
        RECT 103.895 106.965 105.545 107.485 ;
        RECT 99.270 106.745 100.020 106.915 ;
        RECT 99.265 106.195 99.595 106.575 ;
        RECT 99.765 106.455 100.020 106.745 ;
        RECT 100.195 106.195 100.485 106.920 ;
        RECT 100.655 106.195 101.865 106.945 ;
        RECT 102.035 106.195 105.545 106.965 ;
        RECT 105.775 106.195 105.985 107.015 ;
        RECT 106.155 106.995 106.405 107.595 ;
        RECT 106.575 107.185 106.905 107.435 ;
        RECT 107.095 107.135 108.785 107.655 ;
        RECT 106.155 106.365 106.485 106.995 ;
        RECT 106.655 106.195 106.885 107.015 ;
        RECT 108.955 106.965 110.605 107.485 ;
        RECT 107.095 106.195 110.605 106.965 ;
        RECT 110.775 106.870 110.955 107.670 ;
        RECT 111.230 107.645 111.905 107.815 ;
        RECT 112.155 107.655 113.365 108.745 ;
        RECT 111.230 107.500 111.400 107.645 ;
        RECT 111.125 107.170 111.400 107.500 ;
        RECT 111.230 106.915 111.400 107.170 ;
        RECT 111.625 107.095 111.965 107.465 ;
        RECT 112.155 107.115 112.675 107.655 ;
        RECT 112.845 106.945 113.365 107.485 ;
        RECT 110.775 106.365 111.035 106.870 ;
        RECT 111.230 106.745 111.895 106.915 ;
        RECT 111.215 106.195 111.545 106.575 ;
        RECT 111.725 106.365 111.895 106.745 ;
        RECT 112.155 106.195 113.365 106.945 ;
        RECT 15.010 106.025 113.450 106.195 ;
        RECT 19.165 66.070 30.165 66.940 ;
        RECT 19.165 54.930 20.835 66.070 ;
        RECT 21.465 65.555 26.465 65.725 ;
        RECT 21.235 55.300 21.405 65.340 ;
        RECT 26.525 55.300 26.695 65.340 ;
        RECT 27.095 54.930 27.265 66.070 ;
        RECT 27.895 65.555 28.895 65.725 ;
        RECT 27.665 55.300 27.835 65.340 ;
        RECT 28.955 55.300 29.125 65.340 ;
        RECT 29.525 54.930 30.165 66.070 ;
        RECT 19.165 52.860 30.165 54.930 ;
        RECT 19.165 49.370 21.005 52.860 ;
        RECT 22.765 52.780 30.165 52.860 ;
        RECT 21.635 52.350 22.135 52.520 ;
        RECT 21.405 50.095 21.575 52.135 ;
        RECT 22.195 50.095 22.365 52.135 ;
        RECT 21.635 49.710 22.135 49.880 ;
        RECT 22.765 49.370 25.085 52.780 ;
        RECT 25.715 52.270 26.215 52.440 ;
        RECT 19.165 48.650 25.085 49.370 ;
        RECT 19.135 48.040 23.045 48.260 ;
        RECT 19.135 45.640 20.855 48.040 ;
        RECT 21.485 47.530 21.985 47.700 ;
        RECT 21.255 46.320 21.425 47.360 ;
        RECT 22.045 46.320 22.215 47.360 ;
        RECT 21.485 45.980 21.985 46.150 ;
        RECT 22.615 45.640 23.045 48.040 ;
        RECT 24.025 46.290 25.085 48.650 ;
        RECT 25.485 47.015 25.655 52.055 ;
        RECT 26.275 47.015 26.445 52.055 ;
        RECT 25.715 46.630 26.215 46.800 ;
        RECT 26.845 46.290 27.015 52.780 ;
        RECT 27.645 52.270 28.145 52.440 ;
        RECT 27.415 47.015 27.585 52.055 ;
        RECT 28.205 47.015 28.375 52.055 ;
        RECT 27.645 46.630 28.145 46.800 ;
        RECT 28.775 46.290 30.165 52.780 ;
        RECT 30.365 66.080 41.365 66.950 ;
        RECT 30.365 54.940 32.035 66.080 ;
        RECT 32.665 65.565 37.665 65.735 ;
        RECT 32.435 55.310 32.605 65.350 ;
        RECT 37.725 55.310 37.895 65.350 ;
        RECT 38.295 54.940 38.465 66.080 ;
        RECT 39.095 65.565 40.095 65.735 ;
        RECT 38.865 55.310 39.035 65.350 ;
        RECT 40.155 55.310 40.325 65.350 ;
        RECT 40.725 54.940 41.365 66.080 ;
        RECT 30.365 52.870 41.365 54.940 ;
        RECT 30.365 49.380 32.205 52.870 ;
        RECT 33.965 52.790 41.365 52.870 ;
        RECT 32.835 52.360 33.335 52.530 ;
        RECT 32.605 50.105 32.775 52.145 ;
        RECT 33.395 50.105 33.565 52.145 ;
        RECT 32.835 49.720 33.335 49.890 ;
        RECT 33.965 49.380 36.285 52.790 ;
        RECT 36.915 52.280 37.415 52.450 ;
        RECT 30.365 48.660 36.285 49.380 ;
        RECT 24.025 45.800 30.165 46.290 ;
        RECT 30.335 48.050 34.245 48.270 ;
        RECT 19.135 45.370 23.045 45.640 ;
        RECT 30.335 45.650 32.055 48.050 ;
        RECT 32.685 47.540 33.185 47.710 ;
        RECT 32.455 46.330 32.625 47.370 ;
        RECT 33.245 46.330 33.415 47.370 ;
        RECT 32.685 45.990 33.185 46.160 ;
        RECT 33.815 45.650 34.245 48.050 ;
        RECT 35.225 46.300 36.285 48.660 ;
        RECT 36.685 47.025 36.855 52.065 ;
        RECT 37.475 47.025 37.645 52.065 ;
        RECT 36.915 46.640 37.415 46.810 ;
        RECT 38.045 46.300 38.215 52.790 ;
        RECT 38.845 52.280 39.345 52.450 ;
        RECT 38.615 47.025 38.785 52.065 ;
        RECT 39.405 47.025 39.575 52.065 ;
        RECT 38.845 46.640 39.345 46.810 ;
        RECT 39.975 46.300 41.365 52.790 ;
        RECT 41.585 66.050 52.585 66.920 ;
        RECT 41.585 54.910 43.255 66.050 ;
        RECT 43.885 65.535 48.885 65.705 ;
        RECT 43.655 55.280 43.825 65.320 ;
        RECT 48.945 55.280 49.115 65.320 ;
        RECT 49.515 54.910 49.685 66.050 ;
        RECT 50.315 65.535 51.315 65.705 ;
        RECT 50.085 55.280 50.255 65.320 ;
        RECT 51.375 55.280 51.545 65.320 ;
        RECT 51.945 54.910 52.585 66.050 ;
        RECT 41.585 52.840 52.585 54.910 ;
        RECT 41.585 49.350 43.425 52.840 ;
        RECT 45.185 52.760 52.585 52.840 ;
        RECT 44.055 52.330 44.555 52.500 ;
        RECT 43.825 50.075 43.995 52.115 ;
        RECT 44.615 50.075 44.785 52.115 ;
        RECT 44.055 49.690 44.555 49.860 ;
        RECT 45.185 49.350 47.505 52.760 ;
        RECT 48.135 52.250 48.635 52.420 ;
        RECT 41.585 48.630 47.505 49.350 ;
        RECT 35.225 45.810 41.365 46.300 ;
        RECT 41.555 48.020 45.465 48.240 ;
        RECT 30.335 45.380 34.245 45.650 ;
        RECT 41.555 45.620 43.275 48.020 ;
        RECT 43.905 47.510 44.405 47.680 ;
        RECT 43.675 46.300 43.845 47.340 ;
        RECT 44.465 46.300 44.635 47.340 ;
        RECT 43.905 45.960 44.405 46.130 ;
        RECT 45.035 45.620 45.465 48.020 ;
        RECT 46.445 46.270 47.505 48.630 ;
        RECT 47.905 46.995 48.075 52.035 ;
        RECT 48.695 46.995 48.865 52.035 ;
        RECT 48.135 46.610 48.635 46.780 ;
        RECT 49.265 46.270 49.435 52.760 ;
        RECT 50.065 52.250 50.565 52.420 ;
        RECT 49.835 46.995 50.005 52.035 ;
        RECT 50.625 46.995 50.795 52.035 ;
        RECT 50.065 46.610 50.565 46.780 ;
        RECT 51.195 46.270 52.585 52.760 ;
        RECT 52.835 66.030 63.835 66.900 ;
        RECT 52.835 54.890 54.505 66.030 ;
        RECT 55.135 65.515 60.135 65.685 ;
        RECT 54.905 55.260 55.075 65.300 ;
        RECT 60.195 55.260 60.365 65.300 ;
        RECT 60.765 54.890 60.935 66.030 ;
        RECT 61.565 65.515 62.565 65.685 ;
        RECT 61.335 55.260 61.505 65.300 ;
        RECT 62.625 55.260 62.795 65.300 ;
        RECT 63.195 54.890 63.835 66.030 ;
        RECT 52.835 52.820 63.835 54.890 ;
        RECT 52.835 49.330 54.675 52.820 ;
        RECT 56.435 52.740 63.835 52.820 ;
        RECT 55.305 52.310 55.805 52.480 ;
        RECT 55.075 50.055 55.245 52.095 ;
        RECT 55.865 50.055 56.035 52.095 ;
        RECT 55.305 49.670 55.805 49.840 ;
        RECT 56.435 49.330 58.755 52.740 ;
        RECT 59.385 52.230 59.885 52.400 ;
        RECT 52.835 48.610 58.755 49.330 ;
        RECT 46.445 45.780 52.585 46.270 ;
        RECT 52.805 48.000 56.715 48.220 ;
        RECT 41.555 45.350 45.465 45.620 ;
        RECT 52.805 45.600 54.525 48.000 ;
        RECT 55.155 47.490 55.655 47.660 ;
        RECT 54.925 46.280 55.095 47.320 ;
        RECT 55.715 46.280 55.885 47.320 ;
        RECT 55.155 45.940 55.655 46.110 ;
        RECT 56.285 45.600 56.715 48.000 ;
        RECT 57.695 46.250 58.755 48.610 ;
        RECT 59.155 46.975 59.325 52.015 ;
        RECT 59.945 46.975 60.115 52.015 ;
        RECT 59.385 46.590 59.885 46.760 ;
        RECT 60.515 46.250 60.685 52.740 ;
        RECT 61.315 52.230 61.815 52.400 ;
        RECT 61.085 46.975 61.255 52.015 ;
        RECT 61.875 46.975 62.045 52.015 ;
        RECT 61.315 46.590 61.815 46.760 ;
        RECT 62.445 46.250 63.835 52.740 ;
        RECT 64.055 66.020 75.055 66.890 ;
        RECT 64.055 54.880 65.725 66.020 ;
        RECT 66.355 65.505 71.355 65.675 ;
        RECT 66.125 55.250 66.295 65.290 ;
        RECT 71.415 55.250 71.585 65.290 ;
        RECT 71.985 54.880 72.155 66.020 ;
        RECT 72.785 65.505 73.785 65.675 ;
        RECT 72.555 55.250 72.725 65.290 ;
        RECT 73.845 55.250 74.015 65.290 ;
        RECT 74.415 54.880 75.055 66.020 ;
        RECT 64.055 52.810 75.055 54.880 ;
        RECT 64.055 49.320 65.895 52.810 ;
        RECT 67.655 52.730 75.055 52.810 ;
        RECT 66.525 52.300 67.025 52.470 ;
        RECT 66.295 50.045 66.465 52.085 ;
        RECT 67.085 50.045 67.255 52.085 ;
        RECT 66.525 49.660 67.025 49.830 ;
        RECT 67.655 49.320 69.975 52.730 ;
        RECT 70.605 52.220 71.105 52.390 ;
        RECT 64.055 48.600 69.975 49.320 ;
        RECT 57.695 45.760 63.835 46.250 ;
        RECT 64.025 47.990 67.935 48.210 ;
        RECT 52.805 45.330 56.715 45.600 ;
        RECT 64.025 45.590 65.745 47.990 ;
        RECT 66.375 47.480 66.875 47.650 ;
        RECT 66.145 46.270 66.315 47.310 ;
        RECT 66.935 46.270 67.105 47.310 ;
        RECT 66.375 45.930 66.875 46.100 ;
        RECT 67.505 45.590 67.935 47.990 ;
        RECT 68.915 46.240 69.975 48.600 ;
        RECT 70.375 46.965 70.545 52.005 ;
        RECT 71.165 46.965 71.335 52.005 ;
        RECT 70.605 46.580 71.105 46.750 ;
        RECT 71.735 46.240 71.905 52.730 ;
        RECT 72.535 52.220 73.035 52.390 ;
        RECT 72.305 46.965 72.475 52.005 ;
        RECT 73.095 46.965 73.265 52.005 ;
        RECT 72.535 46.580 73.035 46.750 ;
        RECT 73.665 46.240 75.055 52.730 ;
        RECT 75.295 66.010 86.295 66.880 ;
        RECT 75.295 54.870 76.965 66.010 ;
        RECT 77.595 65.495 82.595 65.665 ;
        RECT 77.365 55.240 77.535 65.280 ;
        RECT 82.655 55.240 82.825 65.280 ;
        RECT 83.225 54.870 83.395 66.010 ;
        RECT 84.025 65.495 85.025 65.665 ;
        RECT 83.795 55.240 83.965 65.280 ;
        RECT 85.085 55.240 85.255 65.280 ;
        RECT 85.655 54.870 86.295 66.010 ;
        RECT 75.295 52.800 86.295 54.870 ;
        RECT 75.295 49.310 77.135 52.800 ;
        RECT 78.895 52.720 86.295 52.800 ;
        RECT 77.765 52.290 78.265 52.460 ;
        RECT 77.535 50.035 77.705 52.075 ;
        RECT 78.325 50.035 78.495 52.075 ;
        RECT 77.765 49.650 78.265 49.820 ;
        RECT 78.895 49.310 81.215 52.720 ;
        RECT 81.845 52.210 82.345 52.380 ;
        RECT 75.295 48.590 81.215 49.310 ;
        RECT 68.915 45.750 75.055 46.240 ;
        RECT 75.265 47.980 79.175 48.200 ;
        RECT 64.025 45.320 67.935 45.590 ;
        RECT 75.265 45.580 76.985 47.980 ;
        RECT 77.615 47.470 78.115 47.640 ;
        RECT 77.385 46.260 77.555 47.300 ;
        RECT 78.175 46.260 78.345 47.300 ;
        RECT 77.615 45.920 78.115 46.090 ;
        RECT 78.745 45.580 79.175 47.980 ;
        RECT 80.155 46.230 81.215 48.590 ;
        RECT 81.615 46.955 81.785 51.995 ;
        RECT 82.405 46.955 82.575 51.995 ;
        RECT 81.845 46.570 82.345 46.740 ;
        RECT 82.975 46.230 83.145 52.720 ;
        RECT 83.775 52.210 84.275 52.380 ;
        RECT 83.545 46.955 83.715 51.995 ;
        RECT 84.335 46.955 84.505 51.995 ;
        RECT 83.775 46.570 84.275 46.740 ;
        RECT 84.905 46.230 86.295 52.720 ;
        RECT 86.545 66.020 97.545 66.890 ;
        RECT 131.125 66.880 140.025 66.890 ;
        RECT 86.545 54.880 88.215 66.020 ;
        RECT 88.845 65.505 93.845 65.675 ;
        RECT 88.615 55.250 88.785 65.290 ;
        RECT 93.905 55.250 94.075 65.290 ;
        RECT 94.475 54.880 94.645 66.020 ;
        RECT 95.275 65.505 96.275 65.675 ;
        RECT 95.045 55.250 95.215 65.290 ;
        RECT 96.335 55.250 96.505 65.290 ;
        RECT 96.905 54.880 97.545 66.020 ;
        RECT 86.545 52.810 97.545 54.880 ;
        RECT 86.545 49.320 88.385 52.810 ;
        RECT 90.145 52.730 97.545 52.810 ;
        RECT 89.015 52.300 89.515 52.470 ;
        RECT 88.785 50.045 88.955 52.085 ;
        RECT 89.575 50.045 89.745 52.085 ;
        RECT 89.015 49.660 89.515 49.830 ;
        RECT 90.145 49.320 92.465 52.730 ;
        RECT 93.095 52.220 93.595 52.390 ;
        RECT 86.545 48.600 92.465 49.320 ;
        RECT 80.155 45.740 86.295 46.230 ;
        RECT 86.515 47.990 90.425 48.210 ;
        RECT 75.265 45.310 79.175 45.580 ;
        RECT 86.515 45.590 88.235 47.990 ;
        RECT 88.865 47.480 89.365 47.650 ;
        RECT 88.635 46.270 88.805 47.310 ;
        RECT 89.425 46.270 89.595 47.310 ;
        RECT 88.865 45.930 89.365 46.100 ;
        RECT 89.995 45.590 90.425 47.990 ;
        RECT 91.405 46.240 92.465 48.600 ;
        RECT 92.865 46.965 93.035 52.005 ;
        RECT 93.655 46.965 93.825 52.005 ;
        RECT 93.095 46.580 93.595 46.750 ;
        RECT 94.225 46.240 94.395 52.730 ;
        RECT 95.025 52.220 95.525 52.390 ;
        RECT 94.795 46.965 94.965 52.005 ;
        RECT 95.585 46.965 95.755 52.005 ;
        RECT 95.025 46.580 95.525 46.750 ;
        RECT 96.155 46.240 97.545 52.730 ;
        RECT 97.825 66.010 108.825 66.880 ;
        RECT 97.825 54.870 99.495 66.010 ;
        RECT 100.125 65.495 105.125 65.665 ;
        RECT 99.895 55.240 100.065 65.280 ;
        RECT 105.185 55.240 105.355 65.280 ;
        RECT 105.755 54.870 105.925 66.010 ;
        RECT 106.555 65.495 107.555 65.665 ;
        RECT 106.325 55.240 106.495 65.280 ;
        RECT 107.615 55.240 107.785 65.280 ;
        RECT 108.185 54.870 108.825 66.010 ;
        RECT 97.825 52.800 108.825 54.870 ;
        RECT 97.825 49.310 99.665 52.800 ;
        RECT 101.425 52.720 108.825 52.800 ;
        RECT 100.295 52.290 100.795 52.460 ;
        RECT 100.065 50.035 100.235 52.075 ;
        RECT 100.855 50.035 101.025 52.075 ;
        RECT 100.295 49.650 100.795 49.820 ;
        RECT 101.425 49.310 103.745 52.720 ;
        RECT 104.375 52.210 104.875 52.380 ;
        RECT 97.825 48.590 103.745 49.310 ;
        RECT 91.405 45.750 97.545 46.240 ;
        RECT 97.795 47.980 101.705 48.200 ;
        RECT 86.515 45.320 90.425 45.590 ;
        RECT 97.795 45.580 99.515 47.980 ;
        RECT 100.145 47.470 100.645 47.640 ;
        RECT 99.915 46.260 100.085 47.300 ;
        RECT 100.705 46.260 100.875 47.300 ;
        RECT 100.145 45.920 100.645 46.090 ;
        RECT 101.275 45.580 101.705 47.980 ;
        RECT 102.685 46.230 103.745 48.590 ;
        RECT 104.145 46.955 104.315 51.995 ;
        RECT 104.935 46.955 105.105 51.995 ;
        RECT 104.375 46.570 104.875 46.740 ;
        RECT 105.505 46.230 105.675 52.720 ;
        RECT 106.305 52.210 106.805 52.380 ;
        RECT 106.075 46.955 106.245 51.995 ;
        RECT 106.865 46.955 107.035 51.995 ;
        RECT 106.305 46.570 106.805 46.740 ;
        RECT 107.435 46.230 108.825 52.720 ;
        RECT 109.095 66.010 120.095 66.880 ;
        RECT 109.095 54.870 110.765 66.010 ;
        RECT 111.395 65.495 116.395 65.665 ;
        RECT 111.165 55.240 111.335 65.280 ;
        RECT 116.455 55.240 116.625 65.280 ;
        RECT 117.025 54.870 117.195 66.010 ;
        RECT 117.825 65.495 118.825 65.665 ;
        RECT 117.595 55.240 117.765 65.280 ;
        RECT 118.885 55.240 119.055 65.280 ;
        RECT 119.455 54.870 120.095 66.010 ;
        RECT 109.095 52.800 120.095 54.870 ;
        RECT 109.095 49.310 110.935 52.800 ;
        RECT 112.695 52.720 120.095 52.800 ;
        RECT 111.565 52.290 112.065 52.460 ;
        RECT 111.335 50.035 111.505 52.075 ;
        RECT 112.125 50.035 112.295 52.075 ;
        RECT 111.565 49.650 112.065 49.820 ;
        RECT 112.695 49.310 115.015 52.720 ;
        RECT 115.645 52.210 116.145 52.380 ;
        RECT 109.095 48.590 115.015 49.310 ;
        RECT 102.685 45.740 108.825 46.230 ;
        RECT 109.065 47.980 112.975 48.200 ;
        RECT 97.795 45.310 101.705 45.580 ;
        RECT 109.065 45.580 110.785 47.980 ;
        RECT 111.415 47.470 111.915 47.640 ;
        RECT 111.185 46.260 111.355 47.300 ;
        RECT 111.975 46.260 112.145 47.300 ;
        RECT 111.415 45.920 111.915 46.090 ;
        RECT 112.545 45.580 112.975 47.980 ;
        RECT 113.955 46.230 115.015 48.590 ;
        RECT 115.415 46.955 115.585 51.995 ;
        RECT 116.205 46.955 116.375 51.995 ;
        RECT 115.645 46.570 116.145 46.740 ;
        RECT 116.775 46.230 116.945 52.720 ;
        RECT 117.575 52.210 118.075 52.380 ;
        RECT 117.345 46.955 117.515 51.995 ;
        RECT 118.135 46.955 118.305 51.995 ;
        RECT 117.575 46.570 118.075 46.740 ;
        RECT 118.705 46.230 120.095 52.720 ;
        RECT 120.345 66.010 140.025 66.880 ;
        RECT 120.345 54.870 122.015 66.010 ;
        RECT 122.645 65.495 127.645 65.665 ;
        RECT 122.415 55.240 122.585 65.280 ;
        RECT 127.705 55.240 127.875 65.280 ;
        RECT 128.275 54.870 128.445 66.010 ;
        RECT 130.705 65.980 140.025 66.010 ;
        RECT 129.075 65.495 130.075 65.665 ;
        RECT 128.845 55.240 129.015 65.280 ;
        RECT 130.135 55.240 130.305 65.280 ;
        RECT 130.705 54.870 132.765 65.980 ;
        RECT 133.395 65.465 138.395 65.635 ;
        RECT 133.165 55.210 133.335 65.250 ;
        RECT 138.455 55.210 138.625 65.250 ;
        RECT 120.345 54.840 132.765 54.870 ;
        RECT 139.025 54.840 140.025 65.980 ;
        RECT 120.345 54.720 140.025 54.840 ;
        RECT 120.345 53.550 140.035 54.720 ;
        RECT 120.345 52.800 131.345 53.550 ;
        RECT 120.345 49.310 122.185 52.800 ;
        RECT 123.945 52.720 131.345 52.800 ;
        RECT 122.815 52.290 123.315 52.460 ;
        RECT 122.585 50.035 122.755 52.075 ;
        RECT 123.375 50.035 123.545 52.075 ;
        RECT 122.815 49.650 123.315 49.820 ;
        RECT 123.945 49.310 126.265 52.720 ;
        RECT 126.895 52.210 127.395 52.380 ;
        RECT 120.345 48.590 126.265 49.310 ;
        RECT 113.955 45.740 120.095 46.230 ;
        RECT 120.315 47.980 124.225 48.200 ;
        RECT 109.065 45.310 112.975 45.580 ;
        RECT 120.315 45.580 122.035 47.980 ;
        RECT 122.665 47.470 123.165 47.640 ;
        RECT 122.435 46.260 122.605 47.300 ;
        RECT 123.225 46.260 123.395 47.300 ;
        RECT 122.665 45.920 123.165 46.090 ;
        RECT 123.795 45.580 124.225 47.980 ;
        RECT 125.205 46.230 126.265 48.590 ;
        RECT 126.665 46.955 126.835 51.995 ;
        RECT 127.455 46.955 127.625 51.995 ;
        RECT 126.895 46.570 127.395 46.740 ;
        RECT 128.025 46.230 128.195 52.720 ;
        RECT 128.825 52.210 129.325 52.380 ;
        RECT 128.595 46.955 128.765 51.995 ;
        RECT 129.385 46.955 129.555 51.995 ;
        RECT 128.825 46.570 129.325 46.740 ;
        RECT 129.955 46.230 131.345 52.720 ;
        RECT 125.205 45.740 131.345 46.230 ;
        RECT 120.315 45.310 124.225 45.580 ;
        RECT 25.695 39.770 29.605 40.040 ;
        RECT 18.575 39.120 24.715 39.610 ;
        RECT 18.575 32.630 19.965 39.120 ;
        RECT 20.595 38.610 21.095 38.780 ;
        RECT 20.365 33.355 20.535 38.395 ;
        RECT 21.155 33.355 21.325 38.395 ;
        RECT 20.595 32.970 21.095 33.140 ;
        RECT 21.725 32.630 21.895 39.120 ;
        RECT 22.525 38.610 23.025 38.780 ;
        RECT 22.295 33.355 22.465 38.395 ;
        RECT 23.085 33.355 23.255 38.395 ;
        RECT 23.655 36.760 24.715 39.120 ;
        RECT 25.695 37.370 26.125 39.770 ;
        RECT 26.755 39.260 27.255 39.430 ;
        RECT 26.525 38.050 26.695 39.090 ;
        RECT 27.315 38.050 27.485 39.090 ;
        RECT 26.755 37.710 27.255 37.880 ;
        RECT 27.885 37.370 29.605 39.770 ;
        RECT 36.975 39.770 40.885 40.040 ;
        RECT 25.695 37.150 29.605 37.370 ;
        RECT 29.855 39.120 35.995 39.610 ;
        RECT 23.655 36.040 29.575 36.760 ;
        RECT 22.525 32.970 23.025 33.140 ;
        RECT 23.655 32.630 25.975 36.040 ;
        RECT 26.605 35.530 27.105 35.700 ;
        RECT 26.375 33.275 26.545 35.315 ;
        RECT 27.165 33.275 27.335 35.315 ;
        RECT 26.605 32.890 27.105 33.060 ;
        RECT 18.575 32.550 25.975 32.630 ;
        RECT 27.735 32.550 29.575 36.040 ;
        RECT 18.575 30.480 29.575 32.550 ;
        RECT 18.575 19.340 19.215 30.480 ;
        RECT 19.615 20.070 19.785 30.110 ;
        RECT 20.905 20.070 21.075 30.110 ;
        RECT 19.845 19.685 20.845 19.855 ;
        RECT 21.475 19.340 21.645 30.480 ;
        RECT 22.045 20.070 22.215 30.110 ;
        RECT 27.335 20.070 27.505 30.110 ;
        RECT 22.275 19.685 27.275 19.855 ;
        RECT 27.905 19.340 29.575 30.480 ;
        RECT 18.575 18.470 29.575 19.340 ;
        RECT 29.855 32.630 31.245 39.120 ;
        RECT 31.875 38.610 32.375 38.780 ;
        RECT 31.645 33.355 31.815 38.395 ;
        RECT 32.435 33.355 32.605 38.395 ;
        RECT 31.875 32.970 32.375 33.140 ;
        RECT 33.005 32.630 33.175 39.120 ;
        RECT 33.805 38.610 34.305 38.780 ;
        RECT 33.575 33.355 33.745 38.395 ;
        RECT 34.365 33.355 34.535 38.395 ;
        RECT 34.935 36.760 35.995 39.120 ;
        RECT 36.975 37.370 37.405 39.770 ;
        RECT 38.035 39.260 38.535 39.430 ;
        RECT 37.805 38.050 37.975 39.090 ;
        RECT 38.595 38.050 38.765 39.090 ;
        RECT 38.035 37.710 38.535 37.880 ;
        RECT 39.165 37.370 40.885 39.770 ;
        RECT 48.265 39.750 52.175 40.020 ;
        RECT 36.975 37.150 40.885 37.370 ;
        RECT 41.145 39.100 47.285 39.590 ;
        RECT 34.935 36.040 40.855 36.760 ;
        RECT 33.805 32.970 34.305 33.140 ;
        RECT 34.935 32.630 37.255 36.040 ;
        RECT 37.885 35.530 38.385 35.700 ;
        RECT 37.655 33.275 37.825 35.315 ;
        RECT 38.445 33.275 38.615 35.315 ;
        RECT 37.885 32.890 38.385 33.060 ;
        RECT 29.855 32.550 37.255 32.630 ;
        RECT 39.015 32.550 40.855 36.040 ;
        RECT 29.855 30.480 40.855 32.550 ;
        RECT 29.855 19.340 30.495 30.480 ;
        RECT 30.895 20.070 31.065 30.110 ;
        RECT 32.185 20.070 32.355 30.110 ;
        RECT 31.125 19.685 32.125 19.855 ;
        RECT 32.755 19.340 32.925 30.480 ;
        RECT 33.325 20.070 33.495 30.110 ;
        RECT 38.615 20.070 38.785 30.110 ;
        RECT 33.555 19.685 38.555 19.855 ;
        RECT 39.185 19.340 40.855 30.480 ;
        RECT 29.855 18.470 40.855 19.340 ;
        RECT 41.145 32.610 42.535 39.100 ;
        RECT 43.165 38.590 43.665 38.760 ;
        RECT 42.935 33.335 43.105 38.375 ;
        RECT 43.725 33.335 43.895 38.375 ;
        RECT 43.165 32.950 43.665 33.120 ;
        RECT 44.295 32.610 44.465 39.100 ;
        RECT 45.095 38.590 45.595 38.760 ;
        RECT 44.865 33.335 45.035 38.375 ;
        RECT 45.655 33.335 45.825 38.375 ;
        RECT 46.225 36.740 47.285 39.100 ;
        RECT 48.265 37.350 48.695 39.750 ;
        RECT 49.325 39.240 49.825 39.410 ;
        RECT 49.095 38.030 49.265 39.070 ;
        RECT 49.885 38.030 50.055 39.070 ;
        RECT 49.325 37.690 49.825 37.860 ;
        RECT 50.455 37.350 52.175 39.750 ;
        RECT 59.485 39.750 63.395 40.020 ;
        RECT 48.265 37.130 52.175 37.350 ;
        RECT 52.365 39.100 58.505 39.590 ;
        RECT 46.225 36.020 52.145 36.740 ;
        RECT 45.095 32.950 45.595 33.120 ;
        RECT 46.225 32.610 48.545 36.020 ;
        RECT 49.175 35.510 49.675 35.680 ;
        RECT 48.945 33.255 49.115 35.295 ;
        RECT 49.735 33.255 49.905 35.295 ;
        RECT 49.175 32.870 49.675 33.040 ;
        RECT 41.145 32.530 48.545 32.610 ;
        RECT 50.305 32.530 52.145 36.020 ;
        RECT 41.145 30.460 52.145 32.530 ;
        RECT 41.145 19.320 41.785 30.460 ;
        RECT 42.185 20.050 42.355 30.090 ;
        RECT 43.475 20.050 43.645 30.090 ;
        RECT 42.415 19.665 43.415 19.835 ;
        RECT 44.045 19.320 44.215 30.460 ;
        RECT 44.615 20.050 44.785 30.090 ;
        RECT 49.905 20.050 50.075 30.090 ;
        RECT 44.845 19.665 49.845 19.835 ;
        RECT 50.475 19.320 52.145 30.460 ;
        RECT 41.145 18.450 52.145 19.320 ;
        RECT 52.365 32.610 53.755 39.100 ;
        RECT 54.385 38.590 54.885 38.760 ;
        RECT 54.155 33.335 54.325 38.375 ;
        RECT 54.945 33.335 55.115 38.375 ;
        RECT 54.385 32.950 54.885 33.120 ;
        RECT 55.515 32.610 55.685 39.100 ;
        RECT 56.315 38.590 56.815 38.760 ;
        RECT 56.085 33.335 56.255 38.375 ;
        RECT 56.875 33.335 57.045 38.375 ;
        RECT 57.445 36.740 58.505 39.100 ;
        RECT 59.485 37.350 59.915 39.750 ;
        RECT 60.545 39.240 61.045 39.410 ;
        RECT 60.315 38.030 60.485 39.070 ;
        RECT 61.105 38.030 61.275 39.070 ;
        RECT 60.545 37.690 61.045 37.860 ;
        RECT 61.675 37.350 63.395 39.750 ;
        RECT 70.685 39.750 74.595 40.020 ;
        RECT 59.485 37.130 63.395 37.350 ;
        RECT 63.565 39.100 69.705 39.590 ;
        RECT 57.445 36.020 63.365 36.740 ;
        RECT 56.315 32.950 56.815 33.120 ;
        RECT 57.445 32.610 59.765 36.020 ;
        RECT 60.395 35.510 60.895 35.680 ;
        RECT 60.165 33.255 60.335 35.295 ;
        RECT 60.955 33.255 61.125 35.295 ;
        RECT 60.395 32.870 60.895 33.040 ;
        RECT 52.365 32.530 59.765 32.610 ;
        RECT 61.525 32.530 63.365 36.020 ;
        RECT 52.365 30.460 63.365 32.530 ;
        RECT 52.365 19.320 53.005 30.460 ;
        RECT 53.405 20.050 53.575 30.090 ;
        RECT 54.695 20.050 54.865 30.090 ;
        RECT 53.635 19.665 54.635 19.835 ;
        RECT 55.265 19.320 55.435 30.460 ;
        RECT 55.835 20.050 56.005 30.090 ;
        RECT 61.125 20.050 61.295 30.090 ;
        RECT 56.065 19.665 61.065 19.835 ;
        RECT 61.695 19.320 63.365 30.460 ;
        RECT 52.365 18.450 63.365 19.320 ;
        RECT 63.565 32.610 64.955 39.100 ;
        RECT 65.585 38.590 66.085 38.760 ;
        RECT 65.355 33.335 65.525 38.375 ;
        RECT 66.145 33.335 66.315 38.375 ;
        RECT 65.585 32.950 66.085 33.120 ;
        RECT 66.715 32.610 66.885 39.100 ;
        RECT 67.515 38.590 68.015 38.760 ;
        RECT 67.285 33.335 67.455 38.375 ;
        RECT 68.075 33.335 68.245 38.375 ;
        RECT 68.645 36.740 69.705 39.100 ;
        RECT 70.685 37.350 71.115 39.750 ;
        RECT 71.745 39.240 72.245 39.410 ;
        RECT 71.515 38.030 71.685 39.070 ;
        RECT 72.305 38.030 72.475 39.070 ;
        RECT 71.745 37.690 72.245 37.860 ;
        RECT 72.875 37.350 74.595 39.750 ;
        RECT 81.975 39.740 85.885 40.010 ;
        RECT 70.685 37.130 74.595 37.350 ;
        RECT 74.855 39.090 80.995 39.580 ;
        RECT 68.645 36.020 74.565 36.740 ;
        RECT 67.515 32.950 68.015 33.120 ;
        RECT 68.645 32.610 70.965 36.020 ;
        RECT 71.595 35.510 72.095 35.680 ;
        RECT 71.365 33.255 71.535 35.295 ;
        RECT 72.155 33.255 72.325 35.295 ;
        RECT 71.595 32.870 72.095 33.040 ;
        RECT 63.565 32.530 70.965 32.610 ;
        RECT 72.725 32.530 74.565 36.020 ;
        RECT 63.565 30.460 74.565 32.530 ;
        RECT 63.565 19.320 64.205 30.460 ;
        RECT 64.605 20.050 64.775 30.090 ;
        RECT 65.895 20.050 66.065 30.090 ;
        RECT 64.835 19.665 65.835 19.835 ;
        RECT 66.465 19.320 66.635 30.460 ;
        RECT 67.035 20.050 67.205 30.090 ;
        RECT 72.325 20.050 72.495 30.090 ;
        RECT 67.265 19.665 72.265 19.835 ;
        RECT 72.895 19.320 74.565 30.460 ;
        RECT 63.565 18.450 74.565 19.320 ;
        RECT 74.855 32.600 76.245 39.090 ;
        RECT 76.875 38.580 77.375 38.750 ;
        RECT 76.645 33.325 76.815 38.365 ;
        RECT 77.435 33.325 77.605 38.365 ;
        RECT 76.875 32.940 77.375 33.110 ;
        RECT 78.005 32.600 78.175 39.090 ;
        RECT 78.805 38.580 79.305 38.750 ;
        RECT 78.575 33.325 78.745 38.365 ;
        RECT 79.365 33.325 79.535 38.365 ;
        RECT 79.935 36.730 80.995 39.090 ;
        RECT 81.975 37.340 82.405 39.740 ;
        RECT 83.035 39.230 83.535 39.400 ;
        RECT 82.805 38.020 82.975 39.060 ;
        RECT 83.595 38.020 83.765 39.060 ;
        RECT 83.035 37.680 83.535 37.850 ;
        RECT 84.165 37.340 85.885 39.740 ;
        RECT 93.215 39.760 97.125 40.030 ;
        RECT 81.975 37.120 85.885 37.340 ;
        RECT 86.095 39.110 92.235 39.600 ;
        RECT 79.935 36.010 85.855 36.730 ;
        RECT 78.805 32.940 79.305 33.110 ;
        RECT 79.935 32.600 82.255 36.010 ;
        RECT 82.885 35.500 83.385 35.670 ;
        RECT 82.655 33.245 82.825 35.285 ;
        RECT 83.445 33.245 83.615 35.285 ;
        RECT 82.885 32.860 83.385 33.030 ;
        RECT 74.855 32.520 82.255 32.600 ;
        RECT 84.015 32.520 85.855 36.010 ;
        RECT 74.855 30.450 85.855 32.520 ;
        RECT 74.855 19.310 75.495 30.450 ;
        RECT 75.895 20.040 76.065 30.080 ;
        RECT 77.185 20.040 77.355 30.080 ;
        RECT 76.125 19.655 77.125 19.825 ;
        RECT 77.755 19.310 77.925 30.450 ;
        RECT 78.325 20.040 78.495 30.080 ;
        RECT 83.615 20.040 83.785 30.080 ;
        RECT 78.555 19.655 83.555 19.825 ;
        RECT 84.185 19.310 85.855 30.450 ;
        RECT 74.855 18.440 85.855 19.310 ;
        RECT 86.095 32.620 87.485 39.110 ;
        RECT 88.115 38.600 88.615 38.770 ;
        RECT 87.885 33.345 88.055 38.385 ;
        RECT 88.675 33.345 88.845 38.385 ;
        RECT 88.115 32.960 88.615 33.130 ;
        RECT 89.245 32.620 89.415 39.110 ;
        RECT 90.045 38.600 90.545 38.770 ;
        RECT 89.815 33.345 89.985 38.385 ;
        RECT 90.605 33.345 90.775 38.385 ;
        RECT 91.175 36.750 92.235 39.110 ;
        RECT 93.215 37.360 93.645 39.760 ;
        RECT 94.275 39.250 94.775 39.420 ;
        RECT 94.045 38.040 94.215 39.080 ;
        RECT 94.835 38.040 95.005 39.080 ;
        RECT 94.275 37.700 94.775 37.870 ;
        RECT 95.405 37.360 97.125 39.760 ;
        RECT 104.425 39.780 108.335 40.050 ;
        RECT 93.215 37.140 97.125 37.360 ;
        RECT 97.305 39.130 103.445 39.620 ;
        RECT 91.175 36.030 97.095 36.750 ;
        RECT 90.045 32.960 90.545 33.130 ;
        RECT 91.175 32.620 93.495 36.030 ;
        RECT 94.125 35.520 94.625 35.690 ;
        RECT 93.895 33.265 94.065 35.305 ;
        RECT 94.685 33.265 94.855 35.305 ;
        RECT 94.125 32.880 94.625 33.050 ;
        RECT 86.095 32.540 93.495 32.620 ;
        RECT 95.255 32.540 97.095 36.030 ;
        RECT 86.095 30.470 97.095 32.540 ;
        RECT 86.095 19.330 86.735 30.470 ;
        RECT 87.135 20.060 87.305 30.100 ;
        RECT 88.425 20.060 88.595 30.100 ;
        RECT 87.365 19.675 88.365 19.845 ;
        RECT 88.995 19.330 89.165 30.470 ;
        RECT 89.565 20.060 89.735 30.100 ;
        RECT 94.855 20.060 95.025 30.100 ;
        RECT 89.795 19.675 94.795 19.845 ;
        RECT 95.425 19.330 97.095 30.470 ;
        RECT 86.095 18.460 97.095 19.330 ;
        RECT 97.305 32.640 98.695 39.130 ;
        RECT 99.325 38.620 99.825 38.790 ;
        RECT 99.095 33.365 99.265 38.405 ;
        RECT 99.885 33.365 100.055 38.405 ;
        RECT 99.325 32.980 99.825 33.150 ;
        RECT 100.455 32.640 100.625 39.130 ;
        RECT 101.255 38.620 101.755 38.790 ;
        RECT 101.025 33.365 101.195 38.405 ;
        RECT 101.815 33.365 101.985 38.405 ;
        RECT 102.385 36.770 103.445 39.130 ;
        RECT 104.425 37.380 104.855 39.780 ;
        RECT 105.485 39.270 105.985 39.440 ;
        RECT 105.255 38.060 105.425 39.100 ;
        RECT 106.045 38.060 106.215 39.100 ;
        RECT 105.485 37.720 105.985 37.890 ;
        RECT 106.615 37.380 108.335 39.780 ;
        RECT 115.625 39.820 119.535 40.090 ;
        RECT 104.425 37.160 108.335 37.380 ;
        RECT 108.505 39.170 114.645 39.660 ;
        RECT 102.385 36.050 108.305 36.770 ;
        RECT 101.255 32.980 101.755 33.150 ;
        RECT 102.385 32.640 104.705 36.050 ;
        RECT 105.335 35.540 105.835 35.710 ;
        RECT 105.105 33.285 105.275 35.325 ;
        RECT 105.895 33.285 106.065 35.325 ;
        RECT 105.335 32.900 105.835 33.070 ;
        RECT 97.305 32.560 104.705 32.640 ;
        RECT 106.465 32.560 108.305 36.050 ;
        RECT 97.305 30.490 108.305 32.560 ;
        RECT 97.305 19.350 97.945 30.490 ;
        RECT 98.345 20.080 98.515 30.120 ;
        RECT 99.635 20.080 99.805 30.120 ;
        RECT 98.575 19.695 99.575 19.865 ;
        RECT 100.205 19.350 100.375 30.490 ;
        RECT 100.775 20.080 100.945 30.120 ;
        RECT 106.065 20.080 106.235 30.120 ;
        RECT 101.005 19.695 106.005 19.865 ;
        RECT 106.635 19.350 108.305 30.490 ;
        RECT 97.305 18.480 108.305 19.350 ;
        RECT 108.505 32.680 109.895 39.170 ;
        RECT 110.525 38.660 111.025 38.830 ;
        RECT 110.295 33.405 110.465 38.445 ;
        RECT 111.085 33.405 111.255 38.445 ;
        RECT 110.525 33.020 111.025 33.190 ;
        RECT 111.655 32.680 111.825 39.170 ;
        RECT 112.455 38.660 112.955 38.830 ;
        RECT 112.225 33.405 112.395 38.445 ;
        RECT 113.015 33.405 113.185 38.445 ;
        RECT 113.585 36.810 114.645 39.170 ;
        RECT 115.625 37.420 116.055 39.820 ;
        RECT 116.685 39.310 117.185 39.480 ;
        RECT 116.455 38.100 116.625 39.140 ;
        RECT 117.245 38.100 117.415 39.140 ;
        RECT 116.685 37.760 117.185 37.930 ;
        RECT 117.815 37.420 119.535 39.820 ;
        RECT 126.835 39.840 130.745 40.110 ;
        RECT 115.625 37.200 119.535 37.420 ;
        RECT 119.715 39.190 125.855 39.680 ;
        RECT 113.585 36.090 119.505 36.810 ;
        RECT 112.455 33.020 112.955 33.190 ;
        RECT 113.585 32.680 115.905 36.090 ;
        RECT 116.535 35.580 117.035 35.750 ;
        RECT 116.305 33.325 116.475 35.365 ;
        RECT 117.095 33.325 117.265 35.365 ;
        RECT 116.535 32.940 117.035 33.110 ;
        RECT 108.505 32.600 115.905 32.680 ;
        RECT 117.665 32.600 119.505 36.090 ;
        RECT 108.505 30.530 119.505 32.600 ;
        RECT 108.505 19.390 109.145 30.530 ;
        RECT 109.545 20.120 109.715 30.160 ;
        RECT 110.835 20.120 111.005 30.160 ;
        RECT 109.775 19.735 110.775 19.905 ;
        RECT 111.405 19.390 111.575 30.530 ;
        RECT 111.975 20.120 112.145 30.160 ;
        RECT 117.265 20.120 117.435 30.160 ;
        RECT 112.205 19.735 117.205 19.905 ;
        RECT 117.835 19.390 119.505 30.530 ;
        RECT 108.505 18.520 119.505 19.390 ;
        RECT 119.715 32.700 121.105 39.190 ;
        RECT 121.735 38.680 122.235 38.850 ;
        RECT 121.505 33.425 121.675 38.465 ;
        RECT 122.295 33.425 122.465 38.465 ;
        RECT 121.735 33.040 122.235 33.210 ;
        RECT 122.865 32.700 123.035 39.190 ;
        RECT 123.665 38.680 124.165 38.850 ;
        RECT 123.435 33.425 123.605 38.465 ;
        RECT 124.225 33.425 124.395 38.465 ;
        RECT 124.795 36.830 125.855 39.190 ;
        RECT 126.835 37.440 127.265 39.840 ;
        RECT 127.895 39.330 128.395 39.500 ;
        RECT 127.665 38.120 127.835 39.160 ;
        RECT 128.455 38.120 128.625 39.160 ;
        RECT 127.895 37.780 128.395 37.950 ;
        RECT 129.025 37.440 130.745 39.840 ;
        RECT 126.835 37.220 130.745 37.440 ;
        RECT 124.795 36.110 130.715 36.830 ;
        RECT 123.665 33.040 124.165 33.210 ;
        RECT 124.795 32.700 127.115 36.110 ;
        RECT 127.745 35.600 128.245 35.770 ;
        RECT 127.515 33.345 127.685 35.385 ;
        RECT 128.305 33.345 128.475 35.385 ;
        RECT 127.745 32.960 128.245 33.130 ;
        RECT 119.715 32.620 127.115 32.700 ;
        RECT 128.875 32.620 130.715 36.110 ;
        RECT 119.715 31.140 130.715 32.620 ;
        RECT 119.715 30.550 139.465 31.140 ;
        RECT 119.715 19.410 120.355 30.550 ;
        RECT 120.755 20.140 120.925 30.180 ;
        RECT 122.045 20.140 122.215 30.180 ;
        RECT 120.985 19.755 121.985 19.925 ;
        RECT 122.615 19.410 122.785 30.550 ;
        RECT 129.045 30.520 139.465 30.550 ;
        RECT 123.185 20.140 123.355 30.180 ;
        RECT 128.475 20.140 128.645 30.180 ;
        RECT 123.415 19.755 128.415 19.925 ;
        RECT 129.045 19.410 132.075 30.520 ;
        RECT 132.475 20.110 132.645 30.150 ;
        RECT 137.765 20.110 137.935 30.150 ;
        RECT 132.705 19.725 137.705 19.895 ;
        RECT 119.715 19.380 132.075 19.410 ;
        RECT 138.335 19.380 139.465 30.520 ;
        RECT 119.715 18.540 139.465 19.380 ;
        RECT 131.925 18.520 139.465 18.540 ;
      LAYER met1 ;
        RECT 135.340 223.880 136.790 225.180 ;
        RECT 15.010 203.790 113.450 204.270 ;
        RECT 61.080 202.710 61.400 202.970 ;
        RECT 70.740 202.910 71.060 202.970 ;
        RECT 73.975 202.910 74.265 202.955 ;
        RECT 70.740 202.770 74.265 202.910 ;
        RECT 70.740 202.710 71.060 202.770 ;
        RECT 73.975 202.725 74.265 202.770 ;
        RECT 60.175 201.890 60.465 201.935 ;
        RECT 60.620 201.890 60.940 201.950 ;
        RECT 60.175 201.750 60.940 201.890 ;
        RECT 60.175 201.705 60.465 201.750 ;
        RECT 60.620 201.690 60.940 201.750 ;
        RECT 73.500 201.690 73.820 201.950 ;
        RECT 15.010 201.070 113.450 201.550 ;
        RECT 57.860 200.870 58.180 200.930 ;
        RECT 57.860 200.730 65.910 200.870 ;
        RECT 57.860 200.670 58.180 200.730 ;
        RECT 54.295 200.530 54.585 200.575 ;
        RECT 57.415 200.530 57.705 200.575 ;
        RECT 59.305 200.530 59.595 200.575 ;
        RECT 54.295 200.390 59.595 200.530 ;
        RECT 54.295 200.345 54.585 200.390 ;
        RECT 57.415 200.345 57.705 200.390 ;
        RECT 59.305 200.345 59.595 200.390 ;
        RECT 61.080 200.530 61.400 200.590 ;
        RECT 65.235 200.530 65.525 200.575 ;
        RECT 61.080 200.390 65.525 200.530 ;
        RECT 61.080 200.330 61.400 200.390 ;
        RECT 65.235 200.345 65.525 200.390 ;
        RECT 61.540 200.190 61.860 200.250 ;
        RECT 61.540 200.050 64.070 200.190 ;
        RECT 61.540 199.990 61.860 200.050 ;
        RECT 52.340 199.510 52.660 199.570 ;
        RECT 53.215 199.555 53.505 199.870 ;
        RECT 54.295 199.850 54.585 199.895 ;
        RECT 57.875 199.850 58.165 199.895 ;
        RECT 59.710 199.850 60.000 199.895 ;
        RECT 54.295 199.710 60.000 199.850 ;
        RECT 54.295 199.665 54.585 199.710 ;
        RECT 57.875 199.665 58.165 199.710 ;
        RECT 59.710 199.665 60.000 199.710 ;
        RECT 60.175 199.850 60.465 199.895 ;
        RECT 62.000 199.850 62.320 199.910 ;
        RECT 63.930 199.895 64.070 200.050 ;
        RECT 64.315 200.005 64.605 200.235 ;
        RECT 60.175 199.710 62.320 199.850 ;
        RECT 60.175 199.665 60.465 199.710 ;
        RECT 62.000 199.650 62.320 199.710 ;
        RECT 63.855 199.665 64.145 199.895 ;
        RECT 64.390 199.850 64.530 200.005 ;
        RECT 65.220 199.850 65.540 199.910 ;
        RECT 64.390 199.710 65.540 199.850 ;
        RECT 65.770 199.850 65.910 200.730 ;
        RECT 66.140 200.670 66.460 200.930 ;
        RECT 72.695 200.530 72.985 200.575 ;
        RECT 75.815 200.530 76.105 200.575 ;
        RECT 77.705 200.530 77.995 200.575 ;
        RECT 72.695 200.390 77.995 200.530 ;
        RECT 72.695 200.345 72.985 200.390 ;
        RECT 75.815 200.345 76.105 200.390 ;
        RECT 77.705 200.345 77.995 200.390 ;
        RECT 68.440 200.190 68.760 200.250 ;
        RECT 69.835 200.190 70.125 200.235 ;
        RECT 68.440 200.050 70.125 200.190 ;
        RECT 68.440 199.990 68.760 200.050 ;
        RECT 69.835 200.005 70.125 200.050 ;
        RECT 78.575 200.190 78.865 200.235 ;
        RECT 84.540 200.190 84.860 200.250 ;
        RECT 78.575 200.050 84.860 200.190 ;
        RECT 78.575 200.005 78.865 200.050 ;
        RECT 84.540 199.990 84.860 200.050 ;
        RECT 69.375 199.850 69.665 199.895 ;
        RECT 70.740 199.850 71.060 199.910 ;
        RECT 65.770 199.710 71.060 199.850 ;
        RECT 65.220 199.650 65.540 199.710 ;
        RECT 69.375 199.665 69.665 199.710 ;
        RECT 70.740 199.650 71.060 199.710 ;
        RECT 52.915 199.510 53.505 199.555 ;
        RECT 56.155 199.510 56.805 199.555 ;
        RECT 52.340 199.370 56.805 199.510 ;
        RECT 52.340 199.310 52.660 199.370 ;
        RECT 52.915 199.325 53.205 199.370 ;
        RECT 56.155 199.325 56.805 199.370 ;
        RECT 58.795 199.510 59.085 199.555 ;
        RECT 58.795 199.370 62.230 199.510 ;
        RECT 58.795 199.325 59.085 199.370 ;
        RECT 51.435 199.170 51.725 199.215 ;
        RECT 55.100 199.170 55.420 199.230 ;
        RECT 62.090 199.215 62.230 199.370 ;
        RECT 67.060 199.310 67.380 199.570 ;
        RECT 51.435 199.030 55.420 199.170 ;
        RECT 51.435 198.985 51.725 199.030 ;
        RECT 55.100 198.970 55.420 199.030 ;
        RECT 62.015 198.985 62.305 199.215 ;
        RECT 64.760 199.170 65.080 199.230 ;
        RECT 66.025 199.170 66.315 199.215 ;
        RECT 64.760 199.030 66.315 199.170 ;
        RECT 64.760 198.970 65.080 199.030 ;
        RECT 66.025 198.985 66.315 199.030 ;
        RECT 68.900 198.970 69.220 199.230 ;
        RECT 70.830 199.170 70.970 199.650 ;
        RECT 71.615 199.555 71.905 199.870 ;
        RECT 72.695 199.850 72.985 199.895 ;
        RECT 76.275 199.850 76.565 199.895 ;
        RECT 78.110 199.850 78.400 199.895 ;
        RECT 79.955 199.850 80.245 199.895 ;
        RECT 85.920 199.850 86.240 199.910 ;
        RECT 72.695 199.710 78.400 199.850 ;
        RECT 72.695 199.665 72.985 199.710 ;
        RECT 76.275 199.665 76.565 199.710 ;
        RECT 78.110 199.665 78.400 199.710 ;
        RECT 79.110 199.710 86.240 199.850 ;
        RECT 71.315 199.510 71.905 199.555 ;
        RECT 73.500 199.510 73.820 199.570 ;
        RECT 74.555 199.510 75.205 199.555 ;
        RECT 71.315 199.370 75.205 199.510 ;
        RECT 71.315 199.325 71.605 199.370 ;
        RECT 73.500 199.310 73.820 199.370 ;
        RECT 74.555 199.325 75.205 199.370 ;
        RECT 76.720 199.510 77.040 199.570 ;
        RECT 77.195 199.510 77.485 199.555 ;
        RECT 76.720 199.370 77.485 199.510 ;
        RECT 76.720 199.310 77.040 199.370 ;
        RECT 77.195 199.325 77.485 199.370 ;
        RECT 79.110 199.170 79.250 199.710 ;
        RECT 79.955 199.665 80.245 199.710 ;
        RECT 85.920 199.650 86.240 199.710 ;
        RECT 70.830 199.030 79.250 199.170 ;
        RECT 79.480 198.970 79.800 199.230 ;
        RECT 15.010 198.350 113.450 198.830 ;
        RECT 62.920 197.950 63.240 198.210 ;
        RECT 63.840 197.950 64.160 198.210 ;
        RECT 64.775 198.150 65.065 198.195 ;
        RECT 65.220 198.150 65.540 198.210 ;
        RECT 64.775 198.010 65.540 198.150 ;
        RECT 64.775 197.965 65.065 198.010 ;
        RECT 65.220 197.950 65.540 198.010 ;
        RECT 53.720 197.810 54.040 197.870 ;
        RECT 54.755 197.810 55.045 197.855 ;
        RECT 57.995 197.810 58.645 197.855 ;
        RECT 53.720 197.670 58.645 197.810 ;
        RECT 53.720 197.610 54.040 197.670 ;
        RECT 54.755 197.625 55.345 197.670 ;
        RECT 57.995 197.625 58.645 197.670 ;
        RECT 55.055 197.310 55.345 197.625 ;
        RECT 60.620 197.610 60.940 197.870 ;
        RECT 63.010 197.810 63.150 197.950 ;
        RECT 66.715 197.810 67.005 197.855 ;
        RECT 68.900 197.810 69.220 197.870 ;
        RECT 79.480 197.855 79.800 197.870 ;
        RECT 69.955 197.810 70.605 197.855 ;
        RECT 63.010 197.670 64.990 197.810 ;
        RECT 56.135 197.470 56.425 197.515 ;
        RECT 59.715 197.470 60.005 197.515 ;
        RECT 61.550 197.470 61.840 197.515 ;
        RECT 56.135 197.330 61.840 197.470 ;
        RECT 56.135 197.285 56.425 197.330 ;
        RECT 59.715 197.285 60.005 197.330 ;
        RECT 61.550 197.285 61.840 197.330 ;
        RECT 62.000 197.270 62.320 197.530 ;
        RECT 62.935 197.285 63.225 197.515 ;
        RECT 51.895 197.130 52.185 197.175 ;
        RECT 63.010 197.130 63.150 197.285 ;
        RECT 63.380 197.270 63.700 197.530 ;
        RECT 64.850 197.515 64.990 197.670 ;
        RECT 66.715 197.670 70.605 197.810 ;
        RECT 66.715 197.625 67.305 197.670 ;
        RECT 64.775 197.285 65.065 197.515 ;
        RECT 67.015 197.310 67.305 197.625 ;
        RECT 68.900 197.610 69.220 197.670 ;
        RECT 69.955 197.625 70.605 197.670 ;
        RECT 76.375 197.810 76.665 197.855 ;
        RECT 79.480 197.810 80.265 197.855 ;
        RECT 76.375 197.670 80.265 197.810 ;
        RECT 76.375 197.625 76.965 197.670 ;
        RECT 68.095 197.470 68.385 197.515 ;
        RECT 71.675 197.470 71.965 197.515 ;
        RECT 73.510 197.470 73.800 197.515 ;
        RECT 68.095 197.330 73.800 197.470 ;
        RECT 68.095 197.285 68.385 197.330 ;
        RECT 71.675 197.285 71.965 197.330 ;
        RECT 73.510 197.285 73.800 197.330 ;
        RECT 76.675 197.310 76.965 197.625 ;
        RECT 79.480 197.625 80.265 197.670 ;
        RECT 79.480 197.610 79.800 197.625 ;
        RECT 82.240 197.610 82.560 197.870 ;
        RECT 77.755 197.470 78.045 197.515 ;
        RECT 81.335 197.470 81.625 197.515 ;
        RECT 83.170 197.470 83.460 197.515 ;
        RECT 77.755 197.330 83.460 197.470 ;
        RECT 77.755 197.285 78.045 197.330 ;
        RECT 81.335 197.285 81.625 197.330 ;
        RECT 83.170 197.285 83.460 197.330 ;
        RECT 64.300 197.130 64.620 197.190 ;
        RECT 51.895 196.990 64.620 197.130 ;
        RECT 64.850 197.130 64.990 197.285 ;
        RECT 70.280 197.130 70.600 197.190 ;
        RECT 64.850 196.990 70.600 197.130 ;
        RECT 51.895 196.945 52.185 196.990 ;
        RECT 64.300 196.930 64.620 196.990 ;
        RECT 70.280 196.930 70.600 196.990 ;
        RECT 72.580 196.930 72.900 197.190 ;
        RECT 73.975 197.130 74.265 197.175 ;
        RECT 83.635 197.130 83.925 197.175 ;
        RECT 84.540 197.130 84.860 197.190 ;
        RECT 86.840 197.130 87.160 197.190 ;
        RECT 73.975 196.990 87.160 197.130 ;
        RECT 73.975 196.945 74.265 196.990 ;
        RECT 83.635 196.945 83.925 196.990 ;
        RECT 84.540 196.930 84.860 196.990 ;
        RECT 86.840 196.930 87.160 196.990 ;
        RECT 95.135 197.130 95.425 197.175 ;
        RECT 95.580 197.130 95.900 197.190 ;
        RECT 95.135 196.990 95.900 197.130 ;
        RECT 95.135 196.945 95.425 196.990 ;
        RECT 95.580 196.930 95.900 196.990 ;
        RECT 56.135 196.790 56.425 196.835 ;
        RECT 59.255 196.790 59.545 196.835 ;
        RECT 61.145 196.790 61.435 196.835 ;
        RECT 56.135 196.650 61.435 196.790 ;
        RECT 56.135 196.605 56.425 196.650 ;
        RECT 59.255 196.605 59.545 196.650 ;
        RECT 61.145 196.605 61.435 196.650 ;
        RECT 63.840 196.790 64.160 196.850 ;
        RECT 68.095 196.790 68.385 196.835 ;
        RECT 71.215 196.790 71.505 196.835 ;
        RECT 73.105 196.790 73.395 196.835 ;
        RECT 63.840 196.650 67.750 196.790 ;
        RECT 63.840 196.590 64.160 196.650 ;
        RECT 65.235 196.450 65.525 196.495 ;
        RECT 65.680 196.450 66.000 196.510 ;
        RECT 65.235 196.310 66.000 196.450 ;
        RECT 67.610 196.450 67.750 196.650 ;
        RECT 68.095 196.650 73.395 196.790 ;
        RECT 68.095 196.605 68.385 196.650 ;
        RECT 71.215 196.605 71.505 196.650 ;
        RECT 73.105 196.605 73.395 196.650 ;
        RECT 77.755 196.790 78.045 196.835 ;
        RECT 80.875 196.790 81.165 196.835 ;
        RECT 82.765 196.790 83.055 196.835 ;
        RECT 77.755 196.650 83.055 196.790 ;
        RECT 77.755 196.605 78.045 196.650 ;
        RECT 80.875 196.605 81.165 196.650 ;
        RECT 82.765 196.605 83.055 196.650 ;
        RECT 69.360 196.450 69.680 196.510 ;
        RECT 67.610 196.310 69.680 196.450 ;
        RECT 65.235 196.265 65.525 196.310 ;
        RECT 65.680 196.250 66.000 196.310 ;
        RECT 69.360 196.250 69.680 196.310 ;
        RECT 72.120 196.450 72.440 196.510 ;
        RECT 74.895 196.450 75.185 196.495 ;
        RECT 72.120 196.310 75.185 196.450 ;
        RECT 72.120 196.250 72.440 196.310 ;
        RECT 74.895 196.265 75.185 196.310 ;
        RECT 97.420 196.450 97.740 196.510 ;
        RECT 97.895 196.450 98.185 196.495 ;
        RECT 97.420 196.310 98.185 196.450 ;
        RECT 97.420 196.250 97.740 196.310 ;
        RECT 97.895 196.265 98.185 196.310 ;
        RECT 15.010 195.630 113.450 196.110 ;
        RECT 52.340 195.230 52.660 195.490 ;
        RECT 53.720 195.230 54.040 195.490 ;
        RECT 55.100 195.430 55.420 195.490 ;
        RECT 57.860 195.430 58.180 195.490 ;
        RECT 55.100 195.290 58.180 195.430 ;
        RECT 55.100 195.230 55.420 195.290 ;
        RECT 57.860 195.230 58.180 195.290 ;
        RECT 61.095 195.430 61.385 195.475 ;
        RECT 61.540 195.430 61.860 195.490 ;
        RECT 63.840 195.430 64.160 195.490 ;
        RECT 61.095 195.290 61.860 195.430 ;
        RECT 61.095 195.245 61.385 195.290 ;
        RECT 61.540 195.230 61.860 195.290 ;
        RECT 62.550 195.290 64.160 195.430 ;
        RECT 62.550 195.090 62.690 195.290 ;
        RECT 54.730 194.950 62.690 195.090 ;
        RECT 54.730 194.455 54.870 194.950 ;
        RECT 56.035 194.750 56.325 194.795 ;
        RECT 62.920 194.750 63.240 194.810 ;
        RECT 63.470 194.795 63.610 195.290 ;
        RECT 63.840 195.230 64.160 195.290 ;
        RECT 64.760 195.230 65.080 195.490 ;
        RECT 66.140 195.430 66.460 195.490 ;
        RECT 68.455 195.430 68.745 195.475 ;
        RECT 66.140 195.290 68.745 195.430 ;
        RECT 66.140 195.230 66.460 195.290 ;
        RECT 68.455 195.245 68.745 195.290 ;
        RECT 72.580 195.430 72.900 195.490 ;
        RECT 75.815 195.430 76.105 195.475 ;
        RECT 72.580 195.290 76.105 195.430 ;
        RECT 72.580 195.230 72.900 195.290 ;
        RECT 75.815 195.245 76.105 195.290 ;
        RECT 76.720 195.430 77.040 195.490 ;
        RECT 78.575 195.430 78.865 195.475 ;
        RECT 76.720 195.290 78.865 195.430 ;
        RECT 76.720 195.230 77.040 195.290 ;
        RECT 78.575 195.245 78.865 195.290 ;
        RECT 80.415 195.430 80.705 195.475 ;
        RECT 82.240 195.430 82.560 195.490 ;
        RECT 80.415 195.290 82.560 195.430 ;
        RECT 80.415 195.245 80.705 195.290 ;
        RECT 82.240 195.230 82.560 195.290 ;
        RECT 97.995 195.090 98.285 195.135 ;
        RECT 101.115 195.090 101.405 195.135 ;
        RECT 103.005 195.090 103.295 195.135 ;
        RECT 70.830 194.950 77.410 195.090 ;
        RECT 56.035 194.610 63.240 194.750 ;
        RECT 56.035 194.565 56.325 194.610 ;
        RECT 62.920 194.550 63.240 194.610 ;
        RECT 63.395 194.565 63.685 194.795 ;
        RECT 63.840 194.750 64.160 194.810 ;
        RECT 67.660 194.750 67.950 194.795 ;
        RECT 68.440 194.750 68.760 194.810 ;
        RECT 70.830 194.750 70.970 194.950 ;
        RECT 63.840 194.610 65.910 194.750 ;
        RECT 63.840 194.550 64.160 194.610 ;
        RECT 52.815 194.410 53.105 194.455 ;
        RECT 53.275 194.410 53.565 194.455 ;
        RECT 52.815 194.270 54.410 194.410 ;
        RECT 52.815 194.225 53.105 194.270 ;
        RECT 53.275 194.225 53.565 194.270 ;
        RECT 54.270 194.070 54.410 194.270 ;
        RECT 54.655 194.225 54.945 194.455 ;
        RECT 57.860 194.410 58.180 194.470 ;
        RECT 60.160 194.410 60.480 194.470 ;
        RECT 57.860 194.270 60.480 194.410 ;
        RECT 57.860 194.210 58.180 194.270 ;
        RECT 60.160 194.210 60.480 194.270 ;
        RECT 62.475 194.410 62.765 194.455 ;
        RECT 64.300 194.410 64.620 194.470 ;
        RECT 65.235 194.410 65.525 194.455 ;
        RECT 62.475 194.270 65.525 194.410 ;
        RECT 65.770 194.410 65.910 194.610 ;
        RECT 67.660 194.610 68.760 194.750 ;
        RECT 67.660 194.565 67.950 194.610 ;
        RECT 68.440 194.550 68.760 194.610 ;
        RECT 68.990 194.610 70.970 194.750 ;
        RECT 66.600 194.410 66.920 194.470 ;
        RECT 68.990 194.410 69.130 194.610 ;
        RECT 72.120 194.550 72.440 194.810 ;
        RECT 73.040 194.750 73.360 194.810 ;
        RECT 76.735 194.750 77.025 194.795 ;
        RECT 73.040 194.610 77.025 194.750 ;
        RECT 73.040 194.550 73.360 194.610 ;
        RECT 76.735 194.565 77.025 194.610 ;
        RECT 65.770 194.270 69.130 194.410 ;
        RECT 62.475 194.225 62.765 194.270 ;
        RECT 64.300 194.210 64.620 194.270 ;
        RECT 65.235 194.225 65.525 194.270 ;
        RECT 66.600 194.210 66.920 194.270 ;
        RECT 69.360 194.210 69.680 194.470 ;
        RECT 70.280 194.210 70.600 194.470 ;
        RECT 72.210 194.410 72.350 194.550 ;
        RECT 77.270 194.455 77.410 194.950 ;
        RECT 93.830 194.950 97.650 195.090 ;
        RECT 77.640 194.750 77.960 194.810 ;
        RECT 93.830 194.750 93.970 194.950 ;
        RECT 77.640 194.610 80.170 194.750 ;
        RECT 77.640 194.550 77.960 194.610 ;
        RECT 80.030 194.455 80.170 194.610 ;
        RECT 86.010 194.610 93.970 194.750 ;
        RECT 86.010 194.470 86.150 194.610 ;
        RECT 70.830 194.270 72.350 194.410 ;
        RECT 56.940 194.070 57.260 194.130 ;
        RECT 54.270 193.930 57.260 194.070 ;
        RECT 56.940 193.870 57.260 193.930 ;
        RECT 67.075 194.070 67.365 194.115 ;
        RECT 68.900 194.070 69.220 194.130 ;
        RECT 70.830 194.070 70.970 194.270 ;
        RECT 77.195 194.225 77.485 194.455 ;
        RECT 79.495 194.410 79.785 194.455 ;
        RECT 77.730 194.270 79.785 194.410 ;
        RECT 67.075 193.930 70.970 194.070 ;
        RECT 72.120 194.070 72.440 194.130 ;
        RECT 77.730 194.070 77.870 194.270 ;
        RECT 79.495 194.225 79.785 194.270 ;
        RECT 79.955 194.225 80.245 194.455 ;
        RECT 85.920 194.210 86.240 194.470 ;
        RECT 86.380 194.210 86.700 194.470 ;
        RECT 88.235 194.225 88.525 194.455 ;
        RECT 91.440 194.410 91.760 194.470 ;
        RECT 93.830 194.455 93.970 194.610 ;
        RECT 95.135 194.750 95.425 194.795 ;
        RECT 95.580 194.750 95.900 194.810 ;
        RECT 95.135 194.610 95.900 194.750 ;
        RECT 97.510 194.750 97.650 194.950 ;
        RECT 97.995 194.950 103.295 195.090 ;
        RECT 97.995 194.905 98.285 194.950 ;
        RECT 101.115 194.905 101.405 194.950 ;
        RECT 103.005 194.905 103.295 194.950 ;
        RECT 100.640 194.750 100.960 194.810 ;
        RECT 97.510 194.610 100.960 194.750 ;
        RECT 95.135 194.565 95.425 194.610 ;
        RECT 95.580 194.550 95.900 194.610 ;
        RECT 100.640 194.550 100.960 194.610 ;
        RECT 91.915 194.410 92.205 194.455 ;
        RECT 91.440 194.270 92.205 194.410 ;
        RECT 88.310 194.070 88.450 194.225 ;
        RECT 91.440 194.210 91.760 194.270 ;
        RECT 91.915 194.225 92.205 194.270 ;
        RECT 93.755 194.225 94.045 194.455 ;
        RECT 94.215 194.410 94.505 194.455 ;
        RECT 96.915 194.410 97.205 194.430 ;
        RECT 94.215 194.270 97.205 194.410 ;
        RECT 94.215 194.225 94.505 194.270 ;
        RECT 96.915 194.115 97.205 194.270 ;
        RECT 97.995 194.410 98.285 194.455 ;
        RECT 101.575 194.410 101.865 194.455 ;
        RECT 103.410 194.410 103.700 194.455 ;
        RECT 97.995 194.270 103.700 194.410 ;
        RECT 97.995 194.225 98.285 194.270 ;
        RECT 101.575 194.225 101.865 194.270 ;
        RECT 103.410 194.225 103.700 194.270 ;
        RECT 103.875 194.410 104.165 194.455 ;
        RECT 104.780 194.410 105.100 194.470 ;
        RECT 103.875 194.270 105.100 194.410 ;
        RECT 103.875 194.225 104.165 194.270 ;
        RECT 104.780 194.210 105.100 194.270 ;
        RECT 72.120 193.930 77.870 194.070 ;
        RECT 86.010 193.930 88.450 194.070 ;
        RECT 96.615 194.070 97.205 194.115 ;
        RECT 99.855 194.070 100.505 194.115 ;
        RECT 96.615 193.930 100.505 194.070 ;
        RECT 67.075 193.885 67.365 193.930 ;
        RECT 68.900 193.870 69.220 193.930 ;
        RECT 72.120 193.870 72.440 193.930 ;
        RECT 86.010 193.790 86.150 193.930 ;
        RECT 96.615 193.885 96.905 193.930 ;
        RECT 99.855 193.885 100.505 193.930 ;
        RECT 102.480 193.870 102.800 194.130 ;
        RECT 57.400 193.530 57.720 193.790 ;
        RECT 65.680 193.730 66.000 193.790 ;
        RECT 66.615 193.730 66.905 193.775 ;
        RECT 65.680 193.590 66.905 193.730 ;
        RECT 65.680 193.530 66.000 193.590 ;
        RECT 66.615 193.545 66.905 193.590 ;
        RECT 71.200 193.530 71.520 193.790 ;
        RECT 74.895 193.730 75.185 193.775 ;
        RECT 75.800 193.730 76.120 193.790 ;
        RECT 74.895 193.590 76.120 193.730 ;
        RECT 74.895 193.545 75.185 193.590 ;
        RECT 75.800 193.530 76.120 193.590 ;
        RECT 85.920 193.530 86.240 193.790 ;
        RECT 89.140 193.730 89.460 193.790 ;
        RECT 91.455 193.730 91.745 193.775 ;
        RECT 89.140 193.590 91.745 193.730 ;
        RECT 89.140 193.530 89.460 193.590 ;
        RECT 91.455 193.545 91.745 193.590 ;
        RECT 91.900 193.730 92.220 193.790 ;
        RECT 92.835 193.730 93.125 193.775 ;
        RECT 91.900 193.590 93.125 193.730 ;
        RECT 91.900 193.530 92.220 193.590 ;
        RECT 92.835 193.545 93.125 193.590 ;
        RECT 15.010 192.910 113.450 193.390 ;
        RECT 65.235 192.710 65.525 192.755 ;
        RECT 67.060 192.710 67.380 192.770 ;
        RECT 65.235 192.570 68.210 192.710 ;
        RECT 65.235 192.525 65.525 192.570 ;
        RECT 67.060 192.510 67.380 192.570 ;
        RECT 65.680 192.370 66.000 192.430 ;
        RECT 62.090 192.230 66.000 192.370 ;
        RECT 44.520 192.030 44.840 192.090 ;
        RECT 62.090 192.075 62.230 192.230 ;
        RECT 65.680 192.170 66.000 192.230 ;
        RECT 66.155 192.185 66.445 192.415 ;
        RECT 68.070 192.370 68.210 192.570 ;
        RECT 68.440 192.510 68.760 192.770 ;
        RECT 68.900 192.510 69.220 192.770 ;
        RECT 71.295 192.710 71.585 192.755 ;
        RECT 69.450 192.570 71.585 192.710 ;
        RECT 69.450 192.370 69.590 192.570 ;
        RECT 71.295 192.525 71.585 192.570 ;
        RECT 72.120 192.510 72.440 192.770 ;
        RECT 73.040 192.510 73.360 192.770 ;
        RECT 89.140 192.710 89.460 192.770 ;
        RECT 97.895 192.710 98.185 192.755 ;
        RECT 89.140 192.570 98.185 192.710 ;
        RECT 89.140 192.510 89.460 192.570 ;
        RECT 97.895 192.525 98.185 192.570 ;
        RECT 68.070 192.230 69.590 192.370 ;
        RECT 70.295 192.370 70.585 192.415 ;
        RECT 73.130 192.370 73.270 192.510 ;
        RECT 70.295 192.230 73.270 192.370 ;
        RECT 70.295 192.185 70.585 192.230 ;
        RECT 48.215 192.030 48.505 192.075 ;
        RECT 44.520 191.890 48.505 192.030 ;
        RECT 44.520 191.830 44.840 191.890 ;
        RECT 48.215 191.845 48.505 191.890 ;
        RECT 62.015 191.845 62.305 192.075 ;
        RECT 62.475 192.030 62.765 192.075 ;
        RECT 64.760 192.030 65.080 192.090 ;
        RECT 66.230 192.030 66.370 192.185 ;
        RECT 75.800 192.170 76.120 192.430 ;
        RECT 86.380 192.370 86.700 192.430 ;
        RECT 87.415 192.370 87.705 192.415 ;
        RECT 90.655 192.370 91.305 192.415 ;
        RECT 86.380 192.230 91.305 192.370 ;
        RECT 86.380 192.170 86.700 192.230 ;
        RECT 87.415 192.185 88.005 192.230 ;
        RECT 90.655 192.185 91.305 192.230 ;
        RECT 91.900 192.370 92.220 192.430 ;
        RECT 105.700 192.415 106.020 192.430 ;
        RECT 93.295 192.370 93.585 192.415 ;
        RECT 91.900 192.230 93.585 192.370 ;
        RECT 62.475 191.890 66.370 192.030 ;
        RECT 70.740 192.030 71.060 192.090 ;
        RECT 72.595 192.030 72.885 192.075 ;
        RECT 70.740 191.890 72.885 192.030 ;
        RECT 62.475 191.845 62.765 191.890 ;
        RECT 64.760 191.830 65.080 191.890 ;
        RECT 70.740 191.830 71.060 191.890 ;
        RECT 72.595 191.845 72.885 191.890 ;
        RECT 73.515 191.845 73.805 192.075 ;
        RECT 81.320 192.030 81.640 192.090 ;
        RECT 84.555 192.030 84.845 192.075 ;
        RECT 81.320 191.890 84.845 192.030 ;
        RECT 41.760 191.490 42.080 191.750 ;
        RECT 57.400 191.690 57.720 191.750 ;
        RECT 63.855 191.690 64.145 191.735 ;
        RECT 57.400 191.550 64.145 191.690 ;
        RECT 57.400 191.490 57.720 191.550 ;
        RECT 63.855 191.505 64.145 191.550 ;
        RECT 69.360 191.690 69.680 191.750 ;
        RECT 73.590 191.690 73.730 191.845 ;
        RECT 81.320 191.830 81.640 191.890 ;
        RECT 84.555 191.845 84.845 191.890 ;
        RECT 87.715 191.870 88.005 192.185 ;
        RECT 91.900 192.170 92.220 192.230 ;
        RECT 93.295 192.185 93.585 192.230 ;
        RECT 102.135 192.370 102.425 192.415 ;
        RECT 105.375 192.370 106.025 192.415 ;
        RECT 102.135 192.230 106.025 192.370 ;
        RECT 102.135 192.185 102.725 192.230 ;
        RECT 105.375 192.185 106.025 192.230 ;
        RECT 88.795 192.030 89.085 192.075 ;
        RECT 92.375 192.030 92.665 192.075 ;
        RECT 94.210 192.030 94.500 192.075 ;
        RECT 88.795 191.890 94.500 192.030 ;
        RECT 88.795 191.845 89.085 191.890 ;
        RECT 92.375 191.845 92.665 191.890 ;
        RECT 94.210 191.845 94.500 191.890 ;
        RECT 94.675 192.030 94.965 192.075 ;
        RECT 94.675 191.890 99.950 192.030 ;
        RECT 94.675 191.845 94.965 191.890 ;
        RECT 76.735 191.690 77.025 191.735 ;
        RECT 77.640 191.690 77.960 191.750 ;
        RECT 69.360 191.550 77.960 191.690 ;
        RECT 69.360 191.490 69.680 191.550 ;
        RECT 76.735 191.505 77.025 191.550 ;
        RECT 77.640 191.490 77.960 191.550 ;
        RECT 96.500 191.490 96.820 191.750 ;
        RECT 97.420 191.490 97.740 191.750 ;
        RECT 99.810 191.690 99.950 191.890 ;
        RECT 102.435 191.870 102.725 192.185 ;
        RECT 105.700 192.170 106.020 192.185 ;
        RECT 103.515 192.030 103.805 192.075 ;
        RECT 107.095 192.030 107.385 192.075 ;
        RECT 108.930 192.030 109.220 192.075 ;
        RECT 103.515 191.890 109.220 192.030 ;
        RECT 103.515 191.845 103.805 191.890 ;
        RECT 107.095 191.845 107.385 191.890 ;
        RECT 108.930 191.845 109.220 191.890 ;
        RECT 109.395 191.690 109.685 191.735 ;
        RECT 111.220 191.690 111.540 191.750 ;
        RECT 99.810 191.550 111.540 191.690 ;
        RECT 109.395 191.505 109.685 191.550 ;
        RECT 111.220 191.490 111.540 191.550 ;
        RECT 66.155 191.350 66.445 191.395 ;
        RECT 66.600 191.350 66.920 191.410 ;
        RECT 64.390 191.210 66.920 191.350 ;
        RECT 44.980 190.810 45.300 191.070 ;
        RECT 46.360 191.010 46.680 191.070 ;
        RECT 47.755 191.010 48.045 191.055 ;
        RECT 46.360 190.870 48.045 191.010 ;
        RECT 46.360 190.810 46.680 190.870 ;
        RECT 47.755 190.825 48.045 190.870 ;
        RECT 61.095 191.010 61.385 191.055 ;
        RECT 61.540 191.010 61.860 191.070 ;
        RECT 64.390 191.055 64.530 191.210 ;
        RECT 66.155 191.165 66.445 191.210 ;
        RECT 66.600 191.150 66.920 191.210 ;
        RECT 88.795 191.350 89.085 191.395 ;
        RECT 91.915 191.350 92.205 191.395 ;
        RECT 93.805 191.350 94.095 191.395 ;
        RECT 88.795 191.210 94.095 191.350 ;
        RECT 88.795 191.165 89.085 191.210 ;
        RECT 91.915 191.165 92.205 191.210 ;
        RECT 93.805 191.165 94.095 191.210 ;
        RECT 103.515 191.350 103.805 191.395 ;
        RECT 106.635 191.350 106.925 191.395 ;
        RECT 108.525 191.350 108.815 191.395 ;
        RECT 103.515 191.210 108.815 191.350 ;
        RECT 103.515 191.165 103.805 191.210 ;
        RECT 106.635 191.165 106.925 191.210 ;
        RECT 108.525 191.165 108.815 191.210 ;
        RECT 64.315 191.010 64.605 191.055 ;
        RECT 61.095 190.870 64.605 191.010 ;
        RECT 61.095 190.825 61.385 190.870 ;
        RECT 61.540 190.810 61.860 190.870 ;
        RECT 64.315 190.825 64.605 190.870 ;
        RECT 69.820 190.810 70.140 191.070 ;
        RECT 71.200 190.810 71.520 191.070 ;
        RECT 85.460 190.810 85.780 191.070 ;
        RECT 85.920 190.810 86.240 191.070 ;
        RECT 99.720 190.810 100.040 191.070 ;
        RECT 100.655 191.010 100.945 191.055 ;
        RECT 105.240 191.010 105.560 191.070 ;
        RECT 100.655 190.870 105.560 191.010 ;
        RECT 100.655 190.825 100.945 190.870 ;
        RECT 105.240 190.810 105.560 190.870 ;
        RECT 107.080 191.010 107.400 191.070 ;
        RECT 108.080 191.010 108.370 191.055 ;
        RECT 107.080 190.870 108.370 191.010 ;
        RECT 107.080 190.810 107.400 190.870 ;
        RECT 108.080 190.825 108.370 190.870 ;
        RECT 15.010 190.190 113.450 190.670 ;
        RECT 38.540 189.990 38.860 190.050 ;
        RECT 41.760 189.990 42.080 190.050 ;
        RECT 44.075 189.990 44.365 190.035 ;
        RECT 38.540 189.850 44.365 189.990 ;
        RECT 38.540 189.790 38.860 189.850 ;
        RECT 41.760 189.790 42.080 189.850 ;
        RECT 44.075 189.805 44.365 189.850 ;
        RECT 65.220 189.990 65.540 190.050 ;
        RECT 67.075 189.990 67.365 190.035 ;
        RECT 70.280 189.990 70.600 190.050 ;
        RECT 65.220 189.850 70.600 189.990 ;
        RECT 65.220 189.790 65.540 189.850 ;
        RECT 67.075 189.805 67.365 189.850 ;
        RECT 70.280 189.790 70.600 189.850 ;
        RECT 91.440 189.790 91.760 190.050 ;
        RECT 98.815 189.990 99.105 190.035 ;
        RECT 102.480 189.990 102.800 190.050 ;
        RECT 98.815 189.850 102.800 189.990 ;
        RECT 98.815 189.805 99.105 189.850 ;
        RECT 102.480 189.790 102.800 189.850 ;
        RECT 105.700 189.990 106.020 190.050 ;
        RECT 107.555 189.990 107.845 190.035 ;
        RECT 105.700 189.850 107.845 189.990 ;
        RECT 105.700 189.790 106.020 189.850 ;
        RECT 107.555 189.805 107.845 189.850 ;
        RECT 46.935 189.650 47.225 189.695 ;
        RECT 50.055 189.650 50.345 189.695 ;
        RECT 51.945 189.650 52.235 189.695 ;
        RECT 46.935 189.510 52.235 189.650 ;
        RECT 46.935 189.465 47.225 189.510 ;
        RECT 50.055 189.465 50.345 189.510 ;
        RECT 51.945 189.465 52.235 189.510 ;
        RECT 81.750 189.650 82.040 189.695 ;
        RECT 84.530 189.650 84.820 189.695 ;
        RECT 86.390 189.650 86.680 189.695 ;
        RECT 81.750 189.510 86.680 189.650 ;
        RECT 81.750 189.465 82.040 189.510 ;
        RECT 84.530 189.465 84.820 189.510 ;
        RECT 86.390 189.465 86.680 189.510 ;
        RECT 96.500 189.650 96.820 189.710 ;
        RECT 107.080 189.650 107.400 189.710 ;
        RECT 108.475 189.650 108.765 189.695 ;
        RECT 96.500 189.510 100.410 189.650 ;
        RECT 96.500 189.450 96.820 189.510 ;
        RECT 40.855 189.310 41.145 189.355 ;
        RECT 43.600 189.310 43.920 189.370 ;
        RECT 40.855 189.170 43.920 189.310 ;
        RECT 40.855 189.125 41.145 189.170 ;
        RECT 43.600 189.110 43.920 189.170 ;
        RECT 44.060 189.310 44.380 189.370 ;
        RECT 51.435 189.310 51.725 189.355 ;
        RECT 44.060 189.170 51.725 189.310 ;
        RECT 44.060 189.110 44.380 189.170 ;
        RECT 51.435 189.125 51.725 189.170 ;
        RECT 52.800 189.310 53.120 189.370 ;
        RECT 62.000 189.310 62.320 189.370 ;
        RECT 52.800 189.170 62.320 189.310 ;
        RECT 52.800 189.110 53.120 189.170 ;
        RECT 62.000 189.110 62.320 189.170 ;
        RECT 85.015 189.310 85.305 189.355 ;
        RECT 85.460 189.310 85.780 189.370 ;
        RECT 85.015 189.170 85.780 189.310 ;
        RECT 85.015 189.125 85.305 189.170 ;
        RECT 85.460 189.110 85.780 189.170 ;
        RECT 88.220 189.110 88.540 189.370 ;
        RECT 89.140 189.110 89.460 189.370 ;
        RECT 100.270 189.355 100.410 189.510 ;
        RECT 107.080 189.510 108.765 189.650 ;
        RECT 107.080 189.450 107.400 189.510 ;
        RECT 108.475 189.465 108.765 189.510 ;
        RECT 100.195 189.125 100.485 189.355 ;
        RECT 34.415 188.970 34.705 189.015 ;
        RECT 34.860 188.970 35.180 189.030 ;
        RECT 34.415 188.830 35.180 188.970 ;
        RECT 34.415 188.785 34.705 188.830 ;
        RECT 34.860 188.770 35.180 188.830 ;
        RECT 38.555 188.785 38.845 189.015 ;
        RECT 32.100 188.630 32.420 188.690 ;
        RECT 38.630 188.630 38.770 188.785 ;
        RECT 32.100 188.490 38.770 188.630 ;
        RECT 41.315 188.630 41.605 188.675 ;
        RECT 44.980 188.630 45.300 188.690 ;
        RECT 45.855 188.675 46.145 188.990 ;
        RECT 46.935 188.970 47.225 189.015 ;
        RECT 50.515 188.970 50.805 189.015 ;
        RECT 52.350 188.970 52.640 189.015 ;
        RECT 46.935 188.830 52.640 188.970 ;
        RECT 46.935 188.785 47.225 188.830 ;
        RECT 50.515 188.785 50.805 188.830 ;
        RECT 52.350 188.785 52.640 188.830 ;
        RECT 54.655 188.970 54.945 189.015 ;
        RECT 56.020 188.970 56.340 189.030 ;
        RECT 54.655 188.830 56.340 188.970 ;
        RECT 54.655 188.785 54.945 188.830 ;
        RECT 56.020 188.770 56.340 188.830 ;
        RECT 67.535 188.970 67.825 189.015 ;
        RECT 68.440 188.970 68.760 189.030 ;
        RECT 67.535 188.830 68.760 188.970 ;
        RECT 67.535 188.785 67.825 188.830 ;
        RECT 68.440 188.770 68.760 188.830 ;
        RECT 81.750 188.970 82.040 189.015 ;
        RECT 81.750 188.830 84.285 188.970 ;
        RECT 81.750 188.785 82.040 188.830 ;
        RECT 41.315 188.490 45.300 188.630 ;
        RECT 32.100 188.430 32.420 188.490 ;
        RECT 41.315 188.445 41.605 188.490 ;
        RECT 44.980 188.430 45.300 188.490 ;
        RECT 45.555 188.630 46.145 188.675 ;
        RECT 46.360 188.630 46.680 188.690 ;
        RECT 83.160 188.675 83.480 188.690 ;
        RECT 48.795 188.630 49.445 188.675 ;
        RECT 45.555 188.490 49.445 188.630 ;
        RECT 45.555 188.445 45.845 188.490 ;
        RECT 46.360 188.430 46.680 188.490 ;
        RECT 48.795 188.445 49.445 188.490 ;
        RECT 79.890 188.630 80.180 188.675 ;
        RECT 83.150 188.630 83.480 188.675 ;
        RECT 79.890 188.490 83.480 188.630 ;
        RECT 79.890 188.445 80.180 188.490 ;
        RECT 83.150 188.445 83.480 188.490 ;
        RECT 84.070 188.675 84.285 188.830 ;
        RECT 86.840 188.770 87.160 189.030 ;
        RECT 96.040 188.970 96.360 189.030 ;
        RECT 96.515 188.970 96.805 189.015 ;
        RECT 96.040 188.830 96.805 188.970 ;
        RECT 96.040 188.770 96.360 188.830 ;
        RECT 96.515 188.785 96.805 188.830 ;
        RECT 97.895 188.970 98.185 189.015 ;
        RECT 99.720 188.970 100.040 189.030 ;
        RECT 97.895 188.830 100.040 188.970 ;
        RECT 97.895 188.785 98.185 188.830 ;
        RECT 99.720 188.770 100.040 188.830 ;
        RECT 105.240 188.970 105.560 189.030 ;
        RECT 106.175 188.970 106.465 189.015 ;
        RECT 105.240 188.830 106.465 188.970 ;
        RECT 105.240 188.770 105.560 188.830 ;
        RECT 106.175 188.785 106.465 188.830 ;
        RECT 108.000 188.770 108.320 189.030 ;
        RECT 109.395 188.785 109.685 189.015 ;
        RECT 84.070 188.630 84.360 188.675 ;
        RECT 85.930 188.630 86.220 188.675 ;
        RECT 84.070 188.490 86.220 188.630 ;
        RECT 84.070 188.445 84.360 188.490 ;
        RECT 85.930 188.445 86.220 188.490 ;
        RECT 100.655 188.630 100.945 188.675 ;
        RECT 103.400 188.630 103.720 188.690 ;
        RECT 109.470 188.630 109.610 188.785 ;
        RECT 100.655 188.490 103.720 188.630 ;
        RECT 100.655 188.445 100.945 188.490 ;
        RECT 83.160 188.430 83.480 188.445 ;
        RECT 103.400 188.430 103.720 188.490 ;
        RECT 105.100 188.490 109.610 188.630 ;
        RECT 34.875 188.290 35.165 188.335 ;
        RECT 35.780 188.290 36.100 188.350 ;
        RECT 34.875 188.150 36.100 188.290 ;
        RECT 34.875 188.105 35.165 188.150 ;
        RECT 35.780 188.090 36.100 188.150 ;
        RECT 39.475 188.290 39.765 188.335 ;
        RECT 39.920 188.290 40.240 188.350 ;
        RECT 39.475 188.150 40.240 188.290 ;
        RECT 39.475 188.105 39.765 188.150 ;
        RECT 39.920 188.090 40.240 188.150 ;
        RECT 41.760 188.090 42.080 188.350 ;
        RECT 43.140 188.290 43.460 188.350 ;
        RECT 43.615 188.290 43.905 188.335 ;
        RECT 43.140 188.150 43.905 188.290 ;
        RECT 43.140 188.090 43.460 188.150 ;
        RECT 43.615 188.105 43.905 188.150 ;
        RECT 55.560 188.090 55.880 188.350 ;
        RECT 77.885 188.290 78.175 188.335 ;
        RECT 79.020 188.290 79.340 188.350 ;
        RECT 89.615 188.290 89.905 188.335 ;
        RECT 77.885 188.150 89.905 188.290 ;
        RECT 77.885 188.105 78.175 188.150 ;
        RECT 79.020 188.090 79.340 188.150 ;
        RECT 89.615 188.105 89.905 188.150 ;
        RECT 93.755 188.290 94.045 188.335 ;
        RECT 95.120 188.290 95.440 188.350 ;
        RECT 93.755 188.150 95.440 188.290 ;
        RECT 93.755 188.105 94.045 188.150 ;
        RECT 95.120 188.090 95.440 188.150 ;
        RECT 97.420 188.290 97.740 188.350 ;
        RECT 101.115 188.290 101.405 188.335 ;
        RECT 97.420 188.150 101.405 188.290 ;
        RECT 97.420 188.090 97.740 188.150 ;
        RECT 101.115 188.105 101.405 188.150 ;
        RECT 102.955 188.290 103.245 188.335 ;
        RECT 105.100 188.290 105.240 188.490 ;
        RECT 102.955 188.150 105.240 188.290 ;
        RECT 102.955 188.105 103.245 188.150 ;
        RECT 15.010 187.470 113.450 187.950 ;
        RECT 32.100 187.070 32.420 187.330 ;
        RECT 43.600 187.270 43.920 187.330 ;
        RECT 34.490 187.130 43.920 187.270 ;
        RECT 27.975 186.930 28.265 186.975 ;
        RECT 30.275 186.930 30.565 186.975 ;
        RECT 34.490 186.930 34.630 187.130 ;
        RECT 43.600 187.070 43.920 187.130 ;
        RECT 44.060 187.070 44.380 187.330 ;
        RECT 64.760 187.070 65.080 187.330 ;
        RECT 81.320 187.070 81.640 187.330 ;
        RECT 88.220 187.270 88.540 187.330 ;
        RECT 96.500 187.270 96.820 187.330 ;
        RECT 88.220 187.130 96.820 187.270 ;
        RECT 88.220 187.070 88.540 187.130 ;
        RECT 96.500 187.070 96.820 187.130 ;
        RECT 100.640 187.270 100.960 187.330 ;
        RECT 108.000 187.270 108.320 187.330 ;
        RECT 110.300 187.270 110.620 187.330 ;
        RECT 100.640 187.130 110.620 187.270 ;
        RECT 100.640 187.070 100.960 187.130 ;
        RECT 108.000 187.070 108.320 187.130 ;
        RECT 110.300 187.070 110.620 187.130 ;
        RECT 27.975 186.790 30.565 186.930 ;
        RECT 27.975 186.745 28.265 186.790 ;
        RECT 30.275 186.745 30.565 186.790 ;
        RECT 31.270 186.790 34.630 186.930 ;
        RECT 34.810 186.930 35.100 186.975 ;
        RECT 35.780 186.930 36.100 186.990 ;
        RECT 38.070 186.930 38.360 186.975 ;
        RECT 34.810 186.790 38.360 186.930 ;
        RECT 31.270 186.650 31.410 186.790 ;
        RECT 34.810 186.745 35.100 186.790 ;
        RECT 35.780 186.730 36.100 186.790 ;
        RECT 38.070 186.745 38.360 186.790 ;
        RECT 38.990 186.930 39.280 186.975 ;
        RECT 40.850 186.930 41.140 186.975 ;
        RECT 38.990 186.790 41.140 186.930 ;
        RECT 38.990 186.745 39.280 186.790 ;
        RECT 40.850 186.745 41.140 186.790 ;
        RECT 21.060 186.590 21.380 186.650 ;
        RECT 21.535 186.590 21.825 186.635 ;
        RECT 21.060 186.450 21.825 186.590 ;
        RECT 21.060 186.390 21.380 186.450 ;
        RECT 21.535 186.405 21.825 186.450 ;
        RECT 23.360 186.390 23.680 186.650 ;
        RECT 31.180 186.590 31.500 186.650 ;
        RECT 29.430 186.450 31.500 186.590 ;
        RECT 24.740 186.050 25.060 186.310 ;
        RECT 29.430 186.295 29.570 186.450 ;
        RECT 31.180 186.390 31.500 186.450 ;
        RECT 36.670 186.590 36.960 186.635 ;
        RECT 38.990 186.590 39.205 186.745 ;
        RECT 36.670 186.450 39.205 186.590 ;
        RECT 36.670 186.405 36.960 186.450 ;
        RECT 39.920 186.390 40.240 186.650 ;
        RECT 43.140 186.390 43.460 186.650 ;
        RECT 29.355 186.065 29.645 186.295 ;
        RECT 29.815 186.065 30.105 186.295 ;
        RECT 35.320 186.250 35.640 186.310 ;
        RECT 41.775 186.250 42.065 186.295 ;
        RECT 35.320 186.110 42.065 186.250 ;
        RECT 43.690 186.250 43.830 187.070 ;
        RECT 44.980 186.930 45.300 186.990 ;
        RECT 54.640 186.975 54.960 186.990 ;
        RECT 46.375 186.930 46.665 186.975 ;
        RECT 44.980 186.790 46.665 186.930 ;
        RECT 44.980 186.730 45.300 186.790 ;
        RECT 46.375 186.745 46.665 186.790 ;
        RECT 51.075 186.930 51.365 186.975 ;
        RECT 54.315 186.930 54.965 186.975 ;
        RECT 51.075 186.790 54.965 186.930 ;
        RECT 51.075 186.745 51.665 186.790 ;
        RECT 54.315 186.745 54.965 186.790 ;
        RECT 55.560 186.930 55.880 186.990 ;
        RECT 56.955 186.930 57.245 186.975 ;
        RECT 64.850 186.930 64.990 187.070 ;
        RECT 55.560 186.790 57.245 186.930 ;
        RECT 51.375 186.430 51.665 186.745 ;
        RECT 54.640 186.730 54.960 186.745 ;
        RECT 55.560 186.730 55.880 186.790 ;
        RECT 56.955 186.745 57.245 186.790 ;
        RECT 63.930 186.790 64.990 186.930 ;
        RECT 74.420 186.930 74.740 186.990 ;
        RECT 79.495 186.930 79.785 186.975 ;
        RECT 74.420 186.790 79.785 186.930 ;
        RECT 52.455 186.590 52.745 186.635 ;
        RECT 56.035 186.590 56.325 186.635 ;
        RECT 57.870 186.590 58.160 186.635 ;
        RECT 52.455 186.450 58.160 186.590 ;
        RECT 52.455 186.405 52.745 186.450 ;
        RECT 56.035 186.405 56.325 186.450 ;
        RECT 57.870 186.405 58.160 186.450 ;
        RECT 58.320 186.590 58.640 186.650 ;
        RECT 62.000 186.590 62.320 186.650 ;
        RECT 63.930 186.635 64.070 186.790 ;
        RECT 74.420 186.730 74.740 186.790 ;
        RECT 79.495 186.745 79.785 186.790 ;
        RECT 83.160 186.930 83.480 186.990 ;
        RECT 106.620 186.975 106.940 186.990 ;
        RECT 87.775 186.930 88.065 186.975 ;
        RECT 83.160 186.790 88.065 186.930 ;
        RECT 83.160 186.730 83.480 186.790 ;
        RECT 87.775 186.745 88.065 186.790 ;
        RECT 103.515 186.930 103.805 186.975 ;
        RECT 106.620 186.930 107.405 186.975 ;
        RECT 103.515 186.790 107.405 186.930 ;
        RECT 103.515 186.745 104.105 186.790 ;
        RECT 58.320 186.450 62.320 186.590 ;
        RECT 58.320 186.390 58.640 186.450 ;
        RECT 62.000 186.390 62.320 186.450 ;
        RECT 63.855 186.405 64.145 186.635 ;
        RECT 65.220 186.390 65.540 186.650 ;
        RECT 76.260 186.390 76.580 186.650 ;
        RECT 82.715 186.590 83.005 186.635 ;
        RECT 78.190 186.450 83.005 186.590 ;
        RECT 44.060 186.250 44.380 186.310 ;
        RECT 44.995 186.250 45.285 186.295 ;
        RECT 43.690 186.110 45.285 186.250 ;
        RECT 21.995 185.910 22.285 185.955 ;
        RECT 25.200 185.910 25.520 185.970 ;
        RECT 21.995 185.770 25.520 185.910 ;
        RECT 21.995 185.725 22.285 185.770 ;
        RECT 25.200 185.710 25.520 185.770 ;
        RECT 24.295 185.570 24.585 185.615 ;
        RECT 25.660 185.570 25.980 185.630 ;
        RECT 24.295 185.430 25.980 185.570 ;
        RECT 29.890 185.570 30.030 186.065 ;
        RECT 35.320 186.050 35.640 186.110 ;
        RECT 41.775 186.065 42.065 186.110 ;
        RECT 44.060 186.050 44.380 186.110 ;
        RECT 44.995 186.065 45.285 186.110 ;
        RECT 45.915 186.065 46.205 186.295 ;
        RECT 61.540 186.250 61.860 186.310 ;
        RECT 64.315 186.250 64.605 186.295 ;
        RECT 61.540 186.110 64.605 186.250 ;
        RECT 36.670 185.910 36.960 185.955 ;
        RECT 39.450 185.910 39.740 185.955 ;
        RECT 41.310 185.910 41.600 185.955 ;
        RECT 36.670 185.770 41.600 185.910 ;
        RECT 36.670 185.725 36.960 185.770 ;
        RECT 39.450 185.725 39.740 185.770 ;
        RECT 41.310 185.725 41.600 185.770 ;
        RECT 43.140 185.910 43.460 185.970 ;
        RECT 45.990 185.910 46.130 186.065 ;
        RECT 61.540 186.050 61.860 186.110 ;
        RECT 64.315 186.065 64.605 186.110 ;
        RECT 64.775 186.250 65.065 186.295 ;
        RECT 65.680 186.250 66.000 186.310 ;
        RECT 69.360 186.250 69.680 186.310 ;
        RECT 64.775 186.110 69.680 186.250 ;
        RECT 64.775 186.065 65.065 186.110 ;
        RECT 65.680 186.050 66.000 186.110 ;
        RECT 69.360 186.050 69.680 186.110 ;
        RECT 73.960 186.250 74.280 186.310 ;
        RECT 78.190 186.250 78.330 186.450 ;
        RECT 82.715 186.405 83.005 186.450 ;
        RECT 87.300 186.590 87.620 186.650 ;
        RECT 88.235 186.590 88.525 186.635 ;
        RECT 95.120 186.590 95.440 186.650 ;
        RECT 97.420 186.590 97.740 186.650 ;
        RECT 87.300 186.450 88.525 186.590 ;
        RECT 87.300 186.390 87.620 186.450 ;
        RECT 88.235 186.405 88.525 186.450 ;
        RECT 89.690 186.450 90.750 186.590 ;
        RECT 73.960 186.110 78.330 186.250 ;
        RECT 73.960 186.050 74.280 186.110 ;
        RECT 78.575 186.065 78.865 186.295 ;
        RECT 79.035 186.250 79.325 186.295 ;
        RECT 79.480 186.250 79.800 186.310 ;
        RECT 79.035 186.110 79.800 186.250 ;
        RECT 79.035 186.065 79.325 186.110 ;
        RECT 49.580 185.910 49.900 185.970 ;
        RECT 43.140 185.770 49.900 185.910 ;
        RECT 43.140 185.710 43.460 185.770 ;
        RECT 49.580 185.710 49.900 185.770 ;
        RECT 52.455 185.910 52.745 185.955 ;
        RECT 55.575 185.910 55.865 185.955 ;
        RECT 57.465 185.910 57.755 185.955 ;
        RECT 52.455 185.770 57.755 185.910 ;
        RECT 52.455 185.725 52.745 185.770 ;
        RECT 55.575 185.725 55.865 185.770 ;
        RECT 57.465 185.725 57.755 185.770 ;
        RECT 75.340 185.910 75.660 185.970 ;
        RECT 78.650 185.910 78.790 186.065 ;
        RECT 79.480 186.050 79.800 186.110 ;
        RECT 86.855 186.250 87.145 186.295 ;
        RECT 89.690 186.250 89.830 186.450 ;
        RECT 90.610 186.310 90.750 186.450 ;
        RECT 95.120 186.450 97.740 186.590 ;
        RECT 95.120 186.390 95.440 186.450 ;
        RECT 97.420 186.390 97.740 186.450 ;
        RECT 100.640 186.390 100.960 186.650 ;
        RECT 103.815 186.430 104.105 186.745 ;
        RECT 106.620 186.745 107.405 186.790 ;
        RECT 109.395 186.930 109.685 186.975 ;
        RECT 109.840 186.930 110.160 186.990 ;
        RECT 109.395 186.790 110.160 186.930 ;
        RECT 109.395 186.745 109.685 186.790 ;
        RECT 106.620 186.730 106.940 186.745 ;
        RECT 109.840 186.730 110.160 186.790 ;
        RECT 104.895 186.590 105.185 186.635 ;
        RECT 108.475 186.590 108.765 186.635 ;
        RECT 110.310 186.590 110.600 186.635 ;
        RECT 104.895 186.450 110.600 186.590 ;
        RECT 104.895 186.405 105.185 186.450 ;
        RECT 108.475 186.405 108.765 186.450 ;
        RECT 110.310 186.405 110.600 186.450 ;
        RECT 86.855 186.110 89.830 186.250 ;
        RECT 86.855 186.065 87.145 186.110 ;
        RECT 90.075 186.065 90.365 186.295 ;
        RECT 90.520 186.250 90.840 186.310 ;
        RECT 95.595 186.250 95.885 186.295 ;
        RECT 90.520 186.110 95.885 186.250 ;
        RECT 75.340 185.770 78.790 185.910 ;
        RECT 90.150 185.910 90.290 186.065 ;
        RECT 90.520 186.050 90.840 186.110 ;
        RECT 95.595 186.065 95.885 186.110 ;
        RECT 96.500 186.050 96.820 186.310 ;
        RECT 110.760 186.050 111.080 186.310 ;
        RECT 93.295 185.910 93.585 185.955 ;
        RECT 90.150 185.770 93.585 185.910 ;
        RECT 75.340 185.710 75.660 185.770 ;
        RECT 93.295 185.725 93.585 185.770 ;
        RECT 104.895 185.910 105.185 185.955 ;
        RECT 108.015 185.910 108.305 185.955 ;
        RECT 109.905 185.910 110.195 185.955 ;
        RECT 104.895 185.770 110.195 185.910 ;
        RECT 104.895 185.725 105.185 185.770 ;
        RECT 108.015 185.725 108.305 185.770 ;
        RECT 109.905 185.725 110.195 185.770 ;
        RECT 32.805 185.570 33.095 185.615 ;
        RECT 36.240 185.570 36.560 185.630 ;
        RECT 41.760 185.570 42.080 185.630 ;
        RECT 29.890 185.430 42.080 185.570 ;
        RECT 24.295 185.385 24.585 185.430 ;
        RECT 25.660 185.370 25.980 185.430 ;
        RECT 32.805 185.385 33.095 185.430 ;
        RECT 36.240 185.370 36.560 185.430 ;
        RECT 41.760 185.370 42.080 185.430 ;
        RECT 48.215 185.570 48.505 185.615 ;
        RECT 53.260 185.570 53.580 185.630 ;
        RECT 48.215 185.430 53.580 185.570 ;
        RECT 48.215 185.385 48.505 185.430 ;
        RECT 53.260 185.370 53.580 185.430 ;
        RECT 62.935 185.570 63.225 185.615 ;
        RECT 66.600 185.570 66.920 185.630 ;
        RECT 62.935 185.430 66.920 185.570 ;
        RECT 62.935 185.385 63.225 185.430 ;
        RECT 66.600 185.370 66.920 185.430 ;
        RECT 76.720 185.370 77.040 185.630 ;
        RECT 81.780 185.370 82.100 185.630 ;
        RECT 83.635 185.570 83.925 185.615 ;
        RECT 85.000 185.570 85.320 185.630 ;
        RECT 83.635 185.430 85.320 185.570 ;
        RECT 83.635 185.385 83.925 185.430 ;
        RECT 85.000 185.370 85.320 185.430 ;
        RECT 92.835 185.570 93.125 185.615 ;
        RECT 94.660 185.570 94.980 185.630 ;
        RECT 92.835 185.430 94.980 185.570 ;
        RECT 92.835 185.385 93.125 185.430 ;
        RECT 94.660 185.370 94.980 185.430 ;
        RECT 101.100 185.370 101.420 185.630 ;
        RECT 102.020 185.370 102.340 185.630 ;
        RECT 15.010 184.750 113.450 185.230 ;
        RECT 20.615 184.550 20.905 184.595 ;
        RECT 23.360 184.550 23.680 184.610 ;
        RECT 20.615 184.410 23.680 184.550 ;
        RECT 20.615 184.365 20.905 184.410 ;
        RECT 23.360 184.350 23.680 184.410 ;
        RECT 24.740 184.550 25.060 184.610 ;
        RECT 33.035 184.550 33.325 184.595 ;
        RECT 39.920 184.550 40.240 184.610 ;
        RECT 24.740 184.410 40.240 184.550 ;
        RECT 24.740 184.350 25.060 184.410 ;
        RECT 33.035 184.365 33.325 184.410 ;
        RECT 39.920 184.350 40.240 184.410 ;
        RECT 56.020 184.350 56.340 184.610 ;
        RECT 69.360 184.550 69.680 184.610 ;
        RECT 73.745 184.550 74.035 184.595 ;
        RECT 74.420 184.550 74.740 184.610 ;
        RECT 59.330 184.410 68.210 184.550 ;
        RECT 25.165 184.210 25.455 184.255 ;
        RECT 27.055 184.210 27.345 184.255 ;
        RECT 30.175 184.210 30.465 184.255 ;
        RECT 25.165 184.070 30.465 184.210 ;
        RECT 25.165 184.025 25.455 184.070 ;
        RECT 27.055 184.025 27.345 184.070 ;
        RECT 30.175 184.025 30.465 184.070 ;
        RECT 32.100 184.210 32.420 184.270 ;
        RECT 39.475 184.210 39.765 184.255 ;
        RECT 44.060 184.210 44.380 184.270 ;
        RECT 45.900 184.210 46.220 184.270 ;
        RECT 32.100 184.070 39.765 184.210 ;
        RECT 32.100 184.010 32.420 184.070 ;
        RECT 39.475 184.025 39.765 184.070 ;
        RECT 42.770 184.070 46.220 184.210 ;
        RECT 25.660 183.670 25.980 183.930 ;
        RECT 27.960 183.870 28.280 183.930 ;
        RECT 42.770 183.915 42.910 184.070 ;
        RECT 44.060 184.010 44.380 184.070 ;
        RECT 45.900 184.010 46.220 184.070 ;
        RECT 46.475 184.210 46.765 184.255 ;
        RECT 49.595 184.210 49.885 184.255 ;
        RECT 51.485 184.210 51.775 184.255 ;
        RECT 46.475 184.070 51.775 184.210 ;
        RECT 46.475 184.025 46.765 184.070 ;
        RECT 49.595 184.025 49.885 184.070 ;
        RECT 51.485 184.025 51.775 184.070 ;
        RECT 27.960 183.730 35.550 183.870 ;
        RECT 27.960 183.670 28.280 183.730 ;
        RECT 23.820 183.330 24.140 183.590 ;
        RECT 24.295 183.345 24.585 183.575 ;
        RECT 24.760 183.530 25.050 183.575 ;
        RECT 26.595 183.530 26.885 183.575 ;
        RECT 30.175 183.530 30.465 183.575 ;
        RECT 24.760 183.390 30.465 183.530 ;
        RECT 24.760 183.345 25.050 183.390 ;
        RECT 26.595 183.345 26.885 183.390 ;
        RECT 30.175 183.345 30.465 183.390 ;
        RECT 24.370 183.190 24.510 183.345 ;
        RECT 25.200 183.190 25.520 183.250 ;
        RECT 31.255 183.235 31.545 183.550 ;
        RECT 34.415 183.530 34.705 183.575 ;
        RECT 34.860 183.530 35.180 183.590 ;
        RECT 34.415 183.390 35.180 183.530 ;
        RECT 35.410 183.530 35.550 183.730 ;
        RECT 42.695 183.685 42.985 183.915 ;
        RECT 43.600 183.670 43.920 183.930 ;
        RECT 52.355 183.870 52.645 183.915 ;
        RECT 52.800 183.870 53.120 183.930 ;
        RECT 52.355 183.730 53.120 183.870 ;
        RECT 52.355 183.685 52.645 183.730 ;
        RECT 52.800 183.670 53.120 183.730 ;
        RECT 53.260 183.670 53.580 183.930 ;
        RECT 54.640 183.870 54.960 183.930 ;
        RECT 59.330 183.915 59.470 184.410 ;
        RECT 68.070 184.270 68.210 184.410 ;
        RECT 69.360 184.410 71.890 184.550 ;
        RECT 69.360 184.350 69.680 184.410 ;
        RECT 65.235 184.210 65.525 184.255 ;
        RECT 65.680 184.210 66.000 184.270 ;
        RECT 59.790 184.070 66.000 184.210 ;
        RECT 59.790 183.915 59.930 184.070 ;
        RECT 65.235 184.025 65.525 184.070 ;
        RECT 65.680 184.010 66.000 184.070 ;
        RECT 67.980 184.210 68.300 184.270 ;
        RECT 70.280 184.210 70.600 184.270 ;
        RECT 67.980 184.070 71.430 184.210 ;
        RECT 67.980 184.010 68.300 184.070 ;
        RECT 70.280 184.010 70.600 184.070 ;
        RECT 56.955 183.870 57.245 183.915 ;
        RECT 54.640 183.730 57.245 183.870 ;
        RECT 54.640 183.670 54.960 183.730 ;
        RECT 56.955 183.685 57.245 183.730 ;
        RECT 59.255 183.685 59.545 183.915 ;
        RECT 59.715 183.685 60.005 183.915 ;
        RECT 60.175 183.870 60.465 183.915 ;
        RECT 61.540 183.870 61.860 183.930 ;
        RECT 71.290 183.915 71.430 184.070 ;
        RECT 71.750 183.915 71.890 184.410 ;
        RECT 73.745 184.410 74.740 184.550 ;
        RECT 73.745 184.365 74.035 184.410 ;
        RECT 74.420 184.350 74.740 184.410 ;
        RECT 75.340 184.550 75.660 184.610 ;
        RECT 88.220 184.550 88.540 184.610 ;
        RECT 75.340 184.410 88.540 184.550 ;
        RECT 75.340 184.350 75.660 184.410 ;
        RECT 77.610 184.210 77.900 184.255 ;
        RECT 80.390 184.210 80.680 184.255 ;
        RECT 82.250 184.210 82.540 184.255 ;
        RECT 77.610 184.070 82.540 184.210 ;
        RECT 77.610 184.025 77.900 184.070 ;
        RECT 80.390 184.025 80.680 184.070 ;
        RECT 82.250 184.025 82.540 184.070 ;
        RECT 67.535 183.870 67.825 183.915 ;
        RECT 70.755 183.870 71.045 183.915 ;
        RECT 60.175 183.730 71.045 183.870 ;
        RECT 60.175 183.685 60.465 183.730 ;
        RECT 61.540 183.670 61.860 183.730 ;
        RECT 67.535 183.685 67.825 183.730 ;
        RECT 70.755 183.685 71.045 183.730 ;
        RECT 71.215 183.685 71.505 183.915 ;
        RECT 71.675 183.685 71.965 183.915 ;
        RECT 80.875 183.870 81.165 183.915 ;
        RECT 81.780 183.870 82.100 183.930 ;
        RECT 84.170 183.915 84.310 184.410 ;
        RECT 88.220 184.350 88.540 184.410 ;
        RECT 89.155 184.550 89.445 184.595 ;
        RECT 90.520 184.550 90.840 184.610 ;
        RECT 89.155 184.410 90.840 184.550 ;
        RECT 89.155 184.365 89.445 184.410 ;
        RECT 90.520 184.350 90.840 184.410 ;
        RECT 106.620 184.550 106.940 184.610 ;
        RECT 108.935 184.550 109.225 184.595 ;
        RECT 106.620 184.410 109.225 184.550 ;
        RECT 106.620 184.350 106.940 184.410 ;
        RECT 108.935 184.365 109.225 184.410 ;
        RECT 92.015 184.210 92.305 184.255 ;
        RECT 95.135 184.210 95.425 184.255 ;
        RECT 97.025 184.210 97.315 184.255 ;
        RECT 92.015 184.070 97.315 184.210 ;
        RECT 92.015 184.025 92.305 184.070 ;
        RECT 95.135 184.025 95.425 184.070 ;
        RECT 97.025 184.025 97.315 184.070 ;
        RECT 102.135 184.210 102.425 184.255 ;
        RECT 105.255 184.210 105.545 184.255 ;
        RECT 107.145 184.210 107.435 184.255 ;
        RECT 102.135 184.070 107.435 184.210 ;
        RECT 102.135 184.025 102.425 184.070 ;
        RECT 105.255 184.025 105.545 184.070 ;
        RECT 107.145 184.025 107.435 184.070 ;
        RECT 80.875 183.730 82.100 183.870 ;
        RECT 80.875 183.685 81.165 183.730 ;
        RECT 81.780 183.670 82.100 183.730 ;
        RECT 84.095 183.685 84.385 183.915 ;
        RECT 97.895 183.870 98.185 183.915 ;
        RECT 98.340 183.870 98.660 183.930 ;
        RECT 104.780 183.870 105.100 183.930 ;
        RECT 110.760 183.870 111.080 183.930 ;
        RECT 97.895 183.730 105.100 183.870 ;
        RECT 97.895 183.685 98.185 183.730 ;
        RECT 98.340 183.670 98.660 183.730 ;
        RECT 104.780 183.670 105.100 183.730 ;
        RECT 108.090 183.730 111.080 183.870 ;
        RECT 35.410 183.510 37.850 183.530 ;
        RECT 38.095 183.510 38.385 183.575 ;
        RECT 35.410 183.390 38.385 183.510 ;
        RECT 34.415 183.345 34.705 183.390 ;
        RECT 27.955 183.190 28.605 183.235 ;
        RECT 31.255 183.190 31.845 183.235 ;
        RECT 24.370 183.050 24.970 183.190 ;
        RECT 24.830 182.850 24.970 183.050 ;
        RECT 25.200 183.050 31.845 183.190 ;
        RECT 34.490 183.190 34.630 183.345 ;
        RECT 34.860 183.330 35.180 183.390 ;
        RECT 37.710 183.370 38.385 183.390 ;
        RECT 38.095 183.345 38.385 183.370 ;
        RECT 37.160 183.190 37.480 183.250 ;
        RECT 41.775 183.190 42.065 183.235 ;
        RECT 34.490 183.050 37.480 183.190 ;
        RECT 25.200 182.990 25.520 183.050 ;
        RECT 27.955 183.005 28.605 183.050 ;
        RECT 31.555 183.005 31.845 183.050 ;
        RECT 37.160 182.990 37.480 183.050 ;
        RECT 38.170 183.050 42.065 183.190 ;
        RECT 38.170 182.910 38.310 183.050 ;
        RECT 41.775 183.005 42.065 183.050 ;
        RECT 44.060 183.190 44.380 183.250 ;
        RECT 45.395 183.235 45.685 183.550 ;
        RECT 46.475 183.530 46.765 183.575 ;
        RECT 50.055 183.530 50.345 183.575 ;
        RECT 51.890 183.530 52.180 183.575 ;
        RECT 46.475 183.390 52.180 183.530 ;
        RECT 46.475 183.345 46.765 183.390 ;
        RECT 50.055 183.345 50.345 183.390 ;
        RECT 51.890 183.345 52.180 183.390 ;
        RECT 57.415 183.530 57.705 183.575 ;
        RECT 57.860 183.530 58.180 183.590 ;
        RECT 57.415 183.390 58.180 183.530 ;
        RECT 57.415 183.345 57.705 183.390 ;
        RECT 57.860 183.330 58.180 183.390 ;
        RECT 58.795 183.530 59.085 183.575 ;
        RECT 64.760 183.530 65.080 183.590 ;
        RECT 70.295 183.530 70.585 183.575 ;
        RECT 58.795 183.390 70.585 183.530 ;
        RECT 58.795 183.345 59.085 183.390 ;
        RECT 64.760 183.330 65.080 183.390 ;
        RECT 45.095 183.190 45.685 183.235 ;
        RECT 48.335 183.190 48.985 183.235 ;
        RECT 44.060 183.050 48.985 183.190 ;
        RECT 44.060 182.990 44.380 183.050 ;
        RECT 45.095 183.005 45.385 183.050 ;
        RECT 48.335 183.005 48.985 183.050 ;
        RECT 50.960 182.990 51.280 183.250 ;
        RECT 61.080 182.990 61.400 183.250 ;
        RECT 65.310 183.235 65.450 183.390 ;
        RECT 70.295 183.345 70.585 183.390 ;
        RECT 77.610 183.530 77.900 183.575 ;
        RECT 82.715 183.530 83.005 183.575 ;
        RECT 83.620 183.530 83.940 183.590 ;
        RECT 77.610 183.390 80.145 183.530 ;
        RECT 77.610 183.345 77.900 183.390 ;
        RECT 65.235 183.005 65.525 183.235 ;
        RECT 65.680 183.190 66.000 183.250 ;
        RECT 69.375 183.190 69.665 183.235 ;
        RECT 65.680 183.050 69.665 183.190 ;
        RECT 65.680 182.990 66.000 183.050 ;
        RECT 69.375 183.005 69.665 183.050 ;
        RECT 75.750 183.190 76.040 183.235 ;
        RECT 76.720 183.190 77.040 183.250 ;
        RECT 79.930 183.235 80.145 183.390 ;
        RECT 82.715 183.390 83.940 183.530 ;
        RECT 82.715 183.345 83.005 183.390 ;
        RECT 83.620 183.330 83.940 183.390 ;
        RECT 85.000 183.330 85.320 183.590 ;
        RECT 87.760 183.330 88.080 183.590 ;
        RECT 90.935 183.235 91.225 183.550 ;
        RECT 92.015 183.530 92.305 183.575 ;
        RECT 95.595 183.530 95.885 183.575 ;
        RECT 97.430 183.530 97.720 183.575 ;
        RECT 101.100 183.550 101.420 183.590 ;
        RECT 108.090 183.575 108.230 183.730 ;
        RECT 110.760 183.670 111.080 183.730 ;
        RECT 92.015 183.390 97.720 183.530 ;
        RECT 92.015 183.345 92.305 183.390 ;
        RECT 95.595 183.345 95.885 183.390 ;
        RECT 97.430 183.345 97.720 183.390 ;
        RECT 101.055 183.330 101.420 183.550 ;
        RECT 102.135 183.530 102.425 183.575 ;
        RECT 105.715 183.530 106.005 183.575 ;
        RECT 107.550 183.530 107.840 183.575 ;
        RECT 102.135 183.390 107.840 183.530 ;
        RECT 102.135 183.345 102.425 183.390 ;
        RECT 105.715 183.345 106.005 183.390 ;
        RECT 107.550 183.345 107.840 183.390 ;
        RECT 108.015 183.345 108.305 183.575 ;
        RECT 108.475 183.530 108.765 183.575 ;
        RECT 110.300 183.530 110.620 183.590 ;
        RECT 108.475 183.390 110.620 183.530 ;
        RECT 108.475 183.345 108.765 183.390 ;
        RECT 79.010 183.190 79.300 183.235 ;
        RECT 75.750 183.050 79.300 183.190 ;
        RECT 75.750 183.005 76.040 183.050 ;
        RECT 76.720 182.990 77.040 183.050 ;
        RECT 79.010 183.005 79.300 183.050 ;
        RECT 79.930 183.190 80.220 183.235 ;
        RECT 81.790 183.190 82.080 183.235 ;
        RECT 79.930 183.050 82.080 183.190 ;
        RECT 79.930 183.005 80.220 183.050 ;
        RECT 81.790 183.005 82.080 183.050 ;
        RECT 88.235 183.190 88.525 183.235 ;
        RECT 90.635 183.190 91.225 183.235 ;
        RECT 93.875 183.190 94.525 183.235 ;
        RECT 88.235 183.050 94.525 183.190 ;
        RECT 88.235 183.005 88.525 183.050 ;
        RECT 90.635 183.005 90.925 183.050 ;
        RECT 93.875 183.005 94.525 183.050 ;
        RECT 96.500 182.990 96.820 183.250 ;
        RECT 101.055 183.235 101.345 183.330 ;
        RECT 100.755 183.190 101.345 183.235 ;
        RECT 103.995 183.190 104.645 183.235 ;
        RECT 100.755 183.050 104.645 183.190 ;
        RECT 100.755 183.005 101.045 183.050 ;
        RECT 103.995 183.005 104.645 183.050 ;
        RECT 106.620 182.990 106.940 183.250 ;
        RECT 29.340 182.850 29.660 182.910 ;
        RECT 24.830 182.710 29.660 182.850 ;
        RECT 29.340 182.650 29.660 182.710 ;
        RECT 34.860 182.650 35.180 182.910 ;
        RECT 38.080 182.650 38.400 182.910 ;
        RECT 39.015 182.850 39.305 182.895 ;
        RECT 40.380 182.850 40.700 182.910 ;
        RECT 39.015 182.710 40.700 182.850 ;
        RECT 39.015 182.665 39.305 182.710 ;
        RECT 40.380 182.650 40.700 182.710 ;
        RECT 41.315 182.850 41.605 182.895 ;
        RECT 49.120 182.850 49.440 182.910 ;
        RECT 41.315 182.710 49.440 182.850 ;
        RECT 41.315 182.665 41.605 182.710 ;
        RECT 49.120 182.650 49.440 182.710 ;
        RECT 67.980 182.650 68.300 182.910 ;
        RECT 68.900 182.650 69.220 182.910 ;
        RECT 80.860 182.850 81.180 182.910 ;
        RECT 84.555 182.850 84.845 182.895 ;
        RECT 80.860 182.710 84.845 182.850 ;
        RECT 80.860 182.650 81.180 182.710 ;
        RECT 84.555 182.665 84.845 182.710 ;
        RECT 86.855 182.850 87.145 182.895 ;
        RECT 95.120 182.850 95.440 182.910 ;
        RECT 86.855 182.710 95.440 182.850 ;
        RECT 86.855 182.665 87.145 182.710 ;
        RECT 95.120 182.650 95.440 182.710 ;
        RECT 96.040 182.850 96.360 182.910 ;
        RECT 99.275 182.850 99.565 182.895 ;
        RECT 96.040 182.710 99.565 182.850 ;
        RECT 96.040 182.650 96.360 182.710 ;
        RECT 99.275 182.665 99.565 182.710 ;
        RECT 104.780 182.850 105.100 182.910 ;
        RECT 108.090 182.850 108.230 183.345 ;
        RECT 110.300 183.330 110.620 183.390 ;
        RECT 104.780 182.710 108.230 182.850 ;
        RECT 104.780 182.650 105.100 182.710 ;
        RECT 15.010 182.030 113.450 182.510 ;
        RECT 22.455 181.830 22.745 181.875 ;
        RECT 30.735 181.830 31.025 181.875 ;
        RECT 39.920 181.830 40.240 181.890 ;
        RECT 22.455 181.690 30.490 181.830 ;
        RECT 22.455 181.645 22.745 181.690 ;
        RECT 30.350 181.550 30.490 181.690 ;
        RECT 30.735 181.690 40.240 181.830 ;
        RECT 30.735 181.645 31.025 181.690 ;
        RECT 39.920 181.630 40.240 181.690 ;
        RECT 44.060 181.630 44.380 181.890 ;
        RECT 49.120 181.630 49.440 181.890 ;
        RECT 50.960 181.830 51.280 181.890 ;
        RECT 54.195 181.830 54.485 181.875 ;
        RECT 50.960 181.690 54.485 181.830 ;
        RECT 50.960 181.630 51.280 181.690 ;
        RECT 54.195 181.645 54.485 181.690 ;
        RECT 61.540 181.830 61.860 181.890 ;
        RECT 61.540 181.690 65.910 181.830 ;
        RECT 61.540 181.630 61.860 181.690 ;
        RECT 21.060 181.490 21.380 181.550 ;
        RECT 18.850 181.350 21.380 181.490 ;
        RECT 18.850 181.195 18.990 181.350 ;
        RECT 21.060 181.290 21.380 181.350 ;
        RECT 23.820 181.490 24.140 181.550 ;
        RECT 28.420 181.490 28.740 181.550 ;
        RECT 23.820 181.350 28.740 181.490 ;
        RECT 23.820 181.290 24.140 181.350 ;
        RECT 28.420 181.290 28.740 181.350 ;
        RECT 30.260 181.290 30.580 181.550 ;
        RECT 34.515 181.490 34.805 181.535 ;
        RECT 37.755 181.490 38.405 181.535 ;
        RECT 34.515 181.350 38.405 181.490 ;
        RECT 34.515 181.305 35.105 181.350 ;
        RECT 37.755 181.305 38.405 181.350 ;
        RECT 34.815 181.210 35.105 181.305 ;
        RECT 40.380 181.290 40.700 181.550 ;
        RECT 48.215 181.490 48.505 181.535 ;
        RECT 56.940 181.490 57.260 181.550 ;
        RECT 58.795 181.490 59.085 181.535 ;
        RECT 48.215 181.350 55.330 181.490 ;
        RECT 48.215 181.305 48.505 181.350 ;
        RECT 18.775 180.965 19.065 181.195 ;
        RECT 19.695 181.150 19.985 181.195 ;
        RECT 21.980 181.150 22.300 181.210 ;
        RECT 19.695 181.010 22.300 181.150 ;
        RECT 19.695 180.965 19.985 181.010 ;
        RECT 21.980 180.950 22.300 181.010 ;
        RECT 23.375 180.965 23.665 181.195 ;
        RECT 25.215 181.150 25.505 181.195 ;
        RECT 32.100 181.150 32.420 181.210 ;
        RECT 25.215 181.010 32.420 181.150 ;
        RECT 25.215 180.965 25.505 181.010 ;
        RECT 18.315 180.810 18.605 180.855 ;
        RECT 20.140 180.810 20.460 180.870 ;
        RECT 18.315 180.670 20.460 180.810 ;
        RECT 23.450 180.810 23.590 180.965 ;
        RECT 32.100 180.950 32.420 181.010 ;
        RECT 34.815 180.990 35.180 181.210 ;
        RECT 34.860 180.950 35.180 180.990 ;
        RECT 35.895 181.150 36.185 181.195 ;
        RECT 39.475 181.150 39.765 181.195 ;
        RECT 41.310 181.150 41.600 181.195 ;
        RECT 35.895 181.010 41.600 181.150 ;
        RECT 35.895 180.965 36.185 181.010 ;
        RECT 39.475 180.965 39.765 181.010 ;
        RECT 41.310 180.965 41.600 181.010 ;
        RECT 44.520 181.150 44.840 181.210 ;
        RECT 55.190 181.195 55.330 181.350 ;
        RECT 56.940 181.350 59.085 181.490 ;
        RECT 56.940 181.290 57.260 181.350 ;
        RECT 58.795 181.305 59.085 181.350 ;
        RECT 60.710 181.350 64.530 181.490 ;
        RECT 53.735 181.150 54.025 181.195 ;
        RECT 44.520 181.010 54.025 181.150 ;
        RECT 44.520 180.950 44.840 181.010 ;
        RECT 53.735 180.965 54.025 181.010 ;
        RECT 55.115 180.965 55.405 181.195 ;
        RECT 29.800 180.810 30.120 180.870 ;
        RECT 23.450 180.670 30.120 180.810 ;
        RECT 18.315 180.625 18.605 180.670 ;
        RECT 20.140 180.610 20.460 180.670 ;
        RECT 29.800 180.610 30.120 180.670 ;
        RECT 31.180 180.610 31.500 180.870 ;
        RECT 33.035 180.625 33.325 180.855 ;
        RECT 35.320 180.810 35.640 180.870 ;
        RECT 41.775 180.810 42.065 180.855 ;
        RECT 35.320 180.670 42.065 180.810 ;
        RECT 21.520 180.470 21.840 180.530 ;
        RECT 33.110 180.470 33.250 180.625 ;
        RECT 35.320 180.610 35.640 180.670 ;
        RECT 41.775 180.625 42.065 180.670 ;
        RECT 45.455 180.810 45.745 180.855 ;
        RECT 46.360 180.810 46.680 180.870 ;
        RECT 45.455 180.670 46.680 180.810 ;
        RECT 45.455 180.625 45.745 180.670 ;
        RECT 46.360 180.610 46.680 180.670 ;
        RECT 49.580 180.810 49.900 180.870 ;
        RECT 51.895 180.810 52.185 180.855 ;
        RECT 49.580 180.670 52.185 180.810 ;
        RECT 49.580 180.610 49.900 180.670 ;
        RECT 51.895 180.625 52.185 180.670 ;
        RECT 53.260 180.610 53.580 180.870 ;
        RECT 53.810 180.810 53.950 180.965 ;
        RECT 57.400 180.950 57.720 181.210 ;
        RECT 60.160 181.150 60.480 181.210 ;
        RECT 60.710 181.150 60.850 181.350 ;
        RECT 60.160 181.010 60.850 181.150 ;
        RECT 61.080 181.150 61.400 181.210 ;
        RECT 64.390 181.195 64.530 181.350 ;
        RECT 61.555 181.150 61.845 181.195 ;
        RECT 61.080 181.010 61.845 181.150 ;
        RECT 60.160 180.950 60.480 181.010 ;
        RECT 61.080 180.950 61.400 181.010 ;
        RECT 61.555 180.965 61.845 181.010 ;
        RECT 64.315 180.965 64.605 181.195 ;
        RECT 64.760 180.950 65.080 181.210 ;
        RECT 65.220 180.950 65.540 181.210 ;
        RECT 65.770 181.195 65.910 181.690 ;
        RECT 73.960 181.630 74.280 181.890 ;
        RECT 86.840 181.830 87.160 181.890 ;
        RECT 95.595 181.830 95.885 181.875 ;
        RECT 96.500 181.830 96.820 181.890 ;
        RECT 85.090 181.690 93.050 181.830 ;
        RECT 69.835 181.490 70.125 181.535 ;
        RECT 72.135 181.490 72.425 181.535 ;
        RECT 69.835 181.350 72.425 181.490 ;
        RECT 69.835 181.305 70.125 181.350 ;
        RECT 72.135 181.305 72.425 181.350 ;
        RECT 75.800 181.490 76.120 181.550 ;
        RECT 76.375 181.490 76.665 181.535 ;
        RECT 79.615 181.490 80.265 181.535 ;
        RECT 75.800 181.350 80.265 181.490 ;
        RECT 75.800 181.290 76.120 181.350 ;
        RECT 76.375 181.305 76.965 181.350 ;
        RECT 79.615 181.305 80.265 181.350 ;
        RECT 65.695 180.965 65.985 181.195 ;
        RECT 71.675 181.150 71.965 181.195 ;
        RECT 73.040 181.150 73.360 181.210 ;
        RECT 74.420 181.150 74.740 181.210 ;
        RECT 71.675 181.010 74.740 181.150 ;
        RECT 71.675 180.965 71.965 181.010 ;
        RECT 73.040 180.950 73.360 181.010 ;
        RECT 74.420 180.950 74.740 181.010 ;
        RECT 76.675 180.990 76.965 181.305 ;
        RECT 77.755 181.150 78.045 181.195 ;
        RECT 81.335 181.150 81.625 181.195 ;
        RECT 83.170 181.150 83.460 181.195 ;
        RECT 77.755 181.010 83.460 181.150 ;
        RECT 77.755 180.965 78.045 181.010 ;
        RECT 81.335 180.965 81.625 181.010 ;
        RECT 83.170 180.965 83.460 181.010 ;
        RECT 83.620 181.150 83.940 181.210 ;
        RECT 85.090 181.150 85.230 181.690 ;
        RECT 86.840 181.630 87.160 181.690 ;
        RECT 89.140 181.535 89.460 181.550 ;
        RECT 85.575 181.490 85.865 181.535 ;
        RECT 88.815 181.490 89.465 181.535 ;
        RECT 85.575 181.350 89.465 181.490 ;
        RECT 85.575 181.305 86.165 181.350 ;
        RECT 88.815 181.305 89.465 181.350 ;
        RECT 92.910 181.490 93.050 181.690 ;
        RECT 95.595 181.690 96.820 181.830 ;
        RECT 95.595 181.645 95.885 181.690 ;
        RECT 96.500 181.630 96.820 181.690 ;
        RECT 97.420 181.630 97.740 181.890 ;
        RECT 102.495 181.830 102.785 181.875 ;
        RECT 103.400 181.830 103.720 181.890 ;
        RECT 102.495 181.690 103.720 181.830 ;
        RECT 102.495 181.645 102.785 181.690 ;
        RECT 103.400 181.630 103.720 181.690 ;
        RECT 104.335 181.645 104.625 181.875 ;
        RECT 98.340 181.490 98.660 181.550 ;
        RECT 92.910 181.350 98.660 181.490 ;
        RECT 104.410 181.490 104.550 181.645 ;
        RECT 104.410 181.350 111.450 181.490 ;
        RECT 83.620 181.010 85.230 181.150 ;
        RECT 83.620 180.950 83.940 181.010 ;
        RECT 85.875 180.990 86.165 181.305 ;
        RECT 89.140 181.290 89.460 181.305 ;
        RECT 92.910 181.195 93.050 181.350 ;
        RECT 98.340 181.290 98.660 181.350 ;
        RECT 86.955 181.150 87.245 181.195 ;
        RECT 90.535 181.150 90.825 181.195 ;
        RECT 92.370 181.150 92.660 181.195 ;
        RECT 86.955 181.010 92.660 181.150 ;
        RECT 86.955 180.965 87.245 181.010 ;
        RECT 90.535 180.965 90.825 181.010 ;
        RECT 92.370 180.965 92.660 181.010 ;
        RECT 92.835 180.965 93.125 181.195 ;
        RECT 94.215 180.965 94.505 181.195 ;
        RECT 57.860 180.810 58.180 180.870 ;
        RECT 59.240 180.810 59.560 180.870 ;
        RECT 53.810 180.670 59.560 180.810 ;
        RECT 57.860 180.610 58.180 180.670 ;
        RECT 59.240 180.610 59.560 180.670 ;
        RECT 60.620 180.610 60.940 180.870 ;
        RECT 63.395 180.810 63.685 180.855 ;
        RECT 63.840 180.810 64.160 180.870 ;
        RECT 63.395 180.670 64.160 180.810 ;
        RECT 63.395 180.625 63.685 180.670 ;
        RECT 63.840 180.610 64.160 180.670 ;
        RECT 67.075 180.810 67.365 180.855 ;
        RECT 69.360 180.810 69.680 180.870 ;
        RECT 67.075 180.670 69.680 180.810 ;
        RECT 67.075 180.625 67.365 180.670 ;
        RECT 69.360 180.610 69.680 180.670 ;
        RECT 70.740 180.610 71.060 180.870 ;
        RECT 74.895 180.625 75.185 180.855 ;
        RECT 91.455 180.810 91.745 180.855 ;
        RECT 94.290 180.810 94.430 180.965 ;
        RECT 94.660 180.950 94.980 181.210 ;
        RECT 111.310 181.195 111.450 181.350 ;
        RECT 97.895 181.150 98.185 181.195 ;
        RECT 104.795 181.150 105.085 181.195 ;
        RECT 97.895 181.010 105.085 181.150 ;
        RECT 97.895 180.965 98.185 181.010 ;
        RECT 104.795 180.965 105.085 181.010 ;
        RECT 111.235 180.965 111.525 181.195 ;
        RECT 95.120 180.810 95.440 180.870 ;
        RECT 91.455 180.670 93.510 180.810 ;
        RECT 94.290 180.670 95.440 180.810 ;
        RECT 91.455 180.625 91.745 180.670 ;
        RECT 21.520 180.330 33.250 180.470 ;
        RECT 21.520 180.270 21.840 180.330 ;
        RECT 24.280 179.930 24.600 180.190 ;
        RECT 27.960 179.930 28.280 180.190 ;
        RECT 28.420 179.930 28.740 180.190 ;
        RECT 33.110 180.130 33.250 180.330 ;
        RECT 35.895 180.470 36.185 180.515 ;
        RECT 39.015 180.470 39.305 180.515 ;
        RECT 40.905 180.470 41.195 180.515 ;
        RECT 35.895 180.330 41.195 180.470 ;
        RECT 69.450 180.470 69.590 180.610 ;
        RECT 74.970 180.470 75.110 180.625 ;
        RECT 69.450 180.330 75.110 180.470 ;
        RECT 77.755 180.470 78.045 180.515 ;
        RECT 80.875 180.470 81.165 180.515 ;
        RECT 82.765 180.470 83.055 180.515 ;
        RECT 77.755 180.330 83.055 180.470 ;
        RECT 35.895 180.285 36.185 180.330 ;
        RECT 39.015 180.285 39.305 180.330 ;
        RECT 40.905 180.285 41.195 180.330 ;
        RECT 77.755 180.285 78.045 180.330 ;
        RECT 80.875 180.285 81.165 180.330 ;
        RECT 82.765 180.285 83.055 180.330 ;
        RECT 84.080 180.270 84.400 180.530 ;
        RECT 93.370 180.515 93.510 180.670 ;
        RECT 95.120 180.610 95.440 180.670 ;
        RECT 96.960 180.810 97.280 180.870 ;
        RECT 101.115 180.810 101.405 180.855 ;
        RECT 96.960 180.670 101.405 180.810 ;
        RECT 96.960 180.610 97.280 180.670 ;
        RECT 101.115 180.625 101.405 180.670 ;
        RECT 102.020 180.810 102.340 180.870 ;
        RECT 107.555 180.810 107.845 180.855 ;
        RECT 102.020 180.670 107.845 180.810 ;
        RECT 102.020 180.610 102.340 180.670 ;
        RECT 107.555 180.625 107.845 180.670 ;
        RECT 86.955 180.470 87.245 180.515 ;
        RECT 90.075 180.470 90.365 180.515 ;
        RECT 91.965 180.470 92.255 180.515 ;
        RECT 86.955 180.330 92.255 180.470 ;
        RECT 86.955 180.285 87.245 180.330 ;
        RECT 90.075 180.285 90.365 180.330 ;
        RECT 91.965 180.285 92.255 180.330 ;
        RECT 93.295 180.285 93.585 180.515 ;
        RECT 38.080 180.130 38.400 180.190 ;
        RECT 33.110 179.990 38.400 180.130 ;
        RECT 38.080 179.930 38.400 179.990 ;
        RECT 40.380 180.130 40.700 180.190 ;
        RECT 62.475 180.130 62.765 180.175 ;
        RECT 81.780 180.130 82.100 180.190 ;
        RECT 40.380 179.990 82.100 180.130 ;
        RECT 40.380 179.930 40.700 179.990 ;
        RECT 62.475 179.945 62.765 179.990 ;
        RECT 81.780 179.930 82.100 179.990 ;
        RECT 82.350 180.130 82.640 180.175 ;
        RECT 91.440 180.130 91.760 180.190 ;
        RECT 82.350 179.990 91.760 180.130 ;
        RECT 82.350 179.945 82.640 179.990 ;
        RECT 91.440 179.930 91.760 179.990 ;
        RECT 99.735 180.130 100.025 180.175 ;
        RECT 105.700 180.130 106.020 180.190 ;
        RECT 99.735 179.990 106.020 180.130 ;
        RECT 99.735 179.945 100.025 179.990 ;
        RECT 105.700 179.930 106.020 179.990 ;
        RECT 107.080 180.130 107.400 180.190 ;
        RECT 108.475 180.130 108.765 180.175 ;
        RECT 107.080 179.990 108.765 180.130 ;
        RECT 107.080 179.930 107.400 179.990 ;
        RECT 108.475 179.945 108.765 179.990 ;
        RECT 15.010 179.310 113.450 179.790 ;
        RECT 41.300 179.110 41.620 179.170 ;
        RECT 62.475 179.110 62.765 179.155 ;
        RECT 80.400 179.110 80.720 179.170 ;
        RECT 40.930 178.970 80.720 179.110 ;
        RECT 24.855 178.770 25.145 178.815 ;
        RECT 27.975 178.770 28.265 178.815 ;
        RECT 29.865 178.770 30.155 178.815 ;
        RECT 24.855 178.630 30.155 178.770 ;
        RECT 24.855 178.585 25.145 178.630 ;
        RECT 27.975 178.585 28.265 178.630 ;
        RECT 29.865 178.585 30.155 178.630 ;
        RECT 31.640 178.570 31.960 178.830 ;
        RECT 18.775 178.430 19.065 178.475 ;
        RECT 21.520 178.430 21.840 178.490 ;
        RECT 18.775 178.290 21.840 178.430 ;
        RECT 18.775 178.245 19.065 178.290 ;
        RECT 21.520 178.230 21.840 178.290 ;
        RECT 21.980 178.230 22.300 178.490 ;
        RECT 24.280 178.430 24.600 178.490 ;
        RECT 29.355 178.430 29.645 178.475 ;
        RECT 24.280 178.290 29.645 178.430 ;
        RECT 24.280 178.230 24.600 178.290 ;
        RECT 29.355 178.245 29.645 178.290 ;
        RECT 31.180 178.430 31.500 178.490 ;
        RECT 34.415 178.430 34.705 178.475 ;
        RECT 40.380 178.430 40.700 178.490 ;
        RECT 31.180 178.290 34.705 178.430 ;
        RECT 31.180 178.230 31.500 178.290 ;
        RECT 34.415 178.245 34.705 178.290 ;
        RECT 39.090 178.290 40.700 178.430 ;
        RECT 20.140 177.750 20.460 177.810 ;
        RECT 23.775 177.795 24.065 178.110 ;
        RECT 24.855 178.090 25.145 178.135 ;
        RECT 28.435 178.090 28.725 178.135 ;
        RECT 30.270 178.090 30.560 178.135 ;
        RECT 24.855 177.950 30.560 178.090 ;
        RECT 24.855 177.905 25.145 177.950 ;
        RECT 28.435 177.905 28.725 177.950 ;
        RECT 30.270 177.905 30.560 177.950 ;
        RECT 30.735 177.905 31.025 178.135 ;
        RECT 37.635 177.905 37.925 178.135 ;
        RECT 38.080 178.090 38.400 178.150 ;
        RECT 39.090 178.135 39.230 178.290 ;
        RECT 40.380 178.230 40.700 178.290 ;
        RECT 38.555 178.090 38.845 178.135 ;
        RECT 38.080 177.950 38.845 178.090 ;
        RECT 23.475 177.750 24.065 177.795 ;
        RECT 26.715 177.750 27.365 177.795 ;
        RECT 20.140 177.610 27.365 177.750 ;
        RECT 20.140 177.550 20.460 177.610 ;
        RECT 23.475 177.565 23.765 177.610 ;
        RECT 26.715 177.565 27.365 177.610 ;
        RECT 29.340 177.750 29.660 177.810 ;
        RECT 30.810 177.750 30.950 177.905 ;
        RECT 29.340 177.610 30.950 177.750 ;
        RECT 32.100 177.750 32.420 177.810 ;
        RECT 37.710 177.750 37.850 177.905 ;
        RECT 38.080 177.890 38.400 177.950 ;
        RECT 38.555 177.905 38.845 177.950 ;
        RECT 39.015 177.905 39.305 178.135 ;
        RECT 39.475 178.090 39.765 178.135 ;
        RECT 40.930 178.090 41.070 178.970 ;
        RECT 41.300 178.910 41.620 178.970 ;
        RECT 62.475 178.925 62.765 178.970 ;
        RECT 80.400 178.910 80.720 178.970 ;
        RECT 80.860 178.910 81.180 179.170 ;
        RECT 89.140 179.110 89.460 179.170 ;
        RECT 92.835 179.110 93.125 179.155 ;
        RECT 89.140 178.970 93.125 179.110 ;
        RECT 89.140 178.910 89.460 178.970 ;
        RECT 92.835 178.925 93.125 178.970 ;
        RECT 106.620 178.910 106.940 179.170 ;
        RECT 108.935 179.110 109.225 179.155 ;
        RECT 109.840 179.110 110.160 179.170 ;
        RECT 108.935 178.970 110.160 179.110 ;
        RECT 108.935 178.925 109.225 178.970 ;
        RECT 109.840 178.910 110.160 178.970 ;
        RECT 44.995 178.770 45.285 178.815 ;
        RECT 46.360 178.770 46.680 178.830 ;
        RECT 44.995 178.630 46.680 178.770 ;
        RECT 44.995 178.585 45.285 178.630 ;
        RECT 46.360 178.570 46.680 178.630 ;
        RECT 52.800 178.570 53.120 178.830 ;
        RECT 64.775 178.770 65.065 178.815 ;
        RECT 68.440 178.770 68.760 178.830 ;
        RECT 60.710 178.630 68.760 178.770 ;
        RECT 43.600 178.430 43.920 178.490 ;
        RECT 42.310 178.290 43.920 178.430 ;
        RECT 42.310 178.135 42.450 178.290 ;
        RECT 43.600 178.230 43.920 178.290 ;
        RECT 44.060 178.430 44.380 178.490 ;
        RECT 44.535 178.430 44.825 178.475 ;
        RECT 44.060 178.290 44.825 178.430 ;
        RECT 44.060 178.230 44.380 178.290 ;
        RECT 44.535 178.245 44.825 178.290 ;
        RECT 45.900 178.430 46.220 178.490 ;
        RECT 47.755 178.430 48.045 178.475 ;
        RECT 50.055 178.430 50.345 178.475 ;
        RECT 53.735 178.430 54.025 178.475 ;
        RECT 57.875 178.430 58.165 178.475 ;
        RECT 45.900 178.290 58.165 178.430 ;
        RECT 45.900 178.230 46.220 178.290 ;
        RECT 47.755 178.245 48.045 178.290 ;
        RECT 50.055 178.245 50.345 178.290 ;
        RECT 53.735 178.245 54.025 178.290 ;
        RECT 57.875 178.245 58.165 178.290 ;
        RECT 39.475 177.950 41.070 178.090 ;
        RECT 39.475 177.905 39.765 177.950 ;
        RECT 41.315 177.905 41.605 178.135 ;
        RECT 42.235 177.905 42.525 178.135 ;
        RECT 41.390 177.750 41.530 177.905 ;
        RECT 42.680 177.890 43.000 178.150 ;
        RECT 43.155 177.905 43.445 178.135 ;
        RECT 43.690 178.090 43.830 178.230 ;
        RECT 47.295 178.090 47.585 178.135 ;
        RECT 49.580 178.090 49.900 178.150 ;
        RECT 43.690 177.950 49.900 178.090 ;
        RECT 47.295 177.905 47.585 177.950 ;
        RECT 32.100 177.610 34.170 177.750 ;
        RECT 37.710 177.610 41.530 177.750 ;
        RECT 43.230 177.750 43.370 177.905 ;
        RECT 49.580 177.890 49.900 177.950 ;
        RECT 50.500 178.090 50.820 178.150 ;
        RECT 55.115 178.090 55.405 178.135 ;
        RECT 60.710 178.090 60.850 178.630 ;
        RECT 64.775 178.585 65.065 178.630 ;
        RECT 68.440 178.570 68.760 178.630 ;
        RECT 69.360 178.770 69.680 178.830 ;
        RECT 81.780 178.770 82.100 178.830 ;
        RECT 90.980 178.770 91.300 178.830 ;
        RECT 69.360 178.630 78.330 178.770 ;
        RECT 69.360 178.570 69.680 178.630 ;
        RECT 61.540 178.430 61.860 178.490 ;
        RECT 66.155 178.430 66.445 178.475 ;
        RECT 70.740 178.430 71.060 178.490 ;
        RECT 75.340 178.430 75.660 178.490 ;
        RECT 78.190 178.475 78.330 178.630 ;
        RECT 81.780 178.630 91.300 178.770 ;
        RECT 81.780 178.570 82.100 178.630 ;
        RECT 90.980 178.570 91.300 178.630 ;
        RECT 95.670 178.630 104.550 178.770 ;
        RECT 77.195 178.430 77.485 178.475 ;
        RECT 61.540 178.290 66.445 178.430 ;
        RECT 61.540 178.230 61.860 178.290 ;
        RECT 66.155 178.245 66.445 178.290 ;
        RECT 66.690 178.290 68.210 178.430 ;
        RECT 50.500 177.950 55.405 178.090 ;
        RECT 50.500 177.890 50.820 177.950 ;
        RECT 55.115 177.905 55.405 177.950 ;
        RECT 56.800 177.950 60.850 178.090 ;
        RECT 46.360 177.750 46.680 177.810 ;
        RECT 56.800 177.750 56.940 177.950 ;
        RECT 61.080 177.890 61.400 178.150 ;
        RECT 63.395 178.090 63.685 178.135 ;
        RECT 63.855 178.090 64.145 178.135 ;
        RECT 65.680 178.090 66.000 178.150 ;
        RECT 66.690 178.090 66.830 178.290 ;
        RECT 63.395 177.950 66.000 178.090 ;
        RECT 63.395 177.905 63.685 177.950 ;
        RECT 63.855 177.905 64.145 177.950 ;
        RECT 65.680 177.890 66.000 177.950 ;
        RECT 66.230 177.950 66.830 178.090 ;
        RECT 43.230 177.610 56.940 177.750 ;
        RECT 59.255 177.750 59.545 177.795 ;
        RECT 66.230 177.750 66.370 177.950 ;
        RECT 67.060 177.890 67.380 178.150 ;
        RECT 67.535 177.905 67.825 178.135 ;
        RECT 59.255 177.610 66.370 177.750 ;
        RECT 29.340 177.550 29.660 177.610 ;
        RECT 32.100 177.550 32.420 177.610 ;
        RECT 34.030 177.455 34.170 177.610 ;
        RECT 21.535 177.410 21.825 177.455 ;
        RECT 33.495 177.410 33.785 177.455 ;
        RECT 21.535 177.270 33.785 177.410 ;
        RECT 21.535 177.225 21.825 177.270 ;
        RECT 33.495 177.225 33.785 177.270 ;
        RECT 33.955 177.410 34.245 177.455 ;
        RECT 36.700 177.410 37.020 177.470 ;
        RECT 33.955 177.270 37.020 177.410 ;
        RECT 33.955 177.225 34.245 177.270 ;
        RECT 36.700 177.210 37.020 177.270 ;
        RECT 40.840 177.210 41.160 177.470 ;
        RECT 41.390 177.410 41.530 177.610 ;
        RECT 46.360 177.550 46.680 177.610 ;
        RECT 59.255 177.565 59.545 177.610 ;
        RECT 43.140 177.410 43.460 177.470 ;
        RECT 41.390 177.270 43.460 177.410 ;
        RECT 43.140 177.210 43.460 177.270 ;
        RECT 44.520 177.410 44.840 177.470 ;
        RECT 46.835 177.410 47.125 177.455 ;
        RECT 50.515 177.410 50.805 177.455 ;
        RECT 44.520 177.270 50.805 177.410 ;
        RECT 44.520 177.210 44.840 177.270 ;
        RECT 46.835 177.225 47.125 177.270 ;
        RECT 50.515 177.225 50.805 177.270 ;
        RECT 50.975 177.410 51.265 177.455 ;
        RECT 51.880 177.410 52.200 177.470 ;
        RECT 54.655 177.410 54.945 177.455 ;
        RECT 50.975 177.270 54.945 177.410 ;
        RECT 50.975 177.225 51.265 177.270 ;
        RECT 51.880 177.210 52.200 177.270 ;
        RECT 54.655 177.225 54.945 177.270 ;
        RECT 56.955 177.410 57.245 177.455 ;
        RECT 58.780 177.410 59.100 177.470 ;
        RECT 56.955 177.270 59.100 177.410 ;
        RECT 56.955 177.225 57.245 177.270 ;
        RECT 58.780 177.210 59.100 177.270 ;
        RECT 59.700 177.410 60.020 177.470 ;
        RECT 60.175 177.410 60.465 177.455 ;
        RECT 59.700 177.270 60.465 177.410 ;
        RECT 59.700 177.210 60.020 177.270 ;
        RECT 60.175 177.225 60.465 177.270 ;
        RECT 60.620 177.410 60.940 177.470 ;
        RECT 65.680 177.410 66.000 177.470 ;
        RECT 67.610 177.410 67.750 177.905 ;
        RECT 68.070 177.795 68.210 178.290 ;
        RECT 70.740 178.290 77.485 178.430 ;
        RECT 70.740 178.230 71.060 178.290 ;
        RECT 75.340 178.230 75.660 178.290 ;
        RECT 77.195 178.245 77.485 178.290 ;
        RECT 78.115 178.245 78.405 178.475 ;
        RECT 91.070 178.430 91.210 178.570 ;
        RECT 90.610 178.290 91.210 178.430 ;
        RECT 94.660 178.430 94.980 178.490 ;
        RECT 95.670 178.430 95.810 178.630 ;
        RECT 104.410 178.430 104.550 178.630 ;
        RECT 105.700 178.430 106.020 178.490 ;
        RECT 107.080 178.430 107.400 178.490 ;
        RECT 94.660 178.290 95.810 178.430 ;
        RECT 68.440 178.090 68.760 178.150 ;
        RECT 72.120 178.090 72.440 178.150 ;
        RECT 73.055 178.090 73.345 178.135 ;
        RECT 68.440 177.950 73.345 178.090 ;
        RECT 68.440 177.890 68.760 177.950 ;
        RECT 72.120 177.890 72.440 177.950 ;
        RECT 73.055 177.905 73.345 177.950 ;
        RECT 73.500 177.890 73.820 178.150 ;
        RECT 73.975 177.905 74.265 178.135 ;
        RECT 67.995 177.750 68.285 177.795 ;
        RECT 69.375 177.750 69.665 177.795 ;
        RECT 67.995 177.610 69.665 177.750 ;
        RECT 67.995 177.565 68.285 177.610 ;
        RECT 69.375 177.565 69.665 177.610 ;
        RECT 60.620 177.270 67.750 177.410 ;
        RECT 71.200 177.410 71.520 177.470 ;
        RECT 71.675 177.410 71.965 177.455 ;
        RECT 71.200 177.270 71.965 177.410 ;
        RECT 74.050 177.410 74.190 177.905 ;
        RECT 74.880 177.890 75.200 178.150 ;
        RECT 75.800 177.890 76.120 178.150 ;
        RECT 76.260 177.890 76.580 178.150 ;
        RECT 78.575 178.090 78.865 178.135 ;
        RECT 80.860 178.090 81.180 178.150 ;
        RECT 78.575 177.950 81.180 178.090 ;
        RECT 78.575 177.905 78.865 177.950 ;
        RECT 80.860 177.890 81.180 177.950 ;
        RECT 83.635 178.090 83.925 178.135 ;
        RECT 84.080 178.090 84.400 178.150 ;
        RECT 83.635 177.950 84.400 178.090 ;
        RECT 83.635 177.905 83.925 177.950 ;
        RECT 77.640 177.750 77.960 177.810 ;
        RECT 83.710 177.750 83.850 177.905 ;
        RECT 84.080 177.890 84.400 177.950 ;
        RECT 84.540 177.890 84.860 178.150 ;
        RECT 90.060 178.135 90.380 178.150 ;
        RECT 90.610 178.135 90.750 178.290 ;
        RECT 94.660 178.230 94.980 178.290 ;
        RECT 89.845 177.905 90.380 178.135 ;
        RECT 90.535 177.905 90.825 178.135 ;
        RECT 90.060 177.890 90.380 177.905 ;
        RECT 90.980 177.890 91.300 178.150 ;
        RECT 91.900 178.135 92.220 178.150 ;
        RECT 91.885 178.090 92.220 178.135 ;
        RECT 91.725 177.950 92.220 178.090 ;
        RECT 91.885 177.905 92.220 177.950 ;
        RECT 93.295 178.090 93.585 178.135 ;
        RECT 93.295 177.950 94.890 178.090 ;
        RECT 93.295 177.905 93.585 177.950 ;
        RECT 91.900 177.890 92.220 177.905 ;
        RECT 77.640 177.610 83.850 177.750 ;
        RECT 85.000 177.750 85.320 177.810 ;
        RECT 85.935 177.750 86.225 177.795 ;
        RECT 87.760 177.750 88.080 177.810 ;
        RECT 93.370 177.750 93.510 177.905 ;
        RECT 85.000 177.610 93.510 177.750 ;
        RECT 77.640 177.550 77.960 177.610 ;
        RECT 85.000 177.550 85.320 177.610 ;
        RECT 85.935 177.565 86.225 177.610 ;
        RECT 87.760 177.550 88.080 177.610 ;
        RECT 79.480 177.410 79.800 177.470 ;
        RECT 74.050 177.270 79.800 177.410 ;
        RECT 60.620 177.210 60.940 177.270 ;
        RECT 65.680 177.210 66.000 177.270 ;
        RECT 71.200 177.210 71.520 177.270 ;
        RECT 71.675 177.225 71.965 177.270 ;
        RECT 79.480 177.210 79.800 177.270 ;
        RECT 80.400 177.210 80.720 177.470 ;
        RECT 88.695 177.410 88.985 177.455 ;
        RECT 90.060 177.410 90.380 177.470 ;
        RECT 88.695 177.270 90.380 177.410 ;
        RECT 88.695 177.225 88.985 177.270 ;
        RECT 90.060 177.210 90.380 177.270 ;
        RECT 91.900 177.410 92.220 177.470 ;
        RECT 93.755 177.410 94.045 177.455 ;
        RECT 91.900 177.270 94.045 177.410 ;
        RECT 94.750 177.410 94.890 177.950 ;
        RECT 95.120 177.890 95.440 178.150 ;
        RECT 95.670 178.135 95.810 178.290 ;
        RECT 97.050 178.290 104.090 178.430 ;
        RECT 104.410 178.290 105.010 178.430 ;
        RECT 97.050 178.150 97.190 178.290 ;
        RECT 95.595 177.905 95.885 178.135 ;
        RECT 96.040 177.890 96.360 178.150 ;
        RECT 96.960 177.890 97.280 178.150 ;
        RECT 102.495 178.090 102.785 178.135 ;
        RECT 103.400 178.090 103.720 178.150 ;
        RECT 102.495 177.950 103.720 178.090 ;
        RECT 102.495 177.905 102.785 177.950 ;
        RECT 103.400 177.890 103.720 177.950 ;
        RECT 97.420 177.750 97.740 177.810 ;
        RECT 102.955 177.750 103.245 177.795 ;
        RECT 97.420 177.610 103.245 177.750 ;
        RECT 103.950 177.750 104.090 178.290 ;
        RECT 104.320 177.890 104.640 178.150 ;
        RECT 104.870 178.135 105.010 178.290 ;
        RECT 105.700 178.290 106.850 178.430 ;
        RECT 105.700 178.230 106.020 178.290 ;
        RECT 104.795 177.905 105.085 178.135 ;
        RECT 105.240 177.890 105.560 178.150 ;
        RECT 106.175 177.905 106.465 178.135 ;
        RECT 106.710 178.090 106.850 178.290 ;
        RECT 107.080 178.290 108.230 178.430 ;
        RECT 107.080 178.230 107.400 178.290 ;
        RECT 108.090 178.135 108.230 178.290 ;
        RECT 107.555 178.090 107.845 178.135 ;
        RECT 106.710 177.950 107.845 178.090 ;
        RECT 107.555 177.905 107.845 177.950 ;
        RECT 108.015 177.905 108.305 178.135 ;
        RECT 106.250 177.750 106.390 177.905 ;
        RECT 103.950 177.610 106.390 177.750 ;
        RECT 97.420 177.550 97.740 177.610 ;
        RECT 102.955 177.565 103.245 177.610 ;
        RECT 98.800 177.410 99.120 177.470 ;
        RECT 94.750 177.270 99.120 177.410 ;
        RECT 91.900 177.210 92.220 177.270 ;
        RECT 93.755 177.225 94.045 177.270 ;
        RECT 98.800 177.210 99.120 177.270 ;
        RECT 99.260 177.210 99.580 177.470 ;
        RECT 15.010 176.590 113.450 177.070 ;
        RECT 26.580 176.390 26.900 176.450 ;
        RECT 32.100 176.390 32.420 176.450 ;
        RECT 35.795 176.390 36.085 176.435 ;
        RECT 43.140 176.390 43.460 176.450 ;
        RECT 26.580 176.250 32.420 176.390 ;
        RECT 26.580 176.190 26.900 176.250 ;
        RECT 32.100 176.190 32.420 176.250 ;
        RECT 34.030 176.250 36.085 176.390 ;
        RECT 34.030 176.095 34.170 176.250 ;
        RECT 35.795 176.205 36.085 176.250 ;
        RECT 37.710 176.250 43.460 176.390 ;
        RECT 25.675 176.050 25.965 176.095 ;
        RECT 28.075 176.050 28.365 176.095 ;
        RECT 31.315 176.050 31.965 176.095 ;
        RECT 25.675 175.910 31.965 176.050 ;
        RECT 25.675 175.865 25.965 175.910 ;
        RECT 28.075 175.865 28.665 175.910 ;
        RECT 31.315 175.865 31.965 175.910 ;
        RECT 33.955 175.865 34.245 176.095 ;
        RECT 21.060 175.710 21.380 175.770 ;
        RECT 25.200 175.710 25.520 175.770 ;
        RECT 21.060 175.570 25.520 175.710 ;
        RECT 21.060 175.510 21.380 175.570 ;
        RECT 25.200 175.510 25.520 175.570 ;
        RECT 28.375 175.550 28.665 175.865 ;
        RECT 37.710 175.755 37.850 176.250 ;
        RECT 43.140 176.190 43.460 176.250 ;
        RECT 44.520 176.190 44.840 176.450 ;
        RECT 61.080 176.390 61.400 176.450 ;
        RECT 61.555 176.390 61.845 176.435 ;
        RECT 46.910 176.250 56.940 176.390 ;
        RECT 42.680 176.050 43.000 176.110 ;
        RECT 45.900 176.050 46.220 176.110 ;
        RECT 46.910 176.050 47.050 176.250 ;
        RECT 39.090 175.910 47.050 176.050 ;
        RECT 39.090 175.770 39.230 175.910 ;
        RECT 42.680 175.850 43.000 175.910 ;
        RECT 45.900 175.850 46.220 175.910 ;
        RECT 29.455 175.710 29.745 175.755 ;
        RECT 33.035 175.710 33.325 175.755 ;
        RECT 34.870 175.710 35.160 175.755 ;
        RECT 29.455 175.570 35.160 175.710 ;
        RECT 29.455 175.525 29.745 175.570 ;
        RECT 33.035 175.525 33.325 175.570 ;
        RECT 34.870 175.525 35.160 175.570 ;
        RECT 36.715 175.525 37.005 175.755 ;
        RECT 37.635 175.525 37.925 175.755 ;
        RECT 19.695 175.370 19.985 175.415 ;
        RECT 31.640 175.370 31.960 175.430 ;
        RECT 19.695 175.230 31.960 175.370 ;
        RECT 19.695 175.185 19.985 175.230 ;
        RECT 31.640 175.170 31.960 175.230 ;
        RECT 35.320 175.170 35.640 175.430 ;
        RECT 29.455 175.030 29.745 175.075 ;
        RECT 32.575 175.030 32.865 175.075 ;
        RECT 34.465 175.030 34.755 175.075 ;
        RECT 29.455 174.890 34.755 175.030 ;
        RECT 29.455 174.845 29.745 174.890 ;
        RECT 32.575 174.845 32.865 174.890 ;
        RECT 34.465 174.845 34.755 174.890 ;
        RECT 22.455 174.690 22.745 174.735 ;
        RECT 36.790 174.690 36.930 175.525 ;
        RECT 38.540 175.510 38.860 175.770 ;
        RECT 39.000 175.510 39.320 175.770 ;
        RECT 39.475 175.710 39.765 175.755 ;
        RECT 46.360 175.710 46.680 175.770 ;
        RECT 46.910 175.755 47.050 175.910 ;
        RECT 50.615 176.050 50.905 176.095 ;
        RECT 53.260 176.050 53.580 176.110 ;
        RECT 53.855 176.050 54.505 176.095 ;
        RECT 50.615 175.910 54.505 176.050 ;
        RECT 56.800 176.050 56.940 176.250 ;
        RECT 61.080 176.250 61.845 176.390 ;
        RECT 61.080 176.190 61.400 176.250 ;
        RECT 61.555 176.205 61.845 176.250 ;
        RECT 63.395 176.205 63.685 176.435 ;
        RECT 81.795 176.390 82.085 176.435 ;
        RECT 74.050 176.250 76.950 176.390 ;
        RECT 63.470 176.050 63.610 176.205 ;
        RECT 73.500 176.050 73.820 176.110 ;
        RECT 74.050 176.050 74.190 176.250 ;
        RECT 56.800 175.910 74.190 176.050 ;
        RECT 50.615 175.865 51.205 175.910 ;
        RECT 39.475 175.570 46.680 175.710 ;
        RECT 39.475 175.525 39.765 175.570 ;
        RECT 46.360 175.510 46.680 175.570 ;
        RECT 46.835 175.525 47.125 175.755 ;
        RECT 47.295 175.525 47.585 175.755 ;
        RECT 48.215 175.710 48.505 175.755 ;
        RECT 48.215 175.570 49.810 175.710 ;
        RECT 48.215 175.525 48.505 175.570 ;
        RECT 41.775 175.370 42.065 175.415 ;
        RECT 47.370 175.370 47.510 175.525 ;
        RECT 49.135 175.370 49.425 175.415 ;
        RECT 41.775 175.230 49.425 175.370 ;
        RECT 41.775 175.185 42.065 175.230 ;
        RECT 49.135 175.185 49.425 175.230 ;
        RECT 43.140 175.030 43.460 175.090 ;
        RECT 43.140 174.890 45.670 175.030 ;
        RECT 43.140 174.830 43.460 174.890 ;
        RECT 45.530 174.750 45.670 174.890 ;
        RECT 22.455 174.550 36.930 174.690 ;
        RECT 40.380 174.690 40.700 174.750 ;
        RECT 40.855 174.690 41.145 174.735 ;
        RECT 40.380 174.550 41.145 174.690 ;
        RECT 22.455 174.505 22.745 174.550 ;
        RECT 40.380 174.490 40.700 174.550 ;
        RECT 40.855 174.505 41.145 174.550 ;
        RECT 44.980 174.490 45.300 174.750 ;
        RECT 45.440 174.690 45.760 174.750 ;
        RECT 49.670 174.690 49.810 175.570 ;
        RECT 50.915 175.550 51.205 175.865 ;
        RECT 53.260 175.850 53.580 175.910 ;
        RECT 53.855 175.865 54.505 175.910 ;
        RECT 51.995 175.710 52.285 175.755 ;
        RECT 55.575 175.710 55.865 175.755 ;
        RECT 57.410 175.710 57.700 175.755 ;
        RECT 51.995 175.570 57.700 175.710 ;
        RECT 51.995 175.525 52.285 175.570 ;
        RECT 55.575 175.525 55.865 175.570 ;
        RECT 57.410 175.525 57.700 175.570 ;
        RECT 57.875 175.710 58.165 175.755 ;
        RECT 58.320 175.710 58.640 175.770 ;
        RECT 57.875 175.570 58.640 175.710 ;
        RECT 57.875 175.525 58.165 175.570 ;
        RECT 58.320 175.510 58.640 175.570 ;
        RECT 58.780 175.510 59.100 175.770 ;
        RECT 61.540 175.710 61.860 175.770 ;
        RECT 62.475 175.710 62.765 175.755 ;
        RECT 61.540 175.570 62.765 175.710 ;
        RECT 61.540 175.510 61.860 175.570 ;
        RECT 62.475 175.525 62.765 175.570 ;
        RECT 65.680 175.510 66.000 175.770 ;
        RECT 68.440 175.510 68.760 175.770 ;
        RECT 68.990 175.755 69.130 175.910 ;
        RECT 68.915 175.525 69.205 175.755 ;
        RECT 69.360 175.510 69.680 175.770 ;
        RECT 70.295 175.525 70.585 175.755 ;
        RECT 56.480 175.170 56.800 175.430 ;
        RECT 70.370 175.370 70.510 175.525 ;
        RECT 72.120 175.510 72.440 175.770 ;
        RECT 72.670 175.755 72.810 175.910 ;
        RECT 73.500 175.850 73.820 175.910 ;
        RECT 72.595 175.525 72.885 175.755 ;
        RECT 73.040 175.510 73.360 175.770 ;
        RECT 73.975 175.525 74.265 175.755 ;
        RECT 74.420 175.710 74.740 175.770 ;
        RECT 76.810 175.755 76.950 176.250 ;
        RECT 81.795 176.250 90.290 176.390 ;
        RECT 81.795 176.205 82.085 176.250 ;
        RECT 83.160 176.050 83.480 176.110 ;
        RECT 83.635 176.050 83.925 176.095 ;
        RECT 83.160 175.910 83.925 176.050 ;
        RECT 83.160 175.850 83.480 175.910 ;
        RECT 83.635 175.865 83.925 175.910 ;
        RECT 84.080 176.050 84.400 176.110 ;
        RECT 85.915 176.050 86.565 176.095 ;
        RECT 89.515 176.050 89.805 176.095 ;
        RECT 84.080 175.910 89.805 176.050 ;
        RECT 84.080 175.850 84.400 175.910 ;
        RECT 85.915 175.865 86.565 175.910 ;
        RECT 89.215 175.865 89.805 175.910 ;
        RECT 76.275 175.710 76.565 175.755 ;
        RECT 74.420 175.570 76.565 175.710 ;
        RECT 74.050 175.370 74.190 175.525 ;
        RECT 74.420 175.510 74.740 175.570 ;
        RECT 76.275 175.525 76.565 175.570 ;
        RECT 76.735 175.525 77.025 175.755 ;
        RECT 77.195 175.710 77.485 175.755 ;
        RECT 77.640 175.710 77.960 175.770 ;
        RECT 77.195 175.570 77.960 175.710 ;
        RECT 77.195 175.525 77.485 175.570 ;
        RECT 77.640 175.510 77.960 175.570 ;
        RECT 78.115 175.525 78.405 175.755 ;
        RECT 79.035 175.710 79.325 175.755 ;
        RECT 80.400 175.710 80.720 175.770 ;
        RECT 79.035 175.570 80.720 175.710 ;
        RECT 79.035 175.525 79.325 175.570 ;
        RECT 74.880 175.370 75.200 175.430 ;
        RECT 78.190 175.370 78.330 175.525 ;
        RECT 80.400 175.510 80.720 175.570 ;
        RECT 82.720 175.710 83.010 175.755 ;
        RECT 84.555 175.710 84.845 175.755 ;
        RECT 88.135 175.710 88.425 175.755 ;
        RECT 82.720 175.570 88.425 175.710 ;
        RECT 82.720 175.525 83.010 175.570 ;
        RECT 84.555 175.525 84.845 175.570 ;
        RECT 88.135 175.525 88.425 175.570 ;
        RECT 89.215 175.550 89.505 175.865 ;
        RECT 90.150 175.710 90.290 176.250 ;
        RECT 91.440 176.190 91.760 176.450 ;
        RECT 94.660 176.050 94.980 176.110 ;
        RECT 96.500 176.050 96.820 176.110 ;
        RECT 94.660 175.910 96.820 176.050 ;
        RECT 94.660 175.850 94.980 175.910 ;
        RECT 92.375 175.710 92.665 175.755 ;
        RECT 90.150 175.570 92.665 175.710 ;
        RECT 92.375 175.525 92.665 175.570 ;
        RECT 93.280 175.710 93.600 175.770 ;
        RECT 95.120 175.710 95.440 175.770 ;
        RECT 95.670 175.755 95.810 175.910 ;
        RECT 96.500 175.850 96.820 175.910 ;
        RECT 99.720 176.050 100.040 176.110 ;
        RECT 103.975 176.050 104.265 176.095 ;
        RECT 107.215 176.050 107.865 176.095 ;
        RECT 99.720 175.910 107.865 176.050 ;
        RECT 99.720 175.850 100.040 175.910 ;
        RECT 103.975 175.865 104.565 175.910 ;
        RECT 107.215 175.865 107.865 175.910 ;
        RECT 93.280 175.570 95.440 175.710 ;
        RECT 93.280 175.510 93.600 175.570 ;
        RECT 95.120 175.510 95.440 175.570 ;
        RECT 95.595 175.525 95.885 175.755 ;
        RECT 96.055 175.525 96.345 175.755 ;
        RECT 64.850 175.230 78.330 175.370 ;
        RECT 82.255 175.370 82.545 175.415 ;
        RECT 83.620 175.370 83.940 175.430 ;
        RECT 82.255 175.230 83.940 175.370 ;
        RECT 51.995 175.030 52.285 175.075 ;
        RECT 55.115 175.030 55.405 175.075 ;
        RECT 57.005 175.030 57.295 175.075 ;
        RECT 51.995 174.890 57.295 175.030 ;
        RECT 51.995 174.845 52.285 174.890 ;
        RECT 55.115 174.845 55.405 174.890 ;
        RECT 57.005 174.845 57.295 174.890 ;
        RECT 64.850 174.735 64.990 175.230 ;
        RECT 74.880 175.170 75.200 175.230 ;
        RECT 82.255 175.185 82.545 175.230 ;
        RECT 83.620 175.170 83.940 175.230 ;
        RECT 85.920 175.370 86.240 175.430 ;
        RECT 96.130 175.370 96.270 175.525 ;
        RECT 96.960 175.510 97.280 175.770 ;
        RECT 104.275 175.550 104.565 175.865 ;
        RECT 105.355 175.710 105.645 175.755 ;
        RECT 108.935 175.710 109.225 175.755 ;
        RECT 110.770 175.710 111.060 175.755 ;
        RECT 105.355 175.570 111.060 175.710 ;
        RECT 105.355 175.525 105.645 175.570 ;
        RECT 108.935 175.525 109.225 175.570 ;
        RECT 110.770 175.525 111.060 175.570 ;
        RECT 85.920 175.230 96.270 175.370 ;
        RECT 106.620 175.370 106.940 175.430 ;
        RECT 109.855 175.370 110.145 175.415 ;
        RECT 106.620 175.230 110.145 175.370 ;
        RECT 85.920 175.170 86.240 175.230 ;
        RECT 106.620 175.170 106.940 175.230 ;
        RECT 109.855 175.185 110.145 175.230 ;
        RECT 111.220 175.170 111.540 175.430 ;
        RECT 83.125 175.030 83.415 175.075 ;
        RECT 85.015 175.030 85.305 175.075 ;
        RECT 88.135 175.030 88.425 175.075 ;
        RECT 83.125 174.890 88.425 175.030 ;
        RECT 83.125 174.845 83.415 174.890 ;
        RECT 85.015 174.845 85.305 174.890 ;
        RECT 88.135 174.845 88.425 174.890 ;
        RECT 105.355 175.030 105.645 175.075 ;
        RECT 108.475 175.030 108.765 175.075 ;
        RECT 110.365 175.030 110.655 175.075 ;
        RECT 105.355 174.890 110.655 175.030 ;
        RECT 105.355 174.845 105.645 174.890 ;
        RECT 108.475 174.845 108.765 174.890 ;
        RECT 110.365 174.845 110.655 174.890 ;
        RECT 64.775 174.690 65.065 174.735 ;
        RECT 45.440 174.550 65.065 174.690 ;
        RECT 45.440 174.490 45.760 174.550 ;
        RECT 64.775 174.505 65.065 174.550 ;
        RECT 67.060 174.490 67.380 174.750 ;
        RECT 70.740 174.490 71.060 174.750 ;
        RECT 72.120 174.690 72.440 174.750 ;
        RECT 74.895 174.690 75.185 174.735 ;
        RECT 72.120 174.550 75.185 174.690 ;
        RECT 72.120 174.490 72.440 174.550 ;
        RECT 74.895 174.505 75.185 174.550 ;
        RECT 89.600 174.690 89.920 174.750 ;
        RECT 90.995 174.690 91.285 174.735 ;
        RECT 89.600 174.550 91.285 174.690 ;
        RECT 89.600 174.490 89.920 174.550 ;
        RECT 90.995 174.505 91.285 174.550 ;
        RECT 93.755 174.690 94.045 174.735 ;
        RECT 95.120 174.690 95.440 174.750 ;
        RECT 93.755 174.550 95.440 174.690 ;
        RECT 93.755 174.505 94.045 174.550 ;
        RECT 95.120 174.490 95.440 174.550 ;
        RECT 102.495 174.690 102.785 174.735 ;
        RECT 103.400 174.690 103.720 174.750 ;
        RECT 102.495 174.550 103.720 174.690 ;
        RECT 135.635 174.550 136.775 223.880 ;
        RECT 138.130 223.810 139.580 225.110 ;
        RECT 143.180 223.840 144.630 225.140 ;
        RECT 102.495 174.505 102.785 174.550 ;
        RECT 103.400 174.490 103.720 174.550 ;
        RECT 15.010 173.870 113.450 174.350 ;
        RECT 39.000 173.670 39.320 173.730 ;
        RECT 41.300 173.670 41.620 173.730 ;
        RECT 39.000 173.530 41.620 173.670 ;
        RECT 39.000 173.470 39.320 173.530 ;
        RECT 41.300 173.470 41.620 173.530 ;
        RECT 51.880 173.470 52.200 173.730 ;
        RECT 52.800 173.670 53.120 173.730 ;
        RECT 82.255 173.670 82.545 173.715 ;
        RECT 84.080 173.670 84.400 173.730 ;
        RECT 96.960 173.670 97.280 173.730 ;
        RECT 98.340 173.670 98.660 173.730 ;
        RECT 52.800 173.530 60.850 173.670 ;
        RECT 52.800 173.470 53.120 173.530 ;
        RECT 23.015 173.330 23.305 173.375 ;
        RECT 26.135 173.330 26.425 173.375 ;
        RECT 28.025 173.330 28.315 173.375 ;
        RECT 23.015 173.190 28.315 173.330 ;
        RECT 23.015 173.145 23.305 173.190 ;
        RECT 26.135 173.145 26.425 173.190 ;
        RECT 28.025 173.145 28.315 173.190 ;
        RECT 29.355 173.330 29.645 173.375 ;
        RECT 29.800 173.330 30.120 173.390 ;
        RECT 29.355 173.190 30.120 173.330 ;
        RECT 29.355 173.145 29.645 173.190 ;
        RECT 29.800 173.130 30.120 173.190 ;
        RECT 31.180 173.330 31.500 173.390 ;
        RECT 55.215 173.330 55.505 173.375 ;
        RECT 58.335 173.330 58.625 173.375 ;
        RECT 60.225 173.330 60.515 173.375 ;
        RECT 31.180 173.190 32.330 173.330 ;
        RECT 31.180 173.130 31.500 173.190 ;
        RECT 20.140 172.790 20.460 173.050 ;
        RECT 24.740 172.990 25.060 173.050 ;
        RECT 27.515 172.990 27.805 173.035 ;
        RECT 24.740 172.850 27.805 172.990 ;
        RECT 24.740 172.790 25.060 172.850 ;
        RECT 27.515 172.805 27.805 172.850 ;
        RECT 30.260 172.990 30.580 173.050 ;
        RECT 32.190 173.035 32.330 173.190 ;
        RECT 40.930 173.190 53.030 173.330 ;
        RECT 31.655 172.990 31.945 173.035 ;
        RECT 30.260 172.850 31.945 172.990 ;
        RECT 30.260 172.790 30.580 172.850 ;
        RECT 31.655 172.805 31.945 172.850 ;
        RECT 32.115 172.805 32.405 173.035 ;
        RECT 16.920 172.450 17.240 172.710 ;
        RECT 18.300 172.310 18.620 172.370 ;
        RECT 21.935 172.355 22.225 172.670 ;
        RECT 23.015 172.650 23.305 172.695 ;
        RECT 26.595 172.650 26.885 172.695 ;
        RECT 28.430 172.650 28.720 172.695 ;
        RECT 23.015 172.510 28.720 172.650 ;
        RECT 23.015 172.465 23.305 172.510 ;
        RECT 26.595 172.465 26.885 172.510 ;
        RECT 28.430 172.465 28.720 172.510 ;
        RECT 28.895 172.650 29.185 172.695 ;
        RECT 29.340 172.650 29.660 172.710 ;
        RECT 28.895 172.510 29.660 172.650 ;
        RECT 28.895 172.465 29.185 172.510 ;
        RECT 29.340 172.450 29.660 172.510 ;
        RECT 37.160 172.450 37.480 172.710 ;
        RECT 39.015 172.465 39.305 172.695 ;
        RECT 21.635 172.310 22.225 172.355 ;
        RECT 24.875 172.310 25.525 172.355 ;
        RECT 18.300 172.170 25.525 172.310 ;
        RECT 39.090 172.310 39.230 172.465 ;
        RECT 39.460 172.450 39.780 172.710 ;
        RECT 39.920 172.450 40.240 172.710 ;
        RECT 40.930 172.695 41.070 173.190 ;
        RECT 45.440 172.990 45.760 173.050 ;
        RECT 49.135 172.990 49.425 173.035 ;
        RECT 52.355 172.990 52.645 173.035 ;
        RECT 43.230 172.850 45.760 172.990 ;
        RECT 43.230 172.695 43.370 172.850 ;
        RECT 45.440 172.790 45.760 172.850 ;
        RECT 45.990 172.850 52.645 172.990 ;
        RECT 52.890 172.990 53.030 173.190 ;
        RECT 55.215 173.190 60.515 173.330 ;
        RECT 60.710 173.330 60.850 173.530 ;
        RECT 70.600 173.530 82.010 173.670 ;
        RECT 70.600 173.330 70.740 173.530 ;
        RECT 60.710 173.190 63.150 173.330 ;
        RECT 55.215 173.145 55.505 173.190 ;
        RECT 58.335 173.145 58.625 173.190 ;
        RECT 60.225 173.145 60.515 173.190 ;
        RECT 59.240 172.990 59.560 173.050 ;
        RECT 52.890 172.850 59.560 172.990 ;
        RECT 40.855 172.465 41.145 172.695 ;
        RECT 42.695 172.465 42.985 172.695 ;
        RECT 43.155 172.465 43.445 172.695 ;
        RECT 42.770 172.310 42.910 172.465 ;
        RECT 43.600 172.450 43.920 172.710 ;
        RECT 44.535 172.650 44.825 172.695 ;
        RECT 44.980 172.650 45.300 172.710 ;
        RECT 45.990 172.695 46.130 172.850 ;
        RECT 49.135 172.805 49.425 172.850 ;
        RECT 52.355 172.805 52.645 172.850 ;
        RECT 59.240 172.790 59.560 172.850 ;
        RECT 59.700 172.790 60.020 173.050 ;
        RECT 44.535 172.510 45.300 172.650 ;
        RECT 44.535 172.465 44.825 172.510 ;
        RECT 44.980 172.450 45.300 172.510 ;
        RECT 45.915 172.465 46.205 172.695 ;
        RECT 46.360 172.450 46.680 172.710 ;
        RECT 46.820 172.450 47.140 172.710 ;
        RECT 63.010 172.695 63.150 173.190 ;
        RECT 65.310 173.190 70.740 173.330 ;
        RECT 72.600 173.330 72.890 173.375 ;
        RECT 74.460 173.330 74.750 173.375 ;
        RECT 77.240 173.330 77.530 173.375 ;
        RECT 72.600 173.190 77.530 173.330 ;
        RECT 81.870 173.330 82.010 173.530 ;
        RECT 82.255 173.530 84.400 173.670 ;
        RECT 82.255 173.485 82.545 173.530 ;
        RECT 84.080 173.470 84.400 173.530 ;
        RECT 91.530 173.530 98.660 173.670 ;
        RECT 91.530 173.330 91.670 173.530 ;
        RECT 96.960 173.470 97.280 173.530 ;
        RECT 98.340 173.470 98.660 173.530 ;
        RECT 99.720 173.470 100.040 173.730 ;
        RECT 135.580 173.430 136.830 174.550 ;
        RECT 135.635 173.420 136.775 173.430 ;
        RECT 102.020 173.330 102.340 173.390 ;
        RECT 81.870 173.190 91.670 173.330 ;
        RECT 46.910 172.310 47.050 172.450 ;
        RECT 54.135 172.355 54.425 172.670 ;
        RECT 55.215 172.650 55.505 172.695 ;
        RECT 58.795 172.650 59.085 172.695 ;
        RECT 60.630 172.650 60.920 172.695 ;
        RECT 55.215 172.510 60.920 172.650 ;
        RECT 55.215 172.465 55.505 172.510 ;
        RECT 58.795 172.465 59.085 172.510 ;
        RECT 60.630 172.465 60.920 172.510 ;
        RECT 61.095 172.465 61.385 172.695 ;
        RECT 62.935 172.465 63.225 172.695 ;
        RECT 57.400 172.355 57.720 172.370 ;
        RECT 39.090 172.170 47.050 172.310 ;
        RECT 53.835 172.310 54.425 172.355 ;
        RECT 57.075 172.310 57.725 172.355 ;
        RECT 53.835 172.170 57.725 172.310 ;
        RECT 18.300 172.110 18.620 172.170 ;
        RECT 21.635 172.125 21.925 172.170 ;
        RECT 24.875 172.125 25.525 172.170 ;
        RECT 53.835 172.125 54.125 172.170 ;
        RECT 57.075 172.125 57.725 172.170 ;
        RECT 58.320 172.310 58.640 172.370 ;
        RECT 61.170 172.310 61.310 172.465 ;
        RECT 58.320 172.170 61.310 172.310 ;
        RECT 57.400 172.110 57.720 172.125 ;
        RECT 58.320 172.110 58.640 172.170 ;
        RECT 65.310 172.030 65.450 173.190 ;
        RECT 72.600 173.145 72.890 173.190 ;
        RECT 74.460 173.145 74.750 173.190 ;
        RECT 77.240 173.145 77.530 173.190 ;
        RECT 69.820 172.990 70.140 173.050 ;
        RECT 73.975 172.990 74.265 173.035 ;
        RECT 83.620 172.990 83.940 173.050 ;
        RECT 69.820 172.850 74.265 172.990 ;
        RECT 69.820 172.790 70.140 172.850 ;
        RECT 73.975 172.805 74.265 172.850 ;
        RECT 74.510 172.850 83.940 172.990 ;
        RECT 65.680 172.450 66.000 172.710 ;
        RECT 72.135 172.650 72.425 172.695 ;
        RECT 74.510 172.650 74.650 172.850 ;
        RECT 83.620 172.790 83.940 172.850 ;
        RECT 84.080 172.790 84.400 173.050 ;
        RECT 77.240 172.650 77.530 172.695 ;
        RECT 72.135 172.510 74.650 172.650 ;
        RECT 74.995 172.510 77.530 172.650 ;
        RECT 72.135 172.465 72.425 172.510 ;
        RECT 74.995 172.355 75.210 172.510 ;
        RECT 77.240 172.465 77.530 172.510 ;
        RECT 81.795 172.650 82.085 172.695 ;
        RECT 85.000 172.650 85.320 172.710 ;
        RECT 81.795 172.510 85.320 172.650 ;
        RECT 81.795 172.465 82.085 172.510 ;
        RECT 85.000 172.450 85.320 172.510 ;
        RECT 89.600 172.650 89.920 172.710 ;
        RECT 91.530 172.695 91.670 173.190 ;
        RECT 92.345 173.190 102.340 173.330 ;
        RECT 92.345 172.695 92.485 173.190 ;
        RECT 102.020 173.130 102.340 173.190 ;
        RECT 104.895 173.330 105.185 173.375 ;
        RECT 108.015 173.330 108.305 173.375 ;
        RECT 109.905 173.330 110.195 173.375 ;
        RECT 104.895 173.190 110.195 173.330 ;
        RECT 104.895 173.145 105.185 173.190 ;
        RECT 108.015 173.145 108.305 173.190 ;
        RECT 109.905 173.145 110.195 173.190 ;
        RECT 94.200 172.990 94.520 173.050 ;
        RECT 92.910 172.850 94.520 172.990 ;
        RECT 92.910 172.695 93.050 172.850 ;
        RECT 94.200 172.790 94.520 172.850 ;
        RECT 94.660 172.990 94.980 173.050 ;
        RECT 95.135 172.990 95.425 173.035 ;
        RECT 94.660 172.850 95.425 172.990 ;
        RECT 94.660 172.790 94.980 172.850 ;
        RECT 95.135 172.805 95.425 172.850 ;
        RECT 95.580 172.990 95.900 173.050 ;
        RECT 95.580 172.850 97.650 172.990 ;
        RECT 95.580 172.790 95.900 172.850 ;
        RECT 90.535 172.650 90.825 172.695 ;
        RECT 89.600 172.510 90.825 172.650 ;
        RECT 89.600 172.450 89.920 172.510 ;
        RECT 90.535 172.465 90.825 172.510 ;
        RECT 91.455 172.465 91.745 172.695 ;
        RECT 92.345 172.520 92.665 172.695 ;
        RECT 92.375 172.465 92.665 172.520 ;
        RECT 92.835 172.465 93.125 172.695 ;
        RECT 93.280 172.650 93.600 172.710 ;
        RECT 96.515 172.650 96.805 172.695 ;
        RECT 93.280 172.510 96.805 172.650 ;
        RECT 93.280 172.450 93.600 172.510 ;
        RECT 96.515 172.465 96.805 172.510 ;
        RECT 96.960 172.450 97.280 172.710 ;
        RECT 97.510 172.695 97.650 172.850 ;
        RECT 97.435 172.465 97.725 172.695 ;
        RECT 98.340 172.450 98.660 172.710 ;
        RECT 98.800 172.650 99.120 172.710 ;
        RECT 99.275 172.650 99.565 172.695 ;
        RECT 100.640 172.650 100.960 172.710 ;
        RECT 98.800 172.510 100.960 172.650 ;
        RECT 98.800 172.450 99.120 172.510 ;
        RECT 99.275 172.465 99.565 172.510 ;
        RECT 100.640 172.450 100.960 172.510 ;
        RECT 73.060 172.310 73.350 172.355 ;
        RECT 74.920 172.310 75.210 172.355 ;
        RECT 75.840 172.310 76.130 172.355 ;
        RECT 79.100 172.310 79.390 172.355 ;
        RECT 73.060 172.170 75.210 172.310 ;
        RECT 73.060 172.125 73.350 172.170 ;
        RECT 74.920 172.125 75.210 172.170 ;
        RECT 75.430 172.170 79.390 172.310 ;
        RECT 19.695 171.970 19.985 172.015 ;
        RECT 20.600 171.970 20.920 172.030 ;
        RECT 19.695 171.830 20.920 171.970 ;
        RECT 19.695 171.785 19.985 171.830 ;
        RECT 20.600 171.770 20.920 171.830 ;
        RECT 28.880 171.970 29.200 172.030 ;
        RECT 31.195 171.970 31.485 172.015 ;
        RECT 28.880 171.830 31.485 171.970 ;
        RECT 28.880 171.770 29.200 171.830 ;
        RECT 31.195 171.785 31.485 171.830 ;
        RECT 31.640 171.970 31.960 172.030 ;
        RECT 36.715 171.970 37.005 172.015 ;
        RECT 31.640 171.830 37.005 171.970 ;
        RECT 31.640 171.770 31.960 171.830 ;
        RECT 36.715 171.785 37.005 171.830 ;
        RECT 37.635 171.970 37.925 172.015 ;
        RECT 38.540 171.970 38.860 172.030 ;
        RECT 37.635 171.830 38.860 171.970 ;
        RECT 37.635 171.785 37.925 171.830 ;
        RECT 38.540 171.770 38.860 171.830 ;
        RECT 41.300 171.770 41.620 172.030 ;
        RECT 48.215 171.970 48.505 172.015 ;
        RECT 50.040 171.970 50.360 172.030 ;
        RECT 48.215 171.830 50.360 171.970 ;
        RECT 48.215 171.785 48.505 171.830 ;
        RECT 50.040 171.770 50.360 171.830 ;
        RECT 56.480 171.970 56.800 172.030 ;
        RECT 62.015 171.970 62.305 172.015 ;
        RECT 56.480 171.830 62.305 171.970 ;
        RECT 56.480 171.770 56.800 171.830 ;
        RECT 62.015 171.785 62.305 171.830 ;
        RECT 64.775 171.970 65.065 172.015 ;
        RECT 65.220 171.970 65.540 172.030 ;
        RECT 64.775 171.830 65.540 171.970 ;
        RECT 64.775 171.785 65.065 171.830 ;
        RECT 65.220 171.770 65.540 171.830 ;
        RECT 67.980 171.970 68.300 172.030 ;
        RECT 75.430 171.970 75.570 172.170 ;
        RECT 75.840 172.125 76.130 172.170 ;
        RECT 79.100 172.125 79.390 172.170 ;
        RECT 84.555 172.310 84.845 172.355 ;
        RECT 94.675 172.310 94.965 172.355 ;
        RECT 96.040 172.310 96.360 172.370 ;
        RECT 103.815 172.355 104.105 172.670 ;
        RECT 104.895 172.650 105.185 172.695 ;
        RECT 108.475 172.650 108.765 172.695 ;
        RECT 110.310 172.650 110.600 172.695 ;
        RECT 104.895 172.510 110.600 172.650 ;
        RECT 104.895 172.465 105.185 172.510 ;
        RECT 108.475 172.465 108.765 172.510 ;
        RECT 110.310 172.465 110.600 172.510 ;
        RECT 110.760 172.450 111.080 172.710 ;
        RECT 84.555 172.170 87.990 172.310 ;
        RECT 84.555 172.125 84.845 172.170 ;
        RECT 67.980 171.830 75.570 171.970 ;
        RECT 77.180 171.970 77.500 172.030 ;
        RECT 81.105 171.970 81.395 172.015 ;
        RECT 85.015 171.970 85.305 172.015 ;
        RECT 77.180 171.830 85.305 171.970 ;
        RECT 67.980 171.770 68.300 171.830 ;
        RECT 77.180 171.770 77.500 171.830 ;
        RECT 81.105 171.785 81.395 171.830 ;
        RECT 85.015 171.785 85.305 171.830 ;
        RECT 86.840 171.770 87.160 172.030 ;
        RECT 87.850 172.015 87.990 172.170 ;
        RECT 94.675 172.170 96.360 172.310 ;
        RECT 94.675 172.125 94.965 172.170 ;
        RECT 96.040 172.110 96.360 172.170 ;
        RECT 101.115 172.310 101.405 172.355 ;
        RECT 103.515 172.310 104.105 172.355 ;
        RECT 106.755 172.310 107.405 172.355 ;
        RECT 101.115 172.170 107.405 172.310 ;
        RECT 101.115 172.125 101.405 172.170 ;
        RECT 103.515 172.125 103.805 172.170 ;
        RECT 106.755 172.125 107.405 172.170 ;
        RECT 109.380 172.110 109.700 172.370 ;
        RECT 133.700 172.190 134.930 172.680 ;
        RECT 87.775 171.970 88.065 172.015 ;
        RECT 97.880 171.970 98.200 172.030 ;
        RECT 87.775 171.830 98.200 171.970 ;
        RECT 87.775 171.785 88.065 171.830 ;
        RECT 97.880 171.770 98.200 171.830 ;
        RECT 102.020 171.770 102.340 172.030 ;
        RECT 133.700 171.930 136.690 172.190 ;
        RECT 138.330 171.930 139.470 223.810 ;
        RECT 15.010 171.150 113.450 171.630 ;
        RECT 18.300 170.750 18.620 171.010 ;
        RECT 28.880 170.750 29.200 171.010 ;
        RECT 39.000 170.950 39.320 171.010 ;
        RECT 30.810 170.810 39.320 170.950 ;
        RECT 19.680 170.410 20.000 170.670 ;
        RECT 21.060 170.410 21.380 170.670 ;
        RECT 21.980 170.610 22.300 170.670 ;
        RECT 21.980 170.410 22.440 170.610 ;
        RECT 18.775 170.270 19.065 170.315 ;
        RECT 19.770 170.270 19.910 170.410 ;
        RECT 21.150 170.270 21.290 170.410 ;
        RECT 18.775 170.130 21.290 170.270 ;
        RECT 18.775 170.085 19.065 170.130 ;
        RECT 19.695 169.930 19.985 169.975 ;
        RECT 21.060 169.930 21.380 169.990 ;
        RECT 19.695 169.790 21.380 169.930 ;
        RECT 19.695 169.745 19.985 169.790 ;
        RECT 21.060 169.730 21.380 169.790 ;
        RECT 22.300 169.590 22.440 170.410 ;
        RECT 26.135 170.270 26.425 170.315 ;
        RECT 26.580 170.270 26.900 170.330 ;
        RECT 26.135 170.130 26.900 170.270 ;
        RECT 26.135 170.085 26.425 170.130 ;
        RECT 26.580 170.070 26.900 170.130 ;
        RECT 30.810 169.930 30.950 170.810 ;
        RECT 31.655 170.085 31.945 170.315 ;
        RECT 31.730 169.930 31.870 170.085 ;
        RECT 32.100 170.070 32.420 170.330 ;
        RECT 32.560 170.070 32.880 170.330 ;
        RECT 33.480 170.070 33.800 170.330 ;
        RECT 35.410 170.315 35.550 170.810 ;
        RECT 39.000 170.750 39.320 170.810 ;
        RECT 40.840 170.750 41.160 171.010 ;
        RECT 57.400 170.950 57.720 171.010 ;
        RECT 57.875 170.950 58.165 170.995 ;
        RECT 57.400 170.810 58.165 170.950 ;
        RECT 57.400 170.750 57.720 170.810 ;
        RECT 57.875 170.765 58.165 170.810 ;
        RECT 59.240 170.950 59.560 171.010 ;
        RECT 63.395 170.950 63.685 170.995 ;
        RECT 59.240 170.810 63.685 170.950 ;
        RECT 59.240 170.750 59.560 170.810 ;
        RECT 63.395 170.765 63.685 170.810 ;
        RECT 67.980 170.750 68.300 171.010 ;
        RECT 69.820 170.750 70.140 171.010 ;
        RECT 83.160 170.950 83.480 171.010 ;
        RECT 87.775 170.950 88.065 170.995 ;
        RECT 83.160 170.810 88.065 170.950 ;
        RECT 83.160 170.750 83.480 170.810 ;
        RECT 87.775 170.765 88.065 170.810 ;
        RECT 89.140 170.950 89.460 171.010 ;
        RECT 94.660 170.950 94.980 171.010 ;
        RECT 89.140 170.810 94.980 170.950 ;
        RECT 89.140 170.750 89.460 170.810 ;
        RECT 94.660 170.750 94.980 170.810 ;
        RECT 97.880 170.750 98.200 171.010 ;
        RECT 106.620 170.750 106.940 171.010 ;
        RECT 108.015 170.950 108.305 170.995 ;
        RECT 109.380 170.950 109.700 171.010 ;
        RECT 108.015 170.810 109.700 170.950 ;
        RECT 108.015 170.765 108.305 170.810 ;
        RECT 109.380 170.750 109.700 170.810 ;
        RECT 133.700 170.790 139.470 171.930 ;
        RECT 36.700 170.610 37.020 170.670 ;
        RECT 40.930 170.610 41.070 170.750 ;
        RECT 65.680 170.610 66.000 170.670 ;
        RECT 79.480 170.610 79.800 170.670 ;
        RECT 36.700 170.470 40.150 170.610 ;
        RECT 36.700 170.410 37.020 170.470 ;
        RECT 35.335 170.085 35.625 170.315 ;
        RECT 35.795 170.085 36.085 170.315 ;
        RECT 30.810 169.790 31.870 169.930 ;
        RECT 33.020 169.930 33.340 169.990 ;
        RECT 33.020 169.790 33.710 169.930 ;
        RECT 33.020 169.730 33.340 169.790 ;
        RECT 32.100 169.590 32.420 169.650 ;
        RECT 22.300 169.450 32.420 169.590 ;
        RECT 33.570 169.590 33.710 169.790 ;
        RECT 33.940 169.730 34.260 169.990 ;
        RECT 35.870 169.930 36.010 170.085 ;
        RECT 36.240 170.070 36.560 170.330 ;
        RECT 37.175 170.270 37.465 170.315 ;
        RECT 38.080 170.270 38.400 170.330 ;
        RECT 37.175 170.130 38.400 170.270 ;
        RECT 37.175 170.085 37.465 170.130 ;
        RECT 38.080 170.070 38.400 170.130 ;
        RECT 39.000 170.070 39.320 170.330 ;
        RECT 40.010 170.315 40.150 170.470 ;
        RECT 40.470 170.470 41.070 170.610 ;
        RECT 64.390 170.470 66.000 170.610 ;
        RECT 39.475 170.085 39.765 170.315 ;
        RECT 39.935 170.085 40.225 170.315 ;
        RECT 39.550 169.930 39.690 170.085 ;
        RECT 40.470 169.930 40.610 170.470 ;
        RECT 40.855 170.085 41.145 170.315 ;
        RECT 35.870 169.790 40.610 169.930 ;
        RECT 35.870 169.590 36.010 169.790 ;
        RECT 33.570 169.450 36.010 169.590 ;
        RECT 32.100 169.390 32.420 169.450 ;
        RECT 37.620 169.390 37.940 169.650 ;
        RECT 38.080 169.590 38.400 169.650 ;
        RECT 40.930 169.590 41.070 170.085 ;
        RECT 42.220 170.070 42.540 170.330 ;
        RECT 46.375 170.270 46.665 170.315 ;
        RECT 49.580 170.270 49.900 170.330 ;
        RECT 46.375 170.130 49.900 170.270 ;
        RECT 46.375 170.085 46.665 170.130 ;
        RECT 49.580 170.070 49.900 170.130 ;
        RECT 52.815 170.270 53.105 170.315 ;
        RECT 53.260 170.270 53.580 170.330 ;
        RECT 57.860 170.270 58.180 170.330 ;
        RECT 52.815 170.130 58.180 170.270 ;
        RECT 52.815 170.085 53.105 170.130 ;
        RECT 53.260 170.070 53.580 170.130 ;
        RECT 57.860 170.070 58.180 170.130 ;
        RECT 58.335 170.270 58.625 170.315 ;
        RECT 58.780 170.270 59.100 170.330 ;
        RECT 58.335 170.130 59.100 170.270 ;
        RECT 58.335 170.085 58.625 170.130 ;
        RECT 58.780 170.070 59.100 170.130 ;
        RECT 63.380 170.270 63.700 170.330 ;
        RECT 64.390 170.315 64.530 170.470 ;
        RECT 65.680 170.410 66.000 170.470 ;
        RECT 68.530 170.470 79.800 170.610 ;
        RECT 64.315 170.270 64.605 170.315 ;
        RECT 63.380 170.130 64.605 170.270 ;
        RECT 63.380 170.070 63.700 170.130 ;
        RECT 64.315 170.085 64.605 170.130 ;
        RECT 64.760 170.270 65.080 170.330 ;
        RECT 68.530 170.315 68.670 170.470 ;
        RECT 79.480 170.410 79.800 170.470 ;
        RECT 97.435 170.610 97.725 170.655 ;
        RECT 99.260 170.610 99.580 170.670 ;
        RECT 103.415 170.610 103.705 170.655 ;
        RECT 97.435 170.470 103.705 170.610 ;
        RECT 97.435 170.425 97.725 170.470 ;
        RECT 99.260 170.410 99.580 170.470 ;
        RECT 103.415 170.425 103.705 170.470 ;
        RECT 133.700 170.600 136.690 170.790 ;
        RECT 65.235 170.270 65.525 170.315 ;
        RECT 64.760 170.130 65.525 170.270 ;
        RECT 64.760 170.070 65.080 170.130 ;
        RECT 65.235 170.085 65.525 170.130 ;
        RECT 68.455 170.085 68.745 170.315 ;
        RECT 68.915 170.270 69.205 170.315 ;
        RECT 71.660 170.270 71.980 170.330 ;
        RECT 72.135 170.270 72.425 170.315 ;
        RECT 77.180 170.270 77.500 170.330 ;
        RECT 68.915 170.130 70.510 170.270 ;
        RECT 68.915 170.085 69.205 170.130 ;
        RECT 42.680 169.930 43.000 169.990 ;
        RECT 46.835 169.930 47.125 169.975 ;
        RECT 42.680 169.790 47.125 169.930 ;
        RECT 42.680 169.730 43.000 169.790 ;
        RECT 46.835 169.745 47.125 169.790 ;
        RECT 47.280 169.730 47.600 169.990 ;
        RECT 65.220 169.590 65.540 169.650 ;
        RECT 70.370 169.635 70.510 170.130 ;
        RECT 71.660 170.130 72.425 170.270 ;
        RECT 71.660 170.070 71.980 170.130 ;
        RECT 72.135 170.085 72.425 170.130 ;
        RECT 73.130 170.130 77.500 170.270 ;
        RECT 73.130 169.990 73.270 170.130 ;
        RECT 77.180 170.070 77.500 170.130 ;
        RECT 83.620 170.270 83.940 170.330 ;
        RECT 84.555 170.270 84.845 170.315 ;
        RECT 83.620 170.130 84.845 170.270 ;
        RECT 83.620 170.070 83.940 170.130 ;
        RECT 84.555 170.085 84.845 170.130 ;
        RECT 86.840 170.270 87.160 170.330 ;
        RECT 88.695 170.270 88.985 170.315 ;
        RECT 86.840 170.130 88.985 170.270 ;
        RECT 86.840 170.070 87.160 170.130 ;
        RECT 88.695 170.085 88.985 170.130 ;
        RECT 94.675 170.270 94.965 170.315 ;
        RECT 98.800 170.270 99.120 170.330 ;
        RECT 105.715 170.270 106.005 170.315 ;
        RECT 94.675 170.130 99.120 170.270 ;
        RECT 94.675 170.085 94.965 170.130 ;
        RECT 98.800 170.070 99.120 170.130 ;
        RECT 99.810 170.130 106.005 170.270 ;
        RECT 72.595 169.930 72.885 169.975 ;
        RECT 73.040 169.930 73.360 169.990 ;
        RECT 72.595 169.790 73.360 169.930 ;
        RECT 72.595 169.745 72.885 169.790 ;
        RECT 73.040 169.730 73.360 169.790 ;
        RECT 73.515 169.745 73.805 169.975 ;
        RECT 38.080 169.450 65.540 169.590 ;
        RECT 38.080 169.390 38.400 169.450 ;
        RECT 65.220 169.390 65.540 169.450 ;
        RECT 70.295 169.405 70.585 169.635 ;
        RECT 73.590 169.590 73.730 169.745 ;
        RECT 96.960 169.730 97.280 169.990 ;
        RECT 99.810 169.635 99.950 170.130 ;
        RECT 105.715 170.085 106.005 170.130 ;
        RECT 107.095 170.085 107.385 170.315 ;
        RECT 133.700 170.120 134.930 170.600 ;
        RECT 102.035 169.930 102.325 169.975 ;
        RECT 100.270 169.790 102.325 169.930 ;
        RECT 72.670 169.450 73.730 169.590 ;
        RECT 72.670 169.310 72.810 169.450 ;
        RECT 99.735 169.405 100.025 169.635 ;
        RECT 22.455 169.250 22.745 169.295 ;
        RECT 23.820 169.250 24.140 169.310 ;
        RECT 22.455 169.110 24.140 169.250 ;
        RECT 22.455 169.065 22.745 169.110 ;
        RECT 23.820 169.050 24.140 169.110 ;
        RECT 30.275 169.250 30.565 169.295 ;
        RECT 30.720 169.250 31.040 169.310 ;
        RECT 30.275 169.110 31.040 169.250 ;
        RECT 30.275 169.065 30.565 169.110 ;
        RECT 30.720 169.050 31.040 169.110 ;
        RECT 33.940 169.250 34.260 169.310 ;
        RECT 41.315 169.250 41.605 169.295 ;
        RECT 33.940 169.110 41.605 169.250 ;
        RECT 33.940 169.050 34.260 169.110 ;
        RECT 41.315 169.065 41.605 169.110 ;
        RECT 44.535 169.250 44.825 169.295 ;
        RECT 44.980 169.250 45.300 169.310 ;
        RECT 44.535 169.110 45.300 169.250 ;
        RECT 44.535 169.065 44.825 169.110 ;
        RECT 44.980 169.050 45.300 169.110 ;
        RECT 66.615 169.250 66.905 169.295 ;
        RECT 72.580 169.250 72.900 169.310 ;
        RECT 66.615 169.110 72.900 169.250 ;
        RECT 66.615 169.065 66.905 169.110 ;
        RECT 72.580 169.050 72.900 169.110 ;
        RECT 94.660 169.250 94.980 169.310 ;
        RECT 95.135 169.250 95.425 169.295 ;
        RECT 94.660 169.110 95.425 169.250 ;
        RECT 94.660 169.050 94.980 169.110 ;
        RECT 95.135 169.065 95.425 169.110 ;
        RECT 96.960 169.250 97.280 169.310 ;
        RECT 100.270 169.250 100.410 169.790 ;
        RECT 102.035 169.745 102.325 169.790 ;
        RECT 102.940 169.730 103.260 169.990 ;
        RECT 107.170 169.930 107.310 170.085 ;
        RECT 105.330 169.790 107.310 169.930 ;
        RECT 105.330 169.635 105.470 169.790 ;
        RECT 105.255 169.405 105.545 169.635 ;
        RECT 96.960 169.110 100.410 169.250 ;
        RECT 96.960 169.050 97.280 169.110 ;
        RECT 15.010 168.430 113.450 168.910 ;
        RECT 33.480 168.230 33.800 168.290 ;
        RECT 34.860 168.230 35.180 168.290 ;
        RECT 38.080 168.230 38.400 168.290 ;
        RECT 33.480 168.090 38.400 168.230 ;
        RECT 33.480 168.030 33.800 168.090 ;
        RECT 34.860 168.030 35.180 168.090 ;
        RECT 38.080 168.030 38.400 168.090 ;
        RECT 57.400 168.230 57.720 168.290 ;
        RECT 60.160 168.230 60.480 168.290 ;
        RECT 57.400 168.090 60.480 168.230 ;
        RECT 57.400 168.030 57.720 168.090 ;
        RECT 60.160 168.030 60.480 168.090 ;
        RECT 65.695 168.230 65.985 168.275 ;
        RECT 66.140 168.230 66.460 168.290 ;
        RECT 65.695 168.090 66.460 168.230 ;
        RECT 65.695 168.045 65.985 168.090 ;
        RECT 66.140 168.030 66.460 168.090 ;
        RECT 83.620 168.230 83.940 168.290 ;
        RECT 84.555 168.230 84.845 168.275 ;
        RECT 107.080 168.230 107.400 168.290 ;
        RECT 108.475 168.230 108.765 168.275 ;
        RECT 83.620 168.090 84.845 168.230 ;
        RECT 83.620 168.030 83.940 168.090 ;
        RECT 84.555 168.045 84.845 168.090 ;
        RECT 85.090 168.090 108.765 168.230 ;
        RECT 20.255 167.890 20.545 167.935 ;
        RECT 23.375 167.890 23.665 167.935 ;
        RECT 25.265 167.890 25.555 167.935 ;
        RECT 20.255 167.750 25.555 167.890 ;
        RECT 20.255 167.705 20.545 167.750 ;
        RECT 23.375 167.705 23.665 167.750 ;
        RECT 25.265 167.705 25.555 167.750 ;
        RECT 29.455 167.890 29.745 167.935 ;
        RECT 32.575 167.890 32.865 167.935 ;
        RECT 34.465 167.890 34.755 167.935 ;
        RECT 29.455 167.750 34.755 167.890 ;
        RECT 29.455 167.705 29.745 167.750 ;
        RECT 32.575 167.705 32.865 167.750 ;
        RECT 34.465 167.705 34.755 167.750 ;
        RECT 56.020 167.890 56.340 167.950 ;
        RECT 56.955 167.890 57.245 167.935 ;
        RECT 65.220 167.890 65.540 167.950 ;
        RECT 67.520 167.890 67.840 167.950 ;
        RECT 56.020 167.750 57.245 167.890 ;
        RECT 56.020 167.690 56.340 167.750 ;
        RECT 56.955 167.705 57.245 167.750 ;
        RECT 64.850 167.750 67.840 167.890 ;
        RECT 16.920 167.550 17.240 167.610 ;
        RECT 17.395 167.550 17.685 167.595 ;
        RECT 31.180 167.550 31.500 167.610 ;
        RECT 16.920 167.410 31.500 167.550 ;
        RECT 16.920 167.350 17.240 167.410 ;
        RECT 17.395 167.365 17.685 167.410 ;
        RECT 31.180 167.350 31.500 167.410 ;
        RECT 33.940 167.350 34.260 167.610 ;
        RECT 37.160 167.550 37.480 167.610 ;
        RECT 37.160 167.410 44.290 167.550 ;
        RECT 37.160 167.350 37.480 167.410 ;
        RECT 17.840 166.870 18.160 166.930 ;
        RECT 19.175 166.915 19.465 167.230 ;
        RECT 20.255 167.210 20.545 167.255 ;
        RECT 23.835 167.210 24.125 167.255 ;
        RECT 25.670 167.210 25.960 167.255 ;
        RECT 20.255 167.070 25.960 167.210 ;
        RECT 20.255 167.025 20.545 167.070 ;
        RECT 23.835 167.025 24.125 167.070 ;
        RECT 25.670 167.025 25.960 167.070 ;
        RECT 26.135 167.210 26.425 167.255 ;
        RECT 26.580 167.210 26.900 167.270 ;
        RECT 26.135 167.070 26.900 167.210 ;
        RECT 26.135 167.025 26.425 167.070 ;
        RECT 26.580 167.010 26.900 167.070 ;
        RECT 18.875 166.870 19.465 166.915 ;
        RECT 22.115 166.870 22.765 166.915 ;
        RECT 17.840 166.730 22.765 166.870 ;
        RECT 17.840 166.670 18.160 166.730 ;
        RECT 18.875 166.685 19.165 166.730 ;
        RECT 22.115 166.685 22.765 166.730 ;
        RECT 24.755 166.870 25.045 166.915 ;
        RECT 25.200 166.870 25.520 166.930 ;
        RECT 28.375 166.915 28.665 167.230 ;
        RECT 29.455 167.210 29.745 167.255 ;
        RECT 33.035 167.210 33.325 167.255 ;
        RECT 34.870 167.210 35.160 167.255 ;
        RECT 29.455 167.070 35.160 167.210 ;
        RECT 29.455 167.025 29.745 167.070 ;
        RECT 33.035 167.025 33.325 167.070 ;
        RECT 34.870 167.025 35.160 167.070 ;
        RECT 35.320 167.210 35.640 167.270 ;
        RECT 36.715 167.210 37.005 167.255 ;
        RECT 35.320 167.070 37.005 167.210 ;
        RECT 35.320 167.010 35.640 167.070 ;
        RECT 36.715 167.025 37.005 167.070 ;
        RECT 39.920 167.010 40.240 167.270 ;
        RECT 44.150 167.255 44.290 167.410 ;
        RECT 53.260 167.350 53.580 167.610 ;
        RECT 60.160 167.550 60.480 167.610 ;
        RECT 63.380 167.550 63.700 167.610 ;
        RECT 64.850 167.595 64.990 167.750 ;
        RECT 65.220 167.690 65.540 167.750 ;
        RECT 67.520 167.690 67.840 167.750 ;
        RECT 72.550 167.890 72.840 167.935 ;
        RECT 75.330 167.890 75.620 167.935 ;
        RECT 77.190 167.890 77.480 167.935 ;
        RECT 72.550 167.750 77.480 167.890 ;
        RECT 72.550 167.705 72.840 167.750 ;
        RECT 75.330 167.705 75.620 167.750 ;
        RECT 77.190 167.705 77.480 167.750 ;
        RECT 64.315 167.550 64.605 167.595 ;
        RECT 56.110 167.410 57.170 167.550 ;
        RECT 44.075 167.210 44.365 167.255 ;
        RECT 54.655 167.210 54.945 167.255 ;
        RECT 44.075 167.070 54.945 167.210 ;
        RECT 44.075 167.025 44.365 167.070 ;
        RECT 54.655 167.025 54.945 167.070 ;
        RECT 55.560 167.210 55.880 167.270 ;
        RECT 56.110 167.255 56.250 167.410 ;
        RECT 56.035 167.210 56.325 167.255 ;
        RECT 55.560 167.070 56.325 167.210 ;
        RECT 31.640 166.915 31.960 166.930 ;
        RECT 24.755 166.730 25.520 166.870 ;
        RECT 24.755 166.685 25.045 166.730 ;
        RECT 25.200 166.670 25.520 166.730 ;
        RECT 28.075 166.870 28.665 166.915 ;
        RECT 31.315 166.870 31.965 166.915 ;
        RECT 28.075 166.730 31.965 166.870 ;
        RECT 28.075 166.685 28.365 166.730 ;
        RECT 31.315 166.685 31.965 166.730 ;
        RECT 41.760 166.870 42.080 166.930 ;
        RECT 43.615 166.870 43.905 166.915 ;
        RECT 41.760 166.730 43.905 166.870 ;
        RECT 31.640 166.670 31.960 166.685 ;
        RECT 41.760 166.670 42.080 166.730 ;
        RECT 43.615 166.685 43.905 166.730 ;
        RECT 44.520 166.670 44.840 166.930 ;
        RECT 26.595 166.530 26.885 166.575 ;
        RECT 27.040 166.530 27.360 166.590 ;
        RECT 26.595 166.390 27.360 166.530 ;
        RECT 26.595 166.345 26.885 166.390 ;
        RECT 27.040 166.330 27.360 166.390 ;
        RECT 42.680 166.330 43.000 166.590 ;
        RECT 54.730 166.530 54.870 167.025 ;
        RECT 55.560 167.010 55.880 167.070 ;
        RECT 56.035 167.025 56.325 167.070 ;
        RECT 56.480 167.010 56.800 167.270 ;
        RECT 57.030 167.210 57.170 167.410 ;
        RECT 60.160 167.410 64.605 167.550 ;
        RECT 60.160 167.350 60.480 167.410 ;
        RECT 63.380 167.350 63.700 167.410 ;
        RECT 64.315 167.365 64.605 167.410 ;
        RECT 64.775 167.365 65.065 167.595 ;
        RECT 77.655 167.550 77.945 167.595 ;
        RECT 82.240 167.550 82.560 167.610 ;
        RECT 83.710 167.550 83.850 168.030 ;
        RECT 65.310 167.410 76.490 167.550 ;
        RECT 60.635 167.210 60.925 167.255 ;
        RECT 61.540 167.210 61.860 167.270 ;
        RECT 65.310 167.210 65.450 167.410 ;
        RECT 57.030 167.070 65.450 167.210 ;
        RECT 66.155 167.210 66.445 167.255 ;
        RECT 66.600 167.210 66.920 167.270 ;
        RECT 66.155 167.070 66.920 167.210 ;
        RECT 60.635 167.025 60.925 167.070 ;
        RECT 61.540 167.010 61.860 167.070 ;
        RECT 66.155 167.025 66.445 167.070 ;
        RECT 66.600 167.010 66.920 167.070 ;
        RECT 68.685 167.210 68.975 167.255 ;
        RECT 71.660 167.210 71.980 167.270 ;
        RECT 68.685 167.070 71.980 167.210 ;
        RECT 68.685 167.025 68.975 167.070 ;
        RECT 71.660 167.010 71.980 167.070 ;
        RECT 72.550 167.210 72.840 167.255 ;
        RECT 72.550 167.070 75.085 167.210 ;
        RECT 72.550 167.025 72.840 167.070 ;
        RECT 74.870 166.915 75.085 167.070 ;
        RECT 75.800 167.010 76.120 167.270 ;
        RECT 76.350 167.210 76.490 167.410 ;
        RECT 77.655 167.410 83.850 167.550 ;
        RECT 77.655 167.365 77.945 167.410 ;
        RECT 82.240 167.350 82.560 167.410 ;
        RECT 85.090 167.210 85.230 168.090 ;
        RECT 107.080 168.030 107.400 168.090 ;
        RECT 108.475 168.045 108.765 168.090 ;
        RECT 95.235 167.890 95.525 167.935 ;
        RECT 98.355 167.890 98.645 167.935 ;
        RECT 100.245 167.890 100.535 167.935 ;
        RECT 95.235 167.750 100.535 167.890 ;
        RECT 95.235 167.705 95.525 167.750 ;
        RECT 98.355 167.705 98.645 167.750 ;
        RECT 100.245 167.705 100.535 167.750 ;
        RECT 91.900 167.550 92.220 167.610 ;
        RECT 92.375 167.550 92.665 167.595 ;
        RECT 91.900 167.410 92.665 167.550 ;
        RECT 91.900 167.350 92.220 167.410 ;
        RECT 92.375 167.365 92.665 167.410 ;
        RECT 99.260 167.550 99.580 167.610 ;
        RECT 101.575 167.550 101.865 167.595 ;
        RECT 102.020 167.550 102.340 167.610 ;
        RECT 99.260 167.410 102.340 167.550 ;
        RECT 99.260 167.350 99.580 167.410 ;
        RECT 101.575 167.365 101.865 167.410 ;
        RECT 102.020 167.350 102.340 167.410 ;
        RECT 76.350 167.070 85.230 167.210 ;
        RECT 88.680 167.010 89.000 167.270 ;
        RECT 89.155 167.025 89.445 167.255 ;
        RECT 70.690 166.870 70.980 166.915 ;
        RECT 73.950 166.870 74.240 166.915 ;
        RECT 74.870 166.870 75.160 166.915 ;
        RECT 76.730 166.870 77.020 166.915 ;
        RECT 70.690 166.730 74.650 166.870 ;
        RECT 70.690 166.685 70.980 166.730 ;
        RECT 73.950 166.685 74.240 166.730 ;
        RECT 56.480 166.530 56.800 166.590 ;
        RECT 54.730 166.390 56.800 166.530 ;
        RECT 56.480 166.330 56.800 166.390 ;
        RECT 64.315 166.530 64.605 166.575 ;
        RECT 64.760 166.530 65.080 166.590 ;
        RECT 64.315 166.390 65.080 166.530 ;
        RECT 74.510 166.530 74.650 166.730 ;
        RECT 74.870 166.730 77.020 166.870 ;
        RECT 74.870 166.685 75.160 166.730 ;
        RECT 76.730 166.685 77.020 166.730 ;
        RECT 78.115 166.870 78.405 166.915 ;
        RECT 81.780 166.870 82.100 166.930 ;
        RECT 89.230 166.870 89.370 167.025 ;
        RECT 90.980 167.010 91.300 167.270 ;
        RECT 78.115 166.730 82.100 166.870 ;
        RECT 78.115 166.685 78.405 166.730 ;
        RECT 81.780 166.670 82.100 166.730 ;
        RECT 84.170 166.730 89.370 166.870 ;
        RECT 89.615 166.870 89.905 166.915 ;
        RECT 91.440 166.870 91.760 166.930 ;
        RECT 94.155 166.915 94.445 167.230 ;
        RECT 95.235 167.210 95.525 167.255 ;
        RECT 98.815 167.210 99.105 167.255 ;
        RECT 100.650 167.210 100.940 167.255 ;
        RECT 95.235 167.070 100.940 167.210 ;
        RECT 95.235 167.025 95.525 167.070 ;
        RECT 98.815 167.025 99.105 167.070 ;
        RECT 100.650 167.025 100.940 167.070 ;
        RECT 101.100 167.010 101.420 167.270 ;
        RECT 104.780 167.210 105.100 167.270 ;
        RECT 106.635 167.210 106.925 167.255 ;
        RECT 104.780 167.070 106.925 167.210 ;
        RECT 104.780 167.010 105.100 167.070 ;
        RECT 106.635 167.025 106.925 167.070 ;
        RECT 108.935 167.210 109.225 167.255 ;
        RECT 113.520 167.210 113.840 167.270 ;
        RECT 108.935 167.070 113.840 167.210 ;
        RECT 108.935 167.025 109.225 167.070 ;
        RECT 113.520 167.010 113.840 167.070 ;
        RECT 89.615 166.730 91.760 166.870 ;
        RECT 77.180 166.530 77.500 166.590 ;
        RECT 74.510 166.390 77.500 166.530 ;
        RECT 64.315 166.345 64.605 166.390 ;
        RECT 64.760 166.330 65.080 166.390 ;
        RECT 77.180 166.330 77.500 166.390 ;
        RECT 79.480 166.530 79.800 166.590 ;
        RECT 84.170 166.530 84.310 166.730 ;
        RECT 89.615 166.685 89.905 166.730 ;
        RECT 91.440 166.670 91.760 166.730 ;
        RECT 93.855 166.870 94.445 166.915 ;
        RECT 94.660 166.870 94.980 166.930 ;
        RECT 97.095 166.870 97.745 166.915 ;
        RECT 93.855 166.730 97.745 166.870 ;
        RECT 93.855 166.685 94.145 166.730 ;
        RECT 94.660 166.670 94.980 166.730 ;
        RECT 97.095 166.685 97.745 166.730 ;
        RECT 99.720 166.670 100.040 166.930 ;
        RECT 79.480 166.390 84.310 166.530 ;
        RECT 86.840 166.530 87.160 166.590 ;
        RECT 87.775 166.530 88.065 166.575 ;
        RECT 86.840 166.390 88.065 166.530 ;
        RECT 79.480 166.330 79.800 166.390 ;
        RECT 86.840 166.330 87.160 166.390 ;
        RECT 87.775 166.345 88.065 166.390 ;
        RECT 91.915 166.530 92.205 166.575 ;
        RECT 96.500 166.530 96.820 166.590 ;
        RECT 91.915 166.390 96.820 166.530 ;
        RECT 91.915 166.345 92.205 166.390 ;
        RECT 96.500 166.330 96.820 166.390 ;
        RECT 102.940 166.530 103.260 166.590 ;
        RECT 104.795 166.530 105.085 166.575 ;
        RECT 102.940 166.390 105.085 166.530 ;
        RECT 102.940 166.330 103.260 166.390 ;
        RECT 104.795 166.345 105.085 166.390 ;
        RECT 107.555 166.530 107.845 166.575 ;
        RECT 109.380 166.530 109.700 166.590 ;
        RECT 107.555 166.390 109.700 166.530 ;
        RECT 107.555 166.345 107.845 166.390 ;
        RECT 109.380 166.330 109.700 166.390 ;
        RECT 15.010 165.710 113.450 166.190 ;
        RECT 17.840 165.310 18.160 165.570 ;
        RECT 21.060 165.510 21.380 165.570 ;
        RECT 22.455 165.510 22.745 165.555 ;
        RECT 21.060 165.370 22.745 165.510 ;
        RECT 21.060 165.310 21.380 165.370 ;
        RECT 22.455 165.325 22.745 165.370 ;
        RECT 24.740 165.310 25.060 165.570 ;
        RECT 25.200 165.310 25.520 165.570 ;
        RECT 43.140 165.510 43.460 165.570 ;
        RECT 43.140 165.370 47.510 165.510 ;
        RECT 43.140 165.310 43.460 165.370 ;
        RECT 47.370 165.230 47.510 165.370 ;
        RECT 71.660 165.310 71.980 165.570 ;
        RECT 73.975 165.325 74.265 165.555 ;
        RECT 19.680 164.970 20.000 165.230 ;
        RECT 26.580 165.170 26.900 165.230 ;
        RECT 29.340 165.170 29.660 165.230 ;
        RECT 30.275 165.170 30.565 165.215 ;
        RECT 35.320 165.170 35.640 165.230 ;
        RECT 38.080 165.170 38.400 165.230 ;
        RECT 26.580 165.030 38.400 165.170 ;
        RECT 26.580 164.970 26.900 165.030 ;
        RECT 29.340 164.970 29.660 165.030 ;
        RECT 30.275 164.985 30.565 165.030 ;
        RECT 35.320 164.970 35.640 165.030 ;
        RECT 38.080 164.970 38.400 165.030 ;
        RECT 39.000 164.970 39.320 165.230 ;
        RECT 40.955 165.170 41.245 165.215 ;
        RECT 41.760 165.170 42.080 165.230 ;
        RECT 44.195 165.170 44.845 165.215 ;
        RECT 40.955 165.030 44.845 165.170 ;
        RECT 40.955 164.985 41.545 165.030 ;
        RECT 18.315 164.830 18.605 164.875 ;
        RECT 19.770 164.830 19.910 164.970 ;
        RECT 18.315 164.690 19.910 164.830 ;
        RECT 20.615 164.830 20.905 164.875 ;
        RECT 21.060 164.830 21.380 164.890 ;
        RECT 20.615 164.690 21.380 164.830 ;
        RECT 18.315 164.645 18.605 164.690 ;
        RECT 20.615 164.645 20.905 164.690 ;
        RECT 21.060 164.630 21.380 164.690 ;
        RECT 23.820 164.630 24.140 164.890 ;
        RECT 26.120 164.630 26.440 164.890 ;
        RECT 41.255 164.670 41.545 164.985 ;
        RECT 41.760 164.970 42.080 165.030 ;
        RECT 44.195 164.985 44.845 165.030 ;
        RECT 46.820 164.970 47.140 165.230 ;
        RECT 47.280 165.170 47.600 165.230 ;
        RECT 51.535 165.170 51.825 165.215 ;
        RECT 54.775 165.170 55.425 165.215 ;
        RECT 56.020 165.170 56.340 165.230 ;
        RECT 47.280 165.030 50.730 165.170 ;
        RECT 47.280 164.970 47.600 165.030 ;
        RECT 42.335 164.830 42.625 164.875 ;
        RECT 45.915 164.830 46.205 164.875 ;
        RECT 47.750 164.830 48.040 164.875 ;
        RECT 42.335 164.690 48.040 164.830 ;
        RECT 42.335 164.645 42.625 164.690 ;
        RECT 45.915 164.645 46.205 164.690 ;
        RECT 47.750 164.645 48.040 164.690 ;
        RECT 19.695 164.305 19.985 164.535 ;
        RECT 19.770 163.810 19.910 164.305 ;
        RECT 20.140 164.290 20.460 164.550 ;
        RECT 27.040 164.290 27.360 164.550 ;
        RECT 38.080 164.490 38.400 164.550 ;
        RECT 48.215 164.490 48.505 164.535 ;
        RECT 38.080 164.350 48.505 164.490 ;
        RECT 38.080 164.290 38.400 164.350 ;
        RECT 48.215 164.305 48.505 164.350 ;
        RECT 20.230 164.150 20.370 164.290 ;
        RECT 37.620 164.150 37.940 164.210 ;
        RECT 20.230 164.010 37.940 164.150 ;
        RECT 37.620 163.950 37.940 164.010 ;
        RECT 42.335 164.150 42.625 164.195 ;
        RECT 45.455 164.150 45.745 164.195 ;
        RECT 47.345 164.150 47.635 164.195 ;
        RECT 42.335 164.010 47.635 164.150 ;
        RECT 42.335 163.965 42.625 164.010 ;
        RECT 45.455 163.965 45.745 164.010 ;
        RECT 47.345 163.965 47.635 164.010 ;
        RECT 50.590 163.870 50.730 165.030 ;
        RECT 51.535 165.030 56.340 165.170 ;
        RECT 51.535 164.985 52.125 165.030 ;
        RECT 54.775 164.985 55.425 165.030 ;
        RECT 51.835 164.670 52.125 164.985 ;
        RECT 56.020 164.970 56.340 165.030 ;
        RECT 57.860 165.170 58.180 165.230 ;
        RECT 63.855 165.170 64.145 165.215 ;
        RECT 64.760 165.170 65.080 165.230 ;
        RECT 57.860 165.030 59.010 165.170 ;
        RECT 57.860 164.970 58.180 165.030 ;
        RECT 58.870 164.875 59.010 165.030 ;
        RECT 63.855 165.030 65.080 165.170 ;
        RECT 63.855 164.985 64.145 165.030 ;
        RECT 64.760 164.970 65.080 165.030 ;
        RECT 71.200 165.170 71.520 165.230 ;
        RECT 72.135 165.170 72.425 165.215 ;
        RECT 71.200 165.030 72.425 165.170 ;
        RECT 71.200 164.970 71.520 165.030 ;
        RECT 72.135 164.985 72.425 165.030 ;
        RECT 52.915 164.830 53.205 164.875 ;
        RECT 56.495 164.830 56.785 164.875 ;
        RECT 58.330 164.830 58.620 164.875 ;
        RECT 52.915 164.690 58.620 164.830 ;
        RECT 52.915 164.645 53.205 164.690 ;
        RECT 56.495 164.645 56.785 164.690 ;
        RECT 58.330 164.645 58.620 164.690 ;
        RECT 58.795 164.830 59.085 164.875 ;
        RECT 61.080 164.830 61.400 164.890 ;
        RECT 58.795 164.690 61.400 164.830 ;
        RECT 58.795 164.645 59.085 164.690 ;
        RECT 61.080 164.630 61.400 164.690 ;
        RECT 61.540 164.630 61.860 164.890 ;
        RECT 74.050 164.830 74.190 165.325 ;
        RECT 75.800 165.310 76.120 165.570 ;
        RECT 77.180 165.510 77.500 165.570 ;
        RECT 78.575 165.510 78.865 165.555 ;
        RECT 77.180 165.370 78.865 165.510 ;
        RECT 77.180 165.310 77.500 165.370 ;
        RECT 78.575 165.325 78.865 165.370 ;
        RECT 99.720 165.310 100.040 165.570 ;
        RECT 135.580 165.470 136.830 166.590 ;
        RECT 80.860 165.170 81.180 165.230 ;
        RECT 91.440 165.215 91.760 165.230 ;
        RECT 81.730 165.170 82.020 165.215 ;
        RECT 84.990 165.170 85.280 165.215 ;
        RECT 80.860 165.030 85.280 165.170 ;
        RECT 80.860 164.970 81.180 165.030 ;
        RECT 81.730 164.985 82.020 165.030 ;
        RECT 84.990 164.985 85.280 165.030 ;
        RECT 85.910 165.170 86.200 165.215 ;
        RECT 87.770 165.170 88.060 165.215 ;
        RECT 85.910 165.030 88.060 165.170 ;
        RECT 85.910 164.985 86.200 165.030 ;
        RECT 87.770 164.985 88.060 165.030 ;
        RECT 91.390 165.170 91.760 165.215 ;
        RECT 94.650 165.170 94.940 165.215 ;
        RECT 91.390 165.030 94.940 165.170 ;
        RECT 91.390 164.985 91.760 165.030 ;
        RECT 94.650 164.985 94.940 165.030 ;
        RECT 95.570 165.170 95.860 165.215 ;
        RECT 97.430 165.170 97.720 165.215 ;
        RECT 101.115 165.170 101.405 165.215 ;
        RECT 103.515 165.170 103.805 165.215 ;
        RECT 106.755 165.170 107.405 165.215 ;
        RECT 95.570 165.030 97.720 165.170 ;
        RECT 95.570 164.985 95.860 165.030 ;
        RECT 97.430 164.985 97.720 165.030 ;
        RECT 98.430 165.030 100.410 165.170 ;
        RECT 74.895 164.830 75.185 164.875 ;
        RECT 74.050 164.690 75.185 164.830 ;
        RECT 74.895 164.645 75.185 164.690 ;
        RECT 77.655 164.830 77.945 164.875 ;
        RECT 79.035 164.830 79.325 164.875 ;
        RECT 79.480 164.830 79.800 164.890 ;
        RECT 77.655 164.690 79.800 164.830 ;
        RECT 77.655 164.645 77.945 164.690 ;
        RECT 79.035 164.645 79.325 164.690 ;
        RECT 79.480 164.630 79.800 164.690 ;
        RECT 83.590 164.830 83.880 164.875 ;
        RECT 85.910 164.830 86.125 164.985 ;
        RECT 91.440 164.970 91.760 164.985 ;
        RECT 83.590 164.690 86.125 164.830 ;
        RECT 83.590 164.645 83.880 164.690 ;
        RECT 86.840 164.630 87.160 164.890 ;
        RECT 88.220 164.830 88.540 164.890 ;
        RECT 88.695 164.830 88.985 164.875 ;
        RECT 88.220 164.690 88.985 164.830 ;
        RECT 88.220 164.630 88.540 164.690 ;
        RECT 88.695 164.645 88.985 164.690 ;
        RECT 93.250 164.830 93.540 164.875 ;
        RECT 95.570 164.830 95.785 164.985 ;
        RECT 93.250 164.690 95.785 164.830 ;
        RECT 93.250 164.645 93.540 164.690 ;
        RECT 57.400 164.290 57.720 164.550 ;
        RECT 60.175 164.305 60.465 164.535 ;
        RECT 71.215 164.490 71.505 164.535 ;
        RECT 72.580 164.490 72.900 164.550 ;
        RECT 71.215 164.350 72.900 164.490 ;
        RECT 88.770 164.490 88.910 164.645 ;
        RECT 96.500 164.630 96.820 164.890 ;
        RECT 98.430 164.535 98.570 165.030 ;
        RECT 98.815 164.645 99.105 164.875 ;
        RECT 98.355 164.490 98.645 164.535 ;
        RECT 88.770 164.350 98.645 164.490 ;
        RECT 71.215 164.305 71.505 164.350 ;
        RECT 52.915 164.150 53.205 164.195 ;
        RECT 56.035 164.150 56.325 164.195 ;
        RECT 57.925 164.150 58.215 164.195 ;
        RECT 52.915 164.010 58.215 164.150 ;
        RECT 52.915 163.965 53.205 164.010 ;
        RECT 56.035 163.965 56.325 164.010 ;
        RECT 57.925 163.965 58.215 164.010 ;
        RECT 58.780 164.150 59.100 164.210 ;
        RECT 60.250 164.150 60.390 164.305 ;
        RECT 72.580 164.290 72.900 164.350 ;
        RECT 98.355 164.305 98.645 164.350 ;
        RECT 58.780 164.010 60.390 164.150 ;
        RECT 69.820 164.150 70.140 164.210 ;
        RECT 79.725 164.150 80.015 164.195 ;
        RECT 82.700 164.150 83.020 164.210 ;
        RECT 69.820 164.010 83.020 164.150 ;
        RECT 58.780 163.950 59.100 164.010 ;
        RECT 69.820 163.950 70.140 164.010 ;
        RECT 79.725 163.965 80.015 164.010 ;
        RECT 82.700 163.950 83.020 164.010 ;
        RECT 83.590 164.150 83.880 164.195 ;
        RECT 86.370 164.150 86.660 164.195 ;
        RECT 88.230 164.150 88.520 164.195 ;
        RECT 83.590 164.010 88.520 164.150 ;
        RECT 83.590 163.965 83.880 164.010 ;
        RECT 86.370 163.965 86.660 164.010 ;
        RECT 88.230 163.965 88.520 164.010 ;
        RECT 93.250 164.150 93.540 164.195 ;
        RECT 96.030 164.150 96.320 164.195 ;
        RECT 97.890 164.150 98.180 164.195 ;
        RECT 93.250 164.010 98.180 164.150 ;
        RECT 98.890 164.150 99.030 164.645 ;
        RECT 100.270 164.490 100.410 165.030 ;
        RECT 101.115 165.030 107.405 165.170 ;
        RECT 101.115 164.985 101.405 165.030 ;
        RECT 103.515 164.985 104.105 165.030 ;
        RECT 106.755 164.985 107.405 165.030 ;
        RECT 100.640 164.630 100.960 164.890 ;
        RECT 103.815 164.670 104.105 164.985 ;
        RECT 109.380 164.970 109.700 165.230 ;
        RECT 104.895 164.830 105.185 164.875 ;
        RECT 108.475 164.830 108.765 164.875 ;
        RECT 110.310 164.830 110.600 164.875 ;
        RECT 104.895 164.690 110.600 164.830 ;
        RECT 104.895 164.645 105.185 164.690 ;
        RECT 108.475 164.645 108.765 164.690 ;
        RECT 110.310 164.645 110.600 164.690 ;
        RECT 101.100 164.490 101.420 164.550 ;
        RECT 104.320 164.490 104.640 164.550 ;
        RECT 110.760 164.490 111.080 164.550 ;
        RECT 100.270 164.350 111.080 164.490 ;
        RECT 101.100 164.290 101.420 164.350 ;
        RECT 104.320 164.290 104.640 164.350 ;
        RECT 110.760 164.290 111.080 164.350 ;
        RECT 103.860 164.150 104.180 164.210 ;
        RECT 98.890 164.010 104.180 164.150 ;
        RECT 93.250 163.965 93.540 164.010 ;
        RECT 96.030 163.965 96.320 164.010 ;
        RECT 97.890 163.965 98.180 164.010 ;
        RECT 103.860 163.950 104.180 164.010 ;
        RECT 104.895 164.150 105.185 164.195 ;
        RECT 108.015 164.150 108.305 164.195 ;
        RECT 109.905 164.150 110.195 164.195 ;
        RECT 104.895 164.010 110.195 164.150 ;
        RECT 104.895 163.965 105.185 164.010 ;
        RECT 108.015 163.965 108.305 164.010 ;
        RECT 109.905 163.965 110.195 164.010 ;
        RECT 22.900 163.810 23.220 163.870 ;
        RECT 25.660 163.810 25.980 163.870 ;
        RECT 19.770 163.670 25.980 163.810 ;
        RECT 22.900 163.610 23.220 163.670 ;
        RECT 25.660 163.610 25.980 163.670 ;
        RECT 29.815 163.810 30.105 163.855 ;
        RECT 33.480 163.810 33.800 163.870 ;
        RECT 29.815 163.670 33.800 163.810 ;
        RECT 29.815 163.625 30.105 163.670 ;
        RECT 33.480 163.610 33.800 163.670 ;
        RECT 39.475 163.810 39.765 163.855 ;
        RECT 39.920 163.810 40.240 163.870 ;
        RECT 39.475 163.670 40.240 163.810 ;
        RECT 39.475 163.625 39.765 163.670 ;
        RECT 39.920 163.610 40.240 163.670 ;
        RECT 45.900 163.810 46.220 163.870 ;
        RECT 50.055 163.810 50.345 163.855 ;
        RECT 45.900 163.670 50.345 163.810 ;
        RECT 45.900 163.610 46.220 163.670 ;
        RECT 50.055 163.625 50.345 163.670 ;
        RECT 50.500 163.810 50.820 163.870 ;
        RECT 62.475 163.810 62.765 163.855 ;
        RECT 50.500 163.670 62.765 163.810 ;
        RECT 50.500 163.610 50.820 163.670 ;
        RECT 62.475 163.625 62.765 163.670 ;
        RECT 76.720 163.810 77.040 163.870 ;
        RECT 77.195 163.810 77.485 163.855 ;
        RECT 76.720 163.670 77.485 163.810 ;
        RECT 76.720 163.610 77.040 163.670 ;
        RECT 77.195 163.625 77.485 163.670 ;
        RECT 84.540 163.810 84.860 163.870 ;
        RECT 89.385 163.810 89.675 163.855 ;
        RECT 90.520 163.810 90.840 163.870 ;
        RECT 84.540 163.670 90.840 163.810 ;
        RECT 84.540 163.610 84.860 163.670 ;
        RECT 89.385 163.625 89.675 163.670 ;
        RECT 90.520 163.610 90.840 163.670 ;
        RECT 102.020 163.610 102.340 163.870 ;
        RECT 15.010 162.990 113.450 163.470 ;
        RECT 26.120 162.590 26.440 162.850 ;
        RECT 27.040 162.790 27.360 162.850 ;
        RECT 41.760 162.790 42.080 162.850 ;
        RECT 27.040 162.650 42.080 162.790 ;
        RECT 27.040 162.590 27.360 162.650 ;
        RECT 41.760 162.590 42.080 162.650 ;
        RECT 42.220 162.790 42.540 162.850 ;
        RECT 43.155 162.790 43.445 162.835 ;
        RECT 42.220 162.650 43.445 162.790 ;
        RECT 42.220 162.590 42.540 162.650 ;
        RECT 43.155 162.605 43.445 162.650 ;
        RECT 45.455 162.790 45.745 162.835 ;
        RECT 46.820 162.790 47.140 162.850 ;
        RECT 45.455 162.650 47.140 162.790 ;
        RECT 45.455 162.605 45.745 162.650 ;
        RECT 46.820 162.590 47.140 162.650 ;
        RECT 49.135 162.790 49.425 162.835 ;
        RECT 49.580 162.790 49.900 162.850 ;
        RECT 49.135 162.650 49.900 162.790 ;
        RECT 49.135 162.605 49.425 162.650 ;
        RECT 49.580 162.590 49.900 162.650 ;
        RECT 55.575 162.790 55.865 162.835 ;
        RECT 57.400 162.790 57.720 162.850 ;
        RECT 55.575 162.650 57.720 162.790 ;
        RECT 55.575 162.605 55.865 162.650 ;
        RECT 57.400 162.590 57.720 162.650 ;
        RECT 58.320 162.790 58.640 162.850 ;
        RECT 67.520 162.790 67.840 162.850 ;
        RECT 58.320 162.650 67.840 162.790 ;
        RECT 58.320 162.590 58.640 162.650 ;
        RECT 67.520 162.590 67.840 162.650 ;
        RECT 86.855 162.790 87.145 162.835 ;
        RECT 88.680 162.790 89.000 162.850 ;
        RECT 86.855 162.650 89.000 162.790 ;
        RECT 86.855 162.605 87.145 162.650 ;
        RECT 88.680 162.590 89.000 162.650 ;
        RECT 90.980 162.790 91.300 162.850 ;
        RECT 91.915 162.790 92.205 162.835 ;
        RECT 90.980 162.650 92.205 162.790 ;
        RECT 90.980 162.590 91.300 162.650 ;
        RECT 91.915 162.605 92.205 162.650 ;
        RECT 99.735 162.790 100.025 162.835 ;
        RECT 99.735 162.650 102.710 162.790 ;
        RECT 99.735 162.605 100.025 162.650 ;
        RECT 20.570 162.450 20.860 162.495 ;
        RECT 23.350 162.450 23.640 162.495 ;
        RECT 25.210 162.450 25.500 162.495 ;
        RECT 20.570 162.310 25.500 162.450 ;
        RECT 20.570 162.265 20.860 162.310 ;
        RECT 23.350 162.265 23.640 162.310 ;
        RECT 25.210 162.265 25.500 162.310 ;
        RECT 25.660 162.450 25.980 162.510 ;
        RECT 37.620 162.450 37.940 162.510 ;
        RECT 49.670 162.450 49.810 162.590 ;
        RECT 65.680 162.450 66.000 162.510 ;
        RECT 69.360 162.450 69.680 162.510 ;
        RECT 25.660 162.310 29.570 162.450 ;
        RECT 25.660 162.250 25.980 162.310 ;
        RECT 21.060 162.110 21.380 162.170 ;
        RECT 29.430 162.155 29.570 162.310 ;
        RECT 32.650 162.310 36.010 162.450 ;
        RECT 32.650 162.155 32.790 162.310 ;
        RECT 28.435 162.110 28.725 162.155 ;
        RECT 21.060 161.970 28.725 162.110 ;
        RECT 21.060 161.910 21.380 161.970 ;
        RECT 28.435 161.925 28.725 161.970 ;
        RECT 29.355 162.110 29.645 162.155 ;
        RECT 32.575 162.110 32.865 162.155 ;
        RECT 35.320 162.110 35.640 162.170 ;
        RECT 29.355 161.970 32.865 162.110 ;
        RECT 29.355 161.925 29.645 161.970 ;
        RECT 32.575 161.925 32.865 161.970 ;
        RECT 33.110 161.970 35.640 162.110 ;
        RECT 35.870 162.110 36.010 162.310 ;
        RECT 37.620 162.310 45.670 162.450 ;
        RECT 49.670 162.310 51.190 162.450 ;
        RECT 37.620 162.250 37.940 162.310 ;
        RECT 40.395 162.110 40.685 162.155 ;
        RECT 43.140 162.110 43.460 162.170 ;
        RECT 35.870 161.970 43.460 162.110 ;
        RECT 20.570 161.770 20.860 161.815 ;
        RECT 23.835 161.770 24.125 161.815 ;
        RECT 24.280 161.770 24.600 161.830 ;
        RECT 20.570 161.630 23.105 161.770 ;
        RECT 20.570 161.585 20.860 161.630 ;
        RECT 17.840 161.430 18.160 161.490 ;
        RECT 22.890 161.475 23.105 161.630 ;
        RECT 23.835 161.630 24.600 161.770 ;
        RECT 23.835 161.585 24.125 161.630 ;
        RECT 24.280 161.570 24.600 161.630 ;
        RECT 25.675 161.770 25.965 161.815 ;
        RECT 26.580 161.770 26.900 161.830 ;
        RECT 25.675 161.630 26.900 161.770 ;
        RECT 25.675 161.585 25.965 161.630 ;
        RECT 26.580 161.570 26.900 161.630 ;
        RECT 30.275 161.770 30.565 161.815 ;
        RECT 33.110 161.770 33.250 161.970 ;
        RECT 35.320 161.910 35.640 161.970 ;
        RECT 40.395 161.925 40.685 161.970 ;
        RECT 43.140 161.910 43.460 161.970 ;
        RECT 30.275 161.630 33.250 161.770 ;
        RECT 33.480 161.770 33.800 161.830 ;
        RECT 40.855 161.770 41.145 161.815 ;
        RECT 33.480 161.630 41.145 161.770 ;
        RECT 30.275 161.585 30.565 161.630 ;
        RECT 33.480 161.570 33.800 161.630 ;
        RECT 40.855 161.585 41.145 161.630 ;
        RECT 41.315 161.770 41.605 161.815 ;
        RECT 42.680 161.770 43.000 161.830 ;
        RECT 41.315 161.630 43.000 161.770 ;
        RECT 41.315 161.585 41.605 161.630 ;
        RECT 42.680 161.570 43.000 161.630 ;
        RECT 44.535 161.770 44.825 161.815 ;
        RECT 44.980 161.770 45.300 161.830 ;
        RECT 44.535 161.630 45.300 161.770 ;
        RECT 45.530 161.770 45.670 162.310 ;
        RECT 45.900 161.910 46.220 162.170 ;
        RECT 50.500 161.910 50.820 162.170 ;
        RECT 51.050 162.155 51.190 162.310 ;
        RECT 65.680 162.310 69.680 162.450 ;
        RECT 65.680 162.250 66.000 162.310 ;
        RECT 69.360 162.250 69.680 162.310 ;
        RECT 77.150 162.450 77.440 162.495 ;
        RECT 79.930 162.450 80.220 162.495 ;
        RECT 81.790 162.450 82.080 162.495 ;
        RECT 77.150 162.310 82.080 162.450 ;
        RECT 77.150 162.265 77.440 162.310 ;
        RECT 79.930 162.265 80.220 162.310 ;
        RECT 81.790 162.265 82.080 162.310 ;
        RECT 82.700 162.450 83.020 162.510 ;
        RECT 82.700 162.310 84.770 162.450 ;
        RECT 82.700 162.250 83.020 162.310 ;
        RECT 50.975 161.925 51.265 162.155 ;
        RECT 66.600 162.110 66.920 162.170 ;
        RECT 59.790 161.970 66.920 162.110 ;
        RECT 51.435 161.770 51.725 161.815 ;
        RECT 45.530 161.630 51.725 161.770 ;
        RECT 44.535 161.585 44.825 161.630 ;
        RECT 44.980 161.570 45.300 161.630 ;
        RECT 51.435 161.585 51.725 161.630 ;
        RECT 54.640 161.570 54.960 161.830 ;
        RECT 59.790 161.815 59.930 161.970 ;
        RECT 66.600 161.910 66.920 161.970 ;
        RECT 69.835 162.110 70.125 162.155 ;
        RECT 72.580 162.110 72.900 162.170 ;
        RECT 69.835 161.970 82.010 162.110 ;
        RECT 69.835 161.925 70.125 161.970 ;
        RECT 72.580 161.910 72.900 161.970 ;
        RECT 59.255 161.770 59.545 161.815 ;
        RECT 59.715 161.770 60.005 161.815 ;
        RECT 59.255 161.630 60.005 161.770 ;
        RECT 59.255 161.585 59.545 161.630 ;
        RECT 59.715 161.585 60.005 161.630 ;
        RECT 60.160 161.770 60.480 161.830 ;
        RECT 63.395 161.770 63.685 161.815 ;
        RECT 60.160 161.630 63.685 161.770 ;
        RECT 60.160 161.570 60.480 161.630 ;
        RECT 63.395 161.585 63.685 161.630 ;
        RECT 65.235 161.770 65.525 161.815 ;
        RECT 66.140 161.770 66.460 161.830 ;
        RECT 67.075 161.770 67.365 161.815 ;
        RECT 65.235 161.630 67.365 161.770 ;
        RECT 65.235 161.585 65.525 161.630 ;
        RECT 66.140 161.570 66.460 161.630 ;
        RECT 67.075 161.585 67.365 161.630 ;
        RECT 77.150 161.770 77.440 161.815 ;
        RECT 77.150 161.630 79.685 161.770 ;
        RECT 77.150 161.585 77.440 161.630 ;
        RECT 18.710 161.430 19.000 161.475 ;
        RECT 21.970 161.430 22.260 161.475 ;
        RECT 17.840 161.290 22.260 161.430 ;
        RECT 17.840 161.230 18.160 161.290 ;
        RECT 18.710 161.245 19.000 161.290 ;
        RECT 21.970 161.245 22.260 161.290 ;
        RECT 22.890 161.430 23.180 161.475 ;
        RECT 24.750 161.430 25.040 161.475 ;
        RECT 22.890 161.290 25.040 161.430 ;
        RECT 22.890 161.245 23.180 161.290 ;
        RECT 24.750 161.245 25.040 161.290 ;
        RECT 39.460 161.430 39.780 161.490 ;
        RECT 65.680 161.430 66.000 161.490 ;
        RECT 66.600 161.430 66.920 161.490 ;
        RECT 69.820 161.430 70.140 161.490 ;
        RECT 70.755 161.430 71.045 161.475 ;
        RECT 73.285 161.430 73.575 161.475 ;
        RECT 39.460 161.290 66.370 161.430 ;
        RECT 39.460 161.230 39.780 161.290 ;
        RECT 65.680 161.230 66.000 161.290 ;
        RECT 16.705 161.090 16.995 161.135 ;
        RECT 22.440 161.090 22.760 161.150 ;
        RECT 16.705 160.950 22.760 161.090 ;
        RECT 16.705 160.905 16.995 160.950 ;
        RECT 22.440 160.890 22.760 160.950 ;
        RECT 27.960 160.890 28.280 161.150 ;
        RECT 30.735 161.090 31.025 161.135 ;
        RECT 31.180 161.090 31.500 161.150 ;
        RECT 30.735 160.950 31.500 161.090 ;
        RECT 30.735 160.905 31.025 160.950 ;
        RECT 31.180 160.890 31.500 160.950 ;
        RECT 32.100 161.090 32.420 161.150 ;
        RECT 33.035 161.090 33.325 161.135 ;
        RECT 32.100 160.950 33.325 161.090 ;
        RECT 32.100 160.890 32.420 160.950 ;
        RECT 33.035 160.905 33.325 160.950 ;
        RECT 35.335 161.090 35.625 161.135 ;
        RECT 35.780 161.090 36.100 161.150 ;
        RECT 35.335 160.950 36.100 161.090 ;
        RECT 35.335 160.905 35.625 160.950 ;
        RECT 35.780 160.890 36.100 160.950 ;
        RECT 50.960 161.090 51.280 161.150 ;
        RECT 53.275 161.090 53.565 161.135 ;
        RECT 50.960 160.950 53.565 161.090 ;
        RECT 50.960 160.890 51.280 160.950 ;
        RECT 53.275 160.905 53.565 160.950 ;
        RECT 59.700 161.090 60.020 161.150 ;
        RECT 60.635 161.090 60.925 161.135 ;
        RECT 62.000 161.090 62.320 161.150 ;
        RECT 59.700 160.950 62.320 161.090 ;
        RECT 59.700 160.890 60.020 160.950 ;
        RECT 60.635 160.905 60.925 160.950 ;
        RECT 62.000 160.890 62.320 160.950 ;
        RECT 64.315 161.090 64.605 161.135 ;
        RECT 65.220 161.090 65.540 161.150 ;
        RECT 66.230 161.135 66.370 161.290 ;
        RECT 66.600 161.290 71.045 161.430 ;
        RECT 66.600 161.230 66.920 161.290 ;
        RECT 69.820 161.230 70.140 161.290 ;
        RECT 70.755 161.245 71.045 161.290 ;
        RECT 71.290 161.290 73.575 161.430 ;
        RECT 71.290 161.150 71.430 161.290 ;
        RECT 73.285 161.245 73.575 161.290 ;
        RECT 75.290 161.430 75.580 161.475 ;
        RECT 76.720 161.430 77.040 161.490 ;
        RECT 79.470 161.475 79.685 161.630 ;
        RECT 80.400 161.570 80.720 161.830 ;
        RECT 81.870 161.770 82.010 161.970 ;
        RECT 82.240 161.910 82.560 162.170 ;
        RECT 83.635 162.110 83.925 162.155 ;
        RECT 84.080 162.110 84.400 162.170 ;
        RECT 84.630 162.155 84.770 162.310 ;
        RECT 86.010 162.310 94.890 162.450 ;
        RECT 83.635 161.970 84.400 162.110 ;
        RECT 83.635 161.925 83.925 161.970 ;
        RECT 83.710 161.770 83.850 161.925 ;
        RECT 84.080 161.910 84.400 161.970 ;
        RECT 84.555 161.925 84.845 162.155 ;
        RECT 86.010 161.770 86.150 162.310 ;
        RECT 90.520 162.110 90.840 162.170 ;
        RECT 94.750 162.155 94.890 162.310 ;
        RECT 94.215 162.110 94.505 162.155 ;
        RECT 90.520 161.970 94.505 162.110 ;
        RECT 90.520 161.910 90.840 161.970 ;
        RECT 94.215 161.925 94.505 161.970 ;
        RECT 94.675 162.110 94.965 162.155 ;
        RECT 96.515 162.110 96.805 162.155 ;
        RECT 96.960 162.110 97.280 162.170 ;
        RECT 101.575 162.110 101.865 162.155 ;
        RECT 94.675 161.970 101.865 162.110 ;
        RECT 94.675 161.925 94.965 161.970 ;
        RECT 96.515 161.925 96.805 161.970 ;
        RECT 96.960 161.910 97.280 161.970 ;
        RECT 101.575 161.925 101.865 161.970 ;
        RECT 81.870 161.630 86.150 161.770 ;
        RECT 88.220 161.570 88.540 161.830 ;
        RECT 78.550 161.430 78.840 161.475 ;
        RECT 75.290 161.290 78.840 161.430 ;
        RECT 75.290 161.245 75.580 161.290 ;
        RECT 76.720 161.230 77.040 161.290 ;
        RECT 78.550 161.245 78.840 161.290 ;
        RECT 79.470 161.430 79.760 161.475 ;
        RECT 81.330 161.430 81.620 161.475 ;
        RECT 79.470 161.290 81.620 161.430 ;
        RECT 79.470 161.245 79.760 161.290 ;
        RECT 81.330 161.245 81.620 161.290 ;
        RECT 91.900 161.430 92.220 161.490 ;
        RECT 97.435 161.430 97.725 161.475 ;
        RECT 91.900 161.290 97.725 161.430 ;
        RECT 102.570 161.430 102.710 162.650 ;
        RECT 104.780 162.590 105.100 162.850 ;
        RECT 103.860 162.450 104.180 162.510 ;
        RECT 105.255 162.450 105.545 162.495 ;
        RECT 103.860 162.310 105.545 162.450 ;
        RECT 103.860 162.250 104.180 162.310 ;
        RECT 105.255 162.265 105.545 162.310 ;
        RECT 107.080 162.110 107.400 162.170 ;
        RECT 109.855 162.110 110.145 162.155 ;
        RECT 110.760 162.110 111.080 162.170 ;
        RECT 107.080 161.970 109.150 162.110 ;
        RECT 107.080 161.910 107.400 161.970 ;
        RECT 102.940 161.570 103.260 161.830 ;
        RECT 109.010 161.815 109.150 161.970 ;
        RECT 109.855 161.970 111.080 162.110 ;
        RECT 109.855 161.925 110.145 161.970 ;
        RECT 110.760 161.910 111.080 161.970 ;
        RECT 108.015 161.585 108.305 161.815 ;
        RECT 108.935 161.770 109.225 161.815 ;
        RECT 110.300 161.770 110.620 161.830 ;
        RECT 108.935 161.630 110.620 161.770 ;
        RECT 108.935 161.585 109.225 161.630 ;
        RECT 108.090 161.430 108.230 161.585 ;
        RECT 110.300 161.570 110.620 161.630 ;
        RECT 102.570 161.290 108.230 161.430 ;
        RECT 91.900 161.230 92.220 161.290 ;
        RECT 97.435 161.245 97.725 161.290 ;
        RECT 64.315 160.950 65.540 161.090 ;
        RECT 64.315 160.905 64.605 160.950 ;
        RECT 65.220 160.890 65.540 160.950 ;
        RECT 66.155 160.905 66.445 161.135 ;
        RECT 67.060 161.090 67.380 161.150 ;
        RECT 67.995 161.090 68.285 161.135 ;
        RECT 67.060 160.950 68.285 161.090 ;
        RECT 67.060 160.890 67.380 160.950 ;
        RECT 67.995 160.905 68.285 160.950 ;
        RECT 70.295 161.090 70.585 161.135 ;
        RECT 71.200 161.090 71.520 161.150 ;
        RECT 70.295 160.950 71.520 161.090 ;
        RECT 70.295 160.905 70.585 160.950 ;
        RECT 71.200 160.890 71.520 160.950 ;
        RECT 72.580 160.890 72.900 161.150 ;
        RECT 84.540 161.090 84.860 161.150 ;
        RECT 85.015 161.090 85.305 161.135 ;
        RECT 84.540 160.950 85.305 161.090 ;
        RECT 84.540 160.890 84.860 160.950 ;
        RECT 85.015 160.905 85.305 160.950 ;
        RECT 93.755 161.090 94.045 161.135 ;
        RECT 94.660 161.090 94.980 161.150 ;
        RECT 93.755 160.950 94.980 161.090 ;
        RECT 93.755 160.905 94.045 160.950 ;
        RECT 94.660 160.890 94.980 160.950 ;
        RECT 97.895 161.090 98.185 161.135 ;
        RECT 102.480 161.090 102.800 161.150 ;
        RECT 97.895 160.950 102.800 161.090 ;
        RECT 97.895 160.905 98.185 160.950 ;
        RECT 102.480 160.890 102.800 160.950 ;
        RECT 15.010 160.270 113.450 160.750 ;
        RECT 17.840 159.870 18.160 160.130 ;
        RECT 22.900 160.070 23.220 160.130 ;
        RECT 19.770 159.930 23.220 160.070 ;
        RECT 16.920 159.390 17.240 159.450 ;
        RECT 18.315 159.390 18.605 159.435 ;
        RECT 16.920 159.250 18.605 159.390 ;
        RECT 16.920 159.190 17.240 159.250 ;
        RECT 18.315 159.205 18.605 159.250 ;
        RECT 19.770 159.095 19.910 159.930 ;
        RECT 22.900 159.870 23.220 159.930 ;
        RECT 24.280 159.870 24.600 160.130 ;
        RECT 53.735 160.070 54.025 160.115 ;
        RECT 54.640 160.070 54.960 160.130 ;
        RECT 53.735 159.930 54.960 160.070 ;
        RECT 53.735 159.885 54.025 159.930 ;
        RECT 54.640 159.870 54.960 159.930 ;
        RECT 63.840 160.070 64.160 160.130 ;
        RECT 66.600 160.070 66.920 160.130 ;
        RECT 67.520 160.070 67.840 160.130 ;
        RECT 63.840 159.930 66.920 160.070 ;
        RECT 63.840 159.870 64.160 159.930 ;
        RECT 66.600 159.870 66.920 159.930 ;
        RECT 67.150 159.930 67.840 160.070 ;
        RECT 20.155 159.730 20.445 159.775 ;
        RECT 22.440 159.730 22.760 159.790 ;
        RECT 27.960 159.730 28.280 159.790 ;
        RECT 31.180 159.775 31.500 159.790 ;
        RECT 20.155 159.590 28.280 159.730 ;
        RECT 20.155 159.545 20.445 159.590 ;
        RECT 22.440 159.530 22.760 159.590 ;
        RECT 27.960 159.530 28.280 159.590 ;
        RECT 31.130 159.730 31.500 159.775 ;
        RECT 34.390 159.730 34.680 159.775 ;
        RECT 31.130 159.590 34.680 159.730 ;
        RECT 31.130 159.545 31.500 159.590 ;
        RECT 34.390 159.545 34.680 159.590 ;
        RECT 35.310 159.730 35.600 159.775 ;
        RECT 37.170 159.730 37.460 159.775 ;
        RECT 39.920 159.730 40.240 159.790 ;
        RECT 47.280 159.730 47.600 159.790 ;
        RECT 35.310 159.590 37.460 159.730 ;
        RECT 35.310 159.545 35.600 159.590 ;
        RECT 37.170 159.545 37.460 159.590 ;
        RECT 37.710 159.590 39.690 159.730 ;
        RECT 31.180 159.530 31.500 159.545 ;
        RECT 20.615 159.390 20.905 159.435 ;
        RECT 21.060 159.390 21.380 159.450 ;
        RECT 23.375 159.390 23.665 159.435 ;
        RECT 20.615 159.250 21.380 159.390 ;
        RECT 20.615 159.205 20.905 159.250 ;
        RECT 21.060 159.190 21.380 159.250 ;
        RECT 22.530 159.250 23.665 159.390 ;
        RECT 19.695 158.865 19.985 159.095 ;
        RECT 22.530 158.755 22.670 159.250 ;
        RECT 23.375 159.205 23.665 159.250 ;
        RECT 32.990 159.390 33.280 159.435 ;
        RECT 35.310 159.390 35.525 159.545 ;
        RECT 32.990 159.250 35.525 159.390 ;
        RECT 35.780 159.390 36.100 159.450 ;
        RECT 37.710 159.390 37.850 159.590 ;
        RECT 35.780 159.250 37.850 159.390 ;
        RECT 32.990 159.205 33.280 159.250 ;
        RECT 35.780 159.190 36.100 159.250 ;
        RECT 38.080 159.190 38.400 159.450 ;
        RECT 39.550 159.435 39.690 159.590 ;
        RECT 39.920 159.590 43.830 159.730 ;
        RECT 39.920 159.530 40.240 159.590 ;
        RECT 39.475 159.205 39.765 159.435 ;
        RECT 42.695 159.205 42.985 159.435 ;
        RECT 36.255 159.050 36.545 159.095 ;
        RECT 36.255 158.910 38.770 159.050 ;
        RECT 36.255 158.865 36.545 158.910 ;
        RECT 38.630 158.755 38.770 158.910 ;
        RECT 42.770 158.770 42.910 159.205 ;
        RECT 43.140 159.190 43.460 159.450 ;
        RECT 43.690 159.435 43.830 159.590 ;
        RECT 45.070 159.590 47.600 159.730 ;
        RECT 43.615 159.205 43.905 159.435 ;
        RECT 44.520 159.390 44.840 159.450 ;
        RECT 45.070 159.435 45.210 159.590 ;
        RECT 47.280 159.530 47.600 159.590 ;
        RECT 54.180 159.730 54.500 159.790 ;
        RECT 55.115 159.730 55.405 159.775 ;
        RECT 65.680 159.730 66.000 159.790 ;
        RECT 54.180 159.590 55.405 159.730 ;
        RECT 54.180 159.530 54.500 159.590 ;
        RECT 55.115 159.545 55.405 159.590 ;
        RECT 63.930 159.590 66.000 159.730 ;
        RECT 44.995 159.390 45.285 159.435 ;
        RECT 44.520 159.250 45.285 159.390 ;
        RECT 44.520 159.190 44.840 159.250 ;
        RECT 44.995 159.205 45.285 159.250 ;
        RECT 45.900 159.190 46.220 159.450 ;
        RECT 46.375 159.205 46.665 159.435 ;
        RECT 46.835 159.205 47.125 159.435 ;
        RECT 43.230 159.050 43.370 159.190 ;
        RECT 46.450 159.050 46.590 159.205 ;
        RECT 43.230 158.910 46.590 159.050 ;
        RECT 46.910 159.050 47.050 159.205 ;
        RECT 50.960 159.190 51.280 159.450 ;
        RECT 55.560 159.390 55.880 159.450 ;
        RECT 56.495 159.390 56.785 159.435 ;
        RECT 55.560 159.250 56.785 159.390 ;
        RECT 55.560 159.190 55.880 159.250 ;
        RECT 56.495 159.205 56.785 159.250 ;
        RECT 56.940 159.390 57.260 159.450 ;
        RECT 57.875 159.390 58.165 159.435 ;
        RECT 56.940 159.250 58.165 159.390 ;
        RECT 56.940 159.190 57.260 159.250 ;
        RECT 57.875 159.205 58.165 159.250 ;
        RECT 59.715 159.390 60.005 159.435 ;
        RECT 60.160 159.390 60.480 159.450 ;
        RECT 59.715 159.250 60.480 159.390 ;
        RECT 59.715 159.205 60.005 159.250 ;
        RECT 60.160 159.190 60.480 159.250 ;
        RECT 61.540 159.190 61.860 159.450 ;
        RECT 63.930 159.435 64.070 159.590 ;
        RECT 65.680 159.530 66.000 159.590 ;
        RECT 63.855 159.205 64.145 159.435 ;
        RECT 65.220 159.190 65.540 159.450 ;
        RECT 66.140 159.435 66.460 159.450 ;
        RECT 66.130 159.205 66.460 159.435 ;
        RECT 66.140 159.190 66.460 159.205 ;
        RECT 66.600 159.190 66.920 159.450 ;
        RECT 67.150 159.435 67.290 159.930 ;
        RECT 67.520 159.870 67.840 159.930 ;
        RECT 69.360 160.070 69.680 160.130 ;
        RECT 79.495 160.070 79.785 160.115 ;
        RECT 80.400 160.070 80.720 160.130 ;
        RECT 69.360 159.930 72.350 160.070 ;
        RECT 69.360 159.870 69.680 159.930 ;
        RECT 69.820 159.730 70.140 159.790 ;
        RECT 71.660 159.730 71.980 159.790 ;
        RECT 69.820 159.590 71.980 159.730 ;
        RECT 72.210 159.730 72.350 159.930 ;
        RECT 79.495 159.930 80.720 160.070 ;
        RECT 79.495 159.885 79.785 159.930 ;
        RECT 80.400 159.870 80.720 159.930 ;
        RECT 80.860 159.870 81.180 160.130 ;
        RECT 94.215 160.070 94.505 160.115 ;
        RECT 94.660 160.070 94.980 160.130 ;
        RECT 94.215 159.930 94.980 160.070 ;
        RECT 94.215 159.885 94.505 159.930 ;
        RECT 94.660 159.870 94.980 159.930 ;
        RECT 102.480 160.070 102.800 160.130 ;
        RECT 104.335 160.070 104.625 160.115 ;
        RECT 102.480 159.930 104.625 160.070 ;
        RECT 102.480 159.870 102.800 159.930 ;
        RECT 104.335 159.885 104.625 159.930 ;
        RECT 85.000 159.730 85.320 159.790 ;
        RECT 72.210 159.590 85.320 159.730 ;
        RECT 69.820 159.530 70.140 159.590 ;
        RECT 71.660 159.530 71.980 159.590 ;
        RECT 85.000 159.530 85.320 159.590 ;
        RECT 97.970 159.590 102.250 159.730 ;
        RECT 67.075 159.205 67.365 159.435 ;
        RECT 68.440 159.390 68.760 159.450 ;
        RECT 70.295 159.390 70.585 159.435 ;
        RECT 68.440 159.250 70.585 159.390 ;
        RECT 68.440 159.240 68.900 159.250 ;
        RECT 68.440 159.190 68.760 159.240 ;
        RECT 70.295 159.205 70.585 159.250 ;
        RECT 70.755 159.205 71.045 159.435 ;
        RECT 58.320 159.050 58.640 159.110 ;
        RECT 46.910 158.910 58.640 159.050 ;
        RECT 22.455 158.525 22.745 158.755 ;
        RECT 32.990 158.710 33.280 158.755 ;
        RECT 35.770 158.710 36.060 158.755 ;
        RECT 37.630 158.710 37.920 158.755 ;
        RECT 32.990 158.570 37.920 158.710 ;
        RECT 32.990 158.525 33.280 158.570 ;
        RECT 35.770 158.525 36.060 158.570 ;
        RECT 37.630 158.525 37.920 158.570 ;
        RECT 38.555 158.525 38.845 158.755 ;
        RECT 42.680 158.710 43.000 158.770 ;
        RECT 46.910 158.710 47.050 158.910 ;
        RECT 58.320 158.850 58.640 158.910 ;
        RECT 69.820 159.050 70.140 159.110 ;
        RECT 70.830 159.050 70.970 159.205 ;
        RECT 71.200 159.190 71.520 159.450 ;
        RECT 72.135 159.205 72.425 159.435 ;
        RECT 72.580 159.390 72.900 159.450 ;
        RECT 78.575 159.390 78.865 159.435 ;
        RECT 72.580 159.250 78.865 159.390 ;
        RECT 69.820 158.910 70.970 159.050 ;
        RECT 69.820 158.850 70.140 158.910 ;
        RECT 42.680 158.570 47.050 158.710 ;
        RECT 47.280 158.710 47.600 158.770 ;
        RECT 65.220 158.710 65.540 158.770 ;
        RECT 72.210 158.710 72.350 159.205 ;
        RECT 72.580 159.190 72.900 159.250 ;
        RECT 78.575 159.205 78.865 159.250 ;
        RECT 79.480 159.390 79.800 159.450 ;
        RECT 80.415 159.390 80.705 159.435 ;
        RECT 79.480 159.250 80.705 159.390 ;
        RECT 79.480 159.190 79.800 159.250 ;
        RECT 80.415 159.205 80.705 159.250 ;
        RECT 80.490 159.050 80.630 159.205 ;
        RECT 81.780 159.190 82.100 159.450 ;
        RECT 91.455 159.390 91.745 159.435 ;
        RECT 91.900 159.390 92.220 159.450 ;
        RECT 91.455 159.250 92.220 159.390 ;
        RECT 91.455 159.205 91.745 159.250 ;
        RECT 91.900 159.190 92.220 159.250 ;
        RECT 94.660 159.390 94.980 159.450 ;
        RECT 97.970 159.435 98.110 159.590 ;
        RECT 97.895 159.390 98.185 159.435 ;
        RECT 94.660 159.250 98.185 159.390 ;
        RECT 94.660 159.190 94.980 159.250 ;
        RECT 97.895 159.205 98.185 159.250 ;
        RECT 98.340 159.190 98.660 159.450 ;
        RECT 98.815 159.390 99.105 159.435 ;
        RECT 99.260 159.390 99.580 159.450 ;
        RECT 98.815 159.250 99.580 159.390 ;
        RECT 98.815 159.205 99.105 159.250 ;
        RECT 99.260 159.190 99.580 159.250 ;
        RECT 99.720 159.390 100.040 159.450 ;
        RECT 102.110 159.435 102.250 159.590 ;
        RECT 99.720 159.250 101.790 159.390 ;
        RECT 99.720 159.190 100.040 159.250 ;
        RECT 83.160 159.050 83.480 159.110 ;
        RECT 80.490 158.910 83.480 159.050 ;
        RECT 83.160 158.850 83.480 158.910 ;
        RECT 90.520 159.050 90.840 159.110 ;
        RECT 100.655 159.050 100.945 159.095 ;
        RECT 90.520 158.910 100.945 159.050 ;
        RECT 101.650 159.050 101.790 159.250 ;
        RECT 102.035 159.205 102.325 159.435 ;
        RECT 102.480 159.190 102.800 159.450 ;
        RECT 102.955 159.390 103.245 159.435 ;
        RECT 103.400 159.390 103.720 159.450 ;
        RECT 102.955 159.250 103.720 159.390 ;
        RECT 102.955 159.205 103.245 159.250 ;
        RECT 103.400 159.190 103.720 159.250 ;
        RECT 103.875 159.205 104.165 159.435 ;
        RECT 104.780 159.390 105.100 159.450 ;
        RECT 108.935 159.390 109.225 159.435 ;
        RECT 104.780 159.250 109.225 159.390 ;
        RECT 103.950 159.050 104.090 159.205 ;
        RECT 104.780 159.190 105.100 159.250 ;
        RECT 108.935 159.205 109.225 159.250 ;
        RECT 110.300 159.190 110.620 159.450 ;
        RECT 110.760 159.190 111.080 159.450 ;
        RECT 101.650 158.910 104.090 159.050 ;
        RECT 90.520 158.850 90.840 158.910 ;
        RECT 100.655 158.865 100.945 158.910 ;
        RECT 107.095 158.865 107.385 159.095 ;
        RECT 72.580 158.710 72.900 158.770 ;
        RECT 47.280 158.570 72.900 158.710 ;
        RECT 42.680 158.510 43.000 158.570 ;
        RECT 47.280 158.510 47.600 158.570 ;
        RECT 65.220 158.510 65.540 158.570 ;
        RECT 72.580 158.510 72.900 158.570 ;
        RECT 98.340 158.710 98.660 158.770 ;
        RECT 102.020 158.710 102.340 158.770 ;
        RECT 107.170 158.710 107.310 158.865 ;
        RECT 98.340 158.570 107.310 158.710 ;
        RECT 98.340 158.510 98.660 158.570 ;
        RECT 102.020 158.510 102.340 158.570 ;
        RECT 29.125 158.370 29.415 158.415 ;
        RECT 32.100 158.370 32.420 158.430 ;
        RECT 29.125 158.230 32.420 158.370 ;
        RECT 29.125 158.185 29.415 158.230 ;
        RECT 32.100 158.170 32.420 158.230 ;
        RECT 39.460 158.370 39.780 158.430 ;
        RECT 41.315 158.370 41.605 158.415 ;
        RECT 39.460 158.230 41.605 158.370 ;
        RECT 39.460 158.170 39.780 158.230 ;
        RECT 41.315 158.185 41.605 158.230 ;
        RECT 46.820 158.370 47.140 158.430 ;
        RECT 48.215 158.370 48.505 158.415 ;
        RECT 46.820 158.230 48.505 158.370 ;
        RECT 46.820 158.170 47.140 158.230 ;
        RECT 48.215 158.185 48.505 158.230 ;
        RECT 57.400 158.170 57.720 158.430 ;
        RECT 58.780 158.170 59.100 158.430 ;
        RECT 60.620 158.170 60.940 158.430 ;
        RECT 62.000 158.370 62.320 158.430 ;
        RECT 62.935 158.370 63.225 158.415 ;
        RECT 62.000 158.230 63.225 158.370 ;
        RECT 62.000 158.170 62.320 158.230 ;
        RECT 62.935 158.185 63.225 158.230 ;
        RECT 68.440 158.170 68.760 158.430 ;
        RECT 68.915 158.370 69.205 158.415 ;
        RECT 69.360 158.370 69.680 158.430 ;
        RECT 68.915 158.230 69.680 158.370 ;
        RECT 68.915 158.185 69.205 158.230 ;
        RECT 69.360 158.170 69.680 158.230 ;
        RECT 88.220 158.170 88.540 158.430 ;
        RECT 95.580 158.370 95.900 158.430 ;
        RECT 96.515 158.370 96.805 158.415 ;
        RECT 95.580 158.230 96.805 158.370 ;
        RECT 95.580 158.170 95.900 158.230 ;
        RECT 96.515 158.185 96.805 158.230 ;
        RECT 98.800 158.370 99.120 158.430 ;
        RECT 102.480 158.370 102.800 158.430 ;
        RECT 98.800 158.230 102.800 158.370 ;
        RECT 98.800 158.170 99.120 158.230 ;
        RECT 102.480 158.170 102.800 158.230 ;
        RECT 109.840 158.370 110.160 158.430 ;
        RECT 111.235 158.370 111.525 158.415 ;
        RECT 109.840 158.230 111.525 158.370 ;
        RECT 109.840 158.170 110.160 158.230 ;
        RECT 111.235 158.185 111.525 158.230 ;
        RECT 15.010 157.550 113.450 158.030 ;
        RECT 32.560 157.350 32.880 157.410 ;
        RECT 37.160 157.350 37.480 157.410 ;
        RECT 40.840 157.350 41.160 157.410 ;
        RECT 44.520 157.350 44.840 157.410 ;
        RECT 59.700 157.350 60.020 157.410 ;
        RECT 85.460 157.350 85.780 157.410 ;
        RECT 32.560 157.210 44.840 157.350 ;
        RECT 32.560 157.150 32.880 157.210 ;
        RECT 37.160 157.150 37.480 157.210 ;
        RECT 40.840 157.150 41.160 157.210 ;
        RECT 44.520 157.150 44.840 157.210 ;
        RECT 45.070 157.210 60.020 157.350 ;
        RECT 20.570 157.010 20.860 157.055 ;
        RECT 23.350 157.010 23.640 157.055 ;
        RECT 25.210 157.010 25.500 157.055 ;
        RECT 20.570 156.870 25.500 157.010 ;
        RECT 20.570 156.825 20.860 156.870 ;
        RECT 23.350 156.825 23.640 156.870 ;
        RECT 25.210 156.825 25.500 156.870 ;
        RECT 42.220 157.010 42.540 157.070 ;
        RECT 45.070 157.010 45.210 157.210 ;
        RECT 59.700 157.150 60.020 157.210 ;
        RECT 67.610 157.210 85.780 157.350 ;
        RECT 42.220 156.870 45.210 157.010 ;
        RECT 55.990 157.010 56.280 157.055 ;
        RECT 58.770 157.010 59.060 157.055 ;
        RECT 60.630 157.010 60.920 157.055 ;
        RECT 62.015 157.010 62.305 157.055 ;
        RECT 55.990 156.870 60.920 157.010 ;
        RECT 42.220 156.810 42.540 156.870 ;
        RECT 55.990 156.825 56.280 156.870 ;
        RECT 58.770 156.825 59.060 156.870 ;
        RECT 60.630 156.825 60.920 156.870 ;
        RECT 61.135 156.870 62.305 157.010 ;
        RECT 16.705 156.670 16.995 156.715 ;
        RECT 21.060 156.670 21.380 156.730 ;
        RECT 16.705 156.530 21.380 156.670 ;
        RECT 16.705 156.485 16.995 156.530 ;
        RECT 21.060 156.470 21.380 156.530 ;
        RECT 27.960 156.670 28.280 156.730 ;
        RECT 31.180 156.670 31.500 156.730 ;
        RECT 36.240 156.670 36.560 156.730 ;
        RECT 43.140 156.670 43.460 156.730 ;
        RECT 61.135 156.670 61.275 156.870 ;
        RECT 62.015 156.825 62.305 156.870 ;
        RECT 62.460 157.010 62.780 157.070 ;
        RECT 67.610 157.010 67.750 157.210 ;
        RECT 85.460 157.150 85.780 157.210 ;
        RECT 89.600 157.350 89.920 157.410 ;
        RECT 96.040 157.350 96.360 157.410 ;
        RECT 89.600 157.210 96.360 157.350 ;
        RECT 89.600 157.150 89.920 157.210 ;
        RECT 96.040 157.150 96.360 157.210 ;
        RECT 104.320 157.350 104.640 157.410 ;
        RECT 104.320 157.210 111.450 157.350 ;
        RECT 104.320 157.150 104.640 157.210 ;
        RECT 62.460 156.870 67.750 157.010 ;
        RECT 67.980 157.010 68.300 157.070 ;
        RECT 91.900 157.010 92.220 157.070 ;
        RECT 98.800 157.010 99.120 157.070 ;
        RECT 67.980 156.870 83.850 157.010 ;
        RECT 62.460 156.810 62.780 156.870 ;
        RECT 67.980 156.810 68.300 156.870 ;
        RECT 27.960 156.530 30.950 156.670 ;
        RECT 27.960 156.470 28.280 156.530 ;
        RECT 20.570 156.330 20.860 156.375 ;
        RECT 23.360 156.330 23.680 156.390 ;
        RECT 23.835 156.330 24.125 156.375 ;
        RECT 20.570 156.190 23.105 156.330 ;
        RECT 20.570 156.145 20.860 156.190 ;
        RECT 18.710 155.990 19.000 156.035 ;
        RECT 20.140 155.990 20.460 156.050 ;
        RECT 22.890 156.035 23.105 156.190 ;
        RECT 23.360 156.190 24.125 156.330 ;
        RECT 23.360 156.130 23.680 156.190 ;
        RECT 23.835 156.145 24.125 156.190 ;
        RECT 25.675 156.330 25.965 156.375 ;
        RECT 26.580 156.330 26.900 156.390 ;
        RECT 25.675 156.190 26.900 156.330 ;
        RECT 25.675 156.145 25.965 156.190 ;
        RECT 26.580 156.130 26.900 156.190 ;
        RECT 29.800 156.130 30.120 156.390 ;
        RECT 30.810 156.375 30.950 156.530 ;
        RECT 31.180 156.530 33.250 156.670 ;
        RECT 31.180 156.470 31.500 156.530 ;
        RECT 30.275 156.145 30.565 156.375 ;
        RECT 30.735 156.145 31.025 156.375 ;
        RECT 21.970 155.990 22.260 156.035 ;
        RECT 18.710 155.850 22.260 155.990 ;
        RECT 18.710 155.805 19.000 155.850 ;
        RECT 20.140 155.790 20.460 155.850 ;
        RECT 21.970 155.805 22.260 155.850 ;
        RECT 22.890 155.990 23.180 156.035 ;
        RECT 24.750 155.990 25.040 156.035 ;
        RECT 22.890 155.850 25.040 155.990 ;
        RECT 22.890 155.805 23.180 155.850 ;
        RECT 24.750 155.805 25.040 155.850 ;
        RECT 28.420 155.450 28.740 155.710 ;
        RECT 30.350 155.650 30.490 156.145 ;
        RECT 31.640 156.130 31.960 156.390 ;
        RECT 32.115 156.330 32.405 156.375 ;
        RECT 32.560 156.330 32.880 156.390 ;
        RECT 33.110 156.375 33.250 156.530 ;
        RECT 33.570 156.530 43.460 156.670 ;
        RECT 33.570 156.375 33.710 156.530 ;
        RECT 36.240 156.470 36.560 156.530 ;
        RECT 32.115 156.190 32.880 156.330 ;
        RECT 32.115 156.145 32.405 156.190 ;
        RECT 32.560 156.130 32.880 156.190 ;
        RECT 33.035 156.145 33.325 156.375 ;
        RECT 33.495 156.145 33.785 156.375 ;
        RECT 33.955 156.145 34.245 156.375 ;
        RECT 34.030 155.990 34.170 156.145 ;
        RECT 37.160 156.130 37.480 156.390 ;
        RECT 37.620 156.330 37.940 156.390 ;
        RECT 38.630 156.375 38.770 156.530 ;
        RECT 38.095 156.330 38.385 156.375 ;
        RECT 37.620 156.190 38.385 156.330 ;
        RECT 37.620 156.130 37.940 156.190 ;
        RECT 38.095 156.145 38.385 156.190 ;
        RECT 38.555 156.145 38.845 156.375 ;
        RECT 39.015 156.145 39.305 156.375 ;
        RECT 39.090 155.990 39.230 156.145 ;
        RECT 40.840 156.130 41.160 156.390 ;
        RECT 41.760 156.130 42.080 156.390 ;
        RECT 42.310 156.375 42.450 156.530 ;
        RECT 43.140 156.470 43.460 156.530 ;
        RECT 60.250 156.530 61.275 156.670 ;
        RECT 63.840 156.670 64.160 156.730 ;
        RECT 69.820 156.670 70.140 156.730 ;
        RECT 73.040 156.670 73.360 156.730 ;
        RECT 63.840 156.530 66.830 156.670 ;
        RECT 42.235 156.145 42.525 156.375 ;
        RECT 42.680 156.130 43.000 156.390 ;
        RECT 55.990 156.330 56.280 156.375 ;
        RECT 59.255 156.330 59.545 156.375 ;
        RECT 60.250 156.330 60.390 156.530 ;
        RECT 63.840 156.470 64.160 156.530 ;
        RECT 55.990 156.190 58.525 156.330 ;
        RECT 55.990 156.145 56.280 156.190 ;
        RECT 34.030 155.850 39.230 155.990 ;
        RECT 31.180 155.650 31.500 155.710 ;
        RECT 30.350 155.510 31.500 155.650 ;
        RECT 31.180 155.450 31.500 155.510 ;
        RECT 35.335 155.650 35.625 155.695 ;
        RECT 35.780 155.650 36.100 155.710 ;
        RECT 35.335 155.510 36.100 155.650 ;
        RECT 35.335 155.465 35.625 155.510 ;
        RECT 35.780 155.450 36.100 155.510 ;
        RECT 38.080 155.650 38.400 155.710 ;
        RECT 39.090 155.650 39.230 155.850 ;
        RECT 40.395 155.990 40.685 156.035 ;
        RECT 43.600 155.990 43.920 156.050 ;
        RECT 57.400 156.035 57.720 156.050 ;
        RECT 40.395 155.850 43.920 155.990 ;
        RECT 40.395 155.805 40.685 155.850 ;
        RECT 43.600 155.790 43.920 155.850 ;
        RECT 54.130 155.990 54.420 156.035 ;
        RECT 57.390 155.990 57.720 156.035 ;
        RECT 54.130 155.850 57.720 155.990 ;
        RECT 54.130 155.805 54.420 155.850 ;
        RECT 57.390 155.805 57.720 155.850 ;
        RECT 58.310 156.035 58.525 156.190 ;
        RECT 59.255 156.190 60.390 156.330 ;
        RECT 59.255 156.145 59.545 156.190 ;
        RECT 61.080 156.130 61.400 156.390 ;
        RECT 62.935 156.145 63.225 156.375 ;
        RECT 63.435 156.330 63.725 156.375 ;
        RECT 64.300 156.330 64.620 156.390 ;
        RECT 63.435 156.190 64.620 156.330 ;
        RECT 63.435 156.145 63.725 156.190 ;
        RECT 58.310 155.990 58.600 156.035 ;
        RECT 60.170 155.990 60.460 156.035 ;
        RECT 58.310 155.850 60.460 155.990 ;
        RECT 58.310 155.805 58.600 155.850 ;
        RECT 60.170 155.805 60.460 155.850 ;
        RECT 61.540 155.990 61.860 156.050 ;
        RECT 63.010 155.990 63.150 156.145 ;
        RECT 64.300 156.130 64.620 156.190 ;
        RECT 64.760 156.130 65.080 156.390 ;
        RECT 65.220 156.330 65.540 156.390 ;
        RECT 66.690 156.375 66.830 156.530 ;
        RECT 67.150 156.530 71.430 156.670 ;
        RECT 67.150 156.390 67.290 156.530 ;
        RECT 69.820 156.470 70.140 156.530 ;
        RECT 65.695 156.330 65.985 156.375 ;
        RECT 65.220 156.190 65.985 156.330 ;
        RECT 65.220 156.130 65.540 156.190 ;
        RECT 65.695 156.145 65.985 156.190 ;
        RECT 66.615 156.145 66.905 156.375 ;
        RECT 67.060 156.130 67.380 156.390 ;
        RECT 67.520 156.330 67.840 156.390 ;
        RECT 71.290 156.375 71.430 156.530 ;
        RECT 71.750 156.530 73.360 156.670 ;
        RECT 71.750 156.375 71.890 156.530 ;
        RECT 73.040 156.470 73.360 156.530 ;
        RECT 70.755 156.330 71.045 156.375 ;
        RECT 67.520 156.190 71.045 156.330 ;
        RECT 67.520 156.130 67.840 156.190 ;
        RECT 70.755 156.145 71.045 156.190 ;
        RECT 71.215 156.145 71.505 156.375 ;
        RECT 71.675 156.145 71.965 156.375 ;
        RECT 72.580 156.130 72.900 156.390 ;
        RECT 83.710 156.375 83.850 156.870 ;
        RECT 91.070 156.870 92.220 157.010 ;
        RECT 83.635 156.145 83.925 156.375 ;
        RECT 61.540 155.850 63.150 155.990 ;
        RECT 63.855 155.990 64.145 156.035 ;
        RECT 68.915 155.990 69.205 156.035 ;
        RECT 83.710 155.990 83.850 156.145 ;
        RECT 84.540 156.130 84.860 156.390 ;
        RECT 85.000 156.130 85.320 156.390 ;
        RECT 85.460 156.130 85.780 156.390 ;
        RECT 89.600 156.330 89.920 156.390 ;
        RECT 91.070 156.375 91.210 156.870 ;
        RECT 91.900 156.810 92.220 156.870 ;
        RECT 92.910 156.870 99.120 157.010 ;
        RECT 92.910 156.670 93.050 156.870 ;
        RECT 94.660 156.670 94.980 156.730 ;
        RECT 91.530 156.530 93.050 156.670 ;
        RECT 93.370 156.530 95.350 156.670 ;
        RECT 91.530 156.375 91.670 156.530 ;
        RECT 90.075 156.330 90.365 156.375 ;
        RECT 86.010 156.190 90.365 156.330 ;
        RECT 86.010 155.990 86.150 156.190 ;
        RECT 89.600 156.130 89.920 156.190 ;
        RECT 90.075 156.145 90.365 156.190 ;
        RECT 90.995 156.145 91.285 156.375 ;
        RECT 91.455 156.145 91.745 156.375 ;
        RECT 91.900 156.330 92.220 156.390 ;
        RECT 93.370 156.330 93.510 156.530 ;
        RECT 94.660 156.470 94.980 156.530 ;
        RECT 95.210 156.375 95.350 156.530 ;
        RECT 95.670 156.375 95.810 156.870 ;
        RECT 98.800 156.810 99.120 156.870 ;
        RECT 105.815 157.010 106.105 157.055 ;
        RECT 108.935 157.010 109.225 157.055 ;
        RECT 110.825 157.010 111.115 157.055 ;
        RECT 105.815 156.870 111.115 157.010 ;
        RECT 105.815 156.825 106.105 156.870 ;
        RECT 108.935 156.825 109.225 156.870 ;
        RECT 110.825 156.825 111.115 156.870 ;
        RECT 111.310 156.670 111.450 157.210 ;
        RECT 111.695 156.670 111.985 156.715 ;
        RECT 111.310 156.530 111.985 156.670 ;
        RECT 111.695 156.485 111.985 156.530 ;
        RECT 91.900 156.190 93.510 156.330 ;
        RECT 91.530 155.990 91.670 156.145 ;
        RECT 91.900 156.130 92.220 156.190 ;
        RECT 95.135 156.145 95.425 156.375 ;
        RECT 95.595 156.145 95.885 156.375 ;
        RECT 96.040 156.130 96.360 156.390 ;
        RECT 96.960 156.330 97.280 156.390 ;
        RECT 99.260 156.330 99.580 156.390 ;
        RECT 96.960 156.190 99.580 156.330 ;
        RECT 96.960 156.130 97.280 156.190 ;
        RECT 99.260 156.130 99.580 156.190 ;
        RECT 99.735 156.330 100.025 156.375 ;
        RECT 99.735 156.190 101.330 156.330 ;
        RECT 99.735 156.145 100.025 156.190 ;
        RECT 63.855 155.850 65.910 155.990 ;
        RECT 57.400 155.790 57.720 155.805 ;
        RECT 61.540 155.790 61.860 155.850 ;
        RECT 63.855 155.805 64.145 155.850 ;
        RECT 65.770 155.710 65.910 155.850 ;
        RECT 68.915 155.850 72.810 155.990 ;
        RECT 83.710 155.850 86.150 155.990 ;
        RECT 86.470 155.850 91.670 155.990 ;
        RECT 68.915 155.805 69.205 155.850 ;
        RECT 72.670 155.710 72.810 155.850 ;
        RECT 42.680 155.650 43.000 155.710 ;
        RECT 38.080 155.510 43.000 155.650 ;
        RECT 38.080 155.450 38.400 155.510 ;
        RECT 42.680 155.450 43.000 155.510 ;
        RECT 43.140 155.650 43.460 155.710 ;
        RECT 44.075 155.650 44.365 155.695 ;
        RECT 43.140 155.510 44.365 155.650 ;
        RECT 43.140 155.450 43.460 155.510 ;
        RECT 44.075 155.465 44.365 155.510 ;
        RECT 52.125 155.650 52.415 155.695 ;
        RECT 55.100 155.650 55.420 155.710 ;
        RECT 52.125 155.510 55.420 155.650 ;
        RECT 52.125 155.465 52.415 155.510 ;
        RECT 55.100 155.450 55.420 155.510 ;
        RECT 65.680 155.450 66.000 155.710 ;
        RECT 69.375 155.650 69.665 155.695 ;
        RECT 69.820 155.650 70.140 155.710 ;
        RECT 69.375 155.510 70.140 155.650 ;
        RECT 69.375 155.465 69.665 155.510 ;
        RECT 69.820 155.450 70.140 155.510 ;
        RECT 72.580 155.450 72.900 155.710 ;
        RECT 85.000 155.650 85.320 155.710 ;
        RECT 86.470 155.650 86.610 155.850 ;
        RECT 93.740 155.790 94.060 156.050 ;
        RECT 101.190 155.710 101.330 156.190 ;
        RECT 102.495 155.990 102.785 156.035 ;
        RECT 103.860 155.990 104.180 156.050 ;
        RECT 104.735 156.035 105.025 156.350 ;
        RECT 105.815 156.330 106.105 156.375 ;
        RECT 109.395 156.330 109.685 156.375 ;
        RECT 111.230 156.330 111.520 156.375 ;
        RECT 105.815 156.190 111.520 156.330 ;
        RECT 105.815 156.145 106.105 156.190 ;
        RECT 109.395 156.145 109.685 156.190 ;
        RECT 111.230 156.145 111.520 156.190 ;
        RECT 102.495 155.850 104.180 155.990 ;
        RECT 102.495 155.805 102.785 155.850 ;
        RECT 103.860 155.790 104.180 155.850 ;
        RECT 104.435 155.990 105.025 156.035 ;
        RECT 107.675 155.990 108.325 156.035 ;
        RECT 109.840 155.990 110.160 156.050 ;
        RECT 104.435 155.850 110.160 155.990 ;
        RECT 104.435 155.805 104.725 155.850 ;
        RECT 107.675 155.805 108.325 155.850 ;
        RECT 109.840 155.790 110.160 155.850 ;
        RECT 110.300 155.790 110.620 156.050 ;
        RECT 85.000 155.510 86.610 155.650 ;
        RECT 86.855 155.650 87.145 155.695 ;
        RECT 88.680 155.650 89.000 155.710 ;
        RECT 86.855 155.510 89.000 155.650 ;
        RECT 85.000 155.450 85.320 155.510 ;
        RECT 86.855 155.465 87.145 155.510 ;
        RECT 88.680 155.450 89.000 155.510 ;
        RECT 93.280 155.450 93.600 155.710 ;
        RECT 101.100 155.650 101.420 155.710 ;
        RECT 102.955 155.650 103.245 155.695 ;
        RECT 101.100 155.510 103.245 155.650 ;
        RECT 101.100 155.450 101.420 155.510 ;
        RECT 102.955 155.465 103.245 155.510 ;
        RECT 15.010 154.830 113.450 155.310 ;
        RECT 26.135 154.630 26.425 154.675 ;
        RECT 39.000 154.630 39.320 154.690 ;
        RECT 58.780 154.630 59.100 154.690 ;
        RECT 26.135 154.490 33.710 154.630 ;
        RECT 26.135 154.445 26.425 154.490 ;
        RECT 20.600 154.290 20.920 154.350 ;
        RECT 26.210 154.290 26.350 154.445 ;
        RECT 20.600 154.150 26.350 154.290 ;
        RECT 31.180 154.290 31.500 154.350 ;
        RECT 31.180 154.150 33.250 154.290 ;
        RECT 20.600 154.090 20.920 154.150 ;
        RECT 31.180 154.090 31.500 154.150 ;
        RECT 33.110 154.010 33.250 154.150 ;
        RECT 25.675 153.950 25.965 153.995 ;
        RECT 26.120 153.950 26.440 154.010 ;
        RECT 25.675 153.810 26.440 153.950 ;
        RECT 25.675 153.765 25.965 153.810 ;
        RECT 26.120 153.750 26.440 153.810 ;
        RECT 29.800 153.950 30.120 154.010 ;
        RECT 32.560 153.950 32.880 154.010 ;
        RECT 29.800 153.810 32.880 153.950 ;
        RECT 29.800 153.750 30.120 153.810 ;
        RECT 32.560 153.750 32.880 153.810 ;
        RECT 33.020 153.750 33.340 154.010 ;
        RECT 33.570 153.995 33.710 154.490 ;
        RECT 34.490 154.490 59.100 154.630 ;
        RECT 34.490 153.995 34.630 154.490 ;
        RECT 39.000 154.430 39.320 154.490 ;
        RECT 58.780 154.430 59.100 154.490 ;
        RECT 60.160 154.630 60.480 154.690 ;
        RECT 68.900 154.630 69.220 154.690 ;
        RECT 104.780 154.630 105.100 154.690 ;
        RECT 60.160 154.490 66.830 154.630 ;
        RECT 60.160 154.430 60.480 154.490 ;
        RECT 38.080 154.290 38.400 154.350 ;
        RECT 36.790 154.150 38.400 154.290 ;
        RECT 33.495 153.765 33.785 153.995 ;
        RECT 34.415 153.765 34.705 153.995 ;
        RECT 21.060 153.410 21.380 153.670 ;
        RECT 21.995 153.610 22.285 153.655 ;
        RECT 22.900 153.610 23.220 153.670 ;
        RECT 26.595 153.610 26.885 153.655 ;
        RECT 27.960 153.610 28.280 153.670 ;
        RECT 21.995 153.470 28.280 153.610 ;
        RECT 21.995 153.425 22.285 153.470 ;
        RECT 22.900 153.410 23.220 153.470 ;
        RECT 26.595 153.425 26.885 153.470 ;
        RECT 27.960 153.410 28.280 153.470 ;
        RECT 31.640 153.610 31.960 153.670 ;
        RECT 34.490 153.610 34.630 153.765 ;
        RECT 34.860 153.750 35.180 154.010 ;
        RECT 35.795 153.765 36.085 153.995 ;
        RECT 31.640 153.470 34.630 153.610 ;
        RECT 31.640 153.410 31.960 153.470 ;
        RECT 21.150 153.270 21.290 153.410 ;
        RECT 35.870 153.270 36.010 153.765 ;
        RECT 36.240 153.750 36.560 154.010 ;
        RECT 36.790 153.995 36.930 154.150 ;
        RECT 38.080 154.090 38.400 154.150 ;
        RECT 47.755 154.290 48.045 154.335 ;
        RECT 50.615 154.290 50.905 154.335 ;
        RECT 53.855 154.290 54.505 154.335 ;
        RECT 47.755 154.150 54.505 154.290 ;
        RECT 47.755 154.105 48.045 154.150 ;
        RECT 50.615 154.105 51.205 154.150 ;
        RECT 53.855 154.105 54.505 154.150 ;
        RECT 55.100 154.290 55.420 154.350 ;
        RECT 56.020 154.290 56.340 154.350 ;
        RECT 55.100 154.150 64.530 154.290 ;
        RECT 36.715 153.765 37.005 153.995 ;
        RECT 37.160 153.950 37.480 154.010 ;
        RECT 38.555 153.950 38.845 153.995 ;
        RECT 37.160 153.810 38.845 153.950 ;
        RECT 37.160 153.750 37.480 153.810 ;
        RECT 38.555 153.765 38.845 153.810 ;
        RECT 39.475 153.765 39.765 153.995 ;
        RECT 38.080 153.410 38.400 153.670 ;
        RECT 39.550 153.270 39.690 153.765 ;
        RECT 39.920 153.750 40.240 154.010 ;
        RECT 40.395 153.950 40.685 153.995 ;
        RECT 42.220 153.950 42.540 154.010 ;
        RECT 40.395 153.810 42.540 153.950 ;
        RECT 40.395 153.765 40.685 153.810 ;
        RECT 21.150 153.130 36.010 153.270 ;
        RECT 36.330 153.130 39.690 153.270 ;
        RECT 18.775 152.930 19.065 152.975 ;
        RECT 19.680 152.930 20.000 152.990 ;
        RECT 18.775 152.790 20.000 152.930 ;
        RECT 18.775 152.745 19.065 152.790 ;
        RECT 19.680 152.730 20.000 152.790 ;
        RECT 23.820 152.730 24.140 152.990 ;
        RECT 31.180 152.730 31.500 152.990 ;
        RECT 32.100 152.930 32.420 152.990 ;
        RECT 36.330 152.930 36.470 153.130 ;
        RECT 32.100 152.790 36.470 152.930 ;
        RECT 37.620 152.930 37.940 152.990 ;
        RECT 40.470 152.930 40.610 153.765 ;
        RECT 42.220 153.750 42.540 153.810 ;
        RECT 47.295 153.765 47.585 153.995 ;
        RECT 50.915 153.790 51.205 154.105 ;
        RECT 55.100 154.090 55.420 154.150 ;
        RECT 56.020 154.090 56.340 154.150 ;
        RECT 58.870 153.995 59.010 154.150 ;
        RECT 51.995 153.950 52.285 153.995 ;
        RECT 55.575 153.950 55.865 153.995 ;
        RECT 57.410 153.950 57.700 153.995 ;
        RECT 51.995 153.810 57.700 153.950 ;
        RECT 51.995 153.765 52.285 153.810 ;
        RECT 55.575 153.765 55.865 153.810 ;
        RECT 57.410 153.765 57.700 153.810 ;
        RECT 58.795 153.765 59.085 153.995 ;
        RECT 41.760 153.610 42.080 153.670 ;
        RECT 47.370 153.610 47.510 153.765 ;
        RECT 63.380 153.750 63.700 154.010 ;
        RECT 63.840 153.750 64.160 154.010 ;
        RECT 64.390 153.995 64.530 154.150 ;
        RECT 66.690 154.010 66.830 154.490 ;
        RECT 68.900 154.490 70.740 154.630 ;
        RECT 68.900 154.430 69.220 154.490 ;
        RECT 67.535 154.290 67.825 154.335 ;
        RECT 67.980 154.290 68.300 154.350 ;
        RECT 68.455 154.290 68.745 154.335 ;
        RECT 67.535 154.150 68.745 154.290 ;
        RECT 70.600 154.290 70.740 154.490 ;
        RECT 79.570 154.490 105.100 154.630 ;
        RECT 70.600 154.150 71.430 154.290 ;
        RECT 67.535 154.105 67.825 154.150 ;
        RECT 67.980 154.090 68.300 154.150 ;
        RECT 68.455 154.105 68.745 154.150 ;
        RECT 64.315 153.765 64.605 153.995 ;
        RECT 65.220 153.750 65.540 154.010 ;
        RECT 66.600 153.950 66.920 154.010 ;
        RECT 68.915 153.950 69.205 153.995 ;
        RECT 66.600 153.810 69.205 153.950 ;
        RECT 66.600 153.750 66.920 153.810 ;
        RECT 68.915 153.765 69.205 153.810 ;
        RECT 70.280 153.950 70.600 154.010 ;
        RECT 71.290 153.995 71.430 154.150 ;
        RECT 79.570 153.995 79.710 154.490 ;
        RECT 84.540 154.090 84.860 154.350 ;
        RECT 86.840 154.335 87.160 154.350 ;
        RECT 86.835 154.290 87.485 154.335 ;
        RECT 90.435 154.290 90.725 154.335 ;
        RECT 86.835 154.150 90.725 154.290 ;
        RECT 86.835 154.105 87.485 154.150 ;
        RECT 90.135 154.105 90.725 154.150 ;
        RECT 86.840 154.090 87.160 154.105 ;
        RECT 70.755 153.950 71.045 153.995 ;
        RECT 70.280 153.810 71.045 153.950 ;
        RECT 70.280 153.750 70.600 153.810 ;
        RECT 70.755 153.765 71.045 153.810 ;
        RECT 71.215 153.765 71.505 153.995 ;
        RECT 78.115 153.950 78.405 153.995 ;
        RECT 79.495 153.950 79.785 153.995 ;
        RECT 78.115 153.810 79.785 153.950 ;
        RECT 78.115 153.765 78.405 153.810 ;
        RECT 79.495 153.765 79.785 153.810 ;
        RECT 80.400 153.950 80.720 154.010 ;
        RECT 80.875 153.950 81.165 153.995 ;
        RECT 80.400 153.810 81.165 153.950 ;
        RECT 80.400 153.750 80.720 153.810 ;
        RECT 80.875 153.765 81.165 153.810 ;
        RECT 83.640 153.950 83.930 153.995 ;
        RECT 85.475 153.950 85.765 153.995 ;
        RECT 89.055 153.950 89.345 153.995 ;
        RECT 83.640 153.810 89.345 153.950 ;
        RECT 83.640 153.765 83.930 153.810 ;
        RECT 85.475 153.765 85.765 153.810 ;
        RECT 89.055 153.765 89.345 153.810 ;
        RECT 90.135 153.790 90.425 154.105 ;
        RECT 54.180 153.610 54.500 153.670 ;
        RECT 41.760 153.470 54.500 153.610 ;
        RECT 41.760 153.410 42.080 153.470 ;
        RECT 54.180 153.410 54.500 153.470 ;
        RECT 56.480 153.410 56.800 153.670 ;
        RECT 57.875 153.610 58.165 153.655 ;
        RECT 61.080 153.610 61.400 153.670 ;
        RECT 57.875 153.470 61.400 153.610 ;
        RECT 57.875 153.425 58.165 153.470 ;
        RECT 61.080 153.410 61.400 153.470 ;
        RECT 61.555 153.610 61.845 153.655 ;
        RECT 64.760 153.610 65.080 153.670 ;
        RECT 61.555 153.470 65.080 153.610 ;
        RECT 61.555 153.425 61.845 153.470 ;
        RECT 64.760 153.410 65.080 153.470 ;
        RECT 66.140 153.610 66.460 153.670 ;
        RECT 69.375 153.610 69.665 153.655 ;
        RECT 66.140 153.470 69.665 153.610 ;
        RECT 66.140 153.410 66.460 153.470 ;
        RECT 69.375 153.425 69.665 153.470 ;
        RECT 83.175 153.610 83.465 153.655 ;
        RECT 88.220 153.610 88.540 153.670 ;
        RECT 83.175 153.470 88.540 153.610 ;
        RECT 83.175 153.425 83.465 153.470 ;
        RECT 88.220 153.410 88.540 153.470 ;
        RECT 51.995 153.270 52.285 153.315 ;
        RECT 55.115 153.270 55.405 153.315 ;
        RECT 57.005 153.270 57.295 153.315 ;
        RECT 60.160 153.270 60.480 153.330 ;
        RECT 51.995 153.130 57.295 153.270 ;
        RECT 51.995 153.085 52.285 153.130 ;
        RECT 55.115 153.085 55.405 153.130 ;
        RECT 57.005 153.085 57.295 153.130 ;
        RECT 57.490 153.130 60.480 153.270 ;
        RECT 57.490 152.990 57.630 153.130 ;
        RECT 60.160 153.070 60.480 153.130 ;
        RECT 62.000 153.070 62.320 153.330 ;
        RECT 63.840 153.270 64.160 153.330 ;
        RECT 72.135 153.270 72.425 153.315 ;
        RECT 76.720 153.270 77.040 153.330 ;
        RECT 63.840 153.130 77.040 153.270 ;
        RECT 63.840 153.070 64.160 153.130 ;
        RECT 72.135 153.085 72.425 153.130 ;
        RECT 76.720 153.070 77.040 153.130 ;
        RECT 77.655 153.270 77.945 153.315 ;
        RECT 79.940 153.270 80.260 153.330 ;
        RECT 77.655 153.130 80.260 153.270 ;
        RECT 77.655 153.085 77.945 153.130 ;
        RECT 79.940 153.070 80.260 153.130 ;
        RECT 84.045 153.270 84.335 153.315 ;
        RECT 85.935 153.270 86.225 153.315 ;
        RECT 89.055 153.270 89.345 153.315 ;
        RECT 84.045 153.130 89.345 153.270 ;
        RECT 84.045 153.085 84.335 153.130 ;
        RECT 85.935 153.085 86.225 153.130 ;
        RECT 89.055 153.085 89.345 153.130 ;
        RECT 91.070 152.990 91.210 154.490 ;
        RECT 104.780 154.430 105.100 154.490 ;
        RECT 108.935 154.630 109.225 154.675 ;
        RECT 110.300 154.630 110.620 154.690 ;
        RECT 108.935 154.490 110.620 154.630 ;
        RECT 108.935 154.445 109.225 154.490 ;
        RECT 110.300 154.430 110.620 154.490 ;
        RECT 92.375 154.290 92.665 154.335 ;
        RECT 104.335 154.290 104.625 154.335 ;
        RECT 91.530 154.150 104.625 154.290 ;
        RECT 91.530 153.270 91.670 154.150 ;
        RECT 92.375 154.105 92.665 154.150 ;
        RECT 104.335 154.105 104.625 154.150 ;
        RECT 94.660 153.950 94.980 154.010 ;
        RECT 97.435 153.950 97.725 153.995 ;
        RECT 94.660 153.810 97.725 153.950 ;
        RECT 94.660 153.750 94.980 153.810 ;
        RECT 97.435 153.765 97.725 153.810 ;
        RECT 97.895 153.765 98.185 153.995 ;
        RECT 91.915 153.610 92.205 153.655 ;
        RECT 95.595 153.610 95.885 153.655 ;
        RECT 91.915 153.470 95.885 153.610 ;
        RECT 97.970 153.610 98.110 153.765 ;
        RECT 98.340 153.750 98.660 154.010 ;
        RECT 99.260 153.750 99.580 154.010 ;
        RECT 108.015 153.950 108.305 153.995 ;
        RECT 106.250 153.810 108.305 153.950 ;
        RECT 98.800 153.610 99.120 153.670 ;
        RECT 97.970 153.470 99.120 153.610 ;
        RECT 91.915 153.425 92.205 153.470 ;
        RECT 95.595 153.425 95.885 153.470 ;
        RECT 92.360 153.270 92.680 153.330 ;
        RECT 91.530 153.130 92.680 153.270 ;
        RECT 95.670 153.270 95.810 153.425 ;
        RECT 98.800 153.410 99.120 153.470 ;
        RECT 103.415 153.425 103.705 153.655 ;
        RECT 97.420 153.270 97.740 153.330 ;
        RECT 95.670 153.130 97.740 153.270 ;
        RECT 103.490 153.270 103.630 153.425 ;
        RECT 103.860 153.410 104.180 153.670 ;
        RECT 104.320 153.270 104.640 153.330 ;
        RECT 106.250 153.315 106.390 153.810 ;
        RECT 108.015 153.765 108.305 153.810 ;
        RECT 103.490 153.130 104.640 153.270 ;
        RECT 92.360 153.070 92.680 153.130 ;
        RECT 97.420 153.070 97.740 153.130 ;
        RECT 104.320 153.070 104.640 153.130 ;
        RECT 106.175 153.085 106.465 153.315 ;
        RECT 37.620 152.790 40.610 152.930 ;
        RECT 41.775 152.930 42.065 152.975 ;
        RECT 42.220 152.930 42.540 152.990 ;
        RECT 41.775 152.790 42.540 152.930 ;
        RECT 32.100 152.730 32.420 152.790 ;
        RECT 37.620 152.730 37.940 152.790 ;
        RECT 41.775 152.745 42.065 152.790 ;
        RECT 42.220 152.730 42.540 152.790 ;
        RECT 44.980 152.930 45.300 152.990 ;
        RECT 49.135 152.930 49.425 152.975 ;
        RECT 44.980 152.790 49.425 152.930 ;
        RECT 44.980 152.730 45.300 152.790 ;
        RECT 49.135 152.745 49.425 152.790 ;
        RECT 57.400 152.730 57.720 152.990 ;
        RECT 58.320 152.930 58.640 152.990 ;
        RECT 65.680 152.930 66.000 152.990 ;
        RECT 66.155 152.930 66.445 152.975 ;
        RECT 58.320 152.790 66.445 152.930 ;
        RECT 58.320 152.730 58.640 152.790 ;
        RECT 65.680 152.730 66.000 152.790 ;
        RECT 66.155 152.745 66.445 152.790 ;
        RECT 68.900 152.930 69.220 152.990 ;
        RECT 70.295 152.930 70.585 152.975 ;
        RECT 68.900 152.790 70.585 152.930 ;
        RECT 68.900 152.730 69.220 152.790 ;
        RECT 70.295 152.745 70.585 152.790 ;
        RECT 79.035 152.930 79.325 152.975 ;
        RECT 79.480 152.930 79.800 152.990 ;
        RECT 79.035 152.790 79.800 152.930 ;
        RECT 79.035 152.745 79.325 152.790 ;
        RECT 79.480 152.730 79.800 152.790 ;
        RECT 81.795 152.930 82.085 152.975 ;
        RECT 82.700 152.930 83.020 152.990 ;
        RECT 81.795 152.790 83.020 152.930 ;
        RECT 81.795 152.745 82.085 152.790 ;
        RECT 82.700 152.730 83.020 152.790 ;
        RECT 90.980 152.730 91.300 152.990 ;
        RECT 96.040 152.730 96.360 152.990 ;
        RECT 15.010 152.110 113.450 152.590 ;
        RECT 17.625 151.910 17.915 151.955 ;
        RECT 20.600 151.910 20.920 151.970 ;
        RECT 17.625 151.770 20.920 151.910 ;
        RECT 17.625 151.725 17.915 151.770 ;
        RECT 20.600 151.710 20.920 151.770 ;
        RECT 29.340 151.710 29.660 151.970 ;
        RECT 33.020 151.910 33.340 151.970 ;
        RECT 39.920 151.910 40.240 151.970 ;
        RECT 33.020 151.770 40.240 151.910 ;
        RECT 33.020 151.710 33.340 151.770 ;
        RECT 21.490 151.570 21.780 151.615 ;
        RECT 24.270 151.570 24.560 151.615 ;
        RECT 26.130 151.570 26.420 151.615 ;
        RECT 21.490 151.430 26.420 151.570 ;
        RECT 21.490 151.385 21.780 151.430 ;
        RECT 24.270 151.385 24.560 151.430 ;
        RECT 26.130 151.385 26.420 151.430 ;
        RECT 27.960 151.570 28.280 151.630 ;
        RECT 27.960 151.430 30.950 151.570 ;
        RECT 27.960 151.370 28.280 151.430 ;
        RECT 26.580 151.030 26.900 151.290 ;
        RECT 28.880 151.030 29.200 151.290 ;
        RECT 30.810 151.275 30.950 151.430 ;
        RECT 33.955 151.385 34.245 151.615 ;
        RECT 30.735 151.045 31.025 151.275 ;
        RECT 21.490 150.890 21.780 150.935 ;
        RECT 21.490 150.750 24.025 150.890 ;
        RECT 21.490 150.705 21.780 150.750 ;
        RECT 19.630 150.550 19.920 150.595 ;
        RECT 21.980 150.550 22.300 150.610 ;
        RECT 23.810 150.595 24.025 150.750 ;
        RECT 24.740 150.690 25.060 150.950 ;
        RECT 28.420 150.690 28.740 150.950 ;
        RECT 29.800 150.690 30.120 150.950 ;
        RECT 32.100 150.690 32.420 150.950 ;
        RECT 34.030 150.890 34.170 151.385 ;
        RECT 35.335 150.890 35.625 150.935 ;
        RECT 34.030 150.750 35.625 150.890 ;
        RECT 35.335 150.705 35.625 150.750 ;
        RECT 37.620 150.690 37.940 150.950 ;
        RECT 38.170 150.935 38.310 151.770 ;
        RECT 39.920 151.710 40.240 151.770 ;
        RECT 58.780 151.910 59.100 151.970 ;
        RECT 67.060 151.910 67.380 151.970 ;
        RECT 58.780 151.770 67.380 151.910 ;
        RECT 58.780 151.710 59.100 151.770 ;
        RECT 50.960 151.570 51.280 151.630 ;
        RECT 62.460 151.570 62.780 151.630 ;
        RECT 42.770 151.430 62.780 151.570 ;
        RECT 39.920 151.230 40.240 151.290 ;
        RECT 42.770 151.230 42.910 151.430 ;
        RECT 50.960 151.370 51.280 151.430 ;
        RECT 62.460 151.370 62.780 151.430 ;
        RECT 44.980 151.230 45.300 151.290 ;
        RECT 39.920 151.090 42.910 151.230 ;
        RECT 39.920 151.030 40.240 151.090 ;
        RECT 38.095 150.705 38.385 150.935 ;
        RECT 38.555 150.705 38.845 150.935 ;
        RECT 39.000 150.890 39.320 150.950 ;
        RECT 42.770 150.935 42.910 151.090 ;
        RECT 43.230 151.090 45.300 151.230 ;
        RECT 43.230 150.935 43.370 151.090 ;
        RECT 44.980 151.030 45.300 151.090 ;
        RECT 45.440 151.230 45.760 151.290 ;
        RECT 49.135 151.230 49.425 151.275 ;
        RECT 58.320 151.230 58.640 151.290 ;
        RECT 45.440 151.090 58.640 151.230 ;
        RECT 45.440 151.030 45.760 151.090 ;
        RECT 49.135 151.045 49.425 151.090 ;
        RECT 58.320 151.030 58.640 151.090 ;
        RECT 39.475 150.890 39.765 150.935 ;
        RECT 39.000 150.750 39.765 150.890 ;
        RECT 22.890 150.550 23.180 150.595 ;
        RECT 19.630 150.410 23.180 150.550 ;
        RECT 19.630 150.365 19.920 150.410 ;
        RECT 21.980 150.350 22.300 150.410 ;
        RECT 22.890 150.365 23.180 150.410 ;
        RECT 23.810 150.550 24.100 150.595 ;
        RECT 25.670 150.550 25.960 150.595 ;
        RECT 23.810 150.410 25.960 150.550 ;
        RECT 23.810 150.365 24.100 150.410 ;
        RECT 25.670 150.365 25.960 150.410 ;
        RECT 26.120 150.550 26.440 150.610 ;
        RECT 31.655 150.550 31.945 150.595 ;
        RECT 38.630 150.550 38.770 150.705 ;
        RECT 39.000 150.690 39.320 150.750 ;
        RECT 39.475 150.705 39.765 150.750 ;
        RECT 42.235 150.705 42.525 150.935 ;
        RECT 42.695 150.705 42.985 150.935 ;
        RECT 43.155 150.705 43.445 150.935 ;
        RECT 44.075 150.890 44.365 150.935 ;
        RECT 44.520 150.890 44.840 150.950 ;
        RECT 44.075 150.750 44.840 150.890 ;
        RECT 44.075 150.705 44.365 150.750 ;
        RECT 42.310 150.550 42.450 150.705 ;
        RECT 44.520 150.690 44.840 150.750 ;
        RECT 50.055 150.890 50.345 150.935 ;
        RECT 56.020 150.890 56.340 150.950 ;
        RECT 50.055 150.750 56.340 150.890 ;
        RECT 50.055 150.705 50.345 150.750 ;
        RECT 56.020 150.690 56.340 150.750 ;
        RECT 60.620 150.890 60.940 150.950 ;
        RECT 63.380 150.890 63.700 150.950 ;
        RECT 60.620 150.750 63.700 150.890 ;
        RECT 60.620 150.690 60.940 150.750 ;
        RECT 63.380 150.690 63.700 150.750 ;
        RECT 63.840 150.690 64.160 150.950 ;
        RECT 65.310 150.935 65.450 151.770 ;
        RECT 67.060 151.710 67.380 151.770 ;
        RECT 71.215 151.910 71.505 151.955 ;
        RECT 73.960 151.910 74.280 151.970 ;
        RECT 71.215 151.770 74.280 151.910 ;
        RECT 71.215 151.725 71.505 151.770 ;
        RECT 73.960 151.710 74.280 151.770 ;
        RECT 86.395 151.910 86.685 151.955 ;
        RECT 86.840 151.910 87.160 151.970 ;
        RECT 86.395 151.770 87.160 151.910 ;
        RECT 86.395 151.725 86.685 151.770 ;
        RECT 86.840 151.710 87.160 151.770 ;
        RECT 87.760 151.910 88.080 151.970 ;
        RECT 90.980 151.910 91.300 151.970 ;
        RECT 87.760 151.770 91.300 151.910 ;
        RECT 87.760 151.710 88.080 151.770 ;
        RECT 90.980 151.710 91.300 151.770 ;
        RECT 91.915 151.910 92.205 151.955 ;
        RECT 94.200 151.910 94.520 151.970 ;
        RECT 91.915 151.770 94.520 151.910 ;
        RECT 91.915 151.725 92.205 151.770 ;
        RECT 94.200 151.710 94.520 151.770 ;
        RECT 94.660 151.710 94.980 151.970 ;
        RECT 66.615 151.570 66.905 151.615 ;
        RECT 76.260 151.570 76.580 151.630 ;
        RECT 66.615 151.430 76.580 151.570 ;
        RECT 66.615 151.385 66.905 151.430 ;
        RECT 76.260 151.370 76.580 151.430 ;
        RECT 79.450 151.570 79.740 151.615 ;
        RECT 82.230 151.570 82.520 151.615 ;
        RECT 84.090 151.570 84.380 151.615 ;
        RECT 79.450 151.430 84.380 151.570 ;
        RECT 79.450 151.385 79.740 151.430 ;
        RECT 82.230 151.385 82.520 151.430 ;
        RECT 84.090 151.385 84.380 151.430 ;
        RECT 84.540 151.570 84.860 151.630 ;
        RECT 88.235 151.570 88.525 151.615 ;
        RECT 84.540 151.430 88.525 151.570 ;
        RECT 84.540 151.370 84.860 151.430 ;
        RECT 88.235 151.385 88.525 151.430 ;
        RECT 92.375 151.570 92.665 151.615 ;
        RECT 105.700 151.570 106.020 151.630 ;
        RECT 92.375 151.430 106.020 151.570 ;
        RECT 92.375 151.385 92.665 151.430 ;
        RECT 105.700 151.370 106.020 151.430 ;
        RECT 107.095 151.385 107.385 151.615 ;
        RECT 70.740 151.030 71.060 151.290 ;
        RECT 75.800 151.230 76.120 151.290 ;
        RECT 71.290 151.090 76.120 151.230 ;
        RECT 64.315 150.705 64.605 150.935 ;
        RECT 65.235 150.705 65.525 150.935 ;
        RECT 26.120 150.410 38.770 150.550 ;
        RECT 39.090 150.410 42.450 150.550 ;
        RECT 26.120 150.350 26.440 150.410 ;
        RECT 31.655 150.365 31.945 150.410 ;
        RECT 39.090 150.270 39.230 150.410 ;
        RECT 52.340 150.350 52.660 150.610 ;
        RECT 61.080 150.350 61.400 150.610 ;
        RECT 61.540 150.550 61.860 150.610 ;
        RECT 64.390 150.550 64.530 150.705 ;
        RECT 67.980 150.690 68.300 150.950 ;
        RECT 69.820 150.690 70.140 150.950 ;
        RECT 71.290 150.890 71.430 151.090 ;
        RECT 73.590 150.950 73.730 151.090 ;
        RECT 75.800 151.030 76.120 151.090 ;
        RECT 82.700 151.030 83.020 151.290 ;
        RECT 89.600 151.230 89.920 151.290 ;
        RECT 90.995 151.230 91.285 151.275 ;
        RECT 89.600 151.090 91.285 151.230 ;
        RECT 89.600 151.030 89.920 151.090 ;
        RECT 90.995 151.045 91.285 151.090 ;
        RECT 94.215 151.230 94.505 151.275 ;
        RECT 95.120 151.230 95.440 151.290 ;
        RECT 94.215 151.090 95.440 151.230 ;
        RECT 94.215 151.045 94.505 151.090 ;
        RECT 95.120 151.030 95.440 151.090 ;
        RECT 96.590 151.090 100.410 151.230 ;
        RECT 70.600 150.750 71.430 150.890 ;
        RECT 70.600 150.550 70.740 150.750 ;
        RECT 73.040 150.690 73.360 150.950 ;
        RECT 73.500 150.690 73.820 150.950 ;
        RECT 73.975 150.705 74.265 150.935 ;
        RECT 74.895 150.890 75.185 150.935 ;
        RECT 75.340 150.890 75.660 150.950 ;
        RECT 74.895 150.750 75.660 150.890 ;
        RECT 74.895 150.705 75.185 150.750 ;
        RECT 61.540 150.410 64.530 150.550 ;
        RECT 68.530 150.410 70.740 150.550 ;
        RECT 71.215 150.550 71.505 150.595 ;
        RECT 71.675 150.550 71.965 150.595 ;
        RECT 71.215 150.410 71.965 150.550 ;
        RECT 61.540 150.350 61.860 150.410 ;
        RECT 24.280 150.210 24.600 150.270 ;
        RECT 27.515 150.210 27.805 150.255 ;
        RECT 24.280 150.070 27.805 150.210 ;
        RECT 24.280 150.010 24.600 150.070 ;
        RECT 27.515 150.025 27.805 150.070 ;
        RECT 34.415 150.210 34.705 150.255 ;
        RECT 34.860 150.210 35.180 150.270 ;
        RECT 34.415 150.070 35.180 150.210 ;
        RECT 34.415 150.025 34.705 150.070 ;
        RECT 34.860 150.010 35.180 150.070 ;
        RECT 35.320 150.210 35.640 150.270 ;
        RECT 36.255 150.210 36.545 150.255 ;
        RECT 35.320 150.070 36.545 150.210 ;
        RECT 35.320 150.010 35.640 150.070 ;
        RECT 36.255 150.025 36.545 150.070 ;
        RECT 39.000 150.010 39.320 150.270 ;
        RECT 40.840 150.010 41.160 150.270 ;
        RECT 47.740 150.210 48.060 150.270 ;
        RECT 49.595 150.210 49.885 150.255 ;
        RECT 47.740 150.070 49.885 150.210 ;
        RECT 47.740 150.010 48.060 150.070 ;
        RECT 49.595 150.025 49.885 150.070 ;
        RECT 51.880 150.010 52.200 150.270 ;
        RECT 57.400 150.210 57.720 150.270 ;
        RECT 59.240 150.210 59.560 150.270 ;
        RECT 57.400 150.070 59.560 150.210 ;
        RECT 57.400 150.010 57.720 150.070 ;
        RECT 59.240 150.010 59.560 150.070 ;
        RECT 62.000 150.010 62.320 150.270 ;
        RECT 62.460 150.210 62.780 150.270 ;
        RECT 68.530 150.210 68.670 150.410 ;
        RECT 71.215 150.365 71.505 150.410 ;
        RECT 71.675 150.365 71.965 150.410 ;
        RECT 62.460 150.070 68.670 150.210 ;
        RECT 62.460 150.010 62.780 150.070 ;
        RECT 68.900 150.010 69.220 150.270 ;
        RECT 74.050 150.210 74.190 150.705 ;
        RECT 75.340 150.690 75.660 150.750 ;
        RECT 79.450 150.890 79.740 150.935 ;
        RECT 79.450 150.750 81.985 150.890 ;
        RECT 79.450 150.705 79.740 150.750 ;
        RECT 77.590 150.550 77.880 150.595 ;
        RECT 79.940 150.550 80.260 150.610 ;
        RECT 81.770 150.595 81.985 150.750 ;
        RECT 84.540 150.690 84.860 150.950 ;
        RECT 85.935 150.705 86.225 150.935 ;
        RECT 80.850 150.550 81.140 150.595 ;
        RECT 77.590 150.410 81.140 150.550 ;
        RECT 77.590 150.365 77.880 150.410 ;
        RECT 79.940 150.350 80.260 150.410 ;
        RECT 80.850 150.365 81.140 150.410 ;
        RECT 81.770 150.550 82.060 150.595 ;
        RECT 83.630 150.550 83.920 150.595 ;
        RECT 81.770 150.410 83.920 150.550 ;
        RECT 81.770 150.365 82.060 150.410 ;
        RECT 83.630 150.365 83.920 150.410 ;
        RECT 75.585 150.210 75.875 150.255 ;
        RECT 78.100 150.210 78.420 150.270 ;
        RECT 74.050 150.070 78.420 150.210 ;
        RECT 75.585 150.025 75.875 150.070 ;
        RECT 78.100 150.010 78.420 150.070 ;
        RECT 83.160 150.210 83.480 150.270 ;
        RECT 86.010 150.210 86.150 150.705 ;
        RECT 89.140 150.690 89.460 150.950 ;
        RECT 90.520 150.690 90.840 150.950 ;
        RECT 91.440 150.890 91.760 150.950 ;
        RECT 92.360 150.890 92.680 150.950 ;
        RECT 91.440 150.750 92.680 150.890 ;
        RECT 91.440 150.690 91.760 150.750 ;
        RECT 92.360 150.690 92.680 150.750 ;
        RECT 92.820 150.890 93.140 150.950 ;
        RECT 96.590 150.935 96.730 151.090 ;
        RECT 100.270 150.950 100.410 151.090 ;
        RECT 104.320 151.030 104.640 151.290 ;
        RECT 93.295 150.890 93.585 150.935 ;
        RECT 92.820 150.750 93.585 150.890 ;
        RECT 92.820 150.690 93.140 150.750 ;
        RECT 93.295 150.705 93.585 150.750 ;
        RECT 96.515 150.705 96.805 150.935 ;
        RECT 96.960 150.690 97.280 150.950 ;
        RECT 97.420 150.690 97.740 150.950 ;
        RECT 98.355 150.890 98.645 150.935 ;
        RECT 99.720 150.890 100.040 150.950 ;
        RECT 98.355 150.750 100.040 150.890 ;
        RECT 98.355 150.705 98.645 150.750 ;
        RECT 99.720 150.690 100.040 150.750 ;
        RECT 100.180 150.690 100.500 150.950 ;
        RECT 100.655 150.705 100.945 150.935 ;
        RECT 91.915 150.365 92.205 150.595 ;
        RECT 94.675 150.550 94.965 150.595 ;
        RECT 95.135 150.550 95.425 150.595 ;
        RECT 94.675 150.410 95.425 150.550 ;
        RECT 97.050 150.550 97.190 150.690 ;
        RECT 100.730 150.550 100.870 150.705 ;
        RECT 101.100 150.690 101.420 150.950 ;
        RECT 102.035 150.890 102.325 150.935 ;
        RECT 101.650 150.750 102.325 150.890 ;
        RECT 97.050 150.410 100.870 150.550 ;
        RECT 94.675 150.365 94.965 150.410 ;
        RECT 95.135 150.365 95.425 150.410 ;
        RECT 83.160 150.070 86.150 150.210 ;
        RECT 89.615 150.210 89.905 150.255 ;
        RECT 90.520 150.210 90.840 150.270 ;
        RECT 89.615 150.070 90.840 150.210 ;
        RECT 91.990 150.210 92.130 150.365 ;
        RECT 98.815 150.210 99.105 150.255 ;
        RECT 91.990 150.070 99.105 150.210 ;
        RECT 83.160 150.010 83.480 150.070 ;
        RECT 89.615 150.025 89.905 150.070 ;
        RECT 90.520 150.010 90.840 150.070 ;
        RECT 98.815 150.025 99.105 150.070 ;
        RECT 99.720 150.210 100.040 150.270 ;
        RECT 101.650 150.210 101.790 150.750 ;
        RECT 102.035 150.705 102.325 150.750 ;
        RECT 103.860 150.890 104.180 150.950 ;
        RECT 105.255 150.890 105.545 150.935 ;
        RECT 103.860 150.750 105.545 150.890 ;
        RECT 107.170 150.890 107.310 151.385 ;
        RECT 108.475 150.890 108.765 150.935 ;
        RECT 107.170 150.750 108.765 150.890 ;
        RECT 103.860 150.690 104.180 150.750 ;
        RECT 105.255 150.705 105.545 150.750 ;
        RECT 108.475 150.705 108.765 150.750 ;
        RECT 99.720 150.070 101.790 150.210 ;
        RECT 99.720 150.010 100.040 150.070 ;
        RECT 104.780 150.010 105.100 150.270 ;
        RECT 109.380 150.010 109.700 150.270 ;
        RECT 15.010 149.390 113.450 149.870 ;
        RECT 18.775 149.190 19.065 149.235 ;
        RECT 20.140 149.190 20.460 149.250 ;
        RECT 18.775 149.050 20.460 149.190 ;
        RECT 18.775 149.005 19.065 149.050 ;
        RECT 20.140 148.990 20.460 149.050 ;
        RECT 21.535 149.190 21.825 149.235 ;
        RECT 21.980 149.190 22.300 149.250 ;
        RECT 21.535 149.050 22.300 149.190 ;
        RECT 21.535 149.005 21.825 149.050 ;
        RECT 21.980 148.990 22.300 149.050 ;
        RECT 24.740 148.990 25.060 149.250 ;
        RECT 25.445 149.190 25.735 149.235 ;
        RECT 26.120 149.190 26.440 149.250 ;
        RECT 25.445 149.050 26.440 149.190 ;
        RECT 25.445 149.005 25.735 149.050 ;
        RECT 26.120 148.990 26.440 149.050 ;
        RECT 39.015 149.190 39.305 149.235 ;
        RECT 39.015 149.050 42.910 149.190 ;
        RECT 39.015 149.005 39.305 149.050 ;
        RECT 16.920 148.850 17.240 148.910 ;
        RECT 27.450 148.850 27.740 148.895 ;
        RECT 28.880 148.850 29.200 148.910 ;
        RECT 30.710 148.850 31.000 148.895 ;
        RECT 16.920 148.710 22.210 148.850 ;
        RECT 16.920 148.650 17.240 148.710 ;
        RECT 18.390 148.555 18.530 148.710 ;
        RECT 22.070 148.570 22.210 148.710 ;
        RECT 27.450 148.710 31.000 148.850 ;
        RECT 27.450 148.665 27.740 148.710 ;
        RECT 28.880 148.650 29.200 148.710 ;
        RECT 30.710 148.665 31.000 148.710 ;
        RECT 31.630 148.850 31.920 148.895 ;
        RECT 33.490 148.850 33.780 148.895 ;
        RECT 31.630 148.710 33.780 148.850 ;
        RECT 31.630 148.665 31.920 148.710 ;
        RECT 33.490 148.665 33.780 148.710 ;
        RECT 35.780 148.850 36.100 148.910 ;
        RECT 35.780 148.710 37.850 148.850 ;
        RECT 18.315 148.325 18.605 148.555 ;
        RECT 19.680 148.310 20.000 148.570 ;
        RECT 21.980 148.310 22.300 148.570 ;
        RECT 23.820 148.310 24.140 148.570 ;
        RECT 29.310 148.510 29.600 148.555 ;
        RECT 31.630 148.510 31.845 148.665 ;
        RECT 35.780 148.650 36.100 148.710 ;
        RECT 29.310 148.370 31.845 148.510 ;
        RECT 32.575 148.510 32.865 148.555 ;
        RECT 34.860 148.510 35.180 148.570 ;
        RECT 32.575 148.370 35.180 148.510 ;
        RECT 29.310 148.325 29.600 148.370 ;
        RECT 32.575 148.325 32.865 148.370 ;
        RECT 34.860 148.310 35.180 148.370 ;
        RECT 37.175 148.325 37.465 148.555 ;
        RECT 37.710 148.510 37.850 148.710 ;
        RECT 38.540 148.650 38.860 148.910 ;
        RECT 40.840 148.850 41.160 148.910 ;
        RECT 41.315 148.850 41.605 148.895 ;
        RECT 40.840 148.710 41.605 148.850 ;
        RECT 40.840 148.650 41.160 148.710 ;
        RECT 41.315 148.665 41.605 148.710 ;
        RECT 39.935 148.510 40.225 148.555 ;
        RECT 37.710 148.370 40.225 148.510 ;
        RECT 39.935 148.325 40.225 148.370 ;
        RECT 34.415 148.170 34.705 148.215 ;
        RECT 35.780 148.170 36.100 148.230 ;
        RECT 34.415 148.030 36.100 148.170 ;
        RECT 34.415 147.985 34.705 148.030 ;
        RECT 35.780 147.970 36.100 148.030 ;
        RECT 20.615 147.830 20.905 147.875 ;
        RECT 23.360 147.830 23.680 147.890 ;
        RECT 20.615 147.690 23.680 147.830 ;
        RECT 20.615 147.645 20.905 147.690 ;
        RECT 23.360 147.630 23.680 147.690 ;
        RECT 29.310 147.830 29.600 147.875 ;
        RECT 32.090 147.830 32.380 147.875 ;
        RECT 33.950 147.830 34.240 147.875 ;
        RECT 36.255 147.830 36.545 147.875 ;
        RECT 29.310 147.690 34.240 147.830 ;
        RECT 29.310 147.645 29.600 147.690 ;
        RECT 32.090 147.645 32.380 147.690 ;
        RECT 33.950 147.645 34.240 147.690 ;
        RECT 34.490 147.690 36.545 147.830 ;
        RECT 37.250 147.830 37.390 148.325 ;
        RECT 40.380 148.310 40.700 148.570 ;
        RECT 41.760 148.310 42.080 148.570 ;
        RECT 38.080 147.970 38.400 148.230 ;
        RECT 41.300 148.170 41.620 148.230 ;
        RECT 42.235 148.170 42.525 148.215 ;
        RECT 41.300 148.030 42.525 148.170 ;
        RECT 42.770 148.170 42.910 149.050 ;
        RECT 44.075 149.005 44.365 149.235 ;
        RECT 46.375 149.190 46.665 149.235 ;
        RECT 47.740 149.190 48.060 149.250 ;
        RECT 46.375 149.050 48.060 149.190 ;
        RECT 46.375 149.005 46.665 149.050 ;
        RECT 44.150 148.850 44.290 149.005 ;
        RECT 47.740 148.990 48.060 149.050 ;
        RECT 56.480 149.190 56.800 149.250 ;
        RECT 58.780 149.235 59.100 149.250 ;
        RECT 56.955 149.190 57.245 149.235 ;
        RECT 56.480 149.050 57.245 149.190 ;
        RECT 56.480 148.990 56.800 149.050 ;
        RECT 56.955 149.005 57.245 149.050 ;
        RECT 58.780 149.190 59.315 149.235 ;
        RECT 61.540 149.190 61.860 149.250 ;
        RECT 73.500 149.190 73.820 149.250 ;
        RECT 58.780 149.050 61.860 149.190 ;
        RECT 58.780 149.005 59.315 149.050 ;
        RECT 58.780 148.990 59.100 149.005 ;
        RECT 61.540 148.990 61.860 149.050 ;
        RECT 72.670 149.050 73.820 149.190 ;
        RECT 59.700 148.850 60.020 148.910 ;
        RECT 44.150 148.710 60.020 148.850 ;
        RECT 59.700 148.650 60.020 148.710 ;
        RECT 61.030 148.850 61.320 148.895 ;
        RECT 62.460 148.850 62.780 148.910 ;
        RECT 64.290 148.850 64.580 148.895 ;
        RECT 61.030 148.710 64.580 148.850 ;
        RECT 61.030 148.665 61.320 148.710 ;
        RECT 62.460 148.650 62.780 148.710 ;
        RECT 64.290 148.665 64.580 148.710 ;
        RECT 65.210 148.850 65.500 148.895 ;
        RECT 67.070 148.850 67.360 148.895 ;
        RECT 65.210 148.710 67.360 148.850 ;
        RECT 65.210 148.665 65.500 148.710 ;
        RECT 67.070 148.665 67.360 148.710 ;
        RECT 43.155 148.510 43.445 148.555 ;
        RECT 43.600 148.510 43.920 148.570 ;
        RECT 51.880 148.510 52.200 148.570 ;
        RECT 56.035 148.510 56.325 148.555 ;
        RECT 43.155 148.370 43.920 148.510 ;
        RECT 43.155 148.325 43.445 148.370 ;
        RECT 43.600 148.310 43.920 148.370 ;
        RECT 45.070 148.370 47.970 148.510 ;
        RECT 45.070 148.170 45.210 148.370 ;
        RECT 42.770 148.030 45.210 148.170 ;
        RECT 41.300 147.970 41.620 148.030 ;
        RECT 42.235 147.985 42.525 148.030 ;
        RECT 45.440 147.970 45.760 148.230 ;
        RECT 45.900 147.970 46.220 148.230 ;
        RECT 47.830 148.170 47.970 148.370 ;
        RECT 51.880 148.370 56.325 148.510 ;
        RECT 51.880 148.310 52.200 148.370 ;
        RECT 56.035 148.325 56.325 148.370 ;
        RECT 62.890 148.510 63.180 148.555 ;
        RECT 65.210 148.510 65.425 148.665 ;
        RECT 62.890 148.370 65.425 148.510 ;
        RECT 68.455 148.510 68.745 148.555 ;
        RECT 70.280 148.510 70.600 148.570 ;
        RECT 72.670 148.555 72.810 149.050 ;
        RECT 73.500 148.990 73.820 149.050 ;
        RECT 74.880 149.190 75.200 149.250 ;
        RECT 77.195 149.190 77.485 149.235 ;
        RECT 74.880 149.050 77.485 149.190 ;
        RECT 74.880 148.990 75.200 149.050 ;
        RECT 77.195 149.005 77.485 149.050 ;
        RECT 79.495 149.190 79.785 149.235 ;
        RECT 80.400 149.190 80.720 149.250 ;
        RECT 79.495 149.050 80.720 149.190 ;
        RECT 79.495 149.005 79.785 149.050 ;
        RECT 80.400 148.990 80.720 149.050 ;
        RECT 87.315 149.190 87.605 149.235 ;
        RECT 89.140 149.190 89.460 149.250 ;
        RECT 87.315 149.050 89.460 149.190 ;
        RECT 87.315 149.005 87.605 149.050 ;
        RECT 89.140 148.990 89.460 149.050 ;
        RECT 93.755 149.190 94.045 149.235 ;
        RECT 99.260 149.190 99.580 149.250 ;
        RECT 93.755 149.050 99.580 149.190 ;
        RECT 93.755 149.005 94.045 149.050 ;
        RECT 99.260 148.990 99.580 149.050 ;
        RECT 74.420 148.850 74.740 148.910 ;
        RECT 78.100 148.850 78.420 148.910 ;
        RECT 81.795 148.850 82.085 148.895 ;
        RECT 85.475 148.850 85.765 148.895 ;
        RECT 73.130 148.710 76.950 148.850 ;
        RECT 73.130 148.555 73.270 148.710 ;
        RECT 74.420 148.650 74.740 148.710 ;
        RECT 72.135 148.510 72.425 148.555 ;
        RECT 68.455 148.370 70.600 148.510 ;
        RECT 62.890 148.325 63.180 148.370 ;
        RECT 68.455 148.325 68.745 148.370 ;
        RECT 70.280 148.310 70.600 148.370 ;
        RECT 71.750 148.370 72.425 148.510 ;
        RECT 60.160 148.170 60.480 148.230 ;
        RECT 47.830 148.030 60.480 148.170 ;
        RECT 60.160 147.970 60.480 148.030 ;
        RECT 66.155 148.170 66.445 148.215 ;
        RECT 67.060 148.170 67.380 148.230 ;
        RECT 66.155 148.030 67.380 148.170 ;
        RECT 66.155 147.985 66.445 148.030 ;
        RECT 67.060 147.970 67.380 148.030 ;
        RECT 67.980 147.970 68.300 148.230 ;
        RECT 62.000 147.830 62.320 147.890 ;
        RECT 37.250 147.690 62.320 147.830 ;
        RECT 27.500 147.490 27.820 147.550 ;
        RECT 34.490 147.490 34.630 147.690 ;
        RECT 36.255 147.645 36.545 147.690 ;
        RECT 62.000 147.630 62.320 147.690 ;
        RECT 62.890 147.830 63.180 147.875 ;
        RECT 65.670 147.830 65.960 147.875 ;
        RECT 67.530 147.830 67.820 147.875 ;
        RECT 62.890 147.690 67.820 147.830 ;
        RECT 62.890 147.645 63.180 147.690 ;
        RECT 65.670 147.645 65.960 147.690 ;
        RECT 67.530 147.645 67.820 147.690 ;
        RECT 69.375 147.830 69.665 147.875 ;
        RECT 71.750 147.830 71.890 148.370 ;
        RECT 72.135 148.325 72.425 148.370 ;
        RECT 72.595 148.325 72.885 148.555 ;
        RECT 73.055 148.325 73.345 148.555 ;
        RECT 73.500 148.510 73.820 148.570 ;
        RECT 73.975 148.510 74.265 148.555 ;
        RECT 75.340 148.510 75.660 148.570 ;
        RECT 76.810 148.555 76.950 148.710 ;
        RECT 78.100 148.710 85.765 148.850 ;
        RECT 78.100 148.650 78.420 148.710 ;
        RECT 81.795 148.665 82.085 148.710 ;
        RECT 85.475 148.665 85.765 148.710 ;
        RECT 95.580 148.650 95.900 148.910 ;
        RECT 96.055 148.850 96.345 148.895 ;
        RECT 96.515 148.850 96.805 148.895 ;
        RECT 100.180 148.850 100.500 148.910 ;
        RECT 96.055 148.710 96.805 148.850 ;
        RECT 96.055 148.665 96.345 148.710 ;
        RECT 96.515 148.665 96.805 148.710 ;
        RECT 97.970 148.710 100.500 148.850 ;
        RECT 73.500 148.370 75.660 148.510 ;
        RECT 73.500 148.310 73.820 148.370 ;
        RECT 73.975 148.325 74.265 148.370 ;
        RECT 75.340 148.310 75.660 148.370 ;
        RECT 76.735 148.510 77.025 148.555 ;
        RECT 81.335 148.510 81.625 148.555 ;
        RECT 76.735 148.370 81.625 148.510 ;
        RECT 76.735 148.325 77.025 148.370 ;
        RECT 81.335 148.325 81.625 148.370 ;
        RECT 85.015 148.510 85.305 148.555 ;
        RECT 91.440 148.510 91.760 148.570 ;
        RECT 85.015 148.370 91.760 148.510 ;
        RECT 85.015 148.325 85.305 148.370 ;
        RECT 91.440 148.310 91.760 148.370 ;
        RECT 94.675 148.510 94.965 148.555 ;
        RECT 95.670 148.510 95.810 148.650 ;
        RECT 94.675 148.370 95.810 148.510 ;
        RECT 96.960 148.510 97.280 148.570 ;
        RECT 97.970 148.555 98.110 148.710 ;
        RECT 100.180 148.650 100.500 148.710 ;
        RECT 101.575 148.850 101.865 148.895 ;
        RECT 104.730 148.850 105.020 148.895 ;
        RECT 107.990 148.850 108.280 148.895 ;
        RECT 101.575 148.710 108.280 148.850 ;
        RECT 101.575 148.665 101.865 148.710 ;
        RECT 104.730 148.665 105.020 148.710 ;
        RECT 107.990 148.665 108.280 148.710 ;
        RECT 108.910 148.850 109.200 148.895 ;
        RECT 110.770 148.850 111.060 148.895 ;
        RECT 108.910 148.710 111.060 148.850 ;
        RECT 108.910 148.665 109.200 148.710 ;
        RECT 110.770 148.665 111.060 148.710 ;
        RECT 97.895 148.510 98.185 148.555 ;
        RECT 96.960 148.370 98.185 148.510 ;
        RECT 94.675 148.325 94.965 148.370 ;
        RECT 96.960 148.310 97.280 148.370 ;
        RECT 97.895 148.325 98.185 148.370 ;
        RECT 98.340 148.310 98.660 148.570 ;
        RECT 98.800 148.310 99.120 148.570 ;
        RECT 99.720 148.310 100.040 148.570 ;
        RECT 101.115 148.325 101.405 148.555 ;
        RECT 106.590 148.510 106.880 148.555 ;
        RECT 108.910 148.510 109.125 148.665 ;
        RECT 106.590 148.370 109.125 148.510 ;
        RECT 109.380 148.510 109.700 148.570 ;
        RECT 109.855 148.510 110.145 148.555 ;
        RECT 109.380 148.370 110.145 148.510 ;
        RECT 106.590 148.325 106.880 148.370 ;
        RECT 76.260 148.170 76.580 148.230 ;
        RECT 82.255 148.170 82.545 148.215 ;
        RECT 84.080 148.170 84.400 148.230 ;
        RECT 76.260 148.030 84.400 148.170 ;
        RECT 76.260 147.970 76.580 148.030 ;
        RECT 82.255 147.985 82.545 148.030 ;
        RECT 84.080 147.970 84.400 148.030 ;
        RECT 95.595 148.170 95.885 148.215 ;
        RECT 97.420 148.170 97.740 148.230 ;
        RECT 95.595 148.030 97.740 148.170 ;
        RECT 95.595 147.985 95.885 148.030 ;
        RECT 97.420 147.970 97.740 148.030 ;
        RECT 101.190 147.890 101.330 148.325 ;
        RECT 109.380 148.310 109.700 148.370 ;
        RECT 109.855 148.325 110.145 148.370 ;
        RECT 111.680 147.970 112.000 148.230 ;
        RECT 73.040 147.830 73.360 147.890 ;
        RECT 69.375 147.690 73.360 147.830 ;
        RECT 69.375 147.645 69.665 147.690 ;
        RECT 73.040 147.630 73.360 147.690 ;
        RECT 83.160 147.830 83.480 147.890 ;
        RECT 101.100 147.830 101.420 147.890 ;
        RECT 83.160 147.690 101.420 147.830 ;
        RECT 83.160 147.630 83.480 147.690 ;
        RECT 101.100 147.630 101.420 147.690 ;
        RECT 106.590 147.830 106.880 147.875 ;
        RECT 109.370 147.830 109.660 147.875 ;
        RECT 111.230 147.830 111.520 147.875 ;
        RECT 106.590 147.690 111.520 147.830 ;
        RECT 106.590 147.645 106.880 147.690 ;
        RECT 109.370 147.645 109.660 147.690 ;
        RECT 111.230 147.645 111.520 147.690 ;
        RECT 27.500 147.350 34.630 147.490 ;
        RECT 35.320 147.490 35.640 147.550 ;
        RECT 37.175 147.490 37.465 147.535 ;
        RECT 35.320 147.350 37.465 147.490 ;
        RECT 27.500 147.290 27.820 147.350 ;
        RECT 35.320 147.290 35.640 147.350 ;
        RECT 37.175 147.305 37.465 147.350 ;
        RECT 41.300 147.290 41.620 147.550 ;
        RECT 42.680 147.290 43.000 147.550 ;
        RECT 48.215 147.490 48.505 147.535 ;
        RECT 49.580 147.490 49.900 147.550 ;
        RECT 48.215 147.350 49.900 147.490 ;
        RECT 48.215 147.305 48.505 147.350 ;
        RECT 49.580 147.290 49.900 147.350 ;
        RECT 56.940 147.490 57.260 147.550 ;
        RECT 60.620 147.490 60.940 147.550 ;
        RECT 56.940 147.350 60.940 147.490 ;
        RECT 56.940 147.290 57.260 147.350 ;
        RECT 60.620 147.290 60.940 147.350 ;
        RECT 70.755 147.490 71.045 147.535 ;
        RECT 71.660 147.490 71.980 147.550 ;
        RECT 70.755 147.350 71.980 147.490 ;
        RECT 70.755 147.305 71.045 147.350 ;
        RECT 71.660 147.290 71.980 147.350 ;
        RECT 79.035 147.490 79.325 147.535 ;
        RECT 79.940 147.490 80.260 147.550 ;
        RECT 79.035 147.350 80.260 147.490 ;
        RECT 79.035 147.305 79.325 147.350 ;
        RECT 79.940 147.290 80.260 147.350 ;
        RECT 96.055 147.490 96.345 147.535 ;
        RECT 97.880 147.490 98.200 147.550 ;
        RECT 96.055 147.350 98.200 147.490 ;
        RECT 96.055 147.305 96.345 147.350 ;
        RECT 97.880 147.290 98.200 147.350 ;
        RECT 98.800 147.490 99.120 147.550 ;
        RECT 102.725 147.490 103.015 147.535 ;
        RECT 104.780 147.490 105.100 147.550 ;
        RECT 98.800 147.350 105.100 147.490 ;
        RECT 98.800 147.290 99.120 147.350 ;
        RECT 102.725 147.305 103.015 147.350 ;
        RECT 104.780 147.290 105.100 147.350 ;
        RECT 15.010 146.670 113.450 147.150 ;
        RECT 28.880 146.270 29.200 146.530 ;
        RECT 38.540 146.470 38.860 146.530 ;
        RECT 42.680 146.470 43.000 146.530 ;
        RECT 38.540 146.330 43.000 146.470 ;
        RECT 38.540 146.270 38.860 146.330 ;
        RECT 42.680 146.270 43.000 146.330 ;
        RECT 62.460 146.270 62.780 146.530 ;
        RECT 67.060 146.270 67.380 146.530 ;
        RECT 71.200 146.270 71.520 146.530 ;
        RECT 74.420 146.515 74.740 146.530 ;
        RECT 74.205 146.285 74.740 146.515 ;
        RECT 74.420 146.270 74.740 146.285 ;
        RECT 89.600 146.270 89.920 146.530 ;
        RECT 95.120 146.470 95.440 146.530 ;
        RECT 96.960 146.470 97.280 146.530 ;
        RECT 95.120 146.330 97.280 146.470 ;
        RECT 95.120 146.270 95.440 146.330 ;
        RECT 96.960 146.270 97.280 146.330 ;
        RECT 39.000 146.130 39.320 146.190 ;
        RECT 45.870 146.130 46.160 146.175 ;
        RECT 48.650 146.130 48.940 146.175 ;
        RECT 50.510 146.130 50.800 146.175 ;
        RECT 39.000 145.990 42.910 146.130 ;
        RECT 39.000 145.930 39.320 145.990 ;
        RECT 38.095 145.790 38.385 145.835 ;
        RECT 41.760 145.790 42.080 145.850 ;
        RECT 38.095 145.650 42.080 145.790 ;
        RECT 42.770 145.790 42.910 145.990 ;
        RECT 45.870 145.990 50.800 146.130 ;
        RECT 45.870 145.945 46.160 145.990 ;
        RECT 48.650 145.945 48.940 145.990 ;
        RECT 50.510 145.945 50.800 145.990 ;
        RECT 51.435 145.945 51.725 146.175 ;
        RECT 64.760 146.130 65.080 146.190 ;
        RECT 73.500 146.130 73.820 146.190 ;
        RECT 64.760 145.990 73.820 146.130 ;
        RECT 46.360 145.790 46.680 145.850 ;
        RECT 42.770 145.650 46.680 145.790 ;
        RECT 38.095 145.605 38.385 145.650 ;
        RECT 41.760 145.590 42.080 145.650 ;
        RECT 46.360 145.590 46.680 145.650 ;
        RECT 49.135 145.790 49.425 145.835 ;
        RECT 51.510 145.790 51.650 145.945 ;
        RECT 64.760 145.930 65.080 145.990 ;
        RECT 73.500 145.930 73.820 145.990 ;
        RECT 78.070 146.130 78.360 146.175 ;
        RECT 80.850 146.130 81.140 146.175 ;
        RECT 82.710 146.130 83.000 146.175 ;
        RECT 78.070 145.990 83.000 146.130 ;
        RECT 78.070 145.945 78.360 145.990 ;
        RECT 80.850 145.945 81.140 145.990 ;
        RECT 82.710 145.945 83.000 145.990 ;
        RECT 91.440 146.130 91.760 146.190 ;
        RECT 101.100 146.130 101.420 146.190 ;
        RECT 91.440 145.990 99.950 146.130 ;
        RECT 91.440 145.930 91.760 145.990 ;
        RECT 49.135 145.650 51.650 145.790 ;
        RECT 56.480 145.790 56.800 145.850 ;
        RECT 57.875 145.790 58.165 145.835 ;
        RECT 58.320 145.790 58.640 145.850 ;
        RECT 56.480 145.650 58.640 145.790 ;
        RECT 49.135 145.605 49.425 145.650 ;
        RECT 56.480 145.590 56.800 145.650 ;
        RECT 57.875 145.605 58.165 145.650 ;
        RECT 58.320 145.590 58.640 145.650 ;
        RECT 58.780 145.590 59.100 145.850 ;
        RECT 66.600 145.790 66.920 145.850 ;
        RECT 64.390 145.650 66.920 145.790 ;
        RECT 21.980 145.450 22.300 145.510 ;
        RECT 28.435 145.450 28.725 145.495 ;
        RECT 36.700 145.450 37.020 145.510 ;
        RECT 21.980 145.310 37.020 145.450 ;
        RECT 21.980 145.250 22.300 145.310 ;
        RECT 28.435 145.265 28.725 145.310 ;
        RECT 36.700 145.250 37.020 145.310 ;
        RECT 39.000 145.450 39.320 145.510 ;
        RECT 39.475 145.450 39.765 145.495 ;
        RECT 39.000 145.310 39.765 145.450 ;
        RECT 39.000 145.250 39.320 145.310 ;
        RECT 39.475 145.265 39.765 145.310 ;
        RECT 39.920 145.250 40.240 145.510 ;
        RECT 40.395 145.450 40.685 145.495 ;
        RECT 41.315 145.450 41.605 145.495 ;
        RECT 44.520 145.450 44.840 145.510 ;
        RECT 40.395 145.310 41.070 145.450 ;
        RECT 40.395 145.265 40.685 145.310 ;
        RECT 40.930 144.770 41.070 145.310 ;
        RECT 41.315 145.310 44.840 145.450 ;
        RECT 41.315 145.265 41.605 145.310 ;
        RECT 44.520 145.250 44.840 145.310 ;
        RECT 45.870 145.450 46.160 145.495 ;
        RECT 50.500 145.450 50.820 145.510 ;
        RECT 50.975 145.450 51.265 145.495 ;
        RECT 45.870 145.310 48.405 145.450 ;
        RECT 45.870 145.265 46.160 145.310 ;
        RECT 42.680 145.110 43.000 145.170 ;
        RECT 48.190 145.155 48.405 145.310 ;
        RECT 50.500 145.310 51.265 145.450 ;
        RECT 50.500 145.250 50.820 145.310 ;
        RECT 50.975 145.265 51.265 145.310 ;
        RECT 52.355 145.265 52.645 145.495 ;
        RECT 55.100 145.450 55.420 145.510 ;
        RECT 57.400 145.450 57.720 145.510 ;
        RECT 55.100 145.310 57.720 145.450 ;
        RECT 44.010 145.110 44.300 145.155 ;
        RECT 47.270 145.110 47.560 145.155 ;
        RECT 42.680 144.970 47.560 145.110 ;
        RECT 42.680 144.910 43.000 144.970 ;
        RECT 44.010 144.925 44.300 144.970 ;
        RECT 47.270 144.925 47.560 144.970 ;
        RECT 48.190 145.110 48.480 145.155 ;
        RECT 50.050 145.110 50.340 145.155 ;
        RECT 48.190 144.970 50.340 145.110 ;
        RECT 48.190 144.925 48.480 144.970 ;
        RECT 50.050 144.925 50.340 144.970 ;
        RECT 42.005 144.770 42.295 144.815 ;
        RECT 45.900 144.770 46.220 144.830 ;
        RECT 40.930 144.630 46.220 144.770 ;
        RECT 42.005 144.585 42.295 144.630 ;
        RECT 45.900 144.570 46.220 144.630 ;
        RECT 49.580 144.770 49.900 144.830 ;
        RECT 52.430 144.770 52.570 145.265 ;
        RECT 55.100 145.250 55.420 145.310 ;
        RECT 57.400 145.250 57.720 145.310 ;
        RECT 59.240 145.450 59.560 145.510 ;
        RECT 62.000 145.450 62.320 145.510 ;
        RECT 64.390 145.495 64.530 145.650 ;
        RECT 66.600 145.590 66.920 145.650 ;
        RECT 70.740 145.590 71.060 145.850 ;
        RECT 83.175 145.790 83.465 145.835 ;
        RECT 84.540 145.790 84.860 145.850 ;
        RECT 83.175 145.650 84.860 145.790 ;
        RECT 83.175 145.605 83.465 145.650 ;
        RECT 84.540 145.590 84.860 145.650 ;
        RECT 89.615 145.790 89.905 145.835 ;
        RECT 90.060 145.790 90.380 145.850 ;
        RECT 89.615 145.650 90.380 145.790 ;
        RECT 89.615 145.605 89.905 145.650 ;
        RECT 90.060 145.590 90.380 145.650 ;
        RECT 98.340 145.790 98.660 145.850 ;
        RECT 99.810 145.790 99.950 145.990 ;
        RECT 101.100 145.990 105.240 146.130 ;
        RECT 101.100 145.930 101.420 145.990 ;
        RECT 103.415 145.790 103.705 145.835 ;
        RECT 104.320 145.790 104.640 145.850 ;
        RECT 98.340 145.650 99.490 145.790 ;
        RECT 99.810 145.650 104.640 145.790 ;
        RECT 105.100 145.790 105.240 145.990 ;
        RECT 110.760 145.790 111.080 145.850 ;
        RECT 105.100 145.650 111.080 145.790 ;
        RECT 98.340 145.590 98.660 145.650 ;
        RECT 59.240 145.310 62.320 145.450 ;
        RECT 59.240 145.250 59.560 145.310 ;
        RECT 62.000 145.250 62.320 145.310 ;
        RECT 64.315 145.265 64.605 145.495 ;
        RECT 66.155 145.265 66.445 145.495 ;
        RECT 68.440 145.450 68.760 145.510 ;
        RECT 70.295 145.450 70.585 145.495 ;
        RECT 68.440 145.310 70.585 145.450 ;
        RECT 66.230 145.110 66.370 145.265 ;
        RECT 68.440 145.250 68.760 145.310 ;
        RECT 70.295 145.265 70.585 145.310 ;
        RECT 71.660 145.250 71.980 145.510 ;
        RECT 78.070 145.450 78.360 145.495 ;
        RECT 78.070 145.310 80.605 145.450 ;
        RECT 78.070 145.265 78.360 145.310 ;
        RECT 79.480 145.155 79.800 145.170 ;
        RECT 61.170 144.970 66.370 145.110 ;
        RECT 76.210 145.110 76.500 145.155 ;
        RECT 79.470 145.110 79.800 145.155 ;
        RECT 76.210 144.970 79.800 145.110 ;
        RECT 49.580 144.630 52.570 144.770 ;
        RECT 58.780 144.770 59.100 144.830 ;
        RECT 61.170 144.815 61.310 144.970 ;
        RECT 76.210 144.925 76.500 144.970 ;
        RECT 79.470 144.925 79.800 144.970 ;
        RECT 80.390 145.155 80.605 145.310 ;
        RECT 81.320 145.250 81.640 145.510 ;
        RECT 88.680 145.250 89.000 145.510 ;
        RECT 97.420 145.450 97.740 145.510 ;
        RECT 99.350 145.495 99.490 145.650 ;
        RECT 103.415 145.605 103.705 145.650 ;
        RECT 104.320 145.590 104.640 145.650 ;
        RECT 98.815 145.450 99.105 145.495 ;
        RECT 97.420 145.310 99.105 145.450 ;
        RECT 97.420 145.250 97.740 145.310 ;
        RECT 98.815 145.265 99.105 145.310 ;
        RECT 99.275 145.265 99.565 145.495 ;
        RECT 99.735 145.265 100.025 145.495 ;
        RECT 100.180 145.450 100.500 145.510 ;
        RECT 100.655 145.450 100.945 145.495 ;
        RECT 100.180 145.310 100.945 145.450 ;
        RECT 80.390 145.110 80.680 145.155 ;
        RECT 82.250 145.110 82.540 145.155 ;
        RECT 80.390 144.970 82.540 145.110 ;
        RECT 80.390 144.925 80.680 144.970 ;
        RECT 82.250 144.925 82.540 144.970 ;
        RECT 79.480 144.910 79.800 144.925 ;
        RECT 90.060 144.910 90.380 145.170 ;
        RECT 99.810 145.110 99.950 145.265 ;
        RECT 100.180 145.250 100.500 145.310 ;
        RECT 100.655 145.265 100.945 145.310 ;
        RECT 104.780 145.250 105.100 145.510 ;
        RECT 108.090 145.495 108.230 145.650 ;
        RECT 110.760 145.590 111.080 145.650 ;
        RECT 108.015 145.265 108.305 145.495 ;
        RECT 99.810 144.970 102.710 145.110 ;
        RECT 102.570 144.830 102.710 144.970 ;
        RECT 59.255 144.770 59.545 144.815 ;
        RECT 58.780 144.630 59.545 144.770 ;
        RECT 49.580 144.570 49.900 144.630 ;
        RECT 58.780 144.570 59.100 144.630 ;
        RECT 59.255 144.585 59.545 144.630 ;
        RECT 61.095 144.585 61.385 144.815 ;
        RECT 64.760 144.770 65.080 144.830 ;
        RECT 65.235 144.770 65.525 144.815 ;
        RECT 64.760 144.630 65.525 144.770 ;
        RECT 64.760 144.570 65.080 144.630 ;
        RECT 65.235 144.585 65.525 144.630 ;
        RECT 69.375 144.770 69.665 144.815 ;
        RECT 70.740 144.770 71.060 144.830 ;
        RECT 69.375 144.630 71.060 144.770 ;
        RECT 69.375 144.585 69.665 144.630 ;
        RECT 70.740 144.570 71.060 144.630 ;
        RECT 87.760 144.570 88.080 144.830 ;
        RECT 95.580 144.770 95.900 144.830 ;
        RECT 97.435 144.770 97.725 144.815 ;
        RECT 95.580 144.630 97.725 144.770 ;
        RECT 95.580 144.570 95.900 144.630 ;
        RECT 97.435 144.585 97.725 144.630 ;
        RECT 102.480 144.770 102.800 144.830 ;
        RECT 104.335 144.770 104.625 144.815 ;
        RECT 102.480 144.630 104.625 144.770 ;
        RECT 102.480 144.570 102.800 144.630 ;
        RECT 104.335 144.585 104.625 144.630 ;
        RECT 106.635 144.770 106.925 144.815 ;
        RECT 107.080 144.770 107.400 144.830 ;
        RECT 106.635 144.630 107.400 144.770 ;
        RECT 106.635 144.585 106.925 144.630 ;
        RECT 107.080 144.570 107.400 144.630 ;
        RECT 107.555 144.770 107.845 144.815 ;
        RECT 108.000 144.770 108.320 144.830 ;
        RECT 107.555 144.630 108.320 144.770 ;
        RECT 107.555 144.585 107.845 144.630 ;
        RECT 108.000 144.570 108.320 144.630 ;
        RECT 15.010 143.950 113.450 144.430 ;
        RECT 33.035 143.750 33.325 143.795 ;
        RECT 35.780 143.750 36.100 143.810 ;
        RECT 33.035 143.610 36.100 143.750 ;
        RECT 33.035 143.565 33.325 143.610 ;
        RECT 35.780 143.550 36.100 143.610 ;
        RECT 42.680 143.550 43.000 143.810 ;
        RECT 45.455 143.750 45.745 143.795 ;
        RECT 45.900 143.750 46.220 143.810 ;
        RECT 55.575 143.750 55.865 143.795 ;
        RECT 65.220 143.750 65.540 143.810 ;
        RECT 45.455 143.610 46.220 143.750 ;
        RECT 45.455 143.565 45.745 143.610 ;
        RECT 45.900 143.550 46.220 143.610 ;
        RECT 52.430 143.610 55.865 143.750 ;
        RECT 30.350 143.270 33.250 143.410 ;
        RECT 30.350 143.130 30.490 143.270 ;
        RECT 23.360 142.870 23.680 143.130 ;
        RECT 30.260 142.870 30.580 143.130 ;
        RECT 31.180 142.870 31.500 143.130 ;
        RECT 32.575 142.885 32.865 143.115 ;
        RECT 30.720 142.730 31.040 142.790 ;
        RECT 31.655 142.730 31.945 142.775 ;
        RECT 30.720 142.590 31.945 142.730 ;
        RECT 30.720 142.530 31.040 142.590 ;
        RECT 31.655 142.545 31.945 142.590 ;
        RECT 26.120 142.390 26.440 142.450 ;
        RECT 30.275 142.390 30.565 142.435 ;
        RECT 32.100 142.390 32.420 142.450 ;
        RECT 26.120 142.250 30.565 142.390 ;
        RECT 26.120 142.190 26.440 142.250 ;
        RECT 30.275 142.205 30.565 142.250 ;
        RECT 31.730 142.250 32.420 142.390 ;
        RECT 32.650 142.390 32.790 142.885 ;
        RECT 33.110 142.730 33.250 143.270 ;
        RECT 34.860 143.210 35.180 143.470 ;
        RECT 35.335 143.410 35.625 143.455 ;
        RECT 52.430 143.410 52.570 143.610 ;
        RECT 55.575 143.565 55.865 143.610 ;
        RECT 56.110 143.610 65.540 143.750 ;
        RECT 56.110 143.410 56.250 143.610 ;
        RECT 35.335 143.270 52.570 143.410 ;
        RECT 53.810 143.270 56.250 143.410 ;
        RECT 35.335 143.225 35.625 143.270 ;
        RECT 33.955 143.070 34.245 143.115 ;
        RECT 34.950 143.070 35.090 143.210 ;
        RECT 33.955 142.930 35.090 143.070 ;
        RECT 36.700 143.070 37.020 143.130 ;
        RECT 39.015 143.070 39.305 143.115 ;
        RECT 42.235 143.070 42.525 143.115 ;
        RECT 42.680 143.070 43.000 143.130 ;
        RECT 45.440 143.070 45.760 143.130 ;
        RECT 36.700 142.930 43.000 143.070 ;
        RECT 33.955 142.885 34.245 142.930 ;
        RECT 36.700 142.870 37.020 142.930 ;
        RECT 39.015 142.885 39.305 142.930 ;
        RECT 42.235 142.885 42.525 142.930 ;
        RECT 42.680 142.870 43.000 142.930 ;
        RECT 44.610 142.930 45.760 143.070 ;
        RECT 44.610 142.775 44.750 142.930 ;
        RECT 45.440 142.870 45.760 142.930 ;
        RECT 49.135 143.070 49.425 143.115 ;
        RECT 49.580 143.070 49.900 143.130 ;
        RECT 49.135 142.930 49.900 143.070 ;
        RECT 49.135 142.885 49.425 142.930 ;
        RECT 49.580 142.870 49.900 142.930 ;
        RECT 50.040 142.870 50.360 143.130 ;
        RECT 53.810 143.115 53.950 143.270 ;
        RECT 50.515 142.885 50.805 143.115 ;
        RECT 53.275 142.885 53.565 143.115 ;
        RECT 53.735 142.885 54.025 143.115 ;
        RECT 54.195 142.885 54.485 143.115 ;
        RECT 34.415 142.730 34.705 142.775 ;
        RECT 33.110 142.590 34.705 142.730 ;
        RECT 34.415 142.545 34.705 142.590 ;
        RECT 44.535 142.545 44.825 142.775 ;
        RECT 44.980 142.530 45.300 142.790 ;
        RECT 46.820 142.730 47.140 142.790 ;
        RECT 50.590 142.730 50.730 142.885 ;
        RECT 46.820 142.590 50.730 142.730 ;
        RECT 46.820 142.530 47.140 142.590 ;
        RECT 51.895 142.390 52.185 142.435 ;
        RECT 32.650 142.250 52.185 142.390 ;
        RECT 53.350 142.390 53.490 142.885 ;
        RECT 54.270 142.730 54.410 142.885 ;
        RECT 55.100 142.870 55.420 143.130 ;
        RECT 56.940 142.870 57.260 143.130 ;
        RECT 57.490 143.115 57.630 143.610 ;
        RECT 65.220 143.550 65.540 143.610 ;
        RECT 80.415 143.750 80.705 143.795 ;
        RECT 81.320 143.750 81.640 143.810 ;
        RECT 80.415 143.610 81.640 143.750 ;
        RECT 80.415 143.565 80.705 143.610 ;
        RECT 81.320 143.550 81.640 143.610 ;
        RECT 89.140 143.550 89.460 143.810 ;
        RECT 90.060 143.750 90.380 143.810 ;
        RECT 91.455 143.750 91.745 143.795 ;
        RECT 98.340 143.750 98.660 143.810 ;
        RECT 90.060 143.610 91.745 143.750 ;
        RECT 90.060 143.550 90.380 143.610 ;
        RECT 91.455 143.565 91.745 143.610 ;
        RECT 97.510 143.610 98.660 143.750 ;
        RECT 61.490 143.410 61.780 143.455 ;
        RECT 62.920 143.410 63.240 143.470 ;
        RECT 64.750 143.410 65.040 143.455 ;
        RECT 61.490 143.270 65.040 143.410 ;
        RECT 61.490 143.225 61.780 143.270 ;
        RECT 62.920 143.210 63.240 143.270 ;
        RECT 64.750 143.225 65.040 143.270 ;
        RECT 65.670 143.410 65.960 143.455 ;
        RECT 67.530 143.410 67.820 143.455 ;
        RECT 65.670 143.270 67.820 143.410 ;
        RECT 65.670 143.225 65.960 143.270 ;
        RECT 67.530 143.225 67.820 143.270 ;
        RECT 75.340 143.410 75.660 143.470 ;
        RECT 85.015 143.410 85.305 143.455 ;
        RECT 75.340 143.270 85.305 143.410 ;
        RECT 57.415 142.885 57.705 143.115 ;
        RECT 57.875 143.070 58.165 143.115 ;
        RECT 58.320 143.070 58.640 143.130 ;
        RECT 57.875 142.930 58.640 143.070 ;
        RECT 57.875 142.885 58.165 142.930 ;
        RECT 58.320 142.870 58.640 142.930 ;
        RECT 58.795 143.070 59.085 143.115 ;
        RECT 59.240 143.070 59.560 143.130 ;
        RECT 58.795 142.930 59.560 143.070 ;
        RECT 58.795 142.885 59.085 142.930 ;
        RECT 59.240 142.870 59.560 142.930 ;
        RECT 63.350 143.070 63.640 143.115 ;
        RECT 65.670 143.070 65.885 143.225 ;
        RECT 75.340 143.210 75.660 143.270 ;
        RECT 85.015 143.225 85.305 143.270 ;
        RECT 85.475 143.410 85.765 143.455 ;
        RECT 89.230 143.410 89.370 143.550 ;
        RECT 93.295 143.410 93.585 143.455 ;
        RECT 85.475 143.270 93.585 143.410 ;
        RECT 85.475 143.225 85.765 143.270 ;
        RECT 93.295 143.225 93.585 143.270 ;
        RECT 93.740 143.210 94.060 143.470 ;
        RECT 94.200 143.410 94.520 143.470 ;
        RECT 97.510 143.410 97.650 143.610 ;
        RECT 98.340 143.550 98.660 143.610 ;
        RECT 102.480 143.455 102.800 143.470 ;
        RECT 108.000 143.455 108.320 143.470 ;
        RECT 94.200 143.270 98.110 143.410 ;
        RECT 94.200 143.210 94.520 143.270 ;
        RECT 67.980 143.070 68.300 143.130 ;
        RECT 68.455 143.070 68.745 143.115 ;
        RECT 63.350 142.930 65.885 143.070 ;
        RECT 66.230 142.930 67.750 143.070 ;
        RECT 63.350 142.885 63.640 142.930 ;
        RECT 59.330 142.730 59.470 142.870 ;
        RECT 66.230 142.730 66.370 142.930 ;
        RECT 54.270 142.590 59.010 142.730 ;
        RECT 59.330 142.590 66.370 142.730 ;
        RECT 56.940 142.390 57.260 142.450 ;
        RECT 53.350 142.250 57.260 142.390 ;
        RECT 19.680 142.050 20.000 142.110 ;
        RECT 23.360 142.050 23.680 142.110 ;
        RECT 19.680 141.910 23.680 142.050 ;
        RECT 19.680 141.850 20.000 141.910 ;
        RECT 23.360 141.850 23.680 141.910 ;
        RECT 23.820 141.850 24.140 142.110 ;
        RECT 31.730 142.095 31.870 142.250 ;
        RECT 32.100 142.190 32.420 142.250 ;
        RECT 51.895 142.205 52.185 142.250 ;
        RECT 56.940 142.190 57.260 142.250 ;
        RECT 58.870 142.110 59.010 142.590 ;
        RECT 66.600 142.530 66.920 142.790 ;
        RECT 67.610 142.730 67.750 142.930 ;
        RECT 67.980 142.930 68.745 143.070 ;
        RECT 67.980 142.870 68.300 142.930 ;
        RECT 68.455 142.885 68.745 142.930 ;
        RECT 79.495 143.070 79.785 143.115 ;
        RECT 79.940 143.070 80.260 143.130 ;
        RECT 87.300 143.070 87.620 143.130 ;
        RECT 89.140 143.115 89.460 143.130 ;
        RECT 88.235 143.070 88.525 143.115 ;
        RECT 89.130 143.070 89.460 143.115 ;
        RECT 79.495 142.930 80.260 143.070 ;
        RECT 79.495 142.885 79.785 142.930 ;
        RECT 79.940 142.870 80.260 142.930 ;
        RECT 84.170 142.930 88.525 143.070 ;
        RECT 88.945 142.930 89.460 143.070 ;
        RECT 84.170 142.730 84.310 142.930 ;
        RECT 87.300 142.870 87.620 142.930 ;
        RECT 88.235 142.885 88.525 142.930 ;
        RECT 89.130 142.885 89.460 142.930 ;
        RECT 89.615 142.885 89.905 143.115 ;
        RECT 90.075 143.070 90.365 143.115 ;
        RECT 97.420 143.070 97.740 143.130 ;
        RECT 97.970 143.115 98.110 143.270 ;
        RECT 102.480 143.225 103.015 143.455 ;
        RECT 104.730 143.410 105.020 143.455 ;
        RECT 107.990 143.410 108.320 143.455 ;
        RECT 104.730 143.270 108.320 143.410 ;
        RECT 104.730 143.225 105.020 143.270 ;
        RECT 107.990 143.225 108.320 143.270 ;
        RECT 102.480 143.210 102.800 143.225 ;
        RECT 108.000 143.210 108.320 143.225 ;
        RECT 108.910 143.410 109.200 143.455 ;
        RECT 110.770 143.410 111.060 143.455 ;
        RECT 108.910 143.270 111.060 143.410 ;
        RECT 108.910 143.225 109.200 143.270 ;
        RECT 110.770 143.225 111.060 143.270 ;
        RECT 90.075 142.930 97.740 143.070 ;
        RECT 90.075 142.885 90.365 142.930 ;
        RECT 89.140 142.870 89.460 142.885 ;
        RECT 67.610 142.590 84.310 142.730 ;
        RECT 84.555 142.545 84.845 142.775 ;
        RECT 89.690 142.730 89.830 142.885 ;
        RECT 90.610 142.790 90.750 142.930 ;
        RECT 97.420 142.870 97.740 142.930 ;
        RECT 97.895 142.885 98.185 143.115 ;
        RECT 98.355 143.070 98.645 143.115 ;
        RECT 98.800 143.070 99.120 143.130 ;
        RECT 98.355 142.930 99.120 143.070 ;
        RECT 98.355 142.885 98.645 142.930 ;
        RECT 89.690 142.590 90.290 142.730 ;
        RECT 63.350 142.390 63.640 142.435 ;
        RECT 66.130 142.390 66.420 142.435 ;
        RECT 67.990 142.390 68.280 142.435 ;
        RECT 63.350 142.250 68.280 142.390 ;
        RECT 63.350 142.205 63.640 142.250 ;
        RECT 66.130 142.205 66.420 142.250 ;
        RECT 67.990 142.205 68.280 142.250 ;
        RECT 84.080 142.390 84.400 142.450 ;
        RECT 84.630 142.390 84.770 142.545 ;
        RECT 90.150 142.390 90.290 142.590 ;
        RECT 90.520 142.530 90.840 142.790 ;
        RECT 92.360 142.530 92.680 142.790 ;
        RECT 93.740 142.730 94.060 142.790 ;
        RECT 98.430 142.730 98.570 142.885 ;
        RECT 98.800 142.870 99.120 142.930 ;
        RECT 99.275 143.070 99.565 143.115 ;
        RECT 99.720 143.070 100.040 143.130 ;
        RECT 99.275 142.930 100.040 143.070 ;
        RECT 99.275 142.885 99.565 142.930 ;
        RECT 99.720 142.870 100.040 142.930 ;
        RECT 101.100 142.870 101.420 143.130 ;
        RECT 106.590 143.070 106.880 143.115 ;
        RECT 108.910 143.070 109.125 143.225 ;
        RECT 106.590 142.930 109.125 143.070 ;
        RECT 106.590 142.885 106.880 142.930 ;
        RECT 93.740 142.590 98.570 142.730 ;
        RECT 93.740 142.530 94.060 142.590 ;
        RECT 109.840 142.530 110.160 142.790 ;
        RECT 111.680 142.530 112.000 142.790 ;
        RECT 94.200 142.390 94.520 142.450 ;
        RECT 84.080 142.250 88.220 142.390 ;
        RECT 90.150 142.250 94.520 142.390 ;
        RECT 84.080 142.190 84.400 142.250 ;
        RECT 31.655 141.865 31.945 142.095 ;
        RECT 33.940 141.850 34.260 142.110 ;
        RECT 39.475 142.050 39.765 142.095 ;
        RECT 39.920 142.050 40.240 142.110 ;
        RECT 39.475 141.910 40.240 142.050 ;
        RECT 39.475 141.865 39.765 141.910 ;
        RECT 39.920 141.850 40.240 141.910 ;
        RECT 46.820 142.050 47.140 142.110 ;
        RECT 47.295 142.050 47.585 142.095 ;
        RECT 46.820 141.910 47.585 142.050 ;
        RECT 46.820 141.850 47.140 141.910 ;
        RECT 47.295 141.865 47.585 141.910 ;
        RECT 49.595 142.050 49.885 142.095 ;
        RECT 50.040 142.050 50.360 142.110 ;
        RECT 49.595 141.910 50.360 142.050 ;
        RECT 49.595 141.865 49.885 141.910 ;
        RECT 50.040 141.850 50.360 141.910 ;
        RECT 51.435 142.050 51.725 142.095 ;
        RECT 54.180 142.050 54.500 142.110 ;
        RECT 51.435 141.910 54.500 142.050 ;
        RECT 51.435 141.865 51.725 141.910 ;
        RECT 54.180 141.850 54.500 141.910 ;
        RECT 58.780 142.050 59.100 142.110 ;
        RECT 59.485 142.050 59.775 142.095 ;
        RECT 58.780 141.910 59.775 142.050 ;
        RECT 58.780 141.850 59.100 141.910 ;
        RECT 59.485 141.865 59.775 141.910 ;
        RECT 60.620 142.050 60.940 142.110 ;
        RECT 86.840 142.050 87.160 142.110 ;
        RECT 60.620 141.910 87.160 142.050 ;
        RECT 60.620 141.850 60.940 141.910 ;
        RECT 86.840 141.850 87.160 141.910 ;
        RECT 87.300 141.850 87.620 142.110 ;
        RECT 88.080 142.050 88.220 142.250 ;
        RECT 94.200 142.190 94.520 142.250 ;
        RECT 95.595 142.390 95.885 142.435 ;
        RECT 98.340 142.390 98.660 142.450 ;
        RECT 95.595 142.250 98.660 142.390 ;
        RECT 95.595 142.205 95.885 142.250 ;
        RECT 98.340 142.190 98.660 142.250 ;
        RECT 106.590 142.390 106.880 142.435 ;
        RECT 109.370 142.390 109.660 142.435 ;
        RECT 111.230 142.390 111.520 142.435 ;
        RECT 106.590 142.250 111.520 142.390 ;
        RECT 106.590 142.205 106.880 142.250 ;
        RECT 109.370 142.205 109.660 142.250 ;
        RECT 111.230 142.205 111.520 142.250 ;
        RECT 91.440 142.050 91.760 142.110 ;
        RECT 92.360 142.050 92.680 142.110 ;
        RECT 88.080 141.910 92.680 142.050 ;
        RECT 91.440 141.850 91.760 141.910 ;
        RECT 92.360 141.850 92.680 141.910 ;
        RECT 95.120 142.050 95.440 142.110 ;
        RECT 96.055 142.050 96.345 142.095 ;
        RECT 95.120 141.910 96.345 142.050 ;
        RECT 95.120 141.850 95.440 141.910 ;
        RECT 96.055 141.865 96.345 141.910 ;
        RECT 101.560 141.850 101.880 142.110 ;
        RECT 15.010 141.230 113.450 141.710 ;
        RECT 135.635 141.220 136.775 165.470 ;
        RECT 18.315 141.030 18.605 141.075 ;
        RECT 20.140 141.030 20.460 141.090 ;
        RECT 18.315 140.890 20.460 141.030 ;
        RECT 18.315 140.845 18.605 140.890 ;
        RECT 20.140 140.830 20.460 140.890 ;
        RECT 32.100 141.030 32.420 141.090 ;
        RECT 32.575 141.030 32.865 141.075 ;
        RECT 32.100 140.890 32.865 141.030 ;
        RECT 32.100 140.830 32.420 140.890 ;
        RECT 32.575 140.845 32.865 140.890 ;
        RECT 35.320 140.830 35.640 141.090 ;
        RECT 44.520 141.030 44.840 141.090 ;
        RECT 49.580 141.030 49.900 141.090 ;
        RECT 50.515 141.030 50.805 141.075 ;
        RECT 44.520 140.890 47.510 141.030 ;
        RECT 44.520 140.830 44.840 140.890 ;
        RECT 20.620 140.690 20.910 140.735 ;
        RECT 22.480 140.690 22.770 140.735 ;
        RECT 25.260 140.690 25.550 140.735 ;
        RECT 20.620 140.550 25.550 140.690 ;
        RECT 20.620 140.505 20.910 140.550 ;
        RECT 22.480 140.505 22.770 140.550 ;
        RECT 25.260 140.505 25.550 140.550 ;
        RECT 26.580 140.690 26.900 140.750 ;
        RECT 33.940 140.690 34.260 140.750 ;
        RECT 26.580 140.550 34.260 140.690 ;
        RECT 26.580 140.490 26.900 140.550 ;
        RECT 33.940 140.490 34.260 140.550 ;
        RECT 36.720 140.690 37.010 140.735 ;
        RECT 38.580 140.690 38.870 140.735 ;
        RECT 41.360 140.690 41.650 140.735 ;
        RECT 36.720 140.550 41.650 140.690 ;
        RECT 36.720 140.505 37.010 140.550 ;
        RECT 38.580 140.505 38.870 140.550 ;
        RECT 41.360 140.505 41.650 140.550 ;
        RECT 45.915 140.505 46.205 140.735 ;
        RECT 18.300 140.350 18.620 140.410 ;
        RECT 21.995 140.350 22.285 140.395 ;
        RECT 38.095 140.350 38.385 140.395 ;
        RECT 45.990 140.350 46.130 140.505 ;
        RECT 18.300 140.210 22.285 140.350 ;
        RECT 18.300 140.150 18.620 140.210 ;
        RECT 21.995 140.165 22.285 140.210 ;
        RECT 31.730 140.210 34.630 140.350 ;
        RECT 17.395 140.010 17.685 140.055 ;
        RECT 18.760 140.010 19.080 140.070 ;
        RECT 17.395 139.870 19.080 140.010 ;
        RECT 17.395 139.825 17.685 139.870 ;
        RECT 18.760 139.810 19.080 139.870 ;
        RECT 19.680 139.810 20.000 140.070 ;
        RECT 20.155 140.010 20.445 140.055 ;
        RECT 22.440 140.010 22.760 140.070 ;
        RECT 28.880 140.055 29.200 140.070 ;
        RECT 31.730 140.055 31.870 140.210 ;
        RECT 34.490 140.055 34.630 140.210 ;
        RECT 38.095 140.210 46.130 140.350 ;
        RECT 38.095 140.165 38.385 140.210 ;
        RECT 25.260 140.010 25.550 140.055 ;
        RECT 20.155 139.870 22.760 140.010 ;
        RECT 20.155 139.825 20.445 139.870 ;
        RECT 22.440 139.810 22.760 139.870 ;
        RECT 23.015 139.870 25.550 140.010 ;
        RECT 23.015 139.715 23.230 139.870 ;
        RECT 25.260 139.825 25.550 139.870 ;
        RECT 28.880 140.010 29.415 140.055 ;
        RECT 30.735 140.010 31.025 140.055 ;
        RECT 28.880 139.870 31.025 140.010 ;
        RECT 28.880 139.825 29.415 139.870 ;
        RECT 30.735 139.825 31.025 139.870 ;
        RECT 31.655 139.825 31.945 140.055 ;
        RECT 33.495 139.825 33.785 140.055 ;
        RECT 34.415 140.010 34.705 140.055 ;
        RECT 35.320 140.010 35.640 140.070 ;
        RECT 34.415 139.870 35.640 140.010 ;
        RECT 34.415 139.825 34.705 139.870 ;
        RECT 28.880 139.810 29.200 139.825 ;
        RECT 21.080 139.670 21.370 139.715 ;
        RECT 22.940 139.670 23.230 139.715 ;
        RECT 21.080 139.530 23.230 139.670 ;
        RECT 21.080 139.485 21.370 139.530 ;
        RECT 22.940 139.485 23.230 139.530 ;
        RECT 23.820 139.715 24.140 139.730 ;
        RECT 23.820 139.670 24.150 139.715 ;
        RECT 27.120 139.670 27.410 139.715 ;
        RECT 23.820 139.530 27.410 139.670 ;
        RECT 23.820 139.485 24.150 139.530 ;
        RECT 27.120 139.485 27.410 139.530 ;
        RECT 23.820 139.470 24.140 139.485 ;
        RECT 19.235 139.330 19.525 139.375 ;
        RECT 19.680 139.330 20.000 139.390 ;
        RECT 19.235 139.190 20.000 139.330 ;
        RECT 19.235 139.145 19.525 139.190 ;
        RECT 19.680 139.130 20.000 139.190 ;
        RECT 20.600 139.330 20.920 139.390 ;
        RECT 33.570 139.330 33.710 139.825 ;
        RECT 35.320 139.810 35.640 139.870 ;
        RECT 36.240 139.810 36.560 140.070 ;
        RECT 41.360 140.010 41.650 140.055 ;
        RECT 39.115 139.870 41.650 140.010 ;
        RECT 39.115 139.715 39.330 139.870 ;
        RECT 41.360 139.825 41.650 139.870 ;
        RECT 46.820 139.810 47.140 140.070 ;
        RECT 47.370 140.055 47.510 140.890 ;
        RECT 49.580 140.890 50.805 141.030 ;
        RECT 49.580 140.830 49.900 140.890 ;
        RECT 50.515 140.845 50.805 140.890 ;
        RECT 57.400 141.030 57.720 141.090 ;
        RECT 59.240 141.030 59.560 141.090 ;
        RECT 57.400 140.890 59.560 141.030 ;
        RECT 57.400 140.830 57.720 140.890 ;
        RECT 59.240 140.830 59.560 140.890 ;
        RECT 62.920 141.030 63.240 141.090 ;
        RECT 63.395 141.030 63.685 141.075 ;
        RECT 62.920 140.890 63.685 141.030 ;
        RECT 62.920 140.830 63.240 140.890 ;
        RECT 63.395 140.845 63.685 140.890 ;
        RECT 65.695 141.030 65.985 141.075 ;
        RECT 66.600 141.030 66.920 141.090 ;
        RECT 65.695 140.890 66.920 141.030 ;
        RECT 65.695 140.845 65.985 140.890 ;
        RECT 66.600 140.830 66.920 140.890 ;
        RECT 72.135 140.845 72.425 141.075 ;
        RECT 73.055 141.030 73.345 141.075 ;
        RECT 85.920 141.030 86.240 141.090 ;
        RECT 73.055 140.890 86.240 141.030 ;
        RECT 73.055 140.845 73.345 140.890 ;
        RECT 61.095 140.505 61.385 140.735 ;
        RECT 72.210 140.690 72.350 140.845 ;
        RECT 85.920 140.830 86.240 140.890 ;
        RECT 88.005 141.030 88.295 141.075 ;
        RECT 89.140 141.030 89.460 141.090 ;
        RECT 88.005 140.890 89.460 141.030 ;
        RECT 88.005 140.845 88.295 140.890 ;
        RECT 89.140 140.830 89.460 140.890 ;
        RECT 109.840 140.830 110.160 141.090 ;
        RECT 73.500 140.690 73.820 140.750 ;
        RECT 76.260 140.690 76.580 140.750 ;
        RECT 72.210 140.550 73.820 140.690 ;
        RECT 50.960 140.350 51.280 140.410 ;
        RECT 48.750 140.210 51.280 140.350 ;
        RECT 48.750 140.070 48.890 140.210 ;
        RECT 50.960 140.150 51.280 140.210 ;
        RECT 51.895 140.350 52.185 140.395 ;
        RECT 55.100 140.350 55.420 140.410 ;
        RECT 56.480 140.350 56.800 140.410 ;
        RECT 57.875 140.350 58.165 140.395 ;
        RECT 51.895 140.210 58.165 140.350 ;
        RECT 51.895 140.165 52.185 140.210 ;
        RECT 55.100 140.150 55.420 140.210 ;
        RECT 56.480 140.150 56.800 140.210 ;
        RECT 57.875 140.165 58.165 140.210 ;
        RECT 58.780 140.150 59.100 140.410 ;
        RECT 61.170 140.350 61.310 140.505 ;
        RECT 73.500 140.490 73.820 140.550 ;
        RECT 74.510 140.550 76.580 140.690 ;
        RECT 61.170 140.210 64.990 140.350 ;
        RECT 47.295 140.010 47.585 140.055 ;
        RECT 47.740 140.010 48.060 140.070 ;
        RECT 47.295 139.870 48.060 140.010 ;
        RECT 47.295 139.825 47.585 139.870 ;
        RECT 47.740 139.810 48.060 139.870 ;
        RECT 48.215 139.825 48.505 140.055 ;
        RECT 37.180 139.670 37.470 139.715 ;
        RECT 39.040 139.670 39.330 139.715 ;
        RECT 37.180 139.530 39.330 139.670 ;
        RECT 37.180 139.485 37.470 139.530 ;
        RECT 39.040 139.485 39.330 139.530 ;
        RECT 39.920 139.715 40.240 139.730 ;
        RECT 44.980 139.715 45.300 139.730 ;
        RECT 39.920 139.670 40.250 139.715 ;
        RECT 43.220 139.670 43.510 139.715 ;
        RECT 39.920 139.530 43.510 139.670 ;
        RECT 39.920 139.485 40.250 139.530 ;
        RECT 43.220 139.485 43.510 139.530 ;
        RECT 44.980 139.670 45.515 139.715 ;
        RECT 48.290 139.670 48.430 139.825 ;
        RECT 48.660 139.810 48.980 140.070 ;
        RECT 49.120 139.810 49.440 140.070 ;
        RECT 55.575 140.010 55.865 140.055 ;
        RECT 54.730 139.870 55.865 140.010 ;
        RECT 52.815 139.670 53.105 139.715 ;
        RECT 44.980 139.530 53.105 139.670 ;
        RECT 44.980 139.485 45.515 139.530 ;
        RECT 52.815 139.485 53.105 139.530 ;
        RECT 39.920 139.470 40.240 139.485 ;
        RECT 44.980 139.470 45.300 139.485 ;
        RECT 20.600 139.190 33.710 139.330 ;
        RECT 46.360 139.330 46.680 139.390 ;
        RECT 49.120 139.330 49.440 139.390 ;
        RECT 46.360 139.190 49.440 139.330 ;
        RECT 20.600 139.130 20.920 139.190 ;
        RECT 46.360 139.130 46.680 139.190 ;
        RECT 49.120 139.130 49.440 139.190 ;
        RECT 52.340 139.130 52.660 139.390 ;
        RECT 54.730 139.375 54.870 139.870 ;
        RECT 55.575 139.825 55.865 139.870 ;
        RECT 62.000 140.010 62.320 140.070 ;
        RECT 64.850 140.055 64.990 140.210 ;
        RECT 70.740 140.150 71.060 140.410 ;
        RECT 71.660 140.150 71.980 140.410 ;
        RECT 74.510 140.395 74.650 140.550 ;
        RECT 76.260 140.490 76.580 140.550 ;
        RECT 81.750 140.690 82.040 140.735 ;
        RECT 84.530 140.690 84.820 140.735 ;
        RECT 86.390 140.690 86.680 140.735 ;
        RECT 81.750 140.550 86.680 140.690 ;
        RECT 81.750 140.505 82.040 140.550 ;
        RECT 84.530 140.505 84.820 140.550 ;
        RECT 86.390 140.505 86.680 140.550 ;
        RECT 91.870 140.690 92.160 140.735 ;
        RECT 94.650 140.690 94.940 140.735 ;
        RECT 96.510 140.690 96.800 140.735 ;
        RECT 97.435 140.690 97.725 140.735 ;
        RECT 91.870 140.550 96.800 140.690 ;
        RECT 91.870 140.505 92.160 140.550 ;
        RECT 94.650 140.505 94.940 140.550 ;
        RECT 96.510 140.505 96.800 140.550 ;
        RECT 97.050 140.550 97.725 140.690 ;
        RECT 74.435 140.165 74.725 140.395 ;
        RECT 74.880 140.150 75.200 140.410 ;
        RECT 85.015 140.350 85.305 140.395 ;
        RECT 85.460 140.350 85.780 140.410 ;
        RECT 90.980 140.350 91.300 140.410 ;
        RECT 95.135 140.350 95.425 140.395 ;
        RECT 97.050 140.350 97.190 140.550 ;
        RECT 97.435 140.505 97.725 140.550 ;
        RECT 103.370 140.690 103.660 140.735 ;
        RECT 106.150 140.690 106.440 140.735 ;
        RECT 108.010 140.690 108.300 140.735 ;
        RECT 103.370 140.550 108.300 140.690 ;
        RECT 103.370 140.505 103.660 140.550 ;
        RECT 106.150 140.505 106.440 140.550 ;
        RECT 108.010 140.505 108.300 140.550 ;
        RECT 85.015 140.210 85.780 140.350 ;
        RECT 85.015 140.165 85.305 140.210 ;
        RECT 85.460 140.150 85.780 140.210 ;
        RECT 86.930 140.210 94.890 140.350 ;
        RECT 63.855 140.010 64.145 140.055 ;
        RECT 62.000 139.870 64.145 140.010 ;
        RECT 62.000 139.810 62.320 139.870 ;
        RECT 63.855 139.825 64.145 139.870 ;
        RECT 64.775 139.825 65.065 140.055 ;
        RECT 70.830 140.010 70.970 140.150 ;
        RECT 72.135 140.010 72.425 140.055 ;
        RECT 72.580 140.010 72.900 140.070 ;
        RECT 70.830 139.870 71.890 140.010 ;
        RECT 71.750 139.730 71.890 139.870 ;
        RECT 72.135 139.870 72.900 140.010 ;
        RECT 72.135 139.825 72.425 139.870 ;
        RECT 72.580 139.810 72.900 139.870 ;
        RECT 81.750 140.010 82.040 140.055 ;
        RECT 84.540 140.010 84.860 140.070 ;
        RECT 86.930 140.055 87.070 140.210 ;
        RECT 90.980 140.150 91.300 140.210 ;
        RECT 86.855 140.010 87.145 140.055 ;
        RECT 81.750 139.870 84.285 140.010 ;
        RECT 81.750 139.825 82.040 139.870 ;
        RECT 70.740 139.470 71.060 139.730 ;
        RECT 71.660 139.470 71.980 139.730 ;
        RECT 84.070 139.715 84.285 139.870 ;
        RECT 84.540 139.870 87.145 140.010 ;
        RECT 84.540 139.810 84.860 139.870 ;
        RECT 86.855 139.825 87.145 139.870 ;
        RECT 91.870 140.010 92.160 140.055 ;
        RECT 94.750 140.010 94.890 140.210 ;
        RECT 95.135 140.210 97.190 140.350 ;
        RECT 97.510 140.210 106.390 140.350 ;
        RECT 95.135 140.165 95.425 140.210 ;
        RECT 96.975 140.010 97.265 140.055 ;
        RECT 97.510 140.010 97.650 140.210 ;
        RECT 91.870 139.870 94.405 140.010 ;
        RECT 94.750 139.870 97.650 140.010 ;
        RECT 91.870 139.825 92.160 139.870 ;
        RECT 77.885 139.670 78.175 139.715 ;
        RECT 75.430 139.530 78.175 139.670 ;
        RECT 75.430 139.390 75.570 139.530 ;
        RECT 77.885 139.485 78.175 139.530 ;
        RECT 79.890 139.670 80.180 139.715 ;
        RECT 83.150 139.670 83.440 139.715 ;
        RECT 84.070 139.670 84.360 139.715 ;
        RECT 85.930 139.670 86.220 139.715 ;
        RECT 79.890 139.530 83.850 139.670 ;
        RECT 79.890 139.485 80.180 139.530 ;
        RECT 83.150 139.485 83.440 139.530 ;
        RECT 83.710 139.390 83.850 139.530 ;
        RECT 84.070 139.530 86.220 139.670 ;
        RECT 84.070 139.485 84.360 139.530 ;
        RECT 85.930 139.485 86.220 139.530 ;
        RECT 90.010 139.670 90.300 139.715 ;
        RECT 90.520 139.670 90.840 139.730 ;
        RECT 94.190 139.715 94.405 139.870 ;
        RECT 96.975 139.825 97.265 139.870 ;
        RECT 98.340 139.810 98.660 140.070 ;
        RECT 103.370 140.010 103.660 140.055 ;
        RECT 106.250 140.010 106.390 140.210 ;
        RECT 106.620 140.150 106.940 140.410 ;
        RECT 108.475 140.350 108.765 140.395 ;
        RECT 111.680 140.350 112.000 140.410 ;
        RECT 108.475 140.210 112.000 140.350 ;
        RECT 135.580 140.230 136.830 141.220 ;
        RECT 108.475 140.165 108.765 140.210 ;
        RECT 108.550 140.010 108.690 140.165 ;
        RECT 111.680 140.150 112.000 140.210 ;
        RECT 135.635 140.155 136.775 140.230 ;
        RECT 103.370 139.870 105.905 140.010 ;
        RECT 106.250 139.870 108.690 140.010 ;
        RECT 103.370 139.825 103.660 139.870 ;
        RECT 101.560 139.715 101.880 139.730 ;
        RECT 105.690 139.715 105.905 139.870 ;
        RECT 108.935 139.825 109.225 140.055 ;
        RECT 93.270 139.670 93.560 139.715 ;
        RECT 90.010 139.530 93.560 139.670 ;
        RECT 90.010 139.485 90.300 139.530 ;
        RECT 90.520 139.470 90.840 139.530 ;
        RECT 93.270 139.485 93.560 139.530 ;
        RECT 94.190 139.670 94.480 139.715 ;
        RECT 96.050 139.670 96.340 139.715 ;
        RECT 94.190 139.530 96.340 139.670 ;
        RECT 94.190 139.485 94.480 139.530 ;
        RECT 96.050 139.485 96.340 139.530 ;
        RECT 101.510 139.670 101.880 139.715 ;
        RECT 104.770 139.670 105.060 139.715 ;
        RECT 101.510 139.530 105.060 139.670 ;
        RECT 101.510 139.485 101.880 139.530 ;
        RECT 104.770 139.485 105.060 139.530 ;
        RECT 105.690 139.670 105.980 139.715 ;
        RECT 107.550 139.670 107.840 139.715 ;
        RECT 105.690 139.530 107.840 139.670 ;
        RECT 105.690 139.485 105.980 139.530 ;
        RECT 107.550 139.485 107.840 139.530 ;
        RECT 101.560 139.470 101.880 139.485 ;
        RECT 54.655 139.145 54.945 139.375 ;
        RECT 56.480 139.130 56.800 139.390 ;
        RECT 58.320 139.330 58.640 139.390 ;
        RECT 59.255 139.330 59.545 139.375 ;
        RECT 58.320 139.190 59.545 139.330 ;
        RECT 58.320 139.130 58.640 139.190 ;
        RECT 59.255 139.145 59.545 139.190 ;
        RECT 75.340 139.130 75.660 139.390 ;
        RECT 76.260 139.330 76.580 139.390 ;
        RECT 77.195 139.330 77.485 139.375 ;
        RECT 76.260 139.190 77.485 139.330 ;
        RECT 76.260 139.130 76.580 139.190 ;
        RECT 77.195 139.145 77.485 139.190 ;
        RECT 83.620 139.130 83.940 139.390 ;
        RECT 98.800 139.330 99.120 139.390 ;
        RECT 99.505 139.330 99.795 139.375 ;
        RECT 102.020 139.330 102.340 139.390 ;
        RECT 98.800 139.190 102.340 139.330 ;
        RECT 98.800 139.130 99.120 139.190 ;
        RECT 99.505 139.145 99.795 139.190 ;
        RECT 102.020 139.130 102.340 139.190 ;
        RECT 107.080 139.330 107.400 139.390 ;
        RECT 109.010 139.330 109.150 139.825 ;
        RECT 107.080 139.190 109.150 139.330 ;
        RECT 132.510 139.190 135.210 140.010 ;
        RECT 143.370 139.390 144.510 223.840 ;
        RECT 137.240 139.380 144.510 139.390 ;
        RECT 136.210 139.190 144.510 139.380 ;
        RECT 107.080 139.130 107.400 139.190 ;
        RECT 15.010 138.510 113.450 138.990 ;
        RECT 132.510 138.530 144.510 139.190 ;
        RECT 18.300 138.110 18.620 138.370 ;
        RECT 18.760 138.110 19.080 138.370 ;
        RECT 20.600 138.110 20.920 138.370 ;
        RECT 26.580 138.110 26.900 138.370 ;
        RECT 39.920 138.310 40.240 138.370 ;
        RECT 42.220 138.310 42.540 138.370 ;
        RECT 39.920 138.170 42.540 138.310 ;
        RECT 39.920 138.110 40.240 138.170 ;
        RECT 42.220 138.110 42.540 138.170 ;
        RECT 49.120 138.310 49.440 138.370 ;
        RECT 73.040 138.310 73.360 138.370 ;
        RECT 49.120 138.170 73.360 138.310 ;
        RECT 49.120 138.110 49.440 138.170 ;
        RECT 21.075 137.970 21.365 138.015 ;
        RECT 28.880 137.970 29.200 138.030 ;
        RECT 21.075 137.830 29.200 137.970 ;
        RECT 21.075 137.785 21.365 137.830 ;
        RECT 28.880 137.770 29.200 137.830 ;
        RECT 44.535 137.970 44.825 138.015 ;
        RECT 44.995 137.970 45.285 138.015 ;
        RECT 44.535 137.830 45.285 137.970 ;
        RECT 44.535 137.785 44.825 137.830 ;
        RECT 44.995 137.785 45.285 137.830 ;
        RECT 45.900 137.970 46.220 138.030 ;
        RECT 48.660 137.970 48.980 138.030 ;
        RECT 50.040 137.970 50.360 138.030 ;
        RECT 55.560 138.015 55.880 138.030 ;
        RECT 45.900 137.830 50.360 137.970 ;
        RECT 45.900 137.770 46.220 137.830 ;
        RECT 17.395 137.445 17.685 137.675 ;
        RECT 17.470 136.950 17.610 137.445 ;
        RECT 23.360 137.430 23.680 137.690 ;
        RECT 25.675 137.630 25.965 137.675 ;
        RECT 35.320 137.630 35.640 137.690 ;
        RECT 25.675 137.490 35.640 137.630 ;
        RECT 25.675 137.445 25.965 137.490 ;
        RECT 35.320 137.430 35.640 137.490 ;
        RECT 36.240 137.630 36.560 137.690 ;
        RECT 40.855 137.630 41.145 137.675 ;
        RECT 36.240 137.490 41.145 137.630 ;
        RECT 36.240 137.430 36.560 137.490 ;
        RECT 40.855 137.445 41.145 137.490 ;
        RECT 43.140 137.430 43.460 137.690 ;
        RECT 46.360 137.430 46.680 137.690 ;
        RECT 46.910 137.675 47.050 137.830 ;
        RECT 48.660 137.770 48.980 137.830 ;
        RECT 50.040 137.770 50.360 137.830 ;
        RECT 52.290 137.970 52.580 138.015 ;
        RECT 55.550 137.970 55.880 138.015 ;
        RECT 52.290 137.830 55.880 137.970 ;
        RECT 52.290 137.785 52.580 137.830 ;
        RECT 55.550 137.785 55.880 137.830 ;
        RECT 55.560 137.770 55.880 137.785 ;
        RECT 56.470 137.970 56.760 138.015 ;
        RECT 58.330 137.970 58.620 138.015 ;
        RECT 56.470 137.830 58.620 137.970 ;
        RECT 56.470 137.785 56.760 137.830 ;
        RECT 58.330 137.785 58.620 137.830 ;
        RECT 67.995 137.970 68.285 138.015 ;
        RECT 70.755 137.970 71.045 138.015 ;
        RECT 67.995 137.830 71.045 137.970 ;
        RECT 67.995 137.785 68.285 137.830 ;
        RECT 70.755 137.785 71.045 137.830 ;
        RECT 46.835 137.445 47.125 137.675 ;
        RECT 47.295 137.445 47.585 137.675 ;
        RECT 47.740 137.630 48.060 137.690 ;
        RECT 48.215 137.630 48.505 137.675 ;
        RECT 50.960 137.630 51.280 137.690 ;
        RECT 47.740 137.490 51.280 137.630 ;
        RECT 21.060 137.290 21.380 137.350 ;
        RECT 21.535 137.290 21.825 137.335 ;
        RECT 21.060 137.150 21.825 137.290 ;
        RECT 21.060 137.090 21.380 137.150 ;
        RECT 21.535 137.105 21.825 137.150 ;
        RECT 24.755 137.290 25.045 137.335 ;
        RECT 28.880 137.290 29.200 137.350 ;
        RECT 29.355 137.290 29.645 137.335 ;
        RECT 24.755 137.150 29.645 137.290 ;
        RECT 24.755 137.105 25.045 137.150 ;
        RECT 28.880 137.090 29.200 137.150 ;
        RECT 29.355 137.105 29.645 137.150 ;
        RECT 30.275 137.290 30.565 137.335 ;
        RECT 30.720 137.290 31.040 137.350 ;
        RECT 30.275 137.150 31.040 137.290 ;
        RECT 30.275 137.105 30.565 137.150 ;
        RECT 30.720 137.090 31.040 137.150 ;
        RECT 44.060 137.090 44.380 137.350 ;
        RECT 27.055 136.950 27.345 136.995 ;
        RECT 17.470 136.810 27.345 136.950 ;
        RECT 47.370 136.950 47.510 137.445 ;
        RECT 47.740 137.430 48.060 137.490 ;
        RECT 48.215 137.445 48.505 137.490 ;
        RECT 50.960 137.430 51.280 137.490 ;
        RECT 54.150 137.630 54.440 137.675 ;
        RECT 56.470 137.630 56.685 137.785 ;
        RECT 72.210 137.690 72.350 138.170 ;
        RECT 73.040 138.110 73.360 138.170 ;
        RECT 83.620 138.310 83.940 138.370 ;
        RECT 85.015 138.310 85.305 138.355 ;
        RECT 83.620 138.170 85.305 138.310 ;
        RECT 83.620 138.110 83.940 138.170 ;
        RECT 85.015 138.125 85.305 138.170 ;
        RECT 85.460 138.310 85.780 138.370 ;
        RECT 86.395 138.310 86.685 138.355 ;
        RECT 85.460 138.170 86.685 138.310 ;
        RECT 85.460 138.110 85.780 138.170 ;
        RECT 86.395 138.125 86.685 138.170 ;
        RECT 90.520 138.310 90.840 138.370 ;
        RECT 90.995 138.310 91.285 138.355 ;
        RECT 90.520 138.170 91.285 138.310 ;
        RECT 90.520 138.110 90.840 138.170 ;
        RECT 90.995 138.125 91.285 138.170 ;
        RECT 102.020 138.110 102.340 138.370 ;
        RECT 102.480 138.110 102.800 138.370 ;
        RECT 104.335 138.125 104.625 138.355 ;
        RECT 106.175 138.310 106.465 138.355 ;
        RECT 106.620 138.310 106.940 138.370 ;
        RECT 106.175 138.170 106.940 138.310 ;
        RECT 132.510 138.190 135.210 138.530 ;
        RECT 136.210 138.250 144.510 138.530 ;
        RECT 136.210 138.240 138.350 138.250 ;
        RECT 106.175 138.125 106.465 138.170 ;
        RECT 74.880 138.015 75.200 138.030 ;
        RECT 80.400 138.015 80.720 138.030 ;
        RECT 74.880 137.970 75.415 138.015 ;
        RECT 77.130 137.970 77.420 138.015 ;
        RECT 80.390 137.970 80.720 138.015 ;
        RECT 73.130 137.830 75.635 137.970 ;
        RECT 77.130 137.830 80.720 137.970 ;
        RECT 54.150 137.490 56.685 137.630 ;
        RECT 56.940 137.630 57.260 137.690 ;
        RECT 57.415 137.630 57.705 137.675 ;
        RECT 56.940 137.490 57.705 137.630 ;
        RECT 54.150 137.445 54.440 137.490 ;
        RECT 56.940 137.430 57.260 137.490 ;
        RECT 57.415 137.445 57.705 137.490 ;
        RECT 69.360 137.430 69.680 137.690 ;
        RECT 72.120 137.430 72.440 137.690 ;
        RECT 72.580 137.430 72.900 137.690 ;
        RECT 73.130 137.675 73.270 137.830 ;
        RECT 74.880 137.785 75.415 137.830 ;
        RECT 77.130 137.785 77.420 137.830 ;
        RECT 80.390 137.785 80.720 137.830 ;
        RECT 74.880 137.770 75.200 137.785 ;
        RECT 80.400 137.770 80.720 137.785 ;
        RECT 81.310 137.970 81.600 138.015 ;
        RECT 83.170 137.970 83.460 138.015 ;
        RECT 81.310 137.830 83.460 137.970 ;
        RECT 81.310 137.785 81.600 137.830 ;
        RECT 83.170 137.785 83.460 137.830 ;
        RECT 85.550 137.830 88.450 137.970 ;
        RECT 73.055 137.445 73.345 137.675 ;
        RECT 73.975 137.445 74.265 137.675 ;
        RECT 78.990 137.630 79.280 137.675 ;
        RECT 81.310 137.630 81.525 137.785 ;
        RECT 85.550 137.690 85.690 137.830 ;
        RECT 88.310 137.690 88.450 137.830 ;
        RECT 95.120 137.770 95.440 138.030 ;
        RECT 95.580 137.770 95.900 138.030 ;
        RECT 96.040 137.970 96.360 138.030 ;
        RECT 104.410 137.970 104.550 138.125 ;
        RECT 106.620 138.110 106.940 138.170 ;
        RECT 96.040 137.830 97.190 137.970 ;
        RECT 104.410 137.830 105.470 137.970 ;
        RECT 96.040 137.770 96.360 137.830 ;
        RECT 78.990 137.490 81.525 137.630 ;
        RECT 78.990 137.445 79.280 137.490 ;
        RECT 50.500 137.290 50.820 137.350 ;
        RECT 59.255 137.290 59.545 137.335 ;
        RECT 50.500 137.150 59.545 137.290 ;
        RECT 50.500 137.090 50.820 137.150 ;
        RECT 59.255 137.105 59.545 137.150 ;
        RECT 68.440 137.090 68.760 137.350 ;
        RECT 53.260 136.950 53.580 137.010 ;
        RECT 47.370 136.810 53.580 136.950 ;
        RECT 27.055 136.765 27.345 136.810 ;
        RECT 53.260 136.750 53.580 136.810 ;
        RECT 54.150 136.950 54.440 136.995 ;
        RECT 56.930 136.950 57.220 136.995 ;
        RECT 58.790 136.950 59.080 136.995 ;
        RECT 54.150 136.810 59.080 136.950 ;
        RECT 54.150 136.765 54.440 136.810 ;
        RECT 56.930 136.765 57.220 136.810 ;
        RECT 58.790 136.765 59.080 136.810 ;
        RECT 64.760 136.950 65.080 137.010 ;
        RECT 74.050 136.950 74.190 137.445 ;
        RECT 82.240 137.430 82.560 137.690 ;
        RECT 85.460 137.430 85.780 137.690 ;
        RECT 87.300 137.430 87.620 137.690 ;
        RECT 88.220 137.630 88.540 137.690 ;
        RECT 90.535 137.630 90.825 137.675 ;
        RECT 88.220 137.490 90.825 137.630 ;
        RECT 88.220 137.430 88.540 137.490 ;
        RECT 90.535 137.445 90.825 137.490 ;
        RECT 93.740 137.430 94.060 137.690 ;
        RECT 96.500 137.430 96.820 137.690 ;
        RECT 97.050 137.675 97.190 137.830 ;
        RECT 105.330 137.675 105.470 137.830 ;
        RECT 96.975 137.445 97.265 137.675 ;
        RECT 105.295 137.445 105.585 137.675 ;
        RECT 76.720 137.290 77.040 137.350 ;
        RECT 84.095 137.290 84.385 137.335 ;
        RECT 76.720 137.150 84.385 137.290 ;
        RECT 76.720 137.090 77.040 137.150 ;
        RECT 84.095 137.105 84.385 137.150 ;
        RECT 91.900 137.290 92.220 137.350 ;
        RECT 94.215 137.290 94.505 137.335 ;
        RECT 91.900 137.150 94.505 137.290 ;
        RECT 91.900 137.090 92.220 137.150 ;
        RECT 94.215 137.105 94.505 137.150 ;
        RECT 101.575 137.290 101.865 137.335 ;
        RECT 104.320 137.290 104.640 137.350 ;
        RECT 101.575 137.150 104.640 137.290 ;
        RECT 101.575 137.105 101.865 137.150 ;
        RECT 104.320 137.090 104.640 137.150 ;
        RECT 74.420 136.950 74.740 137.010 ;
        RECT 64.760 136.810 74.740 136.950 ;
        RECT 64.760 136.750 65.080 136.810 ;
        RECT 74.420 136.750 74.740 136.810 ;
        RECT 78.990 136.950 79.280 136.995 ;
        RECT 81.770 136.950 82.060 136.995 ;
        RECT 83.630 136.950 83.920 136.995 ;
        RECT 78.990 136.810 83.920 136.950 ;
        RECT 78.990 136.765 79.280 136.810 ;
        RECT 81.770 136.765 82.060 136.810 ;
        RECT 83.630 136.765 83.920 136.810 ;
        RECT 92.835 136.950 93.125 136.995 ;
        RECT 95.580 136.950 95.900 137.010 ;
        RECT 92.835 136.810 95.900 136.950 ;
        RECT 92.835 136.765 93.125 136.810 ;
        RECT 95.580 136.750 95.900 136.810 ;
        RECT 23.835 136.610 24.125 136.655 ;
        RECT 28.420 136.610 28.740 136.670 ;
        RECT 23.835 136.470 28.740 136.610 ;
        RECT 23.835 136.425 24.125 136.470 ;
        RECT 28.420 136.410 28.740 136.470 ;
        RECT 42.220 136.410 42.540 136.670 ;
        RECT 44.060 136.410 44.380 136.670 ;
        RECT 50.285 136.610 50.575 136.655 ;
        RECT 52.340 136.610 52.660 136.670 ;
        RECT 50.285 136.470 52.660 136.610 ;
        RECT 50.285 136.425 50.575 136.470 ;
        RECT 52.340 136.410 52.660 136.470 ;
        RECT 67.520 136.610 67.840 136.670 ;
        RECT 67.995 136.610 68.285 136.655 ;
        RECT 67.520 136.470 68.285 136.610 ;
        RECT 67.520 136.410 67.840 136.470 ;
        RECT 67.995 136.425 68.285 136.470 ;
        RECT 69.820 136.610 70.140 136.670 ;
        RECT 70.295 136.610 70.585 136.655 ;
        RECT 69.820 136.470 70.585 136.610 ;
        RECT 69.820 136.410 70.140 136.470 ;
        RECT 70.295 136.425 70.585 136.470 ;
        RECT 72.580 136.610 72.900 136.670 ;
        RECT 75.800 136.610 76.120 136.670 ;
        RECT 72.580 136.470 76.120 136.610 ;
        RECT 72.580 136.410 72.900 136.470 ;
        RECT 75.800 136.410 76.120 136.470 ;
        RECT 95.120 136.410 95.440 136.670 ;
        RECT 96.500 136.410 96.820 136.670 ;
        RECT 97.420 136.610 97.740 136.670 ;
        RECT 97.895 136.610 98.185 136.655 ;
        RECT 97.420 136.470 98.185 136.610 ;
        RECT 97.420 136.410 97.740 136.470 ;
        RECT 97.895 136.425 98.185 136.470 ;
        RECT 15.010 135.790 113.450 136.270 ;
        RECT 20.140 135.590 20.460 135.650 ;
        RECT 39.015 135.590 39.305 135.635 ;
        RECT 40.380 135.590 40.700 135.650 ;
        RECT 20.140 135.450 25.890 135.590 ;
        RECT 20.140 135.390 20.460 135.450 ;
        RECT 20.570 135.250 20.860 135.295 ;
        RECT 23.350 135.250 23.640 135.295 ;
        RECT 25.210 135.250 25.500 135.295 ;
        RECT 20.570 135.110 25.500 135.250 ;
        RECT 20.570 135.065 20.860 135.110 ;
        RECT 23.350 135.065 23.640 135.110 ;
        RECT 25.210 135.065 25.500 135.110 ;
        RECT 22.440 134.910 22.760 134.970 ;
        RECT 23.835 134.910 24.125 134.955 ;
        RECT 25.750 134.910 25.890 135.450 ;
        RECT 39.015 135.450 40.700 135.590 ;
        RECT 39.015 135.405 39.305 135.450 ;
        RECT 40.380 135.390 40.700 135.450 ;
        RECT 41.300 135.390 41.620 135.650 ;
        RECT 55.560 135.590 55.880 135.650 ;
        RECT 56.495 135.590 56.785 135.635 ;
        RECT 55.560 135.450 56.785 135.590 ;
        RECT 55.560 135.390 55.880 135.450 ;
        RECT 56.495 135.405 56.785 135.450 ;
        RECT 69.835 135.590 70.125 135.635 ;
        RECT 71.200 135.590 71.520 135.650 ;
        RECT 69.835 135.450 71.520 135.590 ;
        RECT 69.835 135.405 70.125 135.450 ;
        RECT 71.200 135.390 71.520 135.450 ;
        RECT 79.955 135.590 80.245 135.635 ;
        RECT 80.400 135.590 80.720 135.650 ;
        RECT 79.955 135.450 80.720 135.590 ;
        RECT 79.955 135.405 80.245 135.450 ;
        RECT 80.400 135.390 80.720 135.450 ;
        RECT 81.795 135.590 82.085 135.635 ;
        RECT 82.240 135.590 82.560 135.650 ;
        RECT 81.795 135.450 82.560 135.590 ;
        RECT 81.795 135.405 82.085 135.450 ;
        RECT 82.240 135.390 82.560 135.450 ;
        RECT 90.980 135.590 91.300 135.650 ;
        RECT 94.215 135.590 94.505 135.635 ;
        RECT 90.980 135.450 94.505 135.590 ;
        RECT 90.980 135.390 91.300 135.450 ;
        RECT 94.215 135.405 94.505 135.450 ;
        RECT 97.880 135.390 98.200 135.650 ;
        RECT 30.230 135.250 30.520 135.295 ;
        RECT 33.010 135.250 33.300 135.295 ;
        RECT 34.870 135.250 35.160 135.295 ;
        RECT 30.230 135.110 35.160 135.250 ;
        RECT 30.230 135.065 30.520 135.110 ;
        RECT 33.010 135.065 33.300 135.110 ;
        RECT 34.870 135.065 35.160 135.110 ;
        RECT 39.460 135.050 39.780 135.310 ;
        RECT 46.360 135.250 46.680 135.310 ;
        RECT 45.530 135.110 46.680 135.250 ;
        RECT 22.440 134.770 23.590 134.910 ;
        RECT 22.440 134.710 22.760 134.770 ;
        RECT 20.570 134.570 20.860 134.615 ;
        RECT 23.450 134.570 23.590 134.770 ;
        RECT 23.835 134.770 25.890 134.910 ;
        RECT 23.835 134.725 24.125 134.770 ;
        RECT 38.080 134.710 38.400 134.970 ;
        RECT 39.000 134.710 39.320 134.970 ;
        RECT 40.840 134.710 41.160 134.970 ;
        RECT 25.675 134.570 25.965 134.615 ;
        RECT 20.570 134.430 23.105 134.570 ;
        RECT 23.450 134.430 25.965 134.570 ;
        RECT 20.570 134.385 20.860 134.430 ;
        RECT 18.710 134.230 19.000 134.275 ;
        RECT 19.680 134.230 20.000 134.290 ;
        RECT 22.890 134.275 23.105 134.430 ;
        RECT 25.675 134.385 25.965 134.430 ;
        RECT 30.230 134.570 30.520 134.615 ;
        RECT 33.495 134.570 33.785 134.615 ;
        RECT 34.860 134.570 35.180 134.630 ;
        RECT 30.230 134.430 32.765 134.570 ;
        RECT 30.230 134.385 30.520 134.430 ;
        RECT 28.420 134.275 28.740 134.290 ;
        RECT 32.550 134.275 32.765 134.430 ;
        RECT 33.495 134.430 35.180 134.570 ;
        RECT 33.495 134.385 33.785 134.430 ;
        RECT 34.860 134.370 35.180 134.430 ;
        RECT 35.335 134.570 35.625 134.615 ;
        RECT 36.240 134.570 36.560 134.630 ;
        RECT 35.335 134.430 36.560 134.570 ;
        RECT 35.335 134.385 35.625 134.430 ;
        RECT 36.240 134.370 36.560 134.430 ;
        RECT 37.635 134.570 37.925 134.615 ;
        RECT 39.090 134.570 39.230 134.710 ;
        RECT 37.635 134.430 39.230 134.570 ;
        RECT 39.920 134.570 40.240 134.630 ;
        RECT 45.530 134.615 45.670 135.110 ;
        RECT 46.360 135.050 46.680 135.110 ;
        RECT 50.040 135.050 50.360 135.310 ;
        RECT 50.960 135.250 51.280 135.310 ;
        RECT 64.760 135.250 65.080 135.310 ;
        RECT 85.460 135.250 85.780 135.310 ;
        RECT 50.960 135.110 65.080 135.250 ;
        RECT 50.960 135.050 51.280 135.110 ;
        RECT 64.760 135.050 65.080 135.110 ;
        RECT 80.490 135.110 85.780 135.250 ;
        RECT 50.130 134.910 50.270 135.050 ;
        RECT 49.670 134.770 50.270 134.910 ;
        RECT 53.260 134.910 53.580 134.970 ;
        RECT 54.195 134.910 54.485 134.955 ;
        RECT 53.260 134.770 54.485 134.910 ;
        RECT 40.395 134.570 40.685 134.615 ;
        RECT 39.920 134.430 40.685 134.570 ;
        RECT 37.635 134.385 37.925 134.430 ;
        RECT 39.920 134.370 40.240 134.430 ;
        RECT 40.395 134.385 40.685 134.430 ;
        RECT 45.455 134.385 45.745 134.615 ;
        RECT 21.970 134.230 22.260 134.275 ;
        RECT 18.710 134.090 22.260 134.230 ;
        RECT 18.710 134.045 19.000 134.090 ;
        RECT 19.680 134.030 20.000 134.090 ;
        RECT 21.970 134.045 22.260 134.090 ;
        RECT 22.890 134.230 23.180 134.275 ;
        RECT 24.750 134.230 25.040 134.275 ;
        RECT 22.890 134.090 25.040 134.230 ;
        RECT 22.890 134.045 23.180 134.090 ;
        RECT 24.750 134.045 25.040 134.090 ;
        RECT 28.370 134.230 28.740 134.275 ;
        RECT 31.630 134.230 31.920 134.275 ;
        RECT 28.370 134.090 31.920 134.230 ;
        RECT 28.370 134.045 28.740 134.090 ;
        RECT 31.630 134.045 31.920 134.090 ;
        RECT 32.550 134.230 32.840 134.275 ;
        RECT 34.410 134.230 34.700 134.275 ;
        RECT 32.550 134.090 34.700 134.230 ;
        RECT 32.550 134.045 32.840 134.090 ;
        RECT 34.410 134.045 34.700 134.090 ;
        RECT 39.015 134.045 39.305 134.275 ;
        RECT 41.775 134.230 42.065 134.275 ;
        RECT 44.075 134.230 44.365 134.275 ;
        RECT 41.775 134.090 44.365 134.230 ;
        RECT 45.530 134.230 45.670 134.385 ;
        RECT 45.900 134.370 46.220 134.630 ;
        RECT 46.360 134.370 46.680 134.630 ;
        RECT 46.820 134.570 47.140 134.630 ;
        RECT 49.670 134.615 49.810 134.770 ;
        RECT 53.260 134.710 53.580 134.770 ;
        RECT 54.195 134.725 54.485 134.770 ;
        RECT 55.100 134.710 55.420 134.970 ;
        RECT 67.995 134.910 68.285 134.955 ;
        RECT 71.200 134.910 71.520 134.970 ;
        RECT 67.995 134.770 71.520 134.910 ;
        RECT 67.995 134.725 68.285 134.770 ;
        RECT 71.200 134.710 71.520 134.770 ;
        RECT 47.295 134.570 47.585 134.615 ;
        RECT 48.905 134.570 49.195 134.615 ;
        RECT 46.820 134.430 47.585 134.570 ;
        RECT 46.820 134.370 47.140 134.430 ;
        RECT 47.295 134.385 47.585 134.430 ;
        RECT 47.830 134.430 49.195 134.570 ;
        RECT 47.830 134.230 47.970 134.430 ;
        RECT 48.905 134.385 49.195 134.430 ;
        RECT 49.595 134.385 49.885 134.615 ;
        RECT 50.055 134.385 50.345 134.615 ;
        RECT 45.530 134.090 47.970 134.230 ;
        RECT 50.130 134.230 50.270 134.385 ;
        RECT 50.960 134.370 51.280 134.630 ;
        RECT 51.420 134.570 51.740 134.630 ;
        RECT 56.955 134.570 57.245 134.615 ;
        RECT 57.415 134.570 57.705 134.615 ;
        RECT 51.420 134.430 54.410 134.570 ;
        RECT 51.420 134.370 51.740 134.430 ;
        RECT 52.340 134.230 52.660 134.290 ;
        RECT 53.735 134.230 54.025 134.275 ;
        RECT 50.130 134.090 54.025 134.230 ;
        RECT 54.270 134.230 54.410 134.430 ;
        RECT 56.955 134.430 57.705 134.570 ;
        RECT 56.955 134.385 57.245 134.430 ;
        RECT 57.415 134.385 57.705 134.430 ;
        RECT 57.030 134.230 57.170 134.385 ;
        RECT 64.300 134.370 64.620 134.630 ;
        RECT 68.440 134.570 68.760 134.630 ;
        RECT 68.915 134.570 69.205 134.615 ;
        RECT 68.440 134.430 69.205 134.570 ;
        RECT 68.440 134.370 68.760 134.430 ;
        RECT 68.915 134.385 69.205 134.430 ;
        RECT 79.020 134.370 79.340 134.630 ;
        RECT 80.490 134.615 80.630 135.110 ;
        RECT 85.460 135.050 85.780 135.110 ;
        RECT 80.415 134.385 80.705 134.615 ;
        RECT 80.875 134.385 81.165 134.615 ;
        RECT 54.270 134.090 57.170 134.230 ;
        RECT 62.000 134.230 62.320 134.290 ;
        RECT 63.395 134.230 63.685 134.275 ;
        RECT 62.000 134.090 63.685 134.230 ;
        RECT 41.775 134.045 42.065 134.090 ;
        RECT 44.075 134.045 44.365 134.090 ;
        RECT 28.420 134.030 28.740 134.045 ;
        RECT 16.705 133.890 16.995 133.935 ;
        RECT 20.600 133.890 20.920 133.950 ;
        RECT 16.705 133.750 20.920 133.890 ;
        RECT 16.705 133.705 16.995 133.750 ;
        RECT 20.600 133.690 20.920 133.750 ;
        RECT 26.365 133.890 26.655 133.935 ;
        RECT 28.880 133.890 29.200 133.950 ;
        RECT 26.365 133.750 29.200 133.890 ;
        RECT 26.365 133.705 26.655 133.750 ;
        RECT 28.880 133.690 29.200 133.750 ;
        RECT 36.700 133.690 37.020 133.950 ;
        RECT 39.090 133.890 39.230 134.045 ;
        RECT 52.340 134.030 52.660 134.090 ;
        RECT 53.735 134.045 54.025 134.090 ;
        RECT 62.000 134.030 62.320 134.090 ;
        RECT 63.395 134.045 63.685 134.090 ;
        RECT 67.980 134.230 68.300 134.290 ;
        RECT 70.755 134.230 71.045 134.275 ;
        RECT 73.040 134.230 73.360 134.290 ;
        RECT 67.980 134.090 73.360 134.230 ;
        RECT 67.980 134.030 68.300 134.090 ;
        RECT 70.755 134.045 71.045 134.090 ;
        RECT 73.040 134.030 73.360 134.090 ;
        RECT 47.755 133.890 48.045 133.935 ;
        RECT 39.090 133.750 48.045 133.890 ;
        RECT 47.755 133.705 48.045 133.750 ;
        RECT 49.120 133.890 49.440 133.950 ;
        RECT 51.895 133.890 52.185 133.935 ;
        RECT 49.120 133.750 52.185 133.890 ;
        RECT 49.120 133.690 49.440 133.750 ;
        RECT 51.895 133.705 52.185 133.750 ;
        RECT 57.400 133.890 57.720 133.950 ;
        RECT 57.875 133.890 58.165 133.935 ;
        RECT 57.400 133.750 58.165 133.890 ;
        RECT 57.400 133.690 57.720 133.750 ;
        RECT 57.875 133.705 58.165 133.750 ;
        RECT 76.260 133.890 76.580 133.950 ;
        RECT 80.950 133.890 81.090 134.385 ;
        RECT 98.800 134.370 99.120 134.630 ;
        RECT 99.735 134.570 100.025 134.615 ;
        RECT 104.780 134.570 105.100 134.630 ;
        RECT 99.735 134.430 105.100 134.570 ;
        RECT 135.660 134.480 136.800 134.510 ;
        RECT 99.735 134.385 100.025 134.430 ;
        RECT 104.780 134.370 105.100 134.430 ;
        RECT 85.000 134.230 85.320 134.290 ;
        RECT 87.775 134.230 88.065 134.275 ;
        RECT 85.000 134.090 88.065 134.230 ;
        RECT 85.000 134.030 85.320 134.090 ;
        RECT 87.775 134.045 88.065 134.090 ;
        RECT 76.260 133.750 81.090 133.890 ;
        RECT 76.260 133.690 76.580 133.750 ;
        RECT 15.010 133.070 113.450 133.550 ;
        RECT 135.590 133.400 136.850 134.480 ;
        RECT 20.155 132.870 20.445 132.915 ;
        RECT 20.600 132.870 20.920 132.930 ;
        RECT 20.155 132.730 20.920 132.870 ;
        RECT 20.155 132.685 20.445 132.730 ;
        RECT 20.600 132.670 20.920 132.730 ;
        RECT 21.980 132.870 22.300 132.930 ;
        RECT 35.320 132.870 35.640 132.930 ;
        RECT 21.980 132.730 26.810 132.870 ;
        RECT 21.980 132.670 22.300 132.730 ;
        RECT 24.300 132.530 24.590 132.575 ;
        RECT 26.160 132.530 26.450 132.575 ;
        RECT 24.300 132.390 26.450 132.530 ;
        RECT 26.670 132.530 26.810 132.730 ;
        RECT 35.320 132.730 43.370 132.870 ;
        RECT 35.320 132.670 35.640 132.730 ;
        RECT 27.080 132.530 27.370 132.575 ;
        RECT 30.340 132.530 30.630 132.575 ;
        RECT 26.670 132.390 30.630 132.530 ;
        RECT 24.300 132.345 24.590 132.390 ;
        RECT 26.160 132.345 26.450 132.390 ;
        RECT 27.080 132.345 27.370 132.390 ;
        RECT 30.340 132.345 30.630 132.390 ;
        RECT 41.775 132.530 42.065 132.575 ;
        RECT 42.680 132.530 43.000 132.590 ;
        RECT 41.775 132.390 43.000 132.530 ;
        RECT 43.230 132.530 43.370 132.730 ;
        RECT 44.060 132.670 44.380 132.930 ;
        RECT 62.000 132.870 62.320 132.930 ;
        RECT 50.590 132.730 62.320 132.870 ;
        RECT 50.590 132.530 50.730 132.730 ;
        RECT 62.000 132.670 62.320 132.730 ;
        RECT 67.520 132.670 67.840 132.930 ;
        RECT 70.740 132.670 71.060 132.930 ;
        RECT 73.040 132.870 73.360 132.930 ;
        RECT 76.720 132.870 77.040 132.930 ;
        RECT 73.040 132.730 77.040 132.870 ;
        RECT 73.040 132.670 73.360 132.730 ;
        RECT 76.720 132.670 77.040 132.730 ;
        RECT 94.660 132.870 94.980 132.930 ;
        RECT 95.135 132.870 95.425 132.915 ;
        RECT 94.660 132.730 95.425 132.870 ;
        RECT 94.660 132.670 94.980 132.730 ;
        RECT 95.135 132.685 95.425 132.730 ;
        RECT 96.960 132.870 97.280 132.930 ;
        RECT 97.895 132.870 98.185 132.915 ;
        RECT 96.960 132.730 98.185 132.870 ;
        RECT 96.960 132.670 97.280 132.730 ;
        RECT 97.895 132.685 98.185 132.730 ;
        RECT 57.400 132.575 57.720 132.590 ;
        RECT 43.230 132.390 50.730 132.530 ;
        RECT 51.440 132.530 51.730 132.575 ;
        RECT 53.300 132.530 53.590 132.575 ;
        RECT 51.440 132.390 53.590 132.530 ;
        RECT 41.775 132.345 42.065 132.390 ;
        RECT 20.140 132.190 20.460 132.250 ;
        RECT 20.615 132.190 20.905 132.235 ;
        RECT 20.140 132.050 20.905 132.190 ;
        RECT 20.140 131.990 20.460 132.050 ;
        RECT 20.615 132.005 20.905 132.050 ;
        RECT 22.440 132.190 22.760 132.250 ;
        RECT 23.375 132.190 23.665 132.235 ;
        RECT 24.740 132.190 25.060 132.250 ;
        RECT 22.440 132.050 25.060 132.190 ;
        RECT 22.440 131.990 22.760 132.050 ;
        RECT 23.375 132.005 23.665 132.050 ;
        RECT 24.740 131.990 25.060 132.050 ;
        RECT 25.200 131.990 25.520 132.250 ;
        RECT 26.235 132.190 26.450 132.345 ;
        RECT 42.680 132.330 43.000 132.390 ;
        RECT 51.440 132.345 51.730 132.390 ;
        RECT 53.300 132.345 53.590 132.390 ;
        RECT 54.220 132.530 54.510 132.575 ;
        RECT 57.400 132.530 57.770 132.575 ;
        RECT 75.340 132.530 75.660 132.590 ;
        RECT 54.220 132.390 57.770 132.530 ;
        RECT 54.220 132.345 54.510 132.390 ;
        RECT 57.400 132.345 57.770 132.390 ;
        RECT 73.130 132.390 75.660 132.530 ;
        RECT 28.480 132.190 28.770 132.235 ;
        RECT 33.035 132.190 33.325 132.235 ;
        RECT 36.240 132.190 36.560 132.250 ;
        RECT 26.235 132.050 28.770 132.190 ;
        RECT 28.480 132.005 28.770 132.050 ;
        RECT 28.970 132.050 36.560 132.190 ;
        RECT 19.695 131.850 19.985 131.895 ;
        RECT 21.060 131.850 21.380 131.910 ;
        RECT 19.695 131.710 21.380 131.850 ;
        RECT 24.830 131.850 24.970 131.990 ;
        RECT 28.970 131.850 29.110 132.050 ;
        RECT 33.035 132.005 33.325 132.050 ;
        RECT 36.240 131.990 36.560 132.050 ;
        RECT 43.155 132.005 43.445 132.235 ;
        RECT 45.455 132.005 45.745 132.235 ;
        RECT 24.830 131.710 29.110 131.850 ;
        RECT 40.840 131.850 41.160 131.910 ;
        RECT 42.235 131.850 42.525 131.895 ;
        RECT 40.840 131.710 42.525 131.850 ;
        RECT 19.695 131.665 19.985 131.710 ;
        RECT 21.060 131.650 21.380 131.710 ;
        RECT 40.840 131.650 41.160 131.710 ;
        RECT 42.235 131.665 42.525 131.710 ;
        RECT 42.680 131.850 43.000 131.910 ;
        RECT 43.230 131.850 43.370 132.005 ;
        RECT 45.530 131.850 45.670 132.005 ;
        RECT 49.120 131.990 49.440 132.250 ;
        RECT 52.355 132.190 52.645 132.235 ;
        RECT 50.130 132.050 52.645 132.190 ;
        RECT 53.375 132.190 53.590 132.345 ;
        RECT 57.400 132.330 57.720 132.345 ;
        RECT 55.620 132.190 55.910 132.235 ;
        RECT 53.375 132.050 55.910 132.190 ;
        RECT 42.680 131.710 45.670 131.850 ;
        RECT 42.680 131.650 43.000 131.710 ;
        RECT 46.375 131.665 46.665 131.895 ;
        RECT 23.840 131.510 24.130 131.555 ;
        RECT 25.700 131.510 25.990 131.555 ;
        RECT 28.480 131.510 28.770 131.555 ;
        RECT 23.840 131.370 28.770 131.510 ;
        RECT 23.840 131.325 24.130 131.370 ;
        RECT 25.700 131.325 25.990 131.370 ;
        RECT 28.480 131.325 28.770 131.370 ;
        RECT 29.800 131.510 30.120 131.570 ;
        RECT 41.760 131.510 42.080 131.570 ;
        RECT 44.535 131.510 44.825 131.555 ;
        RECT 29.800 131.370 33.250 131.510 ;
        RECT 29.800 131.310 30.120 131.370 ;
        RECT 22.455 131.170 22.745 131.215 ;
        RECT 27.040 131.170 27.360 131.230 ;
        RECT 22.455 131.030 27.360 131.170 ;
        RECT 22.455 130.985 22.745 131.030 ;
        RECT 27.040 130.970 27.360 131.030 ;
        RECT 31.640 131.170 31.960 131.230 ;
        RECT 32.345 131.170 32.635 131.215 ;
        RECT 31.640 131.030 32.635 131.170 ;
        RECT 33.110 131.170 33.250 131.370 ;
        RECT 41.760 131.370 44.825 131.510 ;
        RECT 41.760 131.310 42.080 131.370 ;
        RECT 44.535 131.325 44.825 131.370 ;
        RECT 46.450 131.170 46.590 131.665 ;
        RECT 50.130 131.555 50.270 132.050 ;
        RECT 52.355 132.005 52.645 132.050 ;
        RECT 55.620 132.005 55.910 132.050 ;
        RECT 62.015 132.190 62.305 132.235 ;
        RECT 63.380 132.190 63.700 132.250 ;
        RECT 62.015 132.050 63.700 132.190 ;
        RECT 62.015 132.005 62.305 132.050 ;
        RECT 63.380 131.990 63.700 132.050 ;
        RECT 64.760 132.190 65.080 132.250 ;
        RECT 65.235 132.190 65.525 132.235 ;
        RECT 64.760 132.050 65.525 132.190 ;
        RECT 64.760 131.990 65.080 132.050 ;
        RECT 65.235 132.005 65.525 132.050 ;
        RECT 68.440 132.190 68.760 132.250 ;
        RECT 68.440 132.050 70.970 132.190 ;
        RECT 68.440 131.990 68.760 132.050 ;
        RECT 50.500 131.650 50.820 131.910 ;
        RECT 51.420 131.850 51.740 131.910 ;
        RECT 60.635 131.850 60.925 131.895 ;
        RECT 51.420 131.710 60.925 131.850 ;
        RECT 51.420 131.650 51.740 131.710 ;
        RECT 60.635 131.665 60.925 131.710 ;
        RECT 66.140 131.650 66.460 131.910 ;
        RECT 69.375 131.850 69.665 131.895 ;
        RECT 70.280 131.850 70.600 131.910 ;
        RECT 69.375 131.710 70.600 131.850 ;
        RECT 70.830 131.850 70.970 132.050 ;
        RECT 72.120 131.990 72.440 132.250 ;
        RECT 72.580 131.990 72.900 132.250 ;
        RECT 73.130 132.235 73.270 132.390 ;
        RECT 75.340 132.330 75.660 132.390 ;
        RECT 73.055 132.005 73.345 132.235 ;
        RECT 73.975 132.190 74.265 132.235 ;
        RECT 74.420 132.190 74.740 132.250 ;
        RECT 73.975 132.050 74.740 132.190 ;
        RECT 73.975 132.005 74.265 132.050 ;
        RECT 74.420 131.990 74.740 132.050 ;
        RECT 75.800 131.990 76.120 132.250 ;
        RECT 76.810 132.235 76.950 132.670 ;
        RECT 85.870 132.530 86.160 132.575 ;
        RECT 87.300 132.530 87.620 132.590 ;
        RECT 89.130 132.530 89.420 132.575 ;
        RECT 85.870 132.390 89.420 132.530 ;
        RECT 85.870 132.345 86.160 132.390 ;
        RECT 87.300 132.330 87.620 132.390 ;
        RECT 89.130 132.345 89.420 132.390 ;
        RECT 90.050 132.530 90.340 132.575 ;
        RECT 91.910 132.530 92.200 132.575 ;
        RECT 90.050 132.390 92.200 132.530 ;
        RECT 90.050 132.345 90.340 132.390 ;
        RECT 91.910 132.345 92.200 132.390 ;
        RECT 101.115 132.530 101.405 132.575 ;
        RECT 104.270 132.530 104.560 132.575 ;
        RECT 107.530 132.530 107.820 132.575 ;
        RECT 101.115 132.390 107.820 132.530 ;
        RECT 101.115 132.345 101.405 132.390 ;
        RECT 104.270 132.345 104.560 132.390 ;
        RECT 107.530 132.345 107.820 132.390 ;
        RECT 108.450 132.530 108.740 132.575 ;
        RECT 110.310 132.530 110.600 132.575 ;
        RECT 108.450 132.390 110.600 132.530 ;
        RECT 108.450 132.345 108.740 132.390 ;
        RECT 110.310 132.345 110.600 132.390 ;
        RECT 76.735 132.005 77.025 132.235 ;
        RECT 80.415 132.005 80.705 132.235 ;
        RECT 80.490 131.850 80.630 132.005 ;
        RECT 80.860 131.990 81.180 132.250 ;
        RECT 87.730 132.190 88.020 132.235 ;
        RECT 90.050 132.190 90.265 132.345 ;
        RECT 87.730 132.050 90.265 132.190 ;
        RECT 87.730 132.005 88.020 132.050 ;
        RECT 90.980 131.990 91.300 132.250 ;
        RECT 96.055 132.190 96.345 132.235 ;
        RECT 98.800 132.190 99.120 132.250 ;
        RECT 96.055 132.050 99.120 132.190 ;
        RECT 96.055 132.005 96.345 132.050 ;
        RECT 98.800 131.990 99.120 132.050 ;
        RECT 100.640 131.990 100.960 132.250 ;
        RECT 106.130 132.190 106.420 132.235 ;
        RECT 108.450 132.190 108.665 132.345 ;
        RECT 106.130 132.050 108.665 132.190 ;
        RECT 106.130 132.005 106.420 132.050 ;
        RECT 70.830 131.710 80.630 131.850 ;
        RECT 86.840 131.850 87.160 131.910 ;
        RECT 92.835 131.850 93.125 131.895 ;
        RECT 86.840 131.710 93.125 131.850 ;
        RECT 69.375 131.665 69.665 131.710 ;
        RECT 70.280 131.650 70.600 131.710 ;
        RECT 86.840 131.650 87.160 131.710 ;
        RECT 92.835 131.665 93.125 131.710 ;
        RECT 96.960 131.650 97.280 131.910 ;
        RECT 99.720 131.850 100.040 131.910 ;
        RECT 102.265 131.850 102.555 131.895 ;
        RECT 99.720 131.710 102.555 131.850 ;
        RECT 99.720 131.650 100.040 131.710 ;
        RECT 102.265 131.665 102.555 131.710 ;
        RECT 109.395 131.850 109.685 131.895 ;
        RECT 109.840 131.850 110.160 131.910 ;
        RECT 109.395 131.710 110.160 131.850 ;
        RECT 109.395 131.665 109.685 131.710 ;
        RECT 109.840 131.650 110.160 131.710 ;
        RECT 111.235 131.850 111.525 131.895 ;
        RECT 111.680 131.850 112.000 131.910 ;
        RECT 111.235 131.710 112.000 131.850 ;
        RECT 111.235 131.665 111.525 131.710 ;
        RECT 111.680 131.650 112.000 131.710 ;
        RECT 50.055 131.325 50.345 131.555 ;
        RECT 50.980 131.510 51.270 131.555 ;
        RECT 52.840 131.510 53.130 131.555 ;
        RECT 55.620 131.510 55.910 131.555 ;
        RECT 50.980 131.370 55.910 131.510 ;
        RECT 50.980 131.325 51.270 131.370 ;
        RECT 52.840 131.325 53.130 131.370 ;
        RECT 55.620 131.325 55.910 131.370 ;
        RECT 57.860 131.510 58.180 131.570 ;
        RECT 65.680 131.510 66.000 131.570 ;
        RECT 57.860 131.370 66.000 131.510 ;
        RECT 57.860 131.310 58.180 131.370 ;
        RECT 65.680 131.310 66.000 131.370 ;
        RECT 73.960 131.510 74.280 131.570 ;
        RECT 79.495 131.510 79.785 131.555 ;
        RECT 73.960 131.370 79.785 131.510 ;
        RECT 73.960 131.310 74.280 131.370 ;
        RECT 79.495 131.325 79.785 131.370 ;
        RECT 87.730 131.510 88.020 131.555 ;
        RECT 90.510 131.510 90.800 131.555 ;
        RECT 92.370 131.510 92.660 131.555 ;
        RECT 87.730 131.370 92.660 131.510 ;
        RECT 87.730 131.325 88.020 131.370 ;
        RECT 90.510 131.325 90.800 131.370 ;
        RECT 92.370 131.325 92.660 131.370 ;
        RECT 106.130 131.510 106.420 131.555 ;
        RECT 108.910 131.510 109.200 131.555 ;
        RECT 110.770 131.510 111.060 131.555 ;
        RECT 106.130 131.370 111.060 131.510 ;
        RECT 106.130 131.325 106.420 131.370 ;
        RECT 108.910 131.325 109.200 131.370 ;
        RECT 110.770 131.325 111.060 131.370 ;
        RECT 33.110 131.030 46.590 131.170 ;
        RECT 53.260 131.170 53.580 131.230 ;
        RECT 55.100 131.170 55.420 131.230 ;
        RECT 59.485 131.170 59.775 131.215 ;
        RECT 53.260 131.030 59.775 131.170 ;
        RECT 31.640 130.970 31.960 131.030 ;
        RECT 32.345 130.985 32.635 131.030 ;
        RECT 53.260 130.970 53.580 131.030 ;
        RECT 55.100 130.970 55.420 131.030 ;
        RECT 59.485 130.985 59.775 131.030 ;
        RECT 63.380 131.170 63.700 131.230 ;
        RECT 64.315 131.170 64.605 131.215 ;
        RECT 63.380 131.030 64.605 131.170 ;
        RECT 63.380 130.970 63.700 131.030 ;
        RECT 64.315 130.985 64.605 131.030 ;
        RECT 74.880 130.970 75.200 131.230 ;
        RECT 83.865 131.170 84.155 131.215 ;
        RECT 88.680 131.170 89.000 131.230 ;
        RECT 83.865 131.030 89.000 131.170 ;
        RECT 83.865 130.985 84.155 131.030 ;
        RECT 88.680 130.970 89.000 131.030 ;
        RECT 15.010 130.350 113.450 130.830 ;
        RECT 16.705 130.150 16.995 130.195 ;
        RECT 20.140 130.150 20.460 130.210 ;
        RECT 16.705 130.010 26.350 130.150 ;
        RECT 16.705 129.965 16.995 130.010 ;
        RECT 20.140 129.950 20.460 130.010 ;
        RECT 20.570 129.810 20.860 129.855 ;
        RECT 23.350 129.810 23.640 129.855 ;
        RECT 25.210 129.810 25.500 129.855 ;
        RECT 20.570 129.670 25.500 129.810 ;
        RECT 20.570 129.625 20.860 129.670 ;
        RECT 23.350 129.625 23.640 129.670 ;
        RECT 25.210 129.625 25.500 129.670 ;
        RECT 24.740 129.470 25.060 129.530 ;
        RECT 25.675 129.470 25.965 129.515 ;
        RECT 24.740 129.330 25.965 129.470 ;
        RECT 26.210 129.470 26.350 130.010 ;
        RECT 29.340 129.950 29.660 130.210 ;
        RECT 34.860 130.150 35.180 130.210 ;
        RECT 36.255 130.150 36.545 130.195 ;
        RECT 34.860 130.010 36.545 130.150 ;
        RECT 34.860 129.950 35.180 130.010 ;
        RECT 36.255 129.965 36.545 130.010 ;
        RECT 41.760 130.150 42.080 130.210 ;
        RECT 42.680 130.150 43.000 130.210 ;
        RECT 41.760 130.010 43.000 130.150 ;
        RECT 41.760 129.950 42.080 130.010 ;
        RECT 42.680 129.950 43.000 130.010 ;
        RECT 50.500 130.150 50.820 130.210 ;
        RECT 50.975 130.150 51.265 130.195 ;
        RECT 50.500 130.010 51.265 130.150 ;
        RECT 50.500 129.950 50.820 130.010 ;
        RECT 50.975 129.965 51.265 130.010 ;
        RECT 72.595 130.150 72.885 130.195 ;
        RECT 75.800 130.150 76.120 130.210 ;
        RECT 72.595 130.010 76.120 130.150 ;
        RECT 72.595 129.965 72.885 130.010 ;
        RECT 75.800 129.950 76.120 130.010 ;
        RECT 89.600 130.150 89.920 130.210 ;
        RECT 90.075 130.150 90.365 130.195 ;
        RECT 89.600 130.010 90.365 130.150 ;
        RECT 89.600 129.950 89.920 130.010 ;
        RECT 90.075 129.965 90.365 130.010 ;
        RECT 90.980 130.150 91.300 130.210 ;
        RECT 91.455 130.150 91.745 130.195 ;
        RECT 90.980 130.010 91.745 130.150 ;
        RECT 90.980 129.950 91.300 130.010 ;
        RECT 91.455 129.965 91.745 130.010 ;
        RECT 95.120 129.950 95.440 130.210 ;
        RECT 96.500 129.950 96.820 130.210 ;
        RECT 100.180 130.150 100.500 130.210 ;
        RECT 108.935 130.150 109.225 130.195 ;
        RECT 109.840 130.150 110.160 130.210 ;
        RECT 100.180 130.010 101.790 130.150 ;
        RECT 100.180 129.950 100.500 130.010 ;
        RECT 30.720 129.810 31.040 129.870 ;
        RECT 55.560 129.810 55.880 129.870 ;
        RECT 62.000 129.810 62.320 129.870 ;
        RECT 73.520 129.810 73.810 129.855 ;
        RECT 75.380 129.810 75.670 129.855 ;
        RECT 78.160 129.810 78.450 129.855 ;
        RECT 88.680 129.810 89.000 129.870 ;
        RECT 96.960 129.810 97.280 129.870 ;
        RECT 30.720 129.670 32.790 129.810 ;
        RECT 30.720 129.610 31.040 129.670 ;
        RECT 32.650 129.515 32.790 129.670 ;
        RECT 54.270 129.670 58.090 129.810 ;
        RECT 31.195 129.470 31.485 129.515 ;
        RECT 26.210 129.330 31.485 129.470 ;
        RECT 24.740 129.270 25.060 129.330 ;
        RECT 25.675 129.285 25.965 129.330 ;
        RECT 31.195 129.285 31.485 129.330 ;
        RECT 32.575 129.470 32.865 129.515 ;
        RECT 40.855 129.470 41.145 129.515 ;
        RECT 51.420 129.470 51.740 129.530 ;
        RECT 54.270 129.515 54.410 129.670 ;
        RECT 55.560 129.610 55.880 129.670 ;
        RECT 57.950 129.515 58.090 129.670 ;
        RECT 62.000 129.670 72.810 129.810 ;
        RECT 62.000 129.610 62.320 129.670 ;
        RECT 32.575 129.330 51.740 129.470 ;
        RECT 32.575 129.285 32.865 129.330 ;
        RECT 40.855 129.285 41.145 129.330 ;
        RECT 51.420 129.270 51.740 129.330 ;
        RECT 54.195 129.285 54.485 129.515 ;
        RECT 57.875 129.285 58.165 129.515 ;
        RECT 68.440 129.470 68.760 129.530 ;
        RECT 63.010 129.330 68.760 129.470 ;
        RECT 20.570 129.130 20.860 129.175 ;
        RECT 23.835 129.130 24.125 129.175 ;
        RECT 20.570 128.990 23.105 129.130 ;
        RECT 20.570 128.945 20.860 128.990 ;
        RECT 18.710 128.790 19.000 128.835 ;
        RECT 21.060 128.790 21.380 128.850 ;
        RECT 22.890 128.835 23.105 128.990 ;
        RECT 23.835 128.990 26.350 129.130 ;
        RECT 23.835 128.945 24.125 128.990 ;
        RECT 21.970 128.790 22.260 128.835 ;
        RECT 18.710 128.650 22.260 128.790 ;
        RECT 18.710 128.605 19.000 128.650 ;
        RECT 21.060 128.590 21.380 128.650 ;
        RECT 21.970 128.605 22.260 128.650 ;
        RECT 22.890 128.790 23.180 128.835 ;
        RECT 24.750 128.790 25.040 128.835 ;
        RECT 22.890 128.650 25.040 128.790 ;
        RECT 22.890 128.605 23.180 128.650 ;
        RECT 24.750 128.605 25.040 128.650 ;
        RECT 26.210 128.495 26.350 128.990 ;
        RECT 27.040 128.930 27.360 129.190 ;
        RECT 27.960 128.930 28.280 129.190 ;
        RECT 30.275 129.130 30.565 129.175 ;
        RECT 34.860 129.130 35.180 129.190 ;
        RECT 30.275 128.990 35.180 129.130 ;
        RECT 30.275 128.945 30.565 128.990 ;
        RECT 34.860 128.930 35.180 128.990 ;
        RECT 37.160 128.930 37.480 129.190 ;
        RECT 43.140 129.130 43.460 129.190 ;
        RECT 43.615 129.130 43.905 129.175 ;
        RECT 43.140 128.990 43.905 129.130 ;
        RECT 43.140 128.930 43.460 128.990 ;
        RECT 43.615 128.945 43.905 128.990 ;
        RECT 46.360 129.130 46.680 129.190 ;
        RECT 51.880 129.130 52.200 129.190 ;
        RECT 54.655 129.130 54.945 129.175 ;
        RECT 46.360 128.990 54.945 129.130 ;
        RECT 46.360 128.930 46.680 128.990 ;
        RECT 51.880 128.930 52.200 128.990 ;
        RECT 54.655 128.945 54.945 128.990 ;
        RECT 32.100 128.790 32.420 128.850 ;
        RECT 33.035 128.790 33.325 128.835 ;
        RECT 39.935 128.790 40.225 128.835 ;
        RECT 40.840 128.790 41.160 128.850 ;
        RECT 32.100 128.650 39.690 128.790 ;
        RECT 32.100 128.590 32.420 128.650 ;
        RECT 33.035 128.605 33.325 128.650 ;
        RECT 26.135 128.265 26.425 128.495 ;
        RECT 28.420 128.250 28.740 128.510 ;
        RECT 28.880 128.450 29.200 128.510 ;
        RECT 33.495 128.450 33.785 128.495 ;
        RECT 28.880 128.310 33.785 128.450 ;
        RECT 28.880 128.250 29.200 128.310 ;
        RECT 33.495 128.265 33.785 128.310 ;
        RECT 35.335 128.450 35.625 128.495 ;
        RECT 37.160 128.450 37.480 128.510 ;
        RECT 35.335 128.310 37.480 128.450 ;
        RECT 35.335 128.265 35.625 128.310 ;
        RECT 37.160 128.250 37.480 128.310 ;
        RECT 37.635 128.450 37.925 128.495 ;
        RECT 38.080 128.450 38.400 128.510 ;
        RECT 39.550 128.495 39.690 128.650 ;
        RECT 39.935 128.650 41.160 128.790 ;
        RECT 54.730 128.790 54.870 128.945 ;
        RECT 55.100 128.930 55.420 129.190 ;
        RECT 59.255 128.790 59.545 128.835 ;
        RECT 54.730 128.650 59.545 128.790 ;
        RECT 39.935 128.605 40.225 128.650 ;
        RECT 40.840 128.590 41.160 128.650 ;
        RECT 59.255 128.605 59.545 128.650 ;
        RECT 62.000 128.790 62.320 128.850 ;
        RECT 63.010 128.835 63.150 129.330 ;
        RECT 68.440 129.270 68.760 129.330 ;
        RECT 69.375 129.285 69.665 129.515 ;
        RECT 63.855 129.130 64.145 129.175 ;
        RECT 64.760 129.130 65.080 129.190 ;
        RECT 63.855 128.990 65.080 129.130 ;
        RECT 63.855 128.945 64.145 128.990 ;
        RECT 64.760 128.930 65.080 128.990 ;
        RECT 67.075 129.130 67.365 129.175 ;
        RECT 69.450 129.130 69.590 129.285 ;
        RECT 72.670 129.130 72.810 129.670 ;
        RECT 73.520 129.670 78.450 129.810 ;
        RECT 73.520 129.625 73.810 129.670 ;
        RECT 75.380 129.625 75.670 129.670 ;
        RECT 78.160 129.625 78.450 129.670 ;
        RECT 83.710 129.670 88.450 129.810 ;
        RECT 73.040 129.270 73.360 129.530 ;
        RECT 74.880 129.270 75.200 129.530 ;
        RECT 83.710 129.470 83.850 129.670 ;
        RECT 75.430 129.330 83.850 129.470 ;
        RECT 75.430 129.130 75.570 129.330 ;
        RECT 84.080 129.270 84.400 129.530 ;
        RECT 88.310 129.470 88.450 129.670 ;
        RECT 88.680 129.670 101.330 129.810 ;
        RECT 88.680 129.610 89.000 129.670 ;
        RECT 96.960 129.610 97.280 129.670 ;
        RECT 98.800 129.470 99.120 129.530 ;
        RECT 88.310 129.330 94.430 129.470 ;
        RECT 78.160 129.130 78.450 129.175 ;
        RECT 67.075 128.990 71.890 129.130 ;
        RECT 72.670 128.990 75.570 129.130 ;
        RECT 75.915 128.990 78.450 129.130 ;
        RECT 67.075 128.945 67.365 128.990 ;
        RECT 62.935 128.790 63.225 128.835 ;
        RECT 62.000 128.650 63.225 128.790 ;
        RECT 62.000 128.590 62.320 128.650 ;
        RECT 62.935 128.605 63.225 128.650 ;
        RECT 63.380 128.790 63.700 128.850 ;
        RECT 65.235 128.790 65.525 128.835 ;
        RECT 63.380 128.650 65.525 128.790 ;
        RECT 63.380 128.590 63.700 128.650 ;
        RECT 65.235 128.605 65.525 128.650 ;
        RECT 70.295 128.790 70.585 128.835 ;
        RECT 71.200 128.790 71.520 128.850 ;
        RECT 70.295 128.650 71.520 128.790 ;
        RECT 71.750 128.790 71.890 128.990 ;
        RECT 72.580 128.790 72.900 128.850 ;
        RECT 75.915 128.835 76.130 128.990 ;
        RECT 78.160 128.945 78.450 128.990 ;
        RECT 88.220 128.930 88.540 129.190 ;
        RECT 89.230 129.175 89.370 129.330 ;
        RECT 89.155 128.945 89.445 129.175 ;
        RECT 90.535 128.945 90.825 129.175 ;
        RECT 90.980 129.130 91.300 129.190 ;
        RECT 94.290 129.175 94.430 129.330 ;
        RECT 97.510 129.330 99.120 129.470 ;
        RECT 97.510 129.175 97.650 129.330 ;
        RECT 98.800 129.270 99.120 129.330 ;
        RECT 100.180 129.270 100.500 129.530 ;
        RECT 101.190 129.515 101.330 129.670 ;
        RECT 101.115 129.285 101.405 129.515 ;
        RECT 101.650 129.470 101.790 130.010 ;
        RECT 108.935 130.010 110.160 130.150 ;
        RECT 108.935 129.965 109.225 130.010 ;
        RECT 109.840 129.950 110.160 130.010 ;
        RECT 103.415 129.810 103.705 129.855 ;
        RECT 103.415 129.670 108.230 129.810 ;
        RECT 103.415 129.625 103.705 129.670 ;
        RECT 104.335 129.470 104.625 129.515 ;
        RECT 101.650 129.330 104.625 129.470 ;
        RECT 104.335 129.285 104.625 129.330 ;
        RECT 93.295 129.130 93.585 129.175 ;
        RECT 90.980 128.990 93.585 129.130 ;
        RECT 71.750 128.650 72.900 128.790 ;
        RECT 70.295 128.605 70.585 128.650 ;
        RECT 71.200 128.590 71.520 128.650 ;
        RECT 72.580 128.590 72.900 128.650 ;
        RECT 73.980 128.790 74.270 128.835 ;
        RECT 75.840 128.790 76.130 128.835 ;
        RECT 73.980 128.650 76.130 128.790 ;
        RECT 73.980 128.605 74.270 128.650 ;
        RECT 75.840 128.605 76.130 128.650 ;
        RECT 76.760 128.790 77.050 128.835 ;
        RECT 77.640 128.790 77.960 128.850 ;
        RECT 80.020 128.790 80.310 128.835 ;
        RECT 76.760 128.650 80.310 128.790 ;
        RECT 76.760 128.605 77.050 128.650 ;
        RECT 77.640 128.590 77.960 128.650 ;
        RECT 80.020 128.605 80.310 128.650 ;
        RECT 85.015 128.790 85.305 128.835 ;
        RECT 88.680 128.790 89.000 128.850 ;
        RECT 85.015 128.650 89.000 128.790 ;
        RECT 85.015 128.605 85.305 128.650 ;
        RECT 88.680 128.590 89.000 128.650 ;
        RECT 37.635 128.310 38.400 128.450 ;
        RECT 37.635 128.265 37.925 128.310 ;
        RECT 38.080 128.250 38.400 128.310 ;
        RECT 39.475 128.450 39.765 128.495 ;
        RECT 42.680 128.450 43.000 128.510 ;
        RECT 39.475 128.310 43.000 128.450 ;
        RECT 39.475 128.265 39.765 128.310 ;
        RECT 42.680 128.250 43.000 128.310 ;
        RECT 56.940 128.250 57.260 128.510 ;
        RECT 58.320 128.450 58.640 128.510 ;
        RECT 58.795 128.450 59.085 128.495 ;
        RECT 58.320 128.310 59.085 128.450 ;
        RECT 58.320 128.250 58.640 128.310 ;
        RECT 58.795 128.265 59.085 128.310 ;
        RECT 61.095 128.450 61.385 128.495 ;
        RECT 61.540 128.450 61.860 128.510 ;
        RECT 61.095 128.310 61.860 128.450 ;
        RECT 61.095 128.265 61.385 128.310 ;
        RECT 61.540 128.250 61.860 128.310 ;
        RECT 70.755 128.450 71.045 128.495 ;
        RECT 80.860 128.450 81.180 128.510 ;
        RECT 82.025 128.450 82.315 128.495 ;
        RECT 84.555 128.450 84.845 128.495 ;
        RECT 70.755 128.310 84.845 128.450 ;
        RECT 70.755 128.265 71.045 128.310 ;
        RECT 80.860 128.250 81.180 128.310 ;
        RECT 82.025 128.265 82.315 128.310 ;
        RECT 84.555 128.265 84.845 128.310 ;
        RECT 86.855 128.450 87.145 128.495 ;
        RECT 90.610 128.450 90.750 128.945 ;
        RECT 90.980 128.930 91.300 128.990 ;
        RECT 93.295 128.945 93.585 128.990 ;
        RECT 94.215 129.130 94.505 129.175 ;
        RECT 97.435 129.130 97.725 129.175 ;
        RECT 94.215 128.990 97.725 129.130 ;
        RECT 94.215 128.945 94.505 128.990 ;
        RECT 97.435 128.945 97.725 128.990 ;
        RECT 98.340 128.930 98.660 129.190 ;
        RECT 99.720 129.130 100.040 129.190 ;
        RECT 108.090 129.175 108.230 129.670 ;
        RECT 101.575 129.130 101.865 129.175 ;
        RECT 105.255 129.130 105.545 129.175 ;
        RECT 99.720 128.990 105.545 129.130 ;
        RECT 99.720 128.930 100.040 128.990 ;
        RECT 101.575 128.945 101.865 128.990 ;
        RECT 105.255 128.945 105.545 128.990 ;
        RECT 108.015 128.945 108.305 129.175 ;
        RECT 86.855 128.310 90.750 128.450 ;
        RECT 104.780 128.450 105.100 128.510 ;
        RECT 105.715 128.450 106.005 128.495 ;
        RECT 104.780 128.310 106.005 128.450 ;
        RECT 86.855 128.265 87.145 128.310 ;
        RECT 104.780 128.250 105.100 128.310 ;
        RECT 105.715 128.265 106.005 128.310 ;
        RECT 106.620 128.450 106.940 128.510 ;
        RECT 107.555 128.450 107.845 128.495 ;
        RECT 106.620 128.310 107.845 128.450 ;
        RECT 106.620 128.250 106.940 128.310 ;
        RECT 107.555 128.265 107.845 128.310 ;
        RECT 15.010 127.630 113.450 128.110 ;
        RECT 20.615 127.430 20.905 127.475 ;
        RECT 21.060 127.430 21.380 127.490 ;
        RECT 20.615 127.290 21.380 127.430 ;
        RECT 20.615 127.245 20.905 127.290 ;
        RECT 21.060 127.230 21.380 127.290 ;
        RECT 21.520 127.430 21.840 127.490 ;
        RECT 26.135 127.430 26.425 127.475 ;
        RECT 29.800 127.430 30.120 127.490 ;
        RECT 32.100 127.475 32.420 127.490 ;
        RECT 21.520 127.290 30.120 127.430 ;
        RECT 21.520 127.230 21.840 127.290 ;
        RECT 26.135 127.245 26.425 127.290 ;
        RECT 29.800 127.230 30.120 127.290 ;
        RECT 31.885 127.245 32.420 127.475 ;
        RECT 32.100 127.230 32.420 127.245 ;
        RECT 41.300 127.230 41.620 127.490 ;
        RECT 48.215 127.430 48.505 127.475 ;
        RECT 49.580 127.430 49.900 127.490 ;
        RECT 48.215 127.290 49.900 127.430 ;
        RECT 48.215 127.245 48.505 127.290 ;
        RECT 49.580 127.230 49.900 127.290 ;
        RECT 57.185 127.430 57.475 127.475 ;
        RECT 58.320 127.430 58.640 127.490 ;
        RECT 62.000 127.430 62.320 127.490 ;
        RECT 57.185 127.290 58.640 127.430 ;
        RECT 57.185 127.245 57.475 127.290 ;
        RECT 58.320 127.230 58.640 127.290 ;
        RECT 58.870 127.290 62.320 127.430 ;
        RECT 20.140 127.090 20.460 127.150 ;
        RECT 26.595 127.090 26.885 127.135 ;
        RECT 20.140 126.950 26.885 127.090 ;
        RECT 20.140 126.890 20.460 126.950 ;
        RECT 26.595 126.905 26.885 126.950 ;
        RECT 28.420 127.090 28.740 127.150 ;
        RECT 33.890 127.090 34.180 127.135 ;
        RECT 37.150 127.090 37.440 127.135 ;
        RECT 28.420 126.950 37.440 127.090 ;
        RECT 28.420 126.890 28.740 126.950 ;
        RECT 33.890 126.905 34.180 126.950 ;
        RECT 37.150 126.905 37.440 126.950 ;
        RECT 38.070 127.090 38.360 127.135 ;
        RECT 39.930 127.090 40.220 127.135 ;
        RECT 38.070 126.950 40.220 127.090 ;
        RECT 38.070 126.905 38.360 126.950 ;
        RECT 39.930 126.905 40.220 126.950 ;
        RECT 40.380 127.090 40.700 127.150 ;
        RECT 44.075 127.090 44.365 127.135 ;
        RECT 58.870 127.090 59.010 127.290 ;
        RECT 62.000 127.230 62.320 127.290 ;
        RECT 65.680 127.430 66.000 127.490 ;
        RECT 73.500 127.430 73.820 127.490 ;
        RECT 74.895 127.430 75.185 127.475 ;
        RECT 65.680 127.290 73.270 127.430 ;
        RECT 65.680 127.230 66.000 127.290 ;
        RECT 62.460 127.135 62.780 127.150 ;
        RECT 40.380 126.950 44.365 127.090 ;
        RECT 21.075 126.750 21.365 126.795 ;
        RECT 23.360 126.750 23.680 126.810 ;
        RECT 27.960 126.750 28.280 126.810 ;
        RECT 21.075 126.610 28.280 126.750 ;
        RECT 21.075 126.565 21.365 126.610 ;
        RECT 23.360 126.550 23.680 126.610 ;
        RECT 27.960 126.550 28.280 126.610 ;
        RECT 35.750 126.750 36.040 126.795 ;
        RECT 38.070 126.750 38.285 126.905 ;
        RECT 40.380 126.890 40.700 126.950 ;
        RECT 44.075 126.905 44.365 126.950 ;
        RECT 47.370 126.950 59.010 127.090 ;
        RECT 59.190 127.090 59.480 127.135 ;
        RECT 62.450 127.090 62.780 127.135 ;
        RECT 59.190 126.950 62.780 127.090 ;
        RECT 35.750 126.610 38.285 126.750 ;
        RECT 35.750 126.565 36.040 126.610 ;
        RECT 39.000 126.550 39.320 126.810 ;
        RECT 42.235 126.565 42.525 126.795 ;
        RECT 20.600 126.410 20.920 126.470 ;
        RECT 27.515 126.410 27.805 126.455 ;
        RECT 30.720 126.410 31.040 126.470 ;
        RECT 20.600 126.270 31.040 126.410 ;
        RECT 20.600 126.210 20.920 126.270 ;
        RECT 27.515 126.225 27.805 126.270 ;
        RECT 30.720 126.210 31.040 126.270 ;
        RECT 36.240 126.410 36.560 126.470 ;
        RECT 40.855 126.410 41.145 126.455 ;
        RECT 36.240 126.270 41.145 126.410 ;
        RECT 36.240 126.210 36.560 126.270 ;
        RECT 40.855 126.225 41.145 126.270 ;
        RECT 41.760 126.410 42.080 126.470 ;
        RECT 42.310 126.410 42.450 126.565 ;
        RECT 42.680 126.550 43.000 126.810 ;
        RECT 47.370 126.795 47.510 126.950 ;
        RECT 59.190 126.905 59.480 126.950 ;
        RECT 62.450 126.905 62.780 126.950 ;
        RECT 62.460 126.890 62.780 126.905 ;
        RECT 63.370 127.090 63.660 127.135 ;
        RECT 65.230 127.090 65.520 127.135 ;
        RECT 72.120 127.090 72.440 127.150 ;
        RECT 63.370 126.950 65.520 127.090 ;
        RECT 63.370 126.905 63.660 126.950 ;
        RECT 65.230 126.905 65.520 126.950 ;
        RECT 66.230 126.950 72.440 127.090 ;
        RECT 44.995 126.750 45.285 126.795 ;
        RECT 47.295 126.750 47.585 126.795 ;
        RECT 43.230 126.610 47.585 126.750 ;
        RECT 43.230 126.410 43.370 126.610 ;
        RECT 44.995 126.565 45.285 126.610 ;
        RECT 47.295 126.565 47.585 126.610 ;
        RECT 50.500 126.550 50.820 126.810 ;
        RECT 55.575 126.750 55.865 126.795 ;
        RECT 56.940 126.750 57.260 126.810 ;
        RECT 55.575 126.610 57.260 126.750 ;
        RECT 55.575 126.565 55.865 126.610 ;
        RECT 56.940 126.550 57.260 126.610 ;
        RECT 61.050 126.750 61.340 126.795 ;
        RECT 63.370 126.750 63.585 126.905 ;
        RECT 66.230 126.795 66.370 126.950 ;
        RECT 72.120 126.890 72.440 126.950 ;
        RECT 61.050 126.610 63.585 126.750 ;
        RECT 61.050 126.565 61.340 126.610 ;
        RECT 66.155 126.565 66.445 126.795 ;
        RECT 68.915 126.750 69.205 126.795 ;
        RECT 68.915 126.610 69.590 126.750 ;
        RECT 68.915 126.565 69.205 126.610 ;
        RECT 41.760 126.270 43.370 126.410 ;
        RECT 44.520 126.410 44.840 126.470 ;
        RECT 45.915 126.410 46.205 126.455 ;
        RECT 44.520 126.270 46.205 126.410 ;
        RECT 41.760 126.210 42.080 126.270 ;
        RECT 44.520 126.210 44.840 126.270 ;
        RECT 45.915 126.225 46.205 126.270 ;
        RECT 46.360 126.210 46.680 126.470 ;
        RECT 64.300 126.210 64.620 126.470 ;
        RECT 69.450 126.115 69.590 126.610 ;
        RECT 71.200 126.550 71.520 126.810 ;
        RECT 70.280 126.410 70.600 126.470 ;
        RECT 71.675 126.410 71.965 126.455 ;
        RECT 70.280 126.270 71.965 126.410 ;
        RECT 70.280 126.210 70.600 126.270 ;
        RECT 71.675 126.225 71.965 126.270 ;
        RECT 72.580 126.210 72.900 126.470 ;
        RECT 73.130 126.410 73.270 127.290 ;
        RECT 73.500 127.290 75.185 127.430 ;
        RECT 73.500 127.230 73.820 127.290 ;
        RECT 74.895 127.245 75.185 127.290 ;
        RECT 77.640 127.230 77.960 127.490 ;
        RECT 87.300 127.230 87.620 127.490 ;
        RECT 102.020 127.475 102.340 127.490 ;
        RECT 102.020 127.430 102.555 127.475 ;
        RECT 104.780 127.430 105.100 127.490 ;
        RECT 102.020 127.290 105.100 127.430 ;
        RECT 102.020 127.245 102.555 127.290 ;
        RECT 102.020 127.230 102.340 127.245 ;
        RECT 104.780 127.230 105.100 127.290 ;
        RECT 99.275 127.090 99.565 127.135 ;
        RECT 104.270 127.090 104.560 127.135 ;
        RECT 107.530 127.090 107.820 127.135 ;
        RECT 86.930 126.950 99.030 127.090 ;
        RECT 75.800 126.550 76.120 126.810 ;
        RECT 76.260 126.550 76.580 126.810 ;
        RECT 77.195 126.565 77.485 126.795 ;
        RECT 85.460 126.750 85.780 126.810 ;
        RECT 86.930 126.795 87.070 126.950 ;
        RECT 86.855 126.750 87.145 126.795 ;
        RECT 85.460 126.610 87.145 126.750 ;
        RECT 77.270 126.410 77.410 126.565 ;
        RECT 85.460 126.550 85.780 126.610 ;
        RECT 86.855 126.565 87.145 126.610 ;
        RECT 88.220 126.750 88.540 126.810 ;
        RECT 93.370 126.795 93.510 126.950 ;
        RECT 98.890 126.795 99.030 126.950 ;
        RECT 99.275 126.950 107.820 127.090 ;
        RECT 99.275 126.905 99.565 126.950 ;
        RECT 104.270 126.905 104.560 126.950 ;
        RECT 107.530 126.905 107.820 126.950 ;
        RECT 108.450 127.090 108.740 127.135 ;
        RECT 110.310 127.090 110.600 127.135 ;
        RECT 108.450 126.950 110.600 127.090 ;
        RECT 108.450 126.905 108.740 126.950 ;
        RECT 110.310 126.905 110.600 126.950 ;
        RECT 90.995 126.750 91.285 126.795 ;
        RECT 88.220 126.610 91.285 126.750 ;
        RECT 88.220 126.550 88.540 126.610 ;
        RECT 90.995 126.565 91.285 126.610 ;
        RECT 93.295 126.565 93.585 126.795 ;
        RECT 96.515 126.750 96.805 126.795 ;
        RECT 93.830 126.610 96.805 126.750 ;
        RECT 73.130 126.270 77.410 126.410 ;
        RECT 84.080 126.410 84.400 126.470 ;
        RECT 89.615 126.410 89.905 126.455 ;
        RECT 84.080 126.270 89.905 126.410 ;
        RECT 84.080 126.210 84.400 126.270 ;
        RECT 89.615 126.225 89.905 126.270 ;
        RECT 90.520 126.410 90.840 126.470 ;
        RECT 93.830 126.410 93.970 126.610 ;
        RECT 96.515 126.565 96.805 126.610 ;
        RECT 98.815 126.750 99.105 126.795 ;
        RECT 100.640 126.750 100.960 126.810 ;
        RECT 98.815 126.610 100.960 126.750 ;
        RECT 98.815 126.565 99.105 126.610 ;
        RECT 100.640 126.550 100.960 126.610 ;
        RECT 106.130 126.750 106.420 126.795 ;
        RECT 108.450 126.750 108.665 126.905 ;
        RECT 106.130 126.610 108.665 126.750 ;
        RECT 106.130 126.565 106.420 126.610 ;
        RECT 90.520 126.270 93.970 126.410 ;
        RECT 35.750 126.070 36.040 126.115 ;
        RECT 38.530 126.070 38.820 126.115 ;
        RECT 40.390 126.070 40.680 126.115 ;
        RECT 35.750 125.930 40.680 126.070 ;
        RECT 35.750 125.885 36.040 125.930 ;
        RECT 38.530 125.885 38.820 125.930 ;
        RECT 40.390 125.885 40.680 125.930 ;
        RECT 61.050 126.070 61.340 126.115 ;
        RECT 63.830 126.070 64.120 126.115 ;
        RECT 65.690 126.070 65.980 126.115 ;
        RECT 61.050 125.930 65.980 126.070 ;
        RECT 61.050 125.885 61.340 125.930 ;
        RECT 63.830 125.885 64.120 125.930 ;
        RECT 65.690 125.885 65.980 125.930 ;
        RECT 69.375 125.885 69.665 126.115 ;
        RECT 89.690 126.070 89.830 126.225 ;
        RECT 90.520 126.210 90.840 126.270 ;
        RECT 95.135 126.225 95.425 126.455 ;
        RECT 96.055 126.410 96.345 126.455 ;
        RECT 98.340 126.410 98.660 126.470 ;
        RECT 99.720 126.410 100.040 126.470 ;
        RECT 96.055 126.270 100.040 126.410 ;
        RECT 96.055 126.225 96.345 126.270 ;
        RECT 95.210 126.070 95.350 126.225 ;
        RECT 98.340 126.210 98.660 126.270 ;
        RECT 99.720 126.210 100.040 126.270 ;
        RECT 109.395 126.410 109.685 126.455 ;
        RECT 109.840 126.410 110.160 126.470 ;
        RECT 109.395 126.270 110.160 126.410 ;
        RECT 109.395 126.225 109.685 126.270 ;
        RECT 109.840 126.210 110.160 126.270 ;
        RECT 111.220 126.210 111.540 126.470 ;
        RECT 100.180 126.070 100.500 126.130 ;
        RECT 89.690 125.930 100.500 126.070 ;
        RECT 100.180 125.870 100.500 125.930 ;
        RECT 106.130 126.070 106.420 126.115 ;
        RECT 108.910 126.070 109.200 126.115 ;
        RECT 110.770 126.070 111.060 126.115 ;
        RECT 106.130 125.930 111.060 126.070 ;
        RECT 106.130 125.885 106.420 125.930 ;
        RECT 108.910 125.885 109.200 125.930 ;
        RECT 110.770 125.885 111.060 125.930 ;
        RECT 24.295 125.730 24.585 125.775 ;
        RECT 25.660 125.730 25.980 125.790 ;
        RECT 24.295 125.590 25.980 125.730 ;
        RECT 24.295 125.545 24.585 125.590 ;
        RECT 25.660 125.530 25.980 125.590 ;
        RECT 56.480 125.530 56.800 125.790 ;
        RECT 66.600 125.730 66.920 125.790 ;
        RECT 67.995 125.730 68.285 125.775 ;
        RECT 66.600 125.590 68.285 125.730 ;
        RECT 66.600 125.530 66.920 125.590 ;
        RECT 67.995 125.545 68.285 125.590 ;
        RECT 68.440 125.730 68.760 125.790 ;
        RECT 75.800 125.730 76.120 125.790 ;
        RECT 68.440 125.590 76.120 125.730 ;
        RECT 68.440 125.530 68.760 125.590 ;
        RECT 75.800 125.530 76.120 125.590 ;
        RECT 91.440 125.730 91.760 125.790 ;
        RECT 92.835 125.730 93.125 125.775 ;
        RECT 91.440 125.590 93.125 125.730 ;
        RECT 91.440 125.530 91.760 125.590 ;
        RECT 92.835 125.545 93.125 125.590 ;
        RECT 93.740 125.530 94.060 125.790 ;
        RECT 98.340 125.530 98.660 125.790 ;
        RECT 101.100 125.530 101.420 125.790 ;
        RECT 15.010 124.910 113.450 125.390 ;
        RECT 20.385 124.710 20.675 124.755 ;
        RECT 21.520 124.710 21.840 124.770 ;
        RECT 20.385 124.570 21.840 124.710 ;
        RECT 20.385 124.525 20.675 124.570 ;
        RECT 21.520 124.510 21.840 124.570 ;
        RECT 39.000 124.510 39.320 124.770 ;
        RECT 51.880 124.755 52.200 124.770 ;
        RECT 51.880 124.525 52.415 124.755 ;
        RECT 51.880 124.510 52.200 124.525 ;
        RECT 62.460 124.510 62.780 124.770 ;
        RECT 64.300 124.510 64.620 124.770 ;
        RECT 68.225 124.710 68.515 124.755 ;
        RECT 70.280 124.710 70.600 124.770 ;
        RECT 68.225 124.570 70.600 124.710 ;
        RECT 68.225 124.525 68.515 124.570 ;
        RECT 70.280 124.510 70.600 124.570 ;
        RECT 72.580 124.710 72.900 124.770 ;
        RECT 84.080 124.710 84.400 124.770 ;
        RECT 72.580 124.570 84.400 124.710 ;
        RECT 72.580 124.510 72.900 124.570 ;
        RECT 19.235 124.370 19.525 124.415 ;
        RECT 21.980 124.370 22.300 124.430 ;
        RECT 19.235 124.230 22.300 124.370 ;
        RECT 19.235 124.185 19.525 124.230 ;
        RECT 21.980 124.170 22.300 124.230 ;
        RECT 24.250 124.370 24.540 124.415 ;
        RECT 27.030 124.370 27.320 124.415 ;
        RECT 28.890 124.370 29.180 124.415 ;
        RECT 36.240 124.370 36.560 124.430 ;
        RECT 24.250 124.230 29.180 124.370 ;
        RECT 24.250 124.185 24.540 124.230 ;
        RECT 27.030 124.185 27.320 124.230 ;
        RECT 28.890 124.185 29.180 124.230 ;
        RECT 29.430 124.230 36.560 124.370 ;
        RECT 29.430 124.090 29.570 124.230 ;
        RECT 36.240 124.170 36.560 124.230 ;
        RECT 38.540 124.370 38.860 124.430 ;
        RECT 41.315 124.370 41.605 124.415 ;
        RECT 38.540 124.230 41.605 124.370 ;
        RECT 38.540 124.170 38.860 124.230 ;
        RECT 41.315 124.185 41.605 124.230 ;
        RECT 49.580 124.170 49.900 124.430 ;
        RECT 55.990 124.370 56.280 124.415 ;
        RECT 58.770 124.370 59.060 124.415 ;
        RECT 60.630 124.370 60.920 124.415 ;
        RECT 55.990 124.230 60.920 124.370 ;
        RECT 55.990 124.185 56.280 124.230 ;
        RECT 58.770 124.185 59.060 124.230 ;
        RECT 60.630 124.185 60.920 124.230 ;
        RECT 72.090 124.370 72.380 124.415 ;
        RECT 74.870 124.370 75.160 124.415 ;
        RECT 76.730 124.370 77.020 124.415 ;
        RECT 72.090 124.230 77.020 124.370 ;
        RECT 72.090 124.185 72.380 124.230 ;
        RECT 74.870 124.185 75.160 124.230 ;
        RECT 76.730 124.185 77.020 124.230 ;
        RECT 26.580 124.030 26.900 124.090 ;
        RECT 27.515 124.030 27.805 124.075 ;
        RECT 26.580 123.890 27.805 124.030 ;
        RECT 26.580 123.830 26.900 123.890 ;
        RECT 27.515 123.845 27.805 123.890 ;
        RECT 29.340 123.830 29.660 124.090 ;
        RECT 30.720 123.830 31.040 124.090 ;
        RECT 31.640 124.030 31.960 124.090 ;
        RECT 39.475 124.030 39.765 124.075 ;
        RECT 41.760 124.030 42.080 124.090 ;
        RECT 31.640 123.890 39.765 124.030 ;
        RECT 31.640 123.830 31.960 123.890 ;
        RECT 39.475 123.845 39.765 123.890 ;
        RECT 40.470 123.890 42.080 124.030 ;
        RECT 19.695 123.690 19.985 123.735 ;
        RECT 23.360 123.690 23.680 123.750 ;
        RECT 19.695 123.550 23.680 123.690 ;
        RECT 19.695 123.505 19.985 123.550 ;
        RECT 23.360 123.490 23.680 123.550 ;
        RECT 24.250 123.690 24.540 123.735 ;
        RECT 24.250 123.550 26.785 123.690 ;
        RECT 24.250 123.505 24.540 123.550 ;
        RECT 22.390 123.350 22.680 123.395 ;
        RECT 23.820 123.350 24.140 123.410 ;
        RECT 26.570 123.395 26.785 123.550 ;
        RECT 25.650 123.350 25.940 123.395 ;
        RECT 22.390 123.210 25.940 123.350 ;
        RECT 22.390 123.165 22.680 123.210 ;
        RECT 23.820 123.150 24.140 123.210 ;
        RECT 25.650 123.165 25.940 123.210 ;
        RECT 26.570 123.350 26.860 123.395 ;
        RECT 28.430 123.350 28.720 123.395 ;
        RECT 26.570 123.210 28.720 123.350 ;
        RECT 26.570 123.165 26.860 123.210 ;
        RECT 28.430 123.165 28.720 123.210 ;
        RECT 30.260 123.010 30.580 123.070 ;
        RECT 31.730 123.055 31.870 123.830 ;
        RECT 38.080 123.490 38.400 123.750 ;
        RECT 40.470 123.735 40.610 123.890 ;
        RECT 41.760 123.830 42.080 123.890 ;
        RECT 44.995 124.030 45.285 124.075 ;
        RECT 46.835 124.030 47.125 124.075 ;
        RECT 51.420 124.030 51.740 124.090 ;
        RECT 44.995 123.890 51.740 124.030 ;
        RECT 44.995 123.845 45.285 123.890 ;
        RECT 46.835 123.845 47.125 123.890 ;
        RECT 51.420 123.830 51.740 123.890 ;
        RECT 56.480 124.030 56.800 124.090 ;
        RECT 59.255 124.030 59.545 124.075 ;
        RECT 56.480 123.890 59.545 124.030 ;
        RECT 56.480 123.830 56.800 123.890 ;
        RECT 59.255 123.845 59.545 123.890 ;
        RECT 61.540 124.030 61.860 124.090 ;
        RECT 73.040 124.030 73.360 124.090 ;
        RECT 74.420 124.030 74.740 124.090 ;
        RECT 61.540 123.890 63.610 124.030 ;
        RECT 61.540 123.830 61.860 123.890 ;
        RECT 40.395 123.505 40.685 123.735 ;
        RECT 46.360 123.690 46.680 123.750 ;
        RECT 47.295 123.690 47.585 123.735 ;
        RECT 40.930 123.550 47.585 123.690 ;
        RECT 40.930 123.350 41.070 123.550 ;
        RECT 46.360 123.490 46.680 123.550 ;
        RECT 47.295 123.505 47.585 123.550 ;
        RECT 55.990 123.690 56.280 123.735 ;
        RECT 55.990 123.550 58.525 123.690 ;
        RECT 55.990 123.505 56.280 123.550 ;
        RECT 32.190 123.210 41.070 123.350 ;
        RECT 41.300 123.350 41.620 123.410 ;
        RECT 43.615 123.350 43.905 123.395 ;
        RECT 47.755 123.350 48.045 123.395 ;
        RECT 41.300 123.210 43.905 123.350 ;
        RECT 32.190 123.070 32.330 123.210 ;
        RECT 41.300 123.150 41.620 123.210 ;
        RECT 43.615 123.165 43.905 123.210 ;
        RECT 44.610 123.210 48.045 123.350 ;
        RECT 44.610 123.070 44.750 123.210 ;
        RECT 47.755 123.165 48.045 123.210 ;
        RECT 54.130 123.350 54.420 123.395 ;
        RECT 55.560 123.350 55.880 123.410 ;
        RECT 58.310 123.395 58.525 123.550 ;
        RECT 61.095 123.505 61.385 123.735 ;
        RECT 62.000 123.690 62.320 123.750 ;
        RECT 63.470 123.735 63.610 123.890 ;
        RECT 73.040 123.890 75.110 124.030 ;
        RECT 73.040 123.830 73.360 123.890 ;
        RECT 74.420 123.830 74.740 123.890 ;
        RECT 62.935 123.690 63.225 123.735 ;
        RECT 62.000 123.550 63.225 123.690 ;
        RECT 57.390 123.350 57.680 123.395 ;
        RECT 54.130 123.210 57.680 123.350 ;
        RECT 54.130 123.165 54.420 123.210 ;
        RECT 55.560 123.150 55.880 123.210 ;
        RECT 57.390 123.165 57.680 123.210 ;
        RECT 58.310 123.350 58.600 123.395 ;
        RECT 60.170 123.350 60.460 123.395 ;
        RECT 58.310 123.210 60.460 123.350 ;
        RECT 58.310 123.165 58.600 123.210 ;
        RECT 60.170 123.165 60.460 123.210 ;
        RECT 31.655 123.010 31.945 123.055 ;
        RECT 30.260 122.870 31.945 123.010 ;
        RECT 30.260 122.810 30.580 122.870 ;
        RECT 31.655 122.825 31.945 122.870 ;
        RECT 32.100 122.810 32.420 123.070 ;
        RECT 33.955 123.010 34.245 123.055 ;
        RECT 34.860 123.010 35.180 123.070 ;
        RECT 33.955 122.870 35.180 123.010 ;
        RECT 33.955 122.825 34.245 122.870 ;
        RECT 34.860 122.810 35.180 122.870 ;
        RECT 41.775 123.010 42.065 123.055 ;
        RECT 42.220 123.010 42.540 123.070 ;
        RECT 41.775 122.870 42.540 123.010 ;
        RECT 41.775 122.825 42.065 122.870 ;
        RECT 42.220 122.810 42.540 122.870 ;
        RECT 44.075 123.010 44.365 123.055 ;
        RECT 44.520 123.010 44.840 123.070 ;
        RECT 44.075 122.870 44.840 123.010 ;
        RECT 44.075 122.825 44.365 122.870 ;
        RECT 44.520 122.810 44.840 122.870 ;
        RECT 47.280 123.010 47.600 123.070 ;
        RECT 50.500 123.010 50.820 123.070 ;
        RECT 56.480 123.010 56.800 123.070 ;
        RECT 61.170 123.010 61.310 123.505 ;
        RECT 62.000 123.490 62.320 123.550 ;
        RECT 62.935 123.505 63.225 123.550 ;
        RECT 63.395 123.505 63.685 123.735 ;
        RECT 65.680 123.690 66.000 123.750 ;
        RECT 66.615 123.690 66.905 123.735 ;
        RECT 65.680 123.550 66.905 123.690 ;
        RECT 65.680 123.490 66.000 123.550 ;
        RECT 66.615 123.505 66.905 123.550 ;
        RECT 72.090 123.690 72.380 123.735 ;
        RECT 74.970 123.690 75.110 123.890 ;
        RECT 75.340 123.830 75.660 124.090 ;
        RECT 81.870 124.075 82.010 124.570 ;
        RECT 84.080 124.510 84.400 124.570 ;
        RECT 90.520 124.755 90.840 124.770 ;
        RECT 90.520 124.525 91.055 124.755 ;
        RECT 90.520 124.510 90.840 124.525 ;
        RECT 94.630 124.370 94.920 124.415 ;
        RECT 97.410 124.370 97.700 124.415 ;
        RECT 99.270 124.370 99.560 124.415 ;
        RECT 94.630 124.230 99.560 124.370 ;
        RECT 94.630 124.185 94.920 124.230 ;
        RECT 97.410 124.185 97.700 124.230 ;
        RECT 99.270 124.185 99.560 124.230 ;
        RECT 99.720 124.370 100.040 124.430 ;
        RECT 100.425 124.370 100.715 124.415 ;
        RECT 102.480 124.370 102.800 124.430 ;
        RECT 99.720 124.230 102.800 124.370 ;
        RECT 99.720 124.170 100.040 124.230 ;
        RECT 100.425 124.185 100.715 124.230 ;
        RECT 102.480 124.170 102.800 124.230 ;
        RECT 104.290 124.370 104.580 124.415 ;
        RECT 107.070 124.370 107.360 124.415 ;
        RECT 108.930 124.370 109.220 124.415 ;
        RECT 104.290 124.230 109.220 124.370 ;
        RECT 104.290 124.185 104.580 124.230 ;
        RECT 107.070 124.185 107.360 124.230 ;
        RECT 108.930 124.185 109.220 124.230 ;
        RECT 81.795 123.845 82.085 124.075 ;
        RECT 82.715 124.030 83.005 124.075 ;
        RECT 88.220 124.030 88.540 124.090 ;
        RECT 82.715 123.890 88.540 124.030 ;
        RECT 82.715 123.845 83.005 123.890 ;
        RECT 88.220 123.830 88.540 123.890 ;
        RECT 99.810 123.890 107.310 124.030 ;
        RECT 99.810 123.750 99.950 123.890 ;
        RECT 77.195 123.690 77.485 123.735 ;
        RECT 86.840 123.690 87.160 123.750 ;
        RECT 72.090 123.550 74.625 123.690 ;
        RECT 74.970 123.550 87.160 123.690 ;
        RECT 72.090 123.505 72.380 123.550 ;
        RECT 70.230 123.350 70.520 123.395 ;
        RECT 70.740 123.350 71.060 123.410 ;
        RECT 74.410 123.395 74.625 123.550 ;
        RECT 77.195 123.505 77.485 123.550 ;
        RECT 86.840 123.490 87.160 123.550 ;
        RECT 94.630 123.690 94.920 123.735 ;
        RECT 94.630 123.550 97.165 123.690 ;
        RECT 94.630 123.505 94.920 123.550 ;
        RECT 73.490 123.350 73.780 123.395 ;
        RECT 70.230 123.210 73.780 123.350 ;
        RECT 70.230 123.165 70.520 123.210 ;
        RECT 70.740 123.150 71.060 123.210 ;
        RECT 73.490 123.165 73.780 123.210 ;
        RECT 74.410 123.350 74.700 123.395 ;
        RECT 76.270 123.350 76.560 123.395 ;
        RECT 74.410 123.210 76.560 123.350 ;
        RECT 74.410 123.165 74.700 123.210 ;
        RECT 76.270 123.165 76.560 123.210 ;
        RECT 92.770 123.350 93.060 123.395 ;
        RECT 93.740 123.350 94.060 123.410 ;
        RECT 96.950 123.395 97.165 123.550 ;
        RECT 97.880 123.490 98.200 123.750 ;
        RECT 99.720 123.490 100.040 123.750 ;
        RECT 104.290 123.690 104.580 123.735 ;
        RECT 107.170 123.690 107.310 123.890 ;
        RECT 107.540 123.830 107.860 124.090 ;
        RECT 109.395 123.690 109.685 123.735 ;
        RECT 111.220 123.690 111.540 123.750 ;
        RECT 104.290 123.550 106.825 123.690 ;
        RECT 107.170 123.550 111.540 123.690 ;
        RECT 104.290 123.505 104.580 123.550 ;
        RECT 96.030 123.350 96.320 123.395 ;
        RECT 92.770 123.210 96.320 123.350 ;
        RECT 92.770 123.165 93.060 123.210 ;
        RECT 93.740 123.150 94.060 123.210 ;
        RECT 96.030 123.165 96.320 123.210 ;
        RECT 96.950 123.350 97.240 123.395 ;
        RECT 98.810 123.350 99.100 123.395 ;
        RECT 96.950 123.210 99.100 123.350 ;
        RECT 96.950 123.165 97.240 123.210 ;
        RECT 98.810 123.165 99.100 123.210 ;
        RECT 101.100 123.350 101.420 123.410 ;
        RECT 106.610 123.395 106.825 123.550 ;
        RECT 109.395 123.505 109.685 123.550 ;
        RECT 111.220 123.490 111.540 123.550 ;
        RECT 102.430 123.350 102.720 123.395 ;
        RECT 105.690 123.350 105.980 123.395 ;
        RECT 101.100 123.210 105.980 123.350 ;
        RECT 101.100 123.150 101.420 123.210 ;
        RECT 102.430 123.165 102.720 123.210 ;
        RECT 105.690 123.165 105.980 123.210 ;
        RECT 106.610 123.350 106.900 123.395 ;
        RECT 108.470 123.350 108.760 123.395 ;
        RECT 106.610 123.210 108.760 123.350 ;
        RECT 106.610 123.165 106.900 123.210 ;
        RECT 108.470 123.165 108.760 123.210 ;
        RECT 47.280 122.870 61.310 123.010 ;
        RECT 67.075 123.010 67.365 123.055 ;
        RECT 68.440 123.010 68.760 123.070 ;
        RECT 67.075 122.870 68.760 123.010 ;
        RECT 47.280 122.810 47.600 122.870 ;
        RECT 50.500 122.810 50.820 122.870 ;
        RECT 56.480 122.810 56.800 122.870 ;
        RECT 67.075 122.825 67.365 122.870 ;
        RECT 68.440 122.810 68.760 122.870 ;
        RECT 76.720 123.010 77.040 123.070 ;
        RECT 83.175 123.010 83.465 123.055 ;
        RECT 76.720 122.870 83.465 123.010 ;
        RECT 76.720 122.810 77.040 122.870 ;
        RECT 83.175 122.825 83.465 122.870 ;
        RECT 84.540 123.010 84.860 123.070 ;
        RECT 85.015 123.010 85.305 123.055 ;
        RECT 84.540 122.870 85.305 123.010 ;
        RECT 84.540 122.810 84.860 122.870 ;
        RECT 85.015 122.825 85.305 122.870 ;
        RECT 15.010 122.190 113.450 122.670 ;
        RECT 18.775 121.805 19.065 122.035 ;
        RECT 21.075 121.990 21.365 122.035 ;
        RECT 21.520 121.990 21.840 122.050 ;
        RECT 21.075 121.850 21.840 121.990 ;
        RECT 21.075 121.805 21.365 121.850 ;
        RECT 17.395 121.310 17.685 121.355 ;
        RECT 18.850 121.310 18.990 121.805 ;
        RECT 21.520 121.790 21.840 121.850 ;
        RECT 23.820 121.790 24.140 122.050 ;
        RECT 26.580 121.790 26.900 122.050 ;
        RECT 27.285 121.990 27.575 122.035 ;
        RECT 32.100 121.990 32.420 122.050 ;
        RECT 27.285 121.850 32.420 121.990 ;
        RECT 27.285 121.805 27.575 121.850 ;
        RECT 32.100 121.790 32.420 121.850 ;
        RECT 38.325 121.990 38.615 122.035 ;
        RECT 41.300 121.990 41.620 122.050 ;
        RECT 38.325 121.850 41.620 121.990 ;
        RECT 38.325 121.805 38.615 121.850 ;
        RECT 41.300 121.790 41.620 121.850 ;
        RECT 55.560 121.990 55.880 122.050 ;
        RECT 56.495 121.990 56.785 122.035 ;
        RECT 55.560 121.850 56.785 121.990 ;
        RECT 55.560 121.790 55.880 121.850 ;
        RECT 56.495 121.805 56.785 121.850 ;
        RECT 71.200 121.990 71.520 122.050 ;
        RECT 73.745 121.990 74.035 122.035 ;
        RECT 71.200 121.850 74.035 121.990 ;
        RECT 71.200 121.790 71.520 121.850 ;
        RECT 73.745 121.805 74.035 121.850 ;
        RECT 75.340 121.990 75.660 122.050 ;
        RECT 75.815 121.990 76.105 122.035 ;
        RECT 75.340 121.850 76.105 121.990 ;
        RECT 75.340 121.790 75.660 121.850 ;
        RECT 75.815 121.805 76.105 121.850 ;
        RECT 83.620 121.990 83.940 122.050 ;
        RECT 87.545 121.990 87.835 122.035 ;
        RECT 88.220 121.990 88.540 122.050 ;
        RECT 83.620 121.850 87.070 121.990 ;
        RECT 83.620 121.790 83.940 121.850 ;
        RECT 20.615 121.650 20.905 121.695 ;
        RECT 29.290 121.650 29.580 121.695 ;
        RECT 30.720 121.650 31.040 121.710 ;
        RECT 32.550 121.650 32.840 121.695 ;
        RECT 20.615 121.510 29.110 121.650 ;
        RECT 20.615 121.465 20.905 121.510 ;
        RECT 17.395 121.170 18.990 121.310 ;
        RECT 23.360 121.310 23.680 121.370 ;
        RECT 24.740 121.310 25.060 121.370 ;
        RECT 23.360 121.170 25.060 121.310 ;
        RECT 17.395 121.125 17.685 121.170 ;
        RECT 23.360 121.110 23.680 121.170 ;
        RECT 24.740 121.110 25.060 121.170 ;
        RECT 25.660 121.110 25.980 121.370 ;
        RECT 28.970 121.310 29.110 121.510 ;
        RECT 29.290 121.510 32.840 121.650 ;
        RECT 29.290 121.465 29.580 121.510 ;
        RECT 30.720 121.450 31.040 121.510 ;
        RECT 32.550 121.465 32.840 121.510 ;
        RECT 33.470 121.650 33.760 121.695 ;
        RECT 35.330 121.650 35.620 121.695 ;
        RECT 33.470 121.510 35.620 121.650 ;
        RECT 33.470 121.465 33.760 121.510 ;
        RECT 35.330 121.465 35.620 121.510 ;
        RECT 40.330 121.650 40.620 121.695 ;
        RECT 41.760 121.650 42.080 121.710 ;
        RECT 43.590 121.650 43.880 121.695 ;
        RECT 40.330 121.510 43.880 121.650 ;
        RECT 40.330 121.465 40.620 121.510 ;
        RECT 30.260 121.310 30.580 121.370 ;
        RECT 28.970 121.170 30.580 121.310 ;
        RECT 30.260 121.110 30.580 121.170 ;
        RECT 31.150 121.310 31.440 121.355 ;
        RECT 33.470 121.310 33.685 121.465 ;
        RECT 41.760 121.450 42.080 121.510 ;
        RECT 43.590 121.465 43.880 121.510 ;
        RECT 44.510 121.650 44.800 121.695 ;
        RECT 46.370 121.650 46.660 121.695 ;
        RECT 44.510 121.510 46.660 121.650 ;
        RECT 44.510 121.465 44.800 121.510 ;
        RECT 46.370 121.465 46.660 121.510 ;
        RECT 49.580 121.650 49.900 121.710 ;
        RECT 68.440 121.695 68.760 121.710 ;
        RECT 65.700 121.650 65.990 121.695 ;
        RECT 67.560 121.650 67.850 121.695 ;
        RECT 49.580 121.510 50.730 121.650 ;
        RECT 31.150 121.170 33.685 121.310 ;
        RECT 31.150 121.125 31.440 121.170 ;
        RECT 36.240 121.110 36.560 121.370 ;
        RECT 42.190 121.310 42.480 121.355 ;
        RECT 44.510 121.310 44.725 121.465 ;
        RECT 49.580 121.450 49.900 121.510 ;
        RECT 42.190 121.170 44.725 121.310 ;
        RECT 42.190 121.125 42.480 121.170 ;
        RECT 47.280 121.110 47.600 121.370 ;
        RECT 50.590 121.355 50.730 121.510 ;
        RECT 65.700 121.510 67.850 121.650 ;
        RECT 65.700 121.465 65.990 121.510 ;
        RECT 67.560 121.465 67.850 121.510 ;
        RECT 50.055 121.125 50.345 121.355 ;
        RECT 50.515 121.125 50.805 121.355 ;
        RECT 54.195 121.310 54.485 121.355 ;
        RECT 56.020 121.310 56.340 121.370 ;
        RECT 56.955 121.310 57.245 121.355 ;
        RECT 62.000 121.310 62.320 121.370 ;
        RECT 54.195 121.170 62.320 121.310 ;
        RECT 54.195 121.125 54.485 121.170 ;
        RECT 20.600 120.970 20.920 121.030 ;
        RECT 21.535 120.970 21.825 121.015 ;
        RECT 20.600 120.830 21.825 120.970 ;
        RECT 20.600 120.770 20.920 120.830 ;
        RECT 21.535 120.785 21.825 120.830 ;
        RECT 34.400 120.770 34.720 121.030 ;
        RECT 44.060 120.970 44.380 121.030 ;
        RECT 45.455 120.970 45.745 121.015 ;
        RECT 44.060 120.830 45.745 120.970 ;
        RECT 44.060 120.770 44.380 120.830 ;
        RECT 45.455 120.785 45.745 120.830 ;
        RECT 50.130 120.970 50.270 121.125 ;
        RECT 56.020 121.110 56.340 121.170 ;
        RECT 56.955 121.125 57.245 121.170 ;
        RECT 62.000 121.110 62.320 121.170 ;
        RECT 66.600 121.110 66.920 121.370 ;
        RECT 67.635 121.310 67.850 121.465 ;
        RECT 68.440 121.650 68.770 121.695 ;
        RECT 71.740 121.650 72.030 121.695 ;
        RECT 68.440 121.510 72.030 121.650 ;
        RECT 68.440 121.465 68.770 121.510 ;
        RECT 71.740 121.465 72.030 121.510 ;
        RECT 79.890 121.650 80.180 121.695 ;
        RECT 81.320 121.650 81.640 121.710 ;
        RECT 83.150 121.650 83.440 121.695 ;
        RECT 79.890 121.510 83.440 121.650 ;
        RECT 79.890 121.465 80.180 121.510 ;
        RECT 68.440 121.450 68.760 121.465 ;
        RECT 81.320 121.450 81.640 121.510 ;
        RECT 83.150 121.465 83.440 121.510 ;
        RECT 84.070 121.650 84.360 121.695 ;
        RECT 85.930 121.650 86.220 121.695 ;
        RECT 84.070 121.510 86.220 121.650 ;
        RECT 86.930 121.650 87.070 121.850 ;
        RECT 87.545 121.850 88.540 121.990 ;
        RECT 87.545 121.805 87.835 121.850 ;
        RECT 88.220 121.790 88.540 121.850 ;
        RECT 97.435 121.990 97.725 122.035 ;
        RECT 97.880 121.990 98.200 122.050 ;
        RECT 97.435 121.850 98.200 121.990 ;
        RECT 97.435 121.805 97.725 121.850 ;
        RECT 97.880 121.790 98.200 121.850 ;
        RECT 102.020 121.790 102.340 122.050 ;
        RECT 102.480 121.790 102.800 122.050 ;
        RECT 104.335 121.805 104.625 122.035 ;
        RECT 105.715 121.990 106.005 122.035 ;
        RECT 107.080 121.990 107.400 122.050 ;
        RECT 105.715 121.850 107.400 121.990 ;
        RECT 105.715 121.805 106.005 121.850 ;
        RECT 89.550 121.650 89.840 121.695 ;
        RECT 92.810 121.650 93.100 121.695 ;
        RECT 86.930 121.510 93.100 121.650 ;
        RECT 84.070 121.465 84.360 121.510 ;
        RECT 85.930 121.465 86.220 121.510 ;
        RECT 89.550 121.465 89.840 121.510 ;
        RECT 92.810 121.465 93.100 121.510 ;
        RECT 93.730 121.650 94.020 121.695 ;
        RECT 95.590 121.650 95.880 121.695 ;
        RECT 93.730 121.510 95.880 121.650 ;
        RECT 93.730 121.465 94.020 121.510 ;
        RECT 95.590 121.465 95.880 121.510 ;
        RECT 69.880 121.310 70.170 121.355 ;
        RECT 67.635 121.170 70.170 121.310 ;
        RECT 69.880 121.125 70.170 121.170 ;
        RECT 74.880 121.110 75.200 121.370 ;
        RECT 81.750 121.310 82.040 121.355 ;
        RECT 84.070 121.310 84.285 121.465 ;
        RECT 81.750 121.170 84.285 121.310 ;
        RECT 81.750 121.125 82.040 121.170 ;
        RECT 85.000 121.110 85.320 121.370 ;
        RECT 91.410 121.310 91.700 121.355 ;
        RECT 93.730 121.310 93.945 121.465 ;
        RECT 91.410 121.170 93.945 121.310 ;
        RECT 91.410 121.125 91.700 121.170 ;
        RECT 98.340 121.110 98.660 121.370 ;
        RECT 104.410 121.310 104.550 121.805 ;
        RECT 107.080 121.790 107.400 121.850 ;
        RECT 107.555 121.990 107.845 122.035 ;
        RECT 109.840 121.990 110.160 122.050 ;
        RECT 107.555 121.850 110.160 121.990 ;
        RECT 107.555 121.805 107.845 121.850 ;
        RECT 109.840 121.790 110.160 121.850 ;
        RECT 104.795 121.310 105.085 121.355 ;
        RECT 104.410 121.170 105.085 121.310 ;
        RECT 104.795 121.125 105.085 121.170 ;
        RECT 106.620 121.110 106.940 121.370 ;
        RECT 52.815 120.970 53.105 121.015 ;
        RECT 50.130 120.830 53.105 120.970 ;
        RECT 18.315 120.630 18.605 120.675 ;
        RECT 25.200 120.630 25.520 120.690 ;
        RECT 18.315 120.490 25.520 120.630 ;
        RECT 18.315 120.445 18.605 120.490 ;
        RECT 25.200 120.430 25.520 120.490 ;
        RECT 31.150 120.630 31.440 120.675 ;
        RECT 33.930 120.630 34.220 120.675 ;
        RECT 35.790 120.630 36.080 120.675 ;
        RECT 31.150 120.490 36.080 120.630 ;
        RECT 31.150 120.445 31.440 120.490 ;
        RECT 33.930 120.445 34.220 120.490 ;
        RECT 35.790 120.445 36.080 120.490 ;
        RECT 42.190 120.630 42.480 120.675 ;
        RECT 44.970 120.630 45.260 120.675 ;
        RECT 46.830 120.630 47.120 120.675 ;
        RECT 50.130 120.630 50.270 120.830 ;
        RECT 52.815 120.785 53.105 120.830 ;
        RECT 56.480 120.970 56.800 121.030 ;
        RECT 64.775 120.970 65.065 121.015 ;
        RECT 56.480 120.830 65.065 120.970 ;
        RECT 56.480 120.770 56.800 120.830 ;
        RECT 64.775 120.785 65.065 120.830 ;
        RECT 86.840 120.770 87.160 121.030 ;
        RECT 91.900 120.970 92.220 121.030 ;
        RECT 94.675 120.970 94.965 121.015 ;
        RECT 91.900 120.830 94.965 120.970 ;
        RECT 91.900 120.770 92.220 120.830 ;
        RECT 94.675 120.785 94.965 120.830 ;
        RECT 96.515 120.970 96.805 121.015 ;
        RECT 99.720 120.970 100.040 121.030 ;
        RECT 96.515 120.830 100.040 120.970 ;
        RECT 96.515 120.785 96.805 120.830 ;
        RECT 99.720 120.770 100.040 120.830 ;
        RECT 100.180 120.970 100.500 121.030 ;
        RECT 101.115 120.970 101.405 121.015 ;
        RECT 100.180 120.830 101.405 120.970 ;
        RECT 100.180 120.770 100.500 120.830 ;
        RECT 101.115 120.785 101.405 120.830 ;
        RECT 42.190 120.490 47.120 120.630 ;
        RECT 42.190 120.445 42.480 120.490 ;
        RECT 44.970 120.445 45.260 120.490 ;
        RECT 46.830 120.445 47.120 120.490 ;
        RECT 47.370 120.490 50.270 120.630 ;
        RECT 65.240 120.630 65.530 120.675 ;
        RECT 67.100 120.630 67.390 120.675 ;
        RECT 69.880 120.630 70.170 120.675 ;
        RECT 65.240 120.490 70.170 120.630 ;
        RECT 41.300 120.290 41.620 120.350 ;
        RECT 47.370 120.290 47.510 120.490 ;
        RECT 65.240 120.445 65.530 120.490 ;
        RECT 67.100 120.445 67.390 120.490 ;
        RECT 69.880 120.445 70.170 120.490 ;
        RECT 81.750 120.630 82.040 120.675 ;
        RECT 84.530 120.630 84.820 120.675 ;
        RECT 86.390 120.630 86.680 120.675 ;
        RECT 81.750 120.490 86.680 120.630 ;
        RECT 81.750 120.445 82.040 120.490 ;
        RECT 84.530 120.445 84.820 120.490 ;
        RECT 86.390 120.445 86.680 120.490 ;
        RECT 91.410 120.630 91.700 120.675 ;
        RECT 94.190 120.630 94.480 120.675 ;
        RECT 96.050 120.630 96.340 120.675 ;
        RECT 91.410 120.490 96.340 120.630 ;
        RECT 91.410 120.445 91.700 120.490 ;
        RECT 94.190 120.445 94.480 120.490 ;
        RECT 96.050 120.445 96.340 120.490 ;
        RECT 41.300 120.150 47.510 120.290 ;
        RECT 41.300 120.090 41.620 120.150 ;
        RECT 49.580 120.090 49.900 120.350 ;
        RECT 51.435 120.290 51.725 120.335 ;
        RECT 51.880 120.290 52.200 120.350 ;
        RECT 51.435 120.150 52.200 120.290 ;
        RECT 51.435 120.105 51.725 120.150 ;
        RECT 51.880 120.090 52.200 120.150 ;
        RECT 73.040 120.290 73.360 120.350 ;
        RECT 76.260 120.290 76.580 120.350 ;
        RECT 77.885 120.290 78.175 120.335 ;
        RECT 73.040 120.150 78.175 120.290 ;
        RECT 73.040 120.090 73.360 120.150 ;
        RECT 76.260 120.090 76.580 120.150 ;
        RECT 77.885 120.105 78.175 120.150 ;
        RECT 15.010 119.470 113.450 119.950 ;
        RECT 24.740 119.270 25.060 119.330 ;
        RECT 24.740 119.130 30.490 119.270 ;
        RECT 24.740 119.070 25.060 119.130 ;
        RECT 23.475 118.930 23.765 118.975 ;
        RECT 26.595 118.930 26.885 118.975 ;
        RECT 28.485 118.930 28.775 118.975 ;
        RECT 23.475 118.790 28.775 118.930 ;
        RECT 23.475 118.745 23.765 118.790 ;
        RECT 26.595 118.745 26.885 118.790 ;
        RECT 28.485 118.745 28.775 118.790 ;
        RECT 29.340 118.390 29.660 118.650 ;
        RECT 30.350 118.590 30.490 119.130 ;
        RECT 30.720 119.070 31.040 119.330 ;
        RECT 34.400 119.070 34.720 119.330 ;
        RECT 41.760 119.070 42.080 119.330 ;
        RECT 44.060 119.070 44.380 119.330 ;
        RECT 44.520 119.315 44.840 119.330 ;
        RECT 44.520 119.085 45.055 119.315 ;
        RECT 44.520 119.070 44.840 119.085 ;
        RECT 70.740 119.070 71.060 119.330 ;
        RECT 74.880 119.270 75.200 119.330 ;
        RECT 75.355 119.270 75.645 119.315 ;
        RECT 74.880 119.130 75.645 119.270 ;
        RECT 74.880 119.070 75.200 119.130 ;
        RECT 75.355 119.085 75.645 119.130 ;
        RECT 83.620 119.070 83.940 119.330 ;
        RECT 85.000 119.270 85.320 119.330 ;
        RECT 85.475 119.270 85.765 119.315 ;
        RECT 85.000 119.130 85.765 119.270 ;
        RECT 85.000 119.070 85.320 119.130 ;
        RECT 85.475 119.085 85.765 119.130 ;
        RECT 91.900 119.070 92.220 119.330 ;
        RECT 105.700 119.270 106.020 119.330 ;
        RECT 105.700 119.130 109.150 119.270 ;
        RECT 105.700 119.070 106.020 119.130 ;
        RECT 48.630 118.930 48.920 118.975 ;
        RECT 51.410 118.930 51.700 118.975 ;
        RECT 53.270 118.930 53.560 118.975 ;
        RECT 48.630 118.790 53.560 118.930 ;
        RECT 48.630 118.745 48.920 118.790 ;
        RECT 51.410 118.745 51.700 118.790 ;
        RECT 53.270 118.745 53.560 118.790 ;
        RECT 108.475 118.745 108.765 118.975 ;
        RECT 30.350 118.450 41.530 118.590 ;
        RECT 30.350 118.295 30.490 118.450 ;
        RECT 41.390 118.310 41.530 118.450 ;
        RECT 51.880 118.390 52.200 118.650 ;
        RECT 72.580 118.390 72.900 118.650 ;
        RECT 73.040 118.390 73.360 118.650 ;
        RECT 105.330 118.450 107.310 118.590 ;
        RECT 19.235 117.910 19.525 117.955 ;
        RECT 21.060 117.910 21.380 117.970 ;
        RECT 19.235 117.770 21.380 117.910 ;
        RECT 19.235 117.725 19.525 117.770 ;
        RECT 21.060 117.710 21.380 117.770 ;
        RECT 21.520 117.910 21.840 117.970 ;
        RECT 22.395 117.955 22.685 118.270 ;
        RECT 23.475 118.250 23.765 118.295 ;
        RECT 27.055 118.250 27.345 118.295 ;
        RECT 28.890 118.250 29.180 118.295 ;
        RECT 23.475 118.110 29.180 118.250 ;
        RECT 23.475 118.065 23.765 118.110 ;
        RECT 27.055 118.065 27.345 118.110 ;
        RECT 28.890 118.065 29.180 118.110 ;
        RECT 30.275 118.065 30.565 118.295 ;
        RECT 33.495 118.250 33.785 118.295 ;
        RECT 34.860 118.250 35.180 118.310 ;
        RECT 33.495 118.110 35.180 118.250 ;
        RECT 33.495 118.065 33.785 118.110 ;
        RECT 34.860 118.050 35.180 118.110 ;
        RECT 41.300 118.050 41.620 118.310 ;
        RECT 42.220 118.250 42.540 118.310 ;
        RECT 43.155 118.250 43.445 118.295 ;
        RECT 42.220 118.110 43.445 118.250 ;
        RECT 42.220 118.050 42.540 118.110 ;
        RECT 43.155 118.065 43.445 118.110 ;
        RECT 48.630 118.250 48.920 118.295 ;
        RECT 53.735 118.250 54.025 118.295 ;
        RECT 56.480 118.250 56.800 118.310 ;
        RECT 48.630 118.110 51.165 118.250 ;
        RECT 48.630 118.065 48.920 118.110 ;
        RECT 22.095 117.910 22.685 117.955 ;
        RECT 25.335 117.910 25.985 117.955 ;
        RECT 21.520 117.770 25.985 117.910 ;
        RECT 21.520 117.710 21.840 117.770 ;
        RECT 22.095 117.725 22.385 117.770 ;
        RECT 25.335 117.725 25.985 117.770 ;
        RECT 27.960 117.710 28.280 117.970 ;
        RECT 46.770 117.910 47.060 117.955 ;
        RECT 49.120 117.910 49.440 117.970 ;
        RECT 50.950 117.955 51.165 118.110 ;
        RECT 53.735 118.110 56.800 118.250 ;
        RECT 53.735 118.065 54.025 118.110 ;
        RECT 56.480 118.050 56.800 118.110 ;
        RECT 65.680 118.250 66.000 118.310 ;
        RECT 70.295 118.250 70.585 118.295 ;
        RECT 65.680 118.110 70.585 118.250 ;
        RECT 65.680 118.050 66.000 118.110 ;
        RECT 70.295 118.065 70.585 118.110 ;
        RECT 81.320 118.250 81.640 118.310 ;
        RECT 81.795 118.250 82.085 118.295 ;
        RECT 81.320 118.110 82.085 118.250 ;
        RECT 50.030 117.910 50.320 117.955 ;
        RECT 46.770 117.770 50.320 117.910 ;
        RECT 46.770 117.725 47.060 117.770 ;
        RECT 49.120 117.710 49.440 117.770 ;
        RECT 50.030 117.725 50.320 117.770 ;
        RECT 50.950 117.910 51.240 117.955 ;
        RECT 52.810 117.910 53.100 117.955 ;
        RECT 50.950 117.770 53.100 117.910 ;
        RECT 70.370 117.910 70.510 118.065 ;
        RECT 81.320 118.050 81.640 118.110 ;
        RECT 81.795 118.065 82.085 118.110 ;
        RECT 82.255 118.250 82.545 118.295 ;
        RECT 83.175 118.250 83.465 118.295 ;
        RECT 82.255 118.110 83.465 118.250 ;
        RECT 82.255 118.065 82.545 118.110 ;
        RECT 83.175 118.065 83.465 118.110 ;
        RECT 82.330 117.910 82.470 118.065 ;
        RECT 84.540 118.050 84.860 118.310 ;
        RECT 90.995 118.250 91.285 118.295 ;
        RECT 91.440 118.250 91.760 118.310 ;
        RECT 105.330 118.250 105.470 118.450 ;
        RECT 90.995 118.110 91.760 118.250 ;
        RECT 90.995 118.065 91.285 118.110 ;
        RECT 91.440 118.050 91.760 118.110 ;
        RECT 91.990 118.110 105.470 118.250 ;
        RECT 105.715 118.250 106.005 118.295 ;
        RECT 106.620 118.250 106.940 118.310 ;
        RECT 107.170 118.295 107.310 118.450 ;
        RECT 105.715 118.110 106.940 118.250 ;
        RECT 70.370 117.770 82.470 117.910 ;
        RECT 90.060 117.910 90.380 117.970 ;
        RECT 91.990 117.910 92.130 118.110 ;
        RECT 105.715 118.065 106.005 118.110 ;
        RECT 106.620 118.050 106.940 118.110 ;
        RECT 107.095 118.065 107.385 118.295 ;
        RECT 90.060 117.770 92.130 117.910 ;
        RECT 102.940 117.910 103.260 117.970 ;
        RECT 108.550 117.910 108.690 118.745 ;
        RECT 109.010 118.250 109.150 119.130 ;
        RECT 109.395 118.250 109.685 118.295 ;
        RECT 109.010 118.110 109.685 118.250 ;
        RECT 109.395 118.065 109.685 118.110 ;
        RECT 102.940 117.770 108.690 117.910 ;
        RECT 50.950 117.725 51.240 117.770 ;
        RECT 52.810 117.725 53.100 117.770 ;
        RECT 90.060 117.710 90.380 117.770 ;
        RECT 102.940 117.710 103.260 117.770 ;
        RECT 70.280 117.570 70.600 117.630 ;
        RECT 73.515 117.570 73.805 117.615 ;
        RECT 70.280 117.430 73.805 117.570 ;
        RECT 70.280 117.370 70.600 117.430 ;
        RECT 73.515 117.385 73.805 117.430 ;
        RECT 106.160 117.370 106.480 117.630 ;
        RECT 108.015 117.570 108.305 117.615 ;
        RECT 110.300 117.570 110.620 117.630 ;
        RECT 108.015 117.430 110.620 117.570 ;
        RECT 108.015 117.385 108.305 117.430 ;
        RECT 110.300 117.370 110.620 117.430 ;
        RECT 15.010 116.750 113.450 117.230 ;
        RECT 66.140 116.550 66.460 116.610 ;
        RECT 70.295 116.550 70.585 116.595 ;
        RECT 66.140 116.410 70.585 116.550 ;
        RECT 66.140 116.350 66.460 116.410 ;
        RECT 70.295 116.365 70.585 116.410 ;
        RECT 20.600 116.210 20.920 116.270 ;
        RECT 26.235 116.210 26.525 116.255 ;
        RECT 29.475 116.210 30.125 116.255 ;
        RECT 20.600 116.070 30.125 116.210 ;
        RECT 20.600 116.010 20.920 116.070 ;
        RECT 26.235 116.025 26.825 116.070 ;
        RECT 29.475 116.025 30.125 116.070 ;
        RECT 69.820 116.210 70.140 116.270 ;
        RECT 73.055 116.210 73.345 116.255 ;
        RECT 69.820 116.070 72.810 116.210 ;
        RECT 26.535 115.710 26.825 116.025 ;
        RECT 69.820 116.010 70.140 116.070 ;
        RECT 27.615 115.870 27.905 115.915 ;
        RECT 31.195 115.870 31.485 115.915 ;
        RECT 33.030 115.870 33.320 115.915 ;
        RECT 27.615 115.730 33.320 115.870 ;
        RECT 27.615 115.685 27.905 115.730 ;
        RECT 31.195 115.685 31.485 115.730 ;
        RECT 33.030 115.685 33.320 115.730 ;
        RECT 35.335 115.870 35.625 115.915 ;
        RECT 35.780 115.870 36.100 115.930 ;
        RECT 35.335 115.730 36.100 115.870 ;
        RECT 35.335 115.685 35.625 115.730 ;
        RECT 35.780 115.670 36.100 115.730 ;
        RECT 36.700 115.870 37.020 115.930 ;
        RECT 47.295 115.870 47.585 115.915 ;
        RECT 36.700 115.730 47.585 115.870 ;
        RECT 36.700 115.670 37.020 115.730 ;
        RECT 47.295 115.685 47.585 115.730 ;
        RECT 56.020 115.670 56.340 115.930 ;
        RECT 70.740 115.670 71.060 115.930 ;
        RECT 71.675 115.870 71.965 115.915 ;
        RECT 72.670 115.870 72.810 116.070 ;
        RECT 73.055 116.070 84.310 116.210 ;
        RECT 73.055 116.025 73.345 116.070 ;
        RECT 84.170 115.930 84.310 116.070 ;
        RECT 102.940 116.010 103.260 116.270 ;
        RECT 105.235 116.210 105.885 116.255 ;
        RECT 106.160 116.210 106.480 116.270 ;
        RECT 108.835 116.210 109.125 116.255 ;
        RECT 105.235 116.070 109.125 116.210 ;
        RECT 105.235 116.025 105.885 116.070 ;
        RECT 106.160 116.010 106.480 116.070 ;
        RECT 108.535 116.025 109.125 116.070 ;
        RECT 77.655 115.870 77.945 115.915 ;
        RECT 71.675 115.730 72.350 115.870 ;
        RECT 72.670 115.730 77.945 115.870 ;
        RECT 71.675 115.685 71.965 115.730 ;
        RECT 16.000 115.530 16.320 115.590 ;
        RECT 23.375 115.530 23.665 115.575 ;
        RECT 16.000 115.390 23.665 115.530 ;
        RECT 16.000 115.330 16.320 115.390 ;
        RECT 23.375 115.345 23.665 115.390 ;
        RECT 29.340 115.530 29.660 115.590 ;
        RECT 33.495 115.530 33.785 115.575 ;
        RECT 29.340 115.390 33.785 115.530 ;
        RECT 29.340 115.330 29.660 115.390 ;
        RECT 33.495 115.345 33.785 115.390 ;
        RECT 27.615 115.190 27.905 115.235 ;
        RECT 30.735 115.190 31.025 115.235 ;
        RECT 32.625 115.190 32.915 115.235 ;
        RECT 27.615 115.050 32.915 115.190 ;
        RECT 33.570 115.190 33.710 115.345 ;
        RECT 35.320 115.190 35.640 115.250 ;
        RECT 33.570 115.050 35.640 115.190 ;
        RECT 56.110 115.190 56.250 115.670 ;
        RECT 56.940 115.330 57.260 115.590 ;
        RECT 72.210 115.190 72.350 115.730 ;
        RECT 77.655 115.685 77.945 115.730 ;
        RECT 84.080 115.670 84.400 115.930 ;
        RECT 87.760 115.870 88.080 115.930 ;
        RECT 89.615 115.870 89.905 115.915 ;
        RECT 87.760 115.730 89.905 115.870 ;
        RECT 87.760 115.670 88.080 115.730 ;
        RECT 89.615 115.685 89.905 115.730 ;
        RECT 94.675 115.870 94.965 115.915 ;
        RECT 95.580 115.870 95.900 115.930 ;
        RECT 94.675 115.730 95.900 115.870 ;
        RECT 94.675 115.685 94.965 115.730 ;
        RECT 95.580 115.670 95.900 115.730 ;
        RECT 98.815 115.870 99.105 115.915 ;
        RECT 99.260 115.870 99.580 115.930 ;
        RECT 98.815 115.730 99.580 115.870 ;
        RECT 98.815 115.685 99.105 115.730 ;
        RECT 99.260 115.670 99.580 115.730 ;
        RECT 102.040 115.870 102.330 115.915 ;
        RECT 103.875 115.870 104.165 115.915 ;
        RECT 107.455 115.870 107.745 115.915 ;
        RECT 102.040 115.730 107.745 115.870 ;
        RECT 102.040 115.685 102.330 115.730 ;
        RECT 103.875 115.685 104.165 115.730 ;
        RECT 107.455 115.685 107.745 115.730 ;
        RECT 108.535 115.710 108.825 116.025 ;
        RECT 83.160 115.530 83.480 115.590 ;
        RECT 83.635 115.530 83.925 115.575 ;
        RECT 83.160 115.390 83.925 115.530 ;
        RECT 83.160 115.330 83.480 115.390 ;
        RECT 83.635 115.345 83.925 115.390 ;
        RECT 99.720 115.530 100.040 115.590 ;
        RECT 101.575 115.530 101.865 115.575 ;
        RECT 99.720 115.390 101.865 115.530 ;
        RECT 99.720 115.330 100.040 115.390 ;
        RECT 101.575 115.345 101.865 115.390 ;
        RECT 111.695 115.530 111.985 115.575 ;
        RECT 112.140 115.530 112.460 115.590 ;
        RECT 111.695 115.390 112.460 115.530 ;
        RECT 111.695 115.345 111.985 115.390 ;
        RECT 112.140 115.330 112.460 115.390 ;
        RECT 56.110 115.050 72.350 115.190 ;
        RECT 102.445 115.190 102.735 115.235 ;
        RECT 104.335 115.190 104.625 115.235 ;
        RECT 107.455 115.190 107.745 115.235 ;
        RECT 102.445 115.050 107.745 115.190 ;
        RECT 27.615 115.005 27.905 115.050 ;
        RECT 30.735 115.005 31.025 115.050 ;
        RECT 32.625 115.005 32.915 115.050 ;
        RECT 35.320 114.990 35.640 115.050 ;
        RECT 102.445 115.005 102.735 115.050 ;
        RECT 104.335 115.005 104.625 115.050 ;
        RECT 107.455 115.005 107.745 115.050 ;
        RECT 23.360 114.850 23.680 114.910 ;
        RECT 32.180 114.850 32.470 114.895 ;
        RECT 23.360 114.710 32.470 114.850 ;
        RECT 23.360 114.650 23.680 114.710 ;
        RECT 32.180 114.665 32.470 114.710 ;
        RECT 33.940 114.850 34.260 114.910 ;
        RECT 34.415 114.850 34.705 114.895 ;
        RECT 33.940 114.710 34.705 114.850 ;
        RECT 33.940 114.650 34.260 114.710 ;
        RECT 34.415 114.665 34.705 114.710 ;
        RECT 48.215 114.850 48.505 114.895 ;
        RECT 52.340 114.850 52.660 114.910 ;
        RECT 48.215 114.710 52.660 114.850 ;
        RECT 48.215 114.665 48.505 114.710 ;
        RECT 52.340 114.650 52.660 114.710 ;
        RECT 78.575 114.850 78.865 114.895 ;
        RECT 83.620 114.850 83.940 114.910 ;
        RECT 78.575 114.710 83.940 114.850 ;
        RECT 78.575 114.665 78.865 114.710 ;
        RECT 83.620 114.650 83.940 114.710 ;
        RECT 90.520 114.650 90.840 114.910 ;
        RECT 95.580 114.650 95.900 114.910 ;
        RECT 99.735 114.850 100.025 114.895 ;
        RECT 100.180 114.850 100.500 114.910 ;
        RECT 99.735 114.710 100.500 114.850 ;
        RECT 99.735 114.665 100.025 114.710 ;
        RECT 100.180 114.650 100.500 114.710 ;
        RECT 15.010 114.030 113.450 114.510 ;
        RECT 23.360 113.630 23.680 113.890 ;
        RECT 24.755 113.830 25.045 113.875 ;
        RECT 27.960 113.830 28.280 113.890 ;
        RECT 24.755 113.690 28.280 113.830 ;
        RECT 24.755 113.645 25.045 113.690 ;
        RECT 27.960 113.630 28.280 113.690 ;
        RECT 30.260 113.830 30.580 113.890 ;
        RECT 40.395 113.830 40.685 113.875 ;
        RECT 30.260 113.690 40.685 113.830 ;
        RECT 30.260 113.630 30.580 113.690 ;
        RECT 40.395 113.645 40.685 113.690 ;
        RECT 48.660 113.830 48.980 113.890 ;
        RECT 48.660 113.690 53.950 113.830 ;
        RECT 48.660 113.630 48.980 113.690 ;
        RECT 29.455 113.490 29.745 113.535 ;
        RECT 32.575 113.490 32.865 113.535 ;
        RECT 34.465 113.490 34.755 113.535 ;
        RECT 29.455 113.350 34.755 113.490 ;
        RECT 29.455 113.305 29.745 113.350 ;
        RECT 32.575 113.305 32.865 113.350 ;
        RECT 34.465 113.305 34.755 113.350 ;
        RECT 47.855 113.490 48.145 113.535 ;
        RECT 50.975 113.490 51.265 113.535 ;
        RECT 52.865 113.490 53.155 113.535 ;
        RECT 47.855 113.350 53.155 113.490 ;
        RECT 47.855 113.305 48.145 113.350 ;
        RECT 50.975 113.305 51.265 113.350 ;
        RECT 52.865 113.305 53.155 113.350 ;
        RECT 53.810 113.490 53.950 113.690 ;
        RECT 56.480 113.490 56.800 113.550 ;
        RECT 53.810 113.350 56.800 113.490 ;
        RECT 24.280 113.150 24.600 113.210 ;
        RECT 22.530 113.010 24.600 113.150 ;
        RECT 22.530 112.855 22.670 113.010 ;
        RECT 24.280 112.950 24.600 113.010 ;
        RECT 25.215 113.150 25.505 113.195 ;
        RECT 31.180 113.150 31.500 113.210 ;
        RECT 25.215 113.010 31.500 113.150 ;
        RECT 25.215 112.965 25.505 113.010 ;
        RECT 31.180 112.950 31.500 113.010 ;
        RECT 33.940 112.950 34.260 113.210 ;
        RECT 35.320 112.950 35.640 113.210 ;
        RECT 52.340 112.950 52.660 113.210 ;
        RECT 53.810 113.195 53.950 113.350 ;
        RECT 56.480 113.290 56.800 113.350 ;
        RECT 68.555 113.490 68.845 113.535 ;
        RECT 71.675 113.490 71.965 113.535 ;
        RECT 73.565 113.490 73.855 113.535 ;
        RECT 68.555 113.350 73.855 113.490 ;
        RECT 68.555 113.305 68.845 113.350 ;
        RECT 71.675 113.305 71.965 113.350 ;
        RECT 73.565 113.305 73.855 113.350 ;
        RECT 79.135 113.490 79.425 113.535 ;
        RECT 82.255 113.490 82.545 113.535 ;
        RECT 84.145 113.490 84.435 113.535 ;
        RECT 79.135 113.350 84.435 113.490 ;
        RECT 79.135 113.305 79.425 113.350 ;
        RECT 82.255 113.305 82.545 113.350 ;
        RECT 84.145 113.305 84.435 113.350 ;
        RECT 92.935 113.490 93.225 113.535 ;
        RECT 96.055 113.490 96.345 113.535 ;
        RECT 97.945 113.490 98.235 113.535 ;
        RECT 92.935 113.350 98.235 113.490 ;
        RECT 92.935 113.305 93.225 113.350 ;
        RECT 96.055 113.305 96.345 113.350 ;
        RECT 97.945 113.305 98.235 113.350 ;
        RECT 105.815 113.490 106.105 113.535 ;
        RECT 108.935 113.490 109.225 113.535 ;
        RECT 110.825 113.490 111.115 113.535 ;
        RECT 105.815 113.350 111.115 113.490 ;
        RECT 105.815 113.305 106.105 113.350 ;
        RECT 108.935 113.305 109.225 113.350 ;
        RECT 110.825 113.305 111.115 113.350 ;
        RECT 53.735 112.965 54.025 113.195 ;
        RECT 56.940 113.150 57.260 113.210 ;
        RECT 60.160 113.150 60.480 113.210 ;
        RECT 56.110 113.010 58.090 113.150 ;
        RECT 22.455 112.625 22.745 112.855 ;
        RECT 23.835 112.810 24.125 112.855 ;
        RECT 27.500 112.810 27.820 112.870 ;
        RECT 23.835 112.670 27.820 112.810 ;
        RECT 23.835 112.625 24.125 112.670 ;
        RECT 27.500 112.610 27.820 112.670 ;
        RECT 25.200 112.470 25.520 112.530 ;
        RECT 28.375 112.515 28.665 112.830 ;
        RECT 29.455 112.810 29.745 112.855 ;
        RECT 33.035 112.810 33.325 112.855 ;
        RECT 34.870 112.810 35.160 112.855 ;
        RECT 29.455 112.670 35.160 112.810 ;
        RECT 29.455 112.625 29.745 112.670 ;
        RECT 33.035 112.625 33.325 112.670 ;
        RECT 34.870 112.625 35.160 112.670 ;
        RECT 38.080 112.610 38.400 112.870 ;
        RECT 39.460 112.810 39.780 112.870 ;
        RECT 41.315 112.810 41.605 112.855 ;
        RECT 39.460 112.670 41.605 112.810 ;
        RECT 39.460 112.610 39.780 112.670 ;
        RECT 41.315 112.625 41.605 112.670 ;
        RECT 42.235 112.810 42.525 112.855 ;
        RECT 42.680 112.810 43.000 112.870 ;
        RECT 46.820 112.830 47.140 112.870 ;
        RECT 42.235 112.670 43.000 112.810 ;
        RECT 42.235 112.625 42.525 112.670 ;
        RECT 42.680 112.610 43.000 112.670 ;
        RECT 46.775 112.610 47.140 112.830 ;
        RECT 47.855 112.810 48.145 112.855 ;
        RECT 51.435 112.810 51.725 112.855 ;
        RECT 53.270 112.810 53.560 112.855 ;
        RECT 47.855 112.670 53.560 112.810 ;
        RECT 47.855 112.625 48.145 112.670 ;
        RECT 51.435 112.625 51.725 112.670 ;
        RECT 53.270 112.625 53.560 112.670 ;
        RECT 54.180 112.610 54.500 112.870 ;
        RECT 56.110 112.820 56.250 113.010 ;
        RECT 56.940 112.950 57.260 113.010 ;
        RECT 56.455 112.820 56.745 112.865 ;
        RECT 57.950 112.855 58.090 113.010 ;
        RECT 60.160 113.010 63.150 113.150 ;
        RECT 60.160 112.950 60.480 113.010 ;
        RECT 56.110 112.810 56.745 112.820 ;
        RECT 54.730 112.680 56.745 112.810 ;
        RECT 54.730 112.670 56.250 112.680 ;
        RECT 28.075 112.470 28.665 112.515 ;
        RECT 31.315 112.470 31.965 112.515 ;
        RECT 25.200 112.330 31.965 112.470 ;
        RECT 25.200 112.270 25.520 112.330 ;
        RECT 28.075 112.285 28.365 112.330 ;
        RECT 31.315 112.285 31.965 112.330 ;
        RECT 43.615 112.470 43.905 112.515 ;
        RECT 44.520 112.470 44.840 112.530 ;
        RECT 46.775 112.515 47.065 112.610 ;
        RECT 43.615 112.330 44.840 112.470 ;
        RECT 43.615 112.285 43.905 112.330 ;
        RECT 44.520 112.270 44.840 112.330 ;
        RECT 46.475 112.470 47.065 112.515 ;
        RECT 49.715 112.470 50.365 112.515 ;
        RECT 46.475 112.330 50.365 112.470 ;
        RECT 46.475 112.285 46.765 112.330 ;
        RECT 49.715 112.285 50.365 112.330 ;
        RECT 52.800 112.470 53.120 112.530 ;
        RECT 54.730 112.470 54.870 112.670 ;
        RECT 56.455 112.635 56.745 112.680 ;
        RECT 57.875 112.625 58.165 112.855 ;
        RECT 59.700 112.810 60.020 112.870 ;
        RECT 63.010 112.855 63.150 113.010 ;
        RECT 83.620 112.950 83.940 113.210 ;
        RECT 85.015 113.150 85.305 113.195 ;
        RECT 85.460 113.150 85.780 113.210 ;
        RECT 86.840 113.150 87.160 113.210 ;
        RECT 85.015 113.010 87.160 113.150 ;
        RECT 85.015 112.965 85.305 113.010 ;
        RECT 85.460 112.950 85.780 113.010 ;
        RECT 86.840 112.950 87.160 113.010 ;
        RECT 88.695 113.150 88.985 113.195 ;
        RECT 91.440 113.150 91.760 113.210 ;
        RECT 88.695 113.010 91.760 113.150 ;
        RECT 88.695 112.965 88.985 113.010 ;
        RECT 91.440 112.950 91.760 113.010 ;
        RECT 95.580 113.150 95.900 113.210 ;
        RECT 97.435 113.150 97.725 113.195 ;
        RECT 95.580 113.010 97.725 113.150 ;
        RECT 95.580 112.950 95.900 113.010 ;
        RECT 97.435 112.965 97.725 113.010 ;
        RECT 101.575 113.150 101.865 113.195 ;
        RECT 107.080 113.150 107.400 113.210 ;
        RECT 101.575 113.010 107.400 113.150 ;
        RECT 101.575 112.965 101.865 113.010 ;
        RECT 107.080 112.950 107.400 113.010 ;
        RECT 110.300 112.950 110.620 113.210 ;
        RECT 60.635 112.810 60.925 112.855 ;
        RECT 59.700 112.670 60.925 112.810 ;
        RECT 59.700 112.610 60.020 112.670 ;
        RECT 60.635 112.625 60.925 112.670 ;
        RECT 62.935 112.625 63.225 112.855 ;
        RECT 52.800 112.330 54.870 112.470 ;
        RECT 56.020 112.470 56.340 112.530 ;
        RECT 58.335 112.470 58.625 112.515 ;
        RECT 56.020 112.330 58.625 112.470 ;
        RECT 52.800 112.270 53.120 112.330 ;
        RECT 56.020 112.270 56.340 112.330 ;
        RECT 58.335 112.285 58.625 112.330 ;
        RECT 64.315 112.470 64.605 112.515 ;
        RECT 66.600 112.470 66.920 112.530 ;
        RECT 67.475 112.515 67.765 112.830 ;
        RECT 68.555 112.810 68.845 112.855 ;
        RECT 72.135 112.810 72.425 112.855 ;
        RECT 73.970 112.810 74.260 112.855 ;
        RECT 68.555 112.670 74.260 112.810 ;
        RECT 68.555 112.625 68.845 112.670 ;
        RECT 72.135 112.625 72.425 112.670 ;
        RECT 73.970 112.625 74.260 112.670 ;
        RECT 74.420 112.610 74.740 112.870 ;
        RECT 64.315 112.330 66.920 112.470 ;
        RECT 64.315 112.285 64.605 112.330 ;
        RECT 66.600 112.270 66.920 112.330 ;
        RECT 67.175 112.470 67.765 112.515 ;
        RECT 70.280 112.515 70.600 112.530 ;
        RECT 70.280 112.470 71.065 112.515 ;
        RECT 67.175 112.330 71.065 112.470 ;
        RECT 67.175 112.285 67.465 112.330 ;
        RECT 70.280 112.285 71.065 112.330 ;
        RECT 70.280 112.270 70.600 112.285 ;
        RECT 73.040 112.270 73.360 112.530 ;
        RECT 74.880 112.270 75.200 112.530 ;
        RECT 75.800 112.470 76.120 112.530 ;
        RECT 78.055 112.515 78.345 112.830 ;
        RECT 79.135 112.810 79.425 112.855 ;
        RECT 82.715 112.810 83.005 112.855 ;
        RECT 84.550 112.810 84.840 112.855 ;
        RECT 79.135 112.670 84.840 112.810 ;
        RECT 79.135 112.625 79.425 112.670 ;
        RECT 82.715 112.625 83.005 112.670 ;
        RECT 84.550 112.625 84.840 112.670 ;
        RECT 85.920 112.810 86.240 112.870 ;
        RECT 86.395 112.810 86.685 112.855 ;
        RECT 85.920 112.670 86.685 112.810 ;
        RECT 85.920 112.610 86.240 112.670 ;
        RECT 86.395 112.625 86.685 112.670 ;
        RECT 91.855 112.515 92.145 112.830 ;
        RECT 92.935 112.810 93.225 112.855 ;
        RECT 96.515 112.810 96.805 112.855 ;
        RECT 98.350 112.810 98.640 112.855 ;
        RECT 92.935 112.670 98.640 112.810 ;
        RECT 92.935 112.625 93.225 112.670 ;
        RECT 96.515 112.625 96.805 112.670 ;
        RECT 98.350 112.625 98.640 112.670 ;
        RECT 98.815 112.810 99.105 112.855 ;
        RECT 99.720 112.810 100.040 112.870 ;
        RECT 98.815 112.670 100.040 112.810 ;
        RECT 98.815 112.625 99.105 112.670 ;
        RECT 99.720 112.610 100.040 112.670 ;
        RECT 100.195 112.625 100.485 112.855 ;
        RECT 104.780 112.830 105.100 112.870 ;
        RECT 95.120 112.515 95.440 112.530 ;
        RECT 77.755 112.470 78.345 112.515 ;
        RECT 80.995 112.470 81.645 112.515 ;
        RECT 75.800 112.330 81.645 112.470 ;
        RECT 75.800 112.270 76.120 112.330 ;
        RECT 77.755 112.285 78.045 112.330 ;
        RECT 80.995 112.285 81.645 112.330 ;
        RECT 91.555 112.470 92.145 112.515 ;
        RECT 94.795 112.470 95.445 112.515 ;
        RECT 91.555 112.330 95.445 112.470 ;
        RECT 91.555 112.285 91.845 112.330 ;
        RECT 94.795 112.285 95.445 112.330 ;
        RECT 97.420 112.470 97.740 112.530 ;
        RECT 100.270 112.470 100.410 112.625 ;
        RECT 104.735 112.610 105.100 112.830 ;
        RECT 105.815 112.810 106.105 112.855 ;
        RECT 109.395 112.810 109.685 112.855 ;
        RECT 111.230 112.810 111.520 112.855 ;
        RECT 105.815 112.670 111.520 112.810 ;
        RECT 105.815 112.625 106.105 112.670 ;
        RECT 109.395 112.625 109.685 112.670 ;
        RECT 111.230 112.625 111.520 112.670 ;
        RECT 111.680 112.610 112.000 112.870 ;
        RECT 104.735 112.515 105.025 112.610 ;
        RECT 97.420 112.330 100.410 112.470 ;
        RECT 104.435 112.470 105.025 112.515 ;
        RECT 107.675 112.470 108.325 112.515 ;
        RECT 104.435 112.330 108.325 112.470 ;
        RECT 95.120 112.270 95.440 112.285 ;
        RECT 97.420 112.270 97.740 112.330 ;
        RECT 104.435 112.285 104.725 112.330 ;
        RECT 107.675 112.285 108.325 112.330 ;
        RECT 35.780 112.130 36.100 112.190 ;
        RECT 37.635 112.130 37.925 112.175 ;
        RECT 35.780 111.990 37.925 112.130 ;
        RECT 35.780 111.930 36.100 111.990 ;
        RECT 37.635 111.945 37.925 111.990 ;
        RECT 43.155 112.130 43.445 112.175 ;
        RECT 45.440 112.130 45.760 112.190 ;
        RECT 43.155 111.990 45.760 112.130 ;
        RECT 43.155 111.945 43.445 111.990 ;
        RECT 45.440 111.930 45.760 111.990 ;
        RECT 55.115 112.130 55.405 112.175 ;
        RECT 56.480 112.130 56.800 112.190 ;
        RECT 55.115 111.990 56.800 112.130 ;
        RECT 55.115 111.945 55.405 111.990 ;
        RECT 56.480 111.930 56.800 111.990 ;
        RECT 56.955 112.130 57.245 112.175 ;
        RECT 59.240 112.130 59.560 112.190 ;
        RECT 56.955 111.990 59.560 112.130 ;
        RECT 56.955 111.945 57.245 111.990 ;
        RECT 59.240 111.930 59.560 111.990 ;
        RECT 59.700 111.930 60.020 112.190 ;
        RECT 63.855 112.130 64.145 112.175 ;
        RECT 68.440 112.130 68.760 112.190 ;
        RECT 63.855 111.990 68.760 112.130 ;
        RECT 63.855 111.945 64.145 111.990 ;
        RECT 68.440 111.930 68.760 111.990 ;
        RECT 85.000 112.130 85.320 112.190 ;
        RECT 85.475 112.130 85.765 112.175 ;
        RECT 85.000 111.990 85.765 112.130 ;
        RECT 85.000 111.930 85.320 111.990 ;
        RECT 85.475 111.945 85.765 111.990 ;
        RECT 98.340 112.130 98.660 112.190 ;
        RECT 99.275 112.130 99.565 112.175 ;
        RECT 98.340 111.990 99.565 112.130 ;
        RECT 98.340 111.930 98.660 111.990 ;
        RECT 99.275 111.945 99.565 111.990 ;
        RECT 15.010 111.310 113.450 111.790 ;
        RECT 20.600 110.910 20.920 111.170 ;
        RECT 21.520 111.110 21.840 111.170 ;
        RECT 21.995 111.110 22.285 111.155 ;
        RECT 21.520 110.970 22.285 111.110 ;
        RECT 21.520 110.910 21.840 110.970 ;
        RECT 21.995 110.925 22.285 110.970 ;
        RECT 25.200 110.910 25.520 111.170 ;
        RECT 38.080 111.110 38.400 111.170 ;
        RECT 28.510 110.970 38.400 111.110 ;
        RECT 28.510 110.770 28.650 110.970 ;
        RECT 38.080 110.910 38.400 110.970 ;
        RECT 73.040 110.910 73.360 111.170 ;
        RECT 90.520 111.110 90.840 111.170 ;
        RECT 95.120 111.110 95.440 111.170 ;
        RECT 96.515 111.110 96.805 111.155 ;
        RECT 90.520 110.970 94.430 111.110 ;
        RECT 90.520 110.910 90.840 110.970 ;
        RECT 24.830 110.630 28.650 110.770 ;
        RECT 28.895 110.770 29.185 110.815 ;
        RECT 30.260 110.770 30.580 110.830 ;
        RECT 28.895 110.630 30.580 110.770 ;
        RECT 24.830 110.475 24.970 110.630 ;
        RECT 28.895 110.585 29.185 110.630 ;
        RECT 30.260 110.570 30.580 110.630 ;
        RECT 31.175 110.770 31.825 110.815 ;
        RECT 34.775 110.770 35.065 110.815 ;
        RECT 35.780 110.770 36.100 110.830 ;
        RECT 31.175 110.630 36.100 110.770 ;
        RECT 31.175 110.585 31.825 110.630 ;
        RECT 34.475 110.585 35.065 110.630 ;
        RECT 21.075 110.430 21.365 110.475 ;
        RECT 21.535 110.430 21.825 110.475 ;
        RECT 23.375 110.430 23.665 110.475 ;
        RECT 24.755 110.430 25.045 110.475 ;
        RECT 21.075 110.290 25.045 110.430 ;
        RECT 21.075 110.245 21.365 110.290 ;
        RECT 21.535 110.245 21.825 110.290 ;
        RECT 23.375 110.245 23.665 110.290 ;
        RECT 24.755 110.245 25.045 110.290 ;
        RECT 26.120 110.230 26.440 110.490 ;
        RECT 27.980 110.430 28.270 110.475 ;
        RECT 29.815 110.430 30.105 110.475 ;
        RECT 33.395 110.430 33.685 110.475 ;
        RECT 27.980 110.290 33.685 110.430 ;
        RECT 27.980 110.245 28.270 110.290 ;
        RECT 29.815 110.245 30.105 110.290 ;
        RECT 33.395 110.245 33.685 110.290 ;
        RECT 34.475 110.270 34.765 110.585 ;
        RECT 35.780 110.570 36.100 110.630 ;
        RECT 40.955 110.770 41.245 110.815 ;
        RECT 41.760 110.770 42.080 110.830 ;
        RECT 44.195 110.770 44.845 110.815 ;
        RECT 40.955 110.630 44.845 110.770 ;
        RECT 40.955 110.585 41.545 110.630 ;
        RECT 41.255 110.270 41.545 110.585 ;
        RECT 41.760 110.570 42.080 110.630 ;
        RECT 44.195 110.585 44.845 110.630 ;
        RECT 45.440 110.770 45.760 110.830 ;
        RECT 46.835 110.770 47.125 110.815 ;
        RECT 45.440 110.630 47.125 110.770 ;
        RECT 45.440 110.570 45.760 110.630 ;
        RECT 46.835 110.585 47.125 110.630 ;
        RECT 50.040 110.770 50.360 110.830 ;
        RECT 51.995 110.770 52.285 110.815 ;
        RECT 55.235 110.770 55.885 110.815 ;
        RECT 50.040 110.630 55.885 110.770 ;
        RECT 50.040 110.570 50.360 110.630 ;
        RECT 51.995 110.585 52.585 110.630 ;
        RECT 55.235 110.585 55.885 110.630 ;
        RECT 56.480 110.770 56.800 110.830 ;
        RECT 57.875 110.770 58.165 110.815 ;
        RECT 56.480 110.630 58.165 110.770 ;
        RECT 42.335 110.430 42.625 110.475 ;
        RECT 45.915 110.430 46.205 110.475 ;
        RECT 47.750 110.430 48.040 110.475 ;
        RECT 42.335 110.290 48.040 110.430 ;
        RECT 42.335 110.245 42.625 110.290 ;
        RECT 45.915 110.245 46.205 110.290 ;
        RECT 47.750 110.245 48.040 110.290 ;
        RECT 48.215 110.430 48.505 110.475 ;
        RECT 48.660 110.430 48.980 110.490 ;
        RECT 48.215 110.290 48.980 110.430 ;
        RECT 48.215 110.245 48.505 110.290 ;
        RECT 48.660 110.230 48.980 110.290 ;
        RECT 49.135 110.430 49.425 110.475 ;
        RECT 51.420 110.430 51.740 110.490 ;
        RECT 49.135 110.290 51.740 110.430 ;
        RECT 49.135 110.245 49.425 110.290 ;
        RECT 51.420 110.230 51.740 110.290 ;
        RECT 52.295 110.270 52.585 110.585 ;
        RECT 56.480 110.570 56.800 110.630 ;
        RECT 57.875 110.585 58.165 110.630 ;
        RECT 59.240 110.770 59.560 110.830 ;
        RECT 62.575 110.770 62.865 110.815 ;
        RECT 65.815 110.770 66.465 110.815 ;
        RECT 59.240 110.630 66.465 110.770 ;
        RECT 59.240 110.570 59.560 110.630 ;
        RECT 62.575 110.585 63.165 110.630 ;
        RECT 65.815 110.585 66.465 110.630 ;
        RECT 53.375 110.430 53.665 110.475 ;
        RECT 56.955 110.430 57.245 110.475 ;
        RECT 58.790 110.430 59.080 110.475 ;
        RECT 53.375 110.290 59.080 110.430 ;
        RECT 53.375 110.245 53.665 110.290 ;
        RECT 56.955 110.245 57.245 110.290 ;
        RECT 58.790 110.245 59.080 110.290 ;
        RECT 59.715 110.430 60.005 110.475 ;
        RECT 61.540 110.430 61.860 110.490 ;
        RECT 59.715 110.290 61.860 110.430 ;
        RECT 59.715 110.245 60.005 110.290 ;
        RECT 61.540 110.230 61.860 110.290 ;
        RECT 62.875 110.270 63.165 110.585 ;
        RECT 68.440 110.570 68.760 110.830 ;
        RECT 74.420 110.770 74.740 110.830 ;
        RECT 69.910 110.630 74.740 110.770 ;
        RECT 69.910 110.475 70.050 110.630 ;
        RECT 74.420 110.570 74.740 110.630 ;
        RECT 74.895 110.770 75.185 110.815 ;
        RECT 75.340 110.770 75.660 110.830 ;
        RECT 74.895 110.630 75.660 110.770 ;
        RECT 74.895 110.585 75.185 110.630 ;
        RECT 75.340 110.570 75.660 110.630 ;
        RECT 77.755 110.770 78.045 110.815 ;
        RECT 80.995 110.770 81.645 110.815 ;
        RECT 77.755 110.630 81.645 110.770 ;
        RECT 77.755 110.585 78.345 110.630 ;
        RECT 80.995 110.585 81.645 110.630 ;
        RECT 85.475 110.770 85.765 110.815 ;
        RECT 86.380 110.770 86.700 110.830 ;
        RECT 94.290 110.815 94.430 110.970 ;
        RECT 95.120 110.970 96.805 111.110 ;
        RECT 95.120 110.910 95.440 110.970 ;
        RECT 96.515 110.925 96.805 110.970 ;
        RECT 100.180 111.110 100.500 111.170 ;
        RECT 100.180 110.970 109.610 111.110 ;
        RECT 100.180 110.910 100.500 110.970 ;
        RECT 109.470 110.815 109.610 110.970 ;
        RECT 85.475 110.630 86.700 110.770 ;
        RECT 85.475 110.585 85.765 110.630 ;
        RECT 63.955 110.430 64.245 110.475 ;
        RECT 67.535 110.430 67.825 110.475 ;
        RECT 69.370 110.430 69.660 110.475 ;
        RECT 63.955 110.290 69.660 110.430 ;
        RECT 63.955 110.245 64.245 110.290 ;
        RECT 67.535 110.245 67.825 110.290 ;
        RECT 69.370 110.245 69.660 110.290 ;
        RECT 69.835 110.245 70.125 110.475 ;
        RECT 70.755 110.430 71.045 110.475 ;
        RECT 71.660 110.430 71.980 110.490 ;
        RECT 70.755 110.290 71.980 110.430 ;
        RECT 70.755 110.245 71.045 110.290 ;
        RECT 71.660 110.230 71.980 110.290 ;
        RECT 72.120 110.230 72.440 110.490 ;
        RECT 73.040 110.430 73.360 110.490 ;
        RECT 78.055 110.430 78.345 110.585 ;
        RECT 86.380 110.570 86.700 110.630 ;
        RECT 88.335 110.770 88.625 110.815 ;
        RECT 91.575 110.770 92.225 110.815 ;
        RECT 88.335 110.630 92.225 110.770 ;
        RECT 88.335 110.585 88.925 110.630 ;
        RECT 91.575 110.585 92.225 110.630 ;
        RECT 94.215 110.585 94.505 110.815 ;
        RECT 99.275 110.770 99.565 110.815 ;
        RECT 103.515 110.770 103.805 110.815 ;
        RECT 106.755 110.770 107.405 110.815 ;
        RECT 99.275 110.630 107.405 110.770 ;
        RECT 99.275 110.585 99.565 110.630 ;
        RECT 103.515 110.585 104.105 110.630 ;
        RECT 106.755 110.585 107.405 110.630 ;
        RECT 109.395 110.585 109.685 110.815 ;
        RECT 88.635 110.490 88.925 110.585 ;
        RECT 73.040 110.290 78.345 110.430 ;
        RECT 73.040 110.230 73.360 110.290 ;
        RECT 78.055 110.270 78.345 110.290 ;
        RECT 79.135 110.430 79.425 110.475 ;
        RECT 82.715 110.430 83.005 110.475 ;
        RECT 84.550 110.430 84.840 110.475 ;
        RECT 79.135 110.290 84.840 110.430 ;
        RECT 79.135 110.245 79.425 110.290 ;
        RECT 82.715 110.245 83.005 110.290 ;
        RECT 84.550 110.245 84.840 110.290 ;
        RECT 88.635 110.270 89.000 110.490 ;
        RECT 88.680 110.230 89.000 110.270 ;
        RECT 89.715 110.430 90.005 110.475 ;
        RECT 93.295 110.430 93.585 110.475 ;
        RECT 95.130 110.430 95.420 110.475 ;
        RECT 89.715 110.290 95.420 110.430 ;
        RECT 89.715 110.245 90.005 110.290 ;
        RECT 93.295 110.245 93.585 110.290 ;
        RECT 95.130 110.245 95.420 110.290 ;
        RECT 96.040 110.430 96.360 110.490 ;
        RECT 96.975 110.430 97.265 110.475 ;
        RECT 98.355 110.430 98.645 110.475 ;
        RECT 98.815 110.430 99.105 110.475 ;
        RECT 96.040 110.290 100.410 110.430 ;
        RECT 96.040 110.230 96.360 110.290 ;
        RECT 96.975 110.245 97.265 110.290 ;
        RECT 98.355 110.245 98.645 110.290 ;
        RECT 98.815 110.245 99.105 110.290 ;
        RECT 27.515 110.090 27.805 110.135 ;
        RECT 29.340 110.090 29.660 110.150 ;
        RECT 27.515 109.950 29.660 110.090 ;
        RECT 27.515 109.905 27.805 109.950 ;
        RECT 29.340 109.890 29.660 109.950 ;
        RECT 36.240 110.090 36.560 110.150 ;
        RECT 37.635 110.090 37.925 110.135 ;
        RECT 36.240 109.950 37.925 110.090 ;
        RECT 36.240 109.890 36.560 109.950 ;
        RECT 37.635 109.905 37.925 109.950 ;
        RECT 38.095 109.905 38.385 110.135 ;
        RECT 48.750 110.090 48.890 110.230 ;
        RECT 59.255 110.090 59.545 110.135 ;
        RECT 61.080 110.090 61.400 110.150 ;
        RECT 83.635 110.090 83.925 110.135 ;
        RECT 48.750 109.950 61.400 110.090 ;
        RECT 59.255 109.905 59.545 109.950 ;
        RECT 28.385 109.750 28.675 109.795 ;
        RECT 30.275 109.750 30.565 109.795 ;
        RECT 33.395 109.750 33.685 109.795 ;
        RECT 28.385 109.610 33.685 109.750 ;
        RECT 38.170 109.750 38.310 109.905 ;
        RECT 61.080 109.890 61.400 109.950 ;
        RECT 71.750 109.950 83.925 110.090 ;
        RECT 41.300 109.750 41.620 109.810 ;
        RECT 71.750 109.795 71.890 109.950 ;
        RECT 83.635 109.905 83.925 109.950 ;
        RECT 85.015 110.090 85.305 110.135 ;
        RECT 85.460 110.090 85.780 110.150 ;
        RECT 85.015 109.950 85.780 110.090 ;
        RECT 85.015 109.905 85.305 109.950 ;
        RECT 85.460 109.890 85.780 109.950 ;
        RECT 86.840 110.090 87.160 110.150 ;
        RECT 95.595 110.090 95.885 110.135 ;
        RECT 99.720 110.090 100.040 110.150 ;
        RECT 86.840 109.950 100.040 110.090 ;
        RECT 86.840 109.890 87.160 109.950 ;
        RECT 95.595 109.905 95.885 109.950 ;
        RECT 99.720 109.890 100.040 109.950 ;
        RECT 38.170 109.610 41.620 109.750 ;
        RECT 28.385 109.565 28.675 109.610 ;
        RECT 30.275 109.565 30.565 109.610 ;
        RECT 33.395 109.565 33.685 109.610 ;
        RECT 41.300 109.550 41.620 109.610 ;
        RECT 42.335 109.750 42.625 109.795 ;
        RECT 45.455 109.750 45.745 109.795 ;
        RECT 47.345 109.750 47.635 109.795 ;
        RECT 42.335 109.610 47.635 109.750 ;
        RECT 42.335 109.565 42.625 109.610 ;
        RECT 45.455 109.565 45.745 109.610 ;
        RECT 47.345 109.565 47.635 109.610 ;
        RECT 53.375 109.750 53.665 109.795 ;
        RECT 56.495 109.750 56.785 109.795 ;
        RECT 58.385 109.750 58.675 109.795 ;
        RECT 53.375 109.610 58.675 109.750 ;
        RECT 53.375 109.565 53.665 109.610 ;
        RECT 56.495 109.565 56.785 109.610 ;
        RECT 58.385 109.565 58.675 109.610 ;
        RECT 63.955 109.750 64.245 109.795 ;
        RECT 67.075 109.750 67.365 109.795 ;
        RECT 68.965 109.750 69.255 109.795 ;
        RECT 63.955 109.610 69.255 109.750 ;
        RECT 63.955 109.565 64.245 109.610 ;
        RECT 67.075 109.565 67.365 109.610 ;
        RECT 68.965 109.565 69.255 109.610 ;
        RECT 71.675 109.565 71.965 109.795 ;
        RECT 79.135 109.750 79.425 109.795 ;
        RECT 82.255 109.750 82.545 109.795 ;
        RECT 84.145 109.750 84.435 109.795 ;
        RECT 79.135 109.610 84.435 109.750 ;
        RECT 79.135 109.565 79.425 109.610 ;
        RECT 82.255 109.565 82.545 109.610 ;
        RECT 84.145 109.565 84.435 109.610 ;
        RECT 89.715 109.750 90.005 109.795 ;
        RECT 92.835 109.750 93.125 109.795 ;
        RECT 94.725 109.750 95.015 109.795 ;
        RECT 89.715 109.610 95.015 109.750 ;
        RECT 89.715 109.565 90.005 109.610 ;
        RECT 92.835 109.565 93.125 109.610 ;
        RECT 94.725 109.565 95.015 109.610 ;
        RECT 23.820 109.210 24.140 109.470 ;
        RECT 27.040 109.210 27.360 109.470 ;
        RECT 97.880 109.210 98.200 109.470 ;
        RECT 100.270 109.410 100.410 110.290 ;
        RECT 103.815 110.270 104.105 110.585 ;
        RECT 104.895 110.430 105.185 110.475 ;
        RECT 108.475 110.430 108.765 110.475 ;
        RECT 110.310 110.430 110.600 110.475 ;
        RECT 104.895 110.290 110.600 110.430 ;
        RECT 104.895 110.245 105.185 110.290 ;
        RECT 108.475 110.245 108.765 110.290 ;
        RECT 110.310 110.245 110.600 110.290 ;
        RECT 100.640 109.890 100.960 110.150 ;
        RECT 106.160 110.090 106.480 110.150 ;
        RECT 110.775 110.090 111.065 110.135 ;
        RECT 111.680 110.090 112.000 110.150 ;
        RECT 106.160 109.950 112.000 110.090 ;
        RECT 106.160 109.890 106.480 109.950 ;
        RECT 110.775 109.905 111.065 109.950 ;
        RECT 111.680 109.890 112.000 109.950 ;
        RECT 104.895 109.750 105.185 109.795 ;
        RECT 108.015 109.750 108.305 109.795 ;
        RECT 109.905 109.750 110.195 109.795 ;
        RECT 104.895 109.610 110.195 109.750 ;
        RECT 104.895 109.565 105.185 109.610 ;
        RECT 108.015 109.565 108.305 109.610 ;
        RECT 109.905 109.565 110.195 109.610 ;
        RECT 106.620 109.410 106.940 109.470 ;
        RECT 100.270 109.270 106.940 109.410 ;
        RECT 106.620 109.210 106.940 109.270 ;
        RECT 15.010 108.590 113.450 109.070 ;
        RECT 41.760 108.390 42.080 108.450 ;
        RECT 42.695 108.390 42.985 108.435 ;
        RECT 41.760 108.250 42.985 108.390 ;
        RECT 41.760 108.190 42.080 108.250 ;
        RECT 42.695 108.205 42.985 108.250 ;
        RECT 46.820 108.390 47.140 108.450 ;
        RECT 47.755 108.390 48.045 108.435 ;
        RECT 46.820 108.250 48.045 108.390 ;
        RECT 46.820 108.190 47.140 108.250 ;
        RECT 47.755 108.205 48.045 108.250 ;
        RECT 50.040 108.190 50.360 108.450 ;
        RECT 70.280 108.390 70.600 108.450 ;
        RECT 71.215 108.390 71.505 108.435 ;
        RECT 70.280 108.250 71.505 108.390 ;
        RECT 70.280 108.190 70.600 108.250 ;
        RECT 71.215 108.205 71.505 108.250 ;
        RECT 73.040 108.190 73.360 108.450 ;
        RECT 75.800 108.190 76.120 108.450 ;
        RECT 76.350 108.250 87.990 108.390 ;
        RECT 27.615 108.050 27.905 108.095 ;
        RECT 30.735 108.050 31.025 108.095 ;
        RECT 32.625 108.050 32.915 108.095 ;
        RECT 27.615 107.910 32.915 108.050 ;
        RECT 27.615 107.865 27.905 107.910 ;
        RECT 30.735 107.865 31.025 107.910 ;
        RECT 32.625 107.865 32.915 107.910 ;
        RECT 55.215 108.050 55.505 108.095 ;
        RECT 58.335 108.050 58.625 108.095 ;
        RECT 60.225 108.050 60.515 108.095 ;
        RECT 55.215 107.910 60.515 108.050 ;
        RECT 55.215 107.865 55.505 107.910 ;
        RECT 58.335 107.865 58.625 107.910 ;
        RECT 60.225 107.865 60.515 107.910 ;
        RECT 71.660 108.050 71.980 108.110 ;
        RECT 75.340 108.050 75.660 108.110 ;
        RECT 71.660 107.910 75.660 108.050 ;
        RECT 71.660 107.850 71.980 107.910 ;
        RECT 75.340 107.850 75.660 107.910 ;
        RECT 23.375 107.710 23.665 107.755 ;
        RECT 26.120 107.710 26.440 107.770 ;
        RECT 23.375 107.570 26.440 107.710 ;
        RECT 23.375 107.525 23.665 107.570 ;
        RECT 26.120 107.510 26.440 107.570 ;
        RECT 27.040 107.710 27.360 107.770 ;
        RECT 32.115 107.710 32.405 107.755 ;
        RECT 27.040 107.570 32.405 107.710 ;
        RECT 27.040 107.510 27.360 107.570 ;
        RECT 32.115 107.525 32.405 107.570 ;
        RECT 33.495 107.710 33.785 107.755 ;
        RECT 35.320 107.710 35.640 107.770 ;
        RECT 33.495 107.570 35.640 107.710 ;
        RECT 33.495 107.525 33.785 107.570 ;
        RECT 35.320 107.510 35.640 107.570 ;
        RECT 50.975 107.710 51.265 107.755 ;
        RECT 56.480 107.710 56.800 107.770 ;
        RECT 50.975 107.570 56.800 107.710 ;
        RECT 50.975 107.525 51.265 107.570 ;
        RECT 56.480 107.510 56.800 107.570 ;
        RECT 59.700 107.510 60.020 107.770 ;
        RECT 61.080 107.510 61.400 107.770 ;
        RECT 70.740 107.710 71.060 107.770 ;
        RECT 76.350 107.710 76.490 108.250 ;
        RECT 80.975 108.050 81.265 108.095 ;
        RECT 84.095 108.050 84.385 108.095 ;
        RECT 85.985 108.050 86.275 108.095 ;
        RECT 80.975 107.910 86.275 108.050 ;
        RECT 87.850 108.050 87.990 108.250 ;
        RECT 88.680 108.190 89.000 108.450 ;
        RECT 104.780 108.390 105.100 108.450 ;
        RECT 106.175 108.390 106.465 108.435 ;
        RECT 93.370 108.250 99.490 108.390 ;
        RECT 93.370 108.050 93.510 108.250 ;
        RECT 87.850 107.910 93.510 108.050 ;
        RECT 93.855 108.050 94.145 108.095 ;
        RECT 96.975 108.050 97.265 108.095 ;
        RECT 98.865 108.050 99.155 108.095 ;
        RECT 93.855 107.910 99.155 108.050 ;
        RECT 99.350 108.050 99.490 108.250 ;
        RECT 104.780 108.250 106.465 108.390 ;
        RECT 104.780 108.190 105.100 108.250 ;
        RECT 106.175 108.205 106.465 108.250 ;
        RECT 110.775 108.050 111.065 108.095 ;
        RECT 99.350 107.910 111.065 108.050 ;
        RECT 80.975 107.865 81.265 107.910 ;
        RECT 84.095 107.865 84.385 107.910 ;
        RECT 85.985 107.865 86.275 107.910 ;
        RECT 93.855 107.865 94.145 107.910 ;
        RECT 96.975 107.865 97.265 107.910 ;
        RECT 98.865 107.865 99.155 107.910 ;
        RECT 110.775 107.865 111.065 107.910 ;
        RECT 70.740 107.570 76.490 107.710 ;
        RECT 76.735 107.710 77.025 107.755 ;
        RECT 81.780 107.710 82.100 107.770 ;
        RECT 76.735 107.570 82.100 107.710 ;
        RECT 70.740 107.510 71.060 107.570 ;
        RECT 76.735 107.525 77.025 107.570 ;
        RECT 81.780 107.510 82.100 107.570 ;
        RECT 85.000 107.710 85.320 107.770 ;
        RECT 85.475 107.710 85.765 107.755 ;
        RECT 85.000 107.570 85.765 107.710 ;
        RECT 85.000 107.510 85.320 107.570 ;
        RECT 85.475 107.525 85.765 107.570 ;
        RECT 86.840 107.510 87.160 107.770 ;
        RECT 96.040 107.710 96.360 107.770 ;
        RECT 88.310 107.570 96.360 107.710 ;
        RECT 23.820 107.030 24.140 107.090 ;
        RECT 26.535 107.075 26.825 107.390 ;
        RECT 27.615 107.370 27.905 107.415 ;
        RECT 31.195 107.370 31.485 107.415 ;
        RECT 33.030 107.370 33.320 107.415 ;
        RECT 27.615 107.230 33.320 107.370 ;
        RECT 27.615 107.185 27.905 107.230 ;
        RECT 31.195 107.185 31.485 107.230 ;
        RECT 33.030 107.185 33.320 107.230 ;
        RECT 38.080 107.370 38.400 107.430 ;
        RECT 43.155 107.370 43.445 107.415 ;
        RECT 47.295 107.370 47.585 107.415 ;
        RECT 49.595 107.370 49.885 107.415 ;
        RECT 52.800 107.370 53.120 107.430 ;
        RECT 88.310 107.415 88.450 107.570 ;
        RECT 96.040 107.510 96.360 107.570 ;
        RECT 98.340 107.510 98.660 107.770 ;
        RECT 99.720 107.710 100.040 107.770 ;
        RECT 106.160 107.710 106.480 107.770 ;
        RECT 99.720 107.570 106.480 107.710 ;
        RECT 99.720 107.510 100.040 107.570 ;
        RECT 106.160 107.510 106.480 107.570 ;
        RECT 38.080 107.230 53.120 107.370 ;
        RECT 38.080 107.170 38.400 107.230 ;
        RECT 43.155 107.185 43.445 107.230 ;
        RECT 47.295 107.185 47.585 107.230 ;
        RECT 49.595 107.185 49.885 107.230 ;
        RECT 52.800 107.170 53.120 107.230 ;
        RECT 54.135 107.075 54.425 107.390 ;
        RECT 55.215 107.370 55.505 107.415 ;
        RECT 58.795 107.370 59.085 107.415 ;
        RECT 60.630 107.370 60.920 107.415 ;
        RECT 55.215 107.230 60.920 107.370 ;
        RECT 55.215 107.185 55.505 107.230 ;
        RECT 58.795 107.185 59.085 107.230 ;
        RECT 60.630 107.185 60.920 107.230 ;
        RECT 71.675 107.370 71.965 107.415 ;
        RECT 72.595 107.370 72.885 107.415 ;
        RECT 75.355 107.370 75.645 107.415 ;
        RECT 71.675 107.230 79.250 107.370 ;
        RECT 71.675 107.185 71.965 107.230 ;
        RECT 72.595 107.185 72.885 107.230 ;
        RECT 75.355 107.185 75.645 107.230 ;
        RECT 26.235 107.030 26.825 107.075 ;
        RECT 29.475 107.030 30.125 107.075 ;
        RECT 23.820 106.890 30.125 107.030 ;
        RECT 23.820 106.830 24.140 106.890 ;
        RECT 26.235 106.845 26.525 106.890 ;
        RECT 29.475 106.845 30.125 106.890 ;
        RECT 53.835 107.030 54.425 107.075 ;
        RECT 56.020 107.030 56.340 107.090 ;
        RECT 57.075 107.030 57.725 107.075 ;
        RECT 53.835 106.890 57.725 107.030 ;
        RECT 53.835 106.845 54.125 106.890 ;
        RECT 56.020 106.830 56.340 106.890 ;
        RECT 57.075 106.845 57.725 106.890 ;
        RECT 79.110 106.690 79.250 107.230 ;
        RECT 79.895 107.075 80.185 107.390 ;
        RECT 80.975 107.370 81.265 107.415 ;
        RECT 84.555 107.370 84.845 107.415 ;
        RECT 86.390 107.370 86.680 107.415 ;
        RECT 80.975 107.230 86.680 107.370 ;
        RECT 80.975 107.185 81.265 107.230 ;
        RECT 84.555 107.185 84.845 107.230 ;
        RECT 86.390 107.185 86.680 107.230 ;
        RECT 88.235 107.185 88.525 107.415 ;
        RECT 83.160 107.075 83.480 107.090 ;
        RECT 79.595 107.030 80.185 107.075 ;
        RECT 82.835 107.030 83.485 107.075 ;
        RECT 79.595 106.890 83.485 107.030 ;
        RECT 79.595 106.845 79.885 106.890 ;
        RECT 82.835 106.845 83.485 106.890 ;
        RECT 84.080 107.030 84.400 107.090 ;
        RECT 88.310 107.030 88.450 107.185 ;
        RECT 92.775 107.075 93.065 107.390 ;
        RECT 93.855 107.370 94.145 107.415 ;
        RECT 97.435 107.370 97.725 107.415 ;
        RECT 99.270 107.370 99.560 107.415 ;
        RECT 93.855 107.230 99.560 107.370 ;
        RECT 93.855 107.185 94.145 107.230 ;
        RECT 97.435 107.185 97.725 107.230 ;
        RECT 99.270 107.185 99.560 107.230 ;
        RECT 106.620 107.170 106.940 107.430 ;
        RECT 111.695 107.370 111.985 107.415 ;
        RECT 116.740 107.370 117.060 107.430 ;
        RECT 111.695 107.230 117.060 107.370 ;
        RECT 111.695 107.185 111.985 107.230 ;
        RECT 116.740 107.170 117.060 107.230 ;
        RECT 84.080 106.890 88.450 107.030 ;
        RECT 83.160 106.830 83.480 106.845 ;
        RECT 84.080 106.830 84.400 106.890 ;
        RECT 89.615 106.845 89.905 107.075 ;
        RECT 92.475 107.030 93.065 107.075 ;
        RECT 95.715 107.030 96.365 107.075 ;
        RECT 97.880 107.030 98.200 107.090 ;
        RECT 92.475 106.890 98.200 107.030 ;
        RECT 92.475 106.845 92.765 106.890 ;
        RECT 95.715 106.845 96.365 106.890 ;
        RECT 84.170 106.690 84.310 106.830 ;
        RECT 79.110 106.550 84.310 106.690 ;
        RECT 89.690 106.690 89.830 106.845 ;
        RECT 97.880 106.830 98.200 106.890 ;
        RECT 96.960 106.690 97.280 106.750 ;
        RECT 135.660 106.690 136.800 133.400 ;
        RECT 89.690 106.550 97.280 106.690 ;
        RECT 133.100 106.600 136.850 106.690 ;
        RECT 96.960 106.490 97.280 106.550 ;
        RECT 15.010 105.870 113.450 106.350 ;
        RECT 129.700 105.630 136.850 106.600 ;
        RECT 133.100 105.500 136.850 105.630 ;
        RECT 133.330 76.630 136.060 77.830 ;
        RECT 137.920 77.810 143.450 77.960 ;
        RECT 21.115 74.380 23.065 74.390 ;
        RECT 19.415 73.240 23.065 74.380 ;
        RECT 19.415 73.230 21.125 73.240 ;
        RECT 28.135 73.230 30.305 74.410 ;
        RECT 32.315 74.390 34.265 74.400 ;
        RECT 30.615 73.250 34.265 74.390 ;
        RECT 30.615 73.240 32.325 73.250 ;
        RECT 39.425 73.200 41.595 74.380 ;
        RECT 43.535 74.360 45.485 74.370 ;
        RECT 41.835 73.220 45.485 74.360 ;
        RECT 54.785 74.340 56.735 74.350 ;
        RECT 41.835 73.210 43.545 73.220 ;
        RECT 3.910 73.080 6.100 73.190 ;
        RECT 50.005 73.140 52.175 74.320 ;
        RECT 53.085 73.200 56.735 74.340 ;
        RECT 53.085 73.190 54.795 73.200 ;
        RECT 61.425 73.170 63.595 74.350 ;
        RECT 66.005 74.330 67.955 74.340 ;
        RECT 64.305 73.190 67.955 74.330 ;
        RECT 64.305 73.180 66.015 73.190 ;
        RECT 72.535 73.180 74.705 74.360 ;
        RECT 77.245 74.320 79.195 74.330 ;
        RECT 75.545 73.180 79.195 74.320 ;
        RECT 75.545 73.170 77.255 73.180 ;
        RECT 83.805 73.170 85.975 74.350 ;
        RECT 88.495 74.330 90.445 74.340 ;
        RECT 86.795 73.190 90.445 74.330 ;
        RECT 99.775 74.320 101.725 74.330 ;
        RECT 86.795 73.180 88.505 73.190 ;
        RECT 94.995 73.110 97.165 74.290 ;
        RECT 98.075 73.180 101.725 74.320 ;
        RECT 98.075 73.170 99.785 73.180 ;
        RECT 106.405 73.160 108.575 74.340 ;
        RECT 111.045 74.320 112.995 74.330 ;
        RECT 109.345 73.180 112.995 74.320 ;
        RECT 109.345 73.170 111.055 73.180 ;
        RECT 117.605 73.160 119.775 74.340 ;
        RECT 122.295 74.320 124.245 74.330 ;
        RECT 120.595 73.180 124.245 74.320 ;
        RECT 129.455 73.240 131.625 74.420 ;
        RECT 120.595 73.170 122.305 73.180 ;
        RECT 3.910 72.820 12.240 73.080 ;
        RECT 29.635 72.840 43.235 72.850 ;
        RECT 18.435 72.820 43.235 72.840 ;
        RECT 3.910 72.800 54.455 72.820 ;
        RECT 3.910 72.790 65.705 72.800 ;
        RECT 133.960 72.790 135.640 76.630 ;
        RECT 137.190 76.610 143.450 77.810 ;
        RECT 137.920 75.460 143.450 76.610 ;
        RECT 3.910 72.780 76.925 72.790 ;
        RECT 85.815 72.780 99.415 72.790 ;
        RECT 132.085 72.780 140.600 72.790 ;
        RECT 3.910 71.700 140.600 72.780 ;
        RECT 3.910 71.690 32.035 71.700 ;
        RECT 3.910 71.670 19.135 71.690 ;
        RECT 40.855 71.670 140.600 71.700 ;
        RECT 3.910 71.500 12.240 71.670 ;
        RECT 52.105 71.650 140.600 71.670 ;
        RECT 63.325 71.640 140.600 71.650 ;
        RECT 74.565 71.630 88.165 71.640 ;
        RECT 97.095 71.630 133.215 71.640 ;
        RECT 3.910 71.370 6.100 71.500 ;
        RECT 10.800 71.180 11.950 71.500 ;
        RECT 10.800 69.480 11.915 71.180 ;
        RECT 29.635 71.170 43.285 71.180 ;
        RECT 15.510 71.155 17.040 71.160 ;
        RECT 18.435 71.155 43.285 71.170 ;
        RECT 12.285 71.150 43.285 71.155 ;
        RECT 12.285 71.130 54.505 71.150 ;
        RECT 141.810 71.140 143.230 75.460 ;
        RECT 12.285 71.120 65.755 71.130 ;
        RECT 12.285 71.110 76.975 71.120 ;
        RECT 85.815 71.110 99.465 71.120 ;
        RECT 140.220 71.110 143.240 71.140 ;
        RECT 12.285 70.030 143.240 71.110 ;
        RECT 12.285 70.020 32.085 70.030 ;
        RECT 12.285 70.005 19.375 70.020 ;
        RECT 10.800 13.800 11.950 69.480 ;
        RECT 12.320 15.450 13.470 70.005 ;
        RECT 15.510 68.660 17.040 70.005 ;
        RECT 40.855 70.000 143.240 70.030 ;
        RECT 52.105 69.980 143.240 70.000 ;
        RECT 63.325 69.970 143.240 69.980 ;
        RECT 74.565 69.960 88.215 69.970 ;
        RECT 97.095 69.960 143.240 69.970 ;
        RECT 140.220 69.910 143.240 69.960 ;
        RECT 29.645 69.670 43.315 69.680 ;
        RECT 18.445 69.650 43.315 69.670 ;
        RECT 18.445 69.630 54.535 69.650 ;
        RECT 18.445 69.620 65.785 69.630 ;
        RECT 139.590 69.620 150.610 69.640 ;
        RECT 18.445 69.610 77.005 69.620 ;
        RECT 85.825 69.610 99.495 69.620 ;
        RECT 132.155 69.610 150.610 69.620 ;
        RECT 18.445 69.570 150.610 69.610 ;
        RECT 18.445 68.530 150.740 69.570 ;
        RECT 18.445 68.520 32.115 68.530 ;
        RECT 40.865 68.500 150.740 68.530 ;
        RECT 52.115 68.490 143.320 68.500 ;
        RECT 52.115 68.480 140.670 68.490 ;
        RECT 63.335 68.470 140.670 68.480 ;
        RECT 74.575 68.460 88.245 68.470 ;
        RECT 97.105 68.460 133.295 68.470 ;
        RECT 141.080 68.450 142.300 68.490 ;
        RECT 149.360 68.470 150.740 68.500 ;
        RECT 29.655 68.100 43.325 68.110 ;
        RECT 13.950 68.080 43.325 68.100 ;
        RECT 13.950 68.060 54.545 68.080 ;
        RECT 13.950 68.050 65.795 68.060 ;
        RECT 13.950 68.040 77.015 68.050 ;
        RECT 85.835 68.040 99.505 68.050 ;
        RECT 139.530 68.040 143.320 68.060 ;
        RECT 13.950 66.960 152.870 68.040 ;
        RECT 13.950 66.950 32.125 66.960 ;
        RECT 13.950 18.530 15.100 66.950 ;
        RECT 40.875 66.930 152.870 66.960 ;
        RECT 52.125 66.910 152.870 66.930 ;
        RECT 63.345 66.900 152.870 66.910 ;
        RECT 74.585 66.890 88.255 66.900 ;
        RECT 97.115 66.890 143.320 66.900 ;
        RECT 141.030 66.770 142.490 66.890 ;
        RECT 21.405 65.510 26.555 65.790 ;
        RECT 27.815 65.490 28.965 65.800 ;
        RECT 32.605 65.520 37.755 65.800 ;
        RECT 39.015 65.500 40.165 65.810 ;
        RECT 43.825 65.490 48.975 65.770 ;
        RECT 50.235 65.470 51.385 65.780 ;
        RECT 149.460 65.760 150.600 65.780 ;
        RECT 55.075 65.470 60.225 65.750 ;
        RECT 61.485 65.450 62.635 65.760 ;
        RECT 66.295 65.460 71.445 65.740 ;
        RECT 72.705 65.440 73.855 65.750 ;
        RECT 77.535 65.450 82.685 65.730 ;
        RECT 83.945 65.430 85.095 65.740 ;
        RECT 88.785 65.460 93.935 65.740 ;
        RECT 95.195 65.440 96.345 65.750 ;
        RECT 100.065 65.450 105.215 65.730 ;
        RECT 106.475 65.430 107.625 65.740 ;
        RECT 111.335 65.450 116.485 65.730 ;
        RECT 117.745 65.430 118.895 65.740 ;
        RECT 122.585 65.450 127.735 65.730 ;
        RECT 128.995 65.430 130.145 65.740 ;
        RECT 133.315 65.430 138.455 65.690 ;
        RECT 21.205 65.140 21.435 65.320 ;
        RECT 26.495 65.190 26.725 65.320 ;
        RECT 21.125 55.220 21.485 65.140 ;
        RECT 26.435 55.240 26.805 65.190 ;
        RECT 27.635 65.150 27.865 65.320 ;
        RECT 27.565 55.200 27.935 65.150 ;
        RECT 28.925 65.140 29.155 65.320 ;
        RECT 32.405 65.150 32.635 65.330 ;
        RECT 37.695 65.200 37.925 65.330 ;
        RECT 28.835 55.250 29.255 65.140 ;
        RECT 32.325 55.230 32.685 65.150 ;
        RECT 37.635 55.250 38.005 65.200 ;
        RECT 38.835 65.160 39.065 65.330 ;
        RECT 38.765 55.210 39.135 65.160 ;
        RECT 40.125 65.150 40.355 65.330 ;
        RECT 40.035 55.260 40.455 65.150 ;
        RECT 43.625 65.120 43.855 65.300 ;
        RECT 48.915 65.170 49.145 65.300 ;
        RECT 43.545 55.200 43.905 65.120 ;
        RECT 48.855 55.220 49.225 65.170 ;
        RECT 50.055 65.130 50.285 65.300 ;
        RECT 49.985 55.180 50.355 65.130 ;
        RECT 51.345 65.120 51.575 65.300 ;
        RECT 51.255 55.230 51.675 65.120 ;
        RECT 54.875 65.100 55.105 65.280 ;
        RECT 60.165 65.150 60.395 65.280 ;
        RECT 54.795 55.180 55.155 65.100 ;
        RECT 60.105 55.200 60.475 65.150 ;
        RECT 61.305 65.110 61.535 65.280 ;
        RECT 61.235 55.160 61.605 65.110 ;
        RECT 62.595 65.100 62.825 65.280 ;
        RECT 62.505 55.210 62.925 65.100 ;
        RECT 66.095 65.090 66.325 65.270 ;
        RECT 71.385 65.140 71.615 65.270 ;
        RECT 66.015 55.170 66.375 65.090 ;
        RECT 71.325 55.190 71.695 65.140 ;
        RECT 72.525 65.100 72.755 65.270 ;
        RECT 72.455 55.150 72.825 65.100 ;
        RECT 73.815 65.090 74.045 65.270 ;
        RECT 73.725 55.200 74.145 65.090 ;
        RECT 77.335 65.080 77.565 65.260 ;
        RECT 82.625 65.130 82.855 65.260 ;
        RECT 77.255 55.160 77.615 65.080 ;
        RECT 82.565 55.180 82.935 65.130 ;
        RECT 83.765 65.090 83.995 65.260 ;
        RECT 83.695 55.140 84.065 65.090 ;
        RECT 85.055 65.080 85.285 65.260 ;
        RECT 88.585 65.090 88.815 65.270 ;
        RECT 93.875 65.140 94.105 65.270 ;
        RECT 84.965 55.190 85.385 65.080 ;
        RECT 88.505 55.170 88.865 65.090 ;
        RECT 93.815 55.190 94.185 65.140 ;
        RECT 95.015 65.100 95.245 65.270 ;
        RECT 94.945 55.150 95.315 65.100 ;
        RECT 96.305 65.090 96.535 65.270 ;
        RECT 96.215 55.200 96.635 65.090 ;
        RECT 99.865 65.080 100.095 65.260 ;
        RECT 105.155 65.130 105.385 65.260 ;
        RECT 99.785 55.160 100.145 65.080 ;
        RECT 105.095 55.180 105.465 65.130 ;
        RECT 106.295 65.090 106.525 65.260 ;
        RECT 106.225 55.140 106.595 65.090 ;
        RECT 107.585 65.080 107.815 65.260 ;
        RECT 111.135 65.080 111.365 65.260 ;
        RECT 116.425 65.130 116.655 65.260 ;
        RECT 107.495 55.190 107.915 65.080 ;
        RECT 111.055 55.160 111.415 65.080 ;
        RECT 116.365 55.180 116.735 65.130 ;
        RECT 117.565 65.090 117.795 65.260 ;
        RECT 117.495 55.140 117.865 65.090 ;
        RECT 118.855 65.080 119.085 65.260 ;
        RECT 122.385 65.080 122.615 65.260 ;
        RECT 127.675 65.130 127.905 65.260 ;
        RECT 118.765 55.190 119.185 65.080 ;
        RECT 122.305 55.160 122.665 65.080 ;
        RECT 127.615 55.180 127.985 65.130 ;
        RECT 128.815 65.090 129.045 65.260 ;
        RECT 128.745 55.140 129.115 65.090 ;
        RECT 130.105 65.080 130.335 65.260 ;
        RECT 133.135 65.130 133.365 65.230 ;
        RECT 130.015 55.190 130.435 65.080 ;
        RECT 133.005 55.240 133.405 65.130 ;
        RECT 138.425 65.100 138.655 65.230 ;
        RECT 133.135 55.230 133.365 55.240 ;
        RECT 138.345 55.130 138.725 65.100 ;
        RECT 149.340 64.660 150.720 65.760 ;
        RECT 20.815 54.230 25.555 54.530 ;
        RECT 32.015 54.240 36.755 54.540 ;
        RECT 43.235 54.210 47.975 54.510 ;
        RECT 54.485 54.190 59.225 54.490 ;
        RECT 65.705 54.180 70.445 54.480 ;
        RECT 76.945 54.170 81.685 54.470 ;
        RECT 88.195 54.180 92.935 54.480 ;
        RECT 99.475 54.170 104.215 54.470 ;
        RECT 110.745 54.170 115.485 54.470 ;
        RECT 121.995 54.170 126.735 54.470 ;
        RECT 21.655 52.320 22.115 52.550 ;
        RECT 25.625 52.280 26.255 52.560 ;
        RECT 25.735 52.240 26.195 52.280 ;
        RECT 27.665 52.240 28.125 52.470 ;
        RECT 32.855 52.330 33.315 52.560 ;
        RECT 36.825 52.290 37.455 52.570 ;
        RECT 36.935 52.250 37.395 52.290 ;
        RECT 38.865 52.250 39.325 52.480 ;
        RECT 44.075 52.300 44.535 52.530 ;
        RECT 48.045 52.260 48.675 52.540 ;
        RECT 48.155 52.220 48.615 52.260 ;
        RECT 50.085 52.220 50.545 52.450 ;
        RECT 55.325 52.280 55.785 52.510 ;
        RECT 59.295 52.240 59.925 52.520 ;
        RECT 59.405 52.200 59.865 52.240 ;
        RECT 61.335 52.200 61.795 52.430 ;
        RECT 66.545 52.270 67.005 52.500 ;
        RECT 70.515 52.230 71.145 52.510 ;
        RECT 70.625 52.190 71.085 52.230 ;
        RECT 72.555 52.190 73.015 52.420 ;
        RECT 77.785 52.260 78.245 52.490 ;
        RECT 81.755 52.220 82.385 52.500 ;
        RECT 81.865 52.180 82.325 52.220 ;
        RECT 83.795 52.180 84.255 52.410 ;
        RECT 89.035 52.270 89.495 52.500 ;
        RECT 93.005 52.230 93.635 52.510 ;
        RECT 93.115 52.190 93.575 52.230 ;
        RECT 95.045 52.190 95.505 52.420 ;
        RECT 100.315 52.260 100.775 52.490 ;
        RECT 104.285 52.220 104.915 52.500 ;
        RECT 104.395 52.180 104.855 52.220 ;
        RECT 106.325 52.180 106.785 52.410 ;
        RECT 111.585 52.260 112.045 52.490 ;
        RECT 115.555 52.220 116.185 52.500 ;
        RECT 115.665 52.180 116.125 52.220 ;
        RECT 117.595 52.180 118.055 52.410 ;
        RECT 122.835 52.260 123.295 52.490 ;
        RECT 126.805 52.220 127.435 52.500 ;
        RECT 126.915 52.180 127.375 52.220 ;
        RECT 128.845 52.180 129.305 52.410 ;
        RECT 21.375 52.010 21.605 52.115 ;
        RECT 21.245 50.290 21.615 52.010 ;
        RECT 22.165 51.890 22.395 52.115 ;
        RECT 25.455 51.980 25.685 52.035 ;
        RECT 21.375 50.115 21.605 50.290 ;
        RECT 22.155 50.210 22.525 51.890 ;
        RECT 22.165 50.115 22.395 50.210 ;
        RECT 21.525 49.670 22.245 49.930 ;
        RECT 19.295 46.650 20.065 47.720 ;
        RECT 21.385 47.490 22.105 47.750 ;
        RECT 21.225 47.200 21.455 47.340 ;
        RECT 21.085 46.430 21.475 47.200 ;
        RECT 22.015 47.190 22.245 47.340 ;
        RECT 22.005 46.450 22.375 47.190 ;
        RECT 25.305 47.010 25.735 51.980 ;
        RECT 26.245 51.970 26.475 52.035 ;
        RECT 27.385 51.970 27.615 52.035 ;
        RECT 26.185 46.970 26.585 51.970 ;
        RECT 27.265 46.970 27.665 51.970 ;
        RECT 28.175 51.940 28.405 52.035 ;
        RECT 32.575 52.020 32.805 52.125 ;
        RECT 28.115 46.970 28.545 51.940 ;
        RECT 32.445 50.300 32.815 52.020 ;
        RECT 33.365 51.900 33.595 52.125 ;
        RECT 36.655 51.990 36.885 52.045 ;
        RECT 32.575 50.125 32.805 50.300 ;
        RECT 33.355 50.220 33.725 51.900 ;
        RECT 33.365 50.125 33.595 50.220 ;
        RECT 32.725 49.680 33.445 49.940 ;
        RECT 25.735 46.600 26.195 46.830 ;
        RECT 27.665 46.710 28.125 46.830 ;
        RECT 27.515 46.600 28.125 46.710 ;
        RECT 30.495 46.660 31.265 47.730 ;
        RECT 32.585 47.500 33.305 47.760 ;
        RECT 32.425 47.210 32.655 47.350 ;
        RECT 21.225 46.340 21.455 46.430 ;
        RECT 22.015 46.340 22.245 46.450 ;
        RECT 27.515 46.430 28.095 46.600 ;
        RECT 32.285 46.440 32.675 47.210 ;
        RECT 33.215 47.200 33.445 47.350 ;
        RECT 33.205 46.460 33.575 47.200 ;
        RECT 36.505 47.020 36.935 51.990 ;
        RECT 37.445 51.980 37.675 52.045 ;
        RECT 38.585 51.980 38.815 52.045 ;
        RECT 37.385 46.980 37.785 51.980 ;
        RECT 38.465 46.980 38.865 51.980 ;
        RECT 39.375 51.950 39.605 52.045 ;
        RECT 43.795 51.990 44.025 52.095 ;
        RECT 39.315 46.980 39.745 51.950 ;
        RECT 43.665 50.270 44.035 51.990 ;
        RECT 44.585 51.870 44.815 52.095 ;
        RECT 47.875 51.960 48.105 52.015 ;
        RECT 43.795 50.095 44.025 50.270 ;
        RECT 44.575 50.190 44.945 51.870 ;
        RECT 44.585 50.095 44.815 50.190 ;
        RECT 43.945 49.650 44.665 49.910 ;
        RECT 36.935 46.610 37.395 46.840 ;
        RECT 38.865 46.720 39.325 46.840 ;
        RECT 38.715 46.610 39.325 46.720 ;
        RECT 41.715 46.630 42.485 47.700 ;
        RECT 43.805 47.470 44.525 47.730 ;
        RECT 43.645 47.180 43.875 47.320 ;
        RECT 32.425 46.350 32.655 46.440 ;
        RECT 33.215 46.350 33.445 46.460 ;
        RECT 38.715 46.440 39.295 46.610 ;
        RECT 43.505 46.410 43.895 47.180 ;
        RECT 44.435 47.170 44.665 47.320 ;
        RECT 44.425 46.430 44.795 47.170 ;
        RECT 47.725 46.990 48.155 51.960 ;
        RECT 48.665 51.950 48.895 52.015 ;
        RECT 49.805 51.950 50.035 52.015 ;
        RECT 48.605 46.950 49.005 51.950 ;
        RECT 49.685 46.950 50.085 51.950 ;
        RECT 50.595 51.920 50.825 52.015 ;
        RECT 55.045 51.970 55.275 52.075 ;
        RECT 50.535 46.950 50.965 51.920 ;
        RECT 54.915 50.250 55.285 51.970 ;
        RECT 55.835 51.850 56.065 52.075 ;
        RECT 59.125 51.940 59.355 51.995 ;
        RECT 55.045 50.075 55.275 50.250 ;
        RECT 55.825 50.170 56.195 51.850 ;
        RECT 55.835 50.075 56.065 50.170 ;
        RECT 55.195 49.630 55.915 49.890 ;
        RECT 48.155 46.580 48.615 46.810 ;
        RECT 50.085 46.690 50.545 46.810 ;
        RECT 49.935 46.580 50.545 46.690 ;
        RECT 52.965 46.610 53.735 47.680 ;
        RECT 55.055 47.450 55.775 47.710 ;
        RECT 54.895 47.160 55.125 47.300 ;
        RECT 43.645 46.320 43.875 46.410 ;
        RECT 44.435 46.320 44.665 46.430 ;
        RECT 49.935 46.410 50.515 46.580 ;
        RECT 54.755 46.390 55.145 47.160 ;
        RECT 55.685 47.150 55.915 47.300 ;
        RECT 55.675 46.410 56.045 47.150 ;
        RECT 58.975 46.970 59.405 51.940 ;
        RECT 59.915 51.930 60.145 51.995 ;
        RECT 61.055 51.930 61.285 51.995 ;
        RECT 59.855 46.930 60.255 51.930 ;
        RECT 60.935 46.930 61.335 51.930 ;
        RECT 61.845 51.900 62.075 51.995 ;
        RECT 66.265 51.960 66.495 52.065 ;
        RECT 61.785 46.930 62.215 51.900 ;
        RECT 66.135 50.240 66.505 51.960 ;
        RECT 67.055 51.840 67.285 52.065 ;
        RECT 70.345 51.930 70.575 51.985 ;
        RECT 66.265 50.065 66.495 50.240 ;
        RECT 67.045 50.160 67.415 51.840 ;
        RECT 67.055 50.065 67.285 50.160 ;
        RECT 66.415 49.620 67.135 49.880 ;
        RECT 59.405 46.560 59.865 46.790 ;
        RECT 61.335 46.670 61.795 46.790 ;
        RECT 61.185 46.560 61.795 46.670 ;
        RECT 64.185 46.600 64.955 47.670 ;
        RECT 66.275 47.440 66.995 47.700 ;
        RECT 66.115 47.150 66.345 47.290 ;
        RECT 54.895 46.300 55.125 46.390 ;
        RECT 55.685 46.300 55.915 46.410 ;
        RECT 61.185 46.390 61.765 46.560 ;
        RECT 65.975 46.380 66.365 47.150 ;
        RECT 66.905 47.140 67.135 47.290 ;
        RECT 66.895 46.400 67.265 47.140 ;
        RECT 70.195 46.960 70.625 51.930 ;
        RECT 71.135 51.920 71.365 51.985 ;
        RECT 72.275 51.920 72.505 51.985 ;
        RECT 71.075 46.920 71.475 51.920 ;
        RECT 72.155 46.920 72.555 51.920 ;
        RECT 73.065 51.890 73.295 51.985 ;
        RECT 77.505 51.950 77.735 52.055 ;
        RECT 73.005 46.920 73.435 51.890 ;
        RECT 77.375 50.230 77.745 51.950 ;
        RECT 78.295 51.830 78.525 52.055 ;
        RECT 81.585 51.920 81.815 51.975 ;
        RECT 77.505 50.055 77.735 50.230 ;
        RECT 78.285 50.150 78.655 51.830 ;
        RECT 78.295 50.055 78.525 50.150 ;
        RECT 77.655 49.610 78.375 49.870 ;
        RECT 70.625 46.550 71.085 46.780 ;
        RECT 72.555 46.660 73.015 46.780 ;
        RECT 72.405 46.550 73.015 46.660 ;
        RECT 75.425 46.590 76.195 47.660 ;
        RECT 77.515 47.430 78.235 47.690 ;
        RECT 77.355 47.140 77.585 47.280 ;
        RECT 66.115 46.290 66.345 46.380 ;
        RECT 66.905 46.290 67.135 46.400 ;
        RECT 72.405 46.380 72.985 46.550 ;
        RECT 77.215 46.370 77.605 47.140 ;
        RECT 78.145 47.130 78.375 47.280 ;
        RECT 78.135 46.390 78.505 47.130 ;
        RECT 81.435 46.950 81.865 51.920 ;
        RECT 82.375 51.910 82.605 51.975 ;
        RECT 83.515 51.910 83.745 51.975 ;
        RECT 82.315 46.910 82.715 51.910 ;
        RECT 83.395 46.910 83.795 51.910 ;
        RECT 84.305 51.880 84.535 51.975 ;
        RECT 88.755 51.960 88.985 52.065 ;
        RECT 84.245 46.910 84.675 51.880 ;
        RECT 88.625 50.240 88.995 51.960 ;
        RECT 89.545 51.840 89.775 52.065 ;
        RECT 92.835 51.930 93.065 51.985 ;
        RECT 88.755 50.065 88.985 50.240 ;
        RECT 89.535 50.160 89.905 51.840 ;
        RECT 89.545 50.065 89.775 50.160 ;
        RECT 88.905 49.620 89.625 49.880 ;
        RECT 81.865 46.540 82.325 46.770 ;
        RECT 83.795 46.650 84.255 46.770 ;
        RECT 83.645 46.540 84.255 46.650 ;
        RECT 86.675 46.600 87.445 47.670 ;
        RECT 88.765 47.440 89.485 47.700 ;
        RECT 88.605 47.150 88.835 47.290 ;
        RECT 77.355 46.280 77.585 46.370 ;
        RECT 78.145 46.280 78.375 46.390 ;
        RECT 83.645 46.370 84.225 46.540 ;
        RECT 88.465 46.380 88.855 47.150 ;
        RECT 89.395 47.140 89.625 47.290 ;
        RECT 89.385 46.400 89.755 47.140 ;
        RECT 92.685 46.960 93.115 51.930 ;
        RECT 93.625 51.920 93.855 51.985 ;
        RECT 94.765 51.920 94.995 51.985 ;
        RECT 93.565 46.920 93.965 51.920 ;
        RECT 94.645 46.920 95.045 51.920 ;
        RECT 95.555 51.890 95.785 51.985 ;
        RECT 100.035 51.950 100.265 52.055 ;
        RECT 95.495 46.920 95.925 51.890 ;
        RECT 99.905 50.230 100.275 51.950 ;
        RECT 100.825 51.830 101.055 52.055 ;
        RECT 104.115 51.920 104.345 51.975 ;
        RECT 100.035 50.055 100.265 50.230 ;
        RECT 100.815 50.150 101.185 51.830 ;
        RECT 100.825 50.055 101.055 50.150 ;
        RECT 100.185 49.610 100.905 49.870 ;
        RECT 93.115 46.550 93.575 46.780 ;
        RECT 95.045 46.660 95.505 46.780 ;
        RECT 94.895 46.550 95.505 46.660 ;
        RECT 97.955 46.590 98.725 47.660 ;
        RECT 100.045 47.430 100.765 47.690 ;
        RECT 99.885 47.140 100.115 47.280 ;
        RECT 88.605 46.290 88.835 46.380 ;
        RECT 89.395 46.290 89.625 46.400 ;
        RECT 94.895 46.380 95.475 46.550 ;
        RECT 99.745 46.370 100.135 47.140 ;
        RECT 100.675 47.130 100.905 47.280 ;
        RECT 100.665 46.390 101.035 47.130 ;
        RECT 103.965 46.950 104.395 51.920 ;
        RECT 104.905 51.910 105.135 51.975 ;
        RECT 106.045 51.910 106.275 51.975 ;
        RECT 104.845 46.910 105.245 51.910 ;
        RECT 105.925 46.910 106.325 51.910 ;
        RECT 106.835 51.880 107.065 51.975 ;
        RECT 111.305 51.950 111.535 52.055 ;
        RECT 106.775 46.910 107.205 51.880 ;
        RECT 111.175 50.230 111.545 51.950 ;
        RECT 112.095 51.830 112.325 52.055 ;
        RECT 115.385 51.920 115.615 51.975 ;
        RECT 111.305 50.055 111.535 50.230 ;
        RECT 112.085 50.150 112.455 51.830 ;
        RECT 112.095 50.055 112.325 50.150 ;
        RECT 111.455 49.610 112.175 49.870 ;
        RECT 104.395 46.540 104.855 46.770 ;
        RECT 106.325 46.650 106.785 46.770 ;
        RECT 106.175 46.540 106.785 46.650 ;
        RECT 109.225 46.590 109.995 47.660 ;
        RECT 111.315 47.430 112.035 47.690 ;
        RECT 111.155 47.140 111.385 47.280 ;
        RECT 99.885 46.280 100.115 46.370 ;
        RECT 100.675 46.280 100.905 46.390 ;
        RECT 106.175 46.370 106.755 46.540 ;
        RECT 111.015 46.370 111.405 47.140 ;
        RECT 111.945 47.130 112.175 47.280 ;
        RECT 111.935 46.390 112.305 47.130 ;
        RECT 115.235 46.950 115.665 51.920 ;
        RECT 116.175 51.910 116.405 51.975 ;
        RECT 117.315 51.910 117.545 51.975 ;
        RECT 116.115 46.910 116.515 51.910 ;
        RECT 117.195 46.910 117.595 51.910 ;
        RECT 118.105 51.880 118.335 51.975 ;
        RECT 122.555 51.950 122.785 52.055 ;
        RECT 118.045 46.910 118.475 51.880 ;
        RECT 122.425 50.230 122.795 51.950 ;
        RECT 123.345 51.830 123.575 52.055 ;
        RECT 126.635 51.920 126.865 51.975 ;
        RECT 122.555 50.055 122.785 50.230 ;
        RECT 123.335 50.150 123.705 51.830 ;
        RECT 123.345 50.055 123.575 50.150 ;
        RECT 122.705 49.610 123.425 49.870 ;
        RECT 115.665 46.540 116.125 46.770 ;
        RECT 117.595 46.650 118.055 46.770 ;
        RECT 117.445 46.540 118.055 46.650 ;
        RECT 120.475 46.590 121.245 47.660 ;
        RECT 122.565 47.430 123.285 47.690 ;
        RECT 122.405 47.140 122.635 47.280 ;
        RECT 111.155 46.280 111.385 46.370 ;
        RECT 111.945 46.280 112.175 46.390 ;
        RECT 117.445 46.370 118.025 46.540 ;
        RECT 122.265 46.370 122.655 47.140 ;
        RECT 123.195 47.130 123.425 47.280 ;
        RECT 123.185 46.390 123.555 47.130 ;
        RECT 126.485 46.950 126.915 51.920 ;
        RECT 127.425 51.910 127.655 51.975 ;
        RECT 128.565 51.910 128.795 51.975 ;
        RECT 127.365 46.910 127.765 51.910 ;
        RECT 128.445 46.910 128.845 51.910 ;
        RECT 129.355 51.880 129.585 51.975 ;
        RECT 129.295 46.910 129.725 51.880 ;
        RECT 126.915 46.540 127.375 46.770 ;
        RECT 128.845 46.650 129.305 46.770 ;
        RECT 128.695 46.540 129.305 46.650 ;
        RECT 122.405 46.280 122.635 46.370 ;
        RECT 123.195 46.280 123.425 46.390 ;
        RECT 128.695 46.370 129.275 46.540 ;
        RECT 21.505 45.950 21.965 46.180 ;
        RECT 32.705 45.960 33.165 46.190 ;
        RECT 43.925 45.930 44.385 46.160 ;
        RECT 55.175 45.910 55.635 46.140 ;
        RECT 66.395 45.900 66.855 46.130 ;
        RECT 77.635 45.890 78.095 46.120 ;
        RECT 88.885 45.900 89.345 46.130 ;
        RECT 100.165 45.890 100.625 46.120 ;
        RECT 111.435 45.890 111.895 46.120 ;
        RECT 122.685 45.890 123.145 46.120 ;
        RECT 29.055 45.020 41.225 45.030 ;
        RECT 17.855 45.005 41.225 45.020 ;
        RECT 15.900 45.000 41.225 45.005 ;
        RECT 15.900 44.980 52.445 45.000 ;
        RECT 15.900 44.970 63.695 44.980 ;
        RECT 15.900 44.960 74.915 44.970 ;
        RECT 85.235 44.960 97.405 44.970 ;
        RECT 15.900 43.880 131.205 44.960 ;
        RECT 15.900 43.870 30.025 43.880 ;
        RECT 15.900 43.855 18.690 43.870 ;
        RECT 15.900 41.620 17.050 43.855 ;
        RECT 40.275 43.850 131.205 43.880 ;
        RECT 51.525 43.830 131.205 43.850 ;
        RECT 62.745 43.820 131.205 43.830 ;
        RECT 73.985 43.810 86.155 43.820 ;
        RECT 96.515 43.810 131.205 43.820 ;
        RECT 29.015 43.330 41.185 43.340 ;
        RECT 17.815 43.310 41.185 43.330 ;
        RECT 142.830 43.320 144.150 43.340 ;
        RECT 17.815 43.290 52.405 43.310 ;
        RECT 140.750 43.300 144.150 43.320 ;
        RECT 17.815 43.280 63.655 43.290 ;
        RECT 119.895 43.280 144.150 43.300 ;
        RECT 17.815 43.270 74.875 43.280 ;
        RECT 85.195 43.270 97.365 43.280 ;
        RECT 108.685 43.270 144.150 43.280 ;
        RECT 17.815 42.180 144.150 43.270 ;
        RECT 18.755 42.150 144.150 42.180 ;
        RECT 18.755 42.120 131.165 42.150 ;
        RECT 18.755 42.090 109.655 42.120 ;
        RECT 18.755 42.080 98.445 42.090 ;
        RECT 41.325 42.070 98.445 42.080 ;
        RECT 142.830 42.070 144.150 42.150 ;
        RECT 41.325 42.060 87.205 42.070 ;
        RECT 75.035 42.050 87.205 42.060 ;
        RECT 15.900 41.540 19.685 41.620 ;
        RECT 142.070 41.610 146.210 41.640 ;
        RECT 119.855 41.590 146.210 41.610 ;
        RECT 108.645 41.550 146.210 41.590 ;
        RECT 15.900 41.520 42.165 41.540 ;
        RECT 97.445 41.530 146.210 41.550 ;
        RECT 15.900 41.510 75.875 41.520 ;
        RECT 86.235 41.510 146.210 41.530 ;
        RECT 15.900 40.500 146.210 41.510 ;
        RECT 15.900 40.480 142.320 40.500 ;
        RECT 15.900 40.470 140.920 40.480 ;
        RECT 18.715 40.460 140.920 40.470 ;
        RECT 142.070 40.460 142.250 40.480 ;
        RECT 18.715 40.440 120.815 40.460 ;
        RECT 18.715 40.400 109.615 40.440 ;
        RECT 18.715 40.390 98.405 40.400 ;
        RECT 41.285 40.380 98.405 40.390 ;
        RECT 41.285 40.370 87.165 40.380 ;
        RECT 74.995 40.360 87.165 40.370 ;
        RECT 26.775 39.230 27.235 39.460 ;
        RECT 38.055 39.230 38.515 39.460 ;
        RECT 49.345 39.210 49.805 39.440 ;
        RECT 60.565 39.210 61.025 39.440 ;
        RECT 71.765 39.210 72.225 39.440 ;
        RECT 83.055 39.200 83.515 39.430 ;
        RECT 94.295 39.220 94.755 39.450 ;
        RECT 105.505 39.240 105.965 39.470 ;
        RECT 116.705 39.280 117.165 39.510 ;
        RECT 127.915 39.300 128.375 39.530 ;
        RECT 20.645 38.810 21.225 38.980 ;
        RECT 26.495 38.960 26.725 39.070 ;
        RECT 27.285 38.980 27.515 39.070 ;
        RECT 20.615 38.700 21.225 38.810 ;
        RECT 20.615 38.580 21.075 38.700 ;
        RECT 22.545 38.580 23.005 38.810 ;
        RECT 20.195 33.470 20.625 38.440 ;
        RECT 20.335 33.375 20.565 33.470 ;
        RECT 21.075 33.440 21.475 38.440 ;
        RECT 22.155 33.440 22.555 38.440 ;
        RECT 21.125 33.375 21.355 33.440 ;
        RECT 22.265 33.375 22.495 33.440 ;
        RECT 23.005 33.430 23.435 38.400 ;
        RECT 26.365 38.220 26.735 38.960 ;
        RECT 26.495 38.070 26.725 38.220 ;
        RECT 27.265 38.210 27.655 38.980 ;
        RECT 31.925 38.810 32.505 38.980 ;
        RECT 37.775 38.960 38.005 39.070 ;
        RECT 38.565 38.980 38.795 39.070 ;
        RECT 27.285 38.070 27.515 38.210 ;
        RECT 26.635 37.660 27.355 37.920 ;
        RECT 28.675 37.690 29.445 38.760 ;
        RECT 31.895 38.700 32.505 38.810 ;
        RECT 31.895 38.580 32.355 38.700 ;
        RECT 33.825 38.580 34.285 38.810 ;
        RECT 26.495 35.480 27.215 35.740 ;
        RECT 26.345 35.200 26.575 35.295 ;
        RECT 26.215 33.520 26.585 35.200 ;
        RECT 27.135 35.120 27.365 35.295 ;
        RECT 23.055 33.375 23.285 33.430 ;
        RECT 26.345 33.295 26.575 33.520 ;
        RECT 27.125 33.400 27.495 35.120 ;
        RECT 31.475 33.470 31.905 38.440 ;
        RECT 27.135 33.295 27.365 33.400 ;
        RECT 31.615 33.375 31.845 33.470 ;
        RECT 32.355 33.440 32.755 38.440 ;
        RECT 33.435 33.440 33.835 38.440 ;
        RECT 32.405 33.375 32.635 33.440 ;
        RECT 33.545 33.375 33.775 33.440 ;
        RECT 34.285 33.430 34.715 38.400 ;
        RECT 37.645 38.220 38.015 38.960 ;
        RECT 37.775 38.070 38.005 38.220 ;
        RECT 38.545 38.210 38.935 38.980 ;
        RECT 43.215 38.790 43.795 38.960 ;
        RECT 49.065 38.940 49.295 39.050 ;
        RECT 49.855 38.960 50.085 39.050 ;
        RECT 38.565 38.070 38.795 38.210 ;
        RECT 37.915 37.660 38.635 37.920 ;
        RECT 39.955 37.690 40.725 38.760 ;
        RECT 43.185 38.680 43.795 38.790 ;
        RECT 43.185 38.560 43.645 38.680 ;
        RECT 45.115 38.560 45.575 38.790 ;
        RECT 37.775 35.480 38.495 35.740 ;
        RECT 37.625 35.200 37.855 35.295 ;
        RECT 37.495 33.520 37.865 35.200 ;
        RECT 38.415 35.120 38.645 35.295 ;
        RECT 34.335 33.375 34.565 33.430 ;
        RECT 37.625 33.295 37.855 33.520 ;
        RECT 38.405 33.400 38.775 35.120 ;
        RECT 42.765 33.450 43.195 38.420 ;
        RECT 38.415 33.295 38.645 33.400 ;
        RECT 42.905 33.355 43.135 33.450 ;
        RECT 43.645 33.420 44.045 38.420 ;
        RECT 44.725 33.420 45.125 38.420 ;
        RECT 43.695 33.355 43.925 33.420 ;
        RECT 44.835 33.355 45.065 33.420 ;
        RECT 45.575 33.410 46.005 38.380 ;
        RECT 48.935 38.200 49.305 38.940 ;
        RECT 49.065 38.050 49.295 38.200 ;
        RECT 49.835 38.190 50.225 38.960 ;
        RECT 54.435 38.790 55.015 38.960 ;
        RECT 60.285 38.940 60.515 39.050 ;
        RECT 61.075 38.960 61.305 39.050 ;
        RECT 49.855 38.050 50.085 38.190 ;
        RECT 49.205 37.640 49.925 37.900 ;
        RECT 51.245 37.670 52.015 38.740 ;
        RECT 54.405 38.680 55.015 38.790 ;
        RECT 54.405 38.560 54.865 38.680 ;
        RECT 56.335 38.560 56.795 38.790 ;
        RECT 49.065 35.460 49.785 35.720 ;
        RECT 48.915 35.180 49.145 35.275 ;
        RECT 48.785 33.500 49.155 35.180 ;
        RECT 49.705 35.100 49.935 35.275 ;
        RECT 45.625 33.355 45.855 33.410 ;
        RECT 48.915 33.275 49.145 33.500 ;
        RECT 49.695 33.380 50.065 35.100 ;
        RECT 53.985 33.450 54.415 38.420 ;
        RECT 49.705 33.275 49.935 33.380 ;
        RECT 54.125 33.355 54.355 33.450 ;
        RECT 54.865 33.420 55.265 38.420 ;
        RECT 55.945 33.420 56.345 38.420 ;
        RECT 54.915 33.355 55.145 33.420 ;
        RECT 56.055 33.355 56.285 33.420 ;
        RECT 56.795 33.410 57.225 38.380 ;
        RECT 60.155 38.200 60.525 38.940 ;
        RECT 60.285 38.050 60.515 38.200 ;
        RECT 61.055 38.190 61.445 38.960 ;
        RECT 65.635 38.790 66.215 38.960 ;
        RECT 71.485 38.940 71.715 39.050 ;
        RECT 72.275 38.960 72.505 39.050 ;
        RECT 61.075 38.050 61.305 38.190 ;
        RECT 60.425 37.640 61.145 37.900 ;
        RECT 62.465 37.670 63.235 38.740 ;
        RECT 65.605 38.680 66.215 38.790 ;
        RECT 65.605 38.560 66.065 38.680 ;
        RECT 67.535 38.560 67.995 38.790 ;
        RECT 60.285 35.460 61.005 35.720 ;
        RECT 60.135 35.180 60.365 35.275 ;
        RECT 60.005 33.500 60.375 35.180 ;
        RECT 60.925 35.100 61.155 35.275 ;
        RECT 56.845 33.355 57.075 33.410 ;
        RECT 60.135 33.275 60.365 33.500 ;
        RECT 60.915 33.380 61.285 35.100 ;
        RECT 65.185 33.450 65.615 38.420 ;
        RECT 60.925 33.275 61.155 33.380 ;
        RECT 65.325 33.355 65.555 33.450 ;
        RECT 66.065 33.420 66.465 38.420 ;
        RECT 67.145 33.420 67.545 38.420 ;
        RECT 66.115 33.355 66.345 33.420 ;
        RECT 67.255 33.355 67.485 33.420 ;
        RECT 67.995 33.410 68.425 38.380 ;
        RECT 71.355 38.200 71.725 38.940 ;
        RECT 71.485 38.050 71.715 38.200 ;
        RECT 72.255 38.190 72.645 38.960 ;
        RECT 76.925 38.780 77.505 38.950 ;
        RECT 82.775 38.930 83.005 39.040 ;
        RECT 83.565 38.950 83.795 39.040 ;
        RECT 72.275 38.050 72.505 38.190 ;
        RECT 71.625 37.640 72.345 37.900 ;
        RECT 73.665 37.670 74.435 38.740 ;
        RECT 76.895 38.670 77.505 38.780 ;
        RECT 76.895 38.550 77.355 38.670 ;
        RECT 78.825 38.550 79.285 38.780 ;
        RECT 71.485 35.460 72.205 35.720 ;
        RECT 71.335 35.180 71.565 35.275 ;
        RECT 71.205 33.500 71.575 35.180 ;
        RECT 72.125 35.100 72.355 35.275 ;
        RECT 68.045 33.355 68.275 33.410 ;
        RECT 71.335 33.275 71.565 33.500 ;
        RECT 72.115 33.380 72.485 35.100 ;
        RECT 76.475 33.440 76.905 38.410 ;
        RECT 72.125 33.275 72.355 33.380 ;
        RECT 76.615 33.345 76.845 33.440 ;
        RECT 77.355 33.410 77.755 38.410 ;
        RECT 78.435 33.410 78.835 38.410 ;
        RECT 77.405 33.345 77.635 33.410 ;
        RECT 78.545 33.345 78.775 33.410 ;
        RECT 79.285 33.400 79.715 38.370 ;
        RECT 82.645 38.190 83.015 38.930 ;
        RECT 82.775 38.040 83.005 38.190 ;
        RECT 83.545 38.180 83.935 38.950 ;
        RECT 88.165 38.800 88.745 38.970 ;
        RECT 94.015 38.950 94.245 39.060 ;
        RECT 94.805 38.970 95.035 39.060 ;
        RECT 83.565 38.040 83.795 38.180 ;
        RECT 82.915 37.630 83.635 37.890 ;
        RECT 84.955 37.660 85.725 38.730 ;
        RECT 88.135 38.690 88.745 38.800 ;
        RECT 88.135 38.570 88.595 38.690 ;
        RECT 90.065 38.570 90.525 38.800 ;
        RECT 82.775 35.450 83.495 35.710 ;
        RECT 82.625 35.170 82.855 35.265 ;
        RECT 82.495 33.490 82.865 35.170 ;
        RECT 83.415 35.090 83.645 35.265 ;
        RECT 79.335 33.345 79.565 33.400 ;
        RECT 82.625 33.265 82.855 33.490 ;
        RECT 83.405 33.370 83.775 35.090 ;
        RECT 87.715 33.460 88.145 38.430 ;
        RECT 83.415 33.265 83.645 33.370 ;
        RECT 87.855 33.365 88.085 33.460 ;
        RECT 88.595 33.430 88.995 38.430 ;
        RECT 89.675 33.430 90.075 38.430 ;
        RECT 88.645 33.365 88.875 33.430 ;
        RECT 89.785 33.365 90.015 33.430 ;
        RECT 90.525 33.420 90.955 38.390 ;
        RECT 93.885 38.210 94.255 38.950 ;
        RECT 94.015 38.060 94.245 38.210 ;
        RECT 94.785 38.200 95.175 38.970 ;
        RECT 99.375 38.820 99.955 38.990 ;
        RECT 105.225 38.970 105.455 39.080 ;
        RECT 106.015 38.990 106.245 39.080 ;
        RECT 94.805 38.060 95.035 38.200 ;
        RECT 94.155 37.650 94.875 37.910 ;
        RECT 96.195 37.680 96.965 38.750 ;
        RECT 99.345 38.710 99.955 38.820 ;
        RECT 99.345 38.590 99.805 38.710 ;
        RECT 101.275 38.590 101.735 38.820 ;
        RECT 94.015 35.470 94.735 35.730 ;
        RECT 93.865 35.190 94.095 35.285 ;
        RECT 93.735 33.510 94.105 35.190 ;
        RECT 94.655 35.110 94.885 35.285 ;
        RECT 90.575 33.365 90.805 33.420 ;
        RECT 93.865 33.285 94.095 33.510 ;
        RECT 94.645 33.390 95.015 35.110 ;
        RECT 98.925 33.480 99.355 38.450 ;
        RECT 94.655 33.285 94.885 33.390 ;
        RECT 99.065 33.385 99.295 33.480 ;
        RECT 99.805 33.450 100.205 38.450 ;
        RECT 100.885 33.450 101.285 38.450 ;
        RECT 99.855 33.385 100.085 33.450 ;
        RECT 100.995 33.385 101.225 33.450 ;
        RECT 101.735 33.440 102.165 38.410 ;
        RECT 105.095 38.230 105.465 38.970 ;
        RECT 105.225 38.080 105.455 38.230 ;
        RECT 105.995 38.220 106.385 38.990 ;
        RECT 110.575 38.860 111.155 39.030 ;
        RECT 116.425 39.010 116.655 39.120 ;
        RECT 117.215 39.030 117.445 39.120 ;
        RECT 106.015 38.080 106.245 38.220 ;
        RECT 105.365 37.670 106.085 37.930 ;
        RECT 107.405 37.700 108.175 38.770 ;
        RECT 110.545 38.750 111.155 38.860 ;
        RECT 110.545 38.630 111.005 38.750 ;
        RECT 112.475 38.630 112.935 38.860 ;
        RECT 105.225 35.490 105.945 35.750 ;
        RECT 105.075 35.210 105.305 35.305 ;
        RECT 104.945 33.530 105.315 35.210 ;
        RECT 105.865 35.130 106.095 35.305 ;
        RECT 101.785 33.385 102.015 33.440 ;
        RECT 105.075 33.305 105.305 33.530 ;
        RECT 105.855 33.410 106.225 35.130 ;
        RECT 110.125 33.520 110.555 38.490 ;
        RECT 110.265 33.425 110.495 33.520 ;
        RECT 111.005 33.490 111.405 38.490 ;
        RECT 112.085 33.490 112.485 38.490 ;
        RECT 111.055 33.425 111.285 33.490 ;
        RECT 112.195 33.425 112.425 33.490 ;
        RECT 112.935 33.480 113.365 38.450 ;
        RECT 116.295 38.270 116.665 39.010 ;
        RECT 116.425 38.120 116.655 38.270 ;
        RECT 117.195 38.260 117.585 39.030 ;
        RECT 121.785 38.880 122.365 39.050 ;
        RECT 127.635 39.030 127.865 39.140 ;
        RECT 128.425 39.050 128.655 39.140 ;
        RECT 117.215 38.120 117.445 38.260 ;
        RECT 116.565 37.710 117.285 37.970 ;
        RECT 118.605 37.740 119.375 38.810 ;
        RECT 121.755 38.770 122.365 38.880 ;
        RECT 121.755 38.650 122.215 38.770 ;
        RECT 123.685 38.650 124.145 38.880 ;
        RECT 116.425 35.530 117.145 35.790 ;
        RECT 116.275 35.250 116.505 35.345 ;
        RECT 116.145 33.570 116.515 35.250 ;
        RECT 117.065 35.170 117.295 35.345 ;
        RECT 112.985 33.425 113.215 33.480 ;
        RECT 105.865 33.305 106.095 33.410 ;
        RECT 116.275 33.345 116.505 33.570 ;
        RECT 117.055 33.450 117.425 35.170 ;
        RECT 121.335 33.540 121.765 38.510 ;
        RECT 117.065 33.345 117.295 33.450 ;
        RECT 121.475 33.445 121.705 33.540 ;
        RECT 122.215 33.510 122.615 38.510 ;
        RECT 123.295 33.510 123.695 38.510 ;
        RECT 122.265 33.445 122.495 33.510 ;
        RECT 123.405 33.445 123.635 33.510 ;
        RECT 124.145 33.500 124.575 38.470 ;
        RECT 127.505 38.290 127.875 39.030 ;
        RECT 127.635 38.140 127.865 38.290 ;
        RECT 128.405 38.280 128.795 39.050 ;
        RECT 128.425 38.140 128.655 38.280 ;
        RECT 127.775 37.730 128.495 37.990 ;
        RECT 129.815 37.760 130.585 38.830 ;
        RECT 142.850 37.630 144.170 38.900 ;
        RECT 127.635 35.550 128.355 35.810 ;
        RECT 127.485 35.270 127.715 35.365 ;
        RECT 127.355 33.590 127.725 35.270 ;
        RECT 128.275 35.190 128.505 35.365 ;
        RECT 124.195 33.445 124.425 33.500 ;
        RECT 127.485 33.365 127.715 33.590 ;
        RECT 128.265 33.470 128.635 35.190 ;
        RECT 128.275 33.365 128.505 33.470 ;
        RECT 20.615 32.940 21.075 33.170 ;
        RECT 22.545 33.130 23.005 33.170 ;
        RECT 22.485 32.850 23.115 33.130 ;
        RECT 26.625 32.860 27.085 33.090 ;
        RECT 31.895 32.940 32.355 33.170 ;
        RECT 33.825 33.130 34.285 33.170 ;
        RECT 33.765 32.850 34.395 33.130 ;
        RECT 37.905 32.860 38.365 33.090 ;
        RECT 43.185 32.920 43.645 33.150 ;
        RECT 45.115 33.110 45.575 33.150 ;
        RECT 45.055 32.830 45.685 33.110 ;
        RECT 49.195 32.840 49.655 33.070 ;
        RECT 54.405 32.920 54.865 33.150 ;
        RECT 56.335 33.110 56.795 33.150 ;
        RECT 56.275 32.830 56.905 33.110 ;
        RECT 60.415 32.840 60.875 33.070 ;
        RECT 65.605 32.920 66.065 33.150 ;
        RECT 67.535 33.110 67.995 33.150 ;
        RECT 67.475 32.830 68.105 33.110 ;
        RECT 71.615 32.840 72.075 33.070 ;
        RECT 76.895 32.910 77.355 33.140 ;
        RECT 78.825 33.100 79.285 33.140 ;
        RECT 78.765 32.820 79.395 33.100 ;
        RECT 82.905 32.830 83.365 33.060 ;
        RECT 88.135 32.930 88.595 33.160 ;
        RECT 90.065 33.120 90.525 33.160 ;
        RECT 90.005 32.840 90.635 33.120 ;
        RECT 94.145 32.850 94.605 33.080 ;
        RECT 99.345 32.950 99.805 33.180 ;
        RECT 101.275 33.140 101.735 33.180 ;
        RECT 101.215 32.860 101.845 33.140 ;
        RECT 105.355 32.870 105.815 33.100 ;
        RECT 110.545 32.990 111.005 33.220 ;
        RECT 112.475 33.180 112.935 33.220 ;
        RECT 112.415 32.900 113.045 33.180 ;
        RECT 116.555 32.910 117.015 33.140 ;
        RECT 121.755 33.010 122.215 33.240 ;
        RECT 123.685 33.200 124.145 33.240 ;
        RECT 123.625 32.920 124.255 33.200 ;
        RECT 127.765 32.930 128.225 33.160 ;
        RECT 23.185 30.880 27.925 31.180 ;
        RECT 34.465 30.880 39.205 31.180 ;
        RECT 45.755 30.860 50.495 31.160 ;
        RECT 56.975 30.860 61.715 31.160 ;
        RECT 68.175 30.860 72.915 31.160 ;
        RECT 79.465 30.850 84.205 31.150 ;
        RECT 90.705 30.870 95.445 31.170 ;
        RECT 101.915 30.890 106.655 31.190 ;
        RECT 113.115 30.930 117.855 31.230 ;
        RECT 124.325 30.950 129.065 31.250 ;
        RECT 19.485 20.270 19.905 30.160 ;
        RECT 19.585 20.090 19.815 20.270 ;
        RECT 20.805 20.260 21.175 30.210 ;
        RECT 20.875 20.090 21.105 20.260 ;
        RECT 21.935 20.220 22.305 30.170 ;
        RECT 27.255 20.270 27.615 30.190 ;
        RECT 30.765 20.270 31.185 30.160 ;
        RECT 22.015 20.090 22.245 20.220 ;
        RECT 27.305 20.090 27.535 20.270 ;
        RECT 30.865 20.090 31.095 20.270 ;
        RECT 32.085 20.260 32.455 30.210 ;
        RECT 32.155 20.090 32.385 20.260 ;
        RECT 33.215 20.220 33.585 30.170 ;
        RECT 38.535 20.270 38.895 30.190 ;
        RECT 33.295 20.090 33.525 20.220 ;
        RECT 38.585 20.090 38.815 20.270 ;
        RECT 42.055 20.250 42.475 30.140 ;
        RECT 42.155 20.070 42.385 20.250 ;
        RECT 43.375 20.240 43.745 30.190 ;
        RECT 43.445 20.070 43.675 20.240 ;
        RECT 44.505 20.200 44.875 30.150 ;
        RECT 49.825 20.250 50.185 30.170 ;
        RECT 53.275 20.250 53.695 30.140 ;
        RECT 44.585 20.070 44.815 20.200 ;
        RECT 49.875 20.070 50.105 20.250 ;
        RECT 53.375 20.070 53.605 20.250 ;
        RECT 54.595 20.240 54.965 30.190 ;
        RECT 54.665 20.070 54.895 20.240 ;
        RECT 55.725 20.200 56.095 30.150 ;
        RECT 61.045 20.250 61.405 30.170 ;
        RECT 64.475 20.250 64.895 30.140 ;
        RECT 55.805 20.070 56.035 20.200 ;
        RECT 61.095 20.070 61.325 20.250 ;
        RECT 64.575 20.070 64.805 20.250 ;
        RECT 65.795 20.240 66.165 30.190 ;
        RECT 65.865 20.070 66.095 20.240 ;
        RECT 66.925 20.200 67.295 30.150 ;
        RECT 72.245 20.250 72.605 30.170 ;
        RECT 67.005 20.070 67.235 20.200 ;
        RECT 72.295 20.070 72.525 20.250 ;
        RECT 75.765 20.240 76.185 30.130 ;
        RECT 75.865 20.060 76.095 20.240 ;
        RECT 77.085 20.230 77.455 30.180 ;
        RECT 77.155 20.060 77.385 20.230 ;
        RECT 78.215 20.190 78.585 30.140 ;
        RECT 83.535 20.240 83.895 30.160 ;
        RECT 87.005 20.260 87.425 30.150 ;
        RECT 78.295 20.060 78.525 20.190 ;
        RECT 83.585 20.060 83.815 20.240 ;
        RECT 87.105 20.080 87.335 20.260 ;
        RECT 88.325 20.250 88.695 30.200 ;
        RECT 88.395 20.080 88.625 20.250 ;
        RECT 89.455 20.210 89.825 30.160 ;
        RECT 94.775 20.260 95.135 30.180 ;
        RECT 98.215 20.280 98.635 30.170 ;
        RECT 89.535 20.080 89.765 20.210 ;
        RECT 94.825 20.080 95.055 20.260 ;
        RECT 98.315 20.100 98.545 20.280 ;
        RECT 99.535 20.270 99.905 30.220 ;
        RECT 99.605 20.100 99.835 20.270 ;
        RECT 100.665 20.230 101.035 30.180 ;
        RECT 105.985 20.280 106.345 30.200 ;
        RECT 109.415 20.320 109.835 30.210 ;
        RECT 100.745 20.100 100.975 20.230 ;
        RECT 106.035 20.100 106.265 20.280 ;
        RECT 109.515 20.140 109.745 20.320 ;
        RECT 110.735 20.310 111.105 30.260 ;
        RECT 110.805 20.140 111.035 20.310 ;
        RECT 111.865 20.270 112.235 30.220 ;
        RECT 117.185 20.320 117.545 30.240 ;
        RECT 120.625 20.340 121.045 30.230 ;
        RECT 111.945 20.140 112.175 20.270 ;
        RECT 117.235 20.140 117.465 20.320 ;
        RECT 120.725 20.160 120.955 20.340 ;
        RECT 121.945 20.330 122.315 30.280 ;
        RECT 122.015 20.160 122.245 20.330 ;
        RECT 123.075 20.290 123.445 30.240 ;
        RECT 128.395 20.340 128.755 30.260 ;
        RECT 123.155 20.160 123.385 20.290 ;
        RECT 128.445 20.160 128.675 20.340 ;
        RECT 132.345 20.170 132.755 30.180 ;
        RECT 137.735 30.120 137.965 30.130 ;
        RECT 132.445 20.130 132.675 20.170 ;
        RECT 137.665 20.080 138.055 30.120 ;
        RECT 19.775 19.610 20.925 19.920 ;
        RECT 22.185 19.620 27.335 19.900 ;
        RECT 31.055 19.610 32.205 19.920 ;
        RECT 33.465 19.620 38.615 19.900 ;
        RECT 42.345 19.590 43.495 19.900 ;
        RECT 44.755 19.600 49.905 19.880 ;
        RECT 53.565 19.590 54.715 19.900 ;
        RECT 55.975 19.600 61.125 19.880 ;
        RECT 64.765 19.590 65.915 19.900 ;
        RECT 67.175 19.600 72.325 19.880 ;
        RECT 76.055 19.580 77.205 19.890 ;
        RECT 78.465 19.590 83.615 19.870 ;
        RECT 87.295 19.600 88.445 19.910 ;
        RECT 89.705 19.610 94.855 19.890 ;
        RECT 98.505 19.620 99.655 19.930 ;
        RECT 100.915 19.630 106.065 19.910 ;
        RECT 109.705 19.660 110.855 19.970 ;
        RECT 112.115 19.670 117.265 19.950 ;
        RECT 120.915 19.680 122.065 19.990 ;
        RECT 123.325 19.690 128.475 19.970 ;
        RECT 132.635 19.640 138.025 19.930 ;
        RECT 142.940 19.110 144.080 37.630 ;
        RECT 13.940 18.460 17.635 18.530 ;
        RECT 117.755 18.510 131.425 18.530 ;
        RECT 106.545 18.470 131.425 18.510 ;
        RECT 13.940 18.440 41.565 18.460 ;
        RECT 95.345 18.450 131.425 18.470 ;
        RECT 13.940 18.430 75.275 18.440 ;
        RECT 84.135 18.430 131.425 18.450 ;
        RECT 13.940 17.380 131.425 18.430 ;
        RECT 142.890 17.990 144.140 19.110 ;
        RECT 145.070 18.880 146.210 40.500 ;
        RECT 145.030 17.960 146.250 18.880 ;
        RECT 13.950 17.370 15.100 17.380 ;
        RECT 16.615 17.360 120.215 17.380 ;
        RECT 16.615 17.320 109.015 17.360 ;
        RECT 16.615 17.310 97.805 17.320 ;
        RECT 39.185 17.300 97.805 17.310 ;
        RECT 39.185 17.290 86.565 17.300 ;
        RECT 72.895 17.280 86.565 17.290 ;
        RECT 117.765 16.950 140.620 16.960 ;
        RECT 142.040 16.950 148.010 16.980 ;
        RECT 117.765 16.940 148.010 16.950 ;
        RECT 106.555 16.900 148.010 16.940 ;
        RECT 16.625 16.870 41.575 16.890 ;
        RECT 95.355 16.880 148.010 16.900 ;
        RECT 16.625 16.860 75.285 16.870 ;
        RECT 84.145 16.860 148.010 16.880 ;
        RECT 16.625 15.840 148.010 16.860 ;
        RECT 16.625 15.820 142.660 15.840 ;
        RECT 16.625 15.810 140.620 15.820 ;
        RECT 142.040 15.810 142.660 15.820 ;
        RECT 16.625 15.790 120.225 15.810 ;
        RECT 16.625 15.750 109.025 15.790 ;
        RECT 16.625 15.740 97.815 15.750 ;
        RECT 39.195 15.730 97.815 15.740 ;
        RECT 39.195 15.720 86.575 15.730 ;
        RECT 72.905 15.710 86.575 15.720 ;
        RECT 131.215 15.460 132.585 15.470 ;
        RECT 12.290 15.390 17.625 15.450 ;
        RECT 117.795 15.440 132.785 15.460 ;
        RECT 106.585 15.400 132.785 15.440 ;
        RECT 12.290 15.370 41.585 15.390 ;
        RECT 95.385 15.380 132.785 15.400 ;
        RECT 12.290 15.360 75.295 15.370 ;
        RECT 84.175 15.360 132.785 15.380 ;
        RECT 12.290 14.320 132.785 15.360 ;
        RECT 142.905 15.040 144.045 15.050 ;
        RECT 12.290 14.310 131.445 14.320 ;
        RECT 12.290 14.300 120.235 14.310 ;
        RECT 12.320 14.280 13.470 14.300 ;
        RECT 16.655 14.290 120.235 14.300 ;
        RECT 16.655 14.250 109.035 14.290 ;
        RECT 16.655 14.240 97.825 14.250 ;
        RECT 39.225 14.230 97.825 14.240 ;
        RECT 39.225 14.220 86.585 14.230 ;
        RECT 72.935 14.210 86.585 14.220 ;
        RECT 142.850 13.920 144.100 15.040 ;
        RECT 145.020 14.870 146.160 14.980 ;
        RECT 144.980 13.950 146.200 14.870 ;
        RECT 16.965 13.800 17.435 13.810 ;
        RECT 10.800 13.780 17.435 13.800 ;
        RECT 10.800 13.720 17.555 13.780 ;
        RECT 117.845 13.770 131.445 13.790 ;
        RECT 106.635 13.730 131.445 13.770 ;
        RECT 10.800 13.700 41.585 13.720 ;
        RECT 95.435 13.710 131.445 13.730 ;
        RECT 10.800 13.690 75.295 13.700 ;
        RECT 84.225 13.690 131.445 13.710 ;
        RECT 10.800 12.650 131.445 13.690 ;
        RECT 16.705 12.640 131.445 12.650 ;
        RECT 16.705 12.620 120.235 12.640 ;
        RECT 16.705 12.580 109.035 12.620 ;
        RECT 16.705 12.570 97.825 12.580 ;
        RECT 39.275 12.560 97.825 12.570 ;
        RECT 39.275 12.550 86.585 12.560 ;
        RECT 72.985 12.540 86.585 12.550 ;
        RECT 128.755 12.240 130.465 12.250 ;
        RECT 117.545 12.220 119.255 12.230 ;
        RECT 106.345 12.180 108.055 12.190 ;
        RECT 27.615 12.170 29.325 12.180 ;
        RECT 38.895 12.170 40.605 12.180 ;
        RECT 25.675 11.030 29.325 12.170 ;
        RECT 36.955 11.030 40.605 12.170 ;
        RECT 95.135 12.160 96.845 12.170 ;
        RECT 50.185 12.150 51.895 12.160 ;
        RECT 61.405 12.150 63.115 12.160 ;
        RECT 72.605 12.150 74.315 12.160 ;
        RECT 25.675 11.020 27.625 11.030 ;
        RECT 36.955 11.020 38.905 11.030 ;
        RECT 48.245 11.010 51.895 12.150 ;
        RECT 59.465 11.010 63.115 12.150 ;
        RECT 70.665 11.010 74.315 12.150 ;
        RECT 83.895 12.140 85.605 12.150 ;
        RECT 48.245 11.000 50.195 11.010 ;
        RECT 59.465 11.000 61.415 11.010 ;
        RECT 70.665 11.000 72.615 11.010 ;
        RECT 81.955 11.000 85.605 12.140 ;
        RECT 93.195 11.020 96.845 12.160 ;
        RECT 104.405 11.040 108.055 12.180 ;
        RECT 115.605 11.080 119.255 12.220 ;
        RECT 126.815 11.100 130.465 12.240 ;
        RECT 126.815 11.090 128.765 11.100 ;
        RECT 115.605 11.070 117.555 11.080 ;
        RECT 104.405 11.030 106.355 11.040 ;
        RECT 93.195 11.010 95.145 11.020 ;
        RECT 81.955 10.990 83.905 11.000 ;
        RECT 142.905 8.580 144.045 13.920 ;
        RECT 74.420 7.440 144.045 8.580 ;
        RECT 74.420 1.410 75.560 7.440 ;
        RECT 145.020 6.630 146.160 13.950 ;
        RECT 93.650 5.490 146.160 6.630 ;
        RECT 93.650 1.480 94.790 5.490 ;
        RECT 146.870 4.560 148.010 15.840 ;
        RECT 113.130 3.420 148.010 4.560 ;
        RECT 113.130 1.610 114.270 3.420 ;
        RECT 149.460 2.770 150.600 64.660 ;
        RECT 131.940 1.880 150.600 2.770 ;
        RECT 131.800 1.630 150.600 1.880 ;
        RECT 74.290 0.160 75.680 1.410 ;
        RECT 93.500 0.230 94.890 1.480 ;
        RECT 112.900 0.360 114.290 1.610 ;
        RECT 131.800 1.380 133.490 1.630 ;
        RECT 151.730 1.420 152.870 66.900 ;
        RECT 131.800 0.430 133.540 1.380 ;
        RECT 113.130 0.330 114.270 0.360 ;
        RECT 151.600 0.300 152.970 1.420 ;
        RECT 93.650 0.150 94.790 0.230 ;
      LAYER met2 ;
        RECT 135.390 223.830 136.740 225.230 ;
        RECT 138.180 223.760 139.530 225.160 ;
        RECT 143.230 223.790 144.580 225.190 ;
        RECT 32.510 203.845 34.390 204.215 ;
        RECT 62.510 203.845 64.390 204.215 ;
        RECT 92.510 203.845 94.390 204.215 ;
        RECT 61.110 202.680 61.370 203.000 ;
        RECT 70.770 202.680 71.030 203.000 ;
        RECT 60.650 201.660 60.910 201.980 ;
        RECT 17.510 201.125 19.390 201.495 ;
        RECT 47.510 201.125 49.390 201.495 ;
        RECT 57.890 200.640 58.150 200.960 ;
        RECT 57.950 200.360 58.090 200.640 ;
        RECT 57.490 200.220 58.090 200.360 ;
        RECT 52.370 199.280 52.630 199.600 ;
        RECT 32.510 198.405 34.390 198.775 ;
        RECT 17.510 195.685 19.390 196.055 ;
        RECT 47.510 195.685 49.390 196.055 ;
        RECT 52.430 195.520 52.570 199.280 ;
        RECT 55.130 198.940 55.390 199.260 ;
        RECT 53.750 197.580 54.010 197.900 ;
        RECT 53.810 195.520 53.950 197.580 ;
        RECT 55.190 195.520 55.330 198.940 ;
        RECT 52.370 195.200 52.630 195.520 ;
        RECT 53.750 195.200 54.010 195.520 ;
        RECT 55.130 195.200 55.390 195.520 ;
        RECT 57.490 194.920 57.630 200.220 ;
        RECT 60.710 197.900 60.850 201.660 ;
        RECT 61.170 200.620 61.310 202.680 ;
        RECT 66.170 200.640 66.430 200.960 ;
        RECT 61.110 200.300 61.370 200.620 ;
        RECT 66.230 200.360 66.370 200.640 ;
        RECT 61.570 199.960 61.830 200.280 ;
        RECT 65.310 200.220 66.370 200.360 ;
        RECT 60.650 197.580 60.910 197.900 ;
        RECT 61.630 195.520 61.770 199.960 ;
        RECT 65.310 199.940 65.450 200.220 ;
        RECT 68.470 199.960 68.730 200.280 ;
        RECT 62.030 199.620 62.290 199.940 ;
        RECT 65.250 199.620 65.510 199.940 ;
        RECT 62.090 197.560 62.230 199.620 ;
        RECT 64.790 198.940 65.050 199.260 ;
        RECT 62.510 198.405 64.390 198.775 ;
        RECT 62.950 197.920 63.210 198.240 ;
        RECT 63.870 197.920 64.130 198.240 ;
        RECT 62.030 197.240 62.290 197.560 ;
        RECT 57.890 195.200 58.150 195.520 ;
        RECT 61.570 195.200 61.830 195.520 ;
        RECT 57.030 194.780 57.630 194.920 ;
        RECT 57.030 194.160 57.170 194.780 ;
        RECT 57.950 194.500 58.090 195.200 ;
        RECT 57.890 194.180 58.150 194.500 ;
        RECT 60.190 194.180 60.450 194.500 ;
        RECT 56.970 193.840 57.230 194.160 ;
        RECT 32.510 192.965 34.390 193.335 ;
        RECT 44.550 191.800 44.810 192.120 ;
        RECT 41.790 191.460 42.050 191.780 ;
        RECT 17.510 190.245 19.390 190.615 ;
        RECT 41.850 190.080 41.990 191.460 ;
        RECT 38.570 189.760 38.830 190.080 ;
        RECT 41.790 189.760 42.050 190.080 ;
        RECT 34.890 188.740 35.150 189.060 ;
        RECT 32.130 188.400 32.390 188.720 ;
        RECT 32.190 187.360 32.330 188.400 ;
        RECT 32.510 187.525 34.390 187.895 ;
        RECT 32.130 187.040 32.390 187.360 ;
        RECT 21.090 186.360 21.350 186.680 ;
        RECT 23.390 186.360 23.650 186.680 ;
        RECT 31.210 186.360 31.470 186.680 ;
        RECT 17.510 184.805 19.390 185.175 ;
        RECT 21.150 181.580 21.290 186.360 ;
        RECT 23.450 184.640 23.590 186.360 ;
        RECT 24.770 186.020 25.030 186.340 ;
        RECT 24.830 184.640 24.970 186.020 ;
        RECT 25.230 185.680 25.490 186.000 ;
        RECT 23.390 184.320 23.650 184.640 ;
        RECT 24.770 184.320 25.030 184.640 ;
        RECT 23.850 183.300 24.110 183.620 ;
        RECT 23.910 181.580 24.050 183.300 ;
        RECT 25.290 183.280 25.430 185.680 ;
        RECT 25.690 185.340 25.950 185.660 ;
        RECT 25.750 183.960 25.890 185.340 ;
        RECT 25.690 183.640 25.950 183.960 ;
        RECT 27.990 183.640 28.250 183.960 ;
        RECT 25.230 182.960 25.490 183.280 ;
        RECT 21.090 181.260 21.350 181.580 ;
        RECT 23.850 181.260 24.110 181.580 ;
        RECT 20.170 180.580 20.430 180.900 ;
        RECT 17.510 179.365 19.390 179.735 ;
        RECT 20.230 177.840 20.370 180.580 ;
        RECT 20.170 177.520 20.430 177.840 ;
        RECT 21.150 175.800 21.290 181.260 ;
        RECT 22.010 180.920 22.270 181.240 ;
        RECT 21.550 180.240 21.810 180.560 ;
        RECT 21.610 178.520 21.750 180.240 ;
        RECT 22.070 178.520 22.210 180.920 ;
        RECT 28.050 180.220 28.190 183.640 ;
        RECT 29.370 182.620 29.630 182.940 ;
        RECT 28.450 181.260 28.710 181.580 ;
        RECT 28.510 180.220 28.650 181.260 ;
        RECT 24.310 179.900 24.570 180.220 ;
        RECT 27.990 179.900 28.250 180.220 ;
        RECT 28.450 179.900 28.710 180.220 ;
        RECT 24.370 178.520 24.510 179.900 ;
        RECT 21.550 178.200 21.810 178.520 ;
        RECT 22.010 178.200 22.270 178.520 ;
        RECT 24.310 178.200 24.570 178.520 ;
        RECT 21.090 175.480 21.350 175.800 ;
        RECT 17.510 173.925 19.390 174.295 ;
        RECT 20.170 172.760 20.430 173.080 ;
        RECT 16.950 172.420 17.210 172.740 ;
        RECT 17.010 167.640 17.150 172.420 ;
        RECT 18.330 172.080 18.590 172.400 ;
        RECT 18.390 171.040 18.530 172.080 ;
        RECT 18.330 170.720 18.590 171.040 ;
        RECT 19.710 170.380 19.970 170.700 ;
        RECT 17.510 168.485 19.390 168.855 ;
        RECT 16.950 167.320 17.210 167.640 ;
        RECT 17.870 166.640 18.130 166.960 ;
        RECT 17.930 165.600 18.070 166.640 ;
        RECT 17.870 165.280 18.130 165.600 ;
        RECT 19.770 165.260 19.910 170.380 ;
        RECT 19.710 164.940 19.970 165.260 ;
        RECT 20.230 164.580 20.370 172.760 ;
        RECT 20.630 171.740 20.890 172.060 ;
        RECT 20.690 165.000 20.830 171.740 ;
        RECT 21.150 170.700 21.290 175.480 ;
        RECT 22.070 170.700 22.210 178.200 ;
        RECT 29.430 177.840 29.570 182.620 ;
        RECT 30.290 181.260 30.550 181.580 ;
        RECT 29.830 180.580 30.090 180.900 ;
        RECT 29.370 177.520 29.630 177.840 ;
        RECT 26.610 176.160 26.870 176.480 ;
        RECT 25.220 175.625 25.500 175.995 ;
        RECT 25.230 175.480 25.490 175.625 ;
        RECT 24.770 172.760 25.030 173.080 ;
        RECT 21.090 170.380 21.350 170.700 ;
        RECT 22.010 170.380 22.270 170.700 ;
        RECT 21.090 169.700 21.350 170.020 ;
        RECT 21.150 165.600 21.290 169.700 ;
        RECT 23.850 169.020 24.110 169.340 ;
        RECT 21.090 165.280 21.350 165.600 ;
        RECT 20.690 164.920 21.290 165.000 ;
        RECT 23.910 164.920 24.050 169.020 ;
        RECT 24.830 165.600 24.970 172.760 ;
        RECT 26.670 170.360 26.810 176.160 ;
        RECT 29.430 172.740 29.570 177.520 ;
        RECT 29.890 173.420 30.030 180.580 ;
        RECT 29.830 173.100 30.090 173.420 ;
        RECT 30.350 173.080 30.490 181.260 ;
        RECT 31.270 180.900 31.410 186.360 ;
        RECT 32.130 183.980 32.390 184.300 ;
        RECT 32.190 181.240 32.330 183.980 ;
        RECT 34.950 183.620 35.090 188.740 ;
        RECT 35.810 188.060 36.070 188.380 ;
        RECT 35.870 187.020 36.010 188.060 ;
        RECT 35.810 186.700 36.070 187.020 ;
        RECT 35.350 186.020 35.610 186.340 ;
        RECT 34.890 183.300 35.150 183.620 ;
        RECT 34.890 182.620 35.150 182.940 ;
        RECT 32.510 182.085 34.390 182.455 ;
        RECT 34.950 181.240 35.090 182.620 ;
        RECT 32.130 180.920 32.390 181.240 ;
        RECT 34.890 180.920 35.150 181.240 ;
        RECT 35.410 180.900 35.550 186.020 ;
        RECT 36.270 185.340 36.530 185.660 ;
        RECT 31.210 180.580 31.470 180.900 ;
        RECT 35.350 180.580 35.610 180.900 ;
        RECT 31.270 178.520 31.410 180.580 ;
        RECT 31.670 178.540 31.930 178.860 ;
        RECT 31.210 178.200 31.470 178.520 ;
        RECT 31.270 173.420 31.410 178.200 ;
        RECT 31.730 175.460 31.870 178.540 ;
        RECT 32.130 177.520 32.390 177.840 ;
        RECT 32.190 176.480 32.330 177.520 ;
        RECT 32.510 176.645 34.390 177.015 ;
        RECT 32.130 176.160 32.390 176.480 ;
        RECT 35.410 175.460 35.550 180.580 ;
        RECT 31.670 175.140 31.930 175.460 ;
        RECT 35.350 175.140 35.610 175.460 ;
        RECT 31.210 173.100 31.470 173.420 ;
        RECT 30.290 172.760 30.550 173.080 ;
        RECT 29.370 172.420 29.630 172.740 ;
        RECT 28.910 171.740 29.170 172.060 ;
        RECT 28.970 171.040 29.110 171.740 ;
        RECT 28.910 170.720 29.170 171.040 ;
        RECT 26.610 170.040 26.870 170.360 ;
        RECT 28.900 169.505 29.180 169.875 ;
        RECT 26.610 166.980 26.870 167.300 ;
        RECT 25.230 166.640 25.490 166.960 ;
        RECT 25.290 165.600 25.430 166.640 ;
        RECT 24.770 165.280 25.030 165.600 ;
        RECT 25.230 165.280 25.490 165.600 ;
        RECT 26.670 165.260 26.810 166.980 ;
        RECT 27.070 166.300 27.330 166.620 ;
        RECT 26.610 164.940 26.870 165.260 ;
        RECT 20.690 164.860 21.350 164.920 ;
        RECT 21.090 164.600 21.350 164.860 ;
        RECT 23.850 164.600 24.110 164.920 ;
        RECT 26.150 164.600 26.410 164.920 ;
        RECT 20.170 164.260 20.430 164.580 ;
        RECT 17.510 163.045 19.390 163.415 ;
        RECT 21.150 162.200 21.290 164.600 ;
        RECT 22.930 163.580 23.190 163.900 ;
        RECT 25.690 163.580 25.950 163.900 ;
        RECT 21.090 161.880 21.350 162.200 ;
        RECT 17.870 161.200 18.130 161.520 ;
        RECT 17.930 160.160 18.070 161.200 ;
        RECT 22.470 160.860 22.730 161.180 ;
        RECT 17.870 159.840 18.130 160.160 ;
        RECT 22.530 159.820 22.670 160.860 ;
        RECT 22.990 160.160 23.130 163.580 ;
        RECT 25.750 162.540 25.890 163.580 ;
        RECT 26.210 162.880 26.350 164.600 ;
        RECT 26.150 162.560 26.410 162.880 ;
        RECT 25.690 162.220 25.950 162.540 ;
        RECT 26.670 161.860 26.810 164.940 ;
        RECT 27.130 164.580 27.270 166.300 ;
        RECT 27.070 164.260 27.330 164.580 ;
        RECT 27.130 162.880 27.270 164.260 ;
        RECT 27.070 162.560 27.330 162.880 ;
        RECT 24.310 161.540 24.570 161.860 ;
        RECT 26.610 161.540 26.870 161.860 ;
        RECT 24.370 160.160 24.510 161.540 ;
        RECT 22.930 159.840 23.190 160.160 ;
        RECT 24.310 159.840 24.570 160.160 ;
        RECT 22.470 159.500 22.730 159.820 ;
        RECT 16.950 159.160 17.210 159.480 ;
        RECT 21.090 159.160 21.350 159.480 ;
        RECT 17.010 148.940 17.150 159.160 ;
        RECT 17.510 157.605 19.390 157.975 ;
        RECT 21.150 156.760 21.290 159.160 ;
        RECT 21.090 156.440 21.350 156.760 ;
        RECT 20.170 155.760 20.430 156.080 ;
        RECT 19.710 152.700 19.970 153.020 ;
        RECT 17.510 152.165 19.390 152.535 ;
        RECT 16.950 148.620 17.210 148.940 ;
        RECT 19.770 148.600 19.910 152.700 ;
        RECT 20.230 149.280 20.370 155.760 ;
        RECT 20.630 154.060 20.890 154.380 ;
        RECT 20.690 152.000 20.830 154.060 ;
        RECT 21.150 153.700 21.290 156.440 ;
        RECT 22.990 153.700 23.130 159.840 ;
        RECT 26.670 156.420 26.810 161.540 ;
        RECT 27.990 160.860 28.250 161.180 ;
        RECT 28.050 159.820 28.190 160.860 ;
        RECT 27.990 159.500 28.250 159.820 ;
        RECT 28.050 156.760 28.190 159.500 ;
        RECT 27.990 156.440 28.250 156.760 ;
        RECT 23.390 156.100 23.650 156.420 ;
        RECT 26.610 156.100 26.870 156.420 ;
        RECT 21.090 153.380 21.350 153.700 ;
        RECT 22.930 153.380 23.190 153.700 ;
        RECT 20.630 151.680 20.890 152.000 ;
        RECT 22.010 150.320 22.270 150.640 ;
        RECT 22.070 149.280 22.210 150.320 ;
        RECT 20.170 148.960 20.430 149.280 ;
        RECT 22.010 148.960 22.270 149.280 ;
        RECT 19.710 148.280 19.970 148.600 ;
        RECT 22.010 148.280 22.270 148.600 ;
        RECT 17.510 146.725 19.390 147.095 ;
        RECT 22.070 145.540 22.210 148.280 ;
        RECT 23.450 147.920 23.590 156.100 ;
        RECT 26.150 153.720 26.410 154.040 ;
        RECT 23.850 152.700 24.110 153.020 ;
        RECT 23.910 148.600 24.050 152.700 ;
        RECT 24.770 150.660 25.030 150.980 ;
        RECT 24.310 149.980 24.570 150.300 ;
        RECT 23.850 148.280 24.110 148.600 ;
        RECT 23.390 147.600 23.650 147.920 ;
        RECT 22.010 145.220 22.270 145.540 ;
        RECT 23.390 142.840 23.650 143.160 ;
        RECT 23.450 142.140 23.590 142.840 ;
        RECT 19.710 141.820 19.970 142.140 ;
        RECT 23.390 141.820 23.650 142.140 ;
        RECT 23.850 141.820 24.110 142.140 ;
        RECT 17.510 141.285 19.390 141.655 ;
        RECT 18.330 140.120 18.590 140.440 ;
        RECT 18.390 138.400 18.530 140.120 ;
        RECT 19.770 140.100 19.910 141.820 ;
        RECT 20.170 140.800 20.430 141.120 ;
        RECT 18.790 139.780 19.050 140.100 ;
        RECT 19.710 139.780 19.970 140.100 ;
        RECT 18.850 138.400 18.990 139.780 ;
        RECT 19.710 139.100 19.970 139.420 ;
        RECT 18.330 138.080 18.590 138.400 ;
        RECT 18.790 138.080 19.050 138.400 ;
        RECT 17.510 135.845 19.390 136.215 ;
        RECT 19.770 134.320 19.910 139.100 ;
        RECT 20.230 135.680 20.370 140.800 ;
        RECT 22.470 139.780 22.730 140.100 ;
        RECT 20.630 139.100 20.890 139.420 ;
        RECT 20.690 138.400 20.830 139.100 ;
        RECT 20.630 138.080 20.890 138.400 ;
        RECT 20.170 135.360 20.430 135.680 ;
        RECT 19.710 134.000 19.970 134.320 ;
        RECT 20.690 133.980 20.830 138.080 ;
        RECT 21.090 137.060 21.350 137.380 ;
        RECT 20.630 133.660 20.890 133.980 ;
        RECT 20.690 132.960 20.830 133.660 ;
        RECT 20.630 132.640 20.890 132.960 ;
        RECT 21.150 132.360 21.290 137.060 ;
        RECT 22.530 135.000 22.670 139.780 ;
        RECT 23.450 137.720 23.590 141.820 ;
        RECT 23.910 139.760 24.050 141.820 ;
        RECT 23.850 139.440 24.110 139.760 ;
        RECT 23.390 137.400 23.650 137.720 ;
        RECT 22.470 134.680 22.730 135.000 ;
        RECT 22.010 132.640 22.270 132.960 ;
        RECT 20.170 131.960 20.430 132.280 ;
        RECT 20.690 132.220 21.290 132.360 ;
        RECT 17.510 130.405 19.390 130.775 ;
        RECT 20.230 130.240 20.370 131.960 ;
        RECT 20.170 129.920 20.430 130.240 ;
        RECT 20.230 127.180 20.370 129.920 ;
        RECT 20.170 126.860 20.430 127.180 ;
        RECT 20.690 126.500 20.830 132.220 ;
        RECT 21.150 131.940 21.290 132.220 ;
        RECT 21.090 131.620 21.350 131.940 ;
        RECT 21.090 128.560 21.350 128.880 ;
        RECT 21.150 127.520 21.290 128.560 ;
        RECT 21.090 127.200 21.350 127.520 ;
        RECT 21.550 127.200 21.810 127.520 ;
        RECT 20.630 126.180 20.890 126.500 ;
        RECT 17.510 124.965 19.390 125.335 ;
        RECT 20.690 121.060 20.830 126.180 ;
        RECT 21.610 124.800 21.750 127.200 ;
        RECT 21.550 124.480 21.810 124.800 ;
        RECT 21.610 122.080 21.750 124.480 ;
        RECT 22.070 124.460 22.210 132.640 ;
        RECT 22.530 132.280 22.670 134.680 ;
        RECT 22.470 131.960 22.730 132.280 ;
        RECT 23.450 126.840 23.590 137.400 ;
        RECT 23.390 126.520 23.650 126.840 ;
        RECT 22.010 124.140 22.270 124.460 ;
        RECT 23.450 123.780 23.590 126.520 ;
        RECT 23.390 123.460 23.650 123.780 ;
        RECT 21.550 121.760 21.810 122.080 ;
        RECT 23.450 121.400 23.590 123.460 ;
        RECT 23.850 123.120 24.110 123.440 ;
        RECT 23.910 122.080 24.050 123.120 ;
        RECT 23.850 121.760 24.110 122.080 ;
        RECT 23.390 121.080 23.650 121.400 ;
        RECT 20.630 120.740 20.890 121.060 ;
        RECT 17.510 119.525 19.390 119.895 ;
        RECT 21.090 117.680 21.350 118.000 ;
        RECT 21.550 117.680 21.810 118.000 ;
        RECT 20.630 115.980 20.890 116.300 ;
        RECT 16.030 115.300 16.290 115.620 ;
        RECT 16.090 96.255 16.230 115.300 ;
        RECT 17.510 114.085 19.390 114.455 ;
        RECT 20.690 111.200 20.830 115.980 ;
        RECT 20.630 110.880 20.890 111.200 ;
        RECT 17.510 108.645 19.390 109.015 ;
        RECT 21.150 96.255 21.290 117.680 ;
        RECT 21.610 111.200 21.750 117.680 ;
        RECT 23.390 114.620 23.650 114.940 ;
        RECT 23.450 113.920 23.590 114.620 ;
        RECT 23.390 113.600 23.650 113.920 ;
        RECT 24.370 113.240 24.510 149.980 ;
        RECT 24.830 149.280 24.970 150.660 ;
        RECT 26.210 150.640 26.350 153.720 ;
        RECT 26.670 151.320 26.810 156.100 ;
        RECT 28.450 155.420 28.710 155.740 ;
        RECT 27.990 153.380 28.250 153.700 ;
        RECT 28.050 151.660 28.190 153.380 ;
        RECT 27.990 151.340 28.250 151.660 ;
        RECT 26.610 151.000 26.870 151.320 ;
        RECT 28.510 150.980 28.650 155.420 ;
        RECT 28.970 151.320 29.110 169.505 ;
        RECT 29.430 165.260 29.570 172.420 ;
        RECT 31.670 171.740 31.930 172.060 ;
        RECT 30.280 168.825 30.560 169.195 ;
        RECT 30.750 169.020 31.010 169.340 ;
        RECT 29.370 164.940 29.630 165.260 ;
        RECT 29.830 156.100 30.090 156.420 ;
        RECT 29.890 154.040 30.030 156.100 ;
        RECT 29.830 153.720 30.090 154.040 ;
        RECT 29.820 153.185 30.100 153.555 ;
        RECT 29.370 151.680 29.630 152.000 ;
        RECT 28.910 151.000 29.170 151.320 ;
        RECT 28.450 150.660 28.710 150.980 ;
        RECT 26.150 150.320 26.410 150.640 ;
        RECT 26.210 149.280 26.350 150.320 ;
        RECT 24.770 148.960 25.030 149.280 ;
        RECT 26.150 148.960 26.410 149.280 ;
        RECT 28.910 148.620 29.170 148.940 ;
        RECT 27.530 147.260 27.790 147.580 ;
        RECT 26.150 142.160 26.410 142.480 ;
        RECT 24.770 131.960 25.030 132.280 ;
        RECT 25.230 131.960 25.490 132.280 ;
        RECT 24.830 129.560 24.970 131.960 ;
        RECT 24.770 129.240 25.030 129.560 ;
        RECT 24.770 121.080 25.030 121.400 ;
        RECT 24.830 119.360 24.970 121.080 ;
        RECT 25.290 120.720 25.430 131.960 ;
        RECT 25.690 125.500 25.950 125.820 ;
        RECT 25.750 121.400 25.890 125.500 ;
        RECT 25.690 121.080 25.950 121.400 ;
        RECT 25.230 120.400 25.490 120.720 ;
        RECT 24.770 119.040 25.030 119.360 ;
        RECT 24.310 112.920 24.570 113.240 ;
        RECT 25.230 112.240 25.490 112.560 ;
        RECT 25.290 111.200 25.430 112.240 ;
        RECT 21.550 110.880 21.810 111.200 ;
        RECT 25.230 110.880 25.490 111.200 ;
        RECT 26.210 110.520 26.350 142.160 ;
        RECT 26.610 140.460 26.870 140.780 ;
        RECT 26.670 138.400 26.810 140.460 ;
        RECT 26.610 138.080 26.870 138.400 ;
        RECT 27.070 130.940 27.330 131.260 ;
        RECT 27.130 129.220 27.270 130.940 ;
        RECT 27.070 128.900 27.330 129.220 ;
        RECT 26.610 123.800 26.870 124.120 ;
        RECT 26.670 122.080 26.810 123.800 ;
        RECT 26.610 121.760 26.870 122.080 ;
        RECT 27.590 112.900 27.730 147.260 ;
        RECT 28.970 146.560 29.110 148.620 ;
        RECT 28.910 146.240 29.170 146.560 ;
        RECT 28.910 139.780 29.170 140.100 ;
        RECT 28.970 138.060 29.110 139.780 ;
        RECT 28.910 137.740 29.170 138.060 ;
        RECT 28.910 137.060 29.170 137.380 ;
        RECT 28.450 136.380 28.710 136.700 ;
        RECT 28.510 134.320 28.650 136.380 ;
        RECT 28.450 134.000 28.710 134.320 ;
        RECT 28.970 133.980 29.110 137.060 ;
        RECT 28.910 133.660 29.170 133.980 ;
        RECT 27.990 128.900 28.250 129.220 ;
        RECT 28.050 126.840 28.190 128.900 ;
        RECT 28.970 128.540 29.110 133.660 ;
        RECT 29.430 130.240 29.570 151.680 ;
        RECT 29.890 150.980 30.030 153.185 ;
        RECT 29.830 150.660 30.090 150.980 ;
        RECT 30.350 143.160 30.490 168.825 ;
        RECT 30.290 142.840 30.550 143.160 ;
        RECT 30.810 142.820 30.950 169.020 ;
        RECT 31.210 167.320 31.470 167.640 ;
        RECT 31.270 166.360 31.410 167.320 ;
        RECT 31.730 166.960 31.870 171.740 ;
        RECT 32.510 171.205 34.390 171.575 ;
        RECT 32.190 170.810 33.250 170.950 ;
        RECT 32.190 170.360 32.330 170.810 ;
        RECT 32.130 170.040 32.390 170.360 ;
        RECT 32.590 170.040 32.850 170.360 ;
        RECT 32.130 169.590 32.390 169.680 ;
        RECT 32.650 169.590 32.790 170.040 ;
        RECT 33.110 170.020 33.250 170.810 ;
        RECT 33.510 170.040 33.770 170.360 ;
        RECT 33.050 169.700 33.310 170.020 ;
        RECT 32.130 169.450 32.790 169.590 ;
        RECT 32.130 169.360 32.390 169.450 ;
        RECT 33.570 168.320 33.710 170.040 ;
        RECT 33.970 169.875 34.230 170.020 ;
        RECT 33.960 169.505 34.240 169.875 ;
        RECT 33.970 169.020 34.230 169.340 ;
        RECT 33.510 168.000 33.770 168.320 ;
        RECT 34.030 167.640 34.170 169.020 ;
        RECT 34.890 168.000 35.150 168.320 ;
        RECT 33.970 167.320 34.230 167.640 ;
        RECT 31.670 166.640 31.930 166.960 ;
        RECT 31.270 166.220 31.870 166.360 ;
        RECT 31.210 160.860 31.470 161.180 ;
        RECT 31.270 159.820 31.410 160.860 ;
        RECT 31.210 159.500 31.470 159.820 ;
        RECT 31.730 158.880 31.870 166.220 ;
        RECT 32.510 165.765 34.390 166.135 ;
        RECT 33.510 163.580 33.770 163.900 ;
        RECT 33.570 161.860 33.710 163.580 ;
        RECT 33.510 161.540 33.770 161.860 ;
        RECT 32.130 160.860 32.390 161.180 ;
        RECT 31.270 158.740 31.870 158.880 ;
        RECT 31.270 156.760 31.410 158.740 ;
        RECT 32.190 158.460 32.330 160.860 ;
        RECT 32.510 160.325 34.390 160.695 ;
        RECT 32.130 158.140 32.390 158.460 ;
        RECT 31.210 156.440 31.470 156.760 ;
        RECT 31.670 156.100 31.930 156.420 ;
        RECT 31.210 155.420 31.470 155.740 ;
        RECT 31.270 154.380 31.410 155.420 ;
        RECT 31.210 154.060 31.470 154.380 ;
        RECT 31.730 153.700 31.870 156.100 ;
        RECT 31.670 153.380 31.930 153.700 ;
        RECT 32.190 153.020 32.330 158.140 ;
        RECT 32.590 157.120 32.850 157.440 ;
        RECT 32.650 156.420 32.790 157.120 ;
        RECT 32.590 156.100 32.850 156.420 ;
        RECT 32.510 154.885 34.390 155.255 ;
        RECT 32.580 153.865 32.860 154.235 ;
        RECT 34.950 154.040 35.090 168.000 ;
        RECT 35.410 167.300 35.550 175.140 ;
        RECT 36.330 170.360 36.470 185.340 ;
        RECT 37.190 182.960 37.450 183.280 ;
        RECT 36.730 177.180 36.990 177.500 ;
        RECT 36.790 170.700 36.930 177.180 ;
        RECT 37.250 175.995 37.390 182.960 ;
        RECT 38.110 182.620 38.370 182.940 ;
        RECT 38.170 180.220 38.310 182.620 ;
        RECT 38.110 179.900 38.370 180.220 ;
        RECT 38.170 178.180 38.310 179.900 ;
        RECT 38.110 177.860 38.370 178.180 ;
        RECT 37.180 175.625 37.460 175.995 ;
        RECT 38.630 175.800 38.770 189.760 ;
        RECT 43.630 189.080 43.890 189.400 ;
        RECT 44.090 189.080 44.350 189.400 ;
        RECT 39.950 188.060 40.210 188.380 ;
        RECT 41.790 188.060 42.050 188.380 ;
        RECT 43.170 188.060 43.430 188.380 ;
        RECT 40.010 186.680 40.150 188.060 ;
        RECT 39.950 186.360 40.210 186.680 ;
        RECT 41.850 185.660 41.990 188.060 ;
        RECT 43.230 186.680 43.370 188.060 ;
        RECT 43.690 187.360 43.830 189.080 ;
        RECT 44.150 187.360 44.290 189.080 ;
        RECT 43.630 187.040 43.890 187.360 ;
        RECT 44.090 187.040 44.350 187.360 ;
        RECT 43.170 186.360 43.430 186.680 ;
        RECT 44.090 186.020 44.350 186.340 ;
        RECT 43.170 185.680 43.430 186.000 ;
        RECT 41.790 185.340 42.050 185.660 ;
        RECT 39.950 184.320 40.210 184.640 ;
        RECT 40.010 181.920 40.150 184.320 ;
        RECT 40.410 182.620 40.670 182.940 ;
        RECT 39.950 181.600 40.210 181.920 ;
        RECT 37.250 172.740 37.390 175.625 ;
        RECT 38.570 175.480 38.830 175.800 ;
        RECT 39.030 175.710 39.290 175.800 ;
        RECT 39.030 175.570 39.690 175.710 ;
        RECT 39.030 175.480 39.290 175.570 ;
        RECT 39.030 173.440 39.290 173.760 ;
        RECT 37.190 172.420 37.450 172.740 ;
        RECT 36.730 170.380 36.990 170.700 ;
        RECT 36.270 170.040 36.530 170.360 ;
        RECT 37.250 167.640 37.390 172.420 ;
        RECT 38.570 171.740 38.830 172.060 ;
        RECT 38.110 170.040 38.370 170.360 ;
        RECT 38.170 169.680 38.310 170.040 ;
        RECT 37.650 169.360 37.910 169.680 ;
        RECT 38.110 169.360 38.370 169.680 ;
        RECT 37.710 169.195 37.850 169.360 ;
        RECT 37.640 168.825 37.920 169.195 ;
        RECT 38.170 168.320 38.310 169.360 ;
        RECT 38.110 168.000 38.370 168.320 ;
        RECT 37.190 167.320 37.450 167.640 ;
        RECT 35.350 166.980 35.610 167.300 ;
        RECT 35.410 165.260 35.550 166.980 ;
        RECT 35.350 164.940 35.610 165.260 ;
        RECT 38.110 164.940 38.370 165.260 ;
        RECT 38.170 164.580 38.310 164.940 ;
        RECT 38.110 164.260 38.370 164.580 ;
        RECT 37.650 163.920 37.910 164.240 ;
        RECT 37.710 162.540 37.850 163.920 ;
        RECT 37.650 162.220 37.910 162.540 ;
        RECT 35.350 161.880 35.610 162.200 ;
        RECT 35.410 157.350 35.550 161.880 ;
        RECT 35.810 160.860 36.070 161.180 ;
        RECT 35.870 159.480 36.010 160.860 ;
        RECT 35.810 159.160 36.070 159.480 ;
        RECT 35.410 157.210 36.930 157.350 ;
        RECT 36.270 156.440 36.530 156.760 ;
        RECT 35.810 155.420 36.070 155.740 ;
        RECT 32.590 153.720 32.850 153.865 ;
        RECT 33.050 153.720 33.310 154.040 ;
        RECT 34.890 153.720 35.150 154.040 ;
        RECT 31.210 152.700 31.470 153.020 ;
        RECT 32.130 152.700 32.390 153.020 ;
        RECT 31.270 143.160 31.410 152.700 ;
        RECT 32.190 150.980 32.330 152.700 ;
        RECT 33.110 152.000 33.250 153.720 ;
        RECT 33.050 151.680 33.310 152.000 ;
        RECT 32.130 150.660 32.390 150.980 ;
        RECT 34.890 149.980 35.150 150.300 ;
        RECT 35.350 149.980 35.610 150.300 ;
        RECT 32.510 149.445 34.390 149.815 ;
        RECT 34.950 148.600 35.090 149.980 ;
        RECT 34.890 148.280 35.150 148.600 ;
        RECT 35.410 148.000 35.550 149.980 ;
        RECT 35.870 148.940 36.010 155.420 ;
        RECT 36.330 154.040 36.470 156.440 ;
        RECT 36.790 154.915 36.930 157.210 ;
        RECT 37.190 157.120 37.450 157.440 ;
        RECT 37.250 156.420 37.390 157.120 ;
        RECT 37.710 156.420 37.850 162.220 ;
        RECT 38.170 159.480 38.310 164.260 ;
        RECT 38.110 159.160 38.370 159.480 ;
        RECT 37.190 156.100 37.450 156.420 ;
        RECT 37.650 156.100 37.910 156.420 ;
        RECT 36.720 154.545 37.000 154.915 ;
        RECT 36.270 153.720 36.530 154.040 ;
        RECT 35.810 148.620 36.070 148.940 ;
        RECT 34.950 147.860 35.550 148.000 ;
        RECT 35.810 147.940 36.070 148.260 ;
        RECT 32.510 144.005 34.390 144.375 ;
        RECT 34.950 143.500 35.090 147.860 ;
        RECT 35.350 147.260 35.610 147.580 ;
        RECT 34.890 143.180 35.150 143.500 ;
        RECT 31.210 142.840 31.470 143.160 ;
        RECT 30.750 142.500 31.010 142.820 ;
        RECT 32.130 142.160 32.390 142.480 ;
        RECT 32.190 141.120 32.330 142.160 ;
        RECT 33.970 141.820 34.230 142.140 ;
        RECT 32.130 140.800 32.390 141.120 ;
        RECT 34.030 140.780 34.170 141.820 ;
        RECT 35.410 141.120 35.550 147.260 ;
        RECT 35.870 145.960 36.010 147.940 ;
        RECT 35.870 145.820 36.470 145.960 ;
        RECT 35.810 143.520 36.070 143.840 ;
        RECT 35.350 140.800 35.610 141.120 ;
        RECT 33.970 140.460 34.230 140.780 ;
        RECT 35.350 139.780 35.610 140.100 ;
        RECT 32.510 138.565 34.390 138.935 ;
        RECT 35.410 137.720 35.550 139.780 ;
        RECT 35.350 137.400 35.610 137.720 ;
        RECT 30.750 137.060 31.010 137.380 ;
        RECT 29.830 131.280 30.090 131.600 ;
        RECT 29.370 129.920 29.630 130.240 ;
        RECT 28.450 128.220 28.710 128.540 ;
        RECT 28.910 128.220 29.170 128.540 ;
        RECT 28.510 127.180 28.650 128.220 ;
        RECT 29.890 127.520 30.030 131.280 ;
        RECT 30.810 129.900 30.950 137.060 ;
        RECT 34.890 134.340 35.150 134.660 ;
        RECT 32.510 133.125 34.390 133.495 ;
        RECT 31.670 130.940 31.930 131.260 ;
        RECT 30.750 129.580 31.010 129.900 ;
        RECT 29.830 127.200 30.090 127.520 ;
        RECT 28.450 126.860 28.710 127.180 ;
        RECT 27.990 126.520 28.250 126.840 ;
        RECT 30.810 126.500 30.950 129.580 ;
        RECT 30.750 126.180 31.010 126.500 ;
        RECT 30.810 124.120 30.950 126.180 ;
        RECT 31.730 124.120 31.870 130.940 ;
        RECT 34.950 130.240 35.090 134.340 ;
        RECT 35.410 132.960 35.550 137.400 ;
        RECT 35.350 132.640 35.610 132.960 ;
        RECT 34.890 129.920 35.150 130.240 ;
        RECT 35.410 129.640 35.550 132.640 ;
        RECT 34.950 129.500 35.550 129.640 ;
        RECT 34.950 129.220 35.090 129.500 ;
        RECT 34.890 128.900 35.150 129.220 ;
        RECT 32.130 128.560 32.390 128.880 ;
        RECT 32.190 127.520 32.330 128.560 ;
        RECT 32.510 127.685 34.390 128.055 ;
        RECT 32.130 127.200 32.390 127.520 ;
        RECT 29.370 123.800 29.630 124.120 ;
        RECT 30.750 123.800 31.010 124.120 ;
        RECT 31.670 123.800 31.930 124.120 ;
        RECT 29.430 118.680 29.570 123.800 ;
        RECT 30.290 122.780 30.550 123.100 ;
        RECT 32.130 122.780 32.390 123.100 ;
        RECT 34.890 122.780 35.150 123.100 ;
        RECT 30.350 121.400 30.490 122.780 ;
        RECT 32.190 122.080 32.330 122.780 ;
        RECT 32.510 122.245 34.390 122.615 ;
        RECT 32.130 121.760 32.390 122.080 ;
        RECT 30.750 121.420 31.010 121.740 ;
        RECT 30.290 121.080 30.550 121.400 ;
        RECT 30.810 119.360 30.950 121.420 ;
        RECT 34.430 120.740 34.690 121.060 ;
        RECT 34.490 119.360 34.630 120.740 ;
        RECT 30.750 119.040 31.010 119.360 ;
        RECT 34.430 119.040 34.690 119.360 ;
        RECT 29.370 118.360 29.630 118.680 ;
        RECT 27.990 117.680 28.250 118.000 ;
        RECT 28.050 113.920 28.190 117.680 ;
        RECT 29.430 115.620 29.570 118.360 ;
        RECT 34.950 118.340 35.090 122.780 ;
        RECT 34.890 118.020 35.150 118.340 ;
        RECT 32.510 116.805 34.390 117.175 ;
        RECT 35.870 115.960 36.010 143.520 ;
        RECT 36.330 140.100 36.470 145.820 ;
        RECT 36.790 145.540 36.930 154.545 ;
        RECT 37.250 154.040 37.390 156.100 ;
        RECT 38.110 155.420 38.370 155.740 ;
        RECT 38.170 154.380 38.310 155.420 ;
        RECT 37.190 153.720 37.450 154.040 ;
        RECT 37.640 153.865 37.920 154.235 ;
        RECT 38.110 154.060 38.370 154.380 ;
        RECT 37.710 153.020 37.850 153.865 ;
        RECT 38.110 153.380 38.370 153.700 ;
        RECT 37.650 152.700 37.910 153.020 ;
        RECT 37.710 150.980 37.850 152.700 ;
        RECT 37.650 150.660 37.910 150.980 ;
        RECT 38.170 148.260 38.310 153.380 ;
        RECT 38.630 148.940 38.770 171.740 ;
        RECT 39.090 171.040 39.230 173.440 ;
        RECT 39.550 172.740 39.690 175.570 ;
        RECT 40.010 172.740 40.150 181.600 ;
        RECT 40.470 181.580 40.610 182.620 ;
        RECT 40.410 181.260 40.670 181.580 ;
        RECT 40.410 179.900 40.670 180.220 ;
        RECT 40.470 178.520 40.610 179.900 ;
        RECT 41.330 178.880 41.590 179.200 ;
        RECT 40.410 178.200 40.670 178.520 ;
        RECT 40.470 175.200 40.610 178.200 ;
        RECT 40.870 177.355 41.130 177.500 ;
        RECT 40.860 176.985 41.140 177.355 ;
        RECT 40.470 175.060 41.070 175.200 ;
        RECT 40.410 174.460 40.670 174.780 ;
        RECT 39.490 172.420 39.750 172.740 ;
        RECT 39.950 172.420 40.210 172.740 ;
        RECT 39.030 170.720 39.290 171.040 ;
        RECT 39.090 170.360 39.230 170.720 ;
        RECT 39.030 170.040 39.290 170.360 ;
        RECT 39.950 166.980 40.210 167.300 ;
        RECT 39.020 166.105 39.300 166.475 ;
        RECT 39.090 165.260 39.230 166.105 ;
        RECT 39.030 164.940 39.290 165.260 ;
        RECT 40.010 163.900 40.150 166.980 ;
        RECT 39.950 163.580 40.210 163.900 ;
        RECT 39.490 161.200 39.750 161.520 ;
        RECT 39.550 158.880 39.690 161.200 ;
        RECT 40.010 159.820 40.150 163.580 ;
        RECT 39.950 159.500 40.210 159.820 ;
        RECT 39.550 158.740 40.150 158.880 ;
        RECT 39.490 158.140 39.750 158.460 ;
        RECT 39.030 154.400 39.290 154.720 ;
        RECT 39.090 150.980 39.230 154.400 ;
        RECT 39.030 150.660 39.290 150.980 ;
        RECT 39.030 149.980 39.290 150.300 ;
        RECT 38.570 148.620 38.830 148.940 ;
        RECT 38.110 147.940 38.370 148.260 ;
        RECT 38.570 146.240 38.830 146.560 ;
        RECT 36.730 145.220 36.990 145.540 ;
        RECT 36.790 143.160 36.930 145.220 ;
        RECT 36.730 142.840 36.990 143.160 ;
        RECT 36.270 139.780 36.530 140.100 ;
        RECT 36.330 137.720 36.470 139.780 ;
        RECT 36.270 137.400 36.530 137.720 ;
        RECT 38.100 137.545 38.380 137.915 ;
        RECT 36.330 134.660 36.470 137.400 ;
        RECT 38.170 135.000 38.310 137.545 ;
        RECT 38.110 134.680 38.370 135.000 ;
        RECT 36.270 134.340 36.530 134.660 ;
        RECT 36.330 132.280 36.470 134.340 ;
        RECT 36.730 133.660 36.990 133.980 ;
        RECT 36.270 131.960 36.530 132.280 ;
        RECT 36.330 126.500 36.470 131.960 ;
        RECT 36.270 126.180 36.530 126.500 ;
        RECT 36.330 124.460 36.470 126.180 ;
        RECT 36.270 124.140 36.530 124.460 ;
        RECT 36.330 121.400 36.470 124.140 ;
        RECT 36.270 121.080 36.530 121.400 ;
        RECT 36.790 115.960 36.930 133.660 ;
        RECT 37.190 128.900 37.450 129.220 ;
        RECT 37.250 128.540 37.390 128.900 ;
        RECT 37.190 128.220 37.450 128.540 ;
        RECT 38.110 128.220 38.370 128.540 ;
        RECT 38.170 123.780 38.310 128.220 ;
        RECT 38.630 124.460 38.770 146.240 ;
        RECT 39.090 146.220 39.230 149.980 ;
        RECT 39.030 145.900 39.290 146.220 ;
        RECT 39.090 145.540 39.230 145.900 ;
        RECT 39.030 145.220 39.290 145.540 ;
        RECT 39.550 143.750 39.690 158.140 ;
        RECT 40.010 154.040 40.150 158.740 ;
        RECT 39.950 153.720 40.210 154.040 ;
        RECT 40.010 152.000 40.150 153.720 ;
        RECT 39.950 151.680 40.210 152.000 ;
        RECT 39.950 151.000 40.210 151.320 ;
        RECT 40.010 145.540 40.150 151.000 ;
        RECT 40.470 148.600 40.610 174.460 ;
        RECT 40.930 171.040 41.070 175.060 ;
        RECT 41.390 173.760 41.530 178.880 ;
        RECT 42.710 177.860 42.970 178.180 ;
        RECT 43.230 177.920 43.370 185.680 ;
        RECT 44.150 184.300 44.290 186.020 ;
        RECT 44.090 183.980 44.350 184.300 ;
        RECT 43.630 183.640 43.890 183.960 ;
        RECT 43.690 178.520 43.830 183.640 ;
        RECT 44.090 182.960 44.350 183.280 ;
        RECT 44.150 181.920 44.290 182.960 ;
        RECT 44.090 181.600 44.350 181.920 ;
        RECT 44.610 181.240 44.750 191.800 ;
        RECT 45.010 190.780 45.270 191.100 ;
        RECT 46.390 190.780 46.650 191.100 ;
        RECT 45.070 188.720 45.210 190.780 ;
        RECT 46.450 188.720 46.590 190.780 ;
        RECT 47.510 190.245 49.390 190.615 ;
        RECT 52.830 189.080 53.090 189.400 ;
        RECT 45.010 188.400 45.270 188.720 ;
        RECT 46.390 188.400 46.650 188.720 ;
        RECT 45.070 187.020 45.210 188.400 ;
        RECT 45.010 186.700 45.270 187.020 ;
        RECT 49.610 185.680 49.870 186.000 ;
        RECT 47.510 184.805 49.390 185.175 ;
        RECT 45.930 183.980 46.190 184.300 ;
        RECT 44.550 180.920 44.810 181.240 ;
        RECT 45.990 178.520 46.130 183.980 ;
        RECT 49.150 182.620 49.410 182.940 ;
        RECT 49.210 181.920 49.350 182.620 ;
        RECT 49.150 181.600 49.410 181.920 ;
        RECT 49.670 181.320 49.810 185.680 ;
        RECT 52.890 183.960 53.030 189.080 ;
        RECT 56.050 188.740 56.310 189.060 ;
        RECT 55.590 188.060 55.850 188.380 ;
        RECT 55.650 187.020 55.790 188.060 ;
        RECT 54.670 186.700 54.930 187.020 ;
        RECT 55.590 186.700 55.850 187.020 ;
        RECT 53.290 185.340 53.550 185.660 ;
        RECT 53.350 183.960 53.490 185.340 ;
        RECT 54.730 183.960 54.870 186.700 ;
        RECT 56.110 184.640 56.250 188.740 ;
        RECT 56.050 184.320 56.310 184.640 ;
        RECT 52.830 183.640 53.090 183.960 ;
        RECT 53.290 183.640 53.550 183.960 ;
        RECT 54.670 183.640 54.930 183.960 ;
        RECT 50.990 182.960 51.250 183.280 ;
        RECT 51.050 181.920 51.190 182.960 ;
        RECT 50.990 181.600 51.250 181.920 ;
        RECT 57.030 181.580 57.170 193.840 ;
        RECT 57.430 193.500 57.690 193.820 ;
        RECT 57.490 191.780 57.630 193.500 ;
        RECT 57.430 191.460 57.690 191.780 ;
        RECT 58.350 186.360 58.610 186.680 ;
        RECT 57.890 183.300 58.150 183.620 ;
        RECT 49.670 181.180 50.730 181.320 ;
        RECT 56.970 181.260 57.230 181.580 ;
        RECT 46.390 180.580 46.650 180.900 ;
        RECT 49.610 180.580 49.870 180.900 ;
        RECT 46.450 178.860 46.590 180.580 ;
        RECT 47.510 179.365 49.390 179.735 ;
        RECT 46.390 178.540 46.650 178.860 ;
        RECT 43.630 178.200 43.890 178.520 ;
        RECT 44.090 178.200 44.350 178.520 ;
        RECT 45.930 178.200 46.190 178.520 ;
        RECT 42.770 176.140 42.910 177.860 ;
        RECT 43.230 177.780 43.830 177.920 ;
        RECT 43.170 177.180 43.430 177.500 ;
        RECT 43.230 176.480 43.370 177.180 ;
        RECT 43.170 176.160 43.430 176.480 ;
        RECT 42.710 175.820 42.970 176.140 ;
        RECT 43.230 175.120 43.370 176.160 ;
        RECT 43.170 174.800 43.430 175.120 ;
        RECT 41.330 173.440 41.590 173.760 ;
        RECT 43.690 172.740 43.830 177.780 ;
        RECT 43.630 172.420 43.890 172.740 ;
        RECT 41.330 171.740 41.590 172.060 ;
        RECT 40.870 170.720 41.130 171.040 ;
        RECT 40.870 157.120 41.130 157.440 ;
        RECT 40.930 156.420 41.070 157.120 ;
        RECT 40.870 156.100 41.130 156.420 ;
        RECT 40.870 149.980 41.130 150.300 ;
        RECT 40.930 148.940 41.070 149.980 ;
        RECT 40.870 148.620 41.130 148.940 ;
        RECT 40.410 148.280 40.670 148.600 ;
        RECT 41.390 148.260 41.530 171.740 ;
        RECT 42.250 170.040 42.510 170.360 ;
        RECT 41.790 166.640 42.050 166.960 ;
        RECT 41.850 165.260 41.990 166.640 ;
        RECT 41.790 164.940 42.050 165.260 ;
        RECT 42.310 162.880 42.450 170.040 ;
        RECT 42.710 169.700 42.970 170.020 ;
        RECT 42.770 166.620 42.910 169.700 ;
        RECT 42.710 166.300 42.970 166.620 ;
        RECT 41.790 162.560 42.050 162.880 ;
        RECT 42.250 162.560 42.510 162.880 ;
        RECT 41.850 156.420 41.990 162.560 ;
        RECT 42.770 161.860 42.910 166.300 ;
        RECT 43.170 165.280 43.430 165.600 ;
        RECT 43.230 162.200 43.370 165.280 ;
        RECT 43.170 161.880 43.430 162.200 ;
        RECT 42.710 161.540 42.970 161.860 ;
        RECT 43.170 159.160 43.430 159.480 ;
        RECT 42.710 158.480 42.970 158.800 ;
        RECT 42.250 156.780 42.510 157.100 ;
        RECT 41.790 156.100 42.050 156.420 ;
        RECT 41.780 154.545 42.060 154.915 ;
        RECT 41.850 153.700 41.990 154.545 ;
        RECT 42.310 154.040 42.450 156.780 ;
        RECT 42.770 156.420 42.910 158.480 ;
        RECT 43.230 156.955 43.370 159.160 ;
        RECT 43.160 156.585 43.440 156.955 ;
        RECT 43.170 156.440 43.430 156.585 ;
        RECT 42.710 156.100 42.970 156.420 ;
        RECT 42.770 155.740 42.910 156.100 ;
        RECT 43.630 155.760 43.890 156.080 ;
        RECT 42.710 155.420 42.970 155.740 ;
        RECT 43.170 155.420 43.430 155.740 ;
        RECT 42.250 153.720 42.510 154.040 ;
        RECT 41.790 153.380 42.050 153.700 ;
        RECT 42.250 152.700 42.510 153.020 ;
        RECT 41.790 148.280 42.050 148.600 ;
        RECT 41.330 147.940 41.590 148.260 ;
        RECT 41.330 147.260 41.590 147.580 ;
        RECT 39.950 145.220 40.210 145.540 ;
        RECT 39.090 143.610 39.690 143.750 ;
        RECT 39.090 135.000 39.230 143.610 ;
        RECT 39.950 141.820 40.210 142.140 ;
        RECT 40.010 139.760 40.150 141.820 ;
        RECT 41.390 140.350 41.530 147.260 ;
        RECT 41.850 145.880 41.990 148.280 ;
        RECT 41.790 145.560 42.050 145.880 ;
        RECT 41.390 140.210 41.990 140.350 ;
        RECT 39.950 139.440 40.210 139.760 ;
        RECT 39.950 138.080 40.210 138.400 ;
        RECT 40.860 138.225 41.140 138.595 ;
        RECT 39.490 135.020 39.750 135.340 ;
        RECT 39.030 134.680 39.290 135.000 ;
        RECT 39.030 126.520 39.290 126.840 ;
        RECT 39.090 124.800 39.230 126.520 ;
        RECT 39.030 124.480 39.290 124.800 ;
        RECT 38.570 124.140 38.830 124.460 ;
        RECT 38.110 123.460 38.370 123.780 ;
        RECT 35.810 115.640 36.070 115.960 ;
        RECT 36.730 115.640 36.990 115.960 ;
        RECT 29.370 115.300 29.630 115.620 ;
        RECT 27.990 113.600 28.250 113.920 ;
        RECT 27.530 112.580 27.790 112.900 ;
        RECT 26.150 110.200 26.410 110.520 ;
        RECT 29.430 110.180 29.570 115.300 ;
        RECT 35.350 114.960 35.610 115.280 ;
        RECT 33.970 114.620 34.230 114.940 ;
        RECT 30.290 113.600 30.550 113.920 ;
        RECT 30.350 110.860 30.490 113.600 ;
        RECT 34.030 113.240 34.170 114.620 ;
        RECT 35.410 113.240 35.550 114.960 ;
        RECT 31.210 112.920 31.470 113.240 ;
        RECT 33.970 112.920 34.230 113.240 ;
        RECT 35.350 112.920 35.610 113.240 ;
        RECT 30.290 110.540 30.550 110.860 ;
        RECT 29.370 109.860 29.630 110.180 ;
        RECT 23.850 109.180 24.110 109.500 ;
        RECT 27.070 109.180 27.330 109.500 ;
        RECT 23.910 107.120 24.050 109.180 ;
        RECT 27.130 107.800 27.270 109.180 ;
        RECT 26.150 107.480 26.410 107.800 ;
        RECT 27.070 107.480 27.330 107.800 ;
        RECT 23.850 106.800 24.110 107.120 ;
        RECT 26.210 96.255 26.350 107.480 ;
        RECT 31.270 96.255 31.410 112.920 ;
        RECT 32.510 111.365 34.390 111.735 ;
        RECT 35.410 107.800 35.550 112.920 ;
        RECT 39.550 112.900 39.690 135.020 ;
        RECT 40.010 134.660 40.150 138.080 ;
        RECT 40.410 135.360 40.670 135.680 ;
        RECT 39.950 134.340 40.210 134.660 ;
        RECT 40.470 127.180 40.610 135.360 ;
        RECT 40.930 135.000 41.070 138.225 ;
        RECT 41.330 135.360 41.590 135.680 ;
        RECT 40.870 134.680 41.130 135.000 ;
        RECT 40.870 131.620 41.130 131.940 ;
        RECT 40.930 128.880 41.070 131.620 ;
        RECT 40.870 128.560 41.130 128.880 ;
        RECT 40.410 126.860 40.670 127.180 ;
        RECT 40.930 126.920 41.070 128.560 ;
        RECT 41.390 127.520 41.530 135.360 ;
        RECT 41.850 131.600 41.990 140.210 ;
        RECT 42.310 138.400 42.450 152.700 ;
        RECT 42.710 147.260 42.970 147.580 ;
        RECT 42.770 146.560 42.910 147.260 ;
        RECT 42.710 146.240 42.970 146.560 ;
        RECT 42.710 144.880 42.970 145.200 ;
        RECT 42.770 143.840 42.910 144.880 ;
        RECT 42.710 143.520 42.970 143.840 ;
        RECT 42.710 142.840 42.970 143.160 ;
        RECT 42.770 142.675 42.910 142.840 ;
        RECT 42.700 142.305 42.980 142.675 ;
        RECT 42.250 138.080 42.510 138.400 ;
        RECT 42.700 138.225 42.980 138.595 ;
        RECT 42.250 136.380 42.510 136.700 ;
        RECT 41.790 131.280 42.050 131.600 ;
        RECT 41.790 129.920 42.050 130.240 ;
        RECT 41.330 127.200 41.590 127.520 ;
        RECT 40.930 126.780 41.530 126.920 ;
        RECT 41.390 123.440 41.530 126.780 ;
        RECT 41.850 126.500 41.990 129.920 ;
        RECT 41.790 126.180 42.050 126.500 ;
        RECT 41.850 124.120 41.990 126.180 ;
        RECT 42.310 125.560 42.450 136.380 ;
        RECT 42.770 132.620 42.910 138.225 ;
        RECT 43.230 137.720 43.370 155.420 ;
        RECT 43.690 148.600 43.830 155.760 ;
        RECT 43.630 148.280 43.890 148.600 ;
        RECT 43.170 137.400 43.430 137.720 ;
        RECT 44.150 137.380 44.290 178.200 ;
        RECT 49.670 178.180 49.810 180.580 ;
        RECT 50.590 178.180 50.730 181.180 ;
        RECT 57.430 180.920 57.690 181.240 ;
        RECT 53.290 180.580 53.550 180.900 ;
        RECT 52.830 178.540 53.090 178.860 ;
        RECT 49.610 177.860 49.870 178.180 ;
        RECT 50.530 177.860 50.790 178.180 ;
        RECT 46.390 177.520 46.650 177.840 ;
        RECT 44.550 177.180 44.810 177.500 ;
        RECT 44.610 176.480 44.750 177.180 ;
        RECT 44.550 176.160 44.810 176.480 ;
        RECT 45.930 175.820 46.190 176.140 ;
        RECT 45.010 174.635 45.270 174.780 ;
        RECT 45.000 174.265 45.280 174.635 ;
        RECT 45.470 174.460 45.730 174.780 ;
        RECT 45.530 173.840 45.670 174.460 ;
        RECT 45.070 173.700 45.670 173.840 ;
        RECT 45.070 172.740 45.210 173.700 ;
        RECT 45.990 173.160 46.130 175.820 ;
        RECT 46.450 175.800 46.590 177.520 ;
        RECT 51.910 177.180 52.170 177.500 ;
        RECT 46.390 175.710 46.650 175.800 ;
        RECT 46.390 175.570 47.050 175.710 ;
        RECT 46.390 175.480 46.650 175.570 ;
        RECT 45.530 173.080 46.590 173.160 ;
        RECT 45.470 173.020 46.590 173.080 ;
        RECT 45.470 172.760 45.730 173.020 ;
        RECT 46.450 172.740 46.590 173.020 ;
        RECT 46.910 172.740 47.050 175.570 ;
        RECT 47.510 173.925 49.390 174.295 ;
        RECT 51.970 173.760 52.110 177.180 ;
        RECT 52.890 173.760 53.030 178.540 ;
        RECT 53.350 176.140 53.490 180.580 ;
        RECT 57.490 178.715 57.630 180.920 ;
        RECT 57.950 180.900 58.090 183.300 ;
        RECT 57.890 180.580 58.150 180.900 ;
        RECT 57.420 178.345 57.700 178.715 ;
        RECT 53.290 175.820 53.550 176.140 ;
        RECT 58.410 175.800 58.550 186.360 ;
        RECT 60.250 181.240 60.390 194.180 ;
        RECT 61.570 190.780 61.830 191.100 ;
        RECT 61.630 186.340 61.770 190.780 ;
        RECT 62.090 189.400 62.230 197.240 ;
        RECT 63.010 194.840 63.150 197.920 ;
        RECT 63.410 197.240 63.670 197.560 ;
        RECT 63.470 194.920 63.610 197.240 ;
        RECT 63.930 196.880 64.070 197.920 ;
        RECT 64.330 196.900 64.590 197.220 ;
        RECT 63.870 196.560 64.130 196.880 ;
        RECT 63.930 195.520 64.070 196.560 ;
        RECT 63.870 195.200 64.130 195.520 ;
        RECT 63.470 194.840 64.070 194.920 ;
        RECT 62.950 194.520 63.210 194.840 ;
        RECT 63.470 194.780 64.130 194.840 ;
        RECT 63.870 194.520 64.130 194.780 ;
        RECT 64.390 194.500 64.530 196.900 ;
        RECT 64.850 195.520 64.990 198.940 ;
        RECT 65.310 198.240 65.450 199.620 ;
        RECT 67.090 199.280 67.350 199.600 ;
        RECT 65.250 197.920 65.510 198.240 ;
        RECT 65.710 196.220 65.970 196.540 ;
        RECT 64.790 195.200 65.050 195.520 ;
        RECT 64.330 194.240 64.590 194.500 ;
        RECT 64.330 194.180 64.990 194.240 ;
        RECT 64.390 194.100 64.990 194.180 ;
        RECT 62.510 192.965 64.390 193.335 ;
        RECT 64.850 192.120 64.990 194.100 ;
        RECT 65.770 193.820 65.910 196.220 ;
        RECT 66.170 195.200 66.430 195.520 ;
        RECT 65.710 193.500 65.970 193.820 ;
        RECT 65.770 192.460 65.910 193.500 ;
        RECT 65.710 192.140 65.970 192.460 ;
        RECT 64.790 191.800 65.050 192.120 ;
        RECT 62.030 189.080 62.290 189.400 ;
        RECT 62.090 186.680 62.230 189.080 ;
        RECT 62.510 187.525 64.390 187.895 ;
        RECT 64.850 187.360 64.990 191.800 ;
        RECT 65.250 189.760 65.510 190.080 ;
        RECT 64.790 187.040 65.050 187.360 ;
        RECT 62.030 186.360 62.290 186.680 ;
        RECT 61.570 186.020 61.830 186.340 ;
        RECT 61.630 183.960 61.770 186.020 ;
        RECT 61.570 183.640 61.830 183.960 ;
        RECT 61.110 182.960 61.370 183.280 ;
        RECT 61.170 181.240 61.310 182.960 ;
        RECT 61.630 181.920 61.770 183.640 ;
        RECT 64.850 183.620 64.990 187.040 ;
        RECT 65.310 186.680 65.450 189.760 ;
        RECT 65.250 186.360 65.510 186.680 ;
        RECT 64.790 183.300 65.050 183.620 ;
        RECT 62.510 182.085 64.390 182.455 ;
        RECT 61.570 181.600 61.830 181.920 ;
        RECT 64.850 181.240 64.990 183.300 ;
        RECT 65.310 181.240 65.450 186.360 ;
        RECT 65.710 186.020 65.970 186.340 ;
        RECT 65.770 184.300 65.910 186.020 ;
        RECT 65.710 183.980 65.970 184.300 ;
        RECT 65.710 182.960 65.970 183.280 ;
        RECT 60.190 180.920 60.450 181.240 ;
        RECT 61.110 180.920 61.370 181.240 ;
        RECT 64.790 180.920 65.050 181.240 ;
        RECT 65.250 180.920 65.510 181.240 ;
        RECT 59.270 180.580 59.530 180.900 ;
        RECT 60.650 180.580 60.910 180.900 ;
        RECT 58.810 177.180 59.070 177.500 ;
        RECT 58.870 175.800 59.010 177.180 ;
        RECT 58.350 175.480 58.610 175.800 ;
        RECT 58.810 175.480 59.070 175.800 ;
        RECT 56.510 175.140 56.770 175.460 ;
        RECT 51.910 173.440 52.170 173.760 ;
        RECT 52.830 173.440 53.090 173.760 ;
        RECT 45.010 172.420 45.270 172.740 ;
        RECT 46.390 172.420 46.650 172.740 ;
        RECT 46.850 172.420 47.110 172.740 ;
        RECT 56.570 172.060 56.710 175.140 ;
        RECT 58.410 172.400 58.550 175.480 ;
        RECT 59.330 175.200 59.470 180.580 ;
        RECT 60.180 178.345 60.460 178.715 ;
        RECT 59.730 177.180 59.990 177.500 ;
        RECT 58.870 175.060 59.470 175.200 ;
        RECT 57.430 172.080 57.690 172.400 ;
        RECT 58.350 172.080 58.610 172.400 ;
        RECT 50.070 171.740 50.330 172.060 ;
        RECT 56.510 171.740 56.770 172.060 ;
        RECT 49.610 170.040 49.870 170.360 ;
        RECT 47.310 169.760 47.570 170.020 ;
        RECT 46.910 169.700 47.570 169.760 ;
        RECT 46.910 169.620 47.510 169.700 ;
        RECT 45.010 169.020 45.270 169.340 ;
        RECT 44.540 166.785 44.820 167.155 ;
        RECT 44.550 166.640 44.810 166.785 ;
        RECT 45.070 161.860 45.210 169.020 ;
        RECT 46.910 167.720 47.050 169.620 ;
        RECT 47.510 168.485 49.390 168.855 ;
        RECT 46.910 167.580 47.510 167.720 ;
        RECT 47.370 165.260 47.510 167.580 ;
        RECT 46.850 164.940 47.110 165.260 ;
        RECT 47.310 164.940 47.570 165.260 ;
        RECT 45.930 163.580 46.190 163.900 ;
        RECT 45.990 162.200 46.130 163.580 ;
        RECT 46.910 162.880 47.050 164.940 ;
        RECT 47.510 163.045 49.390 163.415 ;
        RECT 49.670 162.880 49.810 170.040 ;
        RECT 46.850 162.560 47.110 162.880 ;
        RECT 49.610 162.560 49.870 162.880 ;
        RECT 45.930 161.880 46.190 162.200 ;
        RECT 45.010 161.540 45.270 161.860 ;
        RECT 45.990 159.480 46.130 161.880 ;
        RECT 47.310 159.500 47.570 159.820 ;
        RECT 44.550 159.160 44.810 159.480 ;
        RECT 45.930 159.160 46.190 159.480 ;
        RECT 44.610 157.440 44.750 159.160 ;
        RECT 47.370 158.800 47.510 159.500 ;
        RECT 47.310 158.480 47.570 158.800 ;
        RECT 46.850 158.140 47.110 158.460 ;
        RECT 44.550 157.120 44.810 157.440 ;
        RECT 45.010 152.700 45.270 153.020 ;
        RECT 45.070 151.320 45.210 152.700 ;
        RECT 45.010 151.000 45.270 151.320 ;
        RECT 45.470 151.000 45.730 151.320 ;
        RECT 44.550 150.660 44.810 150.980 ;
        RECT 44.610 145.540 44.750 150.660 ;
        RECT 45.530 148.260 45.670 151.000 ;
        RECT 45.470 147.940 45.730 148.260 ;
        RECT 45.930 147.940 46.190 148.260 ;
        RECT 44.550 145.220 44.810 145.540 ;
        RECT 44.610 141.120 44.750 145.220 ;
        RECT 45.530 143.160 45.670 147.940 ;
        RECT 45.990 144.860 46.130 147.940 ;
        RECT 46.390 145.560 46.650 145.880 ;
        RECT 45.930 144.540 46.190 144.860 ;
        RECT 45.990 143.840 46.130 144.540 ;
        RECT 45.930 143.520 46.190 143.840 ;
        RECT 45.470 142.840 45.730 143.160 ;
        RECT 45.010 142.500 45.270 142.820 ;
        RECT 44.550 140.800 44.810 141.120 ;
        RECT 45.070 139.760 45.210 142.500 ;
        RECT 45.010 139.440 45.270 139.760 ;
        RECT 46.450 139.420 46.590 145.560 ;
        RECT 46.910 142.820 47.050 158.140 ;
        RECT 47.510 157.605 49.390 157.975 ;
        RECT 47.510 152.165 49.390 152.535 ;
        RECT 47.770 149.980 48.030 150.300 ;
        RECT 47.830 149.280 47.970 149.980 ;
        RECT 47.770 148.960 48.030 149.280 ;
        RECT 49.610 147.260 49.870 147.580 ;
        RECT 47.510 146.725 49.390 147.095 ;
        RECT 49.670 144.860 49.810 147.260 ;
        RECT 49.610 144.540 49.870 144.860 ;
        RECT 50.130 143.160 50.270 171.740 ;
        RECT 57.490 171.040 57.630 172.080 ;
        RECT 57.430 170.720 57.690 171.040 ;
        RECT 53.290 170.040 53.550 170.360 ;
        RECT 57.890 170.270 58.150 170.360 ;
        RECT 58.410 170.270 58.550 172.080 ;
        RECT 58.870 170.360 59.010 175.060 ;
        RECT 59.790 173.080 59.930 177.180 ;
        RECT 59.270 172.760 59.530 173.080 ;
        RECT 59.730 172.760 59.990 173.080 ;
        RECT 59.330 171.040 59.470 172.760 ;
        RECT 59.270 170.720 59.530 171.040 ;
        RECT 57.890 170.130 58.550 170.270 ;
        RECT 57.890 170.040 58.150 170.130 ;
        RECT 58.810 170.040 59.070 170.360 ;
        RECT 53.350 167.640 53.490 170.040 ;
        RECT 57.430 168.000 57.690 168.320 ;
        RECT 56.050 167.660 56.310 167.980 ;
        RECT 53.290 167.320 53.550 167.640 ;
        RECT 55.590 166.980 55.850 167.300 ;
        RECT 50.530 163.580 50.790 163.900 ;
        RECT 50.590 162.200 50.730 163.580 ;
        RECT 50.530 161.880 50.790 162.200 ;
        RECT 54.670 161.540 54.930 161.860 ;
        RECT 50.990 160.860 51.250 161.180 ;
        RECT 51.050 159.480 51.190 160.860 ;
        RECT 54.730 160.160 54.870 161.540 ;
        RECT 54.670 159.840 54.930 160.160 ;
        RECT 54.210 159.500 54.470 159.820 ;
        RECT 50.990 159.160 51.250 159.480 ;
        RECT 54.270 153.700 54.410 159.500 ;
        RECT 55.650 159.480 55.790 166.980 ;
        RECT 56.110 165.260 56.250 167.660 ;
        RECT 56.510 166.980 56.770 167.300 ;
        RECT 56.570 166.620 56.710 166.980 ;
        RECT 56.510 166.300 56.770 166.620 ;
        RECT 56.050 164.940 56.310 165.260 ;
        RECT 57.490 165.000 57.630 168.000 ;
        RECT 57.950 165.260 58.090 170.040 ;
        RECT 57.030 164.860 57.630 165.000 ;
        RECT 57.890 164.940 58.150 165.260 ;
        RECT 57.030 159.480 57.170 164.860 ;
        RECT 57.430 164.260 57.690 164.580 ;
        RECT 57.490 162.880 57.630 164.260 ;
        RECT 58.870 164.240 59.010 170.040 ;
        RECT 58.810 163.920 59.070 164.240 ;
        RECT 58.870 163.640 59.010 163.920 ;
        RECT 57.950 163.500 59.010 163.640 ;
        RECT 57.430 162.560 57.690 162.880 ;
        RECT 55.590 159.160 55.850 159.480 ;
        RECT 56.970 159.160 57.230 159.480 ;
        RECT 55.130 155.420 55.390 155.740 ;
        RECT 55.190 154.380 55.330 155.420 ;
        RECT 55.130 154.060 55.390 154.380 ;
        RECT 56.050 154.060 56.310 154.380 ;
        RECT 54.210 153.380 54.470 153.700 ;
        RECT 50.990 151.340 51.250 151.660 ;
        RECT 50.530 145.220 50.790 145.540 ;
        RECT 49.610 142.840 49.870 143.160 ;
        RECT 50.070 142.840 50.330 143.160 ;
        RECT 46.850 142.500 47.110 142.820 ;
        RECT 46.850 141.820 47.110 142.140 ;
        RECT 46.910 140.100 47.050 141.820 ;
        RECT 47.510 141.285 49.390 141.655 ;
        RECT 49.670 141.120 49.810 142.840 ;
        RECT 50.070 141.820 50.330 142.140 ;
        RECT 49.610 140.800 49.870 141.120 ;
        RECT 50.130 140.520 50.270 141.820 ;
        RECT 49.670 140.380 50.270 140.520 ;
        RECT 46.850 139.780 47.110 140.100 ;
        RECT 47.770 139.780 48.030 140.100 ;
        RECT 48.690 139.780 48.950 140.100 ;
        RECT 49.150 139.780 49.410 140.100 ;
        RECT 46.390 139.100 46.650 139.420 ;
        RECT 45.930 137.740 46.190 138.060 ;
        RECT 44.090 137.060 44.350 137.380 ;
        RECT 44.090 136.380 44.350 136.700 ;
        RECT 44.150 132.960 44.290 136.380 ;
        RECT 45.990 134.660 46.130 137.740 ;
        RECT 46.450 137.720 46.590 139.100 ;
        RECT 47.830 137.720 47.970 139.780 ;
        RECT 48.750 138.060 48.890 139.780 ;
        RECT 49.210 139.420 49.350 139.780 ;
        RECT 49.150 139.100 49.410 139.420 ;
        RECT 49.210 138.400 49.350 139.100 ;
        RECT 49.150 138.080 49.410 138.400 ;
        RECT 48.690 137.740 48.950 138.060 ;
        RECT 46.390 137.400 46.650 137.720 ;
        RECT 47.770 137.630 48.030 137.720 ;
        RECT 46.910 137.490 48.030 137.630 ;
        RECT 46.450 135.340 46.590 137.400 ;
        RECT 46.390 135.020 46.650 135.340 ;
        RECT 46.910 134.660 47.050 137.490 ;
        RECT 47.770 137.400 48.030 137.490 ;
        RECT 47.510 135.845 49.390 136.215 ;
        RECT 45.930 134.340 46.190 134.660 ;
        RECT 46.390 134.340 46.650 134.660 ;
        RECT 46.850 134.340 47.110 134.660 ;
        RECT 44.090 132.640 44.350 132.960 ;
        RECT 42.710 132.360 42.970 132.620 ;
        RECT 42.710 132.300 43.370 132.360 ;
        RECT 42.770 132.220 43.370 132.300 ;
        RECT 42.710 131.620 42.970 131.940 ;
        RECT 42.770 130.240 42.910 131.620 ;
        RECT 42.710 129.920 42.970 130.240 ;
        RECT 43.230 129.220 43.370 132.220 ;
        RECT 46.450 129.220 46.590 134.340 ;
        RECT 49.150 133.660 49.410 133.980 ;
        RECT 49.210 132.280 49.350 133.660 ;
        RECT 49.150 131.960 49.410 132.280 ;
        RECT 47.510 130.405 49.390 130.775 ;
        RECT 43.170 128.900 43.430 129.220 ;
        RECT 46.390 128.900 46.650 129.220 ;
        RECT 42.710 128.220 42.970 128.540 ;
        RECT 42.770 126.840 42.910 128.220 ;
        RECT 49.670 127.520 49.810 140.380 ;
        RECT 50.070 137.740 50.330 138.060 ;
        RECT 50.130 135.340 50.270 137.740 ;
        RECT 50.590 137.380 50.730 145.220 ;
        RECT 51.050 140.440 51.190 151.340 ;
        RECT 52.360 151.145 52.640 151.515 ;
        RECT 52.430 150.640 52.570 151.145 ;
        RECT 56.110 150.980 56.250 154.060 ;
        RECT 56.510 153.380 56.770 153.700 ;
        RECT 57.030 153.440 57.170 159.160 ;
        RECT 57.430 158.140 57.690 158.460 ;
        RECT 57.490 156.080 57.630 158.140 ;
        RECT 57.430 155.760 57.690 156.080 ;
        RECT 56.050 150.660 56.310 150.980 ;
        RECT 52.370 150.320 52.630 150.640 ;
        RECT 51.910 149.980 52.170 150.300 ;
        RECT 52.430 150.155 52.570 150.320 ;
        RECT 51.970 148.600 52.110 149.980 ;
        RECT 52.360 149.785 52.640 150.155 ;
        RECT 56.570 149.280 56.710 153.380 ;
        RECT 57.030 153.300 57.630 153.440 ;
        RECT 57.490 153.020 57.630 153.300 ;
        RECT 57.430 152.700 57.690 153.020 ;
        RECT 57.430 149.980 57.690 150.300 ;
        RECT 56.510 148.960 56.770 149.280 ;
        RECT 51.910 148.280 52.170 148.600 ;
        RECT 56.970 147.260 57.230 147.580 ;
        RECT 56.510 145.560 56.770 145.880 ;
        RECT 55.130 145.220 55.390 145.540 ;
        RECT 55.190 143.160 55.330 145.220 ;
        RECT 55.130 142.840 55.390 143.160 ;
        RECT 51.440 142.305 51.720 142.675 ;
        RECT 50.990 140.120 51.250 140.440 ;
        RECT 50.990 137.400 51.250 137.720 ;
        RECT 50.530 137.060 50.790 137.380 ;
        RECT 50.070 135.020 50.330 135.340 ;
        RECT 50.590 131.940 50.730 137.060 ;
        RECT 51.050 135.340 51.190 137.400 ;
        RECT 50.990 135.020 51.250 135.340 ;
        RECT 51.050 134.660 51.190 135.020 ;
        RECT 51.510 134.660 51.650 142.305 ;
        RECT 54.210 141.820 54.470 142.140 ;
        RECT 52.370 139.100 52.630 139.420 ;
        RECT 52.430 136.700 52.570 139.100 ;
        RECT 53.290 136.720 53.550 137.040 ;
        RECT 52.370 136.380 52.630 136.700 ;
        RECT 50.990 134.340 51.250 134.660 ;
        RECT 51.450 134.340 51.710 134.660 ;
        RECT 52.430 134.320 52.570 136.380 ;
        RECT 53.350 135.000 53.490 136.720 ;
        RECT 53.290 134.680 53.550 135.000 ;
        RECT 52.370 134.000 52.630 134.320 ;
        RECT 50.530 131.620 50.790 131.940 ;
        RECT 51.450 131.620 51.710 131.940 ;
        RECT 50.590 130.240 50.730 131.620 ;
        RECT 50.530 129.920 50.790 130.240 ;
        RECT 49.610 127.200 49.870 127.520 ;
        RECT 50.590 126.840 50.730 129.920 ;
        RECT 51.510 129.560 51.650 131.620 ;
        RECT 53.350 131.260 53.490 134.680 ;
        RECT 53.290 130.940 53.550 131.260 ;
        RECT 51.450 129.240 51.710 129.560 ;
        RECT 42.710 126.520 42.970 126.840 ;
        RECT 50.530 126.520 50.790 126.840 ;
        RECT 44.550 126.180 44.810 126.500 ;
        RECT 46.390 126.180 46.650 126.500 ;
        RECT 42.310 125.420 42.910 125.560 ;
        RECT 41.790 123.800 42.050 124.120 ;
        RECT 41.330 123.120 41.590 123.440 ;
        RECT 41.390 122.080 41.530 123.120 ;
        RECT 42.250 122.780 42.510 123.100 ;
        RECT 41.330 121.760 41.590 122.080 ;
        RECT 41.790 121.420 42.050 121.740 ;
        RECT 41.330 120.060 41.590 120.380 ;
        RECT 41.390 118.340 41.530 120.060 ;
        RECT 41.850 119.360 41.990 121.420 ;
        RECT 41.790 119.040 42.050 119.360 ;
        RECT 42.310 118.340 42.450 122.780 ;
        RECT 41.330 118.020 41.590 118.340 ;
        RECT 42.250 118.020 42.510 118.340 ;
        RECT 42.770 112.900 42.910 125.420 ;
        RECT 44.610 123.100 44.750 126.180 ;
        RECT 46.450 123.780 46.590 126.180 ;
        RECT 47.510 124.965 49.390 125.335 ;
        RECT 49.610 124.140 49.870 124.460 ;
        RECT 46.390 123.460 46.650 123.780 ;
        RECT 44.550 122.780 44.810 123.100 ;
        RECT 47.310 122.780 47.570 123.100 ;
        RECT 44.090 120.740 44.350 121.060 ;
        RECT 44.150 119.360 44.290 120.740 ;
        RECT 44.610 119.360 44.750 122.780 ;
        RECT 47.370 121.400 47.510 122.780 ;
        RECT 49.670 121.740 49.810 124.140 ;
        RECT 50.590 123.100 50.730 126.520 ;
        RECT 51.510 124.120 51.650 129.240 ;
        RECT 51.910 128.900 52.170 129.220 ;
        RECT 51.970 124.800 52.110 128.900 ;
        RECT 51.910 124.480 52.170 124.800 ;
        RECT 51.450 123.800 51.710 124.120 ;
        RECT 50.530 122.780 50.790 123.100 ;
        RECT 49.610 121.420 49.870 121.740 ;
        RECT 47.310 121.080 47.570 121.400 ;
        RECT 49.610 120.060 49.870 120.380 ;
        RECT 51.910 120.060 52.170 120.380 ;
        RECT 47.510 119.525 49.390 119.895 ;
        RECT 44.090 119.040 44.350 119.360 ;
        RECT 44.550 119.040 44.810 119.360 ;
        RECT 49.670 118.760 49.810 120.060 ;
        RECT 49.210 118.620 49.810 118.760 ;
        RECT 51.970 118.680 52.110 120.060 ;
        RECT 49.210 118.000 49.350 118.620 ;
        RECT 51.910 118.360 52.170 118.680 ;
        RECT 49.150 117.680 49.410 118.000 ;
        RECT 52.370 114.620 52.630 114.940 ;
        RECT 47.510 114.085 49.390 114.455 ;
        RECT 48.690 113.600 48.950 113.920 ;
        RECT 38.110 112.580 38.370 112.900 ;
        RECT 39.490 112.580 39.750 112.900 ;
        RECT 42.710 112.580 42.970 112.900 ;
        RECT 46.850 112.580 47.110 112.900 ;
        RECT 35.810 111.900 36.070 112.220 ;
        RECT 35.870 110.860 36.010 111.900 ;
        RECT 38.170 111.200 38.310 112.580 ;
        RECT 44.550 112.240 44.810 112.560 ;
        RECT 38.110 110.880 38.370 111.200 ;
        RECT 35.810 110.540 36.070 110.860 ;
        RECT 36.270 109.860 36.530 110.180 ;
        RECT 35.350 107.480 35.610 107.800 ;
        RECT 32.510 105.925 34.390 106.295 ;
        RECT 36.330 96.255 36.470 109.860 ;
        RECT 38.170 107.460 38.310 110.880 ;
        RECT 41.790 110.540 42.050 110.860 ;
        RECT 41.330 109.520 41.590 109.840 ;
        RECT 38.110 107.140 38.370 107.460 ;
        RECT 41.390 96.255 41.530 109.520 ;
        RECT 41.850 108.480 41.990 110.540 ;
        RECT 41.790 108.160 42.050 108.480 ;
        RECT 16.020 94.255 16.300 96.255 ;
        RECT 21.080 94.255 21.360 96.255 ;
        RECT 26.140 94.255 26.420 96.255 ;
        RECT 31.200 94.255 31.480 96.255 ;
        RECT 36.260 94.255 36.540 96.255 ;
        RECT 41.320 94.255 41.600 96.255 ;
        RECT 44.610 95.640 44.750 112.240 ;
        RECT 45.470 111.900 45.730 112.220 ;
        RECT 45.530 110.860 45.670 111.900 ;
        RECT 45.470 110.540 45.730 110.860 ;
        RECT 46.910 108.480 47.050 112.580 ;
        RECT 48.750 110.520 48.890 113.600 ;
        RECT 52.430 113.240 52.570 114.620 ;
        RECT 52.370 112.920 52.630 113.240 ;
        RECT 54.270 112.900 54.410 141.820 ;
        RECT 56.570 140.440 56.710 145.560 ;
        RECT 57.030 143.160 57.170 147.260 ;
        RECT 57.490 145.540 57.630 149.980 ;
        RECT 57.430 145.220 57.690 145.540 ;
        RECT 56.970 142.840 57.230 143.160 ;
        RECT 57.030 142.480 57.170 142.840 ;
        RECT 56.970 142.160 57.230 142.480 ;
        RECT 57.490 141.120 57.630 145.220 ;
        RECT 57.430 140.800 57.690 141.120 ;
        RECT 55.130 140.120 55.390 140.440 ;
        RECT 56.510 140.120 56.770 140.440 ;
        RECT 55.190 135.000 55.330 140.120 ;
        RECT 56.510 139.100 56.770 139.420 ;
        RECT 55.590 137.740 55.850 138.060 ;
        RECT 55.650 135.680 55.790 137.740 ;
        RECT 56.570 137.630 56.710 139.100 ;
        RECT 56.970 137.630 57.230 137.720 ;
        RECT 56.570 137.490 57.230 137.630 ;
        RECT 56.970 137.400 57.230 137.490 ;
        RECT 55.590 135.360 55.850 135.680 ;
        RECT 55.130 134.680 55.390 135.000 ;
        RECT 55.190 131.680 55.330 134.680 ;
        RECT 57.430 133.660 57.690 133.980 ;
        RECT 57.490 132.620 57.630 133.660 ;
        RECT 57.430 132.300 57.690 132.620 ;
        RECT 55.190 131.540 55.790 131.680 ;
        RECT 57.950 131.600 58.090 163.500 ;
        RECT 58.350 162.560 58.610 162.880 ;
        RECT 58.410 159.140 58.550 162.560 ;
        RECT 58.350 158.820 58.610 159.140 ;
        RECT 58.810 158.140 59.070 158.460 ;
        RECT 58.870 154.720 59.010 158.140 ;
        RECT 58.810 154.400 59.070 154.720 ;
        RECT 58.350 152.700 58.610 153.020 ;
        RECT 58.410 151.320 58.550 152.700 ;
        RECT 58.870 152.000 59.010 154.400 ;
        RECT 59.330 154.235 59.470 170.720 ;
        RECT 60.250 168.320 60.390 178.345 ;
        RECT 60.710 177.500 60.850 180.580 ;
        RECT 61.170 178.600 61.310 180.920 ;
        RECT 63.870 180.755 64.130 180.900 ;
        RECT 63.860 180.385 64.140 180.755 ;
        RECT 61.170 178.520 61.770 178.600 ;
        RECT 61.170 178.460 61.830 178.520 ;
        RECT 61.570 178.200 61.830 178.460 ;
        RECT 61.110 177.860 61.370 178.180 ;
        RECT 60.650 177.180 60.910 177.500 ;
        RECT 61.170 176.480 61.310 177.860 ;
        RECT 61.110 176.160 61.370 176.480 ;
        RECT 61.630 175.800 61.770 178.200 ;
        RECT 65.770 178.180 65.910 182.960 ;
        RECT 65.710 177.860 65.970 178.180 ;
        RECT 65.710 177.180 65.970 177.500 ;
        RECT 62.510 176.645 64.390 177.015 ;
        RECT 65.770 175.800 65.910 177.180 ;
        RECT 61.570 175.480 61.830 175.800 ;
        RECT 65.710 175.480 65.970 175.800 ;
        RECT 65.770 172.740 65.910 175.480 ;
        RECT 65.710 172.420 65.970 172.740 ;
        RECT 65.250 171.740 65.510 172.060 ;
        RECT 62.510 171.205 64.390 171.575 ;
        RECT 63.410 170.040 63.670 170.360 ;
        RECT 64.790 170.040 65.050 170.360 ;
        RECT 60.190 168.000 60.450 168.320 ;
        RECT 63.470 167.640 63.610 170.040 ;
        RECT 60.190 167.320 60.450 167.640 ;
        RECT 63.410 167.320 63.670 167.640 ;
        RECT 60.250 161.860 60.390 167.320 ;
        RECT 61.570 166.980 61.830 167.300 ;
        RECT 61.630 164.920 61.770 166.980 ;
        RECT 64.850 166.620 64.990 170.040 ;
        RECT 65.310 169.680 65.450 171.740 ;
        RECT 65.770 170.700 65.910 172.420 ;
        RECT 65.710 170.380 65.970 170.700 ;
        RECT 65.250 169.360 65.510 169.680 ;
        RECT 66.230 168.320 66.370 195.200 ;
        RECT 66.630 194.180 66.890 194.500 ;
        RECT 66.690 191.440 66.830 194.180 ;
        RECT 67.150 192.800 67.290 199.280 ;
        RECT 68.530 194.840 68.670 199.960 ;
        RECT 70.830 199.940 70.970 202.680 ;
        RECT 73.530 201.660 73.790 201.980 ;
        RECT 70.770 199.620 71.030 199.940 ;
        RECT 73.590 199.600 73.730 201.660 ;
        RECT 77.510 201.125 79.390 201.495 ;
        RECT 107.510 201.125 109.390 201.495 ;
        RECT 84.570 199.960 84.830 200.280 ;
        RECT 73.530 199.280 73.790 199.600 ;
        RECT 76.750 199.280 77.010 199.600 ;
        RECT 68.930 198.940 69.190 199.260 ;
        RECT 68.990 197.900 69.130 198.940 ;
        RECT 68.930 197.580 69.190 197.900 ;
        RECT 70.310 196.900 70.570 197.220 ;
        RECT 72.610 196.900 72.870 197.220 ;
        RECT 69.390 196.220 69.650 196.540 ;
        RECT 68.470 194.520 68.730 194.840 ;
        RECT 68.530 192.800 68.670 194.520 ;
        RECT 69.450 194.500 69.590 196.220 ;
        RECT 70.370 194.500 70.510 196.900 ;
        RECT 72.150 196.220 72.410 196.540 ;
        RECT 72.210 194.840 72.350 196.220 ;
        RECT 72.670 195.520 72.810 196.900 ;
        RECT 76.810 195.520 76.950 199.280 ;
        RECT 79.510 198.940 79.770 199.260 ;
        RECT 79.570 197.900 79.710 198.940 ;
        RECT 79.510 197.580 79.770 197.900 ;
        RECT 82.270 197.580 82.530 197.900 ;
        RECT 77.510 195.685 79.390 196.055 ;
        RECT 82.330 195.520 82.470 197.580 ;
        RECT 84.630 197.220 84.770 199.960 ;
        RECT 85.950 199.620 86.210 199.940 ;
        RECT 84.570 196.900 84.830 197.220 ;
        RECT 72.610 195.200 72.870 195.520 ;
        RECT 76.750 195.200 77.010 195.520 ;
        RECT 82.270 195.200 82.530 195.520 ;
        RECT 72.150 194.520 72.410 194.840 ;
        RECT 73.070 194.520 73.330 194.840 ;
        RECT 77.670 194.520 77.930 194.840 ;
        RECT 69.390 194.180 69.650 194.500 ;
        RECT 70.310 194.180 70.570 194.500 ;
        RECT 68.930 193.840 69.190 194.160 ;
        RECT 68.990 192.800 69.130 193.840 ;
        RECT 67.090 192.480 67.350 192.800 ;
        RECT 68.470 192.480 68.730 192.800 ;
        RECT 68.930 192.480 69.190 192.800 ;
        RECT 66.630 191.120 66.890 191.440 ;
        RECT 68.530 189.060 68.670 192.480 ;
        RECT 69.450 191.780 69.590 194.180 ;
        RECT 70.370 192.200 70.510 194.180 ;
        RECT 72.150 193.840 72.410 194.160 ;
        RECT 71.230 193.500 71.490 193.820 ;
        RECT 70.370 192.120 70.970 192.200 ;
        RECT 70.370 192.060 71.030 192.120 ;
        RECT 69.390 191.460 69.650 191.780 ;
        RECT 68.470 188.740 68.730 189.060 ;
        RECT 69.450 186.340 69.590 191.460 ;
        RECT 69.850 190.780 70.110 191.100 ;
        RECT 69.390 186.020 69.650 186.340 ;
        RECT 66.630 185.340 66.890 185.660 ;
        RECT 66.170 168.000 66.430 168.320 ;
        RECT 65.250 167.660 65.510 167.980 ;
        RECT 64.790 166.300 65.050 166.620 ;
        RECT 62.510 165.765 64.390 166.135 ;
        RECT 64.850 165.260 64.990 166.300 ;
        RECT 64.790 164.940 65.050 165.260 ;
        RECT 61.110 164.600 61.370 164.920 ;
        RECT 61.570 164.600 61.830 164.920 ;
        RECT 60.190 161.540 60.450 161.860 ;
        RECT 59.730 160.860 59.990 161.180 ;
        RECT 59.790 157.440 59.930 160.860 ;
        RECT 60.250 159.480 60.390 161.540 ;
        RECT 60.190 159.160 60.450 159.480 ;
        RECT 59.730 157.120 59.990 157.440 ;
        RECT 60.250 154.720 60.390 159.160 ;
        RECT 60.650 158.140 60.910 158.460 ;
        RECT 60.190 154.400 60.450 154.720 ;
        RECT 59.260 153.865 59.540 154.235 ;
        RECT 58.810 151.680 59.070 152.000 ;
        RECT 58.350 151.000 58.610 151.320 ;
        RECT 58.410 145.880 58.550 151.000 ;
        RECT 59.330 150.300 59.470 153.865 ;
        RECT 60.190 153.040 60.450 153.360 ;
        RECT 60.250 152.880 60.390 153.040 ;
        RECT 59.790 152.740 60.390 152.880 ;
        RECT 59.270 149.980 59.530 150.300 ;
        RECT 59.790 149.360 59.930 152.740 ;
        RECT 60.710 150.980 60.850 158.140 ;
        RECT 61.170 156.420 61.310 164.600 ;
        RECT 65.310 161.600 65.450 167.660 ;
        RECT 65.710 162.220 65.970 162.540 ;
        RECT 64.850 161.460 65.450 161.600 ;
        RECT 65.770 161.520 65.910 162.220 ;
        RECT 66.230 161.860 66.370 168.000 ;
        RECT 66.690 167.300 66.830 185.340 ;
        RECT 69.450 184.640 69.590 186.020 ;
        RECT 69.390 184.320 69.650 184.640 ;
        RECT 68.010 183.980 68.270 184.300 ;
        RECT 68.070 182.940 68.210 183.980 ;
        RECT 68.010 182.620 68.270 182.940 ;
        RECT 68.930 182.620 69.190 182.940 ;
        RECT 68.470 178.540 68.730 178.860 ;
        RECT 68.530 178.180 68.670 178.540 ;
        RECT 67.090 178.090 67.350 178.180 ;
        RECT 67.090 177.950 67.750 178.090 ;
        RECT 67.090 177.860 67.350 177.950 ;
        RECT 67.090 174.635 67.350 174.780 ;
        RECT 67.080 174.265 67.360 174.635 ;
        RECT 67.610 167.980 67.750 177.950 ;
        RECT 68.470 177.860 68.730 178.180 ;
        RECT 68.530 175.800 68.670 177.860 ;
        RECT 68.470 175.480 68.730 175.800 ;
        RECT 68.010 171.740 68.270 172.060 ;
        RECT 68.070 171.040 68.210 171.740 ;
        RECT 68.010 170.720 68.270 171.040 ;
        RECT 67.550 167.660 67.810 167.980 ;
        RECT 66.630 166.980 66.890 167.300 ;
        RECT 66.690 162.200 66.830 166.980 ;
        RECT 67.550 162.560 67.810 162.880 ;
        RECT 66.630 161.880 66.890 162.200 ;
        RECT 66.170 161.540 66.430 161.860 ;
        RECT 62.030 160.860 62.290 161.180 ;
        RECT 61.560 159.305 61.840 159.675 ;
        RECT 61.570 159.160 61.830 159.305 ;
        RECT 62.090 158.880 62.230 160.860 ;
        RECT 62.510 160.325 64.390 160.695 ;
        RECT 63.870 159.840 64.130 160.160 ;
        RECT 62.090 158.740 62.690 158.880 ;
        RECT 62.030 158.140 62.290 158.460 ;
        RECT 61.110 156.100 61.370 156.420 ;
        RECT 61.170 153.700 61.310 156.100 ;
        RECT 61.570 155.760 61.830 156.080 ;
        RECT 61.110 153.380 61.370 153.700 ;
        RECT 61.630 152.880 61.770 155.760 ;
        RECT 62.090 153.950 62.230 158.140 ;
        RECT 62.550 157.100 62.690 158.740 ;
        RECT 62.490 156.780 62.750 157.100 ;
        RECT 63.930 156.760 64.070 159.840 ;
        RECT 64.850 159.730 64.990 161.460 ;
        RECT 65.710 161.200 65.970 161.520 ;
        RECT 66.630 161.200 66.890 161.520 ;
        RECT 65.250 160.860 65.510 161.180 ;
        RECT 64.390 159.590 64.990 159.730 ;
        RECT 63.870 156.440 64.130 156.760 ;
        RECT 64.390 156.420 64.530 159.590 ;
        RECT 65.310 159.480 65.450 160.860 ;
        RECT 65.700 160.665 65.980 161.035 ;
        RECT 65.770 159.820 65.910 160.665 ;
        RECT 66.160 159.985 66.440 160.355 ;
        RECT 66.690 160.160 66.830 161.200 ;
        RECT 67.090 160.860 67.350 161.180 ;
        RECT 65.710 159.500 65.970 159.820 ;
        RECT 66.230 159.480 66.370 159.985 ;
        RECT 66.630 159.840 66.890 160.160 ;
        RECT 65.250 159.160 65.510 159.480 ;
        RECT 66.170 159.160 66.430 159.480 ;
        RECT 66.630 159.390 66.890 159.480 ;
        RECT 67.150 159.390 67.290 160.860 ;
        RECT 67.610 160.160 67.750 162.560 ;
        RECT 68.990 161.035 69.130 182.620 ;
        RECT 69.390 180.580 69.650 180.900 ;
        RECT 69.450 178.860 69.590 180.580 ;
        RECT 69.390 178.540 69.650 178.860 ;
        RECT 69.450 175.800 69.590 178.540 ;
        RECT 69.390 175.480 69.650 175.800 ;
        RECT 69.910 173.840 70.050 190.780 ;
        RECT 70.370 190.080 70.510 192.060 ;
        RECT 70.770 191.800 71.030 192.060 ;
        RECT 71.290 191.100 71.430 193.500 ;
        RECT 72.210 192.800 72.350 193.840 ;
        RECT 73.130 192.800 73.270 194.520 ;
        RECT 75.830 193.500 76.090 193.820 ;
        RECT 72.150 192.480 72.410 192.800 ;
        RECT 73.070 192.480 73.330 192.800 ;
        RECT 75.890 192.460 76.030 193.500 ;
        RECT 75.830 192.140 76.090 192.460 ;
        RECT 77.730 191.780 77.870 194.520 ;
        RECT 86.010 194.500 86.150 199.620 ;
        RECT 92.510 198.405 94.390 198.775 ;
        RECT 86.870 196.900 87.130 197.220 ;
        RECT 95.610 196.900 95.870 197.220 ;
        RECT 85.950 194.180 86.210 194.500 ;
        RECT 86.410 194.180 86.670 194.500 ;
        RECT 85.950 193.500 86.210 193.820 ;
        RECT 81.350 191.800 81.610 192.120 ;
        RECT 77.670 191.460 77.930 191.780 ;
        RECT 71.230 190.780 71.490 191.100 ;
        RECT 77.510 190.245 79.390 190.615 ;
        RECT 70.310 189.760 70.570 190.080 ;
        RECT 70.370 184.300 70.510 189.760 ;
        RECT 79.050 188.290 79.310 188.380 ;
        RECT 79.050 188.150 79.710 188.290 ;
        RECT 79.050 188.060 79.310 188.150 ;
        RECT 74.450 186.700 74.710 187.020 ;
        RECT 73.990 186.020 74.250 186.340 ;
        RECT 70.310 183.980 70.570 184.300 ;
        RECT 74.050 181.920 74.190 186.020 ;
        RECT 74.510 184.640 74.650 186.700 ;
        RECT 76.280 186.505 76.560 186.875 ;
        RECT 76.290 186.360 76.550 186.505 ;
        RECT 75.370 185.680 75.630 186.000 ;
        RECT 75.430 184.640 75.570 185.680 ;
        RECT 74.450 184.320 74.710 184.640 ;
        RECT 75.370 184.320 75.630 184.640 ;
        RECT 73.990 181.600 74.250 181.920 ;
        RECT 74.510 181.240 74.650 184.320 ;
        RECT 73.070 180.920 73.330 181.240 ;
        RECT 74.450 180.920 74.710 181.240 ;
        RECT 70.770 180.580 71.030 180.900 ;
        RECT 70.830 178.520 70.970 180.580 ;
        RECT 70.770 178.200 71.030 178.520 ;
        RECT 72.150 177.860 72.410 178.180 ;
        RECT 71.230 177.180 71.490 177.500 ;
        RECT 70.770 174.635 71.030 174.780 ;
        RECT 70.760 174.265 71.040 174.635 ;
        RECT 71.290 173.840 71.430 177.180 ;
        RECT 72.210 175.800 72.350 177.860 ;
        RECT 73.130 175.800 73.270 180.920 ;
        RECT 75.430 178.520 75.570 184.320 ;
        RECT 75.830 181.260 76.090 181.580 ;
        RECT 75.370 178.200 75.630 178.520 ;
        RECT 75.890 178.180 76.030 181.260 ;
        RECT 76.350 178.180 76.490 186.360 ;
        RECT 79.570 186.340 79.710 188.150 ;
        RECT 81.410 187.360 81.550 191.800 ;
        RECT 86.010 191.100 86.150 193.500 ;
        RECT 86.470 192.460 86.610 194.180 ;
        RECT 86.410 192.140 86.670 192.460 ;
        RECT 85.490 190.780 85.750 191.100 ;
        RECT 85.950 190.780 86.210 191.100 ;
        RECT 85.550 189.400 85.690 190.780 ;
        RECT 85.490 189.080 85.750 189.400 ;
        RECT 83.190 188.400 83.450 188.720 ;
        RECT 81.350 187.040 81.610 187.360 ;
        RECT 83.250 187.020 83.390 188.400 ;
        RECT 83.190 186.700 83.450 187.020 ;
        RECT 79.510 186.020 79.770 186.340 ;
        RECT 76.750 185.340 77.010 185.660 ;
        RECT 76.810 183.280 76.950 185.340 ;
        RECT 77.510 184.805 79.390 185.175 ;
        RECT 76.750 182.960 77.010 183.280 ;
        RECT 77.510 179.365 79.390 179.735 ;
        RECT 73.530 177.860 73.790 178.180 ;
        RECT 74.910 177.860 75.170 178.180 ;
        RECT 75.830 177.860 76.090 178.180 ;
        RECT 76.290 177.860 76.550 178.180 ;
        RECT 73.590 176.140 73.730 177.860 ;
        RECT 73.530 175.820 73.790 176.140 ;
        RECT 72.150 175.480 72.410 175.800 ;
        RECT 73.070 175.480 73.330 175.800 ;
        RECT 74.450 175.480 74.710 175.800 ;
        RECT 72.210 175.200 72.350 175.480 ;
        RECT 74.510 175.200 74.650 175.480 ;
        RECT 74.970 175.460 75.110 177.860 ;
        RECT 77.670 177.520 77.930 177.840 ;
        RECT 77.730 175.800 77.870 177.520 ;
        RECT 79.570 177.500 79.710 186.020 ;
        RECT 81.810 185.340 82.070 185.660 ;
        RECT 85.030 185.340 85.290 185.660 ;
        RECT 81.870 183.960 82.010 185.340 ;
        RECT 81.810 183.640 82.070 183.960 ;
        RECT 85.090 183.620 85.230 185.340 ;
        RECT 83.650 183.300 83.910 183.620 ;
        RECT 85.030 183.300 85.290 183.620 ;
        RECT 80.890 182.620 81.150 182.940 ;
        RECT 80.950 179.200 81.090 182.620 ;
        RECT 83.710 181.240 83.850 183.300 ;
        RECT 83.650 180.920 83.910 181.240 ;
        RECT 81.810 179.900 82.070 180.220 ;
        RECT 80.430 178.880 80.690 179.200 ;
        RECT 80.890 178.880 81.150 179.200 ;
        RECT 80.490 178.035 80.630 178.880 ;
        RECT 80.950 178.180 81.090 178.880 ;
        RECT 81.870 178.860 82.010 179.900 ;
        RECT 81.810 178.540 82.070 178.860 ;
        RECT 80.420 177.665 80.700 178.035 ;
        RECT 80.890 177.860 81.150 178.180 ;
        RECT 79.510 177.180 79.770 177.500 ;
        RECT 80.430 177.180 80.690 177.500 ;
        RECT 80.490 175.800 80.630 177.180 ;
        RECT 83.190 175.820 83.450 176.140 ;
        RECT 77.670 175.480 77.930 175.800 ;
        RECT 80.430 175.480 80.690 175.800 ;
        RECT 72.210 175.060 74.650 175.200 ;
        RECT 74.910 175.140 75.170 175.460 ;
        RECT 72.150 174.460 72.410 174.780 ;
        RECT 69.910 173.700 70.510 173.840 ;
        RECT 69.850 172.760 70.110 173.080 ;
        RECT 69.910 171.040 70.050 172.760 ;
        RECT 69.850 170.720 70.110 171.040 ;
        RECT 69.850 163.920 70.110 164.240 ;
        RECT 69.390 162.220 69.650 162.540 ;
        RECT 68.920 160.665 69.200 161.035 ;
        RECT 67.550 159.840 67.810 160.160 ;
        RECT 66.630 159.250 67.290 159.390 ;
        RECT 66.630 159.160 66.890 159.250 ;
        RECT 65.310 158.800 65.450 159.160 ;
        RECT 65.250 158.480 65.510 158.800 ;
        RECT 65.310 156.420 65.450 158.480 ;
        RECT 67.150 156.955 67.290 159.250 ;
        RECT 67.610 159.390 67.750 159.840 ;
        RECT 68.470 159.390 68.730 159.480 ;
        RECT 67.610 159.250 68.730 159.390 ;
        RECT 67.080 156.585 67.360 156.955 ;
        RECT 67.150 156.420 67.290 156.585 ;
        RECT 67.610 156.420 67.750 159.250 ;
        RECT 68.470 159.160 68.730 159.250 ;
        RECT 68.470 158.140 68.730 158.460 ;
        RECT 68.010 156.780 68.270 157.100 ;
        RECT 64.330 156.275 64.590 156.420 ;
        RECT 64.320 155.905 64.600 156.275 ;
        RECT 64.790 156.100 65.050 156.420 ;
        RECT 65.250 156.100 65.510 156.420 ;
        RECT 62.510 154.885 64.390 155.255 ;
        RECT 62.090 153.810 62.690 153.950 ;
        RECT 62.020 153.185 62.300 153.555 ;
        RECT 62.030 153.040 62.290 153.185 ;
        RECT 61.630 152.740 62.230 152.880 ;
        RECT 60.650 150.660 60.910 150.980 ;
        RECT 58.810 148.960 59.070 149.280 ;
        RECT 59.330 149.220 59.930 149.360 ;
        RECT 58.870 145.880 59.010 148.960 ;
        RECT 58.350 145.560 58.610 145.880 ;
        RECT 58.810 145.560 59.070 145.880 ;
        RECT 59.330 145.540 59.470 149.220 ;
        RECT 59.730 148.620 59.990 148.940 ;
        RECT 59.270 145.220 59.530 145.540 ;
        RECT 58.810 144.540 59.070 144.860 ;
        RECT 58.350 142.840 58.610 143.160 ;
        RECT 58.410 139.420 58.550 142.840 ;
        RECT 58.870 142.140 59.010 144.540 ;
        RECT 59.270 142.840 59.530 143.160 ;
        RECT 58.810 141.820 59.070 142.140 ;
        RECT 58.870 140.440 59.010 141.820 ;
        RECT 59.330 141.120 59.470 142.840 ;
        RECT 59.270 140.800 59.530 141.120 ;
        RECT 58.810 140.120 59.070 140.440 ;
        RECT 58.350 139.100 58.610 139.420 ;
        RECT 55.130 130.940 55.390 131.260 ;
        RECT 55.190 129.220 55.330 130.940 ;
        RECT 55.650 129.900 55.790 131.540 ;
        RECT 57.890 131.280 58.150 131.600 ;
        RECT 55.590 129.580 55.850 129.900 ;
        RECT 55.130 128.900 55.390 129.220 ;
        RECT 58.410 128.540 58.550 139.100 ;
        RECT 56.970 128.220 57.230 128.540 ;
        RECT 58.350 128.220 58.610 128.540 ;
        RECT 57.030 126.840 57.170 128.220 ;
        RECT 58.410 127.520 58.550 128.220 ;
        RECT 58.350 127.200 58.610 127.520 ;
        RECT 56.970 126.520 57.230 126.840 ;
        RECT 56.510 125.500 56.770 125.820 ;
        RECT 56.570 124.120 56.710 125.500 ;
        RECT 56.510 123.800 56.770 124.120 ;
        RECT 55.590 123.120 55.850 123.440 ;
        RECT 55.650 122.080 55.790 123.120 ;
        RECT 56.510 122.780 56.770 123.100 ;
        RECT 55.590 121.760 55.850 122.080 ;
        RECT 56.050 121.080 56.310 121.400 ;
        RECT 56.110 115.960 56.250 121.080 ;
        RECT 56.570 121.060 56.710 122.780 ;
        RECT 56.510 120.740 56.770 121.060 ;
        RECT 56.570 118.340 56.710 120.740 ;
        RECT 56.510 118.020 56.770 118.340 ;
        RECT 56.050 115.640 56.310 115.960 ;
        RECT 56.570 113.580 56.710 118.020 ;
        RECT 56.970 115.300 57.230 115.620 ;
        RECT 56.510 113.260 56.770 113.580 ;
        RECT 57.030 113.240 57.170 115.300 ;
        RECT 56.970 112.920 57.230 113.240 ;
        RECT 59.790 112.900 59.930 148.620 ;
        RECT 60.190 147.940 60.450 148.260 ;
        RECT 60.250 113.240 60.390 147.940 ;
        RECT 60.710 147.580 60.850 150.660 ;
        RECT 61.110 150.320 61.370 150.640 ;
        RECT 61.570 150.320 61.830 150.640 ;
        RECT 61.170 148.115 61.310 150.320 ;
        RECT 61.630 149.280 61.770 150.320 ;
        RECT 62.090 150.300 62.230 152.740 ;
        RECT 62.550 151.660 62.690 153.810 ;
        RECT 63.410 153.720 63.670 154.040 ;
        RECT 63.870 153.720 64.130 154.040 ;
        RECT 62.490 151.340 62.750 151.660 ;
        RECT 62.550 150.300 62.690 151.340 ;
        RECT 63.470 150.980 63.610 153.720 ;
        RECT 63.930 153.360 64.070 153.720 ;
        RECT 64.850 153.700 64.990 156.100 ;
        RECT 66.160 155.905 66.440 156.275 ;
        RECT 67.090 156.100 67.350 156.420 ;
        RECT 67.550 156.100 67.810 156.420 ;
        RECT 65.710 155.420 65.970 155.740 ;
        RECT 65.240 153.865 65.520 154.235 ;
        RECT 65.250 153.720 65.510 153.865 ;
        RECT 64.790 153.380 65.050 153.700 ;
        RECT 63.870 153.040 64.130 153.360 ;
        RECT 63.930 150.980 64.070 153.040 ;
        RECT 65.770 153.020 65.910 155.420 ;
        RECT 66.230 153.700 66.370 155.905 ;
        RECT 68.070 155.650 68.210 156.780 ;
        RECT 67.610 155.510 68.210 155.650 ;
        RECT 66.630 153.720 66.890 154.040 ;
        RECT 66.170 153.380 66.430 153.700 ;
        RECT 65.710 152.700 65.970 153.020 ;
        RECT 63.410 150.660 63.670 150.980 ;
        RECT 63.870 150.890 64.130 150.980 ;
        RECT 63.870 150.750 65.450 150.890 ;
        RECT 63.870 150.660 64.130 150.750 ;
        RECT 62.030 149.980 62.290 150.300 ;
        RECT 62.490 149.980 62.750 150.300 ;
        RECT 61.570 148.960 61.830 149.280 ;
        RECT 61.100 147.745 61.380 148.115 ;
        RECT 62.090 147.920 62.230 149.980 ;
        RECT 62.510 149.445 64.390 149.815 ;
        RECT 62.490 148.620 62.750 148.940 ;
        RECT 62.030 147.600 62.290 147.920 ;
        RECT 60.650 147.260 60.910 147.580 ;
        RECT 60.710 142.140 60.850 147.260 ;
        RECT 62.550 146.560 62.690 148.620 ;
        RECT 62.490 146.240 62.750 146.560 ;
        RECT 64.790 145.900 65.050 146.220 ;
        RECT 62.030 145.220 62.290 145.540 ;
        RECT 60.650 141.820 60.910 142.140 ;
        RECT 62.090 140.100 62.230 145.220 ;
        RECT 64.850 144.860 64.990 145.900 ;
        RECT 64.790 144.540 65.050 144.860 ;
        RECT 62.510 144.005 64.390 144.375 ;
        RECT 62.950 143.180 63.210 143.500 ;
        RECT 63.010 141.120 63.150 143.180 ;
        RECT 62.950 140.800 63.210 141.120 ;
        RECT 62.030 139.780 62.290 140.100 ;
        RECT 62.090 134.910 62.230 139.780 ;
        RECT 62.510 138.565 64.390 138.935 ;
        RECT 64.850 137.040 64.990 144.540 ;
        RECT 65.310 143.840 65.450 150.750 ;
        RECT 65.250 143.520 65.510 143.840 ;
        RECT 64.790 136.720 65.050 137.040 ;
        RECT 64.850 135.340 64.990 136.720 ;
        RECT 61.170 134.770 62.230 134.910 ;
        RECT 64.320 134.825 64.600 135.195 ;
        RECT 64.790 135.020 65.050 135.340 ;
        RECT 61.170 123.520 61.310 134.770 ;
        RECT 64.390 134.660 64.530 134.825 ;
        RECT 64.330 134.400 64.590 134.660 ;
        RECT 64.330 134.340 64.990 134.400 ;
        RECT 62.030 134.000 62.290 134.320 ;
        RECT 64.390 134.260 64.990 134.340 ;
        RECT 62.090 132.960 62.230 134.000 ;
        RECT 62.510 133.125 64.390 133.495 ;
        RECT 62.030 132.640 62.290 132.960 ;
        RECT 62.090 129.900 62.230 132.640 ;
        RECT 64.850 132.280 64.990 134.260 ;
        RECT 63.410 131.960 63.670 132.280 ;
        RECT 64.790 131.960 65.050 132.280 ;
        RECT 63.470 131.260 63.610 131.960 ;
        RECT 63.410 130.940 63.670 131.260 ;
        RECT 62.030 129.580 62.290 129.900 ;
        RECT 63.470 128.880 63.610 130.940 ;
        RECT 64.850 129.220 64.990 131.960 ;
        RECT 66.230 131.940 66.370 153.380 ;
        RECT 66.690 145.880 66.830 153.720 ;
        RECT 67.610 152.080 67.750 155.510 ;
        RECT 68.010 154.060 68.270 154.380 ;
        RECT 67.150 152.000 67.750 152.080 ;
        RECT 67.090 151.940 67.750 152.000 ;
        RECT 67.090 151.680 67.350 151.940 ;
        RECT 68.070 150.980 68.210 154.060 ;
        RECT 68.010 150.660 68.270 150.980 ;
        RECT 67.090 147.940 67.350 148.260 ;
        RECT 68.010 147.940 68.270 148.260 ;
        RECT 67.150 146.560 67.290 147.940 ;
        RECT 67.090 146.240 67.350 146.560 ;
        RECT 66.630 145.560 66.890 145.880 ;
        RECT 68.070 143.160 68.210 147.940 ;
        RECT 68.530 145.540 68.670 158.140 ;
        RECT 68.990 154.720 69.130 160.665 ;
        RECT 69.450 160.160 69.590 162.220 ;
        RECT 69.910 161.520 70.050 163.920 ;
        RECT 69.850 161.200 70.110 161.520 ;
        RECT 69.390 159.840 69.650 160.160 ;
        RECT 69.840 159.985 70.120 160.355 ;
        RECT 69.910 159.820 70.050 159.985 ;
        RECT 69.850 159.500 70.110 159.820 ;
        RECT 70.370 159.675 70.510 173.700 ;
        RECT 70.830 173.700 71.430 173.840 ;
        RECT 70.300 159.305 70.580 159.675 ;
        RECT 69.850 158.820 70.110 159.140 ;
        RECT 69.390 158.140 69.650 158.460 ;
        RECT 68.930 154.400 69.190 154.720 ;
        RECT 68.990 153.020 69.130 154.400 ;
        RECT 68.930 152.700 69.190 153.020 ;
        RECT 68.930 150.155 69.190 150.300 ;
        RECT 68.920 149.785 69.200 150.155 ;
        RECT 68.470 145.220 68.730 145.540 ;
        RECT 68.010 142.840 68.270 143.160 ;
        RECT 66.630 142.500 66.890 142.820 ;
        RECT 66.690 141.120 66.830 142.500 ;
        RECT 66.630 140.800 66.890 141.120 ;
        RECT 67.550 136.380 67.810 136.700 ;
        RECT 67.610 132.960 67.750 136.380 ;
        RECT 68.070 134.320 68.210 142.840 ;
        RECT 68.460 138.225 68.740 138.595 ;
        RECT 68.530 137.380 68.670 138.225 ;
        RECT 69.450 137.720 69.590 158.140 ;
        RECT 69.910 156.760 70.050 158.820 ;
        RECT 69.850 156.440 70.110 156.760 ;
        RECT 69.850 155.420 70.110 155.740 ;
        RECT 69.910 150.980 70.050 155.420 ;
        RECT 70.370 154.040 70.510 159.305 ;
        RECT 70.310 153.720 70.570 154.040 ;
        RECT 69.850 150.660 70.110 150.980 ;
        RECT 70.370 148.600 70.510 153.720 ;
        RECT 70.830 151.320 70.970 173.700 ;
        RECT 71.690 170.040 71.950 170.360 ;
        RECT 71.750 167.300 71.890 170.040 ;
        RECT 71.690 166.980 71.950 167.300 ;
        RECT 71.750 165.600 71.890 166.980 ;
        RECT 71.690 165.280 71.950 165.600 ;
        RECT 71.230 164.940 71.490 165.260 ;
        RECT 71.290 161.180 71.430 164.940 ;
        RECT 71.230 160.860 71.490 161.180 ;
        RECT 71.290 159.480 71.430 160.860 ;
        RECT 71.750 159.820 71.890 165.280 ;
        RECT 71.690 159.500 71.950 159.820 ;
        RECT 71.230 159.160 71.490 159.480 ;
        RECT 70.770 151.000 71.030 151.320 ;
        RECT 70.310 148.280 70.570 148.600 ;
        RECT 71.690 147.260 71.950 147.580 ;
        RECT 71.230 146.240 71.490 146.560 ;
        RECT 70.760 145.705 71.040 146.075 ;
        RECT 70.770 145.560 71.030 145.705 ;
        RECT 70.770 144.540 71.030 144.860 ;
        RECT 70.830 140.440 70.970 144.540 ;
        RECT 70.770 140.120 71.030 140.440 ;
        RECT 70.770 139.440 71.030 139.760 ;
        RECT 69.390 137.400 69.650 137.720 ;
        RECT 68.470 137.060 68.730 137.380 ;
        RECT 69.850 136.380 70.110 136.700 ;
        RECT 68.470 134.340 68.730 134.660 ;
        RECT 68.010 134.000 68.270 134.320 ;
        RECT 67.550 132.640 67.810 132.960 ;
        RECT 68.530 132.280 68.670 134.340 ;
        RECT 68.470 131.960 68.730 132.280 ;
        RECT 66.170 131.620 66.430 131.940 ;
        RECT 65.710 131.280 65.970 131.600 ;
        RECT 64.790 128.900 65.050 129.220 ;
        RECT 62.030 128.560 62.290 128.880 ;
        RECT 63.410 128.560 63.670 128.880 ;
        RECT 61.570 128.220 61.830 128.540 ;
        RECT 61.630 124.120 61.770 128.220 ;
        RECT 62.090 127.520 62.230 128.560 ;
        RECT 62.510 127.685 64.390 128.055 ;
        RECT 65.770 127.520 65.910 131.280 ;
        RECT 62.030 127.200 62.290 127.520 ;
        RECT 65.710 127.200 65.970 127.520 ;
        RECT 62.490 126.860 62.750 127.180 ;
        RECT 62.550 124.800 62.690 126.860 ;
        RECT 64.330 126.180 64.590 126.500 ;
        RECT 64.390 124.800 64.530 126.180 ;
        RECT 62.490 124.480 62.750 124.800 ;
        RECT 64.330 124.480 64.590 124.800 ;
        RECT 61.570 123.800 61.830 124.120 ;
        RECT 65.770 123.780 65.910 127.200 ;
        RECT 62.030 123.520 62.290 123.780 ;
        RECT 61.170 123.460 62.290 123.520 ;
        RECT 65.710 123.460 65.970 123.780 ;
        RECT 61.170 123.380 62.230 123.460 ;
        RECT 62.090 121.400 62.230 123.380 ;
        RECT 62.510 122.245 64.390 122.615 ;
        RECT 62.030 121.080 62.290 121.400 ;
        RECT 65.770 118.340 65.910 123.460 ;
        RECT 65.710 118.020 65.970 118.340 ;
        RECT 62.510 116.805 64.390 117.175 ;
        RECT 66.230 116.640 66.370 131.620 ;
        RECT 68.530 129.560 68.670 131.960 ;
        RECT 68.470 129.240 68.730 129.560 ;
        RECT 68.530 125.820 68.670 129.240 ;
        RECT 66.630 125.500 66.890 125.820 ;
        RECT 68.470 125.500 68.730 125.820 ;
        RECT 66.690 121.400 66.830 125.500 ;
        RECT 68.470 122.780 68.730 123.100 ;
        RECT 68.530 121.740 68.670 122.780 ;
        RECT 68.470 121.420 68.730 121.740 ;
        RECT 66.630 121.080 66.890 121.400 ;
        RECT 66.170 116.320 66.430 116.640 ;
        RECT 69.910 116.300 70.050 136.380 ;
        RECT 70.830 132.960 70.970 139.440 ;
        RECT 71.290 135.680 71.430 146.240 ;
        RECT 71.750 145.540 71.890 147.260 ;
        RECT 71.690 145.220 71.950 145.540 ;
        RECT 71.690 140.350 71.950 140.440 ;
        RECT 72.210 140.350 72.350 174.460 ;
        RECT 77.510 173.925 79.390 174.295 ;
        RECT 77.210 171.740 77.470 172.060 ;
        RECT 77.270 170.360 77.410 171.740 ;
        RECT 83.250 171.040 83.390 175.820 ;
        RECT 83.710 175.460 83.850 180.920 ;
        RECT 84.110 180.240 84.370 180.560 ;
        RECT 84.170 178.180 84.310 180.240 ;
        RECT 84.560 178.345 84.840 178.715 ;
        RECT 84.630 178.180 84.770 178.345 ;
        RECT 84.110 177.860 84.370 178.180 ;
        RECT 84.570 177.860 84.830 178.180 ;
        RECT 85.030 177.520 85.290 177.840 ;
        RECT 84.110 175.820 84.370 176.140 ;
        RECT 83.650 175.140 83.910 175.460 ;
        RECT 83.710 173.080 83.850 175.140 ;
        RECT 84.170 173.760 84.310 175.820 ;
        RECT 84.110 173.440 84.370 173.760 ;
        RECT 83.650 172.760 83.910 173.080 ;
        RECT 84.110 172.760 84.370 173.080 ;
        RECT 83.190 170.720 83.450 171.040 ;
        RECT 79.510 170.380 79.770 170.700 ;
        RECT 77.210 170.040 77.470 170.360 ;
        RECT 73.070 169.700 73.330 170.020 ;
        RECT 72.610 169.020 72.870 169.340 ;
        RECT 72.670 164.580 72.810 169.020 ;
        RECT 72.610 164.260 72.870 164.580 ;
        RECT 72.670 162.200 72.810 164.260 ;
        RECT 72.610 161.880 72.870 162.200 ;
        RECT 72.610 160.860 72.870 161.180 ;
        RECT 72.670 159.480 72.810 160.860 ;
        RECT 72.610 159.160 72.870 159.480 ;
        RECT 72.610 158.480 72.870 158.800 ;
        RECT 72.670 156.420 72.810 158.480 ;
        RECT 73.130 156.760 73.270 169.700 ;
        RECT 77.510 168.485 79.390 168.855 ;
        RECT 75.830 166.980 76.090 167.300 ;
        RECT 75.890 165.600 76.030 166.980 ;
        RECT 79.570 166.620 79.710 170.380 ;
        RECT 83.710 170.360 83.850 172.760 ;
        RECT 83.650 170.040 83.910 170.360 ;
        RECT 83.710 168.320 83.850 170.040 ;
        RECT 83.650 168.000 83.910 168.320 ;
        RECT 82.270 167.320 82.530 167.640 ;
        RECT 81.810 166.640 82.070 166.960 ;
        RECT 77.210 166.300 77.470 166.620 ;
        RECT 79.510 166.300 79.770 166.620 ;
        RECT 77.270 165.600 77.410 166.300 ;
        RECT 75.830 165.280 76.090 165.600 ;
        RECT 77.210 165.280 77.470 165.600 ;
        RECT 79.570 164.920 79.710 166.300 ;
        RECT 80.890 164.940 81.150 165.260 ;
        RECT 79.510 164.600 79.770 164.920 ;
        RECT 76.750 163.580 77.010 163.900 ;
        RECT 76.810 161.520 76.950 163.580 ;
        RECT 77.510 163.045 79.390 163.415 ;
        RECT 76.750 161.200 77.010 161.520 ;
        RECT 79.570 159.480 79.710 164.600 ;
        RECT 80.430 161.540 80.690 161.860 ;
        RECT 80.490 160.160 80.630 161.540 ;
        RECT 80.950 160.160 81.090 164.940 ;
        RECT 80.430 159.840 80.690 160.160 ;
        RECT 80.890 159.840 81.150 160.160 ;
        RECT 81.870 159.480 82.010 166.640 ;
        RECT 82.330 162.200 82.470 167.320 ;
        RECT 82.730 163.920 82.990 164.240 ;
        RECT 82.790 162.540 82.930 163.920 ;
        RECT 82.730 162.220 82.990 162.540 ;
        RECT 84.170 162.200 84.310 172.760 ;
        RECT 85.090 172.740 85.230 177.520 ;
        RECT 86.010 175.460 86.150 190.780 ;
        RECT 86.930 189.060 87.070 196.900 ;
        RECT 95.670 194.840 95.810 196.900 ;
        RECT 97.450 196.220 97.710 196.540 ;
        RECT 95.610 194.520 95.870 194.840 ;
        RECT 91.470 194.180 91.730 194.500 ;
        RECT 89.170 193.500 89.430 193.820 ;
        RECT 89.230 192.800 89.370 193.500 ;
        RECT 89.170 192.480 89.430 192.800 ;
        RECT 89.230 189.400 89.370 192.480 ;
        RECT 91.530 190.080 91.670 194.180 ;
        RECT 91.930 193.500 92.190 193.820 ;
        RECT 91.990 192.460 92.130 193.500 ;
        RECT 92.510 192.965 94.390 193.335 ;
        RECT 91.930 192.140 92.190 192.460 ;
        RECT 91.470 189.760 91.730 190.080 ;
        RECT 88.250 189.080 88.510 189.400 ;
        RECT 89.170 189.080 89.430 189.400 ;
        RECT 86.870 188.740 87.130 189.060 ;
        RECT 86.930 181.920 87.070 188.740 ;
        RECT 88.310 187.360 88.450 189.080 ;
        RECT 95.150 188.060 95.410 188.380 ;
        RECT 92.510 187.525 94.390 187.895 ;
        RECT 88.250 187.040 88.510 187.360 ;
        RECT 87.320 186.590 87.600 186.875 ;
        RECT 87.320 186.505 87.990 186.590 ;
        RECT 87.330 186.450 87.990 186.505 ;
        RECT 87.330 186.360 87.590 186.450 ;
        RECT 87.850 183.620 87.990 186.450 ;
        RECT 88.310 184.640 88.450 187.040 ;
        RECT 95.210 186.680 95.350 188.060 ;
        RECT 95.150 186.360 95.410 186.680 ;
        RECT 90.550 186.020 90.810 186.340 ;
        RECT 90.610 184.640 90.750 186.020 ;
        RECT 94.690 185.340 94.950 185.660 ;
        RECT 88.250 184.320 88.510 184.640 ;
        RECT 90.550 184.320 90.810 184.640 ;
        RECT 87.790 183.300 88.050 183.620 ;
        RECT 86.870 181.600 87.130 181.920 ;
        RECT 87.850 177.840 87.990 183.300 ;
        RECT 89.170 181.260 89.430 181.580 ;
        RECT 89.230 179.200 89.370 181.260 ;
        RECT 89.170 178.880 89.430 179.200 ;
        RECT 90.090 178.035 90.350 178.180 ;
        RECT 90.610 178.090 90.750 184.320 ;
        RECT 92.510 182.085 94.390 182.455 ;
        RECT 94.750 181.240 94.890 185.340 ;
        RECT 95.150 182.620 95.410 182.940 ;
        RECT 94.690 180.920 94.950 181.240 ;
        RECT 95.210 180.900 95.350 182.620 ;
        RECT 95.150 180.580 95.410 180.900 ;
        RECT 91.470 179.900 91.730 180.220 ;
        RECT 91.000 179.025 91.280 179.395 ;
        RECT 91.070 178.860 91.210 179.025 ;
        RECT 91.010 178.540 91.270 178.860 ;
        RECT 91.010 178.090 91.270 178.180 ;
        RECT 87.790 177.520 88.050 177.840 ;
        RECT 90.080 177.665 90.360 178.035 ;
        RECT 90.610 177.950 91.270 178.090 ;
        RECT 91.010 177.860 91.270 177.950 ;
        RECT 90.090 177.180 90.350 177.500 ;
        RECT 85.950 175.140 86.210 175.460 ;
        RECT 89.630 174.460 89.890 174.780 ;
        RECT 89.690 172.740 89.830 174.460 ;
        RECT 85.030 172.420 85.290 172.740 ;
        RECT 89.630 172.420 89.890 172.740 ;
        RECT 86.870 171.740 87.130 172.060 ;
        RECT 86.930 170.360 87.070 171.740 ;
        RECT 89.170 170.720 89.430 171.040 ;
        RECT 86.870 170.040 87.130 170.360 ;
        RECT 88.710 166.980 88.970 167.300 ;
        RECT 86.870 166.300 87.130 166.620 ;
        RECT 86.930 164.920 87.070 166.300 ;
        RECT 86.870 164.600 87.130 164.920 ;
        RECT 88.250 164.600 88.510 164.920 ;
        RECT 84.570 163.580 84.830 163.900 ;
        RECT 82.270 161.880 82.530 162.200 ;
        RECT 84.110 161.880 84.370 162.200 ;
        RECT 84.630 161.180 84.770 163.580 ;
        RECT 88.310 161.860 88.450 164.600 ;
        RECT 88.770 162.880 88.910 166.980 ;
        RECT 88.710 162.560 88.970 162.880 ;
        RECT 88.250 161.540 88.510 161.860 ;
        RECT 84.570 160.860 84.830 161.180 ;
        RECT 79.510 159.160 79.770 159.480 ;
        RECT 81.810 159.160 82.070 159.480 ;
        RECT 81.870 158.995 82.010 159.160 ;
        RECT 81.800 158.625 82.080 158.995 ;
        RECT 83.190 158.820 83.450 159.140 ;
        RECT 77.510 157.605 79.390 157.975 ;
        RECT 73.070 156.440 73.330 156.760 ;
        RECT 72.610 156.100 72.870 156.420 ;
        RECT 72.610 155.420 72.870 155.740 ;
        RECT 71.690 140.210 72.350 140.350 ;
        RECT 71.690 140.120 71.950 140.210 ;
        RECT 72.670 140.100 72.810 155.420 ;
        RECT 80.430 153.720 80.690 154.040 ;
        RECT 76.750 153.040 77.010 153.360 ;
        RECT 79.970 153.040 80.230 153.360 ;
        RECT 73.990 151.680 74.250 152.000 ;
        RECT 73.070 150.660 73.330 150.980 ;
        RECT 73.530 150.660 73.790 150.980 ;
        RECT 73.130 147.920 73.270 150.660 ;
        RECT 73.590 149.280 73.730 150.660 ;
        RECT 73.530 148.960 73.790 149.280 ;
        RECT 73.530 148.280 73.790 148.600 ;
        RECT 73.070 147.600 73.330 147.920 ;
        RECT 72.610 139.780 72.870 140.100 ;
        RECT 71.690 139.440 71.950 139.760 ;
        RECT 71.230 135.360 71.490 135.680 ;
        RECT 71.230 134.680 71.490 135.000 ;
        RECT 70.770 132.640 71.030 132.960 ;
        RECT 70.310 131.620 70.570 131.940 ;
        RECT 70.370 126.500 70.510 131.620 ;
        RECT 71.290 128.880 71.430 134.680 ;
        RECT 71.230 128.560 71.490 128.880 ;
        RECT 71.290 126.840 71.430 128.560 ;
        RECT 71.230 126.520 71.490 126.840 ;
        RECT 70.310 126.180 70.570 126.500 ;
        RECT 70.370 124.800 70.510 126.180 ;
        RECT 70.310 124.480 70.570 124.800 ;
        RECT 70.370 117.660 70.510 124.480 ;
        RECT 70.770 123.120 71.030 123.440 ;
        RECT 70.830 119.360 70.970 123.120 ;
        RECT 71.290 122.080 71.430 126.520 ;
        RECT 71.230 121.760 71.490 122.080 ;
        RECT 70.770 119.040 71.030 119.360 ;
        RECT 70.310 117.340 70.570 117.660 ;
        RECT 69.850 115.980 70.110 116.300 ;
        RECT 70.770 115.640 71.030 115.960 ;
        RECT 60.190 112.920 60.450 113.240 ;
        RECT 54.210 112.580 54.470 112.900 ;
        RECT 59.730 112.580 59.990 112.900 ;
        RECT 52.830 112.240 53.090 112.560 ;
        RECT 56.050 112.240 56.310 112.560 ;
        RECT 66.630 112.240 66.890 112.560 ;
        RECT 70.310 112.240 70.570 112.560 ;
        RECT 50.070 110.540 50.330 110.860 ;
        RECT 48.690 110.200 48.950 110.520 ;
        RECT 47.510 108.645 49.390 109.015 ;
        RECT 50.130 108.480 50.270 110.540 ;
        RECT 51.450 110.200 51.710 110.520 ;
        RECT 46.850 108.160 47.110 108.480 ;
        RECT 50.070 108.160 50.330 108.480 ;
        RECT 51.510 96.255 51.650 110.200 ;
        RECT 52.890 107.460 53.030 112.240 ;
        RECT 52.830 107.140 53.090 107.460 ;
        RECT 56.110 107.120 56.250 112.240 ;
        RECT 56.510 111.900 56.770 112.220 ;
        RECT 59.270 111.900 59.530 112.220 ;
        RECT 59.730 111.900 59.990 112.220 ;
        RECT 56.570 110.860 56.710 111.900 ;
        RECT 59.330 110.860 59.470 111.900 ;
        RECT 56.510 110.540 56.770 110.860 ;
        RECT 59.270 110.540 59.530 110.860 ;
        RECT 59.790 107.800 59.930 111.900 ;
        RECT 62.510 111.365 64.390 111.735 ;
        RECT 61.570 110.200 61.830 110.520 ;
        RECT 61.110 109.860 61.370 110.180 ;
        RECT 61.170 107.800 61.310 109.860 ;
        RECT 56.510 107.480 56.770 107.800 ;
        RECT 59.730 107.480 59.990 107.800 ;
        RECT 61.110 107.480 61.370 107.800 ;
        RECT 56.050 106.800 56.310 107.120 ;
        RECT 56.570 96.255 56.710 107.480 ;
        RECT 61.630 96.255 61.770 110.200 ;
        RECT 62.510 105.925 64.390 106.295 ;
        RECT 66.690 96.255 66.830 112.240 ;
        RECT 68.470 111.900 68.730 112.220 ;
        RECT 68.530 110.860 68.670 111.900 ;
        RECT 68.470 110.540 68.730 110.860 ;
        RECT 70.370 108.480 70.510 112.240 ;
        RECT 70.310 108.160 70.570 108.480 ;
        RECT 70.830 107.800 70.970 115.640 ;
        RECT 71.750 110.520 71.890 139.440 ;
        RECT 73.130 138.400 73.270 147.600 ;
        RECT 73.590 146.220 73.730 148.280 ;
        RECT 73.530 145.900 73.790 146.220 ;
        RECT 73.530 140.460 73.790 140.780 ;
        RECT 73.070 138.080 73.330 138.400 ;
        RECT 72.150 137.400 72.410 137.720 ;
        RECT 72.610 137.400 72.870 137.720 ;
        RECT 72.210 132.280 72.350 137.400 ;
        RECT 72.670 136.700 72.810 137.400 ;
        RECT 72.610 136.380 72.870 136.700 ;
        RECT 72.670 132.280 72.810 136.380 ;
        RECT 73.070 134.000 73.330 134.320 ;
        RECT 73.130 132.960 73.270 134.000 ;
        RECT 73.070 132.640 73.330 132.960 ;
        RECT 72.150 131.960 72.410 132.280 ;
        RECT 72.610 131.960 72.870 132.280 ;
        RECT 73.130 129.640 73.270 132.640 ;
        RECT 72.210 129.560 73.270 129.640 ;
        RECT 72.210 129.500 73.330 129.560 ;
        RECT 72.210 127.180 72.350 129.500 ;
        RECT 73.070 129.240 73.330 129.500 ;
        RECT 72.610 128.560 72.870 128.880 ;
        RECT 72.150 126.860 72.410 127.180 ;
        RECT 72.670 126.500 72.810 128.560 ;
        RECT 72.610 126.180 72.870 126.500 ;
        RECT 72.670 124.800 72.810 126.180 ;
        RECT 72.610 124.480 72.870 124.800 ;
        RECT 72.670 118.680 72.810 124.480 ;
        RECT 73.130 124.120 73.270 129.240 ;
        RECT 73.590 127.520 73.730 140.460 ;
        RECT 74.050 131.600 74.190 151.680 ;
        RECT 76.290 151.340 76.550 151.660 ;
        RECT 75.830 151.000 76.090 151.320 ;
        RECT 75.370 150.660 75.630 150.980 ;
        RECT 74.910 148.960 75.170 149.280 ;
        RECT 74.450 148.620 74.710 148.940 ;
        RECT 74.510 146.560 74.650 148.620 ;
        RECT 74.450 146.240 74.710 146.560 ;
        RECT 74.970 140.440 75.110 148.960 ;
        RECT 75.430 148.600 75.570 150.660 ;
        RECT 75.370 148.280 75.630 148.600 ;
        RECT 75.370 143.180 75.630 143.500 ;
        RECT 74.910 140.120 75.170 140.440 ;
        RECT 74.970 138.060 75.110 140.120 ;
        RECT 75.430 139.420 75.570 143.180 ;
        RECT 75.370 139.100 75.630 139.420 ;
        RECT 74.910 137.740 75.170 138.060 ;
        RECT 74.450 136.720 74.710 137.040 ;
        RECT 74.510 132.280 74.650 136.720 ;
        RECT 75.430 132.620 75.570 139.100 ;
        RECT 75.890 136.700 76.030 151.000 ;
        RECT 76.350 148.260 76.490 151.340 ;
        RECT 76.810 150.835 76.950 153.040 ;
        RECT 79.510 152.700 79.770 153.020 ;
        RECT 77.510 152.165 79.390 152.535 ;
        RECT 76.740 150.465 77.020 150.835 ;
        RECT 78.130 149.980 78.390 150.300 ;
        RECT 78.190 148.940 78.330 149.980 ;
        RECT 78.130 148.620 78.390 148.940 ;
        RECT 76.290 147.940 76.550 148.260 ;
        RECT 76.350 140.780 76.490 147.940 ;
        RECT 77.510 146.725 79.390 147.095 ;
        RECT 79.570 145.200 79.710 152.700 ;
        RECT 80.030 150.640 80.170 153.040 ;
        RECT 79.970 150.320 80.230 150.640 ;
        RECT 80.490 149.280 80.630 153.720 ;
        RECT 82.730 152.700 82.990 153.020 ;
        RECT 82.790 151.320 82.930 152.700 ;
        RECT 82.730 151.000 82.990 151.320 ;
        RECT 83.250 150.300 83.390 158.820 ;
        RECT 84.630 156.420 84.770 160.860 ;
        RECT 85.030 159.500 85.290 159.820 ;
        RECT 85.090 156.420 85.230 159.500 ;
        RECT 88.310 158.460 88.450 161.540 ;
        RECT 88.250 158.140 88.510 158.460 ;
        RECT 85.490 157.120 85.750 157.440 ;
        RECT 85.550 156.420 85.690 157.120 ;
        RECT 84.570 156.100 84.830 156.420 ;
        RECT 85.030 156.100 85.290 156.420 ;
        RECT 85.490 156.275 85.750 156.420 ;
        RECT 85.090 155.740 85.230 156.100 ;
        RECT 85.480 155.905 85.760 156.275 ;
        RECT 85.030 155.420 85.290 155.740 ;
        RECT 84.570 154.060 84.830 154.380 ;
        RECT 86.870 154.060 87.130 154.380 ;
        RECT 84.630 151.660 84.770 154.060 ;
        RECT 86.930 152.000 87.070 154.060 ;
        RECT 88.310 153.700 88.450 158.140 ;
        RECT 88.710 155.420 88.970 155.740 ;
        RECT 88.250 153.380 88.510 153.700 ;
        RECT 86.870 151.680 87.130 152.000 ;
        RECT 87.790 151.680 88.050 152.000 ;
        RECT 84.570 151.340 84.830 151.660 ;
        RECT 84.570 150.660 84.830 150.980 ;
        RECT 83.190 149.980 83.450 150.300 ;
        RECT 80.430 148.960 80.690 149.280 ;
        RECT 83.250 147.920 83.390 149.980 ;
        RECT 84.110 147.940 84.370 148.260 ;
        RECT 83.190 147.600 83.450 147.920 ;
        RECT 79.970 147.260 80.230 147.580 ;
        RECT 79.510 144.880 79.770 145.200 ;
        RECT 80.030 143.160 80.170 147.260 ;
        RECT 81.350 145.220 81.610 145.540 ;
        RECT 81.410 143.840 81.550 145.220 ;
        RECT 81.350 143.520 81.610 143.840 ;
        RECT 79.970 142.840 80.230 143.160 ;
        RECT 84.170 142.480 84.310 147.940 ;
        RECT 84.630 145.880 84.770 150.660 ;
        RECT 84.570 145.560 84.830 145.880 ;
        RECT 84.110 142.160 84.370 142.480 ;
        RECT 77.510 141.285 79.390 141.655 ;
        RECT 76.290 140.460 76.550 140.780 ;
        RECT 84.630 140.100 84.770 145.560 ;
        RECT 87.850 145.280 87.990 151.680 ;
        RECT 88.770 145.540 88.910 155.420 ;
        RECT 89.230 152.880 89.370 170.720 ;
        RECT 89.690 157.440 89.830 172.420 ;
        RECT 89.630 157.120 89.890 157.440 ;
        RECT 89.620 156.585 89.900 156.955 ;
        RECT 89.690 156.420 89.830 156.585 ;
        RECT 89.630 156.100 89.890 156.420 ;
        RECT 89.230 152.740 89.830 152.880 ;
        RECT 89.690 151.320 89.830 152.740 ;
        RECT 89.630 151.000 89.890 151.320 ;
        RECT 89.170 150.660 89.430 150.980 ;
        RECT 89.230 149.280 89.370 150.660 ;
        RECT 89.170 148.960 89.430 149.280 ;
        RECT 89.630 146.240 89.890 146.560 ;
        RECT 87.850 145.140 88.450 145.280 ;
        RECT 88.710 145.220 88.970 145.540 ;
        RECT 87.790 144.540 88.050 144.860 ;
        RECT 87.320 142.985 87.600 143.355 ;
        RECT 87.330 142.840 87.590 142.985 ;
        RECT 86.860 142.305 87.140 142.675 ;
        RECT 86.930 142.140 87.070 142.305 ;
        RECT 86.870 141.820 87.130 142.140 ;
        RECT 87.330 141.820 87.590 142.140 ;
        RECT 85.950 140.800 86.210 141.120 ;
        RECT 85.490 140.120 85.750 140.440 ;
        RECT 84.570 139.780 84.830 140.100 ;
        RECT 76.290 139.100 76.550 139.420 ;
        RECT 83.650 139.100 83.910 139.420 ;
        RECT 75.830 136.380 76.090 136.700 ;
        RECT 76.350 133.980 76.490 139.100 ;
        RECT 83.710 138.400 83.850 139.100 ;
        RECT 85.550 138.400 85.690 140.120 ;
        RECT 83.650 138.080 83.910 138.400 ;
        RECT 85.490 138.080 85.750 138.400 ;
        RECT 80.430 137.740 80.690 138.060 ;
        RECT 76.750 137.060 77.010 137.380 ;
        RECT 76.290 133.660 76.550 133.980 ;
        RECT 76.810 132.960 76.950 137.060 ;
        RECT 77.510 135.845 79.390 136.215 ;
        RECT 80.490 135.680 80.630 137.740 ;
        RECT 82.270 137.400 82.530 137.720 ;
        RECT 85.490 137.400 85.750 137.720 ;
        RECT 82.330 135.680 82.470 137.400 ;
        RECT 80.430 135.360 80.690 135.680 ;
        RECT 82.270 135.360 82.530 135.680 ;
        RECT 85.550 135.340 85.690 137.400 ;
        RECT 79.040 134.825 79.320 135.195 ;
        RECT 85.020 134.825 85.300 135.195 ;
        RECT 85.490 135.020 85.750 135.340 ;
        RECT 79.110 134.660 79.250 134.825 ;
        RECT 79.050 134.340 79.310 134.660 ;
        RECT 85.090 134.320 85.230 134.825 ;
        RECT 85.030 134.000 85.290 134.320 ;
        RECT 76.750 132.640 77.010 132.960 ;
        RECT 75.370 132.300 75.630 132.620 ;
        RECT 74.450 131.960 74.710 132.280 ;
        RECT 75.830 131.960 76.090 132.280 ;
        RECT 80.890 131.960 81.150 132.280 ;
        RECT 73.990 131.280 74.250 131.600 ;
        RECT 74.910 130.940 75.170 131.260 ;
        RECT 74.970 129.560 75.110 130.940 ;
        RECT 75.890 130.240 76.030 131.960 ;
        RECT 77.510 130.405 79.390 130.775 ;
        RECT 75.830 129.920 76.090 130.240 ;
        RECT 74.910 129.240 75.170 129.560 ;
        RECT 77.670 128.560 77.930 128.880 ;
        RECT 77.730 127.520 77.870 128.560 ;
        RECT 80.950 128.540 81.090 131.960 ;
        RECT 84.110 129.240 84.370 129.560 ;
        RECT 80.890 128.220 81.150 128.540 ;
        RECT 73.530 127.200 73.790 127.520 ;
        RECT 77.670 127.200 77.930 127.520 ;
        RECT 75.830 126.520 76.090 126.840 ;
        RECT 76.290 126.520 76.550 126.840 ;
        RECT 75.890 125.820 76.030 126.520 ;
        RECT 75.830 125.500 76.090 125.820 ;
        RECT 73.070 123.800 73.330 124.120 ;
        RECT 74.450 123.800 74.710 124.120 ;
        RECT 75.370 123.800 75.630 124.120 ;
        RECT 73.070 120.060 73.330 120.380 ;
        RECT 73.130 118.680 73.270 120.060 ;
        RECT 72.610 118.360 72.870 118.680 ;
        RECT 73.070 118.360 73.330 118.680 ;
        RECT 74.510 112.900 74.650 123.800 ;
        RECT 75.430 122.080 75.570 123.800 ;
        RECT 76.350 123.010 76.490 126.520 ;
        RECT 84.170 126.500 84.310 129.240 ;
        RECT 85.550 126.840 85.690 135.020 ;
        RECT 85.490 126.520 85.750 126.840 ;
        RECT 84.110 126.180 84.370 126.500 ;
        RECT 77.510 124.965 79.390 125.335 ;
        RECT 84.170 124.800 84.310 126.180 ;
        RECT 84.110 124.480 84.370 124.800 ;
        RECT 76.750 123.010 77.010 123.100 ;
        RECT 76.350 122.870 77.010 123.010 ;
        RECT 75.370 121.760 75.630 122.080 ;
        RECT 74.910 121.080 75.170 121.400 ;
        RECT 74.970 119.360 75.110 121.080 ;
        RECT 76.350 120.380 76.490 122.870 ;
        RECT 76.750 122.780 77.010 122.870 ;
        RECT 84.570 122.780 84.830 123.100 ;
        RECT 83.650 121.760 83.910 122.080 ;
        RECT 81.350 121.420 81.610 121.740 ;
        RECT 76.290 120.060 76.550 120.380 ;
        RECT 77.510 119.525 79.390 119.895 ;
        RECT 74.910 119.040 75.170 119.360 ;
        RECT 81.410 118.340 81.550 121.420 ;
        RECT 83.710 119.360 83.850 121.760 ;
        RECT 83.650 119.040 83.910 119.360 ;
        RECT 84.630 118.340 84.770 122.780 ;
        RECT 85.030 121.080 85.290 121.400 ;
        RECT 85.090 119.360 85.230 121.080 ;
        RECT 85.030 119.040 85.290 119.360 ;
        RECT 81.350 118.020 81.610 118.340 ;
        RECT 84.570 118.020 84.830 118.340 ;
        RECT 84.110 115.640 84.370 115.960 ;
        RECT 83.190 115.300 83.450 115.620 ;
        RECT 77.510 114.085 79.390 114.455 ;
        RECT 74.450 112.580 74.710 112.900 ;
        RECT 73.070 112.240 73.330 112.560 ;
        RECT 72.140 111.025 72.420 111.395 ;
        RECT 73.130 111.200 73.270 112.240 ;
        RECT 72.210 110.520 72.350 111.025 ;
        RECT 73.070 110.880 73.330 111.200 ;
        RECT 74.510 110.860 74.650 112.580 ;
        RECT 74.910 112.240 75.170 112.560 ;
        RECT 75.830 112.240 76.090 112.560 ;
        RECT 74.450 110.540 74.710 110.860 ;
        RECT 71.690 110.200 71.950 110.520 ;
        RECT 72.150 110.200 72.410 110.520 ;
        RECT 73.070 110.200 73.330 110.520 ;
        RECT 73.130 108.480 73.270 110.200 ;
        RECT 73.070 108.160 73.330 108.480 ;
        RECT 71.690 107.820 71.950 108.140 ;
        RECT 70.770 107.480 71.030 107.800 ;
        RECT 71.750 96.255 71.890 107.820 ;
        RECT 46.380 95.640 46.660 96.255 ;
        RECT 44.610 95.500 46.660 95.640 ;
        RECT 46.380 94.255 46.660 95.500 ;
        RECT 51.440 94.255 51.720 96.255 ;
        RECT 56.500 94.255 56.780 96.255 ;
        RECT 61.560 94.255 61.840 96.255 ;
        RECT 66.620 94.255 66.900 96.255 ;
        RECT 71.680 94.255 71.960 96.255 ;
        RECT 74.970 95.640 75.110 112.240 ;
        RECT 75.370 110.540 75.630 110.860 ;
        RECT 75.430 108.140 75.570 110.540 ;
        RECT 75.890 108.480 76.030 112.240 ;
        RECT 77.510 108.645 79.390 109.015 ;
        RECT 75.830 108.160 76.090 108.480 ;
        RECT 75.370 107.820 75.630 108.140 ;
        RECT 81.810 107.480 82.070 107.800 ;
        RECT 81.870 96.255 82.010 107.480 ;
        RECT 83.250 107.120 83.390 115.300 ;
        RECT 83.650 114.620 83.910 114.940 ;
        RECT 83.710 113.240 83.850 114.620 ;
        RECT 83.650 112.920 83.910 113.240 ;
        RECT 84.170 107.120 84.310 115.640 ;
        RECT 85.490 112.920 85.750 113.240 ;
        RECT 85.030 111.900 85.290 112.220 ;
        RECT 85.090 107.800 85.230 111.900 ;
        RECT 85.550 110.180 85.690 112.920 ;
        RECT 86.010 112.900 86.150 140.800 ;
        RECT 87.390 137.720 87.530 141.820 ;
        RECT 87.330 137.400 87.590 137.720 ;
        RECT 87.330 132.300 87.590 132.620 ;
        RECT 86.870 131.620 87.130 131.940 ;
        RECT 86.930 123.780 87.070 131.620 ;
        RECT 87.390 127.520 87.530 132.300 ;
        RECT 87.330 127.200 87.590 127.520 ;
        RECT 86.870 123.460 87.130 123.780 ;
        RECT 86.930 121.060 87.070 123.460 ;
        RECT 86.870 120.740 87.130 121.060 ;
        RECT 86.930 113.240 87.070 120.740 ;
        RECT 87.850 115.960 87.990 144.540 ;
        RECT 88.310 137.720 88.450 145.140 ;
        RECT 89.170 143.520 89.430 143.840 ;
        RECT 89.230 143.160 89.370 143.520 ;
        RECT 89.170 142.840 89.430 143.160 ;
        RECT 89.230 141.120 89.370 142.840 ;
        RECT 89.170 140.800 89.430 141.120 ;
        RECT 88.250 137.400 88.510 137.720 ;
        RECT 88.710 130.940 88.970 131.260 ;
        RECT 88.770 129.900 88.910 130.940 ;
        RECT 89.690 130.240 89.830 146.240 ;
        RECT 90.150 145.880 90.290 177.180 ;
        RECT 91.530 176.480 91.670 179.900 ;
        RECT 94.680 179.025 94.960 179.395 ;
        RECT 91.920 178.345 92.200 178.715 ;
        RECT 94.750 178.520 94.890 179.025 ;
        RECT 91.990 178.180 92.130 178.345 ;
        RECT 94.690 178.200 94.950 178.520 ;
        RECT 91.930 177.860 92.190 178.180 ;
        RECT 91.930 177.180 92.190 177.500 ;
        RECT 91.470 176.160 91.730 176.480 ;
        RECT 91.990 170.950 92.130 177.180 ;
        RECT 92.510 176.645 94.390 177.015 ;
        RECT 94.750 176.140 94.890 178.200 ;
        RECT 95.150 178.035 95.410 178.180 ;
        RECT 95.140 177.665 95.420 178.035 ;
        RECT 94.690 176.050 94.950 176.140 ;
        RECT 94.290 175.910 94.950 176.050 ;
        RECT 93.310 175.480 93.570 175.800 ;
        RECT 93.370 172.740 93.510 175.480 ;
        RECT 94.290 173.080 94.430 175.910 ;
        RECT 94.690 175.820 94.950 175.910 ;
        RECT 95.210 175.800 95.350 177.665 ;
        RECT 95.150 175.480 95.410 175.800 ;
        RECT 95.150 174.460 95.410 174.780 ;
        RECT 94.230 172.760 94.490 173.080 ;
        RECT 94.690 172.760 94.950 173.080 ;
        RECT 93.310 172.420 93.570 172.740 ;
        RECT 92.510 171.205 94.390 171.575 ;
        RECT 94.750 171.040 94.890 172.760 ;
        RECT 91.990 170.810 92.590 170.950 ;
        RECT 91.930 167.320 92.190 167.640 ;
        RECT 91.010 166.980 91.270 167.300 ;
        RECT 90.550 163.580 90.810 163.900 ;
        RECT 90.610 162.200 90.750 163.580 ;
        RECT 91.070 162.880 91.210 166.980 ;
        RECT 91.470 166.640 91.730 166.960 ;
        RECT 91.530 165.260 91.670 166.640 ;
        RECT 91.470 164.940 91.730 165.260 ;
        RECT 91.990 164.490 92.130 167.320 ;
        RECT 92.450 166.795 92.590 170.810 ;
        RECT 94.690 170.720 94.950 171.040 ;
        RECT 94.690 169.020 94.950 169.340 ;
        RECT 94.750 166.960 94.890 169.020 ;
        RECT 92.380 166.425 92.660 166.795 ;
        RECT 94.690 166.640 94.950 166.960 ;
        RECT 92.510 165.765 94.390 166.135 ;
        RECT 91.460 164.065 91.740 164.435 ;
        RECT 91.990 164.350 92.590 164.490 ;
        RECT 91.010 162.560 91.270 162.880 ;
        RECT 90.550 161.880 90.810 162.200 ;
        RECT 90.550 158.820 90.810 159.140 ;
        RECT 90.610 150.980 90.750 158.820 ;
        RECT 91.010 152.700 91.270 153.020 ;
        RECT 91.070 152.000 91.210 152.700 ;
        RECT 91.010 151.680 91.270 152.000 ;
        RECT 91.530 151.400 91.670 164.065 ;
        RECT 92.450 161.600 92.590 164.350 ;
        RECT 91.990 161.520 92.590 161.600 ;
        RECT 91.930 161.460 92.590 161.520 ;
        RECT 91.930 161.200 92.190 161.460 ;
        RECT 91.990 159.480 92.130 161.200 ;
        RECT 94.690 160.860 94.950 161.180 ;
        RECT 92.510 160.325 94.390 160.695 ;
        RECT 94.750 160.160 94.890 160.860 ;
        RECT 94.690 159.840 94.950 160.160 ;
        RECT 91.930 159.160 92.190 159.480 ;
        RECT 94.690 159.160 94.950 159.480 ;
        RECT 91.990 157.100 92.130 159.160 ;
        RECT 91.930 156.780 92.190 157.100 ;
        RECT 94.750 156.760 94.890 159.160 ;
        RECT 92.450 156.530 93.970 156.670 ;
        RECT 91.930 156.275 92.190 156.420 ;
        RECT 91.920 155.905 92.200 156.275 ;
        RECT 92.450 155.650 92.590 156.530 ;
        RECT 93.300 155.905 93.580 156.275 ;
        RECT 93.830 156.080 93.970 156.530 ;
        RECT 94.690 156.440 94.950 156.760 ;
        RECT 93.370 155.740 93.510 155.905 ;
        RECT 93.770 155.760 94.030 156.080 ;
        RECT 91.990 155.510 92.590 155.650 ;
        RECT 91.990 154.630 92.130 155.510 ;
        RECT 93.310 155.420 93.570 155.740 ;
        RECT 92.510 154.885 94.390 155.255 ;
        RECT 91.990 154.490 93.050 154.630 ;
        RECT 92.390 153.040 92.650 153.360 ;
        RECT 91.530 151.260 92.130 151.400 ;
        RECT 90.550 150.660 90.810 150.980 ;
        RECT 91.470 150.660 91.730 150.980 ;
        RECT 90.550 149.980 90.810 150.300 ;
        RECT 90.090 145.560 90.350 145.880 ;
        RECT 90.090 144.880 90.350 145.200 ;
        RECT 90.150 143.840 90.290 144.880 ;
        RECT 90.090 143.520 90.350 143.840 ;
        RECT 90.610 143.240 90.750 149.980 ;
        RECT 91.530 148.600 91.670 150.660 ;
        RECT 91.470 148.280 91.730 148.600 ;
        RECT 91.470 145.900 91.730 146.220 ;
        RECT 90.150 143.100 90.750 143.240 ;
        RECT 89.630 129.920 89.890 130.240 ;
        RECT 88.710 129.580 88.970 129.900 ;
        RECT 88.250 128.900 88.510 129.220 ;
        RECT 88.310 126.840 88.450 128.900 ;
        RECT 88.770 128.880 88.910 129.580 ;
        RECT 88.710 128.560 88.970 128.880 ;
        RECT 88.250 126.520 88.510 126.840 ;
        RECT 88.310 124.120 88.450 126.520 ;
        RECT 88.250 123.800 88.510 124.120 ;
        RECT 88.310 122.080 88.450 123.800 ;
        RECT 88.250 121.760 88.510 122.080 ;
        RECT 90.150 118.000 90.290 143.100 ;
        RECT 90.550 142.675 90.810 142.820 ;
        RECT 90.540 142.305 90.820 142.675 ;
        RECT 91.530 142.140 91.670 145.900 ;
        RECT 91.470 141.820 91.730 142.140 ;
        RECT 91.010 140.120 91.270 140.440 ;
        RECT 90.550 139.440 90.810 139.760 ;
        RECT 90.610 138.400 90.750 139.440 ;
        RECT 90.550 138.080 90.810 138.400 ;
        RECT 91.070 135.680 91.210 140.120 ;
        RECT 91.990 137.380 92.130 151.260 ;
        RECT 92.450 150.980 92.590 153.040 ;
        RECT 92.910 150.980 93.050 154.490 ;
        RECT 94.750 154.040 94.890 156.440 ;
        RECT 94.690 153.720 94.950 154.040 ;
        RECT 93.830 152.620 94.890 152.760 ;
        RECT 92.390 150.660 92.650 150.980 ;
        RECT 92.850 150.660 93.110 150.980 ;
        RECT 93.830 150.210 93.970 152.620 ;
        RECT 94.750 152.000 94.890 152.620 ;
        RECT 94.230 151.680 94.490 152.000 ;
        RECT 94.690 151.680 94.950 152.000 ;
        RECT 94.290 150.720 94.430 151.680 ;
        RECT 95.210 151.320 95.350 174.460 ;
        RECT 95.670 173.080 95.810 194.520 ;
        RECT 97.510 191.780 97.650 196.220 ;
        RECT 107.510 195.685 109.390 196.055 ;
        RECT 100.670 194.520 100.930 194.840 ;
        RECT 96.530 191.460 96.790 191.780 ;
        RECT 97.450 191.460 97.710 191.780 ;
        RECT 96.590 189.740 96.730 191.460 ;
        RECT 96.530 189.420 96.790 189.740 ;
        RECT 96.070 188.740 96.330 189.060 ;
        RECT 96.130 182.940 96.270 188.740 ;
        RECT 96.590 187.360 96.730 189.420 ;
        RECT 97.510 188.380 97.650 191.460 ;
        RECT 99.750 190.780 100.010 191.100 ;
        RECT 99.810 189.060 99.950 190.780 ;
        RECT 99.750 188.740 100.010 189.060 ;
        RECT 97.450 188.060 97.710 188.380 ;
        RECT 100.730 187.360 100.870 194.520 ;
        RECT 104.810 194.180 105.070 194.500 ;
        RECT 102.510 193.840 102.770 194.160 ;
        RECT 102.570 190.080 102.710 193.840 ;
        RECT 102.510 189.760 102.770 190.080 ;
        RECT 103.430 188.400 103.690 188.720 ;
        RECT 96.530 187.040 96.790 187.360 ;
        RECT 100.670 187.040 100.930 187.360 ;
        RECT 96.590 186.340 96.730 187.040 ;
        RECT 100.730 186.680 100.870 187.040 ;
        RECT 97.450 186.360 97.710 186.680 ;
        RECT 100.670 186.360 100.930 186.680 ;
        RECT 96.530 186.020 96.790 186.340 ;
        RECT 96.590 184.040 96.730 186.020 ;
        RECT 96.590 183.900 97.190 184.040 ;
        RECT 96.530 182.960 96.790 183.280 ;
        RECT 96.070 182.620 96.330 182.940 ;
        RECT 96.130 178.180 96.270 182.620 ;
        RECT 96.590 181.920 96.730 182.960 ;
        RECT 96.530 181.600 96.790 181.920 ;
        RECT 97.050 180.900 97.190 183.900 ;
        RECT 97.510 181.920 97.650 186.360 ;
        RECT 101.130 185.340 101.390 185.660 ;
        RECT 102.050 185.340 102.310 185.660 ;
        RECT 98.370 183.640 98.630 183.960 ;
        RECT 97.450 181.600 97.710 181.920 ;
        RECT 98.430 181.580 98.570 183.640 ;
        RECT 101.190 183.620 101.330 185.340 ;
        RECT 101.130 183.300 101.390 183.620 ;
        RECT 98.370 181.260 98.630 181.580 ;
        RECT 102.110 180.900 102.250 185.340 ;
        RECT 103.490 181.920 103.630 188.400 ;
        RECT 104.870 183.960 105.010 194.180 ;
        RECT 105.730 192.140 105.990 192.460 ;
        RECT 105.270 190.780 105.530 191.100 ;
        RECT 105.330 189.060 105.470 190.780 ;
        RECT 105.790 190.080 105.930 192.140 ;
        RECT 111.250 191.460 111.510 191.780 ;
        RECT 107.110 190.780 107.370 191.100 ;
        RECT 105.730 189.760 105.990 190.080 ;
        RECT 107.170 189.740 107.310 190.780 ;
        RECT 107.510 190.245 109.390 190.615 ;
        RECT 107.110 189.420 107.370 189.740 ;
        RECT 105.270 188.740 105.530 189.060 ;
        RECT 108.030 188.740 108.290 189.060 ;
        RECT 104.810 183.640 105.070 183.960 ;
        RECT 104.870 182.940 105.010 183.640 ;
        RECT 104.810 182.620 105.070 182.940 ;
        RECT 103.430 181.600 103.690 181.920 ;
        RECT 96.990 180.580 97.250 180.900 ;
        RECT 102.050 180.580 102.310 180.900 ;
        RECT 96.980 178.345 97.260 178.715 ;
        RECT 97.050 178.180 97.190 178.345 ;
        RECT 96.070 177.860 96.330 178.180 ;
        RECT 96.990 177.860 97.250 178.180 ;
        RECT 96.530 175.820 96.790 176.140 ;
        RECT 95.610 172.760 95.870 173.080 ;
        RECT 96.590 172.650 96.730 175.820 ;
        RECT 97.050 175.800 97.190 177.860 ;
        RECT 97.450 177.520 97.710 177.840 ;
        RECT 96.990 175.480 97.250 175.800 ;
        RECT 97.050 173.760 97.190 175.480 ;
        RECT 96.990 173.440 97.250 173.760 ;
        RECT 96.990 172.650 97.250 172.740 ;
        RECT 96.590 172.510 97.250 172.650 ;
        RECT 96.990 172.420 97.250 172.510 ;
        RECT 96.070 172.080 96.330 172.400 ;
        RECT 96.130 163.640 96.270 172.080 ;
        RECT 97.510 170.440 97.650 177.520 ;
        RECT 98.830 177.180 99.090 177.500 ;
        RECT 99.290 177.180 99.550 177.500 ;
        RECT 98.370 173.440 98.630 173.760 ;
        RECT 98.430 172.740 98.570 173.440 ;
        RECT 98.890 172.740 99.030 177.180 ;
        RECT 98.370 172.420 98.630 172.740 ;
        RECT 98.830 172.420 99.090 172.740 ;
        RECT 97.910 171.740 98.170 172.060 ;
        RECT 97.970 171.040 98.110 171.740 ;
        RECT 97.910 170.720 98.170 171.040 ;
        RECT 97.510 170.300 98.110 170.440 ;
        RECT 98.890 170.360 99.030 172.420 ;
        RECT 99.350 170.700 99.490 177.180 ;
        RECT 99.750 175.820 100.010 176.140 ;
        RECT 99.810 173.760 99.950 175.820 ;
        RECT 99.750 173.440 100.010 173.760 ;
        RECT 102.110 173.420 102.250 180.580 ;
        RECT 105.330 178.180 105.470 188.740 ;
        RECT 108.090 187.360 108.230 188.740 ;
        RECT 108.030 187.040 108.290 187.360 ;
        RECT 110.330 187.040 110.590 187.360 ;
        RECT 106.650 186.700 106.910 187.020 ;
        RECT 109.870 186.700 110.130 187.020 ;
        RECT 106.710 184.640 106.850 186.700 ;
        RECT 107.510 184.805 109.390 185.175 ;
        RECT 106.650 184.320 106.910 184.640 ;
        RECT 106.650 182.960 106.910 183.280 ;
        RECT 105.730 179.900 105.990 180.220 ;
        RECT 105.790 178.520 105.930 179.900 ;
        RECT 106.710 179.200 106.850 182.960 ;
        RECT 107.110 179.900 107.370 180.220 ;
        RECT 106.650 178.880 106.910 179.200 ;
        RECT 107.170 178.520 107.310 179.900 ;
        RECT 107.510 179.365 109.390 179.735 ;
        RECT 109.930 179.200 110.070 186.700 ;
        RECT 110.390 183.620 110.530 187.040 ;
        RECT 110.790 186.020 111.050 186.340 ;
        RECT 110.850 183.960 110.990 186.020 ;
        RECT 110.790 183.640 111.050 183.960 ;
        RECT 110.330 183.300 110.590 183.620 ;
        RECT 109.870 178.880 110.130 179.200 ;
        RECT 105.730 178.200 105.990 178.520 ;
        RECT 107.110 178.200 107.370 178.520 ;
        RECT 103.430 177.860 103.690 178.180 ;
        RECT 104.350 178.035 104.610 178.180 ;
        RECT 103.490 174.780 103.630 177.860 ;
        RECT 104.340 177.665 104.620 178.035 ;
        RECT 105.270 177.860 105.530 178.180 ;
        RECT 111.310 175.460 111.450 191.460 ;
        RECT 106.650 175.140 106.910 175.460 ;
        RECT 111.250 175.370 111.510 175.460 ;
        RECT 110.850 175.230 111.510 175.370 ;
        RECT 103.430 174.460 103.690 174.780 ;
        RECT 102.050 173.100 102.310 173.420 ;
        RECT 100.670 172.420 100.930 172.740 ;
        RECT 99.290 170.380 99.550 170.700 ;
        RECT 96.990 169.700 97.250 170.020 ;
        RECT 97.050 169.340 97.190 169.700 ;
        RECT 96.990 169.020 97.250 169.340 ;
        RECT 96.530 166.300 96.790 166.620 ;
        RECT 96.590 164.920 96.730 166.300 ;
        RECT 96.530 164.600 96.790 164.920 ;
        RECT 96.130 163.500 96.730 163.640 ;
        RECT 95.610 158.140 95.870 158.460 ;
        RECT 95.150 151.000 95.410 151.320 ;
        RECT 94.290 150.580 95.350 150.720 ;
        RECT 93.830 150.070 94.890 150.210 ;
        RECT 92.510 149.445 94.390 149.815 ;
        RECT 92.510 144.005 94.390 144.375 ;
        RECT 93.770 143.180 94.030 143.500 ;
        RECT 94.230 143.180 94.490 143.500 ;
        RECT 93.830 142.820 93.970 143.180 ;
        RECT 92.390 142.500 92.650 142.820 ;
        RECT 93.770 142.500 94.030 142.820 ;
        RECT 92.450 142.140 92.590 142.500 ;
        RECT 94.290 142.480 94.430 143.180 ;
        RECT 94.230 142.160 94.490 142.480 ;
        RECT 92.390 141.820 92.650 142.140 ;
        RECT 92.510 138.565 94.390 138.935 ;
        RECT 93.760 137.545 94.040 137.915 ;
        RECT 93.770 137.400 94.030 137.545 ;
        RECT 91.930 137.060 92.190 137.380 ;
        RECT 91.010 135.360 91.270 135.680 ;
        RECT 92.510 133.125 94.390 133.495 ;
        RECT 94.750 132.960 94.890 150.070 ;
        RECT 95.210 146.560 95.350 150.580 ;
        RECT 95.670 148.940 95.810 158.140 ;
        RECT 96.070 157.120 96.330 157.440 ;
        RECT 96.130 156.420 96.270 157.120 ;
        RECT 96.070 156.100 96.330 156.420 ;
        RECT 96.070 152.700 96.330 153.020 ;
        RECT 95.610 148.620 95.870 148.940 ;
        RECT 95.150 146.240 95.410 146.560 ;
        RECT 95.610 144.540 95.870 144.860 ;
        RECT 95.150 141.820 95.410 142.140 ;
        RECT 95.210 138.060 95.350 141.820 ;
        RECT 95.670 138.060 95.810 144.540 ;
        RECT 96.130 138.060 96.270 152.700 ;
        RECT 95.150 137.740 95.410 138.060 ;
        RECT 95.610 137.740 95.870 138.060 ;
        RECT 96.070 137.740 96.330 138.060 ;
        RECT 96.590 137.720 96.730 163.500 ;
        RECT 97.050 162.200 97.190 169.020 ;
        RECT 96.990 161.880 97.250 162.200 ;
        RECT 96.980 156.585 97.260 156.955 ;
        RECT 97.050 156.420 97.190 156.585 ;
        RECT 96.990 156.100 97.250 156.420 ;
        RECT 97.450 153.040 97.710 153.360 ;
        RECT 97.510 150.980 97.650 153.040 ;
        RECT 96.990 150.835 97.250 150.980 ;
        RECT 96.980 150.465 97.260 150.835 ;
        RECT 97.450 150.660 97.710 150.980 ;
        RECT 97.970 150.040 98.110 170.300 ;
        RECT 98.830 170.040 99.090 170.360 ;
        RECT 99.290 167.320 99.550 167.640 ;
        RECT 99.350 159.480 99.490 167.320 ;
        RECT 99.750 166.640 100.010 166.960 ;
        RECT 99.810 165.600 99.950 166.640 ;
        RECT 99.750 165.280 100.010 165.600 ;
        RECT 100.730 164.920 100.870 172.420 ;
        RECT 102.050 171.740 102.310 172.060 ;
        RECT 102.110 167.640 102.250 171.740 ;
        RECT 102.970 169.700 103.230 170.020 ;
        RECT 102.050 167.320 102.310 167.640 ;
        RECT 101.130 166.980 101.390 167.300 ;
        RECT 100.670 164.600 100.930 164.920 ;
        RECT 101.190 164.580 101.330 166.980 ;
        RECT 103.030 166.620 103.170 169.700 ;
        RECT 102.970 166.300 103.230 166.620 ;
        RECT 101.130 164.260 101.390 164.580 ;
        RECT 102.050 163.580 102.310 163.900 ;
        RECT 98.370 159.390 98.630 159.480 ;
        RECT 98.370 159.250 99.030 159.390 ;
        RECT 98.370 159.160 98.630 159.250 ;
        RECT 98.370 158.480 98.630 158.800 ;
        RECT 98.430 154.040 98.570 158.480 ;
        RECT 98.890 158.460 99.030 159.250 ;
        RECT 99.290 159.160 99.550 159.480 ;
        RECT 99.750 159.160 100.010 159.480 ;
        RECT 98.830 158.140 99.090 158.460 ;
        RECT 98.890 157.100 99.030 158.140 ;
        RECT 98.830 156.780 99.090 157.100 ;
        RECT 98.370 153.720 98.630 154.040 ;
        RECT 98.890 153.700 99.030 156.780 ;
        RECT 99.290 156.330 99.550 156.420 ;
        RECT 99.810 156.330 99.950 159.160 ;
        RECT 102.110 158.800 102.250 163.580 ;
        RECT 103.030 161.860 103.170 166.300 ;
        RECT 102.970 161.540 103.230 161.860 ;
        RECT 102.510 160.860 102.770 161.180 ;
        RECT 102.570 160.160 102.710 160.860 ;
        RECT 102.510 159.840 102.770 160.160 ;
        RECT 103.490 159.480 103.630 174.460 ;
        RECT 106.710 171.040 106.850 175.140 ;
        RECT 107.510 173.925 109.390 174.295 ;
        RECT 110.850 172.740 110.990 175.230 ;
        RECT 111.250 175.140 111.510 175.230 ;
        RECT 135.630 173.380 136.780 174.600 ;
        RECT 110.790 172.420 111.050 172.740 ;
        RECT 109.410 172.080 109.670 172.400 ;
        RECT 109.470 171.040 109.610 172.080 ;
        RECT 106.650 170.720 106.910 171.040 ;
        RECT 109.410 170.720 109.670 171.040 ;
        RECT 107.510 168.485 109.390 168.855 ;
        RECT 107.110 168.000 107.370 168.320 ;
        RECT 104.810 166.980 105.070 167.300 ;
        RECT 104.350 164.260 104.610 164.580 ;
        RECT 103.890 163.920 104.150 164.240 ;
        RECT 103.950 162.540 104.090 163.920 ;
        RECT 103.890 162.220 104.150 162.540 ;
        RECT 102.510 159.160 102.770 159.480 ;
        RECT 103.430 159.160 103.690 159.480 ;
        RECT 102.050 158.480 102.310 158.800 ;
        RECT 102.570 158.460 102.710 159.160 ;
        RECT 102.510 158.140 102.770 158.460 ;
        RECT 104.410 157.440 104.550 164.260 ;
        RECT 104.870 162.880 105.010 166.980 ;
        RECT 104.810 162.560 105.070 162.880 ;
        RECT 107.170 162.200 107.310 168.000 ;
        RECT 109.410 166.300 109.670 166.620 ;
        RECT 109.470 165.260 109.610 166.300 ;
        RECT 109.410 164.940 109.670 165.260 ;
        RECT 110.850 164.580 110.990 172.420 ;
        RECT 133.750 170.070 134.880 172.730 ;
        RECT 113.540 169.505 113.820 169.875 ;
        RECT 113.610 167.300 113.750 169.505 ;
        RECT 113.550 166.980 113.810 167.300 ;
        RECT 135.630 166.640 136.740 173.380 ;
        RECT 135.630 165.420 136.780 166.640 ;
        RECT 110.790 164.260 111.050 164.580 ;
        RECT 107.510 163.045 109.390 163.415 ;
        RECT 107.110 161.880 107.370 162.200 ;
        RECT 110.790 161.880 111.050 162.200 ;
        RECT 110.330 161.540 110.590 161.860 ;
        RECT 110.390 159.480 110.530 161.540 ;
        RECT 110.850 159.480 110.990 161.880 ;
        RECT 104.810 159.160 105.070 159.480 ;
        RECT 110.330 159.160 110.590 159.480 ;
        RECT 110.790 159.160 111.050 159.480 ;
        RECT 104.350 157.120 104.610 157.440 ;
        RECT 99.290 156.190 99.950 156.330 ;
        RECT 99.290 156.100 99.550 156.190 ;
        RECT 99.350 154.040 99.490 156.100 ;
        RECT 103.890 155.760 104.150 156.080 ;
        RECT 101.130 155.420 101.390 155.740 ;
        RECT 99.290 153.720 99.550 154.040 ;
        RECT 98.830 153.380 99.090 153.700 ;
        RECT 101.190 150.980 101.330 155.420 ;
        RECT 103.950 153.700 104.090 155.760 ;
        RECT 104.870 154.720 105.010 159.160 ;
        RECT 109.870 158.140 110.130 158.460 ;
        RECT 107.510 157.605 109.390 157.975 ;
        RECT 109.930 156.080 110.070 158.140 ;
        RECT 109.870 155.760 110.130 156.080 ;
        RECT 110.330 155.760 110.590 156.080 ;
        RECT 110.390 154.720 110.530 155.760 ;
        RECT 104.810 154.400 105.070 154.720 ;
        RECT 110.330 154.400 110.590 154.720 ;
        RECT 103.890 153.380 104.150 153.700 ;
        RECT 103.950 150.980 104.090 153.380 ;
        RECT 104.350 153.040 104.610 153.360 ;
        RECT 104.410 151.320 104.550 153.040 ;
        RECT 107.510 152.165 109.390 152.535 ;
        RECT 105.730 151.340 105.990 151.660 ;
        RECT 104.350 151.000 104.610 151.320 ;
        RECT 98.360 150.465 98.640 150.835 ;
        RECT 99.750 150.660 100.010 150.980 ;
        RECT 100.210 150.660 100.470 150.980 ;
        RECT 101.130 150.660 101.390 150.980 ;
        RECT 103.890 150.660 104.150 150.980 ;
        RECT 97.510 149.900 98.110 150.040 ;
        RECT 96.990 148.280 97.250 148.600 ;
        RECT 97.050 147.490 97.190 148.280 ;
        RECT 97.510 148.260 97.650 149.900 ;
        RECT 98.430 148.600 98.570 150.465 ;
        RECT 99.810 150.300 99.950 150.660 ;
        RECT 99.750 149.980 100.010 150.300 ;
        RECT 99.290 148.960 99.550 149.280 ;
        RECT 98.370 148.280 98.630 148.600 ;
        RECT 98.830 148.280 99.090 148.600 ;
        RECT 97.450 147.940 97.710 148.260 ;
        RECT 97.050 147.350 97.650 147.490 ;
        RECT 96.990 146.240 97.250 146.560 ;
        RECT 96.530 137.400 96.790 137.720 ;
        RECT 95.610 136.720 95.870 137.040 ;
        RECT 95.150 136.380 95.410 136.700 ;
        RECT 94.690 132.640 94.950 132.960 ;
        RECT 91.010 131.960 91.270 132.280 ;
        RECT 91.070 130.240 91.210 131.960 ;
        RECT 95.210 130.240 95.350 136.380 ;
        RECT 91.010 129.920 91.270 130.240 ;
        RECT 95.150 129.920 95.410 130.240 ;
        RECT 91.010 129.130 91.270 129.220 ;
        RECT 90.610 128.990 91.270 129.130 ;
        RECT 90.610 126.500 90.750 128.990 ;
        RECT 91.010 128.900 91.270 128.990 ;
        RECT 92.510 127.685 94.390 128.055 ;
        RECT 90.550 126.180 90.810 126.500 ;
        RECT 90.610 124.800 90.750 126.180 ;
        RECT 91.470 125.500 91.730 125.820 ;
        RECT 93.770 125.500 94.030 125.820 ;
        RECT 90.550 124.480 90.810 124.800 ;
        RECT 91.530 118.340 91.670 125.500 ;
        RECT 93.830 123.440 93.970 125.500 ;
        RECT 93.770 123.120 94.030 123.440 ;
        RECT 92.510 122.245 94.390 122.615 ;
        RECT 91.930 120.740 92.190 121.060 ;
        RECT 91.990 119.360 92.130 120.740 ;
        RECT 91.930 119.040 92.190 119.360 ;
        RECT 91.470 118.020 91.730 118.340 ;
        RECT 90.090 117.680 90.350 118.000 ;
        RECT 92.510 116.805 94.390 117.175 ;
        RECT 95.670 115.960 95.810 136.720 ;
        RECT 96.530 136.380 96.790 136.700 ;
        RECT 96.590 130.240 96.730 136.380 ;
        RECT 97.050 132.960 97.190 146.240 ;
        RECT 97.510 145.540 97.650 147.350 ;
        RECT 97.910 147.260 98.170 147.580 ;
        RECT 97.450 145.220 97.710 145.540 ;
        RECT 97.510 143.160 97.650 145.220 ;
        RECT 97.450 142.840 97.710 143.160 ;
        RECT 97.450 136.380 97.710 136.700 ;
        RECT 96.990 132.640 97.250 132.960 ;
        RECT 96.990 131.620 97.250 131.940 ;
        RECT 96.530 129.920 96.790 130.240 ;
        RECT 97.050 129.900 97.190 131.620 ;
        RECT 96.990 129.580 97.250 129.900 ;
        RECT 87.790 115.640 88.050 115.960 ;
        RECT 95.610 115.640 95.870 115.960 ;
        RECT 90.550 114.620 90.810 114.940 ;
        RECT 95.610 114.620 95.870 114.940 ;
        RECT 86.870 112.920 87.130 113.240 ;
        RECT 85.950 112.580 86.210 112.900 ;
        RECT 90.610 111.200 90.750 114.620 ;
        RECT 95.670 113.240 95.810 114.620 ;
        RECT 91.470 112.920 91.730 113.240 ;
        RECT 95.610 112.920 95.870 113.240 ;
        RECT 90.550 110.880 90.810 111.200 ;
        RECT 86.410 110.540 86.670 110.860 ;
        RECT 85.490 109.860 85.750 110.180 ;
        RECT 85.030 107.480 85.290 107.800 ;
        RECT 83.190 106.800 83.450 107.120 ;
        RECT 84.110 106.800 84.370 107.120 ;
        RECT 86.470 104.580 86.610 110.540 ;
        RECT 88.710 110.200 88.970 110.520 ;
        RECT 86.870 109.860 87.130 110.180 ;
        RECT 86.930 107.800 87.070 109.860 ;
        RECT 88.770 108.480 88.910 110.200 ;
        RECT 88.710 108.160 88.970 108.480 ;
        RECT 86.870 107.480 87.130 107.800 ;
        RECT 86.470 104.440 87.070 104.580 ;
        RECT 86.930 96.255 87.070 104.440 ;
        RECT 76.740 95.640 77.020 96.255 ;
        RECT 74.970 95.500 77.020 95.640 ;
        RECT 76.740 94.255 77.020 95.500 ;
        RECT 81.800 94.255 82.080 96.255 ;
        RECT 86.860 94.255 87.140 96.255 ;
        RECT 91.530 95.640 91.670 112.920 ;
        RECT 97.510 112.560 97.650 136.380 ;
        RECT 97.970 135.680 98.110 147.260 ;
        RECT 98.430 145.880 98.570 148.280 ;
        RECT 98.890 147.580 99.030 148.280 ;
        RECT 98.830 147.260 99.090 147.580 ;
        RECT 98.370 145.560 98.630 145.880 ;
        RECT 98.430 143.840 98.570 145.560 ;
        RECT 98.370 143.520 98.630 143.840 ;
        RECT 98.830 142.840 99.090 143.160 ;
        RECT 98.370 142.160 98.630 142.480 ;
        RECT 98.430 140.100 98.570 142.160 ;
        RECT 98.370 139.780 98.630 140.100 ;
        RECT 98.890 139.420 99.030 142.840 ;
        RECT 98.830 139.100 99.090 139.420 ;
        RECT 97.910 135.360 98.170 135.680 ;
        RECT 98.830 134.340 99.090 134.660 ;
        RECT 98.890 132.280 99.030 134.340 ;
        RECT 98.830 131.960 99.090 132.280 ;
        RECT 98.890 129.560 99.030 131.960 ;
        RECT 98.830 129.240 99.090 129.560 ;
        RECT 98.370 128.900 98.630 129.220 ;
        RECT 98.430 126.500 98.570 128.900 ;
        RECT 98.370 126.180 98.630 126.500 ;
        RECT 98.370 125.500 98.630 125.820 ;
        RECT 97.910 123.460 98.170 123.780 ;
        RECT 97.970 122.080 98.110 123.460 ;
        RECT 97.910 121.760 98.170 122.080 ;
        RECT 98.430 121.400 98.570 125.500 ;
        RECT 98.370 121.080 98.630 121.400 ;
        RECT 99.350 115.960 99.490 148.960 ;
        RECT 99.810 148.600 99.950 149.980 ;
        RECT 100.270 148.940 100.410 150.660 ;
        RECT 100.210 148.620 100.470 148.940 ;
        RECT 99.750 148.280 100.010 148.600 ;
        RECT 99.810 145.450 99.950 148.280 ;
        RECT 101.130 147.600 101.390 147.920 ;
        RECT 101.190 146.220 101.330 147.600 ;
        RECT 101.130 145.900 101.390 146.220 ;
        RECT 100.210 145.450 100.470 145.540 ;
        RECT 99.810 145.310 100.470 145.450 ;
        RECT 99.810 143.355 99.950 145.310 ;
        RECT 100.210 145.220 100.470 145.310 ;
        RECT 99.740 142.985 100.020 143.355 ;
        RECT 101.190 143.160 101.330 145.900 ;
        RECT 104.410 145.880 104.550 151.000 ;
        RECT 104.810 149.980 105.070 150.300 ;
        RECT 104.870 147.580 105.010 149.980 ;
        RECT 104.810 147.260 105.070 147.580 ;
        RECT 104.350 145.560 104.610 145.880 ;
        RECT 102.510 144.540 102.770 144.860 ;
        RECT 102.570 143.500 102.710 144.540 ;
        RECT 102.510 143.180 102.770 143.500 ;
        RECT 99.750 142.840 100.010 142.985 ;
        RECT 101.130 142.840 101.390 143.160 ;
        RECT 101.590 141.820 101.850 142.140 ;
        RECT 101.650 139.760 101.790 141.820 ;
        RECT 101.590 139.440 101.850 139.760 ;
        RECT 102.050 139.100 102.310 139.420 ;
        RECT 102.110 138.400 102.250 139.100 ;
        RECT 102.570 138.400 102.710 143.180 ;
        RECT 102.050 138.080 102.310 138.400 ;
        RECT 102.510 138.080 102.770 138.400 ;
        RECT 104.410 137.380 104.550 145.560 ;
        RECT 104.870 145.540 105.010 147.260 ;
        RECT 104.810 145.220 105.070 145.540 ;
        RECT 104.350 137.060 104.610 137.380 ;
        RECT 104.810 134.340 105.070 134.660 ;
        RECT 100.670 131.960 100.930 132.280 ;
        RECT 99.750 131.620 100.010 131.940 ;
        RECT 99.810 129.220 99.950 131.620 ;
        RECT 100.210 129.920 100.470 130.240 ;
        RECT 100.270 129.560 100.410 129.920 ;
        RECT 100.210 129.240 100.470 129.560 ;
        RECT 99.750 128.900 100.010 129.220 ;
        RECT 99.750 126.180 100.010 126.500 ;
        RECT 99.810 124.460 99.950 126.180 ;
        RECT 100.270 126.160 100.410 129.240 ;
        RECT 100.730 126.840 100.870 131.960 ;
        RECT 104.870 128.540 105.010 134.340 ;
        RECT 104.810 128.220 105.070 128.540 ;
        RECT 104.870 127.520 105.010 128.220 ;
        RECT 102.050 127.200 102.310 127.520 ;
        RECT 104.810 127.200 105.070 127.520 ;
        RECT 100.670 126.520 100.930 126.840 ;
        RECT 100.210 125.840 100.470 126.160 ;
        RECT 99.750 124.140 100.010 124.460 ;
        RECT 99.750 123.460 100.010 123.780 ;
        RECT 99.810 121.060 99.950 123.460 ;
        RECT 100.270 121.060 100.410 125.840 ;
        RECT 101.130 125.500 101.390 125.820 ;
        RECT 101.190 123.440 101.330 125.500 ;
        RECT 101.130 123.120 101.390 123.440 ;
        RECT 102.110 122.080 102.250 127.200 ;
        RECT 102.510 124.140 102.770 124.460 ;
        RECT 102.570 122.080 102.710 124.140 ;
        RECT 102.050 121.760 102.310 122.080 ;
        RECT 102.510 121.760 102.770 122.080 ;
        RECT 99.750 120.740 100.010 121.060 ;
        RECT 100.210 120.740 100.470 121.060 ;
        RECT 99.290 115.640 99.550 115.960 ;
        RECT 99.810 115.620 99.950 120.740 ;
        RECT 105.790 119.360 105.930 151.340 ;
        RECT 109.410 149.980 109.670 150.300 ;
        RECT 109.470 148.600 109.610 149.980 ;
        RECT 109.410 148.280 109.670 148.600 ;
        RECT 107.510 146.725 109.390 147.095 ;
        RECT 110.850 145.880 110.990 159.160 ;
        RECT 111.710 147.940 111.970 148.260 ;
        RECT 110.790 145.560 111.050 145.880 ;
        RECT 107.110 144.540 107.370 144.860 ;
        RECT 108.030 144.540 108.290 144.860 ;
        RECT 106.650 140.120 106.910 140.440 ;
        RECT 106.710 138.400 106.850 140.120 ;
        RECT 107.170 139.420 107.310 144.540 ;
        RECT 108.090 143.500 108.230 144.540 ;
        RECT 108.030 143.180 108.290 143.500 ;
        RECT 111.770 142.820 111.910 147.940 ;
        RECT 109.870 142.500 110.130 142.820 ;
        RECT 111.710 142.500 111.970 142.820 ;
        RECT 107.510 141.285 109.390 141.655 ;
        RECT 109.930 141.120 110.070 142.500 ;
        RECT 109.870 140.800 110.130 141.120 ;
        RECT 111.770 140.440 111.910 142.500 ;
        RECT 135.630 141.200 136.780 141.270 ;
        RECT 111.710 140.120 111.970 140.440 ;
        RECT 135.630 140.180 136.800 141.200 ;
        RECT 107.110 139.100 107.370 139.420 ;
        RECT 106.650 138.080 106.910 138.400 ;
        RECT 107.510 135.845 109.390 136.215 ;
        RECT 111.770 131.940 111.910 140.120 ;
        RECT 132.560 138.140 135.160 140.060 ;
        RECT 135.640 133.320 136.800 140.180 ;
        RECT 109.870 131.620 110.130 131.940 ;
        RECT 111.710 131.680 111.970 131.940 ;
        RECT 111.310 131.620 111.970 131.680 ;
        RECT 107.510 130.405 109.390 130.775 ;
        RECT 109.930 130.240 110.070 131.620 ;
        RECT 111.310 131.540 111.910 131.620 ;
        RECT 109.870 129.920 110.130 130.240 ;
        RECT 106.650 128.220 106.910 128.540 ;
        RECT 106.710 121.400 106.850 128.220 ;
        RECT 111.310 126.500 111.450 131.540 ;
        RECT 109.870 126.180 110.130 126.500 ;
        RECT 111.250 126.180 111.510 126.500 ;
        RECT 107.510 124.965 109.390 125.335 ;
        RECT 107.570 123.800 107.830 124.120 ;
        RECT 107.630 123.520 107.770 123.800 ;
        RECT 107.170 123.380 107.770 123.520 ;
        RECT 107.170 122.080 107.310 123.380 ;
        RECT 109.930 122.080 110.070 126.180 ;
        RECT 111.310 123.780 111.450 126.180 ;
        RECT 111.250 123.460 111.510 123.780 ;
        RECT 107.110 121.760 107.370 122.080 ;
        RECT 109.870 121.760 110.130 122.080 ;
        RECT 106.650 121.080 106.910 121.400 ;
        RECT 107.510 119.525 109.390 119.895 ;
        RECT 105.730 119.040 105.990 119.360 ;
        RECT 106.650 118.020 106.910 118.340 ;
        RECT 102.970 117.680 103.230 118.000 ;
        RECT 103.030 116.300 103.170 117.680 ;
        RECT 106.190 117.340 106.450 117.660 ;
        RECT 106.250 116.300 106.390 117.340 ;
        RECT 102.970 115.980 103.230 116.300 ;
        RECT 106.190 115.980 106.450 116.300 ;
        RECT 99.750 115.300 100.010 115.620 ;
        RECT 99.810 112.900 99.950 115.300 ;
        RECT 100.210 114.620 100.470 114.940 ;
        RECT 99.750 112.580 100.010 112.900 ;
        RECT 95.150 112.240 95.410 112.560 ;
        RECT 97.450 112.240 97.710 112.560 ;
        RECT 92.510 111.365 94.390 111.735 ;
        RECT 95.210 111.200 95.350 112.240 ;
        RECT 98.370 111.900 98.630 112.220 ;
        RECT 95.150 110.880 95.410 111.200 ;
        RECT 96.070 110.200 96.330 110.520 ;
        RECT 96.130 107.800 96.270 110.200 ;
        RECT 97.910 109.180 98.170 109.500 ;
        RECT 96.070 107.480 96.330 107.800 ;
        RECT 97.970 107.120 98.110 109.180 ;
        RECT 98.430 107.800 98.570 111.900 ;
        RECT 99.810 110.180 99.950 112.580 ;
        RECT 100.270 111.200 100.410 114.620 ;
        RECT 104.810 112.580 105.070 112.900 ;
        RECT 100.210 110.880 100.470 111.200 ;
        RECT 99.750 109.860 100.010 110.180 ;
        RECT 100.670 109.860 100.930 110.180 ;
        RECT 99.810 107.800 99.950 109.860 ;
        RECT 98.370 107.480 98.630 107.800 ;
        RECT 99.750 107.480 100.010 107.800 ;
        RECT 97.910 106.800 98.170 107.120 ;
        RECT 96.990 106.460 97.250 106.780 ;
        RECT 92.510 105.925 94.390 106.295 ;
        RECT 97.050 96.255 97.190 106.460 ;
        RECT 91.920 95.640 92.200 96.255 ;
        RECT 91.530 95.500 92.200 95.640 ;
        RECT 91.920 94.255 92.200 95.500 ;
        RECT 96.980 94.255 97.260 96.255 ;
        RECT 100.730 95.640 100.870 109.860 ;
        RECT 104.870 108.480 105.010 112.580 ;
        RECT 106.190 109.860 106.450 110.180 ;
        RECT 104.810 108.160 105.070 108.480 ;
        RECT 106.250 107.800 106.390 109.860 ;
        RECT 106.710 109.500 106.850 118.020 ;
        RECT 110.330 117.340 110.590 117.660 ;
        RECT 107.510 114.085 109.390 114.455 ;
        RECT 110.390 113.240 110.530 117.340 ;
        RECT 112.170 115.300 112.430 115.620 ;
        RECT 107.110 112.920 107.370 113.240 ;
        RECT 110.330 112.920 110.590 113.240 ;
        RECT 106.650 109.180 106.910 109.500 ;
        RECT 106.190 107.480 106.450 107.800 ;
        RECT 106.710 107.460 106.850 109.180 ;
        RECT 106.650 107.140 106.910 107.460 ;
        RECT 107.170 96.255 107.310 112.920 ;
        RECT 111.710 112.580 111.970 112.900 ;
        RECT 111.770 110.180 111.910 112.580 ;
        RECT 111.710 109.860 111.970 110.180 ;
        RECT 107.510 108.645 109.390 109.015 ;
        RECT 112.230 96.255 112.370 115.300 ;
        RECT 116.760 109.665 117.040 110.035 ;
        RECT 116.830 107.460 116.970 109.665 ;
        RECT 116.770 107.140 117.030 107.460 ;
        RECT 129.750 105.580 133.160 106.650 ;
        RECT 102.040 95.640 102.320 96.255 ;
        RECT 100.730 95.500 102.320 95.640 ;
        RECT 102.040 94.255 102.320 95.500 ;
        RECT 107.100 94.255 107.380 96.255 ;
        RECT 112.160 94.255 112.440 96.255 ;
        RECT 13.920 85.550 15.140 89.420 ;
        RECT 19.910 85.980 21.130 89.850 ;
        RECT 67.730 89.640 68.670 89.840 ;
        RECT 25.730 85.120 26.950 88.990 ;
        RECT 31.780 85.510 33.000 89.380 ;
        RECT 37.750 88.780 38.970 89.290 ;
        RECT 37.680 88.620 38.970 88.780 ;
        RECT 43.810 88.630 45.030 89.530 ;
        RECT 49.740 88.640 50.960 89.040 ;
        RECT 37.680 86.810 39.070 88.620 ;
        RECT 37.750 85.420 38.970 86.810 ;
        RECT 43.810 86.720 45.140 88.630 ;
        RECT 49.740 86.920 51.010 88.640 ;
        RECT 43.810 85.660 45.030 86.720 ;
        RECT 49.740 85.170 50.960 86.920 ;
        RECT 55.530 85.320 56.750 89.190 ;
        RECT 61.720 88.640 62.940 88.870 ;
        RECT 61.720 86.600 63.130 88.640 ;
        RECT 61.720 85.000 62.940 86.600 ;
        RECT 67.580 85.770 68.800 89.640 ;
        RECT 73.850 84.290 75.070 88.160 ;
        RECT 79.730 84.310 80.950 88.180 ;
        RECT 74.090 80.440 74.370 84.290 ;
        RECT 20.140 80.160 74.370 80.440 ;
        RECT 20.140 75.650 20.420 80.160 ;
        RECT 80.070 79.800 80.350 84.310 ;
        RECT 85.470 84.100 86.690 87.970 ;
        RECT 91.460 84.500 92.680 88.320 ;
        RECT 97.600 84.630 98.820 88.240 ;
        RECT 103.650 84.740 104.870 88.610 ;
        RECT 109.620 85.420 110.840 89.290 ;
        RECT 115.740 85.700 116.960 89.570 ;
        RECT 121.520 85.700 122.740 89.570 ;
        RECT 31.380 79.520 80.350 79.800 ;
        RECT 31.380 75.850 31.660 79.520 ;
        RECT 86.050 79.170 86.330 84.100 ;
        RECT 42.510 78.890 86.330 79.170 ;
        RECT 3.960 71.320 6.050 73.240 ;
        RECT 19.330 73.120 21.890 75.650 ;
        RECT 28.185 73.180 30.255 74.460 ;
        RECT 30.670 73.320 33.230 75.850 ;
        RECT 42.510 75.750 42.790 78.890 ;
        RECT 92.030 78.570 92.310 84.500 ;
        RECT 53.830 78.290 92.310 78.570 ;
        RECT 53.830 75.820 54.110 78.290 ;
        RECT 98.010 77.990 98.290 84.630 ;
        RECT 64.900 77.710 98.290 77.990 ;
        RECT 19.005 71.800 19.865 72.640 ;
        RECT 15.560 68.610 16.990 71.210 ;
        RECT 19.305 68.570 19.845 71.800 ;
        RECT 20.145 70.600 20.555 73.120 ;
        RECT 30.205 71.810 31.065 72.650 ;
        RECT 19.325 47.770 19.825 68.570 ;
        RECT 20.165 49.090 20.555 70.600 ;
        RECT 20.955 70.010 21.845 70.740 ;
        RECT 21.055 65.190 21.315 70.010 ;
        RECT 22.695 68.620 25.405 69.470 ;
        RECT 22.895 65.840 24.825 68.620 ;
        RECT 30.505 68.580 31.045 71.810 ;
        RECT 31.345 70.610 31.755 73.320 ;
        RECT 39.475 73.150 41.545 74.430 ;
        RECT 41.910 73.220 44.470 75.750 ;
        RECT 41.425 71.780 42.285 72.620 ;
        RECT 27.795 67.130 28.915 67.810 ;
        RECT 28.075 65.850 28.745 67.130 ;
        RECT 21.455 65.460 26.505 65.840 ;
        RECT 27.865 65.440 28.915 65.850 ;
        RECT 21.055 63.640 21.435 65.190 ;
        RECT 21.175 55.800 21.435 63.640 ;
        RECT 26.485 63.200 26.755 65.240 ;
        RECT 27.615 63.200 27.885 65.200 ;
        RECT 26.485 56.510 27.885 63.200 ;
        RECT 21.085 55.290 21.445 55.800 ;
        RECT 21.065 54.860 21.445 55.290 ;
        RECT 26.485 55.190 26.755 56.510 ;
        RECT 27.615 55.150 27.885 56.510 ;
        RECT 28.885 55.260 29.205 65.190 ;
        RECT 28.885 55.200 29.215 55.260 ;
        RECT 21.065 54.580 21.315 54.860 ;
        RECT 20.865 54.180 25.505 54.580 ;
        RECT 26.405 54.290 27.535 54.300 ;
        RECT 28.895 54.290 29.215 55.200 ;
        RECT 21.065 52.060 21.315 54.180 ;
        RECT 25.765 53.490 26.125 54.110 ;
        RECT 25.845 52.610 26.105 53.490 ;
        RECT 26.385 53.240 29.215 54.290 ;
        RECT 25.675 52.230 26.205 52.610 ;
        RECT 21.065 51.970 21.565 52.060 ;
        RECT 21.055 51.240 21.565 51.970 ;
        RECT 21.295 50.240 21.565 51.240 ;
        RECT 22.205 50.990 22.475 51.940 ;
        RECT 22.205 50.840 22.675 50.990 ;
        RECT 22.205 50.160 22.765 50.840 ;
        RECT 22.285 50.150 22.765 50.160 ;
        RECT 21.575 49.620 22.195 49.980 ;
        RECT 21.615 49.090 22.045 49.620 ;
        RECT 20.165 48.670 22.045 49.090 ;
        RECT 22.535 48.960 22.765 50.150 ;
        RECT 21.615 47.800 22.045 48.670 ;
        RECT 22.455 48.360 22.835 48.960 ;
        RECT 19.325 47.060 20.015 47.770 ;
        RECT 21.435 47.440 22.055 47.800 ;
        RECT 21.135 47.060 21.425 47.250 ;
        RECT 19.325 46.620 21.425 47.060 ;
        RECT 19.325 46.600 20.015 46.620 ;
        RECT 21.135 46.380 21.425 46.620 ;
        RECT 22.055 46.990 22.325 47.240 ;
        RECT 22.535 46.990 22.765 48.360 ;
        RECT 25.355 47.010 25.685 52.030 ;
        RECT 26.405 52.020 27.535 53.240 ;
        RECT 28.895 53.220 29.215 53.240 ;
        RECT 22.055 46.880 22.765 46.990 ;
        RECT 25.345 46.960 25.685 47.010 ;
        RECT 26.235 47.780 27.615 52.020 ;
        RECT 22.055 46.570 22.715 46.880 ;
        RECT 22.055 46.400 22.325 46.570 ;
        RECT 25.345 45.000 25.625 46.960 ;
        RECT 26.235 46.920 26.535 47.780 ;
        RECT 27.315 46.920 27.615 47.780 ;
        RECT 28.165 46.920 28.495 51.990 ;
        RECT 27.565 46.380 28.045 46.760 ;
        RECT 27.665 45.760 27.915 46.380 ;
        RECT 27.565 45.160 27.945 45.760 ;
        RECT 24.825 44.230 25.925 45.000 ;
        RECT 28.215 44.930 28.495 46.920 ;
        RECT 30.525 47.780 31.025 68.580 ;
        RECT 31.365 49.100 31.755 70.610 ;
        RECT 32.155 70.020 33.045 70.750 ;
        RECT 32.255 65.200 32.515 70.020 ;
        RECT 33.895 68.630 36.605 69.480 ;
        RECT 34.095 65.850 36.025 68.630 ;
        RECT 41.725 68.550 42.265 71.780 ;
        RECT 42.565 70.580 42.975 73.220 ;
        RECT 50.055 73.090 52.125 74.370 ;
        RECT 53.150 73.290 55.710 75.820 ;
        RECT 64.900 75.810 65.180 77.710 ;
        RECT 103.990 77.230 104.270 84.740 ;
        RECT 76.140 76.950 104.270 77.230 ;
        RECT 52.675 71.760 53.535 72.600 ;
        RECT 38.995 67.140 40.115 67.820 ;
        RECT 39.275 65.860 39.945 67.140 ;
        RECT 32.655 65.470 37.705 65.850 ;
        RECT 39.065 65.450 40.115 65.860 ;
        RECT 32.255 63.650 32.635 65.200 ;
        RECT 32.375 55.810 32.635 63.650 ;
        RECT 37.685 63.210 37.955 65.250 ;
        RECT 38.815 63.210 39.085 65.210 ;
        RECT 37.685 56.520 39.085 63.210 ;
        RECT 32.285 55.300 32.645 55.810 ;
        RECT 32.265 54.870 32.645 55.300 ;
        RECT 37.685 55.200 37.955 56.520 ;
        RECT 38.815 55.160 39.085 56.520 ;
        RECT 40.085 55.270 40.405 65.200 ;
        RECT 40.085 55.210 40.415 55.270 ;
        RECT 32.265 54.590 32.515 54.870 ;
        RECT 32.065 54.190 36.705 54.590 ;
        RECT 37.605 54.300 38.735 54.310 ;
        RECT 40.095 54.300 40.415 55.210 ;
        RECT 32.265 52.070 32.515 54.190 ;
        RECT 36.965 53.500 37.325 54.120 ;
        RECT 37.045 52.620 37.305 53.500 ;
        RECT 37.585 53.250 40.415 54.300 ;
        RECT 36.875 52.240 37.405 52.620 ;
        RECT 32.265 51.980 32.765 52.070 ;
        RECT 32.255 51.250 32.765 51.980 ;
        RECT 32.495 50.250 32.765 51.250 ;
        RECT 33.405 51.000 33.675 51.950 ;
        RECT 33.405 50.850 33.875 51.000 ;
        RECT 33.405 50.170 33.965 50.850 ;
        RECT 33.485 50.160 33.965 50.170 ;
        RECT 32.775 49.630 33.395 49.990 ;
        RECT 32.815 49.100 33.245 49.630 ;
        RECT 31.365 48.680 33.245 49.100 ;
        RECT 33.735 48.970 33.965 50.160 ;
        RECT 32.815 47.810 33.245 48.680 ;
        RECT 33.655 48.370 34.035 48.970 ;
        RECT 30.525 47.070 31.215 47.780 ;
        RECT 32.635 47.450 33.255 47.810 ;
        RECT 32.335 47.070 32.625 47.260 ;
        RECT 30.525 46.630 32.625 47.070 ;
        RECT 30.525 46.610 31.215 46.630 ;
        RECT 32.335 46.390 32.625 46.630 ;
        RECT 33.255 47.000 33.525 47.250 ;
        RECT 33.735 47.000 33.965 48.370 ;
        RECT 36.555 47.020 36.885 52.040 ;
        RECT 37.605 52.030 38.735 53.250 ;
        RECT 40.095 53.230 40.415 53.250 ;
        RECT 33.255 46.890 33.965 47.000 ;
        RECT 36.545 46.970 36.885 47.020 ;
        RECT 37.435 47.790 38.815 52.030 ;
        RECT 33.255 46.580 33.915 46.890 ;
        RECT 33.255 46.410 33.525 46.580 ;
        RECT 36.545 45.010 36.825 46.970 ;
        RECT 37.435 46.930 37.735 47.790 ;
        RECT 38.515 46.930 38.815 47.790 ;
        RECT 39.365 46.930 39.695 52.000 ;
        RECT 38.765 46.390 39.245 46.770 ;
        RECT 38.865 45.770 39.115 46.390 ;
        RECT 38.765 45.170 39.145 45.770 ;
        RECT 28.215 43.200 28.515 44.930 ;
        RECT 36.025 44.240 37.125 45.010 ;
        RECT 39.415 44.940 39.695 46.930 ;
        RECT 41.745 47.750 42.245 68.550 ;
        RECT 42.585 49.070 42.975 70.580 ;
        RECT 43.375 69.990 44.265 70.720 ;
        RECT 43.475 65.170 43.735 69.990 ;
        RECT 45.115 68.600 47.825 69.450 ;
        RECT 45.315 65.820 47.245 68.600 ;
        RECT 52.975 68.530 53.515 71.760 ;
        RECT 53.815 70.560 54.225 73.290 ;
        RECT 61.475 73.120 63.545 74.400 ;
        RECT 64.400 73.280 66.960 75.810 ;
        RECT 76.140 75.740 76.420 76.950 ;
        RECT 109.970 76.610 110.250 85.420 ;
        RECT 87.580 76.330 110.250 76.610 ;
        RECT 87.580 75.760 87.860 76.330 ;
        RECT 115.950 76.030 116.230 85.700 ;
        RECT 98.850 75.840 116.230 76.030 ;
        RECT 63.895 71.750 64.755 72.590 ;
        RECT 50.215 67.110 51.335 67.790 ;
        RECT 50.495 65.830 51.165 67.110 ;
        RECT 43.875 65.440 48.925 65.820 ;
        RECT 50.285 65.420 51.335 65.830 ;
        RECT 43.475 63.620 43.855 65.170 ;
        RECT 43.595 55.780 43.855 63.620 ;
        RECT 48.905 63.180 49.175 65.220 ;
        RECT 50.035 63.180 50.305 65.180 ;
        RECT 48.905 56.490 50.305 63.180 ;
        RECT 43.505 55.270 43.865 55.780 ;
        RECT 43.485 54.840 43.865 55.270 ;
        RECT 48.905 55.170 49.175 56.490 ;
        RECT 50.035 55.130 50.305 56.490 ;
        RECT 51.305 55.240 51.625 65.170 ;
        RECT 51.305 55.180 51.635 55.240 ;
        RECT 43.485 54.560 43.735 54.840 ;
        RECT 43.285 54.160 47.925 54.560 ;
        RECT 48.825 54.270 49.955 54.280 ;
        RECT 51.315 54.270 51.635 55.180 ;
        RECT 43.485 52.040 43.735 54.160 ;
        RECT 48.185 53.470 48.545 54.090 ;
        RECT 48.265 52.590 48.525 53.470 ;
        RECT 48.805 53.220 51.635 54.270 ;
        RECT 48.095 52.210 48.625 52.590 ;
        RECT 43.485 51.950 43.985 52.040 ;
        RECT 43.475 51.220 43.985 51.950 ;
        RECT 43.715 50.220 43.985 51.220 ;
        RECT 44.625 50.970 44.895 51.920 ;
        RECT 44.625 50.820 45.095 50.970 ;
        RECT 44.625 50.140 45.185 50.820 ;
        RECT 44.705 50.130 45.185 50.140 ;
        RECT 43.995 49.600 44.615 49.960 ;
        RECT 44.035 49.070 44.465 49.600 ;
        RECT 42.585 48.650 44.465 49.070 ;
        RECT 44.955 48.940 45.185 50.130 ;
        RECT 44.035 47.780 44.465 48.650 ;
        RECT 44.875 48.340 45.255 48.940 ;
        RECT 41.745 47.040 42.435 47.750 ;
        RECT 43.855 47.420 44.475 47.780 ;
        RECT 43.555 47.040 43.845 47.230 ;
        RECT 41.745 46.600 43.845 47.040 ;
        RECT 41.745 46.580 42.435 46.600 ;
        RECT 43.555 46.360 43.845 46.600 ;
        RECT 44.475 46.970 44.745 47.220 ;
        RECT 44.955 46.970 45.185 48.340 ;
        RECT 47.775 46.990 48.105 52.010 ;
        RECT 48.825 52.000 49.955 53.220 ;
        RECT 51.315 53.200 51.635 53.220 ;
        RECT 44.475 46.860 45.185 46.970 ;
        RECT 47.765 46.940 48.105 46.990 ;
        RECT 48.655 47.760 50.035 52.000 ;
        RECT 44.475 46.550 45.135 46.860 ;
        RECT 44.475 46.380 44.745 46.550 ;
        RECT 47.765 44.980 48.045 46.940 ;
        RECT 48.655 46.900 48.955 47.760 ;
        RECT 49.735 46.900 50.035 47.760 ;
        RECT 50.585 46.900 50.915 51.970 ;
        RECT 49.985 46.360 50.465 46.740 ;
        RECT 50.085 45.740 50.335 46.360 ;
        RECT 49.985 45.140 50.365 45.740 ;
        RECT 39.415 43.210 39.715 44.940 ;
        RECT 47.245 44.210 48.345 44.980 ;
        RECT 50.635 44.910 50.915 46.900 ;
        RECT 52.995 47.730 53.495 68.530 ;
        RECT 53.835 49.050 54.225 70.560 ;
        RECT 54.625 69.970 55.515 70.700 ;
        RECT 54.725 65.150 54.985 69.970 ;
        RECT 56.365 68.580 59.075 69.430 ;
        RECT 56.565 65.800 58.495 68.580 ;
        RECT 64.195 68.520 64.735 71.750 ;
        RECT 65.035 70.550 65.445 73.280 ;
        RECT 72.585 73.130 74.655 74.410 ;
        RECT 75.550 73.210 78.110 75.740 ;
        RECT 75.135 71.740 75.995 72.580 ;
        RECT 61.465 67.090 62.585 67.770 ;
        RECT 61.745 65.810 62.415 67.090 ;
        RECT 55.125 65.420 60.175 65.800 ;
        RECT 61.535 65.400 62.585 65.810 ;
        RECT 54.725 63.600 55.105 65.150 ;
        RECT 54.845 55.760 55.105 63.600 ;
        RECT 60.155 63.160 60.425 65.200 ;
        RECT 61.285 63.160 61.555 65.160 ;
        RECT 60.155 56.470 61.555 63.160 ;
        RECT 54.755 55.250 55.115 55.760 ;
        RECT 54.735 54.820 55.115 55.250 ;
        RECT 60.155 55.150 60.425 56.470 ;
        RECT 61.285 55.110 61.555 56.470 ;
        RECT 62.555 55.220 62.875 65.150 ;
        RECT 62.555 55.160 62.885 55.220 ;
        RECT 54.735 54.540 54.985 54.820 ;
        RECT 54.535 54.140 59.175 54.540 ;
        RECT 60.075 54.250 61.205 54.260 ;
        RECT 62.565 54.250 62.885 55.160 ;
        RECT 54.735 52.020 54.985 54.140 ;
        RECT 59.435 53.450 59.795 54.070 ;
        RECT 59.515 52.570 59.775 53.450 ;
        RECT 60.055 53.200 62.885 54.250 ;
        RECT 59.345 52.190 59.875 52.570 ;
        RECT 54.735 51.930 55.235 52.020 ;
        RECT 54.725 51.200 55.235 51.930 ;
        RECT 54.965 50.200 55.235 51.200 ;
        RECT 55.875 50.950 56.145 51.900 ;
        RECT 55.875 50.800 56.345 50.950 ;
        RECT 55.875 50.120 56.435 50.800 ;
        RECT 55.955 50.110 56.435 50.120 ;
        RECT 55.245 49.580 55.865 49.940 ;
        RECT 55.285 49.050 55.715 49.580 ;
        RECT 53.835 48.630 55.715 49.050 ;
        RECT 56.205 48.920 56.435 50.110 ;
        RECT 55.285 47.760 55.715 48.630 ;
        RECT 56.125 48.320 56.505 48.920 ;
        RECT 52.995 47.020 53.685 47.730 ;
        RECT 55.105 47.400 55.725 47.760 ;
        RECT 54.805 47.020 55.095 47.210 ;
        RECT 52.995 46.580 55.095 47.020 ;
        RECT 52.995 46.560 53.685 46.580 ;
        RECT 54.805 46.340 55.095 46.580 ;
        RECT 55.725 46.950 55.995 47.200 ;
        RECT 56.205 46.950 56.435 48.320 ;
        RECT 59.025 46.970 59.355 51.990 ;
        RECT 60.075 51.980 61.205 53.200 ;
        RECT 62.565 53.180 62.885 53.200 ;
        RECT 55.725 46.840 56.435 46.950 ;
        RECT 59.015 46.920 59.355 46.970 ;
        RECT 59.905 47.740 61.285 51.980 ;
        RECT 55.725 46.530 56.385 46.840 ;
        RECT 55.725 46.360 55.995 46.530 ;
        RECT 59.015 44.960 59.295 46.920 ;
        RECT 59.905 46.880 60.205 47.740 ;
        RECT 60.985 46.880 61.285 47.740 ;
        RECT 61.835 46.880 62.165 51.950 ;
        RECT 61.235 46.340 61.715 46.720 ;
        RECT 61.335 45.720 61.585 46.340 ;
        RECT 61.235 45.120 61.615 45.720 ;
        RECT 19.865 42.210 21.245 42.780 ;
        RECT 27.495 42.630 28.875 43.200 ;
        RECT 31.145 42.210 32.525 42.780 ;
        RECT 38.695 42.640 40.075 43.210 ;
        RECT 50.635 43.180 50.935 44.910 ;
        RECT 58.495 44.190 59.595 44.960 ;
        RECT 61.885 44.890 62.165 46.880 ;
        RECT 64.215 47.720 64.715 68.520 ;
        RECT 65.055 49.040 65.445 70.550 ;
        RECT 65.845 69.960 66.735 70.690 ;
        RECT 65.945 65.140 66.205 69.960 ;
        RECT 67.585 68.570 70.295 69.420 ;
        RECT 67.785 65.790 69.715 68.570 ;
        RECT 75.435 68.510 75.975 71.740 ;
        RECT 76.275 70.540 76.685 73.210 ;
        RECT 83.855 73.120 85.925 74.400 ;
        RECT 86.850 73.230 89.410 75.760 ;
        RECT 98.150 75.750 116.230 75.840 ;
        RECT 86.385 71.750 87.245 72.590 ;
        RECT 72.685 67.080 73.805 67.760 ;
        RECT 72.965 65.800 73.635 67.080 ;
        RECT 66.345 65.410 71.395 65.790 ;
        RECT 72.755 65.390 73.805 65.800 ;
        RECT 65.945 63.590 66.325 65.140 ;
        RECT 66.065 55.750 66.325 63.590 ;
        RECT 71.375 63.150 71.645 65.190 ;
        RECT 72.505 63.150 72.775 65.150 ;
        RECT 71.375 56.460 72.775 63.150 ;
        RECT 65.975 55.240 66.335 55.750 ;
        RECT 65.955 54.810 66.335 55.240 ;
        RECT 71.375 55.140 71.645 56.460 ;
        RECT 72.505 55.100 72.775 56.460 ;
        RECT 73.775 55.210 74.095 65.140 ;
        RECT 73.775 55.150 74.105 55.210 ;
        RECT 65.955 54.530 66.205 54.810 ;
        RECT 65.755 54.130 70.395 54.530 ;
        RECT 71.295 54.240 72.425 54.250 ;
        RECT 73.785 54.240 74.105 55.150 ;
        RECT 65.955 52.010 66.205 54.130 ;
        RECT 70.655 53.440 71.015 54.060 ;
        RECT 70.735 52.560 70.995 53.440 ;
        RECT 71.275 53.190 74.105 54.240 ;
        RECT 70.565 52.180 71.095 52.560 ;
        RECT 65.955 51.920 66.455 52.010 ;
        RECT 65.945 51.190 66.455 51.920 ;
        RECT 66.185 50.190 66.455 51.190 ;
        RECT 67.095 50.940 67.365 51.890 ;
        RECT 67.095 50.790 67.565 50.940 ;
        RECT 67.095 50.110 67.655 50.790 ;
        RECT 67.175 50.100 67.655 50.110 ;
        RECT 66.465 49.570 67.085 49.930 ;
        RECT 66.505 49.040 66.935 49.570 ;
        RECT 65.055 48.620 66.935 49.040 ;
        RECT 67.425 48.910 67.655 50.100 ;
        RECT 66.505 47.750 66.935 48.620 ;
        RECT 67.345 48.310 67.725 48.910 ;
        RECT 64.215 47.010 64.905 47.720 ;
        RECT 66.325 47.390 66.945 47.750 ;
        RECT 66.025 47.010 66.315 47.200 ;
        RECT 64.215 46.570 66.315 47.010 ;
        RECT 64.215 46.550 64.905 46.570 ;
        RECT 66.025 46.330 66.315 46.570 ;
        RECT 66.945 46.940 67.215 47.190 ;
        RECT 67.425 46.940 67.655 48.310 ;
        RECT 70.245 46.960 70.575 51.980 ;
        RECT 71.295 51.970 72.425 53.190 ;
        RECT 73.785 53.170 74.105 53.190 ;
        RECT 66.945 46.830 67.655 46.940 ;
        RECT 70.235 46.910 70.575 46.960 ;
        RECT 71.125 47.730 72.505 51.970 ;
        RECT 66.945 46.520 67.605 46.830 ;
        RECT 66.945 46.350 67.215 46.520 ;
        RECT 70.235 44.950 70.515 46.910 ;
        RECT 71.125 46.870 71.425 47.730 ;
        RECT 72.205 46.870 72.505 47.730 ;
        RECT 73.055 46.870 73.385 51.940 ;
        RECT 72.455 46.330 72.935 46.710 ;
        RECT 72.555 45.710 72.805 46.330 ;
        RECT 72.455 45.110 72.835 45.710 ;
        RECT 20.225 40.480 20.525 42.210 ;
        RECT 20.245 38.490 20.525 40.480 ;
        RECT 22.815 40.410 23.915 41.180 ;
        RECT 31.505 40.480 31.805 42.210 ;
        RECT 42.435 42.190 43.815 42.760 ;
        RECT 49.915 42.610 51.295 43.180 ;
        RECT 61.885 43.160 62.185 44.890 ;
        RECT 69.715 44.180 70.815 44.950 ;
        RECT 73.105 44.880 73.385 46.870 ;
        RECT 75.455 47.710 75.955 68.510 ;
        RECT 76.295 49.030 76.685 70.540 ;
        RECT 77.085 69.950 77.975 70.680 ;
        RECT 77.185 65.130 77.445 69.950 ;
        RECT 78.825 68.560 81.535 69.410 ;
        RECT 79.025 65.780 80.955 68.560 ;
        RECT 86.685 68.520 87.225 71.750 ;
        RECT 87.525 70.550 87.935 73.230 ;
        RECT 95.045 73.060 97.115 74.340 ;
        RECT 98.150 73.310 100.710 75.750 ;
        RECT 109.390 75.480 111.950 75.560 ;
        RECT 121.930 75.480 122.210 85.700 ;
        RECT 127.550 85.510 128.770 89.380 ;
        RECT 127.910 76.040 128.190 85.510 ;
        RECT 133.380 76.580 136.010 77.880 ;
        RECT 137.240 76.560 139.870 77.860 ;
        RECT 109.390 75.200 122.210 75.480 ;
        RECT 97.665 71.740 98.525 72.580 ;
        RECT 83.925 67.070 85.045 67.750 ;
        RECT 84.205 65.790 84.875 67.070 ;
        RECT 77.585 65.400 82.635 65.780 ;
        RECT 83.995 65.380 85.045 65.790 ;
        RECT 77.185 63.580 77.565 65.130 ;
        RECT 77.305 55.740 77.565 63.580 ;
        RECT 82.615 63.140 82.885 65.180 ;
        RECT 83.745 63.140 84.015 65.140 ;
        RECT 82.615 56.450 84.015 63.140 ;
        RECT 77.215 55.230 77.575 55.740 ;
        RECT 77.195 54.800 77.575 55.230 ;
        RECT 82.615 55.130 82.885 56.450 ;
        RECT 83.745 55.090 84.015 56.450 ;
        RECT 85.015 55.200 85.335 65.130 ;
        RECT 85.015 55.140 85.345 55.200 ;
        RECT 77.195 54.520 77.445 54.800 ;
        RECT 76.995 54.120 81.635 54.520 ;
        RECT 82.535 54.230 83.665 54.240 ;
        RECT 85.025 54.230 85.345 55.140 ;
        RECT 77.195 52.000 77.445 54.120 ;
        RECT 81.895 53.430 82.255 54.050 ;
        RECT 81.975 52.550 82.235 53.430 ;
        RECT 82.515 53.180 85.345 54.230 ;
        RECT 81.805 52.170 82.335 52.550 ;
        RECT 77.195 51.910 77.695 52.000 ;
        RECT 77.185 51.180 77.695 51.910 ;
        RECT 77.425 50.180 77.695 51.180 ;
        RECT 78.335 50.930 78.605 51.880 ;
        RECT 78.335 50.780 78.805 50.930 ;
        RECT 78.335 50.100 78.895 50.780 ;
        RECT 78.415 50.090 78.895 50.100 ;
        RECT 77.705 49.560 78.325 49.920 ;
        RECT 77.745 49.030 78.175 49.560 ;
        RECT 76.295 48.610 78.175 49.030 ;
        RECT 78.665 48.900 78.895 50.090 ;
        RECT 77.745 47.740 78.175 48.610 ;
        RECT 78.585 48.300 78.965 48.900 ;
        RECT 75.455 47.000 76.145 47.710 ;
        RECT 77.565 47.380 78.185 47.740 ;
        RECT 77.265 47.000 77.555 47.190 ;
        RECT 75.455 46.560 77.555 47.000 ;
        RECT 75.455 46.540 76.145 46.560 ;
        RECT 77.265 46.320 77.555 46.560 ;
        RECT 78.185 46.930 78.455 47.180 ;
        RECT 78.665 46.930 78.895 48.300 ;
        RECT 81.485 46.950 81.815 51.970 ;
        RECT 82.535 51.960 83.665 53.180 ;
        RECT 85.025 53.160 85.345 53.180 ;
        RECT 78.185 46.820 78.895 46.930 ;
        RECT 81.475 46.900 81.815 46.950 ;
        RECT 82.365 47.720 83.745 51.960 ;
        RECT 78.185 46.510 78.845 46.820 ;
        RECT 78.185 46.340 78.455 46.510 ;
        RECT 81.475 44.940 81.755 46.900 ;
        RECT 82.365 46.860 82.665 47.720 ;
        RECT 83.445 46.860 83.745 47.720 ;
        RECT 84.295 46.860 84.625 51.930 ;
        RECT 83.695 46.320 84.175 46.700 ;
        RECT 83.795 45.700 84.045 46.320 ;
        RECT 83.695 45.100 84.075 45.700 ;
        RECT 53.655 42.190 55.035 42.760 ;
        RECT 61.165 42.590 62.545 43.160 ;
        RECT 73.105 43.150 73.405 44.880 ;
        RECT 80.955 44.170 82.055 44.940 ;
        RECT 84.345 44.870 84.625 46.860 ;
        RECT 86.705 47.720 87.205 68.520 ;
        RECT 87.545 49.040 87.935 70.550 ;
        RECT 88.335 69.960 89.225 70.690 ;
        RECT 88.435 65.140 88.695 69.960 ;
        RECT 90.075 68.570 92.785 69.420 ;
        RECT 90.275 65.790 92.205 68.570 ;
        RECT 97.965 68.510 98.505 71.740 ;
        RECT 98.805 70.540 99.215 73.310 ;
        RECT 106.455 73.110 108.525 74.390 ;
        RECT 109.390 73.030 111.950 75.200 ;
        RECT 125.760 74.810 128.190 76.040 ;
        RECT 121.290 74.790 128.190 74.810 ;
        RECT 120.600 74.530 128.190 74.790 ;
        RECT 117.655 73.110 119.725 74.390 ;
        RECT 120.600 73.180 128.160 74.530 ;
        RECT 129.505 73.190 131.575 74.470 ;
        RECT 120.600 73.110 126.160 73.180 ;
        RECT 108.935 71.740 109.795 72.580 ;
        RECT 95.175 67.080 96.295 67.760 ;
        RECT 95.455 65.800 96.125 67.080 ;
        RECT 88.835 65.410 93.885 65.790 ;
        RECT 95.245 65.390 96.295 65.800 ;
        RECT 88.435 63.590 88.815 65.140 ;
        RECT 88.555 55.750 88.815 63.590 ;
        RECT 93.865 63.150 94.135 65.190 ;
        RECT 94.995 63.150 95.265 65.150 ;
        RECT 93.865 56.460 95.265 63.150 ;
        RECT 88.465 55.240 88.825 55.750 ;
        RECT 88.445 54.810 88.825 55.240 ;
        RECT 93.865 55.140 94.135 56.460 ;
        RECT 94.995 55.100 95.265 56.460 ;
        RECT 96.265 55.210 96.585 65.140 ;
        RECT 96.265 55.150 96.595 55.210 ;
        RECT 88.445 54.530 88.695 54.810 ;
        RECT 88.245 54.130 92.885 54.530 ;
        RECT 93.785 54.240 94.915 54.250 ;
        RECT 96.275 54.240 96.595 55.150 ;
        RECT 88.445 52.010 88.695 54.130 ;
        RECT 93.145 53.440 93.505 54.060 ;
        RECT 93.225 52.560 93.485 53.440 ;
        RECT 93.765 53.190 96.595 54.240 ;
        RECT 93.055 52.180 93.585 52.560 ;
        RECT 88.445 51.920 88.945 52.010 ;
        RECT 88.435 51.190 88.945 51.920 ;
        RECT 88.675 50.190 88.945 51.190 ;
        RECT 89.585 50.940 89.855 51.890 ;
        RECT 89.585 50.790 90.055 50.940 ;
        RECT 89.585 50.110 90.145 50.790 ;
        RECT 89.665 50.100 90.145 50.110 ;
        RECT 88.955 49.570 89.575 49.930 ;
        RECT 88.995 49.040 89.425 49.570 ;
        RECT 87.545 48.620 89.425 49.040 ;
        RECT 89.915 48.910 90.145 50.100 ;
        RECT 88.995 47.750 89.425 48.620 ;
        RECT 89.835 48.310 90.215 48.910 ;
        RECT 86.705 47.010 87.395 47.720 ;
        RECT 88.815 47.390 89.435 47.750 ;
        RECT 88.515 47.010 88.805 47.200 ;
        RECT 86.705 46.570 88.805 47.010 ;
        RECT 86.705 46.550 87.395 46.570 ;
        RECT 88.515 46.330 88.805 46.570 ;
        RECT 89.435 46.940 89.705 47.190 ;
        RECT 89.915 46.940 90.145 48.310 ;
        RECT 92.735 46.960 93.065 51.980 ;
        RECT 93.785 51.970 94.915 53.190 ;
        RECT 96.275 53.170 96.595 53.190 ;
        RECT 89.435 46.830 90.145 46.940 ;
        RECT 92.725 46.910 93.065 46.960 ;
        RECT 93.615 47.730 94.995 51.970 ;
        RECT 89.435 46.520 90.095 46.830 ;
        RECT 89.435 46.350 89.705 46.520 ;
        RECT 92.725 44.950 93.005 46.910 ;
        RECT 93.615 46.870 93.915 47.730 ;
        RECT 94.695 46.870 94.995 47.730 ;
        RECT 95.545 46.870 95.875 51.940 ;
        RECT 94.945 46.330 95.425 46.710 ;
        RECT 95.045 45.710 95.295 46.330 ;
        RECT 94.945 45.110 95.325 45.710 ;
        RECT 64.855 42.190 66.235 42.760 ;
        RECT 72.385 42.580 73.765 43.150 ;
        RECT 84.345 43.140 84.645 44.870 ;
        RECT 92.205 44.180 93.305 44.950 ;
        RECT 95.595 44.880 95.875 46.870 ;
        RECT 97.985 47.710 98.485 68.510 ;
        RECT 98.825 49.030 99.215 70.540 ;
        RECT 99.615 69.950 100.505 70.680 ;
        RECT 99.715 65.130 99.975 69.950 ;
        RECT 101.355 68.560 104.065 69.410 ;
        RECT 101.555 65.780 103.485 68.560 ;
        RECT 109.235 68.510 109.775 71.740 ;
        RECT 110.075 70.540 110.485 73.030 ;
        RECT 120.185 71.740 121.045 72.580 ;
        RECT 106.455 67.070 107.575 67.750 ;
        RECT 106.735 65.790 107.405 67.070 ;
        RECT 100.115 65.400 105.165 65.780 ;
        RECT 106.525 65.380 107.575 65.790 ;
        RECT 99.715 63.580 100.095 65.130 ;
        RECT 99.835 55.740 100.095 63.580 ;
        RECT 105.145 63.140 105.415 65.180 ;
        RECT 106.275 63.140 106.545 65.140 ;
        RECT 105.145 56.450 106.545 63.140 ;
        RECT 99.745 55.230 100.105 55.740 ;
        RECT 99.725 54.800 100.105 55.230 ;
        RECT 105.145 55.130 105.415 56.450 ;
        RECT 106.275 55.090 106.545 56.450 ;
        RECT 107.545 55.200 107.865 65.130 ;
        RECT 107.545 55.140 107.875 55.200 ;
        RECT 99.725 54.520 99.975 54.800 ;
        RECT 99.525 54.120 104.165 54.520 ;
        RECT 105.065 54.230 106.195 54.240 ;
        RECT 107.555 54.230 107.875 55.140 ;
        RECT 99.725 52.000 99.975 54.120 ;
        RECT 104.425 53.430 104.785 54.050 ;
        RECT 104.505 52.550 104.765 53.430 ;
        RECT 105.045 53.180 107.875 54.230 ;
        RECT 104.335 52.170 104.865 52.550 ;
        RECT 99.725 51.910 100.225 52.000 ;
        RECT 99.715 51.180 100.225 51.910 ;
        RECT 99.955 50.180 100.225 51.180 ;
        RECT 100.865 50.930 101.135 51.880 ;
        RECT 100.865 50.780 101.335 50.930 ;
        RECT 100.865 50.100 101.425 50.780 ;
        RECT 100.945 50.090 101.425 50.100 ;
        RECT 100.235 49.560 100.855 49.920 ;
        RECT 100.275 49.030 100.705 49.560 ;
        RECT 98.825 48.610 100.705 49.030 ;
        RECT 101.195 48.900 101.425 50.090 ;
        RECT 100.275 47.740 100.705 48.610 ;
        RECT 101.115 48.300 101.495 48.900 ;
        RECT 97.985 47.000 98.675 47.710 ;
        RECT 100.095 47.380 100.715 47.740 ;
        RECT 99.795 47.000 100.085 47.190 ;
        RECT 97.985 46.560 100.085 47.000 ;
        RECT 97.985 46.540 98.675 46.560 ;
        RECT 99.795 46.320 100.085 46.560 ;
        RECT 100.715 46.930 100.985 47.180 ;
        RECT 101.195 46.930 101.425 48.300 ;
        RECT 104.015 46.950 104.345 51.970 ;
        RECT 105.065 51.960 106.195 53.180 ;
        RECT 107.555 53.160 107.875 53.180 ;
        RECT 100.715 46.820 101.425 46.930 ;
        RECT 104.005 46.900 104.345 46.950 ;
        RECT 104.895 47.720 106.275 51.960 ;
        RECT 100.715 46.510 101.375 46.820 ;
        RECT 100.715 46.340 100.985 46.510 ;
        RECT 104.005 44.940 104.285 46.900 ;
        RECT 104.895 46.860 105.195 47.720 ;
        RECT 105.975 46.860 106.275 47.720 ;
        RECT 106.825 46.860 107.155 51.930 ;
        RECT 106.225 46.320 106.705 46.700 ;
        RECT 106.325 45.700 106.575 46.320 ;
        RECT 106.225 45.100 106.605 45.700 ;
        RECT 95.595 43.150 95.895 44.880 ;
        RECT 103.485 44.170 104.585 44.940 ;
        RECT 106.875 44.870 107.155 46.860 ;
        RECT 109.255 47.710 109.755 68.510 ;
        RECT 110.095 49.030 110.485 70.540 ;
        RECT 110.885 69.950 111.775 70.680 ;
        RECT 110.985 65.130 111.245 69.950 ;
        RECT 112.625 68.560 115.335 69.410 ;
        RECT 112.825 65.780 114.755 68.560 ;
        RECT 120.485 68.510 121.025 71.740 ;
        RECT 121.325 70.540 121.735 73.110 ;
        RECT 132.925 70.810 133.225 70.900 ;
        RECT 117.725 67.070 118.845 67.750 ;
        RECT 118.005 65.790 118.675 67.070 ;
        RECT 111.385 65.400 116.435 65.780 ;
        RECT 117.795 65.380 118.845 65.790 ;
        RECT 110.985 63.580 111.365 65.130 ;
        RECT 111.105 55.740 111.365 63.580 ;
        RECT 116.415 63.140 116.685 65.180 ;
        RECT 117.545 63.140 117.815 65.140 ;
        RECT 116.415 56.450 117.815 63.140 ;
        RECT 111.015 55.230 111.375 55.740 ;
        RECT 110.995 54.800 111.375 55.230 ;
        RECT 116.415 55.130 116.685 56.450 ;
        RECT 117.545 55.090 117.815 56.450 ;
        RECT 118.815 55.200 119.135 65.130 ;
        RECT 118.815 55.140 119.145 55.200 ;
        RECT 110.995 54.520 111.245 54.800 ;
        RECT 110.795 54.120 115.435 54.520 ;
        RECT 116.335 54.230 117.465 54.240 ;
        RECT 118.825 54.230 119.145 55.140 ;
        RECT 110.995 52.000 111.245 54.120 ;
        RECT 115.695 53.430 116.055 54.050 ;
        RECT 115.775 52.550 116.035 53.430 ;
        RECT 116.315 53.180 119.145 54.230 ;
        RECT 115.605 52.170 116.135 52.550 ;
        RECT 110.995 51.910 111.495 52.000 ;
        RECT 110.985 51.180 111.495 51.910 ;
        RECT 111.225 50.180 111.495 51.180 ;
        RECT 112.135 50.930 112.405 51.880 ;
        RECT 112.135 50.780 112.605 50.930 ;
        RECT 112.135 50.100 112.695 50.780 ;
        RECT 112.215 50.090 112.695 50.100 ;
        RECT 111.505 49.560 112.125 49.920 ;
        RECT 111.545 49.030 111.975 49.560 ;
        RECT 110.095 48.610 111.975 49.030 ;
        RECT 112.465 48.900 112.695 50.090 ;
        RECT 111.545 47.740 111.975 48.610 ;
        RECT 112.385 48.300 112.765 48.900 ;
        RECT 109.255 47.000 109.945 47.710 ;
        RECT 111.365 47.380 111.985 47.740 ;
        RECT 111.065 47.000 111.355 47.190 ;
        RECT 109.255 46.560 111.355 47.000 ;
        RECT 109.255 46.540 109.945 46.560 ;
        RECT 111.065 46.320 111.355 46.560 ;
        RECT 111.985 46.930 112.255 47.180 ;
        RECT 112.465 46.930 112.695 48.300 ;
        RECT 115.285 46.950 115.615 51.970 ;
        RECT 116.335 51.960 117.465 53.180 ;
        RECT 118.825 53.160 119.145 53.180 ;
        RECT 111.985 46.820 112.695 46.930 ;
        RECT 115.275 46.900 115.615 46.950 ;
        RECT 116.165 47.720 117.545 51.960 ;
        RECT 111.985 46.510 112.645 46.820 ;
        RECT 111.985 46.340 112.255 46.510 ;
        RECT 115.275 44.940 115.555 46.900 ;
        RECT 116.165 46.860 116.465 47.720 ;
        RECT 117.245 46.860 117.545 47.720 ;
        RECT 118.095 46.860 118.425 51.930 ;
        RECT 117.495 46.320 117.975 46.700 ;
        RECT 117.595 45.700 117.845 46.320 ;
        RECT 117.495 45.100 117.875 45.700 ;
        RECT 20.795 39.650 21.175 40.250 ;
        RECT 20.825 39.030 21.075 39.650 ;
        RECT 20.695 38.650 21.175 39.030 ;
        RECT 20.245 33.420 20.575 38.490 ;
        RECT 21.125 37.630 21.425 38.490 ;
        RECT 22.205 37.630 22.505 38.490 ;
        RECT 23.115 38.450 23.395 40.410 ;
        RECT 26.415 38.840 26.685 39.010 ;
        RECT 26.025 38.530 26.685 38.840 ;
        RECT 21.125 33.390 22.505 37.630 ;
        RECT 23.055 38.400 23.395 38.450 ;
        RECT 25.975 38.420 26.685 38.530 ;
        RECT 19.525 32.170 19.845 32.190 ;
        RECT 21.205 32.170 22.335 33.390 ;
        RECT 23.055 33.380 23.385 38.400 ;
        RECT 25.975 37.050 26.205 38.420 ;
        RECT 26.415 38.170 26.685 38.420 ;
        RECT 27.315 38.790 27.605 39.030 ;
        RECT 28.725 38.790 29.415 38.810 ;
        RECT 27.315 38.350 29.415 38.790 ;
        RECT 27.315 38.160 27.605 38.350 ;
        RECT 26.685 37.610 27.305 37.970 ;
        RECT 28.725 37.640 29.415 38.350 ;
        RECT 25.905 36.450 26.285 37.050 ;
        RECT 26.695 36.740 27.125 37.610 ;
        RECT 25.975 35.260 26.205 36.450 ;
        RECT 26.695 36.320 28.575 36.740 ;
        RECT 26.695 35.790 27.125 36.320 ;
        RECT 26.545 35.430 27.165 35.790 ;
        RECT 25.975 35.250 26.455 35.260 ;
        RECT 25.975 34.570 26.535 35.250 ;
        RECT 26.065 34.420 26.535 34.570 ;
        RECT 26.265 33.470 26.535 34.420 ;
        RECT 27.175 34.170 27.445 35.170 ;
        RECT 27.175 33.440 27.685 34.170 ;
        RECT 27.175 33.350 27.675 33.440 ;
        RECT 22.535 32.800 23.065 33.180 ;
        RECT 19.525 31.120 22.355 32.170 ;
        RECT 22.635 31.920 22.895 32.800 ;
        RECT 22.615 31.300 22.975 31.920 ;
        RECT 27.425 31.230 27.675 33.350 ;
        RECT 19.525 30.210 19.845 31.120 ;
        RECT 21.205 31.110 22.335 31.120 ;
        RECT 23.235 30.830 27.875 31.230 ;
        RECT 27.425 30.550 27.675 30.830 ;
        RECT 19.525 30.150 19.855 30.210 ;
        RECT 19.535 20.220 19.855 30.150 ;
        RECT 20.855 28.900 21.125 30.260 ;
        RECT 21.985 28.900 22.255 30.220 ;
        RECT 27.295 30.120 27.675 30.550 ;
        RECT 27.295 29.610 27.655 30.120 ;
        RECT 20.855 22.210 22.255 28.900 ;
        RECT 20.855 20.210 21.125 22.210 ;
        RECT 21.985 20.170 22.255 22.210 ;
        RECT 27.305 21.770 27.565 29.610 ;
        RECT 27.305 20.220 27.685 21.770 ;
        RECT 19.825 19.560 20.875 19.970 ;
        RECT 22.235 19.570 27.285 19.950 ;
        RECT 19.995 18.280 20.665 19.560 ;
        RECT 19.825 17.600 20.945 18.280 ;
        RECT 23.915 16.790 25.845 19.570 ;
        RECT 23.335 15.940 26.045 16.790 ;
        RECT 27.425 15.400 27.685 20.220 ;
        RECT 26.895 14.670 27.785 15.400 ;
        RECT 28.185 14.810 28.575 36.320 ;
        RECT 28.915 16.840 29.415 37.640 ;
        RECT 31.525 38.490 31.805 40.480 ;
        RECT 34.095 40.410 35.195 41.180 ;
        RECT 42.795 40.460 43.095 42.190 ;
        RECT 32.075 39.650 32.455 40.250 ;
        RECT 32.105 39.030 32.355 39.650 ;
        RECT 31.975 38.650 32.455 39.030 ;
        RECT 31.525 33.420 31.855 38.490 ;
        RECT 32.405 37.630 32.705 38.490 ;
        RECT 33.485 37.630 33.785 38.490 ;
        RECT 34.395 38.450 34.675 40.410 ;
        RECT 37.695 38.840 37.965 39.010 ;
        RECT 37.305 38.530 37.965 38.840 ;
        RECT 32.405 33.390 33.785 37.630 ;
        RECT 34.335 38.400 34.675 38.450 ;
        RECT 37.255 38.420 37.965 38.530 ;
        RECT 30.805 32.170 31.125 32.190 ;
        RECT 32.485 32.170 33.615 33.390 ;
        RECT 34.335 33.380 34.665 38.400 ;
        RECT 37.255 37.050 37.485 38.420 ;
        RECT 37.695 38.170 37.965 38.420 ;
        RECT 38.595 38.790 38.885 39.030 ;
        RECT 40.005 38.790 40.695 38.810 ;
        RECT 38.595 38.350 40.695 38.790 ;
        RECT 38.595 38.160 38.885 38.350 ;
        RECT 37.965 37.610 38.585 37.970 ;
        RECT 40.005 37.640 40.695 38.350 ;
        RECT 37.185 36.450 37.565 37.050 ;
        RECT 37.975 36.740 38.405 37.610 ;
        RECT 37.255 35.260 37.485 36.450 ;
        RECT 37.975 36.320 39.855 36.740 ;
        RECT 37.975 35.790 38.405 36.320 ;
        RECT 37.825 35.430 38.445 35.790 ;
        RECT 37.255 35.250 37.735 35.260 ;
        RECT 37.255 34.570 37.815 35.250 ;
        RECT 37.345 34.420 37.815 34.570 ;
        RECT 37.545 33.470 37.815 34.420 ;
        RECT 38.455 34.170 38.725 35.170 ;
        RECT 38.455 33.440 38.965 34.170 ;
        RECT 38.455 33.350 38.955 33.440 ;
        RECT 33.815 32.800 34.345 33.180 ;
        RECT 30.805 31.120 33.635 32.170 ;
        RECT 33.915 31.920 34.175 32.800 ;
        RECT 33.895 31.300 34.255 31.920 ;
        RECT 38.705 31.230 38.955 33.350 ;
        RECT 30.805 30.210 31.125 31.120 ;
        RECT 32.485 31.110 33.615 31.120 ;
        RECT 34.515 30.830 39.155 31.230 ;
        RECT 38.705 30.550 38.955 30.830 ;
        RECT 30.805 30.150 31.135 30.210 ;
        RECT 30.815 20.220 31.135 30.150 ;
        RECT 32.135 28.900 32.405 30.260 ;
        RECT 33.265 28.900 33.535 30.220 ;
        RECT 38.575 30.120 38.955 30.550 ;
        RECT 38.575 29.610 38.935 30.120 ;
        RECT 32.135 22.210 33.535 28.900 ;
        RECT 32.135 20.210 32.405 22.210 ;
        RECT 33.265 20.170 33.535 22.210 ;
        RECT 38.585 21.770 38.845 29.610 ;
        RECT 38.585 20.220 38.965 21.770 ;
        RECT 31.105 19.560 32.155 19.970 ;
        RECT 33.515 19.570 38.565 19.950 ;
        RECT 31.275 18.280 31.945 19.560 ;
        RECT 31.105 17.600 32.225 18.280 ;
        RECT 28.185 12.290 28.595 14.810 ;
        RECT 28.895 13.610 29.435 16.840 ;
        RECT 35.195 16.790 37.125 19.570 ;
        RECT 34.615 15.940 37.325 16.790 ;
        RECT 38.705 15.400 38.965 20.220 ;
        RECT 38.175 14.670 39.065 15.400 ;
        RECT 39.465 14.810 39.855 36.320 ;
        RECT 40.195 16.840 40.695 37.640 ;
        RECT 42.815 38.470 43.095 40.460 ;
        RECT 45.385 40.390 46.485 41.160 ;
        RECT 54.015 40.460 54.315 42.190 ;
        RECT 43.365 39.630 43.745 40.230 ;
        RECT 43.395 39.010 43.645 39.630 ;
        RECT 43.265 38.630 43.745 39.010 ;
        RECT 42.815 33.400 43.145 38.470 ;
        RECT 43.695 37.610 43.995 38.470 ;
        RECT 44.775 37.610 45.075 38.470 ;
        RECT 45.685 38.430 45.965 40.390 ;
        RECT 48.985 38.820 49.255 38.990 ;
        RECT 48.595 38.510 49.255 38.820 ;
        RECT 43.695 33.370 45.075 37.610 ;
        RECT 45.625 38.380 45.965 38.430 ;
        RECT 48.545 38.400 49.255 38.510 ;
        RECT 42.095 32.150 42.415 32.170 ;
        RECT 43.775 32.150 44.905 33.370 ;
        RECT 45.625 33.360 45.955 38.380 ;
        RECT 48.545 37.030 48.775 38.400 ;
        RECT 48.985 38.150 49.255 38.400 ;
        RECT 49.885 38.770 50.175 39.010 ;
        RECT 51.295 38.770 51.985 38.790 ;
        RECT 49.885 38.330 51.985 38.770 ;
        RECT 49.885 38.140 50.175 38.330 ;
        RECT 49.255 37.590 49.875 37.950 ;
        RECT 51.295 37.620 51.985 38.330 ;
        RECT 48.475 36.430 48.855 37.030 ;
        RECT 49.265 36.720 49.695 37.590 ;
        RECT 48.545 35.240 48.775 36.430 ;
        RECT 49.265 36.300 51.145 36.720 ;
        RECT 49.265 35.770 49.695 36.300 ;
        RECT 49.115 35.410 49.735 35.770 ;
        RECT 48.545 35.230 49.025 35.240 ;
        RECT 48.545 34.550 49.105 35.230 ;
        RECT 48.635 34.400 49.105 34.550 ;
        RECT 48.835 33.450 49.105 34.400 ;
        RECT 49.745 34.150 50.015 35.150 ;
        RECT 49.745 33.420 50.255 34.150 ;
        RECT 49.745 33.330 50.245 33.420 ;
        RECT 45.105 32.780 45.635 33.160 ;
        RECT 42.095 31.100 44.925 32.150 ;
        RECT 45.205 31.900 45.465 32.780 ;
        RECT 45.185 31.280 45.545 31.900 ;
        RECT 49.995 31.210 50.245 33.330 ;
        RECT 42.095 30.190 42.415 31.100 ;
        RECT 43.775 31.090 44.905 31.100 ;
        RECT 45.805 30.810 50.445 31.210 ;
        RECT 49.995 30.530 50.245 30.810 ;
        RECT 42.095 30.130 42.425 30.190 ;
        RECT 42.105 20.200 42.425 30.130 ;
        RECT 43.425 28.880 43.695 30.240 ;
        RECT 44.555 28.880 44.825 30.200 ;
        RECT 49.865 30.100 50.245 30.530 ;
        RECT 49.865 29.590 50.225 30.100 ;
        RECT 43.425 22.190 44.825 28.880 ;
        RECT 43.425 20.190 43.695 22.190 ;
        RECT 44.555 20.150 44.825 22.190 ;
        RECT 49.875 21.750 50.135 29.590 ;
        RECT 49.875 20.200 50.255 21.750 ;
        RECT 42.395 19.540 43.445 19.950 ;
        RECT 44.805 19.550 49.855 19.930 ;
        RECT 42.565 18.260 43.235 19.540 ;
        RECT 42.395 17.580 43.515 18.260 ;
        RECT 28.875 12.770 29.735 13.610 ;
        RECT 28.185 11.950 30.415 12.290 ;
        RECT 39.465 11.990 39.875 14.810 ;
        RECT 40.175 13.610 40.715 16.840 ;
        RECT 46.485 16.770 48.415 19.550 ;
        RECT 45.905 15.920 48.615 16.770 ;
        RECT 49.995 15.380 50.255 20.200 ;
        RECT 49.465 14.650 50.355 15.380 ;
        RECT 50.755 14.790 51.145 36.300 ;
        RECT 51.485 16.820 51.985 37.620 ;
        RECT 54.035 38.470 54.315 40.460 ;
        RECT 56.605 40.390 57.705 41.160 ;
        RECT 65.215 40.460 65.515 42.190 ;
        RECT 76.145 42.180 77.525 42.750 ;
        RECT 83.625 42.570 85.005 43.140 ;
        RECT 87.385 42.200 88.765 42.770 ;
        RECT 94.875 42.580 96.255 43.150 ;
        RECT 106.875 43.140 107.175 44.870 ;
        RECT 114.755 44.170 115.855 44.940 ;
        RECT 118.145 44.870 118.425 46.860 ;
        RECT 120.505 47.710 121.005 68.510 ;
        RECT 121.345 49.030 121.735 70.540 ;
        RECT 122.135 69.950 123.025 70.680 ;
        RECT 132.615 70.040 134.265 70.810 ;
        RECT 122.235 65.130 122.495 69.950 ;
        RECT 123.875 68.560 126.585 69.410 ;
        RECT 124.075 65.780 126.005 68.560 ;
        RECT 128.975 67.070 130.095 67.750 ;
        RECT 129.255 65.790 129.925 67.070 ;
        RECT 122.635 65.400 127.685 65.780 ;
        RECT 129.045 65.380 130.095 65.790 ;
        RECT 132.925 65.180 133.225 70.040 ;
        RECT 137.675 68.690 139.075 69.460 ;
        RECT 138.385 65.740 138.645 68.690 ;
        RECT 149.410 68.420 150.690 69.620 ;
        RECT 149.480 65.810 150.640 68.420 ;
        RECT 133.365 65.380 138.645 65.740 ;
        RECT 122.235 63.580 122.615 65.130 ;
        RECT 122.355 55.740 122.615 63.580 ;
        RECT 127.665 63.140 127.935 65.180 ;
        RECT 128.795 63.140 129.065 65.140 ;
        RECT 127.665 56.450 129.065 63.140 ;
        RECT 122.265 55.230 122.625 55.740 ;
        RECT 122.245 54.800 122.625 55.230 ;
        RECT 127.665 55.130 127.935 56.450 ;
        RECT 128.795 55.090 129.065 56.450 ;
        RECT 130.065 55.200 130.385 65.130 ;
        RECT 132.925 61.010 133.355 65.180 ;
        RECT 138.385 65.150 138.645 65.380 ;
        RECT 138.385 64.770 138.675 65.150 ;
        RECT 130.065 55.140 130.395 55.200 ;
        RECT 133.055 55.190 133.355 61.010 ;
        RECT 122.245 54.520 122.495 54.800 ;
        RECT 122.045 54.120 126.685 54.520 ;
        RECT 127.585 54.230 128.715 54.240 ;
        RECT 130.075 54.230 130.395 55.140 ;
        RECT 138.395 55.080 138.675 64.770 ;
        RECT 149.390 64.610 150.670 65.810 ;
        RECT 122.245 52.000 122.495 54.120 ;
        RECT 126.945 53.430 127.305 54.050 ;
        RECT 127.025 52.550 127.285 53.430 ;
        RECT 127.565 53.180 130.395 54.230 ;
        RECT 126.855 52.170 127.385 52.550 ;
        RECT 122.245 51.910 122.745 52.000 ;
        RECT 122.235 51.180 122.745 51.910 ;
        RECT 122.475 50.180 122.745 51.180 ;
        RECT 123.385 50.930 123.655 51.880 ;
        RECT 123.385 50.780 123.855 50.930 ;
        RECT 123.385 50.100 123.945 50.780 ;
        RECT 123.465 50.090 123.945 50.100 ;
        RECT 122.755 49.560 123.375 49.920 ;
        RECT 122.795 49.030 123.225 49.560 ;
        RECT 121.345 48.610 123.225 49.030 ;
        RECT 123.715 48.900 123.945 50.090 ;
        RECT 122.795 47.740 123.225 48.610 ;
        RECT 123.635 48.300 124.015 48.900 ;
        RECT 120.505 47.000 121.195 47.710 ;
        RECT 122.615 47.380 123.235 47.740 ;
        RECT 122.315 47.000 122.605 47.190 ;
        RECT 120.505 46.560 122.605 47.000 ;
        RECT 120.505 46.540 121.195 46.560 ;
        RECT 122.315 46.320 122.605 46.560 ;
        RECT 123.235 46.930 123.505 47.180 ;
        RECT 123.715 46.930 123.945 48.300 ;
        RECT 126.535 46.950 126.865 51.970 ;
        RECT 127.585 51.960 128.715 53.180 ;
        RECT 130.075 53.160 130.395 53.180 ;
        RECT 123.235 46.820 123.945 46.930 ;
        RECT 126.525 46.900 126.865 46.950 ;
        RECT 127.415 47.720 128.795 51.960 ;
        RECT 123.235 46.510 123.895 46.820 ;
        RECT 123.235 46.340 123.505 46.510 ;
        RECT 126.525 44.940 126.805 46.900 ;
        RECT 127.415 46.860 127.715 47.720 ;
        RECT 128.495 46.860 128.795 47.720 ;
        RECT 129.345 46.860 129.675 51.930 ;
        RECT 128.745 46.320 129.225 46.700 ;
        RECT 128.845 45.700 129.095 46.320 ;
        RECT 128.745 45.100 129.125 45.700 ;
        RECT 118.145 43.140 118.445 44.870 ;
        RECT 126.005 44.170 127.105 44.940 ;
        RECT 129.395 44.870 129.675 46.860 ;
        RECT 129.395 43.140 129.695 44.870 ;
        RECT 98.595 42.220 99.975 42.790 ;
        RECT 106.155 42.570 107.535 43.140 ;
        RECT 109.795 42.260 111.175 42.830 ;
        RECT 117.425 42.570 118.805 43.140 ;
        RECT 121.005 42.280 122.385 42.850 ;
        RECT 128.675 42.570 130.055 43.140 ;
        RECT 54.585 39.630 54.965 40.230 ;
        RECT 54.615 39.010 54.865 39.630 ;
        RECT 54.485 38.630 54.965 39.010 ;
        RECT 54.035 33.400 54.365 38.470 ;
        RECT 54.915 37.610 55.215 38.470 ;
        RECT 55.995 37.610 56.295 38.470 ;
        RECT 56.905 38.430 57.185 40.390 ;
        RECT 60.205 38.820 60.475 38.990 ;
        RECT 59.815 38.510 60.475 38.820 ;
        RECT 54.915 33.370 56.295 37.610 ;
        RECT 56.845 38.380 57.185 38.430 ;
        RECT 59.765 38.400 60.475 38.510 ;
        RECT 53.315 32.150 53.635 32.170 ;
        RECT 54.995 32.150 56.125 33.370 ;
        RECT 56.845 33.360 57.175 38.380 ;
        RECT 59.765 37.030 59.995 38.400 ;
        RECT 60.205 38.150 60.475 38.400 ;
        RECT 61.105 38.770 61.395 39.010 ;
        RECT 62.515 38.770 63.205 38.790 ;
        RECT 61.105 38.330 63.205 38.770 ;
        RECT 61.105 38.140 61.395 38.330 ;
        RECT 60.475 37.590 61.095 37.950 ;
        RECT 62.515 37.620 63.205 38.330 ;
        RECT 59.695 36.430 60.075 37.030 ;
        RECT 60.485 36.720 60.915 37.590 ;
        RECT 59.765 35.240 59.995 36.430 ;
        RECT 60.485 36.300 62.365 36.720 ;
        RECT 60.485 35.770 60.915 36.300 ;
        RECT 60.335 35.410 60.955 35.770 ;
        RECT 59.765 35.230 60.245 35.240 ;
        RECT 59.765 34.550 60.325 35.230 ;
        RECT 59.855 34.400 60.325 34.550 ;
        RECT 60.055 33.450 60.325 34.400 ;
        RECT 60.965 34.150 61.235 35.150 ;
        RECT 60.965 33.420 61.475 34.150 ;
        RECT 60.965 33.330 61.465 33.420 ;
        RECT 56.325 32.780 56.855 33.160 ;
        RECT 53.315 31.100 56.145 32.150 ;
        RECT 56.425 31.900 56.685 32.780 ;
        RECT 56.405 31.280 56.765 31.900 ;
        RECT 61.215 31.210 61.465 33.330 ;
        RECT 53.315 30.190 53.635 31.100 ;
        RECT 54.995 31.090 56.125 31.100 ;
        RECT 57.025 30.810 61.665 31.210 ;
        RECT 61.215 30.530 61.465 30.810 ;
        RECT 53.315 30.130 53.645 30.190 ;
        RECT 53.325 20.200 53.645 30.130 ;
        RECT 54.645 28.880 54.915 30.240 ;
        RECT 55.775 28.880 56.045 30.200 ;
        RECT 61.085 30.100 61.465 30.530 ;
        RECT 61.085 29.590 61.445 30.100 ;
        RECT 54.645 22.190 56.045 28.880 ;
        RECT 54.645 20.190 54.915 22.190 ;
        RECT 55.775 20.150 56.045 22.190 ;
        RECT 61.095 21.750 61.355 29.590 ;
        RECT 61.095 20.200 61.475 21.750 ;
        RECT 53.615 19.540 54.665 19.950 ;
        RECT 56.025 19.550 61.075 19.930 ;
        RECT 53.785 18.260 54.455 19.540 ;
        RECT 53.615 17.580 54.735 18.260 ;
        RECT 40.155 12.770 41.015 13.610 ;
        RECT 50.755 12.170 51.165 14.790 ;
        RECT 51.465 13.590 52.005 16.820 ;
        RECT 57.705 16.770 59.635 19.550 ;
        RECT 57.125 15.920 59.835 16.770 ;
        RECT 61.215 15.380 61.475 20.200 ;
        RECT 60.685 14.650 61.575 15.380 ;
        RECT 61.975 14.790 62.365 36.300 ;
        RECT 62.705 16.820 63.205 37.620 ;
        RECT 65.235 38.470 65.515 40.460 ;
        RECT 67.805 40.390 68.905 41.160 ;
        RECT 76.505 40.450 76.805 42.180 ;
        RECT 65.785 39.630 66.165 40.230 ;
        RECT 65.815 39.010 66.065 39.630 ;
        RECT 65.685 38.630 66.165 39.010 ;
        RECT 65.235 33.400 65.565 38.470 ;
        RECT 66.115 37.610 66.415 38.470 ;
        RECT 67.195 37.610 67.495 38.470 ;
        RECT 68.105 38.430 68.385 40.390 ;
        RECT 71.405 38.820 71.675 38.990 ;
        RECT 71.015 38.510 71.675 38.820 ;
        RECT 66.115 33.370 67.495 37.610 ;
        RECT 68.045 38.380 68.385 38.430 ;
        RECT 70.965 38.400 71.675 38.510 ;
        RECT 64.515 32.150 64.835 32.170 ;
        RECT 66.195 32.150 67.325 33.370 ;
        RECT 68.045 33.360 68.375 38.380 ;
        RECT 70.965 37.030 71.195 38.400 ;
        RECT 71.405 38.150 71.675 38.400 ;
        RECT 72.305 38.770 72.595 39.010 ;
        RECT 73.715 38.770 74.405 38.790 ;
        RECT 72.305 38.330 74.405 38.770 ;
        RECT 72.305 38.140 72.595 38.330 ;
        RECT 71.675 37.590 72.295 37.950 ;
        RECT 73.715 37.620 74.405 38.330 ;
        RECT 70.895 36.430 71.275 37.030 ;
        RECT 71.685 36.720 72.115 37.590 ;
        RECT 70.965 35.240 71.195 36.430 ;
        RECT 71.685 36.300 73.565 36.720 ;
        RECT 71.685 35.770 72.115 36.300 ;
        RECT 71.535 35.410 72.155 35.770 ;
        RECT 70.965 35.230 71.445 35.240 ;
        RECT 70.965 34.550 71.525 35.230 ;
        RECT 71.055 34.400 71.525 34.550 ;
        RECT 71.255 33.450 71.525 34.400 ;
        RECT 72.165 34.150 72.435 35.150 ;
        RECT 72.165 33.420 72.675 34.150 ;
        RECT 72.165 33.330 72.665 33.420 ;
        RECT 67.525 32.780 68.055 33.160 ;
        RECT 64.515 31.100 67.345 32.150 ;
        RECT 67.625 31.900 67.885 32.780 ;
        RECT 67.605 31.280 67.965 31.900 ;
        RECT 72.415 31.210 72.665 33.330 ;
        RECT 64.515 30.190 64.835 31.100 ;
        RECT 66.195 31.090 67.325 31.100 ;
        RECT 68.225 30.810 72.865 31.210 ;
        RECT 72.415 30.530 72.665 30.810 ;
        RECT 64.515 30.130 64.845 30.190 ;
        RECT 64.525 20.200 64.845 30.130 ;
        RECT 65.845 28.880 66.115 30.240 ;
        RECT 66.975 28.880 67.245 30.200 ;
        RECT 72.285 30.100 72.665 30.530 ;
        RECT 72.285 29.590 72.645 30.100 ;
        RECT 65.845 22.190 67.245 28.880 ;
        RECT 65.845 20.190 66.115 22.190 ;
        RECT 66.975 20.150 67.245 22.190 ;
        RECT 72.295 21.750 72.555 29.590 ;
        RECT 72.295 20.200 72.675 21.750 ;
        RECT 64.815 19.540 65.865 19.950 ;
        RECT 67.225 19.550 72.275 19.930 ;
        RECT 64.985 18.260 65.655 19.540 ;
        RECT 64.815 17.580 65.935 18.260 ;
        RECT 51.445 12.750 52.305 13.590 ;
        RECT 27.865 11.130 30.415 11.950 ;
        RECT 28.395 11.090 30.415 11.130 ;
        RECT 39.115 10.980 41.565 11.990 ;
        RECT 50.335 10.970 52.355 12.170 ;
        RECT 61.975 12.160 62.385 14.790 ;
        RECT 62.685 13.590 63.225 16.820 ;
        RECT 68.905 16.770 70.835 19.550 ;
        RECT 68.325 15.920 71.035 16.770 ;
        RECT 72.415 15.380 72.675 20.200 ;
        RECT 71.885 14.650 72.775 15.380 ;
        RECT 73.175 14.790 73.565 36.300 ;
        RECT 73.905 16.820 74.405 37.620 ;
        RECT 76.525 38.460 76.805 40.450 ;
        RECT 79.095 40.380 80.195 41.150 ;
        RECT 87.745 40.470 88.045 42.200 ;
        RECT 77.075 39.620 77.455 40.220 ;
        RECT 77.105 39.000 77.355 39.620 ;
        RECT 76.975 38.620 77.455 39.000 ;
        RECT 76.525 33.390 76.855 38.460 ;
        RECT 77.405 37.600 77.705 38.460 ;
        RECT 78.485 37.600 78.785 38.460 ;
        RECT 79.395 38.420 79.675 40.380 ;
        RECT 82.695 38.810 82.965 38.980 ;
        RECT 82.305 38.500 82.965 38.810 ;
        RECT 77.405 33.360 78.785 37.600 ;
        RECT 79.335 38.370 79.675 38.420 ;
        RECT 82.255 38.390 82.965 38.500 ;
        RECT 75.805 32.140 76.125 32.160 ;
        RECT 77.485 32.140 78.615 33.360 ;
        RECT 79.335 33.350 79.665 38.370 ;
        RECT 82.255 37.020 82.485 38.390 ;
        RECT 82.695 38.140 82.965 38.390 ;
        RECT 83.595 38.760 83.885 39.000 ;
        RECT 85.005 38.760 85.695 38.780 ;
        RECT 83.595 38.320 85.695 38.760 ;
        RECT 83.595 38.130 83.885 38.320 ;
        RECT 82.965 37.580 83.585 37.940 ;
        RECT 85.005 37.610 85.695 38.320 ;
        RECT 82.185 36.420 82.565 37.020 ;
        RECT 82.975 36.710 83.405 37.580 ;
        RECT 82.255 35.230 82.485 36.420 ;
        RECT 82.975 36.290 84.855 36.710 ;
        RECT 82.975 35.760 83.405 36.290 ;
        RECT 82.825 35.400 83.445 35.760 ;
        RECT 82.255 35.220 82.735 35.230 ;
        RECT 82.255 34.540 82.815 35.220 ;
        RECT 82.345 34.390 82.815 34.540 ;
        RECT 82.545 33.440 82.815 34.390 ;
        RECT 83.455 34.140 83.725 35.140 ;
        RECT 83.455 33.410 83.965 34.140 ;
        RECT 83.455 33.320 83.955 33.410 ;
        RECT 78.815 32.770 79.345 33.150 ;
        RECT 75.805 31.090 78.635 32.140 ;
        RECT 78.915 31.890 79.175 32.770 ;
        RECT 78.895 31.270 79.255 31.890 ;
        RECT 83.705 31.200 83.955 33.320 ;
        RECT 75.805 30.180 76.125 31.090 ;
        RECT 77.485 31.080 78.615 31.090 ;
        RECT 79.515 30.800 84.155 31.200 ;
        RECT 83.705 30.520 83.955 30.800 ;
        RECT 75.805 30.120 76.135 30.180 ;
        RECT 75.815 20.190 76.135 30.120 ;
        RECT 77.135 28.870 77.405 30.230 ;
        RECT 78.265 28.870 78.535 30.190 ;
        RECT 83.575 30.090 83.955 30.520 ;
        RECT 83.575 29.580 83.935 30.090 ;
        RECT 77.135 22.180 78.535 28.870 ;
        RECT 77.135 20.180 77.405 22.180 ;
        RECT 78.265 20.140 78.535 22.180 ;
        RECT 83.585 21.740 83.845 29.580 ;
        RECT 83.585 20.190 83.965 21.740 ;
        RECT 76.105 19.530 77.155 19.940 ;
        RECT 78.515 19.540 83.565 19.920 ;
        RECT 76.275 18.250 76.945 19.530 ;
        RECT 76.105 17.570 77.225 18.250 ;
        RECT 62.665 12.750 63.525 13.590 ;
        RECT 73.175 12.190 73.585 14.790 ;
        RECT 73.885 13.590 74.425 16.820 ;
        RECT 80.195 16.760 82.125 19.540 ;
        RECT 79.615 15.910 82.325 16.760 ;
        RECT 83.705 15.370 83.965 20.190 ;
        RECT 83.175 14.640 84.065 15.370 ;
        RECT 84.465 14.780 84.855 36.290 ;
        RECT 85.195 16.810 85.695 37.610 ;
        RECT 87.765 38.480 88.045 40.470 ;
        RECT 90.335 40.400 91.435 41.170 ;
        RECT 98.955 40.490 99.255 42.220 ;
        RECT 88.315 39.640 88.695 40.240 ;
        RECT 88.345 39.020 88.595 39.640 ;
        RECT 88.215 38.640 88.695 39.020 ;
        RECT 87.765 33.410 88.095 38.480 ;
        RECT 88.645 37.620 88.945 38.480 ;
        RECT 89.725 37.620 90.025 38.480 ;
        RECT 90.635 38.440 90.915 40.400 ;
        RECT 93.935 38.830 94.205 39.000 ;
        RECT 93.545 38.520 94.205 38.830 ;
        RECT 88.645 33.380 90.025 37.620 ;
        RECT 90.575 38.390 90.915 38.440 ;
        RECT 93.495 38.410 94.205 38.520 ;
        RECT 87.045 32.160 87.365 32.180 ;
        RECT 88.725 32.160 89.855 33.380 ;
        RECT 90.575 33.370 90.905 38.390 ;
        RECT 93.495 37.040 93.725 38.410 ;
        RECT 93.935 38.160 94.205 38.410 ;
        RECT 94.835 38.780 95.125 39.020 ;
        RECT 96.245 38.780 96.935 38.800 ;
        RECT 94.835 38.340 96.935 38.780 ;
        RECT 94.835 38.150 95.125 38.340 ;
        RECT 94.205 37.600 94.825 37.960 ;
        RECT 96.245 37.630 96.935 38.340 ;
        RECT 93.425 36.440 93.805 37.040 ;
        RECT 94.215 36.730 94.645 37.600 ;
        RECT 93.495 35.250 93.725 36.440 ;
        RECT 94.215 36.310 96.095 36.730 ;
        RECT 94.215 35.780 94.645 36.310 ;
        RECT 94.065 35.420 94.685 35.780 ;
        RECT 93.495 35.240 93.975 35.250 ;
        RECT 93.495 34.560 94.055 35.240 ;
        RECT 93.585 34.410 94.055 34.560 ;
        RECT 93.785 33.460 94.055 34.410 ;
        RECT 94.695 34.160 94.965 35.160 ;
        RECT 94.695 33.430 95.205 34.160 ;
        RECT 94.695 33.340 95.195 33.430 ;
        RECT 90.055 32.790 90.585 33.170 ;
        RECT 87.045 31.110 89.875 32.160 ;
        RECT 90.155 31.910 90.415 32.790 ;
        RECT 90.135 31.290 90.495 31.910 ;
        RECT 94.945 31.220 95.195 33.340 ;
        RECT 87.045 30.200 87.365 31.110 ;
        RECT 88.725 31.100 89.855 31.110 ;
        RECT 90.755 30.820 95.395 31.220 ;
        RECT 94.945 30.540 95.195 30.820 ;
        RECT 87.045 30.140 87.375 30.200 ;
        RECT 87.055 20.210 87.375 30.140 ;
        RECT 88.375 28.890 88.645 30.250 ;
        RECT 89.505 28.890 89.775 30.210 ;
        RECT 94.815 30.110 95.195 30.540 ;
        RECT 94.815 29.600 95.175 30.110 ;
        RECT 88.375 22.200 89.775 28.890 ;
        RECT 88.375 20.200 88.645 22.200 ;
        RECT 89.505 20.160 89.775 22.200 ;
        RECT 94.825 21.760 95.085 29.600 ;
        RECT 94.825 20.210 95.205 21.760 ;
        RECT 87.345 19.550 88.395 19.960 ;
        RECT 89.755 19.560 94.805 19.940 ;
        RECT 87.515 18.270 88.185 19.550 ;
        RECT 87.345 17.590 88.465 18.270 ;
        RECT 73.865 12.750 74.725 13.590 ;
        RECT 61.415 10.960 63.435 12.160 ;
        RECT 72.725 10.990 74.745 12.190 ;
        RECT 84.465 12.180 84.875 14.780 ;
        RECT 85.175 13.580 85.715 16.810 ;
        RECT 91.435 16.780 93.365 19.560 ;
        RECT 90.855 15.930 93.565 16.780 ;
        RECT 94.945 15.390 95.205 20.210 ;
        RECT 94.415 14.660 95.305 15.390 ;
        RECT 95.705 14.800 96.095 36.310 ;
        RECT 96.435 16.830 96.935 37.630 ;
        RECT 98.975 38.500 99.255 40.490 ;
        RECT 101.545 40.420 102.645 41.190 ;
        RECT 110.155 40.530 110.455 42.260 ;
        RECT 99.525 39.660 99.905 40.260 ;
        RECT 99.555 39.040 99.805 39.660 ;
        RECT 99.425 38.660 99.905 39.040 ;
        RECT 98.975 33.430 99.305 38.500 ;
        RECT 99.855 37.640 100.155 38.500 ;
        RECT 100.935 37.640 101.235 38.500 ;
        RECT 101.845 38.460 102.125 40.420 ;
        RECT 105.145 38.850 105.415 39.020 ;
        RECT 104.755 38.540 105.415 38.850 ;
        RECT 99.855 33.400 101.235 37.640 ;
        RECT 101.785 38.410 102.125 38.460 ;
        RECT 104.705 38.430 105.415 38.540 ;
        RECT 98.255 32.180 98.575 32.200 ;
        RECT 99.935 32.180 101.065 33.400 ;
        RECT 101.785 33.390 102.115 38.410 ;
        RECT 104.705 37.060 104.935 38.430 ;
        RECT 105.145 38.180 105.415 38.430 ;
        RECT 106.045 38.800 106.335 39.040 ;
        RECT 107.455 38.800 108.145 38.820 ;
        RECT 106.045 38.360 108.145 38.800 ;
        RECT 106.045 38.170 106.335 38.360 ;
        RECT 105.415 37.620 106.035 37.980 ;
        RECT 107.455 37.650 108.145 38.360 ;
        RECT 104.635 36.460 105.015 37.060 ;
        RECT 105.425 36.750 105.855 37.620 ;
        RECT 104.705 35.270 104.935 36.460 ;
        RECT 105.425 36.330 107.305 36.750 ;
        RECT 105.425 35.800 105.855 36.330 ;
        RECT 105.275 35.440 105.895 35.800 ;
        RECT 104.705 35.260 105.185 35.270 ;
        RECT 104.705 34.580 105.265 35.260 ;
        RECT 104.795 34.430 105.265 34.580 ;
        RECT 104.995 33.480 105.265 34.430 ;
        RECT 105.905 34.180 106.175 35.180 ;
        RECT 105.905 33.450 106.415 34.180 ;
        RECT 105.905 33.360 106.405 33.450 ;
        RECT 101.265 32.810 101.795 33.190 ;
        RECT 98.255 31.130 101.085 32.180 ;
        RECT 101.365 31.930 101.625 32.810 ;
        RECT 101.345 31.310 101.705 31.930 ;
        RECT 106.155 31.240 106.405 33.360 ;
        RECT 98.255 30.220 98.575 31.130 ;
        RECT 99.935 31.120 101.065 31.130 ;
        RECT 101.965 30.840 106.605 31.240 ;
        RECT 106.155 30.560 106.405 30.840 ;
        RECT 98.255 30.160 98.585 30.220 ;
        RECT 98.265 20.230 98.585 30.160 ;
        RECT 99.585 28.910 99.855 30.270 ;
        RECT 100.715 28.910 100.985 30.230 ;
        RECT 106.025 30.130 106.405 30.560 ;
        RECT 106.025 29.620 106.385 30.130 ;
        RECT 99.585 22.220 100.985 28.910 ;
        RECT 99.585 20.220 99.855 22.220 ;
        RECT 100.715 20.180 100.985 22.220 ;
        RECT 106.035 21.780 106.295 29.620 ;
        RECT 106.035 20.230 106.415 21.780 ;
        RECT 98.555 19.570 99.605 19.980 ;
        RECT 100.965 19.580 106.015 19.960 ;
        RECT 98.725 18.290 99.395 19.570 ;
        RECT 98.555 17.610 99.675 18.290 ;
        RECT 85.155 12.740 86.015 13.580 ;
        RECT 95.705 12.180 96.115 14.800 ;
        RECT 96.415 13.600 96.955 16.830 ;
        RECT 102.645 16.800 104.575 19.580 ;
        RECT 102.065 15.950 104.775 16.800 ;
        RECT 106.155 15.410 106.415 20.230 ;
        RECT 105.625 14.680 106.515 15.410 ;
        RECT 106.915 14.820 107.305 36.330 ;
        RECT 107.645 16.850 108.145 37.650 ;
        RECT 110.175 38.540 110.455 40.530 ;
        RECT 112.745 40.460 113.845 41.230 ;
        RECT 121.365 40.550 121.665 42.280 ;
        RECT 142.880 42.020 144.100 43.390 ;
        RECT 110.725 39.700 111.105 40.300 ;
        RECT 110.755 39.080 111.005 39.700 ;
        RECT 110.625 38.700 111.105 39.080 ;
        RECT 110.175 33.470 110.505 38.540 ;
        RECT 111.055 37.680 111.355 38.540 ;
        RECT 112.135 37.680 112.435 38.540 ;
        RECT 113.045 38.500 113.325 40.460 ;
        RECT 116.345 38.890 116.615 39.060 ;
        RECT 115.955 38.580 116.615 38.890 ;
        RECT 111.055 33.440 112.435 37.680 ;
        RECT 112.985 38.450 113.325 38.500 ;
        RECT 115.905 38.470 116.615 38.580 ;
        RECT 109.455 32.220 109.775 32.240 ;
        RECT 111.135 32.220 112.265 33.440 ;
        RECT 112.985 33.430 113.315 38.450 ;
        RECT 115.905 37.100 116.135 38.470 ;
        RECT 116.345 38.220 116.615 38.470 ;
        RECT 117.245 38.840 117.535 39.080 ;
        RECT 118.655 38.840 119.345 38.860 ;
        RECT 117.245 38.400 119.345 38.840 ;
        RECT 117.245 38.210 117.535 38.400 ;
        RECT 116.615 37.660 117.235 38.020 ;
        RECT 118.655 37.690 119.345 38.400 ;
        RECT 115.835 36.500 116.215 37.100 ;
        RECT 116.625 36.790 117.055 37.660 ;
        RECT 115.905 35.310 116.135 36.500 ;
        RECT 116.625 36.370 118.505 36.790 ;
        RECT 116.625 35.840 117.055 36.370 ;
        RECT 116.475 35.480 117.095 35.840 ;
        RECT 115.905 35.300 116.385 35.310 ;
        RECT 115.905 34.620 116.465 35.300 ;
        RECT 115.995 34.470 116.465 34.620 ;
        RECT 116.195 33.520 116.465 34.470 ;
        RECT 117.105 34.220 117.375 35.220 ;
        RECT 117.105 33.490 117.615 34.220 ;
        RECT 117.105 33.400 117.605 33.490 ;
        RECT 112.465 32.850 112.995 33.230 ;
        RECT 109.455 31.170 112.285 32.220 ;
        RECT 112.565 31.970 112.825 32.850 ;
        RECT 112.545 31.350 112.905 31.970 ;
        RECT 117.355 31.280 117.605 33.400 ;
        RECT 109.455 30.260 109.775 31.170 ;
        RECT 111.135 31.160 112.265 31.170 ;
        RECT 113.165 30.880 117.805 31.280 ;
        RECT 117.355 30.600 117.605 30.880 ;
        RECT 109.455 30.200 109.785 30.260 ;
        RECT 109.465 20.270 109.785 30.200 ;
        RECT 110.785 28.950 111.055 30.310 ;
        RECT 111.915 28.950 112.185 30.270 ;
        RECT 117.225 30.170 117.605 30.600 ;
        RECT 117.225 29.660 117.585 30.170 ;
        RECT 110.785 22.260 112.185 28.950 ;
        RECT 110.785 20.260 111.055 22.260 ;
        RECT 111.915 20.220 112.185 22.260 ;
        RECT 117.235 21.820 117.495 29.660 ;
        RECT 117.235 20.270 117.615 21.820 ;
        RECT 109.755 19.610 110.805 20.020 ;
        RECT 112.165 19.620 117.215 20.000 ;
        RECT 109.925 18.330 110.595 19.610 ;
        RECT 109.755 17.650 110.875 18.330 ;
        RECT 96.395 12.760 97.255 13.600 ;
        RECT 106.915 12.230 107.325 14.820 ;
        RECT 107.625 13.620 108.165 16.850 ;
        RECT 113.845 16.840 115.775 19.620 ;
        RECT 113.265 15.990 115.975 16.840 ;
        RECT 117.355 15.450 117.615 20.270 ;
        RECT 116.825 14.720 117.715 15.450 ;
        RECT 118.115 14.860 118.505 36.370 ;
        RECT 118.845 16.890 119.345 37.690 ;
        RECT 121.385 38.560 121.665 40.550 ;
        RECT 123.955 40.480 125.055 41.250 ;
        RECT 121.935 39.720 122.315 40.320 ;
        RECT 121.965 39.100 122.215 39.720 ;
        RECT 121.835 38.720 122.315 39.100 ;
        RECT 121.385 33.490 121.715 38.560 ;
        RECT 122.265 37.700 122.565 38.560 ;
        RECT 123.345 37.700 123.645 38.560 ;
        RECT 124.255 38.520 124.535 40.480 ;
        RECT 127.555 38.910 127.825 39.080 ;
        RECT 127.165 38.600 127.825 38.910 ;
        RECT 122.265 33.460 123.645 37.700 ;
        RECT 124.195 38.470 124.535 38.520 ;
        RECT 127.115 38.490 127.825 38.600 ;
        RECT 120.665 32.240 120.985 32.260 ;
        RECT 122.345 32.240 123.475 33.460 ;
        RECT 124.195 33.450 124.525 38.470 ;
        RECT 127.115 37.120 127.345 38.490 ;
        RECT 127.555 38.240 127.825 38.490 ;
        RECT 128.455 38.860 128.745 39.100 ;
        RECT 142.940 38.950 144.100 42.020 ;
        RECT 129.865 38.860 130.555 38.880 ;
        RECT 128.455 38.420 130.555 38.860 ;
        RECT 128.455 38.230 128.745 38.420 ;
        RECT 127.825 37.680 128.445 38.040 ;
        RECT 129.865 37.710 130.555 38.420 ;
        RECT 127.045 36.520 127.425 37.120 ;
        RECT 127.835 36.810 128.265 37.680 ;
        RECT 127.115 35.330 127.345 36.520 ;
        RECT 127.835 36.390 129.715 36.810 ;
        RECT 127.835 35.860 128.265 36.390 ;
        RECT 127.685 35.500 128.305 35.860 ;
        RECT 127.115 35.320 127.595 35.330 ;
        RECT 127.115 34.640 127.675 35.320 ;
        RECT 127.205 34.490 127.675 34.640 ;
        RECT 127.405 33.540 127.675 34.490 ;
        RECT 128.315 34.240 128.585 35.240 ;
        RECT 128.315 33.510 128.825 34.240 ;
        RECT 128.315 33.420 128.815 33.510 ;
        RECT 123.675 32.870 124.205 33.250 ;
        RECT 120.665 31.190 123.495 32.240 ;
        RECT 123.775 31.990 124.035 32.870 ;
        RECT 123.755 31.370 124.115 31.990 ;
        RECT 128.565 31.300 128.815 33.420 ;
        RECT 120.665 30.280 120.985 31.190 ;
        RECT 122.345 31.180 123.475 31.190 ;
        RECT 124.375 30.900 129.015 31.300 ;
        RECT 128.565 30.620 128.815 30.900 ;
        RECT 120.665 30.220 120.995 30.280 ;
        RECT 120.675 20.290 120.995 30.220 ;
        RECT 121.995 28.970 122.265 30.330 ;
        RECT 123.125 28.970 123.395 30.290 ;
        RECT 128.435 30.190 128.815 30.620 ;
        RECT 128.435 29.680 128.795 30.190 ;
        RECT 121.995 22.280 123.395 28.970 ;
        RECT 121.995 20.280 122.265 22.280 ;
        RECT 123.125 20.240 123.395 22.280 ;
        RECT 128.445 21.840 128.705 29.680 ;
        RECT 128.445 20.290 128.825 21.840 ;
        RECT 120.965 19.630 122.015 20.040 ;
        RECT 123.375 19.640 128.425 20.020 ;
        RECT 121.135 18.350 121.805 19.630 ;
        RECT 120.965 17.670 122.085 18.350 ;
        RECT 107.605 12.780 108.465 13.620 ;
        RECT 118.115 12.230 118.525 14.860 ;
        RECT 118.825 13.660 119.365 16.890 ;
        RECT 125.055 16.860 126.985 19.640 ;
        RECT 124.475 16.010 127.185 16.860 ;
        RECT 128.565 15.470 128.825 20.290 ;
        RECT 128.035 14.740 128.925 15.470 ;
        RECT 129.325 14.880 129.715 36.390 ;
        RECT 130.055 16.910 130.555 37.710 ;
        RECT 142.900 37.580 144.120 38.950 ;
        RECT 132.395 24.340 132.705 30.230 ;
        RECT 132.195 20.120 132.705 24.340 ;
        RECT 118.805 12.820 119.665 13.660 ;
        RECT 129.325 12.260 129.735 14.880 ;
        RECT 130.035 13.680 130.575 16.910 ;
        RECT 132.195 15.510 132.505 20.120 ;
        RECT 137.715 19.980 138.005 30.170 ;
        RECT 132.685 19.590 138.005 19.980 ;
        RECT 137.715 16.940 138.005 19.590 ;
        RECT 142.940 17.940 144.090 19.160 ;
        RECT 145.080 18.760 146.200 18.930 ;
        RECT 137.395 15.890 138.295 16.940 ;
        RECT 137.715 15.720 138.005 15.890 ;
        RECT 131.975 14.270 132.735 15.510 ;
        RECT 142.940 15.090 144.050 17.940 ;
        RECT 142.900 13.870 144.050 15.090 ;
        RECT 145.070 14.920 146.200 18.760 ;
        RECT 145.030 13.970 146.200 14.920 ;
        RECT 145.030 13.900 146.150 13.970 ;
        RECT 130.015 12.840 130.875 13.680 ;
        RECT 83.845 10.980 85.865 12.180 ;
        RECT 95.145 10.980 97.165 12.180 ;
        RECT 106.335 11.030 108.355 12.230 ;
        RECT 117.565 11.030 119.585 12.230 ;
        RECT 128.865 11.060 130.885 12.260 ;
        RECT 74.340 0.110 75.630 1.460 ;
        RECT 93.550 0.180 94.840 1.530 ;
        RECT 112.950 0.310 114.240 1.660 ;
        RECT 131.850 0.380 133.490 1.930 ;
        RECT 151.650 0.250 152.920 1.470 ;
      LAYER met3 ;
        RECT 135.340 223.855 136.790 225.205 ;
        RECT 138.130 223.785 139.580 225.135 ;
        RECT 143.180 223.815 144.630 225.165 ;
        RECT 32.460 203.865 34.440 204.195 ;
        RECT 62.460 203.865 64.440 204.195 ;
        RECT 92.460 203.865 94.440 204.195 ;
        RECT 17.460 201.145 19.440 201.475 ;
        RECT 47.460 201.145 49.440 201.475 ;
        RECT 77.460 201.145 79.440 201.475 ;
        RECT 107.460 201.145 109.440 201.475 ;
        RECT 32.460 198.425 34.440 198.755 ;
        RECT 62.460 198.425 64.440 198.755 ;
        RECT 92.460 198.425 94.440 198.755 ;
        RECT 17.460 195.705 19.440 196.035 ;
        RECT 47.460 195.705 49.440 196.035 ;
        RECT 77.460 195.705 79.440 196.035 ;
        RECT 107.460 195.705 109.440 196.035 ;
        RECT 32.460 192.985 34.440 193.315 ;
        RECT 62.460 192.985 64.440 193.315 ;
        RECT 92.460 192.985 94.440 193.315 ;
        RECT 17.460 190.265 19.440 190.595 ;
        RECT 47.460 190.265 49.440 190.595 ;
        RECT 77.460 190.265 79.440 190.595 ;
        RECT 107.460 190.265 109.440 190.595 ;
        RECT 32.460 187.545 34.440 187.875 ;
        RECT 62.460 187.545 64.440 187.875 ;
        RECT 92.460 187.545 94.440 187.875 ;
        RECT 76.255 186.840 76.585 186.855 ;
        RECT 87.295 186.840 87.625 186.855 ;
        RECT 76.255 186.540 87.625 186.840 ;
        RECT 76.255 186.525 76.585 186.540 ;
        RECT 87.295 186.525 87.625 186.540 ;
        RECT 17.460 184.825 19.440 185.155 ;
        RECT 47.460 184.825 49.440 185.155 ;
        RECT 77.460 184.825 79.440 185.155 ;
        RECT 107.460 184.825 109.440 185.155 ;
        RECT 32.460 182.105 34.440 182.435 ;
        RECT 62.460 182.105 64.440 182.435 ;
        RECT 92.460 182.105 94.440 182.435 ;
        RECT 63.835 180.720 64.165 180.735 ;
        RECT 65.880 180.720 66.260 180.730 ;
        RECT 63.835 180.420 66.260 180.720 ;
        RECT 63.835 180.405 64.165 180.420 ;
        RECT 65.880 180.410 66.260 180.420 ;
        RECT 17.460 179.385 19.440 179.715 ;
        RECT 47.460 179.385 49.440 179.715 ;
        RECT 77.460 179.385 79.440 179.715 ;
        RECT 107.460 179.385 109.440 179.715 ;
        RECT 90.975 179.360 91.305 179.375 ;
        RECT 94.655 179.360 94.985 179.375 ;
        RECT 90.975 179.060 94.985 179.360 ;
        RECT 90.975 179.045 91.305 179.060 ;
        RECT 94.655 179.045 94.985 179.060 ;
        RECT 57.395 178.680 57.725 178.695 ;
        RECT 60.155 178.680 60.485 178.695 ;
        RECT 84.535 178.680 84.865 178.695 ;
        RECT 57.395 178.380 84.865 178.680 ;
        RECT 57.395 178.365 57.725 178.380 ;
        RECT 60.155 178.365 60.485 178.380 ;
        RECT 84.535 178.365 84.865 178.380 ;
        RECT 91.895 178.680 92.225 178.695 ;
        RECT 96.955 178.680 97.285 178.695 ;
        RECT 91.895 178.380 97.285 178.680 ;
        RECT 91.895 178.365 92.225 178.380 ;
        RECT 96.955 178.365 97.285 178.380 ;
        RECT 80.395 178.000 80.725 178.015 ;
        RECT 90.055 178.000 90.385 178.015 ;
        RECT 95.115 178.000 95.445 178.015 ;
        RECT 104.315 178.000 104.645 178.015 ;
        RECT 80.395 177.700 104.645 178.000 ;
        RECT 80.395 177.685 80.725 177.700 ;
        RECT 90.055 177.685 90.385 177.700 ;
        RECT 95.115 177.685 95.445 177.700 ;
        RECT 104.315 177.685 104.645 177.700 ;
        RECT 40.835 177.330 41.165 177.335 ;
        RECT 40.835 177.320 41.420 177.330 ;
        RECT 40.610 177.020 41.420 177.320 ;
        RECT 40.835 177.010 41.420 177.020 ;
        RECT 40.835 177.005 41.165 177.010 ;
        RECT 32.460 176.665 34.440 176.995 ;
        RECT 62.460 176.665 64.440 176.995 ;
        RECT 92.460 176.665 94.440 176.995 ;
        RECT 25.195 175.960 25.525 175.975 ;
        RECT 37.155 175.960 37.485 175.975 ;
        RECT 25.195 175.660 37.485 175.960 ;
        RECT 25.195 175.645 25.525 175.660 ;
        RECT 37.155 175.645 37.485 175.660 ;
        RECT 41.960 174.600 42.340 174.610 ;
        RECT 44.975 174.600 45.305 174.615 ;
        RECT 41.960 174.300 45.305 174.600 ;
        RECT 41.960 174.290 42.340 174.300 ;
        RECT 44.975 174.285 45.305 174.300 ;
        RECT 67.055 174.600 67.385 174.615 ;
        RECT 70.735 174.610 71.065 174.615 ;
        RECT 67.720 174.600 68.100 174.610 ;
        RECT 67.055 174.300 68.100 174.600 ;
        RECT 67.055 174.285 67.385 174.300 ;
        RECT 67.720 174.290 68.100 174.300 ;
        RECT 70.480 174.600 71.065 174.610 ;
        RECT 70.480 174.300 71.290 174.600 ;
        RECT 70.480 174.290 71.065 174.300 ;
        RECT 70.735 174.285 71.065 174.290 ;
        RECT 17.460 173.945 19.440 174.275 ;
        RECT 47.460 173.945 49.440 174.275 ;
        RECT 77.460 173.945 79.440 174.275 ;
        RECT 107.460 173.945 109.440 174.275 ;
        RECT 133.700 172.500 134.930 172.705 ;
        RECT 32.460 171.225 34.440 171.555 ;
        RECT 62.460 171.225 64.440 171.555 ;
        RECT 92.460 171.225 94.440 171.555 ;
        RECT 129.030 170.130 134.930 172.500 ;
        RECT 133.700 170.095 134.930 170.130 ;
        RECT 28.875 169.840 29.205 169.855 ;
        RECT 33.935 169.840 34.265 169.855 ;
        RECT 28.875 169.540 34.265 169.840 ;
        RECT 28.875 169.525 29.205 169.540 ;
        RECT 33.935 169.525 34.265 169.540 ;
        RECT 113.515 169.840 113.845 169.855 ;
        RECT 116.970 169.840 118.970 169.990 ;
        RECT 113.515 169.540 118.970 169.840 ;
        RECT 113.515 169.525 113.845 169.540 ;
        RECT 116.970 169.390 118.970 169.540 ;
        RECT 30.255 169.160 30.585 169.175 ;
        RECT 37.615 169.160 37.945 169.175 ;
        RECT 30.255 168.860 37.945 169.160 ;
        RECT 30.255 168.845 30.585 168.860 ;
        RECT 37.615 168.845 37.945 168.860 ;
        RECT 17.460 168.505 19.440 168.835 ;
        RECT 47.460 168.505 49.440 168.835 ;
        RECT 77.460 168.505 79.440 168.835 ;
        RECT 107.460 168.505 109.440 168.835 ;
        RECT 42.880 167.120 43.260 167.130 ;
        RECT 44.515 167.120 44.845 167.135 ;
        RECT 42.880 166.820 44.845 167.120 ;
        RECT 42.880 166.810 43.260 166.820 ;
        RECT 38.995 166.440 39.325 166.455 ;
        RECT 42.920 166.440 43.220 166.810 ;
        RECT 44.515 166.805 44.845 166.820 ;
        RECT 92.355 166.760 92.685 166.775 ;
        RECT 38.995 166.140 43.220 166.440 ;
        RECT 91.680 166.460 92.685 166.760 ;
        RECT 38.995 166.125 39.325 166.140 ;
        RECT 32.460 165.785 34.440 166.115 ;
        RECT 62.460 165.785 64.440 166.115 ;
        RECT 91.680 164.415 91.980 166.460 ;
        RECT 92.355 166.445 92.685 166.460 ;
        RECT 92.460 165.785 94.440 166.115 ;
        RECT 91.435 164.100 91.980 164.415 ;
        RECT 91.435 164.085 91.765 164.100 ;
        RECT 17.460 163.065 19.440 163.395 ;
        RECT 47.460 163.065 49.440 163.395 ;
        RECT 77.460 163.065 79.440 163.395 ;
        RECT 107.460 163.065 109.440 163.395 ;
        RECT 65.675 161.000 66.005 161.015 ;
        RECT 68.895 161.000 69.225 161.015 ;
        RECT 65.675 160.700 69.225 161.000 ;
        RECT 65.675 160.685 66.005 160.700 ;
        RECT 68.895 160.685 69.225 160.700 ;
        RECT 32.460 160.345 34.440 160.675 ;
        RECT 62.460 160.345 64.440 160.675 ;
        RECT 92.460 160.345 94.440 160.675 ;
        RECT 66.135 160.320 66.465 160.335 ;
        RECT 69.815 160.320 70.145 160.335 ;
        RECT 66.135 160.020 70.145 160.320 ;
        RECT 66.135 160.005 66.465 160.020 ;
        RECT 69.815 160.005 70.145 160.020 ;
        RECT 61.535 159.640 61.865 159.655 ;
        RECT 70.275 159.640 70.605 159.655 ;
        RECT 61.535 159.340 70.605 159.640 ;
        RECT 61.535 159.325 61.865 159.340 ;
        RECT 70.275 159.325 70.605 159.340 ;
        RECT 81.775 158.970 82.105 158.975 ;
        RECT 81.520 158.960 82.105 158.970 ;
        RECT 81.520 158.660 82.330 158.960 ;
        RECT 81.520 158.650 82.105 158.660 ;
        RECT 81.775 158.645 82.105 158.650 ;
        RECT 17.460 157.625 19.440 157.955 ;
        RECT 47.460 157.625 49.440 157.955 ;
        RECT 77.460 157.625 79.440 157.955 ;
        RECT 107.460 157.625 109.440 157.955 ;
        RECT 43.135 156.920 43.465 156.935 ;
        RECT 67.055 156.920 67.385 156.935 ;
        RECT 43.135 156.620 67.385 156.920 ;
        RECT 43.135 156.605 43.465 156.620 ;
        RECT 67.055 156.605 67.385 156.620 ;
        RECT 89.595 156.920 89.925 156.935 ;
        RECT 96.955 156.920 97.285 156.935 ;
        RECT 89.595 156.620 97.285 156.920 ;
        RECT 89.595 156.605 89.925 156.620 ;
        RECT 96.955 156.605 97.285 156.620 ;
        RECT 64.295 156.240 64.625 156.255 ;
        RECT 66.135 156.240 66.465 156.255 ;
        RECT 64.295 155.940 66.465 156.240 ;
        RECT 64.295 155.925 64.625 155.940 ;
        RECT 66.135 155.925 66.465 155.940 ;
        RECT 85.455 156.240 85.785 156.255 ;
        RECT 91.895 156.240 92.225 156.255 ;
        RECT 85.455 155.940 92.225 156.240 ;
        RECT 85.455 155.925 85.785 155.940 ;
        RECT 91.895 155.925 92.225 155.940 ;
        RECT 93.275 156.240 93.605 156.255 ;
        RECT 95.320 156.240 95.700 156.250 ;
        RECT 93.275 155.940 95.700 156.240 ;
        RECT 93.275 155.925 93.605 155.940 ;
        RECT 95.320 155.930 95.700 155.940 ;
        RECT 32.460 154.905 34.440 155.235 ;
        RECT 62.460 154.905 64.440 155.235 ;
        RECT 92.460 154.905 94.440 155.235 ;
        RECT 36.695 154.880 37.025 154.895 ;
        RECT 41.755 154.880 42.085 154.895 ;
        RECT 36.695 154.580 42.085 154.880 ;
        RECT 36.695 154.565 37.025 154.580 ;
        RECT 41.755 154.565 42.085 154.580 ;
        RECT 32.555 154.200 32.885 154.215 ;
        RECT 37.615 154.200 37.945 154.215 ;
        RECT 32.555 153.900 37.945 154.200 ;
        RECT 32.555 153.885 32.885 153.900 ;
        RECT 37.615 153.885 37.945 153.900 ;
        RECT 59.235 154.200 59.565 154.215 ;
        RECT 65.215 154.200 65.545 154.215 ;
        RECT 59.235 153.900 65.545 154.200 ;
        RECT 59.235 153.885 59.565 153.900 ;
        RECT 65.215 153.885 65.545 153.900 ;
        RECT 29.795 153.520 30.125 153.535 ;
        RECT 61.995 153.520 62.325 153.535 ;
        RECT 29.795 153.220 62.325 153.520 ;
        RECT 29.795 153.205 30.125 153.220 ;
        RECT 61.995 153.205 62.325 153.220 ;
        RECT 17.460 152.185 19.440 152.515 ;
        RECT 47.460 152.185 49.440 152.515 ;
        RECT 77.460 152.185 79.440 152.515 ;
        RECT 107.460 152.185 109.440 152.515 ;
        RECT 52.335 151.480 52.665 151.495 ;
        RECT 81.520 151.480 81.900 151.490 ;
        RECT 52.335 151.180 81.900 151.480 ;
        RECT 52.335 151.165 52.665 151.180 ;
        RECT 81.520 151.170 81.900 151.180 ;
        RECT 76.715 150.800 77.045 150.815 ;
        RECT 96.955 150.800 97.285 150.815 ;
        RECT 98.335 150.800 98.665 150.815 ;
        RECT 76.715 150.500 98.665 150.800 ;
        RECT 76.715 150.485 77.045 150.500 ;
        RECT 96.955 150.485 97.285 150.500 ;
        RECT 98.335 150.485 98.665 150.500 ;
        RECT 42.880 150.120 43.260 150.130 ;
        RECT 52.335 150.120 52.665 150.135 ;
        RECT 42.880 149.820 52.665 150.120 ;
        RECT 42.880 149.810 43.260 149.820 ;
        RECT 52.335 149.805 52.665 149.820 ;
        RECT 68.895 150.120 69.225 150.135 ;
        RECT 71.400 150.120 71.780 150.130 ;
        RECT 68.895 149.820 71.780 150.120 ;
        RECT 68.895 149.805 69.225 149.820 ;
        RECT 71.400 149.810 71.780 149.820 ;
        RECT 32.460 149.465 34.440 149.795 ;
        RECT 62.460 149.465 64.440 149.795 ;
        RECT 92.460 149.465 94.440 149.795 ;
        RECT 61.075 148.080 61.405 148.095 ;
        RECT 98.080 148.080 98.460 148.090 ;
        RECT 61.075 147.780 98.460 148.080 ;
        RECT 61.075 147.765 61.405 147.780 ;
        RECT 98.080 147.770 98.460 147.780 ;
        RECT 17.460 146.745 19.440 147.075 ;
        RECT 47.460 146.745 49.440 147.075 ;
        RECT 77.460 146.745 79.440 147.075 ;
        RECT 107.460 146.745 109.440 147.075 ;
        RECT 70.735 146.050 71.065 146.055 ;
        RECT 70.480 146.040 71.065 146.050 ;
        RECT 70.280 145.740 71.065 146.040 ;
        RECT 70.480 145.730 71.065 145.740 ;
        RECT 70.735 145.725 71.065 145.730 ;
        RECT 32.460 144.025 34.440 144.355 ;
        RECT 62.460 144.025 64.440 144.355 ;
        RECT 92.460 144.025 94.440 144.355 ;
        RECT 87.295 143.320 87.625 143.335 ;
        RECT 99.715 143.320 100.045 143.335 ;
        RECT 87.295 143.020 100.045 143.320 ;
        RECT 87.295 143.005 87.625 143.020 ;
        RECT 99.715 143.005 100.045 143.020 ;
        RECT 42.675 142.640 43.005 142.655 ;
        RECT 51.415 142.640 51.745 142.655 ;
        RECT 42.675 142.340 51.745 142.640 ;
        RECT 42.675 142.325 43.005 142.340 ;
        RECT 51.415 142.325 51.745 142.340 ;
        RECT 86.835 142.640 87.165 142.655 ;
        RECT 90.515 142.640 90.845 142.655 ;
        RECT 86.835 142.340 90.845 142.640 ;
        RECT 86.835 142.325 87.165 142.340 ;
        RECT 90.515 142.325 90.845 142.340 ;
        RECT 17.460 141.305 19.440 141.635 ;
        RECT 47.460 141.305 49.440 141.635 ;
        RECT 77.460 141.305 79.440 141.635 ;
        RECT 107.460 141.305 109.440 141.635 ;
        RECT 98.080 139.920 98.460 139.930 ;
        RECT 116.970 139.920 118.970 140.070 ;
        RECT 98.080 139.620 118.970 139.920 ;
        RECT 98.080 139.610 98.460 139.620 ;
        RECT 116.970 139.470 118.970 139.620 ;
        RECT 32.460 138.585 34.440 138.915 ;
        RECT 62.460 138.585 64.440 138.915 ;
        RECT 92.460 138.585 94.440 138.915 ;
        RECT 40.835 138.570 41.165 138.575 ;
        RECT 42.675 138.570 43.005 138.575 ;
        RECT 40.835 138.560 41.420 138.570 ;
        RECT 42.675 138.560 43.260 138.570 ;
        RECT 67.720 138.560 68.100 138.570 ;
        RECT 68.435 138.560 68.765 138.575 ;
        RECT 40.835 138.260 41.620 138.560 ;
        RECT 42.675 138.260 43.460 138.560 ;
        RECT 67.720 138.260 68.765 138.560 ;
        RECT 40.835 138.250 41.420 138.260 ;
        RECT 42.675 138.250 43.260 138.260 ;
        RECT 67.720 138.250 68.100 138.260 ;
        RECT 40.835 138.245 41.165 138.250 ;
        RECT 42.675 138.245 43.005 138.250 ;
        RECT 68.435 138.245 68.765 138.260 ;
        RECT 132.510 138.165 135.210 140.035 ;
        RECT 38.075 137.880 38.405 137.895 ;
        RECT 41.960 137.880 42.340 137.890 ;
        RECT 38.075 137.580 42.340 137.880 ;
        RECT 38.075 137.565 38.405 137.580 ;
        RECT 41.960 137.570 42.340 137.580 ;
        RECT 93.735 137.880 94.065 137.895 ;
        RECT 95.320 137.880 95.700 137.890 ;
        RECT 93.735 137.580 95.700 137.880 ;
        RECT 93.735 137.565 94.065 137.580 ;
        RECT 95.320 137.570 95.700 137.580 ;
        RECT 17.460 135.865 19.440 136.195 ;
        RECT 47.460 135.865 49.440 136.195 ;
        RECT 77.460 135.865 79.440 136.195 ;
        RECT 107.460 135.865 109.440 136.195 ;
        RECT 64.295 135.160 64.625 135.175 ;
        RECT 65.880 135.160 66.260 135.170 ;
        RECT 64.295 134.860 66.260 135.160 ;
        RECT 64.295 134.845 64.625 134.860 ;
        RECT 65.880 134.850 66.260 134.860 ;
        RECT 79.015 135.160 79.345 135.175 ;
        RECT 81.520 135.160 81.900 135.170 ;
        RECT 84.995 135.160 85.325 135.175 ;
        RECT 79.015 134.860 85.325 135.160 ;
        RECT 79.015 134.845 79.345 134.860 ;
        RECT 81.520 134.850 81.900 134.860 ;
        RECT 84.995 134.845 85.325 134.860 ;
        RECT 32.460 133.145 34.440 133.475 ;
        RECT 62.460 133.145 64.440 133.475 ;
        RECT 92.460 133.145 94.440 133.475 ;
        RECT 17.460 130.425 19.440 130.755 ;
        RECT 47.460 130.425 49.440 130.755 ;
        RECT 77.460 130.425 79.440 130.755 ;
        RECT 107.460 130.425 109.440 130.755 ;
        RECT 32.460 127.705 34.440 128.035 ;
        RECT 62.460 127.705 64.440 128.035 ;
        RECT 92.460 127.705 94.440 128.035 ;
        RECT 17.460 124.985 19.440 125.315 ;
        RECT 47.460 124.985 49.440 125.315 ;
        RECT 77.460 124.985 79.440 125.315 ;
        RECT 107.460 124.985 109.440 125.315 ;
        RECT 32.460 122.265 34.440 122.595 ;
        RECT 62.460 122.265 64.440 122.595 ;
        RECT 92.460 122.265 94.440 122.595 ;
        RECT 17.460 119.545 19.440 119.875 ;
        RECT 47.460 119.545 49.440 119.875 ;
        RECT 77.460 119.545 79.440 119.875 ;
        RECT 107.460 119.545 109.440 119.875 ;
        RECT 32.460 116.825 34.440 117.155 ;
        RECT 62.460 116.825 64.440 117.155 ;
        RECT 92.460 116.825 94.440 117.155 ;
        RECT 17.460 114.105 19.440 114.435 ;
        RECT 47.460 114.105 49.440 114.435 ;
        RECT 77.460 114.105 79.440 114.435 ;
        RECT 107.460 114.105 109.440 114.435 ;
        RECT 32.460 111.385 34.440 111.715 ;
        RECT 62.460 111.385 64.440 111.715 ;
        RECT 92.460 111.385 94.440 111.715 ;
        RECT 71.400 111.360 71.780 111.370 ;
        RECT 72.115 111.360 72.445 111.375 ;
        RECT 71.400 111.060 72.445 111.360 ;
        RECT 71.400 111.050 71.780 111.060 ;
        RECT 72.115 111.045 72.445 111.060 ;
        RECT 116.970 110.015 118.970 110.150 ;
        RECT 116.735 109.685 118.970 110.015 ;
        RECT 116.970 109.550 118.970 109.685 ;
        RECT 17.460 108.665 19.440 108.995 ;
        RECT 47.460 108.665 49.440 108.995 ;
        RECT 77.460 108.665 79.440 108.995 ;
        RECT 107.460 108.665 109.440 108.995 ;
        RECT 32.460 105.945 34.440 106.275 ;
        RECT 62.460 105.945 64.440 106.275 ;
        RECT 92.460 105.945 94.440 106.275 ;
        RECT 129.700 105.605 133.210 106.625 ;
        RECT 37.630 88.620 38.970 88.755 ;
        RECT 13.950 87.980 14.980 88.515 ;
        RECT 13.950 87.500 14.990 87.980 ;
        RECT 13.950 87.175 14.980 87.500 ;
        RECT 14.070 86.570 14.810 87.175 ;
        RECT 20.050 87.105 20.920 88.515 ;
        RECT 14.070 75.715 14.700 86.570 ;
        RECT 20.170 77.115 20.800 87.105 ;
        RECT 25.910 87.055 26.860 88.515 ;
        RECT 26.070 78.385 26.700 87.055 ;
        RECT 31.730 86.965 32.910 88.585 ;
        RECT 32.005 79.615 32.635 86.965 ;
        RECT 37.630 86.835 39.120 88.620 ;
        RECT 38.060 81.125 38.690 86.835 ;
        RECT 43.790 86.745 45.190 88.605 ;
        RECT 49.710 86.945 51.060 88.615 ;
        RECT 44.175 82.625 44.805 86.745 ;
        RECT 50.070 83.875 50.700 86.945 ;
        RECT 55.530 86.785 56.750 88.545 ;
        RECT 55.825 85.115 56.455 86.785 ;
        RECT 61.670 86.625 63.180 88.615 ;
        RECT 67.680 88.305 68.720 89.815 ;
        RECT 67.885 87.225 68.515 88.305 ;
        RECT 62.110 86.175 62.740 86.625 ;
        RECT 67.885 86.595 130.605 87.225 ;
        RECT 62.110 85.545 118.855 86.175 ;
        RECT 55.825 84.485 107.605 85.115 ;
        RECT 50.070 83.245 96.285 83.875 ;
        RECT 44.175 81.995 85.055 82.625 ;
        RECT 38.060 80.495 73.765 81.125 ;
        RECT 32.005 78.985 62.635 79.615 ;
        RECT 26.070 77.755 51.245 78.385 ;
        RECT 20.170 76.485 40.645 77.115 ;
        RECT 14.070 75.660 29.295 75.715 ;
        RECT 40.015 75.710 40.645 76.485 ;
        RECT 14.070 75.085 30.410 75.660 ;
        RECT 27.850 74.670 30.410 75.085 ;
        RECT 3.910 71.345 6.100 73.215 ;
        RECT 27.850 73.120 30.450 74.670 ;
        RECT 39.060 74.510 41.620 75.710 ;
        RECT 50.615 75.580 51.245 77.755 ;
        RECT 62.005 75.690 62.635 78.985 ;
        RECT 49.930 74.650 52.490 75.580 ;
        RECT 0.970 70.330 3.070 70.430 ;
        RECT 15.510 70.330 17.040 71.185 ;
        RECT 0.960 68.750 17.040 70.330 ;
        RECT 0.970 68.710 3.070 68.750 ;
        RECT 15.510 68.635 17.040 68.750 ;
        RECT 20.145 54.060 20.605 54.135 ;
        RECT 25.715 54.060 26.175 54.085 ;
        RECT 20.145 53.620 26.175 54.060 ;
        RECT 20.145 53.565 20.605 53.620 ;
        RECT 25.715 53.515 26.175 53.620 ;
        RECT 22.405 48.870 22.885 48.935 ;
        RECT 22.405 48.550 24.205 48.870 ;
        RECT 22.405 48.385 22.885 48.550 ;
        RECT 23.635 45.710 24.195 48.550 ;
        RECT 27.515 45.710 27.995 45.735 ;
        RECT 23.635 45.290 27.995 45.710 ;
        RECT 23.635 45.280 24.195 45.290 ;
        RECT 27.515 45.185 27.995 45.290 ;
        RECT 20.745 40.120 21.225 40.225 ;
        RECT 24.545 40.120 25.105 40.130 ;
        RECT 20.745 39.700 25.105 40.120 ;
        RECT 20.745 39.675 21.225 39.700 ;
        RECT 24.545 36.860 25.105 39.700 ;
        RECT 25.855 36.860 26.335 37.025 ;
        RECT 24.535 36.540 26.335 36.860 ;
        RECT 25.855 36.475 26.335 36.540 ;
        RECT 22.565 31.790 23.025 31.895 ;
        RECT 28.135 31.790 28.595 31.845 ;
        RECT 22.565 31.350 28.595 31.790 ;
        RECT 22.565 31.325 23.025 31.350 ;
        RECT 28.135 31.275 28.595 31.350 ;
        RECT 29.765 12.265 30.255 73.120 ;
        RECT 38.960 73.080 41.730 74.510 ;
        RECT 31.345 54.070 31.805 54.145 ;
        RECT 36.915 54.070 37.375 54.095 ;
        RECT 31.345 53.630 37.375 54.070 ;
        RECT 31.345 53.575 31.805 53.630 ;
        RECT 36.915 53.525 37.375 53.630 ;
        RECT 33.605 48.880 34.085 48.945 ;
        RECT 33.605 48.560 35.405 48.880 ;
        RECT 33.605 48.395 34.085 48.560 ;
        RECT 34.835 45.720 35.395 48.560 ;
        RECT 38.715 45.720 39.195 45.745 ;
        RECT 34.835 45.300 39.195 45.720 ;
        RECT 34.835 45.290 35.395 45.300 ;
        RECT 38.715 45.195 39.195 45.300 ;
        RECT 32.025 40.120 32.505 40.225 ;
        RECT 35.825 40.120 36.385 40.130 ;
        RECT 32.025 39.700 36.385 40.120 ;
        RECT 32.025 39.675 32.505 39.700 ;
        RECT 35.825 36.860 36.385 39.700 ;
        RECT 37.135 36.860 37.615 37.025 ;
        RECT 35.815 36.540 37.615 36.860 ;
        RECT 37.135 36.475 37.615 36.540 ;
        RECT 33.845 31.790 34.305 31.895 ;
        RECT 39.415 31.790 39.875 31.845 ;
        RECT 33.845 31.350 39.875 31.790 ;
        RECT 33.845 31.325 34.305 31.350 ;
        RECT 39.415 31.275 39.875 31.350 ;
        RECT 41.055 12.360 41.545 73.080 ;
        RECT 49.930 73.030 52.530 74.650 ;
        RECT 61.330 74.530 63.890 75.690 ;
        RECT 73.135 75.580 73.765 80.495 ;
        RECT 84.425 75.690 85.055 81.995 ;
        RECT 72.340 74.980 74.900 75.580 ;
        RECT 42.565 54.040 43.025 54.115 ;
        RECT 48.135 54.040 48.595 54.065 ;
        RECT 42.565 53.600 48.595 54.040 ;
        RECT 42.565 53.545 43.025 53.600 ;
        RECT 48.135 53.495 48.595 53.600 ;
        RECT 44.825 48.850 45.305 48.915 ;
        RECT 44.825 48.530 46.625 48.850 ;
        RECT 44.825 48.365 45.305 48.530 ;
        RECT 46.055 45.690 46.615 48.530 ;
        RECT 49.935 45.690 50.415 45.715 ;
        RECT 46.055 45.270 50.415 45.690 ;
        RECT 46.055 45.260 46.615 45.270 ;
        RECT 49.935 45.165 50.415 45.270 ;
        RECT 43.315 40.100 43.795 40.205 ;
        RECT 47.115 40.100 47.675 40.110 ;
        RECT 43.315 39.680 47.675 40.100 ;
        RECT 43.315 39.655 43.795 39.680 ;
        RECT 47.115 36.840 47.675 39.680 ;
        RECT 48.425 36.840 48.905 37.005 ;
        RECT 47.105 36.520 48.905 36.840 ;
        RECT 48.425 36.455 48.905 36.520 ;
        RECT 45.135 31.770 45.595 31.875 ;
        RECT 50.705 31.770 51.165 31.825 ;
        RECT 45.135 31.330 51.165 31.770 ;
        RECT 45.135 31.305 45.595 31.330 ;
        RECT 50.705 31.255 51.165 31.330 ;
        RECT 41.055 12.350 41.555 12.360 ;
        RECT 28.345 11.115 30.465 12.265 ;
        RECT 41.065 11.965 41.555 12.350 ;
        RECT 51.635 12.145 52.125 73.030 ;
        RECT 61.260 73.010 64.060 74.530 ;
        RECT 72.340 73.050 75.020 74.980 ;
        RECT 83.730 74.540 86.290 75.690 ;
        RECT 95.655 75.580 96.285 83.245 ;
        RECT 106.975 75.640 107.605 84.485 ;
        RECT 118.225 75.650 118.855 85.545 ;
        RECT 129.975 75.650 130.605 86.595 ;
        RECT 133.330 76.605 136.060 77.855 ;
        RECT 137.190 76.585 139.920 77.835 ;
        RECT 53.815 54.020 54.275 54.095 ;
        RECT 59.385 54.020 59.845 54.045 ;
        RECT 53.815 53.580 59.845 54.020 ;
        RECT 53.815 53.525 54.275 53.580 ;
        RECT 59.385 53.475 59.845 53.580 ;
        RECT 56.075 48.830 56.555 48.895 ;
        RECT 56.075 48.510 57.875 48.830 ;
        RECT 56.075 48.345 56.555 48.510 ;
        RECT 57.305 45.670 57.865 48.510 ;
        RECT 61.185 45.670 61.665 45.695 ;
        RECT 57.305 45.250 61.665 45.670 ;
        RECT 57.305 45.240 57.865 45.250 ;
        RECT 61.185 45.145 61.665 45.250 ;
        RECT 54.535 40.100 55.015 40.205 ;
        RECT 58.335 40.100 58.895 40.110 ;
        RECT 54.535 39.680 58.895 40.100 ;
        RECT 54.535 39.655 55.015 39.680 ;
        RECT 58.335 36.840 58.895 39.680 ;
        RECT 59.645 36.840 60.125 37.005 ;
        RECT 58.325 36.520 60.125 36.840 ;
        RECT 59.645 36.455 60.125 36.520 ;
        RECT 56.355 31.770 56.815 31.875 ;
        RECT 61.925 31.770 62.385 31.825 ;
        RECT 56.355 31.330 62.385 31.770 ;
        RECT 56.355 31.305 56.815 31.330 ;
        RECT 61.925 31.255 62.385 31.330 ;
        RECT 29.765 11.100 30.255 11.115 ;
        RECT 39.065 11.005 41.615 11.965 ;
        RECT 50.285 10.995 52.405 12.145 ;
        RECT 62.915 12.135 63.405 73.010 ;
        RECT 65.035 54.010 65.495 54.085 ;
        RECT 70.605 54.010 71.065 54.035 ;
        RECT 65.035 53.570 71.065 54.010 ;
        RECT 65.035 53.515 65.495 53.570 ;
        RECT 70.605 53.465 71.065 53.570 ;
        RECT 67.295 48.820 67.775 48.885 ;
        RECT 67.295 48.500 69.095 48.820 ;
        RECT 67.295 48.335 67.775 48.500 ;
        RECT 68.525 45.660 69.085 48.500 ;
        RECT 72.405 45.660 72.885 45.685 ;
        RECT 68.525 45.240 72.885 45.660 ;
        RECT 68.525 45.230 69.085 45.240 ;
        RECT 72.405 45.135 72.885 45.240 ;
        RECT 65.735 40.100 66.215 40.205 ;
        RECT 69.535 40.100 70.095 40.110 ;
        RECT 65.735 39.680 70.095 40.100 ;
        RECT 65.735 39.655 66.215 39.680 ;
        RECT 69.535 36.840 70.095 39.680 ;
        RECT 70.845 36.840 71.325 37.005 ;
        RECT 69.525 36.520 71.325 36.840 ;
        RECT 70.845 36.455 71.325 36.520 ;
        RECT 67.555 31.770 68.015 31.875 ;
        RECT 73.125 31.770 73.585 31.825 ;
        RECT 67.555 31.330 73.585 31.770 ;
        RECT 67.555 31.305 68.015 31.330 ;
        RECT 73.125 31.255 73.585 31.330 ;
        RECT 74.055 12.165 74.545 73.050 ;
        RECT 83.690 73.000 86.290 74.540 ;
        RECT 94.960 74.710 97.520 75.580 ;
        RECT 94.960 73.020 97.570 74.710 ;
        RECT 106.340 74.460 108.900 75.640 ;
        RECT 117.470 74.720 120.030 75.650 ;
        RECT 76.275 54.000 76.735 54.075 ;
        RECT 81.845 54.000 82.305 54.025 ;
        RECT 76.275 53.560 82.305 54.000 ;
        RECT 76.275 53.505 76.735 53.560 ;
        RECT 81.845 53.455 82.305 53.560 ;
        RECT 78.535 48.810 79.015 48.875 ;
        RECT 78.535 48.490 80.335 48.810 ;
        RECT 78.535 48.325 79.015 48.490 ;
        RECT 79.765 45.650 80.325 48.490 ;
        RECT 83.645 45.650 84.125 45.675 ;
        RECT 79.765 45.230 84.125 45.650 ;
        RECT 79.765 45.220 80.325 45.230 ;
        RECT 83.645 45.125 84.125 45.230 ;
        RECT 77.025 40.090 77.505 40.195 ;
        RECT 80.825 40.090 81.385 40.100 ;
        RECT 77.025 39.670 81.385 40.090 ;
        RECT 77.025 39.645 77.505 39.670 ;
        RECT 80.825 36.830 81.385 39.670 ;
        RECT 82.135 36.830 82.615 36.995 ;
        RECT 80.815 36.510 82.615 36.830 ;
        RECT 82.135 36.445 82.615 36.510 ;
        RECT 78.845 31.760 79.305 31.865 ;
        RECT 84.415 31.760 84.875 31.815 ;
        RECT 78.845 31.320 84.875 31.760 ;
        RECT 78.845 31.295 79.305 31.320 ;
        RECT 84.415 31.245 84.875 31.320 ;
        RECT 61.365 10.985 63.485 12.135 ;
        RECT 72.675 11.015 74.795 12.165 ;
        RECT 85.375 12.155 85.865 73.000 ;
        RECT 87.525 54.010 87.985 54.085 ;
        RECT 93.095 54.010 93.555 54.035 ;
        RECT 87.525 53.570 93.555 54.010 ;
        RECT 87.525 53.515 87.985 53.570 ;
        RECT 93.095 53.465 93.555 53.570 ;
        RECT 89.785 48.820 90.265 48.885 ;
        RECT 89.785 48.500 91.585 48.820 ;
        RECT 89.785 48.335 90.265 48.500 ;
        RECT 91.015 45.660 91.575 48.500 ;
        RECT 94.895 45.660 95.375 45.685 ;
        RECT 91.015 45.240 95.375 45.660 ;
        RECT 91.015 45.230 91.575 45.240 ;
        RECT 94.895 45.135 95.375 45.240 ;
        RECT 88.265 40.110 88.745 40.215 ;
        RECT 92.065 40.110 92.625 40.120 ;
        RECT 88.265 39.690 92.625 40.110 ;
        RECT 88.265 39.665 88.745 39.690 ;
        RECT 92.065 36.850 92.625 39.690 ;
        RECT 93.375 36.850 93.855 37.015 ;
        RECT 92.055 36.530 93.855 36.850 ;
        RECT 93.375 36.465 93.855 36.530 ;
        RECT 90.085 31.780 90.545 31.885 ;
        RECT 95.655 31.780 96.115 31.835 ;
        RECT 90.085 31.340 96.115 31.780 ;
        RECT 90.085 31.315 90.545 31.340 ;
        RECT 95.655 31.265 96.115 31.340 ;
        RECT 96.605 12.155 97.095 73.020 ;
        RECT 106.150 73.000 109.060 74.460 ;
        RECT 117.470 73.070 120.000 74.720 ;
        RECT 129.290 74.650 131.850 75.650 ;
        RECT 129.300 73.140 131.820 74.650 ;
        RECT 98.805 54.000 99.265 54.075 ;
        RECT 104.375 54.000 104.835 54.025 ;
        RECT 98.805 53.560 104.835 54.000 ;
        RECT 98.805 53.505 99.265 53.560 ;
        RECT 104.375 53.455 104.835 53.560 ;
        RECT 101.065 48.810 101.545 48.875 ;
        RECT 101.065 48.490 102.865 48.810 ;
        RECT 101.065 48.325 101.545 48.490 ;
        RECT 102.295 45.650 102.855 48.490 ;
        RECT 106.175 45.650 106.655 45.675 ;
        RECT 102.295 45.230 106.655 45.650 ;
        RECT 102.295 45.220 102.855 45.230 ;
        RECT 106.175 45.125 106.655 45.230 ;
        RECT 99.475 40.130 99.955 40.235 ;
        RECT 103.275 40.130 103.835 40.140 ;
        RECT 99.475 39.710 103.835 40.130 ;
        RECT 99.475 39.685 99.955 39.710 ;
        RECT 103.275 36.870 103.835 39.710 ;
        RECT 104.585 36.870 105.065 37.035 ;
        RECT 103.265 36.550 105.065 36.870 ;
        RECT 104.585 36.485 105.065 36.550 ;
        RECT 101.295 31.800 101.755 31.905 ;
        RECT 106.865 31.800 107.325 31.855 ;
        RECT 101.295 31.360 107.325 31.800 ;
        RECT 101.295 31.335 101.755 31.360 ;
        RECT 106.865 31.285 107.325 31.360 ;
        RECT 107.865 12.205 108.355 73.000 ;
        RECT 110.075 54.000 110.535 54.075 ;
        RECT 115.645 54.000 116.105 54.025 ;
        RECT 110.075 53.560 116.105 54.000 ;
        RECT 110.075 53.505 110.535 53.560 ;
        RECT 115.645 53.455 116.105 53.560 ;
        RECT 112.335 48.810 112.815 48.875 ;
        RECT 112.335 48.490 114.135 48.810 ;
        RECT 112.335 48.325 112.815 48.490 ;
        RECT 113.565 45.650 114.125 48.490 ;
        RECT 117.445 45.650 117.925 45.675 ;
        RECT 113.565 45.230 117.925 45.650 ;
        RECT 113.565 45.220 114.125 45.230 ;
        RECT 117.445 45.125 117.925 45.230 ;
        RECT 110.675 40.170 111.155 40.275 ;
        RECT 114.475 40.170 115.035 40.180 ;
        RECT 110.675 39.750 115.035 40.170 ;
        RECT 110.675 39.725 111.155 39.750 ;
        RECT 114.475 36.910 115.035 39.750 ;
        RECT 115.785 36.910 116.265 37.075 ;
        RECT 114.465 36.590 116.265 36.910 ;
        RECT 115.785 36.525 116.265 36.590 ;
        RECT 112.495 31.840 112.955 31.945 ;
        RECT 118.065 31.840 118.525 31.895 ;
        RECT 112.495 31.400 118.525 31.840 ;
        RECT 112.495 31.375 112.955 31.400 ;
        RECT 118.065 31.325 118.525 31.400 ;
        RECT 119.085 12.205 119.575 73.070 ;
        RECT 121.325 54.000 121.785 54.075 ;
        RECT 126.895 54.000 127.355 54.025 ;
        RECT 121.325 53.560 127.355 54.000 ;
        RECT 121.325 53.505 121.785 53.560 ;
        RECT 126.895 53.455 127.355 53.560 ;
        RECT 123.585 48.810 124.065 48.875 ;
        RECT 123.585 48.490 125.385 48.810 ;
        RECT 123.585 48.325 124.065 48.490 ;
        RECT 124.815 45.650 125.375 48.490 ;
        RECT 128.695 45.650 129.175 45.675 ;
        RECT 124.815 45.230 129.175 45.650 ;
        RECT 124.815 45.220 125.375 45.230 ;
        RECT 128.695 45.125 129.175 45.230 ;
        RECT 121.885 40.190 122.365 40.295 ;
        RECT 125.685 40.190 126.245 40.200 ;
        RECT 121.885 39.770 126.245 40.190 ;
        RECT 121.885 39.745 122.365 39.770 ;
        RECT 125.685 36.930 126.245 39.770 ;
        RECT 126.995 36.930 127.475 37.095 ;
        RECT 125.675 36.610 127.475 36.930 ;
        RECT 126.995 36.545 127.475 36.610 ;
        RECT 123.705 31.860 124.165 31.965 ;
        RECT 129.275 31.860 129.735 31.915 ;
        RECT 123.705 31.420 129.735 31.860 ;
        RECT 123.705 31.395 124.165 31.420 ;
        RECT 129.275 31.345 129.735 31.420 ;
        RECT 130.335 12.235 130.825 73.140 ;
        RECT 74.055 11.010 74.545 11.015 ;
        RECT 83.795 11.005 85.915 12.155 ;
        RECT 95.095 11.005 97.215 12.155 ;
        RECT 106.285 11.055 108.405 12.205 ;
        RECT 117.515 11.055 119.635 12.205 ;
        RECT 128.815 11.085 130.935 12.235 ;
        RECT 107.865 11.010 108.355 11.055 ;
        RECT 119.085 11.050 119.575 11.055 ;
        RECT 85.375 11.000 85.865 11.005 ;
        RECT 96.605 10.980 97.095 11.005 ;
        RECT 74.290 0.135 75.680 1.435 ;
        RECT 93.500 0.205 94.890 1.505 ;
        RECT 112.900 0.335 114.290 1.635 ;
        RECT 131.800 0.405 133.540 1.905 ;
        RECT 151.600 0.275 152.970 1.445 ;
      LAYER met4 ;
        RECT 30.420 225.130 30.670 225.140 ;
        RECT 30.300 224.760 30.670 225.130 ;
        RECT 30.970 224.760 33.430 225.140 ;
        RECT 33.730 224.760 36.190 225.140 ;
        RECT 36.490 224.760 38.950 225.140 ;
        RECT 39.250 224.760 41.710 225.140 ;
        RECT 42.010 224.760 44.470 225.140 ;
        RECT 44.770 224.760 47.230 225.140 ;
        RECT 47.530 224.760 49.990 225.140 ;
        RECT 50.290 224.760 52.750 225.140 ;
        RECT 53.050 224.760 55.510 225.140 ;
        RECT 55.810 224.760 58.270 225.140 ;
        RECT 58.570 224.760 61.030 225.140 ;
        RECT 61.330 224.760 63.790 225.140 ;
        RECT 64.090 224.760 66.550 225.140 ;
        RECT 66.850 224.760 69.310 225.140 ;
        RECT 69.610 224.760 72.070 225.140 ;
        RECT 72.370 224.760 74.830 225.140 ;
        RECT 75.130 224.760 77.590 225.140 ;
        RECT 77.890 224.760 80.350 225.140 ;
        RECT 80.650 224.760 83.110 225.140 ;
        RECT 83.410 224.760 85.870 225.140 ;
        RECT 86.170 224.760 88.630 225.140 ;
        RECT 88.930 224.760 91.390 225.140 ;
        RECT 91.690 224.760 94.150 225.140 ;
        RECT 94.450 224.760 96.910 225.140 ;
        RECT 97.210 224.760 99.670 225.140 ;
        RECT 99.970 224.760 102.430 225.140 ;
        RECT 102.730 224.760 105.190 225.140 ;
        RECT 105.490 224.760 107.950 225.140 ;
        RECT 108.250 224.760 110.710 225.140 ;
        RECT 111.010 224.760 113.470 225.140 ;
        RECT 113.770 224.760 116.230 225.140 ;
        RECT 116.530 224.760 118.990 225.140 ;
        RECT 119.290 224.760 121.750 225.140 ;
        RECT 122.050 224.760 124.510 225.140 ;
        RECT 124.810 224.760 127.270 225.140 ;
        RECT 127.570 224.760 130.030 225.140 ;
        RECT 130.330 224.760 132.790 225.140 ;
        RECT 133.090 224.760 133.520 225.140 ;
        RECT 30.300 224.240 133.520 224.760 ;
        RECT 135.385 224.760 135.550 225.185 ;
        RECT 135.850 224.760 136.745 225.185 ;
        RECT 30.300 219.100 31.660 224.240 ;
        RECT 135.385 223.875 136.745 224.760 ;
        RECT 138.175 224.760 138.310 225.115 ;
        RECT 138.610 224.760 139.535 225.115 ;
        RECT 138.175 223.805 139.535 224.760 ;
        RECT 143.225 224.760 143.830 225.145 ;
        RECT 144.130 224.760 144.585 225.145 ;
        RECT 143.225 223.835 144.585 224.760 ;
        RECT 6.000 218.040 31.660 219.100 ;
        RECT 30.300 217.960 31.660 218.040 ;
        RECT 17.450 105.870 19.450 204.270 ;
        RECT 32.450 105.870 34.450 204.270 ;
        RECT 41.065 177.005 41.395 177.335 ;
        RECT 41.080 138.575 41.380 177.005 ;
        RECT 41.985 174.285 42.315 174.615 ;
        RECT 41.065 138.245 41.395 138.575 ;
        RECT 42.000 137.895 42.300 174.285 ;
        RECT 42.905 166.805 43.235 167.135 ;
        RECT 42.920 150.135 43.220 166.805 ;
        RECT 42.905 149.805 43.235 150.135 ;
        RECT 42.920 138.575 43.220 149.805 ;
        RECT 42.905 138.245 43.235 138.575 ;
        RECT 41.985 137.565 42.315 137.895 ;
        RECT 47.450 105.870 49.450 204.270 ;
        RECT 62.450 105.870 64.450 204.270 ;
        RECT 65.905 180.405 66.235 180.735 ;
        RECT 65.920 135.175 66.220 180.405 ;
        RECT 67.745 174.285 68.075 174.615 ;
        RECT 70.505 174.285 70.835 174.615 ;
        RECT 67.760 138.575 68.060 174.285 ;
        RECT 70.520 146.055 70.820 174.285 ;
        RECT 71.425 149.805 71.755 150.135 ;
        RECT 70.505 145.725 70.835 146.055 ;
        RECT 67.745 138.245 68.075 138.575 ;
        RECT 65.905 134.845 66.235 135.175 ;
        RECT 71.440 111.375 71.740 149.805 ;
        RECT 71.425 111.045 71.755 111.375 ;
        RECT 77.450 105.870 79.450 204.270 ;
        RECT 81.545 158.645 81.875 158.975 ;
        RECT 81.560 151.495 81.860 158.645 ;
        RECT 81.545 151.165 81.875 151.495 ;
        RECT 81.560 135.175 81.860 151.165 ;
        RECT 81.545 134.845 81.875 135.175 ;
        RECT 92.450 105.870 94.450 204.270 ;
        RECT 95.345 155.925 95.675 156.255 ;
        RECT 95.360 137.895 95.660 155.925 ;
        RECT 98.105 147.765 98.435 148.095 ;
        RECT 98.120 139.935 98.420 147.765 ;
        RECT 98.105 139.605 98.435 139.935 ;
        RECT 95.345 137.565 95.675 137.895 ;
        RECT 107.450 105.870 109.450 204.270 ;
        RECT 118.110 97.700 120.130 99.670 ;
        RECT 121.810 97.750 123.830 99.720 ;
        RECT 118.130 93.980 120.130 97.700 ;
        RECT 121.820 96.830 123.820 97.750 ;
        RECT 121.820 94.830 139.410 96.830 ;
        RECT 118.130 91.980 135.580 93.980 ;
        RECT 133.580 77.835 135.580 91.980 ;
        RECT 133.375 76.625 136.015 77.835 ;
        RECT 137.410 77.815 139.410 94.830 ;
        RECT 137.235 76.605 139.875 77.815 ;
        RECT 3.955 71.365 4.000 73.195 ;
        RECT 6.000 71.365 6.055 73.195 ;
        RECT 3.000 68.705 3.025 70.435 ;
        RECT 15.555 68.655 16.995 71.165 ;
        RECT 74.335 1.000 75.635 1.415 ;
        RECT 74.335 0.155 74.530 1.000 ;
        RECT 75.430 0.155 75.635 1.000 ;
        RECT 93.545 1.000 94.845 1.485 ;
        RECT 93.545 0.225 93.850 1.000 ;
        RECT 94.750 0.225 94.845 1.000 ;
        RECT 112.945 1.000 114.245 1.615 ;
        RECT 112.945 0.355 113.170 1.000 ;
        RECT 114.070 0.355 114.245 1.000 ;
        RECT 131.845 1.000 133.495 1.885 ;
        RECT 131.845 0.425 132.490 1.000 ;
        RECT 133.390 0.425 133.495 1.000 ;
        RECT 151.645 1.000 152.925 1.425 ;
        RECT 151.645 0.295 151.810 1.000 ;
        RECT 152.710 0.295 152.925 1.000 ;
  END
END tt_um_08_sws
END LIBRARY

