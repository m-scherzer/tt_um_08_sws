MACRO sky130_fd_sc_hd__fill_2
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_hd__fill_2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 0.920 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 -0.085 0.920 0.000 ;
      LAYER met1 ;
        RECT 0.100 0.000 0.365 0.090 ;
        RECT 0.000 -0.240 0.920 0.000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.155 -0.050 0.315 0.060 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190 2.720 1.110 2.910 ;
        RECT -0.190 1.305 0.000 2.720 ;
        RECT 0.140 2.675 0.310 2.720 ;
        RECT 0.920 1.305 1.110 2.720 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 0.000 2.720 0.920 2.805 ;
      LAYER met1 ;
        RECT 0.000 2.720 0.920 2.960 ;
        RECT 0.105 2.650 0.365 2.720 ;
    END
  END VPWR
  OBS
      LAYER nwell ;
        RECT 0.000 2.675 0.140 2.720 ;
        RECT 0.310 2.675 0.920 2.720 ;
        RECT 0.000 1.305 0.920 2.675 ;
      LAYER li1 ;
        RECT 0.000 2.635 0.920 2.720 ;
        RECT 0.000 0.000 0.920 0.085 ;
      LAYER met1 ;
        RECT 0.000 2.650 0.105 2.720 ;
        RECT 0.365 2.650 0.920 2.720 ;
        RECT 0.000 2.480 0.920 2.650 ;
        RECT 0.000 0.090 0.920 0.240 ;
        RECT 0.000 0.000 0.100 0.090 ;
        RECT 0.365 0.000 0.920 0.090 ;
  END
END sky130_fd_sc_hd__fill_2
END LIBRARY

