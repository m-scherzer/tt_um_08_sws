VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_08_sws
  CLASS BLOCK ;
  FOREIGN tt_um_08_sws ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ua[0]
    ANTENNAGATEAREA 200.000000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    ANTENNAGATEAREA 550.000000 ;
    ANTENNADIFFAREA 2.900000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    ANTENNADIFFAREA 29.000000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    PORT
      LAYER met4 ;
        RECT 55.210 0.000 56.110 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    PORT
      LAYER met4 ;
        RECT 35.890 0.000 36.790 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    PORT
      LAYER met4 ;
        RECT 16.570 0.000 17.470 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    ANTENNADIFFAREA 36.399998 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    ANTENNADIFFAREA 394.109192 ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 18.310 193.515 18.480 193.705 ;
        RECT 19.745 193.565 19.865 193.675 ;
        RECT 21.530 193.515 21.700 193.705 ;
        RECT 23.370 193.515 23.540 193.705 ;
        RECT 28.890 193.515 29.060 193.705 ;
        RECT 34.410 193.515 34.580 193.705 ;
        RECT 36.250 193.515 36.420 193.705 ;
        RECT 41.770 193.515 41.940 193.705 ;
        RECT 47.290 193.515 47.460 193.705 ;
        RECT 49.130 193.515 49.300 193.705 ;
        RECT 54.650 193.515 54.820 193.705 ;
        RECT 60.170 193.515 60.340 193.705 ;
        RECT 62.010 193.515 62.180 193.705 ;
        RECT 67.530 193.515 67.700 193.705 ;
        RECT 73.050 193.515 73.220 193.705 ;
        RECT 74.890 193.515 75.060 193.705 ;
        RECT 80.410 193.515 80.580 193.705 ;
        RECT 85.930 193.515 86.100 193.705 ;
        RECT 87.770 193.515 87.940 193.705 ;
        RECT 93.290 193.515 93.460 193.705 ;
        RECT 98.810 193.515 98.980 193.705 ;
        RECT 99.785 193.565 99.905 193.675 ;
        RECT 105.250 193.515 105.420 193.705 ;
        RECT 110.770 193.515 110.940 193.705 ;
        RECT 112.150 193.515 112.320 193.705 ;
        RECT 18.170 192.705 19.540 193.515 ;
        RECT 20.010 192.705 21.840 193.515 ;
        RECT 21.860 192.645 22.290 193.430 ;
        RECT 22.310 192.705 23.680 193.515 ;
        RECT 23.690 192.705 29.200 193.515 ;
        RECT 29.210 192.705 34.720 193.515 ;
        RECT 34.740 192.645 35.170 193.430 ;
        RECT 35.190 192.705 36.560 193.515 ;
        RECT 36.570 192.705 42.080 193.515 ;
        RECT 42.090 192.705 47.600 193.515 ;
        RECT 47.620 192.645 48.050 193.430 ;
        RECT 48.070 192.705 49.440 193.515 ;
        RECT 49.450 192.705 54.960 193.515 ;
        RECT 54.970 192.705 60.480 193.515 ;
        RECT 60.500 192.645 60.930 193.430 ;
        RECT 60.950 192.705 62.320 193.515 ;
        RECT 62.330 192.705 67.840 193.515 ;
        RECT 67.850 192.705 73.360 193.515 ;
        RECT 73.380 192.645 73.810 193.430 ;
        RECT 73.830 192.705 75.200 193.515 ;
        RECT 75.210 192.705 80.720 193.515 ;
        RECT 80.730 192.705 86.240 193.515 ;
        RECT 86.260 192.645 86.690 193.430 ;
        RECT 86.710 192.705 88.080 193.515 ;
        RECT 88.090 192.705 93.600 193.515 ;
        RECT 93.610 192.705 99.120 193.515 ;
        RECT 99.140 192.645 99.570 193.430 ;
        RECT 100.050 192.705 105.560 193.515 ;
        RECT 105.570 192.705 111.080 193.515 ;
        RECT 111.090 192.705 112.460 193.515 ;
      LAYER nwell ;
        RECT 17.975 189.485 112.655 192.315 ;
      LAYER pwell ;
        RECT 18.170 188.285 19.540 189.095 ;
        RECT 20.010 188.285 23.680 189.095 ;
        RECT 23.690 188.285 29.200 189.095 ;
        RECT 29.210 188.285 34.720 189.095 ;
        RECT 34.740 188.370 35.170 189.155 ;
        RECT 35.650 188.285 38.400 189.095 ;
        RECT 38.410 188.285 43.920 189.095 ;
        RECT 43.930 188.285 49.440 189.095 ;
        RECT 49.450 188.285 54.960 189.095 ;
        RECT 54.970 188.285 60.480 189.095 ;
        RECT 60.500 188.370 60.930 189.155 ;
        RECT 60.950 188.285 62.780 189.095 ;
        RECT 62.790 188.285 68.300 189.095 ;
        RECT 68.320 188.285 69.670 189.195 ;
        RECT 69.690 188.285 75.200 189.095 ;
        RECT 75.210 188.285 80.720 189.095 ;
        RECT 80.730 188.285 86.240 189.095 ;
        RECT 86.260 188.370 86.690 189.155 ;
        RECT 87.170 188.285 89.000 189.095 ;
        RECT 89.010 188.285 94.520 189.095 ;
        RECT 94.530 188.285 100.040 189.095 ;
        RECT 100.050 188.285 105.560 189.095 ;
        RECT 105.570 188.285 111.080 189.095 ;
        RECT 111.090 188.285 112.460 189.095 ;
        RECT 18.310 188.075 18.480 188.285 ;
        RECT 19.745 188.125 19.865 188.235 ;
        RECT 21.530 188.075 21.700 188.265 ;
        RECT 22.505 188.125 22.625 188.235 ;
        RECT 23.370 188.095 23.540 188.285 ;
        RECT 25.210 188.075 25.380 188.265 ;
        RECT 28.890 188.095 29.060 188.285 ;
        RECT 30.730 188.075 30.900 188.265 ;
        RECT 34.410 188.095 34.580 188.285 ;
        RECT 35.385 188.125 35.505 188.235 ;
        RECT 36.250 188.075 36.420 188.265 ;
        RECT 38.090 188.095 38.260 188.285 ;
        RECT 41.770 188.075 41.940 188.265 ;
        RECT 43.610 188.095 43.780 188.285 ;
        RECT 47.290 188.075 47.460 188.265 ;
        RECT 49.130 188.095 49.300 188.285 ;
        RECT 50.510 188.075 50.680 188.265 ;
        RECT 54.650 188.095 54.820 188.285 ;
        RECT 56.030 188.075 56.200 188.265 ;
        RECT 57.410 188.075 57.580 188.265 ;
        RECT 57.870 188.075 58.040 188.265 ;
        RECT 60.170 188.095 60.340 188.285 ;
        RECT 62.470 188.095 62.640 188.285 ;
        RECT 67.990 188.075 68.160 188.285 ;
        RECT 69.370 188.095 69.540 188.285 ;
        RECT 71.210 188.075 71.380 188.265 ;
        RECT 73.050 188.075 73.220 188.265 ;
        RECT 74.430 188.120 74.590 188.230 ;
        RECT 74.890 188.095 75.060 188.285 ;
        RECT 78.110 188.075 78.280 188.265 ;
        RECT 80.410 188.095 80.580 188.285 ;
        RECT 83.630 188.075 83.800 188.265 ;
        RECT 85.930 188.095 86.100 188.285 ;
        RECT 86.905 188.125 87.025 188.235 ;
        RECT 88.690 188.095 88.860 188.285 ;
        RECT 89.150 188.075 89.320 188.265 ;
        RECT 94.210 188.095 94.380 188.285 ;
        RECT 94.670 188.075 94.840 188.265 ;
        RECT 95.130 188.075 95.300 188.265 ;
        RECT 98.810 188.075 98.980 188.265 ;
        RECT 99.730 188.235 99.900 188.285 ;
        RECT 99.730 188.125 99.905 188.235 ;
        RECT 99.730 188.095 99.900 188.125 ;
        RECT 105.250 188.075 105.420 188.285 ;
        RECT 110.770 188.075 110.940 188.285 ;
        RECT 112.150 188.075 112.320 188.285 ;
        RECT 18.170 187.265 19.540 188.075 ;
        RECT 20.010 187.265 21.840 188.075 ;
        RECT 21.860 187.205 22.290 187.990 ;
        RECT 22.770 187.265 25.520 188.075 ;
        RECT 25.530 187.265 31.040 188.075 ;
        RECT 31.050 187.265 36.560 188.075 ;
        RECT 36.570 187.265 42.080 188.075 ;
        RECT 42.090 187.265 47.600 188.075 ;
        RECT 47.620 187.205 48.050 187.990 ;
        RECT 48.070 187.265 50.820 188.075 ;
        RECT 50.830 187.265 56.340 188.075 ;
        RECT 56.360 187.165 57.710 188.075 ;
        RECT 57.740 187.165 59.090 188.075 ;
        RECT 59.110 187.395 68.300 188.075 ;
        RECT 59.110 187.165 60.030 187.395 ;
        RECT 62.860 187.175 63.790 187.395 ;
        RECT 68.310 187.165 71.420 188.075 ;
        RECT 71.530 187.265 73.360 188.075 ;
        RECT 73.380 187.205 73.810 187.990 ;
        RECT 74.750 187.265 78.420 188.075 ;
        RECT 78.430 187.265 83.940 188.075 ;
        RECT 83.950 187.265 89.460 188.075 ;
        RECT 89.470 187.265 94.980 188.075 ;
        RECT 95.000 187.165 96.350 188.075 ;
        RECT 96.370 187.265 99.120 188.075 ;
        RECT 99.140 187.205 99.570 187.990 ;
        RECT 100.050 187.265 105.560 188.075 ;
        RECT 105.570 187.265 111.080 188.075 ;
        RECT 111.090 187.265 112.460 188.075 ;
      LAYER nwell ;
        RECT 17.975 184.045 112.655 186.875 ;
      LAYER pwell ;
        RECT 18.170 182.845 19.540 183.655 ;
        RECT 20.010 182.845 23.680 183.655 ;
        RECT 23.690 182.845 29.200 183.655 ;
        RECT 29.210 182.845 34.720 183.655 ;
        RECT 34.740 182.930 35.170 183.715 ;
        RECT 35.190 182.845 36.560 183.655 ;
        RECT 36.570 182.845 40.240 183.655 ;
        RECT 40.250 182.845 45.760 183.655 ;
        RECT 45.770 182.845 51.280 183.655 ;
        RECT 55.800 183.525 56.730 183.745 ;
        RECT 59.560 183.525 60.480 183.755 ;
        RECT 51.290 182.845 60.480 183.525 ;
        RECT 60.500 182.930 60.930 183.715 ;
        RECT 61.435 183.525 62.780 183.755 ;
        RECT 60.950 182.845 62.780 183.525 ;
        RECT 63.710 182.845 65.080 183.625 ;
        RECT 65.090 183.525 66.010 183.755 ;
        RECT 68.840 183.525 69.770 183.745 ;
        RECT 65.090 182.845 74.280 183.525 ;
        RECT 74.300 182.845 75.650 183.755 ;
        RECT 75.670 182.845 78.420 183.655 ;
        RECT 78.440 182.845 79.790 183.755 ;
        RECT 83.010 183.525 83.940 183.755 ;
        RECT 80.040 182.845 83.940 183.525 ;
        RECT 83.950 182.845 85.320 183.625 ;
        RECT 86.260 182.930 86.690 183.715 ;
        RECT 86.720 182.845 88.070 183.755 ;
        RECT 92.600 183.525 93.530 183.745 ;
        RECT 96.360 183.525 97.280 183.755 ;
        RECT 88.090 182.845 97.280 183.525 ;
        RECT 97.290 183.525 98.210 183.755 ;
        RECT 101.040 183.525 101.970 183.745 ;
        RECT 97.290 182.845 106.480 183.525 ;
        RECT 107.410 182.845 111.080 183.655 ;
        RECT 111.090 182.845 112.460 183.655 ;
        RECT 18.310 182.635 18.480 182.845 ;
        RECT 19.745 182.685 19.865 182.795 ;
        RECT 21.530 182.635 21.700 182.825 ;
        RECT 22.505 182.685 22.625 182.795 ;
        RECT 23.370 182.655 23.540 182.845 ;
        RECT 25.210 182.635 25.380 182.825 ;
        RECT 28.890 182.655 29.060 182.845 ;
        RECT 30.730 182.635 30.900 182.825 ;
        RECT 34.410 182.655 34.580 182.845 ;
        RECT 36.250 182.635 36.420 182.845 ;
        RECT 39.930 182.655 40.100 182.845 ;
        RECT 41.770 182.635 41.940 182.825 ;
        RECT 45.450 182.655 45.620 182.845 ;
        RECT 47.290 182.635 47.460 182.825 ;
        RECT 50.970 182.655 51.140 182.845 ;
        RECT 51.430 182.635 51.600 182.845 ;
        RECT 56.950 182.635 57.120 182.825 ;
        RECT 57.410 182.635 57.580 182.825 ;
        RECT 61.090 182.635 61.260 182.845 ;
        RECT 63.390 182.690 63.550 182.800 ;
        RECT 64.770 182.655 64.940 182.845 ;
        RECT 65.690 182.635 65.860 182.825 ;
        RECT 67.530 182.655 67.700 182.825 ;
        RECT 67.535 182.635 67.700 182.655 ;
        RECT 71.670 182.635 71.840 182.825 ;
        RECT 73.050 182.635 73.220 182.825 ;
        RECT 73.970 182.655 74.140 182.845 ;
        RECT 74.430 182.655 74.600 182.845 ;
        RECT 76.270 182.635 76.440 182.825 ;
        RECT 76.730 182.635 76.900 182.825 ;
        RECT 78.110 182.655 78.280 182.845 ;
        RECT 78.570 182.655 78.740 182.845 ;
        RECT 83.355 182.655 83.525 182.845 ;
        RECT 84.090 182.655 84.260 182.845 ;
        RECT 85.930 182.690 86.090 182.800 ;
        RECT 86.850 182.635 87.020 182.845 ;
        RECT 87.365 182.685 87.485 182.795 ;
        RECT 88.230 182.655 88.400 182.845 ;
        RECT 89.150 182.635 89.320 182.825 ;
        RECT 90.530 182.635 90.700 182.825 ;
        RECT 91.265 182.635 91.435 182.825 ;
        RECT 98.535 182.635 98.705 182.825 ;
        RECT 99.730 182.635 99.900 182.825 ;
        RECT 101.570 182.680 101.730 182.790 ;
        RECT 105.250 182.635 105.420 182.825 ;
        RECT 106.170 182.655 106.340 182.845 ;
        RECT 107.090 182.690 107.250 182.800 ;
        RECT 110.770 182.635 110.940 182.845 ;
        RECT 112.150 182.635 112.320 182.845 ;
        RECT 18.170 181.825 19.540 182.635 ;
        RECT 20.010 181.825 21.840 182.635 ;
        RECT 21.860 181.765 22.290 182.550 ;
        RECT 22.770 181.825 25.520 182.635 ;
        RECT 25.530 181.825 31.040 182.635 ;
        RECT 31.050 181.825 36.560 182.635 ;
        RECT 36.570 181.825 42.080 182.635 ;
        RECT 42.090 181.825 47.600 182.635 ;
        RECT 47.620 181.765 48.050 182.550 ;
        RECT 48.070 181.825 51.740 182.635 ;
        RECT 51.750 181.825 57.260 182.635 ;
        RECT 57.270 181.955 60.940 182.635 ;
        RECT 60.950 182.405 62.520 182.635 ;
        RECT 64.610 182.595 65.530 182.635 ;
        RECT 64.610 182.405 65.540 182.595 ;
        RECT 60.950 182.045 65.540 182.405 ;
        RECT 60.950 181.955 65.530 182.045 ;
        RECT 65.550 181.955 67.380 182.635 ;
        RECT 67.535 181.955 69.370 182.635 ;
        RECT 60.010 181.725 60.940 181.955 ;
        RECT 62.530 181.725 65.530 181.955 ;
        RECT 68.440 181.725 69.370 181.955 ;
        RECT 69.690 181.955 71.980 182.635 ;
        RECT 69.690 181.725 70.610 181.955 ;
        RECT 71.990 181.825 73.360 182.635 ;
        RECT 73.380 181.765 73.810 182.550 ;
        RECT 73.830 181.825 76.580 182.635 ;
        RECT 76.600 181.725 77.950 182.635 ;
        RECT 77.970 181.955 87.160 182.635 ;
        RECT 77.970 181.725 78.890 181.955 ;
        RECT 81.720 181.735 82.650 181.955 ;
        RECT 87.630 181.825 89.460 182.635 ;
        RECT 89.470 181.855 90.840 182.635 ;
        RECT 90.850 181.955 94.750 182.635 ;
        RECT 95.220 181.955 99.120 182.635 ;
        RECT 90.850 181.725 91.780 181.955 ;
        RECT 98.190 181.725 99.120 181.955 ;
        RECT 99.140 181.765 99.570 182.550 ;
        RECT 99.590 181.855 100.960 182.635 ;
        RECT 101.890 181.825 105.560 182.635 ;
        RECT 105.570 181.825 111.080 182.635 ;
        RECT 111.090 181.825 112.460 182.635 ;
      LAYER nwell ;
        RECT 17.975 178.605 112.655 181.435 ;
      LAYER pwell ;
        RECT 18.170 177.405 19.540 178.215 ;
        RECT 20.010 177.405 23.680 178.215 ;
        RECT 23.690 177.405 29.200 178.215 ;
        RECT 29.210 177.405 34.720 178.215 ;
        RECT 34.740 177.490 35.170 178.275 ;
        RECT 35.190 177.405 37.020 178.215 ;
        RECT 37.030 177.405 42.540 178.215 ;
        RECT 42.560 177.405 43.910 178.315 ;
        RECT 44.300 178.205 45.220 178.315 ;
        RECT 44.300 178.085 46.635 178.205 ;
        RECT 51.300 178.085 52.220 178.305 ;
        RECT 44.300 177.405 53.580 178.085 ;
        RECT 53.590 177.405 54.960 178.215 ;
        RECT 54.970 177.405 58.640 178.215 ;
        RECT 58.650 177.405 60.480 178.085 ;
        RECT 60.500 177.490 60.930 178.275 ;
        RECT 63.240 178.085 64.160 178.315 ;
        RECT 61.870 177.405 64.160 178.085 ;
        RECT 64.170 177.405 67.090 178.315 ;
        RECT 67.390 177.405 68.760 178.185 ;
        RECT 68.790 177.405 70.140 178.315 ;
        RECT 71.070 177.405 74.740 178.215 ;
        RECT 75.120 178.205 76.040 178.315 ;
        RECT 75.120 178.085 77.455 178.205 ;
        RECT 82.120 178.085 83.040 178.305 ;
        RECT 75.120 177.405 84.400 178.085 ;
        RECT 84.410 177.405 85.780 178.185 ;
        RECT 86.260 177.490 86.690 178.275 ;
        RECT 86.710 177.405 92.220 178.215 ;
        RECT 92.240 177.405 93.590 178.315 ;
        RECT 93.610 178.085 94.530 178.315 ;
        RECT 97.360 178.085 98.290 178.305 ;
        RECT 93.610 177.405 102.800 178.085 ;
        RECT 102.810 177.405 104.180 178.185 ;
        RECT 104.190 177.405 105.560 178.215 ;
        RECT 105.570 177.405 111.080 178.215 ;
        RECT 111.090 177.405 112.460 178.215 ;
        RECT 18.310 177.195 18.480 177.405 ;
        RECT 19.745 177.245 19.865 177.355 ;
        RECT 21.530 177.195 21.700 177.385 ;
        RECT 22.910 177.240 23.070 177.350 ;
        RECT 23.370 177.215 23.540 177.405 ;
        RECT 26.590 177.195 26.760 177.385 ;
        RECT 28.890 177.215 29.060 177.405 ;
        RECT 32.110 177.195 32.280 177.385 ;
        RECT 34.410 177.215 34.580 177.405 ;
        RECT 36.710 177.215 36.880 177.405 ;
        RECT 37.630 177.195 37.800 177.385 ;
        RECT 42.230 177.215 42.400 177.405 ;
        RECT 43.610 177.215 43.780 177.405 ;
        RECT 47.290 177.195 47.460 177.385 ;
        RECT 49.130 177.195 49.300 177.385 ;
        RECT 50.050 177.240 50.210 177.350 ;
        RECT 50.510 177.195 50.680 177.385 ;
        RECT 52.810 177.195 52.980 177.385 ;
        RECT 53.270 177.215 53.440 177.405 ;
        RECT 54.190 177.195 54.360 177.385 ;
        RECT 54.650 177.355 54.820 177.405 ;
        RECT 54.650 177.245 54.825 177.355 ;
        RECT 54.650 177.215 54.820 177.245 ;
        RECT 58.330 177.215 58.500 177.405 ;
        RECT 58.790 177.215 58.960 177.405 ;
        RECT 61.550 177.250 61.710 177.360 ;
        RECT 62.010 177.215 62.180 177.405 ;
        RECT 64.315 177.215 64.485 177.405 ;
        RECT 65.230 177.195 65.400 177.385 ;
        RECT 18.170 176.385 19.540 177.195 ;
        RECT 20.010 176.385 21.840 177.195 ;
        RECT 21.860 176.325 22.290 177.110 ;
        RECT 23.230 176.385 26.900 177.195 ;
        RECT 26.910 176.385 32.420 177.195 ;
        RECT 32.430 176.385 37.940 177.195 ;
        RECT 38.320 176.515 47.600 177.195 ;
        RECT 38.320 176.395 40.655 176.515 ;
        RECT 38.320 176.285 39.240 176.395 ;
        RECT 45.320 176.295 46.240 176.515 ;
        RECT 47.620 176.325 48.050 177.110 ;
        RECT 48.080 176.285 49.430 177.195 ;
        RECT 50.370 176.415 51.740 177.195 ;
        RECT 51.760 176.285 53.110 177.195 ;
        RECT 53.130 176.415 54.500 177.195 ;
        RECT 55.170 176.515 65.540 177.195 ;
        RECT 65.690 177.165 65.860 177.385 ;
        RECT 68.450 177.215 68.620 177.405 ;
        RECT 68.905 177.355 69.075 177.405 ;
        RECT 68.905 177.245 69.085 177.355 ;
        RECT 70.750 177.250 70.910 177.360 ;
        RECT 68.905 177.215 69.075 177.245 ;
        RECT 72.775 177.195 72.945 177.385 ;
        RECT 74.430 177.215 74.600 177.405 ;
        RECT 83.170 177.195 83.340 177.385 ;
        RECT 83.685 177.245 83.805 177.355 ;
        RECT 84.090 177.215 84.260 177.405 ;
        RECT 85.470 177.195 85.640 177.405 ;
        RECT 85.930 177.355 86.100 177.385 ;
        RECT 85.930 177.245 86.105 177.355 ;
        RECT 87.365 177.245 87.485 177.355 ;
        RECT 85.930 177.195 86.100 177.245 ;
        RECT 87.770 177.195 87.940 177.385 ;
        RECT 91.910 177.215 92.080 177.405 ;
        RECT 92.370 177.215 92.540 177.405 ;
        RECT 97.890 177.195 98.060 177.385 ;
        RECT 98.810 177.240 98.970 177.350 ;
        RECT 99.785 177.245 99.905 177.355 ;
        RECT 101.570 177.195 101.740 177.385 ;
        RECT 102.030 177.195 102.200 177.385 ;
        RECT 102.490 177.215 102.660 177.405 ;
        RECT 103.870 177.215 104.040 177.405 ;
        RECT 104.330 177.195 104.500 177.385 ;
        RECT 105.250 177.215 105.420 177.405 ;
        RECT 110.770 177.195 110.940 177.405 ;
        RECT 112.150 177.195 112.320 177.405 ;
        RECT 67.815 177.165 68.760 177.195 ;
        RECT 65.690 176.965 68.760 177.165 ;
        RECT 55.170 176.285 57.380 176.515 ;
        RECT 60.100 176.295 61.030 176.515 ;
        RECT 65.550 176.485 68.760 176.965 ;
        RECT 69.460 176.515 73.360 177.195 ;
        RECT 65.550 176.285 66.480 176.485 ;
        RECT 67.815 176.285 68.760 176.485 ;
        RECT 72.430 176.285 73.360 176.515 ;
        RECT 73.380 176.325 73.810 177.110 ;
        RECT 74.200 176.515 83.480 177.195 ;
        RECT 74.200 176.395 76.535 176.515 ;
        RECT 74.200 176.285 75.120 176.395 ;
        RECT 81.200 176.295 82.120 176.515 ;
        RECT 83.950 176.385 85.780 177.195 ;
        RECT 85.800 176.285 87.150 177.195 ;
        RECT 87.630 176.415 89.000 177.195 ;
        RECT 89.010 176.515 98.200 177.195 ;
        RECT 89.010 176.285 89.930 176.515 ;
        RECT 92.760 176.295 93.690 176.515 ;
        RECT 99.140 176.325 99.570 177.110 ;
        RECT 100.050 176.385 101.880 177.195 ;
        RECT 101.900 176.285 103.250 177.195 ;
        RECT 103.280 176.285 104.630 177.195 ;
        RECT 105.570 176.385 111.080 177.195 ;
        RECT 111.090 176.385 112.460 177.195 ;
      LAYER nwell ;
        RECT 17.975 173.165 112.655 175.995 ;
      LAYER pwell ;
        RECT 18.170 171.965 19.540 172.775 ;
        RECT 20.010 171.965 23.680 172.775 ;
        RECT 23.690 171.965 29.200 172.775 ;
        RECT 29.210 171.965 34.720 172.775 ;
        RECT 34.740 172.050 35.170 172.835 ;
        RECT 35.650 171.965 38.400 172.775 ;
        RECT 38.420 171.965 39.770 172.875 ;
        RECT 42.990 172.645 43.920 172.875 ;
        RECT 47.130 172.645 48.060 172.875 ;
        RECT 40.020 171.965 43.920 172.645 ;
        RECT 44.160 171.965 48.060 172.645 ;
        RECT 48.440 172.765 49.360 172.875 ;
        RECT 48.440 172.645 50.775 172.765 ;
        RECT 55.440 172.645 56.360 172.865 ;
        RECT 48.440 171.965 57.720 172.645 ;
        RECT 57.730 171.965 59.100 172.775 ;
        RECT 59.120 171.965 60.470 172.875 ;
        RECT 60.500 172.050 60.930 172.835 ;
        RECT 61.880 171.965 63.230 172.875 ;
        RECT 64.170 172.675 65.100 172.875 ;
        RECT 66.435 172.675 67.380 172.875 ;
        RECT 64.170 172.195 67.380 172.675 ;
        RECT 64.310 171.995 67.380 172.195 ;
        RECT 18.310 171.755 18.480 171.965 ;
        RECT 19.745 171.805 19.865 171.915 ;
        RECT 21.530 171.755 21.700 171.945 ;
        RECT 22.505 171.805 22.625 171.915 ;
        RECT 23.370 171.775 23.540 171.965 ;
        RECT 25.210 171.755 25.380 171.945 ;
        RECT 25.670 171.755 25.840 171.945 ;
        RECT 27.050 171.755 27.220 171.945 ;
        RECT 28.430 171.755 28.600 171.945 ;
        RECT 28.890 171.775 29.060 171.965 ;
        RECT 29.815 171.755 29.985 171.945 ;
        RECT 33.490 171.755 33.660 171.945 ;
        RECT 34.410 171.775 34.580 171.965 ;
        RECT 35.385 171.805 35.505 171.915 ;
        RECT 38.090 171.775 38.260 171.965 ;
        RECT 38.550 171.775 38.720 171.965 ;
        RECT 42.745 171.805 42.865 171.915 ;
        RECT 43.335 171.775 43.505 171.965 ;
        RECT 45.450 171.755 45.620 171.945 ;
        RECT 46.830 171.755 47.000 171.945 ;
        RECT 47.345 171.805 47.465 171.915 ;
        RECT 47.475 171.775 47.645 171.965 ;
        RECT 48.265 171.805 48.385 171.915 ;
        RECT 48.670 171.755 48.840 171.945 ;
        RECT 53.455 171.755 53.625 171.945 ;
        RECT 54.190 171.755 54.360 171.945 ;
        RECT 55.570 171.755 55.740 171.945 ;
        RECT 57.410 171.775 57.580 171.965 ;
        RECT 58.790 171.775 58.960 171.965 ;
        RECT 60.170 171.775 60.340 171.965 ;
        RECT 61.550 171.810 61.710 171.920 ;
        RECT 62.930 171.775 63.100 171.965 ;
        RECT 63.850 171.810 64.010 171.920 ;
        RECT 64.310 171.775 64.480 171.995 ;
        RECT 66.435 171.965 67.380 171.995 ;
        RECT 67.390 171.965 70.500 172.875 ;
        RECT 70.610 171.965 72.900 172.875 ;
        RECT 73.840 171.965 75.190 172.875 ;
        RECT 78.410 172.645 79.340 172.875 ;
        RECT 75.440 171.965 79.340 172.645 ;
        RECT 80.270 171.965 81.640 172.745 ;
        RECT 81.650 171.965 83.020 172.745 ;
        RECT 83.030 171.965 84.860 172.775 ;
        RECT 84.880 171.965 86.230 172.875 ;
        RECT 86.260 172.050 86.690 172.835 ;
        RECT 86.710 172.645 87.630 172.875 ;
        RECT 90.460 172.645 91.390 172.865 ;
        RECT 99.110 172.645 100.040 172.875 ;
        RECT 86.710 171.965 95.900 172.645 ;
        RECT 96.140 171.965 100.040 172.645 ;
        RECT 100.970 172.645 101.890 172.875 ;
        RECT 104.720 172.645 105.650 172.865 ;
        RECT 100.970 171.965 110.160 172.645 ;
        RECT 111.090 171.965 112.460 172.775 ;
        RECT 67.990 171.755 68.160 171.945 ;
        RECT 68.455 171.755 68.625 171.945 ;
        RECT 70.290 171.775 70.460 171.965 ;
        RECT 70.755 171.775 70.925 171.965 ;
        RECT 71.265 171.805 71.385 171.915 ;
        RECT 73.050 171.755 73.220 171.945 ;
        RECT 73.510 171.810 73.670 171.920 ;
        RECT 73.970 171.775 74.140 171.965 ;
        RECT 74.430 171.800 74.590 171.910 ;
        RECT 74.890 171.755 75.060 171.945 ;
        RECT 78.755 171.775 78.925 171.965 ;
        RECT 79.950 171.810 80.110 171.920 ;
        RECT 81.330 171.775 81.500 171.965 ;
        RECT 82.710 171.775 82.880 171.965 ;
        RECT 84.550 171.775 84.720 171.965 ;
        RECT 85.010 171.755 85.180 171.965 ;
        RECT 85.525 171.805 85.645 171.915 ;
        RECT 87.310 171.755 87.480 171.945 ;
        RECT 88.045 171.755 88.215 171.945 ;
        RECT 92.370 171.800 92.530 171.910 ;
        RECT 95.590 171.775 95.760 171.965 ;
        RECT 96.235 171.755 96.405 171.945 ;
        RECT 97.890 171.755 98.060 171.945 ;
        RECT 98.810 171.800 98.970 171.910 ;
        RECT 99.455 171.775 99.625 171.965 ;
        RECT 100.190 171.800 100.350 171.910 ;
        RECT 100.650 171.810 100.810 171.920 ;
        RECT 109.390 171.755 109.560 171.945 ;
        RECT 109.850 171.775 110.020 171.965 ;
        RECT 110.770 171.755 110.940 171.945 ;
        RECT 112.150 171.755 112.320 171.965 ;
        RECT 18.170 170.945 19.540 171.755 ;
        RECT 20.010 170.945 21.840 171.755 ;
        RECT 21.860 170.885 22.290 171.670 ;
        RECT 22.770 170.945 25.520 171.755 ;
        RECT 25.540 170.845 26.890 171.755 ;
        RECT 26.920 170.845 28.270 171.755 ;
        RECT 28.290 170.975 29.660 171.755 ;
        RECT 29.670 170.845 33.145 171.755 ;
        RECT 33.350 171.075 42.540 171.755 ;
        RECT 37.860 170.855 38.790 171.075 ;
        RECT 41.620 170.845 42.540 171.075 ;
        RECT 43.010 170.945 45.760 171.755 ;
        RECT 45.770 170.975 47.140 171.755 ;
        RECT 47.620 170.885 48.050 171.670 ;
        RECT 48.540 170.845 49.890 171.755 ;
        RECT 50.140 171.075 54.040 171.755 ;
        RECT 53.110 170.845 54.040 171.075 ;
        RECT 54.050 170.975 55.420 171.755 ;
        RECT 55.540 171.075 59.005 171.755 ;
        RECT 58.085 170.845 59.005 171.075 ;
        RECT 59.110 171.075 68.300 171.755 ;
        RECT 59.110 170.845 60.030 171.075 ;
        RECT 62.860 170.855 63.790 171.075 ;
        RECT 68.310 170.845 70.920 171.755 ;
        RECT 71.530 170.945 73.360 171.755 ;
        RECT 73.380 170.885 73.810 171.670 ;
        RECT 74.760 170.845 76.110 171.755 ;
        RECT 76.130 171.075 85.320 171.755 ;
        RECT 76.130 170.845 77.050 171.075 ;
        RECT 79.880 170.855 80.810 171.075 ;
        RECT 85.790 170.945 87.620 171.755 ;
        RECT 87.630 171.075 91.530 171.755 ;
        RECT 92.920 171.075 96.820 171.755 ;
        RECT 87.630 170.845 88.560 171.075 ;
        RECT 95.890 170.845 96.820 171.075 ;
        RECT 96.830 170.975 98.200 171.755 ;
        RECT 99.140 170.885 99.570 171.670 ;
        RECT 100.510 171.075 109.700 171.755 ;
        RECT 100.510 170.845 101.430 171.075 ;
        RECT 104.260 170.855 105.190 171.075 ;
        RECT 109.710 170.975 111.080 171.755 ;
        RECT 111.090 170.945 112.460 171.755 ;
      LAYER nwell ;
        RECT 17.975 167.725 112.655 170.555 ;
      LAYER pwell ;
        RECT 18.170 166.525 19.540 167.335 ;
        RECT 20.010 166.525 25.520 167.335 ;
        RECT 30.040 167.205 30.970 167.425 ;
        RECT 33.800 167.205 34.720 167.435 ;
        RECT 25.530 166.525 34.720 167.205 ;
        RECT 34.740 166.610 35.170 167.395 ;
        RECT 35.190 166.525 36.560 167.305 ;
        RECT 36.570 167.205 37.490 167.435 ;
        RECT 40.320 167.205 41.250 167.425 ;
        RECT 36.570 166.525 45.760 167.205 ;
        RECT 45.770 166.525 49.245 167.435 ;
        RECT 53.570 167.205 54.500 167.435 ;
        RECT 50.600 166.525 54.500 167.205 ;
        RECT 54.970 166.525 56.340 167.305 ;
        RECT 56.810 166.525 60.480 167.335 ;
        RECT 60.500 166.610 60.930 167.395 ;
        RECT 60.950 166.525 64.620 167.335 ;
        RECT 64.630 166.525 70.140 167.335 ;
        RECT 70.150 166.525 72.760 167.435 ;
        RECT 72.910 167.205 73.830 167.435 ;
        RECT 76.660 167.205 77.590 167.425 ;
        RECT 85.310 167.205 86.240 167.435 ;
        RECT 72.910 166.525 82.100 167.205 ;
        RECT 82.340 166.525 86.240 167.205 ;
        RECT 86.260 166.610 86.690 167.395 ;
        RECT 86.710 166.525 88.080 167.305 ;
        RECT 88.100 166.525 89.450 167.435 ;
        RECT 90.400 166.525 91.750 167.435 ;
        RECT 96.280 167.205 97.210 167.425 ;
        RECT 100.040 167.205 100.960 167.435 ;
        RECT 104.170 167.205 105.100 167.435 ;
        RECT 91.770 166.525 100.960 167.205 ;
        RECT 101.200 166.525 105.100 167.205 ;
        RECT 105.570 166.525 106.940 167.305 ;
        RECT 107.410 166.525 111.080 167.335 ;
        RECT 111.090 166.525 112.460 167.335 ;
        RECT 18.310 166.315 18.480 166.525 ;
        RECT 19.745 166.365 19.865 166.475 ;
        RECT 21.530 166.315 21.700 166.505 ;
        RECT 22.450 166.315 22.620 166.505 ;
        RECT 23.830 166.315 24.000 166.505 ;
        RECT 25.210 166.335 25.380 166.525 ;
        RECT 25.670 166.335 25.840 166.525 ;
        RECT 33.030 166.315 33.200 166.505 ;
        RECT 36.250 166.335 36.420 166.525 ;
        RECT 36.985 166.315 37.155 166.505 ;
        RECT 44.255 166.315 44.425 166.505 ;
        RECT 45.450 166.335 45.620 166.525 ;
        RECT 45.915 166.505 46.085 166.525 ;
        RECT 45.910 166.335 46.085 166.505 ;
        RECT 45.910 166.315 46.080 166.335 ;
        RECT 46.370 166.315 46.540 166.505 ;
        RECT 49.590 166.315 49.760 166.505 ;
        RECT 50.050 166.370 50.210 166.480 ;
        RECT 53.915 166.335 54.085 166.525 ;
        RECT 54.705 166.365 54.825 166.475 ;
        RECT 55.110 166.335 55.280 166.525 ;
        RECT 56.545 166.365 56.665 166.475 ;
        RECT 59.250 166.315 59.420 166.505 ;
        RECT 60.170 166.335 60.340 166.525 ;
        RECT 60.630 166.315 60.800 166.505 ;
        RECT 64.310 166.315 64.480 166.525 ;
        RECT 64.770 166.315 64.940 166.505 ;
        RECT 66.150 166.335 66.320 166.505 ;
        RECT 69.830 166.335 70.000 166.525 ;
        RECT 70.295 166.335 70.465 166.525 ;
        RECT 72.130 166.335 72.300 166.505 ;
        RECT 73.050 166.360 73.210 166.470 ;
        RECT 74.430 166.360 74.590 166.470 ;
        RECT 66.250 166.315 66.320 166.335 ;
        RECT 72.130 166.315 72.200 166.335 ;
        RECT 74.890 166.315 75.060 166.505 ;
        RECT 79.675 166.315 79.845 166.505 ;
        RECT 81.790 166.335 81.960 166.525 ;
        RECT 83.170 166.335 83.340 166.505 ;
        RECT 84.550 166.315 84.720 166.505 ;
        RECT 85.065 166.365 85.185 166.475 ;
        RECT 85.655 166.335 85.825 166.525 ;
        RECT 87.770 166.335 87.940 166.525 ;
        RECT 89.150 166.335 89.320 166.525 ;
        RECT 90.070 166.370 90.230 166.480 ;
        RECT 90.530 166.335 90.700 166.525 ;
        RECT 91.910 166.335 92.080 166.525 ;
        RECT 94.210 166.315 94.380 166.505 ;
        RECT 94.945 166.315 95.115 166.505 ;
        RECT 98.865 166.365 98.985 166.475 ;
        RECT 99.785 166.365 99.905 166.475 ;
        RECT 103.595 166.315 103.765 166.505 ;
        RECT 104.330 166.315 104.500 166.505 ;
        RECT 104.515 166.335 104.685 166.525 ;
        RECT 105.305 166.365 105.425 166.475 ;
        RECT 105.710 166.335 105.880 166.525 ;
        RECT 106.170 166.360 106.330 166.470 ;
        RECT 106.630 166.315 106.800 166.505 ;
        RECT 107.145 166.365 107.265 166.475 ;
        RECT 108.065 166.365 108.185 166.475 ;
        RECT 110.770 166.315 110.940 166.525 ;
        RECT 112.150 166.315 112.320 166.525 ;
        RECT 18.170 165.505 19.540 166.315 ;
        RECT 20.010 165.505 21.840 166.315 ;
        RECT 21.860 165.445 22.290 166.230 ;
        RECT 22.310 165.535 23.680 166.315 ;
        RECT 23.690 165.635 32.880 166.315 ;
        RECT 33.000 165.635 36.465 166.315 ;
        RECT 28.200 165.415 29.130 165.635 ;
        RECT 31.960 165.405 32.880 165.635 ;
        RECT 35.545 165.405 36.465 165.635 ;
        RECT 36.570 165.635 40.470 166.315 ;
        RECT 40.940 165.635 44.840 166.315 ;
        RECT 36.570 165.405 37.500 165.635 ;
        RECT 43.910 165.405 44.840 165.635 ;
        RECT 44.850 165.505 46.220 166.315 ;
        RECT 46.240 165.405 47.590 166.315 ;
        RECT 47.620 165.445 48.050 166.230 ;
        RECT 48.070 165.505 49.900 166.315 ;
        RECT 50.280 165.635 59.560 166.315 ;
        RECT 50.280 165.515 52.615 165.635 ;
        RECT 50.280 165.405 51.200 165.515 ;
        RECT 57.280 165.415 58.200 165.635 ;
        RECT 59.580 165.405 60.930 166.315 ;
        RECT 60.950 165.505 64.620 166.315 ;
        RECT 64.640 165.405 65.990 166.315 ;
        RECT 66.250 166.085 68.520 166.315 ;
        RECT 69.930 166.085 72.200 166.315 ;
        RECT 66.250 165.405 69.005 166.085 ;
        RECT 69.445 165.405 72.200 166.085 ;
        RECT 73.380 165.445 73.810 166.230 ;
        RECT 74.760 165.405 76.110 166.315 ;
        RECT 76.360 165.635 80.260 166.315 ;
        RECT 80.650 165.635 83.075 166.315 ;
        RECT 79.330 165.405 80.260 165.635 ;
        RECT 83.500 165.405 84.850 166.315 ;
        RECT 85.330 165.635 94.520 166.315 ;
        RECT 94.530 165.635 98.430 166.315 ;
        RECT 85.330 165.405 86.250 165.635 ;
        RECT 89.080 165.415 90.010 165.635 ;
        RECT 94.530 165.405 95.460 165.635 ;
        RECT 99.140 165.445 99.570 166.230 ;
        RECT 100.280 165.635 104.180 166.315 ;
        RECT 103.250 165.405 104.180 165.635 ;
        RECT 104.200 165.405 105.550 166.315 ;
        RECT 106.490 165.535 107.860 166.315 ;
        RECT 108.330 165.505 111.080 166.315 ;
        RECT 111.090 165.505 112.460 166.315 ;
      LAYER nwell ;
        RECT 17.975 162.285 112.655 165.115 ;
      LAYER pwell ;
        RECT 18.170 161.085 19.540 161.895 ;
        RECT 19.550 161.085 21.380 161.895 ;
        RECT 21.400 161.085 22.750 161.995 ;
        RECT 22.780 161.085 24.130 161.995 ;
        RECT 24.150 161.085 25.520 161.895 ;
        RECT 25.530 161.765 26.450 161.995 ;
        RECT 29.280 161.765 30.210 161.985 ;
        RECT 25.530 161.085 34.720 161.765 ;
        RECT 34.740 161.170 35.170 161.955 ;
        RECT 35.190 161.765 36.120 161.995 ;
        RECT 35.190 161.085 39.090 161.765 ;
        RECT 40.445 161.085 43.920 161.995 ;
        RECT 43.930 161.085 47.405 161.995 ;
        RECT 47.980 161.885 48.900 161.995 ;
        RECT 47.980 161.765 50.315 161.885 ;
        RECT 54.980 161.765 55.900 161.985 ;
        RECT 47.980 161.085 57.260 161.765 ;
        RECT 57.730 161.085 59.100 161.865 ;
        RECT 59.110 161.085 60.480 161.865 ;
        RECT 60.500 161.170 60.930 161.955 ;
        RECT 61.650 161.315 64.405 161.995 ;
        RECT 66.210 161.765 69.210 161.995 ;
        RECT 85.310 161.765 86.240 161.995 ;
        RECT 64.630 161.675 69.210 161.765 ;
        RECT 64.630 161.315 69.220 161.675 ;
        RECT 61.650 161.085 63.920 161.315 ;
        RECT 64.630 161.085 66.200 161.315 ;
        RECT 68.290 161.125 69.220 161.315 ;
        RECT 68.290 161.085 69.210 161.125 ;
        RECT 69.230 161.085 71.970 161.765 ;
        RECT 71.990 161.085 81.095 161.765 ;
        RECT 82.340 161.085 86.240 161.765 ;
        RECT 86.260 161.170 86.690 161.955 ;
        RECT 86.720 161.085 88.070 161.995 ;
        RECT 89.010 161.085 90.375 161.765 ;
        RECT 90.850 161.085 92.220 161.865 ;
        RECT 92.690 161.085 95.440 161.895 ;
        RECT 95.450 161.085 96.820 161.865 ;
        RECT 100.030 161.765 100.960 161.995 ;
        RECT 97.060 161.085 100.960 161.765 ;
        RECT 100.970 161.765 101.890 161.995 ;
        RECT 104.720 161.765 105.650 161.985 ;
        RECT 100.970 161.085 110.160 161.765 ;
        RECT 111.090 161.085 112.460 161.895 ;
        RECT 18.310 160.875 18.480 161.085 ;
        RECT 20.150 160.920 20.310 161.030 ;
        RECT 20.610 160.875 20.780 161.065 ;
        RECT 21.070 160.895 21.240 161.085 ;
        RECT 21.530 160.895 21.700 161.085 ;
        RECT 22.505 160.925 22.625 161.035 ;
        RECT 23.830 160.895 24.000 161.085 ;
        RECT 25.210 161.065 25.380 161.085 ;
        RECT 25.205 160.895 25.380 161.065 ;
        RECT 25.205 160.875 25.375 160.895 ;
        RECT 25.945 160.875 26.115 161.065 ;
        RECT 29.865 160.925 29.985 161.035 ;
        RECT 31.650 160.875 31.820 161.065 ;
        RECT 34.410 160.895 34.580 161.085 ;
        RECT 35.605 160.895 35.775 161.085 ;
        RECT 43.605 161.065 43.775 161.085 ;
        RECT 39.930 160.930 40.090 161.040 ;
        RECT 40.850 160.875 41.020 161.065 ;
        RECT 43.605 160.895 43.780 161.065 ;
        RECT 43.610 160.875 43.780 160.895 ;
        RECT 44.075 160.875 44.245 161.085 ;
        RECT 51.615 160.875 51.785 161.065 ;
        RECT 52.355 160.875 52.525 161.065 ;
        RECT 56.950 160.895 57.120 161.085 ;
        RECT 57.410 161.035 57.580 161.065 ;
        RECT 57.410 160.925 57.585 161.035 ;
        RECT 57.925 160.925 58.045 161.035 ;
        RECT 57.410 160.875 57.580 160.925 ;
        RECT 58.790 160.895 58.960 161.085 ;
        RECT 59.250 160.895 59.420 161.085 ;
        RECT 61.650 161.065 61.720 161.085 ;
        RECT 59.710 160.875 59.880 161.065 ;
        RECT 61.145 160.925 61.265 161.035 ;
        RECT 61.550 160.875 61.720 161.065 ;
        RECT 62.010 160.875 62.180 161.065 ;
        RECT 63.390 160.875 63.560 161.065 ;
        RECT 64.770 160.895 64.940 161.085 ;
        RECT 66.150 160.895 66.320 161.065 ;
        RECT 69.370 160.895 69.540 161.085 ;
        RECT 66.250 160.875 66.320 160.895 ;
        RECT 70.290 160.875 70.460 161.065 ;
        RECT 70.750 160.875 70.920 161.065 ;
        RECT 72.130 160.895 72.300 161.085 ;
        RECT 74.430 160.920 74.590 161.030 ;
        RECT 81.790 160.930 81.950 161.040 ;
        RECT 84.090 160.875 84.260 161.065 ;
        RECT 85.470 160.875 85.640 161.065 ;
        RECT 85.655 160.895 85.825 161.085 ;
        RECT 87.770 160.895 87.940 161.085 ;
        RECT 88.690 160.930 88.850 161.040 ;
        RECT 89.145 160.875 89.315 161.065 ;
        RECT 90.530 160.895 90.700 161.065 ;
        RECT 90.990 160.895 91.160 161.085 ;
        RECT 92.425 160.925 92.545 161.035 ;
        RECT 93.015 160.875 93.185 161.065 ;
        RECT 93.750 160.875 93.920 161.065 ;
        RECT 95.130 161.035 95.300 161.085 ;
        RECT 95.130 160.925 95.305 161.035 ;
        RECT 95.130 160.895 95.300 160.925 ;
        RECT 95.595 160.875 95.765 161.065 ;
        RECT 96.510 160.895 96.680 161.085 ;
        RECT 100.375 160.895 100.545 161.085 ;
        RECT 102.945 160.875 103.115 161.065 ;
        RECT 103.870 160.920 104.030 161.030 ;
        RECT 104.330 160.875 104.500 161.065 ;
        RECT 106.630 160.875 106.800 161.065 ;
        RECT 108.470 160.875 108.640 161.065 ;
        RECT 108.985 160.925 109.105 161.035 ;
        RECT 109.850 160.895 110.020 161.085 ;
        RECT 110.770 160.875 110.940 161.065 ;
        RECT 112.150 160.875 112.320 161.085 ;
        RECT 18.170 160.065 19.540 160.875 ;
        RECT 20.470 160.095 21.840 160.875 ;
        RECT 21.860 160.005 22.290 160.790 ;
        RECT 22.910 159.965 25.520 160.875 ;
        RECT 25.530 160.195 29.430 160.875 ;
        RECT 25.530 159.965 26.460 160.195 ;
        RECT 30.130 160.065 31.960 160.875 ;
        RECT 31.970 160.195 41.160 160.875 ;
        RECT 41.180 160.195 43.920 160.875 ;
        RECT 31.970 159.965 32.890 160.195 ;
        RECT 35.720 159.975 36.650 160.195 ;
        RECT 43.930 159.965 47.405 160.875 ;
        RECT 47.620 160.005 48.050 160.790 ;
        RECT 48.300 160.195 52.200 160.875 ;
        RECT 51.270 159.965 52.200 160.195 ;
        RECT 52.210 159.965 54.820 160.875 ;
        RECT 54.980 160.195 57.720 160.875 ;
        RECT 58.190 160.195 60.020 160.875 ;
        RECT 60.030 160.195 61.860 160.875 ;
        RECT 58.190 159.965 59.535 160.195 ;
        RECT 60.030 159.965 61.375 160.195 ;
        RECT 61.870 160.095 63.240 160.875 ;
        RECT 63.250 159.965 65.970 160.875 ;
        RECT 66.250 160.645 68.520 160.875 ;
        RECT 66.250 159.965 69.005 160.645 ;
        RECT 69.230 160.065 70.600 160.875 ;
        RECT 70.610 160.195 73.350 160.875 ;
        RECT 73.380 160.005 73.810 160.790 ;
        RECT 75.120 160.195 84.400 160.875 ;
        RECT 75.120 160.075 77.455 160.195 ;
        RECT 75.120 159.965 76.040 160.075 ;
        RECT 82.120 159.975 83.040 160.195 ;
        RECT 84.410 160.095 85.780 160.875 ;
        RECT 85.985 159.965 89.460 160.875 ;
        RECT 89.700 160.195 93.600 160.875 ;
        RECT 92.670 159.965 93.600 160.195 ;
        RECT 93.610 160.095 94.980 160.875 ;
        RECT 95.450 159.965 98.925 160.875 ;
        RECT 99.140 160.005 99.570 160.790 ;
        RECT 99.785 159.965 103.260 160.875 ;
        RECT 104.200 159.965 105.550 160.875 ;
        RECT 105.570 160.065 106.940 160.875 ;
        RECT 106.950 160.195 108.780 160.875 ;
        RECT 109.250 160.065 111.080 160.875 ;
        RECT 111.090 160.065 112.460 160.875 ;
      LAYER nwell ;
        RECT 17.975 156.845 112.655 159.675 ;
      LAYER pwell ;
        RECT 18.170 155.645 19.540 156.455 ;
        RECT 19.550 156.325 20.470 156.555 ;
        RECT 23.300 156.325 24.230 156.545 ;
        RECT 19.550 155.645 28.740 156.325 ;
        RECT 29.220 155.645 30.570 156.555 ;
        RECT 33.790 156.325 34.720 156.555 ;
        RECT 30.820 155.645 34.720 156.325 ;
        RECT 34.740 155.730 35.170 156.515 ;
        RECT 35.190 155.645 36.560 156.455 ;
        RECT 36.765 155.645 40.240 156.555 ;
        RECT 40.445 155.645 43.920 156.555 ;
        RECT 44.015 155.645 53.120 156.325 ;
        RECT 53.130 155.645 56.290 156.555 ;
        RECT 56.350 156.325 57.695 156.555 ;
        RECT 56.350 155.645 58.180 156.325 ;
        RECT 59.110 155.645 60.480 156.425 ;
        RECT 60.500 155.730 60.930 156.515 ;
        RECT 62.355 156.325 63.700 156.555 ;
        RECT 61.870 155.645 63.700 156.325 ;
        RECT 64.630 156.325 65.975 156.555 ;
        RECT 64.630 155.645 66.460 156.325 ;
        RECT 66.510 155.645 71.060 156.555 ;
        RECT 74.270 156.325 75.200 156.555 ;
        RECT 71.300 155.645 75.200 156.325 ;
        RECT 75.580 156.445 76.500 156.555 ;
        RECT 75.580 156.325 77.915 156.445 ;
        RECT 82.580 156.325 83.500 156.545 ;
        RECT 75.580 155.645 84.860 156.325 ;
        RECT 84.870 155.645 86.240 156.425 ;
        RECT 86.260 155.730 86.690 156.515 ;
        RECT 87.080 156.445 88.000 156.555 ;
        RECT 87.080 156.325 89.415 156.445 ;
        RECT 94.080 156.325 95.000 156.545 ;
        RECT 100.030 156.325 100.960 156.555 ;
        RECT 87.080 155.645 96.360 156.325 ;
        RECT 97.060 155.645 100.960 156.325 ;
        RECT 101.340 156.445 102.260 156.555 ;
        RECT 101.340 156.325 103.675 156.445 ;
        RECT 108.340 156.325 109.260 156.545 ;
        RECT 101.340 155.645 110.620 156.325 ;
        RECT 111.090 155.645 112.460 156.455 ;
        RECT 18.310 155.435 18.480 155.645 ;
        RECT 19.745 155.485 19.865 155.595 ;
        RECT 21.530 155.435 21.700 155.625 ;
        RECT 22.505 155.485 22.625 155.595 ;
        RECT 22.910 155.435 23.080 155.625 ;
        RECT 24.565 155.435 24.735 155.625 ;
        RECT 28.430 155.455 28.600 155.645 ;
        RECT 28.945 155.485 29.065 155.595 ;
        RECT 29.810 155.435 29.980 155.625 ;
        RECT 30.270 155.455 30.440 155.645 ;
        RECT 34.135 155.455 34.305 155.645 ;
        RECT 36.250 155.455 36.420 155.645 ;
        RECT 39.010 155.435 39.180 155.625 ;
        RECT 39.525 155.485 39.645 155.595 ;
        RECT 39.925 155.455 40.095 155.645 ;
        RECT 41.310 155.435 41.480 155.625 ;
        RECT 41.775 155.435 41.945 155.625 ;
        RECT 43.605 155.455 43.775 155.645 ;
        RECT 45.505 155.485 45.625 155.595 ;
        RECT 47.290 155.435 47.460 155.625 ;
        RECT 48.215 155.435 48.385 155.625 ;
        RECT 52.810 155.435 52.980 155.645 ;
        RECT 56.030 155.455 56.200 155.645 ;
        RECT 57.870 155.455 58.040 155.645 ;
        RECT 58.790 155.490 58.950 155.600 ;
        RECT 59.250 155.455 59.420 155.645 ;
        RECT 61.550 155.490 61.710 155.600 ;
        RECT 62.010 155.455 62.180 155.645 ;
        RECT 62.470 155.435 62.640 155.625 ;
        RECT 62.930 155.435 63.100 155.625 ;
        RECT 64.310 155.490 64.470 155.600 ;
        RECT 65.690 155.435 65.860 155.625 ;
        RECT 66.150 155.455 66.320 155.645 ;
        RECT 69.365 155.435 69.535 155.625 ;
        RECT 70.750 155.455 70.920 155.645 ;
        RECT 73.045 155.435 73.215 155.625 ;
        RECT 74.615 155.455 74.785 155.645 ;
        RECT 76.270 155.435 76.440 155.625 ;
        RECT 80.135 155.435 80.305 155.625 ;
        RECT 81.330 155.480 81.490 155.590 ;
        RECT 81.790 155.435 81.960 155.625 ;
        RECT 84.550 155.455 84.720 155.645 ;
        RECT 85.930 155.455 86.100 155.645 ;
        RECT 90.995 155.435 91.165 155.625 ;
        RECT 95.130 155.480 95.290 155.590 ;
        RECT 96.050 155.455 96.220 155.645 ;
        RECT 96.565 155.485 96.685 155.595 ;
        RECT 98.805 155.435 98.975 155.625 ;
        RECT 100.375 155.455 100.545 155.645 ;
        RECT 102.945 155.435 103.115 155.625 ;
        RECT 105.705 155.435 105.875 155.625 ;
        RECT 106.170 155.435 106.340 155.625 ;
        RECT 110.310 155.455 110.480 155.645 ;
        RECT 110.770 155.595 110.940 155.625 ;
        RECT 110.770 155.485 110.945 155.595 ;
        RECT 110.770 155.435 110.940 155.485 ;
        RECT 112.150 155.435 112.320 155.645 ;
        RECT 18.170 154.625 19.540 155.435 ;
        RECT 20.010 154.625 21.840 155.435 ;
        RECT 21.860 154.565 22.290 155.350 ;
        RECT 22.770 154.655 24.140 155.435 ;
        RECT 24.150 154.755 28.050 155.435 ;
        RECT 24.150 154.525 25.080 154.755 ;
        RECT 28.290 154.625 30.120 155.435 ;
        RECT 30.215 154.755 39.320 155.435 ;
        RECT 39.790 154.625 41.620 155.435 ;
        RECT 41.630 154.525 45.105 155.435 ;
        RECT 45.770 154.625 47.600 155.435 ;
        RECT 47.620 154.565 48.050 155.350 ;
        RECT 48.070 154.525 51.545 155.435 ;
        RECT 51.750 154.625 53.120 155.435 ;
        RECT 53.500 154.755 62.780 155.435 ;
        RECT 53.500 154.635 55.835 154.755 ;
        RECT 53.500 154.525 54.420 154.635 ;
        RECT 60.500 154.535 61.420 154.755 ;
        RECT 62.790 154.655 64.160 155.435 ;
        RECT 64.170 154.755 66.000 155.435 ;
        RECT 64.170 154.525 65.515 154.755 ;
        RECT 66.205 154.525 69.680 155.435 ;
        RECT 69.885 154.525 73.360 155.435 ;
        RECT 73.380 154.565 73.810 155.350 ;
        RECT 73.840 154.755 76.580 155.435 ;
        RECT 76.820 154.755 80.720 155.435 ;
        RECT 81.650 154.755 90.755 155.435 ;
        RECT 79.790 154.525 80.720 154.755 ;
        RECT 90.850 154.525 94.325 155.435 ;
        RECT 95.645 154.525 99.120 155.435 ;
        RECT 99.140 154.565 99.570 155.350 ;
        RECT 99.785 154.525 103.260 155.435 ;
        RECT 103.410 154.525 106.020 155.435 ;
        RECT 106.030 154.655 107.400 155.435 ;
        RECT 107.410 154.625 111.080 155.435 ;
        RECT 111.090 154.625 112.460 155.435 ;
      LAYER nwell ;
        RECT 17.975 151.405 112.655 154.235 ;
      LAYER pwell ;
        RECT 18.170 150.205 19.540 151.015 ;
        RECT 19.560 150.205 20.910 151.115 ;
        RECT 25.440 150.885 26.370 151.105 ;
        RECT 29.200 150.885 30.120 151.115 ;
        RECT 33.790 150.885 34.720 151.115 ;
        RECT 20.930 150.205 30.120 150.885 ;
        RECT 30.820 150.205 34.720 150.885 ;
        RECT 34.740 150.290 35.170 151.075 ;
        RECT 38.850 150.885 39.780 151.115 ;
        RECT 35.880 150.205 39.780 150.885 ;
        RECT 39.790 150.205 41.160 150.985 ;
        RECT 41.630 150.205 45.105 151.115 ;
        RECT 45.505 150.205 48.980 151.115 ;
        RECT 48.990 150.205 50.820 151.015 ;
        RECT 51.200 151.005 52.120 151.115 ;
        RECT 51.200 150.885 53.535 151.005 ;
        RECT 58.200 150.885 59.120 151.105 ;
        RECT 51.200 150.205 60.480 150.885 ;
        RECT 60.500 150.290 60.930 151.075 ;
        RECT 60.950 150.205 62.320 150.985 ;
        RECT 62.340 150.205 63.690 151.115 ;
        RECT 64.655 150.885 66.000 151.115 ;
        RECT 66.495 150.885 67.840 151.115 ;
        RECT 64.170 150.205 66.000 150.885 ;
        RECT 66.010 150.205 67.840 150.885 ;
        RECT 68.770 150.205 72.245 151.115 ;
        RECT 72.450 150.205 75.925 151.115 ;
        RECT 76.500 151.005 77.420 151.115 ;
        RECT 76.500 150.885 78.835 151.005 ;
        RECT 83.500 150.885 84.420 151.105 ;
        RECT 76.500 150.205 85.780 150.885 ;
        RECT 86.260 150.290 86.690 151.075 ;
        RECT 87.640 150.205 88.990 151.115 ;
        RECT 89.205 150.205 92.680 151.115 ;
        RECT 92.885 150.205 96.360 151.115 ;
        RECT 97.485 150.205 100.960 151.115 ;
        RECT 101.430 150.885 102.350 151.115 ;
        RECT 105.180 150.885 106.110 151.105 ;
        RECT 101.430 150.205 110.620 150.885 ;
        RECT 111.090 150.205 112.460 151.015 ;
        RECT 18.310 149.995 18.480 150.205 ;
        RECT 19.745 150.045 19.865 150.155 ;
        RECT 20.610 150.015 20.780 150.205 ;
        RECT 21.070 150.015 21.240 150.205 ;
        RECT 21.530 149.995 21.700 150.185 ;
        RECT 22.450 149.995 22.620 150.185 ;
        RECT 24.750 149.995 24.920 150.185 ;
        RECT 25.485 149.995 25.655 150.185 ;
        RECT 29.350 149.995 29.520 150.185 ;
        RECT 30.325 150.045 30.445 150.155 ;
        RECT 30.730 149.995 30.900 150.185 ;
        RECT 34.135 150.015 34.305 150.205 ;
        RECT 35.385 150.045 35.505 150.155 ;
        RECT 39.195 150.015 39.365 150.205 ;
        RECT 40.850 150.015 41.020 150.205 ;
        RECT 41.365 150.045 41.485 150.155 ;
        RECT 41.775 150.015 41.945 150.205 ;
        RECT 48.665 150.185 48.835 150.205 ;
        RECT 43.150 149.995 43.320 150.185 ;
        RECT 43.665 150.045 43.785 150.155 ;
        RECT 44.075 149.995 44.245 150.185 ;
        RECT 48.265 150.045 48.385 150.155 ;
        RECT 48.665 150.015 48.845 150.185 ;
        RECT 50.510 150.015 50.680 150.205 ;
        RECT 48.675 149.995 48.845 150.015 ;
        RECT 55.755 149.995 55.925 150.185 ;
        RECT 59.895 149.995 60.065 150.185 ;
        RECT 60.170 150.015 60.340 150.205 ;
        RECT 61.550 149.995 61.720 150.185 ;
        RECT 62.010 149.995 62.180 150.205 ;
        RECT 63.390 149.995 63.560 150.205 ;
        RECT 63.905 150.045 64.025 150.155 ;
        RECT 64.310 150.015 64.480 150.205 ;
        RECT 65.230 149.995 65.400 150.185 ;
        RECT 66.150 150.015 66.320 150.205 ;
        RECT 68.450 150.050 68.610 150.160 ;
        RECT 68.915 150.015 69.085 150.205 ;
        RECT 69.830 149.995 70.000 150.185 ;
        RECT 70.290 149.995 70.460 150.185 ;
        RECT 72.595 150.015 72.765 150.205 ;
        RECT 73.050 149.995 73.220 150.185 ;
        RECT 74.025 150.045 74.145 150.155 ;
        RECT 77.650 149.995 77.820 150.185 ;
        RECT 79.030 149.995 79.200 150.185 ;
        RECT 79.490 149.995 79.660 150.185 ;
        RECT 84.275 149.995 84.445 150.185 ;
        RECT 85.470 150.015 85.640 150.205 ;
        RECT 85.930 150.155 86.100 150.185 ;
        RECT 85.930 150.045 86.105 150.155 ;
        RECT 87.310 150.050 87.470 150.160 ;
        RECT 85.930 149.995 86.100 150.045 ;
        RECT 87.770 150.015 87.940 150.205 ;
        RECT 88.690 149.995 88.860 150.185 ;
        RECT 89.155 149.995 89.325 150.185 ;
        RECT 92.365 150.015 92.535 150.205 ;
        RECT 96.045 149.995 96.215 150.205 ;
        RECT 18.170 149.185 19.540 149.995 ;
        RECT 20.010 149.185 21.840 149.995 ;
        RECT 21.860 149.125 22.290 149.910 ;
        RECT 22.320 149.085 23.670 149.995 ;
        RECT 23.690 149.215 25.060 149.995 ;
        RECT 25.070 149.315 28.970 149.995 ;
        RECT 25.070 149.085 26.000 149.315 ;
        RECT 29.220 149.085 30.570 149.995 ;
        RECT 30.590 149.315 39.870 149.995 ;
        RECT 31.950 149.095 32.870 149.315 ;
        RECT 37.535 149.195 39.870 149.315 ;
        RECT 38.950 149.085 39.870 149.195 ;
        RECT 40.250 149.085 43.410 149.995 ;
        RECT 43.930 149.085 47.405 149.995 ;
        RECT 47.620 149.125 48.050 149.910 ;
        RECT 48.530 149.085 52.005 149.995 ;
        RECT 52.440 149.315 56.340 149.995 ;
        RECT 56.580 149.315 60.480 149.995 ;
        RECT 55.410 149.085 56.340 149.315 ;
        RECT 59.550 149.085 60.480 149.315 ;
        RECT 60.490 149.215 61.860 149.995 ;
        RECT 61.880 149.085 63.230 149.995 ;
        RECT 63.250 149.315 65.080 149.995 ;
        RECT 63.735 149.085 65.080 149.315 ;
        RECT 65.090 149.085 68.300 149.995 ;
        RECT 68.310 149.315 70.140 149.995 ;
        RECT 70.150 149.315 71.980 149.995 ;
        RECT 68.310 149.085 69.655 149.315 ;
        RECT 70.635 149.085 71.980 149.315 ;
        RECT 71.990 149.215 73.360 149.995 ;
        RECT 73.380 149.125 73.810 149.910 ;
        RECT 74.290 149.185 77.960 149.995 ;
        RECT 77.980 149.085 79.330 149.995 ;
        RECT 79.360 149.085 80.710 149.995 ;
        RECT 80.960 149.315 84.860 149.995 ;
        RECT 83.930 149.085 84.860 149.315 ;
        RECT 84.870 149.215 86.240 149.995 ;
        RECT 86.250 149.185 89.000 149.995 ;
        RECT 89.010 149.085 92.485 149.995 ;
        RECT 92.885 149.085 96.360 149.995 ;
        RECT 96.515 149.965 96.685 150.185 ;
        RECT 96.970 150.050 97.130 150.160 ;
        RECT 99.785 150.045 99.905 150.155 ;
        RECT 100.190 149.995 100.360 150.185 ;
        RECT 100.645 150.015 100.815 150.205 ;
        RECT 101.165 150.045 101.285 150.155 ;
        RECT 110.310 150.015 110.480 150.205 ;
        RECT 110.770 150.155 110.940 150.185 ;
        RECT 110.770 150.045 110.945 150.155 ;
        RECT 110.770 149.995 110.940 150.045 ;
        RECT 112.150 149.995 112.320 150.205 ;
        RECT 98.175 149.965 99.120 149.995 ;
        RECT 96.370 149.285 99.120 149.965 ;
        RECT 98.175 149.085 99.120 149.285 ;
        RECT 99.140 149.125 99.570 149.910 ;
        RECT 100.060 149.085 101.410 149.995 ;
        RECT 101.800 149.315 111.080 149.995 ;
        RECT 101.800 149.195 104.135 149.315 ;
        RECT 101.800 149.085 102.720 149.195 ;
        RECT 108.800 149.095 109.720 149.315 ;
        RECT 111.090 149.185 112.460 149.995 ;
      LAYER nwell ;
        RECT 17.975 145.965 112.655 148.795 ;
      LAYER pwell ;
        RECT 18.170 144.765 19.540 145.575 ;
        RECT 19.550 144.765 20.920 145.575 ;
        RECT 20.930 145.445 21.850 145.675 ;
        RECT 24.680 145.445 25.610 145.665 ;
        RECT 20.930 144.765 30.120 145.445 ;
        RECT 30.130 144.765 31.500 145.545 ;
        RECT 31.980 144.765 33.330 145.675 ;
        RECT 33.350 144.765 34.720 145.545 ;
        RECT 34.740 144.850 35.170 145.635 ;
        RECT 35.190 145.445 36.120 145.675 ;
        RECT 35.190 144.765 39.090 145.445 ;
        RECT 39.330 144.765 41.160 145.575 ;
        RECT 41.170 144.765 44.645 145.675 ;
        RECT 44.850 144.765 48.325 145.675 ;
        RECT 48.990 144.765 52.465 145.675 ;
        RECT 55.325 145.445 56.245 145.675 ;
        RECT 59.550 145.445 60.480 145.675 ;
        RECT 52.780 144.765 56.245 145.445 ;
        RECT 56.580 144.765 60.480 145.445 ;
        RECT 60.500 144.850 60.930 145.635 ;
        RECT 61.320 145.565 62.240 145.675 ;
        RECT 61.320 145.445 63.655 145.565 ;
        RECT 68.320 145.445 69.240 145.665 ;
        RECT 61.320 144.765 70.600 145.445 ;
        RECT 71.530 144.765 77.040 145.575 ;
        RECT 77.050 145.445 77.970 145.675 ;
        RECT 80.800 145.445 81.730 145.665 ;
        RECT 77.050 144.765 86.240 145.445 ;
        RECT 86.260 144.850 86.690 145.635 ;
        RECT 87.365 144.765 90.840 145.675 ;
        RECT 90.850 144.765 92.680 145.575 ;
        RECT 92.885 144.765 96.360 145.675 ;
        RECT 96.370 144.765 97.740 145.575 ;
        RECT 97.750 144.765 101.225 145.675 ;
        RECT 104.630 145.445 105.560 145.675 ;
        RECT 101.660 144.765 105.560 145.445 ;
        RECT 105.580 144.765 106.930 145.675 ;
        RECT 106.950 144.765 108.320 145.545 ;
        RECT 108.330 144.765 109.700 145.545 ;
        RECT 109.710 144.765 111.080 145.575 ;
        RECT 111.090 144.765 112.460 145.575 ;
        RECT 18.310 144.555 18.480 144.765 ;
        RECT 19.745 144.605 19.865 144.715 ;
        RECT 20.610 144.575 20.780 144.765 ;
        RECT 21.530 144.555 21.700 144.745 ;
        RECT 24.750 144.555 24.920 144.745 ;
        RECT 28.615 144.555 28.785 144.745 ;
        RECT 29.810 144.575 29.980 144.765 ;
        RECT 30.270 144.555 30.440 144.745 ;
        RECT 31.190 144.575 31.360 144.765 ;
        RECT 31.705 144.605 31.825 144.715 ;
        RECT 32.110 144.575 32.280 144.765 ;
        RECT 34.410 144.575 34.580 144.765 ;
        RECT 35.605 144.575 35.775 144.765 ;
        RECT 40.390 144.555 40.560 144.745 ;
        RECT 40.850 144.715 41.020 144.765 ;
        RECT 40.850 144.605 41.025 144.715 ;
        RECT 40.850 144.575 41.020 144.605 ;
        RECT 41.315 144.575 41.485 144.765 ;
        RECT 18.170 143.745 19.540 144.555 ;
        RECT 20.010 143.745 21.840 144.555 ;
        RECT 21.860 143.685 22.290 144.470 ;
        RECT 22.310 143.745 25.060 144.555 ;
        RECT 25.300 143.875 29.200 144.555 ;
        RECT 28.270 143.645 29.200 143.875 ;
        RECT 30.140 143.645 31.490 144.555 ;
        RECT 31.510 143.875 40.700 144.555 ;
        RECT 41.170 144.525 42.115 144.555 ;
        RECT 43.605 144.525 43.775 144.745 ;
        RECT 44.995 144.575 45.165 144.765 ;
        RECT 47.285 144.555 47.455 144.745 ;
        RECT 48.265 144.605 48.385 144.715 ;
        RECT 48.675 144.555 48.845 144.745 ;
        RECT 49.135 144.575 49.305 144.765 ;
        RECT 52.355 144.555 52.525 144.745 ;
        RECT 52.810 144.575 52.980 144.765 ;
        RECT 56.085 144.605 56.205 144.715 ;
        RECT 59.895 144.575 60.065 144.765 ;
        RECT 65.230 144.555 65.400 144.745 ;
        RECT 66.610 144.555 66.780 144.745 ;
        RECT 69.370 144.555 69.540 144.745 ;
        RECT 69.830 144.555 70.000 144.745 ;
        RECT 70.290 144.575 70.460 144.765 ;
        RECT 71.210 144.610 71.370 144.720 ;
        RECT 73.050 144.600 73.210 144.710 ;
        RECT 73.970 144.555 74.140 144.745 ;
        RECT 76.730 144.575 76.900 144.765 ;
        RECT 79.030 144.555 79.200 144.745 ;
        RECT 82.895 144.555 83.065 144.745 ;
        RECT 83.630 144.555 83.800 144.745 ;
        RECT 85.065 144.605 85.185 144.715 ;
        RECT 85.930 144.575 86.100 144.765 ;
        RECT 86.905 144.605 87.025 144.715 ;
        RECT 87.770 144.555 87.940 144.745 ;
        RECT 31.510 143.645 32.430 143.875 ;
        RECT 35.260 143.655 36.190 143.875 ;
        RECT 41.170 143.845 43.920 144.525 ;
        RECT 41.170 143.645 42.115 143.845 ;
        RECT 44.125 143.645 47.600 144.555 ;
        RECT 47.620 143.685 48.050 144.470 ;
        RECT 48.530 143.645 52.005 144.555 ;
        RECT 52.210 143.645 55.685 144.555 ;
        RECT 56.435 143.875 65.540 144.555 ;
        RECT 65.550 143.745 66.920 144.555 ;
        RECT 66.940 143.875 69.680 144.555 ;
        RECT 69.690 143.645 72.410 144.555 ;
        RECT 73.380 143.685 73.810 144.470 ;
        RECT 73.830 143.875 76.570 144.555 ;
        RECT 76.590 143.745 79.340 144.555 ;
        RECT 79.580 143.875 83.480 144.555 ;
        RECT 82.550 143.645 83.480 143.875 ;
        RECT 83.490 143.775 84.860 144.555 ;
        RECT 85.330 143.745 88.080 144.555 ;
        RECT 88.235 144.525 88.405 144.745 ;
        RECT 90.525 144.575 90.695 144.765 ;
        RECT 90.995 144.555 91.165 144.745 ;
        RECT 92.370 144.575 92.540 144.765 ;
        RECT 95.130 144.600 95.290 144.710 ;
        RECT 96.045 144.575 96.215 144.765 ;
        RECT 97.430 144.575 97.600 144.765 ;
        RECT 97.895 144.575 98.065 144.765 ;
        RECT 98.805 144.555 98.975 144.745 ;
        RECT 89.895 144.525 90.840 144.555 ;
        RECT 88.090 143.845 90.840 144.525 ;
        RECT 89.895 143.645 90.840 143.845 ;
        RECT 90.850 143.645 94.325 144.555 ;
        RECT 95.645 143.645 99.120 144.555 ;
        RECT 99.735 144.525 99.905 144.745 ;
        RECT 104.975 144.575 105.145 144.765 ;
        RECT 105.895 144.555 106.065 144.745 ;
        RECT 106.630 144.575 106.800 144.765 ;
        RECT 107.090 144.575 107.260 144.765 ;
        RECT 108.470 144.575 108.640 144.765 ;
        RECT 110.770 144.555 110.940 144.765 ;
        RECT 112.150 144.555 112.320 144.765 ;
        RECT 101.395 144.525 102.340 144.555 ;
        RECT 99.140 143.685 99.570 144.470 ;
        RECT 99.590 143.845 102.340 144.525 ;
        RECT 102.580 143.875 106.480 144.555 ;
        RECT 101.395 143.645 102.340 143.845 ;
        RECT 105.550 143.645 106.480 143.875 ;
        RECT 107.410 143.745 111.080 144.555 ;
        RECT 111.090 143.745 112.460 144.555 ;
      LAYER nwell ;
        RECT 17.975 140.525 112.655 143.355 ;
      LAYER pwell ;
        RECT 18.170 139.325 19.540 140.135 ;
        RECT 19.550 140.005 20.470 140.235 ;
        RECT 23.300 140.005 24.230 140.225 ;
        RECT 31.405 140.005 32.325 140.235 ;
        RECT 19.550 139.325 28.740 140.005 ;
        RECT 28.860 139.325 32.325 140.005 ;
        RECT 33.350 139.325 34.720 140.105 ;
        RECT 34.740 139.410 35.170 140.195 ;
        RECT 36.110 139.325 37.480 140.105 ;
        RECT 37.630 139.325 40.240 140.235 ;
        RECT 42.055 140.035 43.000 140.235 ;
        RECT 40.250 139.355 43.000 140.035 ;
        RECT 18.310 139.115 18.480 139.325 ;
        RECT 20.150 139.160 20.310 139.270 ;
        RECT 21.530 139.115 21.700 139.305 ;
        RECT 23.370 139.115 23.540 139.305 ;
        RECT 27.235 139.115 27.405 139.305 ;
        RECT 28.430 139.135 28.600 139.325 ;
        RECT 28.890 139.115 29.060 139.325 ;
        RECT 30.730 139.115 30.900 139.305 ;
        RECT 31.190 139.115 31.360 139.305 ;
        RECT 33.030 139.170 33.190 139.280 ;
        RECT 34.410 139.135 34.580 139.325 ;
        RECT 35.790 139.170 35.950 139.280 ;
        RECT 36.250 139.135 36.420 139.325 ;
        RECT 39.925 139.135 40.095 139.325 ;
        RECT 40.395 139.135 40.565 139.355 ;
        RECT 42.055 139.325 43.000 139.355 ;
        RECT 43.010 139.325 46.485 140.235 ;
        RECT 47.160 139.325 48.510 140.235 ;
        RECT 50.335 140.035 51.280 140.235 ;
        RECT 48.530 139.355 51.280 140.035 ;
        RECT 18.170 138.305 19.540 139.115 ;
        RECT 20.480 138.205 21.830 139.115 ;
        RECT 21.860 138.245 22.290 139.030 ;
        RECT 22.320 138.205 23.670 139.115 ;
        RECT 23.920 138.435 27.820 139.115 ;
        RECT 26.890 138.205 27.820 138.435 ;
        RECT 27.830 138.335 29.200 139.115 ;
        RECT 29.210 138.305 31.040 139.115 ;
        RECT 31.050 138.435 40.240 139.115 ;
        RECT 35.560 138.215 36.490 138.435 ;
        RECT 39.320 138.205 40.240 138.435 ;
        RECT 40.250 139.085 41.195 139.115 ;
        RECT 42.685 139.085 42.855 139.305 ;
        RECT 43.155 139.135 43.325 139.325 ;
        RECT 46.825 139.275 46.995 139.305 ;
        RECT 47.290 139.275 47.460 139.325 ;
        RECT 46.825 139.165 47.005 139.275 ;
        RECT 47.290 139.165 47.465 139.275 ;
        RECT 48.265 139.165 48.385 139.275 ;
        RECT 46.825 139.115 46.995 139.165 ;
        RECT 47.290 139.135 47.460 139.165 ;
        RECT 48.675 139.115 48.845 139.355 ;
        RECT 50.335 139.325 51.280 139.355 ;
        RECT 51.290 140.005 52.210 140.235 ;
        RECT 55.040 140.005 55.970 140.225 ;
        RECT 51.290 139.325 60.480 140.005 ;
        RECT 60.500 139.410 60.930 140.195 ;
        RECT 61.410 140.005 62.755 140.235 ;
        RECT 63.250 140.005 64.595 140.235 ;
        RECT 65.575 140.005 66.920 140.235 ;
        RECT 67.415 140.005 68.760 140.235 ;
        RECT 61.410 139.325 63.240 140.005 ;
        RECT 63.250 139.325 65.080 140.005 ;
        RECT 65.090 139.325 66.920 140.005 ;
        RECT 66.930 139.325 68.760 140.005 ;
        RECT 68.770 139.325 72.245 140.235 ;
        RECT 72.450 139.325 75.925 140.235 ;
        RECT 76.960 140.125 77.880 140.235 ;
        RECT 76.960 140.005 79.295 140.125 ;
        RECT 83.960 140.005 84.880 140.225 ;
        RECT 76.960 139.325 86.240 140.005 ;
        RECT 86.260 139.410 86.690 140.195 ;
        RECT 86.710 139.325 88.080 140.135 ;
        RECT 88.090 140.035 89.035 140.235 ;
        RECT 88.090 139.355 90.840 140.035 ;
        RECT 88.090 139.325 89.035 139.355 ;
        RECT 60.170 139.135 60.340 139.325 ;
        RECT 61.145 139.165 61.265 139.275 ;
        RECT 61.550 139.115 61.720 139.305 ;
        RECT 62.930 139.115 63.100 139.325 ;
        RECT 64.770 139.115 64.940 139.325 ;
        RECT 65.230 139.115 65.400 139.325 ;
        RECT 67.070 139.115 67.240 139.325 ;
        RECT 68.915 139.135 69.085 139.325 ;
        RECT 69.370 139.160 69.530 139.270 ;
        RECT 69.835 139.115 70.005 139.305 ;
        RECT 72.595 139.135 72.765 139.325 ;
        RECT 73.975 139.115 74.145 139.305 ;
        RECT 76.325 139.165 76.445 139.275 ;
        RECT 77.705 139.165 77.825 139.275 ;
        RECT 79.490 139.115 79.660 139.305 ;
        RECT 83.355 139.115 83.525 139.305 ;
        RECT 85.010 139.115 85.180 139.305 ;
        RECT 85.930 139.135 86.100 139.325 ;
        RECT 86.390 139.115 86.560 139.305 ;
        RECT 87.770 139.115 87.940 139.325 ;
        RECT 90.525 139.135 90.695 139.355 ;
        RECT 90.850 139.325 94.325 140.235 ;
        RECT 94.530 139.325 95.900 140.135 ;
        RECT 95.910 139.325 99.385 140.235 ;
        RECT 101.395 140.035 102.340 140.235 ;
        RECT 99.590 139.355 102.340 140.035 ;
        RECT 105.550 140.005 106.480 140.235 ;
        RECT 90.995 139.135 91.165 139.325 ;
        RECT 93.290 139.115 93.460 139.305 ;
        RECT 40.250 138.405 43.000 139.085 ;
        RECT 40.250 138.205 41.195 138.405 ;
        RECT 43.665 138.205 47.140 139.115 ;
        RECT 47.620 138.245 48.050 139.030 ;
        RECT 48.530 138.205 52.005 139.115 ;
        RECT 52.580 138.435 61.860 139.115 ;
        RECT 52.580 138.315 54.915 138.435 ;
        RECT 52.580 138.205 53.500 138.315 ;
        RECT 59.580 138.215 60.500 138.435 ;
        RECT 61.870 138.335 63.240 139.115 ;
        RECT 63.250 138.435 65.080 139.115 ;
        RECT 65.090 138.435 66.920 139.115 ;
        RECT 66.930 138.435 68.760 139.115 ;
        RECT 63.250 138.205 64.595 138.435 ;
        RECT 65.575 138.205 66.920 138.435 ;
        RECT 67.415 138.205 68.760 138.435 ;
        RECT 69.690 138.205 73.165 139.115 ;
        RECT 73.380 138.245 73.810 139.030 ;
        RECT 73.830 138.205 77.305 139.115 ;
        RECT 77.970 138.305 79.800 139.115 ;
        RECT 80.040 138.435 83.940 139.115 ;
        RECT 83.010 138.205 83.940 138.435 ;
        RECT 83.960 138.205 85.310 139.115 ;
        RECT 85.330 138.335 86.700 139.115 ;
        RECT 86.710 138.305 88.080 139.115 ;
        RECT 88.090 138.305 93.600 139.115 ;
        RECT 93.755 139.085 93.925 139.305 ;
        RECT 95.590 139.135 95.760 139.325 ;
        RECT 96.055 139.135 96.225 139.325 ;
        RECT 96.515 139.115 96.685 139.305 ;
        RECT 99.735 139.135 99.905 139.355 ;
        RECT 101.395 139.325 102.340 139.355 ;
        RECT 102.580 139.325 106.480 140.005 ;
        RECT 106.500 139.325 107.850 140.235 ;
        RECT 107.870 139.325 109.240 140.105 ;
        RECT 109.250 139.325 111.080 140.135 ;
        RECT 111.090 139.325 112.460 140.135 ;
        RECT 100.190 139.115 100.360 139.305 ;
        RECT 105.895 139.135 106.065 139.325 ;
        RECT 106.630 139.135 106.800 139.325 ;
        RECT 108.010 139.135 108.180 139.325 ;
        RECT 110.770 139.115 110.940 139.325 ;
        RECT 112.150 139.115 112.320 139.325 ;
        RECT 95.415 139.085 96.360 139.115 ;
        RECT 93.610 138.405 96.360 139.085 ;
        RECT 95.415 138.205 96.360 138.405 ;
        RECT 96.370 138.205 98.980 139.115 ;
        RECT 99.140 138.245 99.570 139.030 ;
        RECT 100.060 138.205 101.410 139.115 ;
        RECT 101.800 138.435 111.080 139.115 ;
        RECT 101.800 138.315 104.135 138.435 ;
        RECT 101.800 138.205 102.720 138.315 ;
        RECT 108.800 138.215 109.720 138.435 ;
        RECT 111.090 138.305 112.460 139.115 ;
      LAYER nwell ;
        RECT 17.975 135.085 112.655 137.915 ;
      LAYER pwell ;
        RECT 18.170 133.885 19.540 134.695 ;
        RECT 20.010 134.565 20.930 134.795 ;
        RECT 23.760 134.565 24.690 134.785 ;
        RECT 20.010 133.885 29.200 134.565 ;
        RECT 29.220 133.885 30.570 134.795 ;
        RECT 33.790 134.565 34.720 134.795 ;
        RECT 30.820 133.885 34.720 134.565 ;
        RECT 34.740 133.970 35.170 134.755 ;
        RECT 35.190 134.565 36.120 134.795 ;
        RECT 39.790 134.595 40.735 134.795 ;
        RECT 35.190 133.885 39.090 134.565 ;
        RECT 39.790 133.915 42.540 134.595 ;
        RECT 39.790 133.885 40.735 133.915 ;
        RECT 18.310 133.675 18.480 133.885 ;
        RECT 19.745 133.725 19.865 133.835 ;
        RECT 21.530 133.675 21.700 133.865 ;
        RECT 22.505 133.725 22.625 133.835 ;
        RECT 22.910 133.675 23.080 133.865 ;
        RECT 24.290 133.675 24.460 133.865 ;
        RECT 28.890 133.695 29.060 133.885 ;
        RECT 29.350 133.695 29.520 133.885 ;
        RECT 34.135 133.695 34.305 133.885 ;
        RECT 34.410 133.675 34.580 133.865 ;
        RECT 35.605 133.695 35.775 133.885 ;
        RECT 35.790 133.675 35.960 133.865 ;
        RECT 37.630 133.675 37.800 133.865 ;
        RECT 38.090 133.695 38.260 133.865 ;
        RECT 39.525 133.725 39.645 133.835 ;
        RECT 38.110 133.675 38.260 133.695 ;
        RECT 18.170 132.865 19.540 133.675 ;
        RECT 20.010 132.865 21.840 133.675 ;
        RECT 21.860 132.805 22.290 133.590 ;
        RECT 22.780 132.765 24.130 133.675 ;
        RECT 24.150 132.895 25.520 133.675 ;
        RECT 25.530 132.995 34.720 133.675 ;
        RECT 25.530 132.765 26.450 132.995 ;
        RECT 29.280 132.775 30.210 132.995 ;
        RECT 34.730 132.895 36.100 133.675 ;
        RECT 36.110 132.865 37.940 133.675 ;
        RECT 38.110 132.855 40.040 133.675 ;
        RECT 40.395 133.645 40.565 133.865 ;
        RECT 42.225 133.695 42.395 133.915 ;
        RECT 42.550 133.885 46.025 134.795 ;
        RECT 46.230 133.885 49.705 134.795 ;
        RECT 50.370 133.885 53.845 134.795 ;
        RECT 54.980 133.885 56.330 134.795 ;
        RECT 59.550 134.565 60.480 134.795 ;
        RECT 56.580 133.885 60.480 134.565 ;
        RECT 60.500 133.970 60.930 134.755 ;
        RECT 61.870 133.885 63.240 134.665 ;
        RECT 63.260 133.885 64.610 134.795 ;
        RECT 64.630 133.885 66.000 134.665 ;
        RECT 66.470 133.885 67.840 134.665 ;
        RECT 67.850 133.885 71.520 134.695 ;
        RECT 71.530 134.595 72.475 134.795 ;
        RECT 71.530 133.915 74.280 134.595 ;
        RECT 71.530 133.885 72.475 133.915 ;
        RECT 42.695 133.695 42.865 133.885 ;
        RECT 43.155 133.675 43.325 133.865 ;
        RECT 46.375 133.695 46.545 133.885 ;
        RECT 47.290 133.720 47.450 133.830 ;
        RECT 50.105 133.725 50.225 133.835 ;
        RECT 50.515 133.695 50.685 133.885 ;
        RECT 51.430 133.675 51.600 133.865 ;
        RECT 51.895 133.675 52.065 133.865 ;
        RECT 54.650 133.730 54.810 133.840 ;
        RECT 55.110 133.695 55.280 133.885 ;
        RECT 58.975 133.675 59.145 133.865 ;
        RECT 59.895 133.695 60.065 133.885 ;
        RECT 61.550 133.730 61.710 133.840 ;
        RECT 62.930 133.695 63.100 133.885 ;
        RECT 64.310 133.695 64.480 133.885 ;
        RECT 64.770 133.695 64.940 133.885 ;
        RECT 66.205 133.725 66.325 133.835 ;
        RECT 66.610 133.695 66.780 133.885 ;
        RECT 68.910 133.675 69.080 133.865 ;
        RECT 70.290 133.675 70.460 133.865 ;
        RECT 42.055 133.645 43.000 133.675 ;
        RECT 40.250 132.965 43.000 133.645 ;
        RECT 39.090 132.765 40.040 132.855 ;
        RECT 42.055 132.765 43.000 132.965 ;
        RECT 43.010 132.765 46.485 133.675 ;
        RECT 47.620 132.805 48.050 133.590 ;
        RECT 48.070 132.865 51.740 133.675 ;
        RECT 51.750 132.765 55.225 133.675 ;
        RECT 55.660 132.995 59.560 133.675 ;
        RECT 58.630 132.765 59.560 132.995 ;
        RECT 59.940 132.995 69.220 133.675 ;
        RECT 59.940 132.875 62.275 132.995 ;
        RECT 59.940 132.765 60.860 132.875 ;
        RECT 66.940 132.775 67.860 132.995 ;
        RECT 69.230 132.895 70.600 133.675 ;
        RECT 70.755 133.645 70.925 133.865 ;
        RECT 71.210 133.695 71.380 133.885 ;
        RECT 73.965 133.835 74.135 133.915 ;
        RECT 74.290 133.885 77.765 134.795 ;
        RECT 78.430 133.885 80.260 134.695 ;
        RECT 83.470 134.565 84.400 134.795 ;
        RECT 80.500 133.885 84.400 134.565 ;
        RECT 84.870 133.885 86.240 134.665 ;
        RECT 86.260 133.970 86.690 134.755 ;
        RECT 87.170 133.885 89.920 134.695 ;
        RECT 89.940 133.885 91.290 134.795 ;
        RECT 94.510 134.565 95.440 134.795 ;
        RECT 99.110 134.565 100.040 134.795 ;
        RECT 91.540 133.885 95.440 134.565 ;
        RECT 96.140 133.885 100.040 134.565 ;
        RECT 101.340 134.685 102.260 134.795 ;
        RECT 101.340 134.565 103.675 134.685 ;
        RECT 108.340 134.565 109.260 134.785 ;
        RECT 101.340 133.885 110.620 134.565 ;
        RECT 111.090 133.885 112.460 134.695 ;
        RECT 73.965 133.725 74.145 133.835 ;
        RECT 73.965 133.695 74.135 133.725 ;
        RECT 74.435 133.675 74.605 133.885 ;
        RECT 78.165 133.725 78.285 133.835 ;
        RECT 79.030 133.675 79.200 133.865 ;
        RECT 79.950 133.695 80.120 133.885 ;
        RECT 83.815 133.695 83.985 133.885 ;
        RECT 84.605 133.725 84.725 133.835 ;
        RECT 85.010 133.695 85.180 133.885 ;
        RECT 86.905 133.725 87.025 133.835 ;
        RECT 88.690 133.675 88.860 133.865 ;
        RECT 89.205 133.725 89.325 133.835 ;
        RECT 89.610 133.695 89.780 133.885 ;
        RECT 90.070 133.695 90.240 133.885 ;
        RECT 94.855 133.695 95.025 133.885 ;
        RECT 95.645 133.725 95.765 133.835 ;
        RECT 98.810 133.675 98.980 133.865 ;
        RECT 99.455 133.695 99.625 133.885 ;
        RECT 100.650 133.675 100.820 133.865 ;
        RECT 101.165 133.725 101.285 133.835 ;
        RECT 104.975 133.675 105.145 133.865 ;
        RECT 106.170 133.720 106.330 133.830 ;
        RECT 106.630 133.675 106.800 133.865 ;
        RECT 108.065 133.725 108.185 133.835 ;
        RECT 110.310 133.695 110.480 133.885 ;
        RECT 110.770 133.835 110.940 133.865 ;
        RECT 110.770 133.725 110.945 133.835 ;
        RECT 110.770 133.675 110.940 133.725 ;
        RECT 112.150 133.675 112.320 133.885 ;
        RECT 72.415 133.645 73.360 133.675 ;
        RECT 70.610 132.965 73.360 133.645 ;
        RECT 72.415 132.765 73.360 132.965 ;
        RECT 73.380 132.805 73.810 133.590 ;
        RECT 74.290 132.765 77.765 133.675 ;
        RECT 77.980 132.765 79.330 133.675 ;
        RECT 79.720 132.995 89.000 133.675 ;
        RECT 89.840 132.995 99.120 133.675 ;
        RECT 79.720 132.875 82.055 132.995 ;
        RECT 79.720 132.765 80.640 132.875 ;
        RECT 86.720 132.775 87.640 132.995 ;
        RECT 89.840 132.875 92.175 132.995 ;
        RECT 89.840 132.765 90.760 132.875 ;
        RECT 96.840 132.775 97.760 132.995 ;
        RECT 99.140 132.805 99.570 133.590 ;
        RECT 99.600 132.765 100.950 133.675 ;
        RECT 101.660 132.995 105.560 133.675 ;
        RECT 104.630 132.765 105.560 132.995 ;
        RECT 106.490 132.895 107.860 133.675 ;
        RECT 108.330 132.865 111.080 133.675 ;
        RECT 111.090 132.865 112.460 133.675 ;
      LAYER nwell ;
        RECT 17.975 129.645 112.655 132.475 ;
      LAYER pwell ;
        RECT 18.170 128.445 19.540 129.255 ;
        RECT 22.205 129.125 23.125 129.355 ;
        RECT 19.660 128.445 23.125 129.125 ;
        RECT 23.230 128.445 24.600 129.255 ;
        RECT 24.610 129.125 25.540 129.355 ;
        RECT 24.610 128.445 28.510 129.125 ;
        RECT 28.750 128.445 30.120 129.255 ;
        RECT 30.140 128.445 31.490 129.355 ;
        RECT 31.970 128.445 34.720 129.255 ;
        RECT 34.740 128.530 35.170 129.315 ;
        RECT 38.170 129.265 39.120 129.355 ;
        RECT 35.650 128.445 37.020 129.225 ;
        RECT 37.190 128.445 39.120 129.265 ;
        RECT 41.135 129.155 42.080 129.355 ;
        RECT 43.895 129.155 44.840 129.355 ;
        RECT 39.330 128.475 42.080 129.155 ;
        RECT 42.090 128.475 44.840 129.155 ;
        RECT 18.310 128.235 18.480 128.445 ;
        RECT 19.690 128.255 19.860 128.445 ;
        RECT 20.150 128.280 20.310 128.390 ;
        RECT 21.530 128.235 21.700 128.425 ;
        RECT 24.290 128.255 24.460 128.445 ;
        RECT 25.025 128.255 25.195 128.445 ;
        RECT 29.810 128.255 29.980 128.445 ;
        RECT 31.190 128.255 31.360 128.445 ;
        RECT 31.650 128.395 31.820 128.425 ;
        RECT 31.650 128.285 31.825 128.395 ;
        RECT 31.650 128.235 31.820 128.285 ;
        RECT 34.410 128.255 34.580 128.445 ;
        RECT 35.385 128.285 35.505 128.395 ;
        RECT 35.515 128.235 35.685 128.425 ;
        RECT 36.305 128.285 36.425 128.395 ;
        RECT 36.710 128.235 36.880 128.445 ;
        RECT 37.190 128.425 37.340 128.445 ;
        RECT 37.170 128.255 37.340 128.425 ;
        RECT 38.365 128.235 38.535 128.425 ;
        RECT 39.475 128.255 39.645 128.475 ;
        RECT 41.135 128.445 42.080 128.475 ;
        RECT 42.235 128.255 42.405 128.475 ;
        RECT 43.895 128.445 44.840 128.475 ;
        RECT 44.850 129.155 45.795 129.355 ;
        RECT 44.850 128.475 47.600 129.155 ;
        RECT 44.850 128.445 45.795 128.475 ;
        RECT 42.690 128.255 42.860 128.425 ;
        RECT 42.710 128.235 42.860 128.255 ;
        RECT 18.170 127.425 19.540 128.235 ;
        RECT 20.480 127.325 21.830 128.235 ;
        RECT 21.860 127.365 22.290 128.150 ;
        RECT 22.680 127.555 31.960 128.235 ;
        RECT 32.200 127.555 36.100 128.235 ;
        RECT 22.680 127.435 25.015 127.555 ;
        RECT 22.680 127.325 23.600 127.435 ;
        RECT 29.680 127.335 30.600 127.555 ;
        RECT 35.170 127.325 36.100 127.555 ;
        RECT 36.570 127.455 37.940 128.235 ;
        RECT 37.950 127.555 41.850 128.235 ;
        RECT 37.950 127.325 38.880 127.555 ;
        RECT 42.710 127.415 44.640 128.235 ;
        RECT 43.690 127.325 44.640 127.415 ;
        RECT 44.850 128.205 45.795 128.235 ;
        RECT 47.285 128.205 47.455 128.475 ;
        RECT 48.070 128.445 51.545 129.355 ;
        RECT 51.750 128.445 55.225 129.355 ;
        RECT 59.550 129.125 60.480 129.355 ;
        RECT 56.580 128.445 60.480 129.125 ;
        RECT 60.500 128.530 60.930 129.315 ;
        RECT 61.320 129.245 62.240 129.355 ;
        RECT 61.320 129.125 63.655 129.245 ;
        RECT 68.320 129.125 69.240 129.345 ;
        RECT 70.810 129.265 71.760 129.355 ;
        RECT 61.320 128.445 70.600 129.125 ;
        RECT 70.810 128.445 72.740 129.265 ;
        RECT 72.910 128.445 76.385 129.355 ;
        RECT 76.960 129.245 77.880 129.355 ;
        RECT 76.960 129.125 79.295 129.245 ;
        RECT 83.960 129.125 84.880 129.345 ;
        RECT 76.960 128.445 86.240 129.125 ;
        RECT 86.260 128.530 86.690 129.315 ;
        RECT 86.720 128.445 88.070 129.355 ;
        RECT 88.460 129.245 89.380 129.355 ;
        RECT 88.460 129.125 90.795 129.245 ;
        RECT 95.460 129.125 96.380 129.345 ;
        RECT 88.460 128.445 97.740 129.125 ;
        RECT 97.750 128.445 99.120 129.225 ;
        RECT 99.590 128.445 100.960 129.225 ;
        RECT 101.890 128.445 105.560 129.255 ;
        RECT 105.570 128.445 111.080 129.255 ;
        RECT 111.090 128.445 112.460 129.255 ;
        RECT 47.805 128.285 47.925 128.395 ;
        RECT 48.215 128.255 48.385 128.445 ;
        RECT 48.670 128.280 48.830 128.390 ;
        RECT 51.430 128.235 51.600 128.425 ;
        RECT 51.895 128.235 52.065 128.445 ;
        RECT 56.030 128.290 56.190 128.400 ;
        RECT 59.895 128.255 60.065 128.445 ;
        RECT 64.770 128.235 64.940 128.425 ;
        RECT 65.230 128.235 65.400 128.425 ;
        RECT 44.850 127.525 47.600 128.205 ;
        RECT 44.850 127.325 45.795 127.525 ;
        RECT 47.620 127.365 48.050 128.150 ;
        RECT 49.000 127.555 51.740 128.235 ;
        RECT 51.750 127.325 55.225 128.235 ;
        RECT 55.800 127.555 65.080 128.235 ;
        RECT 65.090 127.555 66.920 128.235 ;
        RECT 66.930 128.205 67.875 128.235 ;
        RECT 69.365 128.205 69.535 128.425 ;
        RECT 69.835 128.235 70.005 128.425 ;
        RECT 70.290 128.255 70.460 128.445 ;
        RECT 72.590 128.425 72.740 128.445 ;
        RECT 72.590 128.255 72.760 128.425 ;
        RECT 73.055 128.255 73.225 128.445 ;
        RECT 74.430 128.280 74.590 128.390 ;
        RECT 76.730 128.255 76.900 128.425 ;
        RECT 76.730 128.235 76.880 128.255 ;
        RECT 80.595 128.235 80.765 128.425 ;
        RECT 81.385 128.285 81.505 128.395 ;
        RECT 81.790 128.235 81.960 128.425 ;
        RECT 85.930 128.255 86.100 128.445 ;
        RECT 87.770 128.255 87.940 128.445 ;
        RECT 91.910 128.235 92.080 128.425 ;
        RECT 92.425 128.285 92.545 128.395 ;
        RECT 94.210 128.235 94.380 128.425 ;
        RECT 94.670 128.255 94.840 128.425 ;
        RECT 96.970 128.255 97.140 128.425 ;
        RECT 97.430 128.255 97.600 128.445 ;
        RECT 98.810 128.255 98.980 128.445 ;
        RECT 99.325 128.285 99.445 128.395 ;
        RECT 94.690 128.235 94.840 128.255 ;
        RECT 96.990 128.235 97.140 128.255 ;
        RECT 100.650 128.235 100.820 128.445 ;
        RECT 101.570 128.290 101.730 128.400 ;
        RECT 104.330 128.235 104.500 128.425 ;
        RECT 104.790 128.235 104.960 128.425 ;
        RECT 105.250 128.255 105.420 128.445 ;
        RECT 106.630 128.280 106.790 128.390 ;
        RECT 107.090 128.235 107.260 128.425 ;
        RECT 110.770 128.235 110.940 128.445 ;
        RECT 112.150 128.235 112.320 128.445 ;
        RECT 55.800 127.435 58.135 127.555 ;
        RECT 55.800 127.325 56.720 127.435 ;
        RECT 62.800 127.335 63.720 127.555 ;
        RECT 66.930 127.525 69.680 128.205 ;
        RECT 66.930 127.325 67.875 127.525 ;
        RECT 69.690 127.325 73.165 128.235 ;
        RECT 73.380 127.365 73.810 128.150 ;
        RECT 74.950 127.415 76.880 128.235 ;
        RECT 77.280 127.555 81.180 128.235 ;
        RECT 81.650 127.555 90.755 128.235 ;
        RECT 74.950 127.325 75.900 127.415 ;
        RECT 80.250 127.325 81.180 127.555 ;
        RECT 90.850 127.455 92.220 128.235 ;
        RECT 92.690 127.425 94.520 128.235 ;
        RECT 94.690 127.415 96.620 128.235 ;
        RECT 96.990 127.415 98.920 128.235 ;
        RECT 95.670 127.325 96.620 127.415 ;
        RECT 97.970 127.325 98.920 127.415 ;
        RECT 99.140 127.365 99.570 128.150 ;
        RECT 99.590 127.425 100.960 128.235 ;
        RECT 100.970 127.425 104.640 128.235 ;
        RECT 104.660 127.325 106.010 128.235 ;
        RECT 106.950 127.455 108.320 128.235 ;
        RECT 108.330 127.425 111.080 128.235 ;
        RECT 111.090 127.425 112.460 128.235 ;
      LAYER nwell ;
        RECT 17.975 124.205 112.655 127.035 ;
      LAYER pwell ;
        RECT 18.170 123.005 19.540 123.815 ;
        RECT 19.550 123.005 20.920 123.785 ;
        RECT 20.930 123.685 21.860 123.915 ;
        RECT 25.440 123.805 26.360 123.915 ;
        RECT 25.440 123.685 27.775 123.805 ;
        RECT 32.440 123.685 33.360 123.905 ;
        RECT 20.930 123.005 24.830 123.685 ;
        RECT 25.440 123.005 34.720 123.685 ;
        RECT 34.740 123.090 35.170 123.875 ;
        RECT 44.590 123.825 45.540 123.915 ;
        RECT 46.890 123.825 47.840 123.915 ;
        RECT 35.275 123.005 44.380 123.685 ;
        RECT 44.590 123.005 46.520 123.825 ;
        RECT 46.890 123.005 48.820 123.825 ;
        RECT 48.990 123.685 49.920 123.915 ;
        RECT 48.990 123.005 52.890 123.685 ;
        RECT 53.130 123.005 56.290 123.915 ;
        RECT 56.350 123.685 57.280 123.915 ;
        RECT 56.350 123.005 60.250 123.685 ;
        RECT 60.500 123.090 60.930 123.875 ;
        RECT 61.610 123.825 62.560 123.915 ;
        RECT 64.850 123.825 65.800 123.915 ;
        RECT 61.610 123.005 63.540 123.825 ;
        RECT 18.310 122.795 18.480 123.005 ;
        RECT 19.690 122.815 19.860 123.005 ;
        RECT 20.150 122.840 20.310 122.950 ;
        RECT 20.610 122.795 20.780 122.985 ;
        RECT 21.345 122.815 21.515 123.005 ;
        RECT 31.650 122.795 31.820 122.985 ;
        RECT 34.410 122.815 34.580 123.005 ;
        RECT 41.310 122.795 41.480 122.985 ;
        RECT 42.690 122.815 42.860 122.985 ;
        RECT 43.205 122.845 43.325 122.955 ;
        RECT 44.070 122.815 44.240 123.005 ;
        RECT 46.370 122.985 46.520 123.005 ;
        RECT 48.670 122.985 48.820 123.005 ;
        RECT 45.450 122.815 45.620 122.985 ;
        RECT 45.965 122.845 46.085 122.955 ;
        RECT 45.450 122.795 45.600 122.815 ;
        RECT 46.370 122.795 46.540 122.985 ;
        RECT 48.210 122.795 48.380 122.985 ;
        RECT 48.670 122.815 48.840 122.985 ;
        RECT 49.405 122.815 49.575 123.005 ;
        RECT 56.030 122.815 56.200 123.005 ;
        RECT 56.765 122.815 56.935 123.005 ;
        RECT 63.390 122.985 63.540 123.005 ;
        RECT 63.870 123.005 65.800 123.825 ;
        RECT 66.010 123.715 66.955 123.915 ;
        RECT 66.010 123.035 68.760 123.715 ;
        RECT 66.010 123.005 66.955 123.035 ;
        RECT 63.870 122.985 64.020 123.005 ;
        RECT 57.465 122.845 57.585 122.955 ;
        RECT 61.145 122.845 61.265 122.955 ;
        RECT 63.390 122.815 63.560 122.985 ;
        RECT 63.850 122.815 64.020 122.985 ;
        RECT 67.070 122.795 67.240 122.985 ;
        RECT 67.530 122.795 67.700 122.985 ;
        RECT 68.445 122.815 68.615 123.035 ;
        RECT 68.770 123.005 71.510 123.685 ;
        RECT 71.615 123.005 80.720 123.685 ;
        RECT 80.730 123.005 82.100 123.785 ;
        RECT 85.310 123.685 86.240 123.915 ;
        RECT 82.340 123.005 86.240 123.685 ;
        RECT 86.260 123.090 86.690 123.875 ;
        RECT 88.310 123.825 89.260 123.915 ;
        RECT 87.330 123.005 89.260 123.825 ;
        RECT 89.670 123.825 90.620 123.915 ;
        RECT 93.370 123.825 94.320 123.915 ;
        RECT 89.670 123.005 91.600 123.825 ;
        RECT 68.910 122.815 69.080 123.005 ;
        RECT 72.775 122.795 72.945 122.985 ;
        RECT 76.730 122.815 76.900 122.985 ;
        RECT 77.190 122.795 77.360 122.985 ;
        RECT 80.410 122.815 80.580 123.005 ;
        RECT 81.790 122.815 81.960 123.005 ;
        RECT 85.655 122.815 85.825 123.005 ;
        RECT 87.330 122.985 87.480 123.005 ;
        RECT 91.450 122.985 91.600 123.005 ;
        RECT 92.390 123.005 94.320 123.825 ;
        RECT 94.730 123.825 95.680 123.915 ;
        RECT 94.730 123.005 96.660 123.825 ;
        RECT 100.490 123.685 101.420 123.915 ;
        RECT 97.520 123.005 101.420 123.685 ;
        RECT 101.800 123.805 102.720 123.915 ;
        RECT 101.800 123.685 104.135 123.805 ;
        RECT 108.800 123.685 109.720 123.905 ;
        RECT 101.800 123.005 111.080 123.685 ;
        RECT 111.090 123.005 112.460 123.815 ;
        RECT 92.390 122.985 92.540 123.005 ;
        RECT 96.510 122.985 96.660 123.005 ;
        RECT 86.905 122.845 87.025 122.955 ;
        RECT 87.310 122.815 87.480 122.985 ;
        RECT 87.770 122.795 87.940 122.985 ;
        RECT 91.450 122.815 91.620 122.985 ;
        RECT 91.635 122.795 91.805 122.985 ;
        RECT 91.965 122.845 92.085 122.955 ;
        RECT 92.370 122.815 92.540 122.985 ;
        RECT 93.290 122.795 93.460 122.985 ;
        RECT 93.750 122.795 93.920 122.985 ;
        RECT 96.510 122.815 96.680 122.985 ;
        RECT 97.025 122.845 97.145 122.955 ;
        RECT 98.535 122.795 98.705 122.985 ;
        RECT 100.650 122.795 100.820 122.985 ;
        RECT 100.835 122.815 101.005 123.005 ;
        RECT 110.310 122.795 110.480 122.985 ;
        RECT 110.770 122.955 110.940 123.005 ;
        RECT 110.770 122.845 110.945 122.955 ;
        RECT 110.770 122.815 110.940 122.845 ;
        RECT 112.150 122.795 112.320 123.005 ;
        RECT 18.170 121.985 19.540 122.795 ;
        RECT 20.470 122.015 21.840 122.795 ;
        RECT 21.860 121.925 22.290 122.710 ;
        RECT 22.680 122.115 31.960 122.795 ;
        RECT 32.340 122.115 41.620 122.795 ;
        RECT 41.630 122.115 42.585 122.795 ;
        RECT 22.680 121.995 25.015 122.115 ;
        RECT 22.680 121.885 23.600 121.995 ;
        RECT 29.680 121.895 30.600 122.115 ;
        RECT 32.340 121.995 34.675 122.115 ;
        RECT 32.340 121.885 33.260 121.995 ;
        RECT 39.340 121.895 40.260 122.115 ;
        RECT 43.670 121.975 45.600 122.795 ;
        RECT 46.230 122.015 47.600 122.795 ;
        RECT 43.670 121.885 44.620 121.975 ;
        RECT 47.620 121.925 48.050 122.710 ;
        RECT 48.070 122.115 57.175 122.795 ;
        RECT 58.100 122.115 67.380 122.795 ;
        RECT 67.390 122.115 69.220 122.795 ;
        RECT 69.460 122.115 73.360 122.795 ;
        RECT 58.100 121.995 60.435 122.115 ;
        RECT 58.100 121.885 59.020 121.995 ;
        RECT 65.100 121.895 66.020 122.115 ;
        RECT 72.430 121.885 73.360 122.115 ;
        RECT 73.380 121.925 73.810 122.710 ;
        RECT 74.210 122.115 76.635 122.795 ;
        RECT 77.050 122.115 86.330 122.795 ;
        RECT 78.410 121.895 79.330 122.115 ;
        RECT 83.995 121.995 86.330 122.115 ;
        RECT 85.410 121.885 86.330 121.995 ;
        RECT 86.710 121.985 88.080 122.795 ;
        RECT 88.320 122.115 92.220 122.795 ;
        RECT 91.290 121.885 92.220 122.115 ;
        RECT 92.240 121.885 93.590 122.795 ;
        RECT 93.610 122.015 94.980 122.795 ;
        RECT 95.220 122.115 99.120 122.795 ;
        RECT 98.190 121.885 99.120 122.115 ;
        RECT 99.140 121.925 99.570 122.710 ;
        RECT 99.600 121.885 100.950 122.795 ;
        RECT 101.340 122.115 110.620 122.795 ;
        RECT 101.340 121.995 103.675 122.115 ;
        RECT 101.340 121.885 102.260 121.995 ;
        RECT 108.340 121.895 109.260 122.115 ;
        RECT 111.090 121.985 112.460 122.795 ;
      LAYER nwell ;
        RECT 17.975 118.765 112.655 121.595 ;
      LAYER pwell ;
        RECT 18.170 117.565 19.540 118.375 ;
        RECT 19.550 117.565 21.380 118.375 ;
        RECT 21.400 117.565 22.750 118.475 ;
        RECT 22.770 118.245 23.700 118.475 ;
        RECT 30.110 118.245 31.040 118.475 ;
        RECT 22.770 117.565 26.670 118.245 ;
        RECT 27.140 117.565 31.040 118.245 ;
        RECT 31.060 117.565 32.410 118.475 ;
        RECT 33.570 118.385 34.520 118.475 ;
        RECT 32.590 117.565 34.520 118.385 ;
        RECT 34.740 117.650 35.170 118.435 ;
        RECT 36.790 118.385 37.740 118.475 ;
        RECT 40.010 118.385 40.960 118.475 ;
        RECT 35.810 117.565 37.740 118.385 ;
        RECT 39.030 117.565 40.960 118.385 ;
        RECT 41.370 118.385 42.320 118.475 ;
        RECT 41.370 117.565 43.300 118.385 ;
        RECT 46.670 118.245 47.600 118.475 ;
        RECT 51.270 118.245 52.200 118.475 ;
        RECT 43.700 117.565 47.600 118.245 ;
        RECT 48.300 117.565 52.200 118.245 ;
        RECT 52.210 117.565 53.580 118.345 ;
        RECT 53.590 117.565 54.960 118.345 ;
        RECT 54.980 117.565 56.330 118.475 ;
        RECT 59.550 118.245 60.480 118.475 ;
        RECT 56.580 117.565 60.480 118.245 ;
        RECT 60.500 117.650 60.930 118.435 ;
        RECT 60.950 118.245 61.880 118.475 ;
        RECT 60.950 117.565 64.850 118.245 ;
        RECT 65.100 117.565 66.450 118.475 ;
        RECT 66.480 117.565 67.830 118.475 ;
        RECT 69.140 118.365 70.060 118.475 ;
        RECT 69.140 118.245 71.475 118.365 ;
        RECT 76.140 118.245 77.060 118.465 ;
        RECT 78.630 118.385 79.580 118.475 ;
        RECT 69.140 117.565 78.420 118.245 ;
        RECT 78.630 117.565 80.560 118.385 ;
        RECT 80.730 117.565 82.100 118.345 ;
        RECT 85.310 118.245 86.240 118.475 ;
        RECT 82.340 117.565 86.240 118.245 ;
        RECT 86.260 117.650 86.690 118.435 ;
        RECT 88.000 118.365 88.920 118.475 ;
        RECT 88.000 118.245 90.335 118.365 ;
        RECT 95.000 118.245 95.920 118.465 ;
        RECT 100.490 118.245 101.420 118.475 ;
        RECT 104.630 118.245 105.560 118.475 ;
        RECT 88.000 117.565 97.280 118.245 ;
        RECT 97.520 117.565 101.420 118.245 ;
        RECT 101.660 117.565 105.560 118.245 ;
        RECT 105.580 117.565 106.930 118.475 ;
        RECT 106.950 117.565 108.320 118.345 ;
        RECT 108.330 117.565 111.080 118.375 ;
        RECT 111.090 117.565 112.460 118.375 ;
        RECT 18.310 117.355 18.480 117.565 ;
        RECT 20.150 117.400 20.310 117.510 ;
        RECT 21.070 117.375 21.240 117.565 ;
        RECT 21.530 117.355 21.700 117.565 ;
        RECT 22.450 117.355 22.620 117.545 ;
        RECT 23.185 117.375 23.355 117.565 ;
        RECT 30.455 117.375 30.625 117.565 ;
        RECT 31.190 117.375 31.360 117.565 ;
        RECT 32.590 117.545 32.740 117.565 ;
        RECT 35.810 117.545 35.960 117.565 ;
        RECT 39.030 117.545 39.180 117.565 ;
        RECT 32.165 117.405 32.285 117.515 ;
        RECT 32.570 117.355 32.740 117.545 ;
        RECT 34.225 117.355 34.395 117.545 ;
        RECT 35.385 117.405 35.505 117.515 ;
        RECT 35.790 117.375 35.960 117.545 ;
        RECT 38.550 117.410 38.710 117.520 ;
        RECT 39.010 117.375 39.180 117.545 ;
        RECT 43.150 117.545 43.300 117.565 ;
        RECT 43.150 117.375 43.320 117.545 ;
        RECT 47.015 117.375 47.185 117.565 ;
        RECT 47.290 117.355 47.460 117.545 ;
        RECT 47.805 117.405 47.925 117.515 ;
        RECT 51.615 117.375 51.785 117.565 ;
        RECT 52.350 117.375 52.520 117.565 ;
        RECT 53.730 117.375 53.900 117.565 ;
        RECT 55.110 117.375 55.280 117.565 ;
        RECT 57.410 117.355 57.580 117.545 ;
        RECT 57.870 117.355 58.040 117.545 ;
        RECT 59.895 117.375 60.065 117.565 ;
        RECT 61.365 117.375 61.535 117.565 ;
        RECT 65.230 117.375 65.400 117.565 ;
        RECT 67.530 117.375 67.700 117.565 ;
        RECT 68.450 117.355 68.620 117.545 ;
        RECT 68.965 117.405 69.085 117.515 ;
        RECT 69.370 117.355 69.540 117.545 ;
        RECT 70.750 117.355 70.920 117.545 ;
        RECT 72.130 117.355 72.300 117.545 ;
        RECT 74.245 117.355 74.415 117.545 ;
        RECT 78.110 117.515 78.280 117.565 ;
        RECT 80.410 117.545 80.560 117.565 ;
        RECT 78.110 117.405 78.285 117.515 ;
        RECT 78.110 117.375 78.280 117.405 ;
        RECT 80.410 117.375 80.580 117.545 ;
        RECT 81.790 117.375 81.960 117.565 ;
        RECT 85.655 117.375 85.825 117.565 ;
        RECT 87.310 117.410 87.470 117.520 ;
        RECT 87.770 117.355 87.940 117.545 ;
        RECT 89.150 117.355 89.320 117.545 ;
        RECT 96.970 117.375 97.140 117.565 ;
        RECT 98.810 117.355 98.980 117.545 ;
        RECT 99.785 117.405 99.905 117.515 ;
        RECT 100.835 117.375 101.005 117.565 ;
        RECT 101.110 117.355 101.280 117.545 ;
        RECT 104.975 117.375 105.145 117.565 ;
        RECT 105.710 117.375 105.880 117.565 ;
        RECT 107.090 117.375 107.260 117.565 ;
        RECT 110.770 117.355 110.940 117.565 ;
        RECT 112.150 117.355 112.320 117.565 ;
        RECT 18.170 116.545 19.540 117.355 ;
        RECT 20.480 116.445 21.830 117.355 ;
        RECT 21.860 116.485 22.290 117.270 ;
        RECT 22.310 116.675 31.590 117.355 ;
        RECT 23.670 116.455 24.590 116.675 ;
        RECT 29.255 116.555 31.590 116.675 ;
        RECT 30.670 116.445 31.590 116.555 ;
        RECT 32.440 116.445 33.790 117.355 ;
        RECT 33.810 116.675 37.710 117.355 ;
        RECT 38.320 116.675 47.600 117.355 ;
        RECT 33.810 116.445 34.740 116.675 ;
        RECT 38.320 116.555 40.655 116.675 ;
        RECT 38.320 116.445 39.240 116.555 ;
        RECT 45.320 116.455 46.240 116.675 ;
        RECT 47.620 116.485 48.050 117.270 ;
        RECT 48.440 116.675 57.720 117.355 ;
        RECT 57.730 116.675 67.010 117.355 ;
        RECT 48.440 116.555 50.775 116.675 ;
        RECT 48.440 116.445 49.360 116.555 ;
        RECT 55.440 116.455 56.360 116.675 ;
        RECT 59.090 116.455 60.010 116.675 ;
        RECT 64.675 116.555 67.010 116.675 ;
        RECT 67.390 116.575 68.760 117.355 ;
        RECT 69.230 116.575 70.600 117.355 ;
        RECT 66.090 116.445 67.010 116.555 ;
        RECT 70.620 116.445 71.970 117.355 ;
        RECT 72.000 116.445 73.350 117.355 ;
        RECT 73.380 116.485 73.810 117.270 ;
        RECT 73.830 116.675 77.730 117.355 ;
        RECT 78.800 116.675 88.080 117.355 ;
        RECT 73.830 116.445 74.760 116.675 ;
        RECT 78.800 116.555 81.135 116.675 ;
        RECT 78.800 116.445 79.720 116.555 ;
        RECT 85.800 116.455 86.720 116.675 ;
        RECT 88.090 116.575 89.460 117.355 ;
        RECT 89.840 116.675 99.120 117.355 ;
        RECT 89.840 116.555 92.175 116.675 ;
        RECT 89.840 116.445 90.760 116.555 ;
        RECT 96.840 116.455 97.760 116.675 ;
        RECT 99.140 116.485 99.570 117.270 ;
        RECT 100.050 116.575 101.420 117.355 ;
        RECT 101.800 116.675 111.080 117.355 ;
        RECT 101.800 116.555 104.135 116.675 ;
        RECT 101.800 116.445 102.720 116.555 ;
        RECT 108.800 116.455 109.720 116.675 ;
        RECT 111.090 116.545 112.460 117.355 ;
      LAYER nwell ;
        RECT 17.975 113.325 112.655 116.155 ;
      LAYER pwell ;
        RECT 18.170 112.125 19.540 112.935 ;
        RECT 19.550 112.125 20.920 112.905 ;
        RECT 20.940 112.125 22.290 113.035 ;
        RECT 22.680 112.925 23.600 113.035 ;
        RECT 22.680 112.805 25.015 112.925 ;
        RECT 29.680 112.805 30.600 113.025 ;
        RECT 22.680 112.125 31.960 112.805 ;
        RECT 31.970 112.125 33.340 112.905 ;
        RECT 33.350 112.125 34.720 112.905 ;
        RECT 34.740 112.210 35.170 112.995 ;
        RECT 36.550 112.805 37.470 113.025 ;
        RECT 43.550 112.925 44.470 113.035 ;
        RECT 42.135 112.805 44.470 112.925 ;
        RECT 35.190 112.125 44.470 112.805 ;
        RECT 45.770 112.125 47.140 112.905 ;
        RECT 47.160 112.125 48.510 113.035 ;
        RECT 48.900 112.925 49.820 113.035 ;
        RECT 48.900 112.805 51.235 112.925 ;
        RECT 55.900 112.805 56.820 113.025 ;
        RECT 48.900 112.125 58.180 112.805 ;
        RECT 58.650 112.125 60.480 112.935 ;
        RECT 60.500 112.210 60.930 112.995 ;
        RECT 61.420 112.125 62.770 113.035 ;
        RECT 63.250 112.125 68.760 112.935 ;
        RECT 68.780 112.125 70.130 113.035 ;
        RECT 71.510 112.805 72.430 113.025 ;
        RECT 78.510 112.925 79.430 113.035 ;
        RECT 77.095 112.805 79.430 112.925 ;
        RECT 70.150 112.125 79.430 112.805 ;
        RECT 79.810 112.125 81.180 112.905 ;
        RECT 81.200 112.125 82.550 113.035 ;
        RECT 82.580 112.125 83.930 113.035 ;
        RECT 84.880 112.125 86.230 113.035 ;
        RECT 86.260 112.210 86.690 112.995 ;
        RECT 87.080 112.925 88.000 113.035 ;
        RECT 87.080 112.805 89.415 112.925 ;
        RECT 94.080 112.805 95.000 113.025 ;
        RECT 87.080 112.125 96.360 112.805 ;
        RECT 96.370 112.125 97.740 112.905 ;
        RECT 98.670 112.125 104.180 112.935 ;
        RECT 104.200 112.125 105.550 113.035 ;
        RECT 106.030 112.125 107.400 112.905 ;
        RECT 107.410 112.125 111.080 112.935 ;
        RECT 111.090 112.125 112.460 112.935 ;
        RECT 18.310 111.915 18.480 112.125 ;
        RECT 19.690 111.935 19.860 112.125 ;
        RECT 20.150 111.960 20.310 112.070 ;
        RECT 20.610 111.915 20.780 112.105 ;
        RECT 21.990 111.935 22.160 112.125 ;
        RECT 22.910 111.960 23.070 112.070 ;
        RECT 23.645 111.915 23.815 112.105 ;
        RECT 27.510 111.915 27.680 112.105 ;
        RECT 31.650 111.935 31.820 112.125 ;
        RECT 33.030 111.935 33.200 112.125 ;
        RECT 33.490 111.935 33.660 112.125 ;
        RECT 35.330 111.935 35.500 112.125 ;
        RECT 39.010 111.915 39.180 112.105 ;
        RECT 41.770 111.915 41.940 112.105 ;
        RECT 45.450 111.970 45.610 112.080 ;
        RECT 46.830 111.935 47.000 112.125 ;
        RECT 47.290 111.915 47.460 112.125 ;
        RECT 48.670 111.960 48.830 112.070 ;
        RECT 49.130 111.915 49.300 112.105 ;
        RECT 50.510 111.915 50.680 112.105 ;
        RECT 51.890 111.915 52.060 112.105 ;
        RECT 55.565 111.915 55.735 112.105 ;
        RECT 57.870 111.935 58.040 112.125 ;
        RECT 58.385 111.965 58.505 112.075 ;
        RECT 60.170 111.935 60.340 112.125 ;
        RECT 61.145 111.965 61.265 112.075 ;
        RECT 61.550 111.935 61.720 112.125 ;
        RECT 62.985 111.965 63.105 112.075 ;
        RECT 66.150 111.915 66.320 112.105 ;
        RECT 66.665 111.965 66.785 112.075 ;
        RECT 68.450 111.935 68.620 112.125 ;
        RECT 69.830 111.935 70.000 112.125 ;
        RECT 70.290 111.915 70.460 112.125 ;
        RECT 73.045 111.915 73.215 112.105 ;
        RECT 73.970 111.915 74.140 112.105 ;
        RECT 75.405 111.965 75.525 112.075 ;
        RECT 75.810 111.915 75.980 112.105 ;
        RECT 77.190 111.915 77.360 112.105 ;
        RECT 79.030 111.960 79.190 112.070 ;
        RECT 80.870 111.935 81.040 112.125 ;
        RECT 82.250 111.935 82.420 112.125 ;
        RECT 82.710 111.915 82.880 112.105 ;
        RECT 83.170 111.915 83.340 112.105 ;
        RECT 83.630 111.935 83.800 112.125 ;
        RECT 84.550 111.970 84.710 112.080 ;
        RECT 85.010 111.935 85.180 112.125 ;
        RECT 85.470 111.915 85.640 112.105 ;
        RECT 89.150 111.915 89.320 112.105 ;
        RECT 89.610 111.915 89.780 112.105 ;
        RECT 94.395 111.915 94.565 112.105 ;
        RECT 95.185 111.965 95.305 112.075 ;
        RECT 96.050 111.935 96.220 112.125 ;
        RECT 96.970 111.915 97.140 112.105 ;
        RECT 97.430 111.935 97.600 112.125 ;
        RECT 98.350 111.915 98.520 112.105 ;
        RECT 98.865 111.965 98.985 112.075 ;
        RECT 100.650 111.915 100.820 112.105 ;
        RECT 101.110 111.915 101.280 112.105 ;
        RECT 102.490 111.915 102.660 112.105 ;
        RECT 103.870 111.915 104.040 112.125 ;
        RECT 104.330 111.935 104.500 112.125 ;
        RECT 105.765 111.965 105.885 112.075 ;
        RECT 106.170 111.915 106.340 112.125 ;
        RECT 110.770 112.105 110.940 112.125 ;
        RECT 106.630 111.915 106.800 112.105 ;
        RECT 109.390 111.915 109.560 112.105 ;
        RECT 110.760 111.935 110.940 112.105 ;
        RECT 110.760 111.915 110.930 111.935 ;
        RECT 112.150 111.915 112.320 112.125 ;
        RECT 18.170 111.105 19.540 111.915 ;
        RECT 20.470 111.135 21.840 111.915 ;
        RECT 21.860 111.045 22.290 111.830 ;
        RECT 23.230 111.235 27.130 111.915 ;
        RECT 23.230 111.005 24.160 111.235 ;
        RECT 27.380 111.005 28.730 111.915 ;
        RECT 28.950 111.235 39.320 111.915 ;
        RECT 28.950 111.005 31.160 111.235 ;
        RECT 33.880 111.015 34.810 111.235 ;
        RECT 39.330 111.105 42.080 111.915 ;
        RECT 42.090 111.105 47.600 111.915 ;
        RECT 47.620 111.045 48.050 111.830 ;
        RECT 48.990 111.135 50.360 111.915 ;
        RECT 50.380 111.005 51.730 111.915 ;
        RECT 51.750 111.135 53.120 111.915 ;
        RECT 53.270 111.005 55.880 111.915 ;
        RECT 56.090 111.235 66.460 111.915 ;
        RECT 56.090 111.005 58.300 111.235 ;
        RECT 61.020 111.015 61.950 111.235 ;
        RECT 66.930 111.105 70.600 111.915 ;
        RECT 70.750 111.005 73.360 111.915 ;
        RECT 73.380 111.045 73.810 111.830 ;
        RECT 73.830 111.135 75.200 111.915 ;
        RECT 75.680 111.005 77.030 111.915 ;
        RECT 77.050 111.135 78.420 111.915 ;
        RECT 79.350 111.105 83.020 111.915 ;
        RECT 83.030 111.135 84.400 111.915 ;
        RECT 84.410 111.105 85.780 111.915 ;
        RECT 85.790 111.105 89.460 111.915 ;
        RECT 89.470 111.135 90.840 111.915 ;
        RECT 91.080 111.235 94.980 111.915 ;
        RECT 94.050 111.005 94.980 111.235 ;
        RECT 95.450 111.105 97.280 111.915 ;
        RECT 97.290 111.135 98.660 111.915 ;
        RECT 99.140 111.045 99.570 111.830 ;
        RECT 99.590 111.105 100.960 111.915 ;
        RECT 100.970 111.135 102.340 111.915 ;
        RECT 102.360 111.005 103.710 111.915 ;
        RECT 103.740 111.005 105.090 111.915 ;
        RECT 105.110 111.135 106.480 111.915 ;
        RECT 106.490 111.135 107.860 111.915 ;
        RECT 107.870 111.105 109.700 111.915 ;
        RECT 109.710 111.135 111.080 111.915 ;
        RECT 111.090 111.105 112.460 111.915 ;
      LAYER nwell ;
        RECT 17.975 107.885 112.655 110.715 ;
      LAYER pwell ;
        RECT 18.170 106.685 19.540 107.495 ;
        RECT 19.550 106.685 23.220 107.495 ;
        RECT 23.430 107.365 25.640 107.595 ;
        RECT 28.360 107.365 29.290 107.585 ;
        RECT 23.430 106.685 33.800 107.365 ;
        RECT 34.740 106.770 35.170 107.555 ;
        RECT 35.650 106.685 37.020 107.465 ;
        RECT 37.500 106.685 38.850 107.595 ;
        RECT 39.340 106.685 40.690 107.595 ;
        RECT 40.710 106.685 42.080 107.465 ;
        RECT 42.550 106.685 43.920 107.465 ;
        RECT 43.930 106.685 45.300 107.465 ;
        RECT 45.310 106.685 46.680 107.465 ;
        RECT 46.890 107.365 49.100 107.595 ;
        RECT 51.820 107.365 52.750 107.585 ;
        RECT 46.890 106.685 57.260 107.365 ;
        RECT 57.730 106.685 60.340 107.595 ;
        RECT 60.500 106.770 60.930 107.555 ;
        RECT 60.960 106.685 62.310 107.595 ;
        RECT 62.330 106.685 63.700 107.465 ;
        RECT 63.710 106.685 65.080 107.465 ;
        RECT 65.290 107.365 67.500 107.595 ;
        RECT 70.220 107.365 71.150 107.585 ;
        RECT 75.870 107.365 78.080 107.595 ;
        RECT 80.800 107.365 81.730 107.585 ;
        RECT 65.290 106.685 75.660 107.365 ;
        RECT 75.870 106.685 86.240 107.365 ;
        RECT 86.260 106.770 86.690 107.555 ;
        RECT 87.830 107.365 90.040 107.595 ;
        RECT 92.760 107.365 93.690 107.585 ;
        RECT 87.830 106.685 98.200 107.365 ;
        RECT 98.210 106.685 99.580 107.465 ;
        RECT 100.710 107.365 102.920 107.595 ;
        RECT 105.640 107.365 106.570 107.585 ;
        RECT 100.710 106.685 111.080 107.365 ;
        RECT 111.090 106.685 112.460 107.495 ;
        RECT 18.310 106.475 18.480 106.685 ;
        RECT 19.745 106.525 19.865 106.635 ;
        RECT 21.530 106.475 21.700 106.665 ;
        RECT 22.910 106.495 23.080 106.685 ;
        RECT 23.370 106.475 23.540 106.665 ;
        RECT 23.830 106.475 24.000 106.665 ;
        RECT 25.210 106.475 25.380 106.665 ;
        RECT 26.590 106.475 26.760 106.665 ;
        RECT 33.490 106.495 33.660 106.685 ;
        RECT 34.410 106.530 34.570 106.640 ;
        RECT 35.385 106.525 35.505 106.635 ;
        RECT 36.710 106.495 36.880 106.685 ;
        RECT 37.170 106.635 37.340 106.665 ;
        RECT 37.170 106.525 37.345 106.635 ;
        RECT 37.170 106.475 37.340 106.525 ;
        RECT 38.550 106.495 38.720 106.685 ;
        RECT 39.065 106.525 39.185 106.635 ;
        RECT 39.470 106.495 39.640 106.685 ;
        RECT 41.770 106.495 41.940 106.685 ;
        RECT 42.285 106.525 42.405 106.635 ;
        RECT 43.610 106.495 43.780 106.685 ;
        RECT 44.990 106.495 45.160 106.685 ;
        RECT 45.450 106.495 45.620 106.685 ;
        RECT 49.130 106.475 49.300 106.665 ;
        RECT 49.590 106.475 49.760 106.665 ;
        RECT 56.950 106.495 57.120 106.685 ;
        RECT 57.465 106.525 57.585 106.635 ;
        RECT 57.875 106.495 58.045 106.685 ;
        RECT 61.090 106.475 61.260 106.685 ;
        RECT 62.470 106.495 62.640 106.685 ;
        RECT 63.850 106.495 64.020 106.685 ;
        RECT 71.670 106.475 71.840 106.665 ;
        RECT 72.130 106.475 72.300 106.665 ;
        RECT 75.350 106.495 75.520 106.685 ;
        RECT 84.090 106.475 84.260 106.665 ;
        RECT 85.930 106.495 86.100 106.685 ;
        RECT 87.310 106.530 87.470 106.640 ;
        RECT 94.670 106.475 94.840 106.665 ;
        RECT 96.050 106.475 96.220 106.665 ;
        RECT 97.430 106.475 97.600 106.665 ;
        RECT 97.890 106.475 98.060 106.685 ;
        RECT 99.270 106.495 99.440 106.685 ;
        RECT 100.190 106.530 100.350 106.640 ;
        RECT 109.850 106.475 110.020 106.665 ;
        RECT 110.770 106.495 110.940 106.685 ;
        RECT 112.150 106.475 112.320 106.685 ;
        RECT 18.170 105.665 19.540 106.475 ;
        RECT 20.010 105.665 21.840 106.475 ;
        RECT 21.860 105.605 22.290 106.390 ;
        RECT 22.320 105.565 23.670 106.475 ;
        RECT 23.700 105.565 25.050 106.475 ;
        RECT 25.080 105.565 26.430 106.475 ;
        RECT 26.450 105.795 36.820 106.475 ;
        RECT 37.030 105.795 47.400 106.475 ;
        RECT 30.960 105.575 31.890 105.795 ;
        RECT 34.610 105.565 36.820 105.795 ;
        RECT 41.540 105.575 42.470 105.795 ;
        RECT 45.190 105.565 47.400 105.795 ;
        RECT 47.620 105.605 48.050 106.390 ;
        RECT 48.080 105.565 49.430 106.475 ;
        RECT 49.460 105.565 50.810 106.475 ;
        RECT 51.030 105.795 61.400 106.475 ;
        RECT 61.610 105.795 71.980 106.475 ;
        RECT 51.030 105.565 53.240 105.795 ;
        RECT 55.960 105.575 56.890 105.795 ;
        RECT 61.610 105.565 63.820 105.795 ;
        RECT 66.540 105.575 67.470 105.795 ;
        RECT 71.990 105.695 73.360 106.475 ;
        RECT 73.380 105.605 73.810 106.390 ;
        RECT 74.030 105.795 84.400 106.475 ;
        RECT 84.610 105.795 94.980 106.475 ;
        RECT 74.030 105.565 76.240 105.795 ;
        RECT 78.960 105.575 79.890 105.795 ;
        RECT 84.610 105.565 86.820 105.795 ;
        RECT 89.540 105.575 90.470 105.795 ;
        RECT 95.000 105.565 96.350 106.475 ;
        RECT 96.380 105.565 97.730 106.475 ;
        RECT 97.760 105.565 99.110 106.475 ;
        RECT 99.140 105.605 99.570 106.390 ;
        RECT 99.790 105.795 110.160 106.475 ;
        RECT 99.790 105.565 102.000 105.795 ;
        RECT 104.720 105.575 105.650 105.795 ;
        RECT 111.090 105.665 112.460 106.475 ;
      LAYER nwell ;
        RECT 17.975 102.445 112.655 105.275 ;
      LAYER pwell ;
        RECT 18.170 101.245 19.540 102.055 ;
        RECT 20.010 101.245 21.840 102.055 ;
        RECT 21.860 101.330 22.290 102.115 ;
        RECT 22.510 101.925 24.720 102.155 ;
        RECT 27.440 101.925 28.370 102.145 ;
        RECT 22.510 101.245 32.880 101.925 ;
        RECT 32.890 101.245 34.720 102.055 ;
        RECT 34.740 101.330 35.170 102.115 ;
        RECT 35.190 101.245 37.020 102.055 ;
        RECT 37.230 101.925 39.440 102.155 ;
        RECT 42.160 101.925 43.090 102.145 ;
        RECT 37.230 101.245 47.600 101.925 ;
        RECT 47.620 101.330 48.050 102.115 ;
        RECT 48.070 101.245 49.900 102.055 ;
        RECT 49.910 101.245 55.420 102.055 ;
        RECT 55.440 101.245 56.790 102.155 ;
        RECT 56.810 101.245 58.180 102.025 ;
        RECT 59.120 101.245 60.470 102.155 ;
        RECT 60.500 101.330 60.930 102.115 ;
        RECT 61.410 101.245 65.080 102.055 ;
        RECT 65.090 101.245 70.600 102.055 ;
        RECT 70.620 101.245 71.970 102.155 ;
        RECT 72.000 101.245 73.350 102.155 ;
        RECT 73.380 101.330 73.810 102.115 ;
        RECT 74.030 101.925 76.240 102.155 ;
        RECT 78.960 101.925 79.890 102.145 ;
        RECT 74.030 101.245 84.400 101.925 ;
        RECT 84.420 101.245 85.770 102.155 ;
        RECT 86.260 101.330 86.690 102.115 ;
        RECT 86.720 101.245 88.070 102.155 ;
        RECT 88.750 101.925 90.960 102.155 ;
        RECT 93.680 101.925 94.610 102.145 ;
        RECT 88.750 101.245 99.120 101.925 ;
        RECT 99.140 101.330 99.570 102.115 ;
        RECT 105.020 101.925 105.950 102.145 ;
        RECT 108.670 101.925 110.880 102.155 ;
        RECT 100.510 101.245 110.880 101.925 ;
        RECT 111.090 101.245 112.460 102.055 ;
        RECT 18.310 101.055 18.480 101.245 ;
        RECT 19.745 101.085 19.865 101.195 ;
        RECT 21.530 101.055 21.700 101.245 ;
        RECT 32.570 101.055 32.740 101.245 ;
        RECT 34.410 101.055 34.580 101.245 ;
        RECT 36.710 101.055 36.880 101.245 ;
        RECT 47.290 101.055 47.460 101.245 ;
        RECT 49.590 101.055 49.760 101.245 ;
        RECT 55.110 101.055 55.280 101.245 ;
        RECT 56.490 101.055 56.660 101.245 ;
        RECT 56.950 101.055 57.120 101.245 ;
        RECT 58.790 101.090 58.950 101.200 ;
        RECT 59.250 101.055 59.420 101.245 ;
        RECT 61.145 101.085 61.265 101.195 ;
        RECT 64.770 101.055 64.940 101.245 ;
        RECT 70.290 101.055 70.460 101.245 ;
        RECT 71.670 101.055 71.840 101.245 ;
        RECT 72.130 101.055 72.300 101.245 ;
        RECT 84.090 101.055 84.260 101.245 ;
        RECT 85.470 101.055 85.640 101.245 ;
        RECT 85.985 101.085 86.105 101.195 ;
        RECT 86.850 101.055 87.020 101.245 ;
        RECT 88.285 101.085 88.405 101.195 ;
        RECT 98.810 101.055 98.980 101.245 ;
        RECT 100.190 101.090 100.350 101.200 ;
        RECT 100.650 101.055 100.820 101.245 ;
        RECT 112.150 101.055 112.320 101.245 ;
      LAYER nwell ;
        RECT 20.485 54.580 29.875 66.420 ;
        RECT 31.685 54.590 41.075 66.430 ;
        RECT 42.905 54.560 52.295 66.400 ;
        RECT 54.155 54.540 63.545 66.380 ;
        RECT 65.375 54.530 74.765 66.370 ;
        RECT 76.615 54.520 86.005 66.360 ;
        RECT 87.865 54.530 97.255 66.370 ;
        RECT 99.145 54.520 108.535 66.360 ;
        RECT 110.415 54.520 119.805 66.360 ;
        RECT 121.665 54.520 131.055 66.360 ;
        RECT 132.415 54.490 139.375 66.330 ;
        RECT 20.655 49.020 23.115 53.210 ;
      LAYER pwell ;
        RECT 20.555 45.340 22.915 48.340 ;
      LAYER nwell ;
        RECT 24.735 45.940 29.125 53.130 ;
        RECT 31.855 49.030 34.315 53.220 ;
      LAYER pwell ;
        RECT 31.755 45.350 34.115 48.350 ;
      LAYER nwell ;
        RECT 35.935 45.950 40.325 53.140 ;
        RECT 43.075 49.000 45.535 53.190 ;
      LAYER pwell ;
        RECT 42.975 45.320 45.335 48.320 ;
      LAYER nwell ;
        RECT 47.155 45.920 51.545 53.110 ;
        RECT 54.325 48.980 56.785 53.170 ;
      LAYER pwell ;
        RECT 54.225 45.300 56.585 48.300 ;
      LAYER nwell ;
        RECT 58.405 45.900 62.795 53.090 ;
        RECT 65.545 48.970 68.005 53.160 ;
      LAYER pwell ;
        RECT 65.445 45.290 67.805 48.290 ;
      LAYER nwell ;
        RECT 69.625 45.890 74.015 53.080 ;
        RECT 76.785 48.960 79.245 53.150 ;
      LAYER pwell ;
        RECT 76.685 45.280 79.045 48.280 ;
      LAYER nwell ;
        RECT 80.865 45.880 85.255 53.070 ;
        RECT 88.035 48.970 90.495 53.160 ;
      LAYER pwell ;
        RECT 87.935 45.290 90.295 48.290 ;
      LAYER nwell ;
        RECT 92.115 45.890 96.505 53.080 ;
        RECT 99.315 48.960 101.775 53.150 ;
      LAYER pwell ;
        RECT 99.215 45.280 101.575 48.280 ;
      LAYER nwell ;
        RECT 103.395 45.880 107.785 53.070 ;
        RECT 110.585 48.960 113.045 53.150 ;
      LAYER pwell ;
        RECT 110.485 45.280 112.845 48.280 ;
      LAYER nwell ;
        RECT 114.665 45.880 119.055 53.070 ;
        RECT 121.835 48.960 124.295 53.150 ;
      LAYER pwell ;
        RECT 121.735 45.280 124.095 48.280 ;
      LAYER nwell ;
        RECT 125.915 45.880 130.305 53.070 ;
        RECT 19.615 32.280 24.005 39.470 ;
      LAYER pwell ;
        RECT 25.825 37.070 28.185 40.070 ;
      LAYER nwell ;
        RECT 25.625 32.200 28.085 36.390 ;
        RECT 30.895 32.280 35.285 39.470 ;
      LAYER pwell ;
        RECT 37.105 37.070 39.465 40.070 ;
      LAYER nwell ;
        RECT 36.905 32.200 39.365 36.390 ;
        RECT 42.185 32.260 46.575 39.450 ;
      LAYER pwell ;
        RECT 48.395 37.050 50.755 40.050 ;
      LAYER nwell ;
        RECT 48.195 32.180 50.655 36.370 ;
        RECT 53.405 32.260 57.795 39.450 ;
      LAYER pwell ;
        RECT 59.615 37.050 61.975 40.050 ;
      LAYER nwell ;
        RECT 59.415 32.180 61.875 36.370 ;
        RECT 64.605 32.260 68.995 39.450 ;
      LAYER pwell ;
        RECT 70.815 37.050 73.175 40.050 ;
      LAYER nwell ;
        RECT 70.615 32.180 73.075 36.370 ;
        RECT 75.895 32.250 80.285 39.440 ;
      LAYER pwell ;
        RECT 82.105 37.040 84.465 40.040 ;
      LAYER nwell ;
        RECT 81.905 32.170 84.365 36.360 ;
        RECT 87.135 32.270 91.525 39.460 ;
      LAYER pwell ;
        RECT 93.345 37.060 95.705 40.060 ;
      LAYER nwell ;
        RECT 93.145 32.190 95.605 36.380 ;
        RECT 98.345 32.290 102.735 39.480 ;
      LAYER pwell ;
        RECT 104.555 37.080 106.915 40.080 ;
      LAYER nwell ;
        RECT 104.355 32.210 106.815 36.400 ;
        RECT 109.545 32.330 113.935 39.520 ;
      LAYER pwell ;
        RECT 115.755 37.120 118.115 40.120 ;
      LAYER nwell ;
        RECT 115.555 32.250 118.015 36.440 ;
        RECT 120.755 32.350 125.145 39.540 ;
      LAYER pwell ;
        RECT 126.965 37.140 129.325 40.140 ;
      LAYER nwell ;
        RECT 126.765 32.270 129.225 36.460 ;
        RECT 18.865 18.990 28.255 30.830 ;
        RECT 30.145 18.990 39.535 30.830 ;
        RECT 41.435 18.970 50.825 30.810 ;
        RECT 52.655 18.970 62.045 30.810 ;
        RECT 63.855 18.970 73.245 30.810 ;
        RECT 75.145 18.960 84.535 30.800 ;
        RECT 86.385 18.980 95.775 30.820 ;
        RECT 97.595 19.000 106.985 30.840 ;
        RECT 108.795 19.040 118.185 30.880 ;
        RECT 120.005 19.060 129.395 30.900 ;
        RECT 131.725 19.030 138.685 30.870 ;
      LAYER li1 ;
        RECT 18.165 193.535 112.465 193.705 ;
        RECT 18.250 192.785 19.460 193.535 ;
        RECT 18.250 192.245 18.770 192.785 ;
        RECT 20.090 192.765 21.760 193.535 ;
        RECT 21.930 192.810 22.220 193.535 ;
        RECT 22.390 192.785 23.600 193.535 ;
        RECT 23.775 192.990 29.120 193.535 ;
        RECT 29.295 192.990 34.640 193.535 ;
        RECT 18.940 192.075 19.460 192.615 ;
        RECT 18.250 190.985 19.460 192.075 ;
        RECT 20.090 192.075 20.840 192.595 ;
        RECT 21.010 192.245 21.760 192.765 ;
        RECT 20.090 190.985 21.760 192.075 ;
        RECT 21.930 190.985 22.220 192.150 ;
        RECT 22.390 192.075 22.910 192.615 ;
        RECT 23.080 192.245 23.600 192.785 ;
        RECT 22.390 190.985 23.600 192.075 ;
        RECT 25.365 191.420 25.715 192.670 ;
        RECT 27.195 192.160 27.535 192.990 ;
        RECT 30.885 191.420 31.235 192.670 ;
        RECT 32.715 192.160 33.055 192.990 ;
        RECT 34.810 192.810 35.100 193.535 ;
        RECT 35.270 192.785 36.480 193.535 ;
        RECT 36.655 192.990 42.000 193.535 ;
        RECT 42.175 192.990 47.520 193.535 ;
        RECT 23.775 190.985 29.120 191.420 ;
        RECT 29.295 190.985 34.640 191.420 ;
        RECT 34.810 190.985 35.100 192.150 ;
        RECT 35.270 192.075 35.790 192.615 ;
        RECT 35.960 192.245 36.480 192.785 ;
        RECT 35.270 190.985 36.480 192.075 ;
        RECT 38.245 191.420 38.595 192.670 ;
        RECT 40.075 192.160 40.415 192.990 ;
        RECT 43.765 191.420 44.115 192.670 ;
        RECT 45.595 192.160 45.935 192.990 ;
        RECT 47.690 192.810 47.980 193.535 ;
        RECT 48.150 192.785 49.360 193.535 ;
        RECT 49.535 192.990 54.880 193.535 ;
        RECT 55.055 192.990 60.400 193.535 ;
        RECT 36.655 190.985 42.000 191.420 ;
        RECT 42.175 190.985 47.520 191.420 ;
        RECT 47.690 190.985 47.980 192.150 ;
        RECT 48.150 192.075 48.670 192.615 ;
        RECT 48.840 192.245 49.360 192.785 ;
        RECT 48.150 190.985 49.360 192.075 ;
        RECT 51.125 191.420 51.475 192.670 ;
        RECT 52.955 192.160 53.295 192.990 ;
        RECT 56.645 191.420 56.995 192.670 ;
        RECT 58.475 192.160 58.815 192.990 ;
        RECT 60.570 192.810 60.860 193.535 ;
        RECT 61.030 192.785 62.240 193.535 ;
        RECT 62.415 192.990 67.760 193.535 ;
        RECT 67.935 192.990 73.280 193.535 ;
        RECT 49.535 190.985 54.880 191.420 ;
        RECT 55.055 190.985 60.400 191.420 ;
        RECT 60.570 190.985 60.860 192.150 ;
        RECT 61.030 192.075 61.550 192.615 ;
        RECT 61.720 192.245 62.240 192.785 ;
        RECT 61.030 190.985 62.240 192.075 ;
        RECT 64.005 191.420 64.355 192.670 ;
        RECT 65.835 192.160 66.175 192.990 ;
        RECT 69.525 191.420 69.875 192.670 ;
        RECT 71.355 192.160 71.695 192.990 ;
        RECT 73.450 192.810 73.740 193.535 ;
        RECT 73.910 192.785 75.120 193.535 ;
        RECT 75.295 192.990 80.640 193.535 ;
        RECT 80.815 192.990 86.160 193.535 ;
        RECT 62.415 190.985 67.760 191.420 ;
        RECT 67.935 190.985 73.280 191.420 ;
        RECT 73.450 190.985 73.740 192.150 ;
        RECT 73.910 192.075 74.430 192.615 ;
        RECT 74.600 192.245 75.120 192.785 ;
        RECT 73.910 190.985 75.120 192.075 ;
        RECT 76.885 191.420 77.235 192.670 ;
        RECT 78.715 192.160 79.055 192.990 ;
        RECT 82.405 191.420 82.755 192.670 ;
        RECT 84.235 192.160 84.575 192.990 ;
        RECT 86.330 192.810 86.620 193.535 ;
        RECT 86.790 192.785 88.000 193.535 ;
        RECT 88.175 192.990 93.520 193.535 ;
        RECT 93.695 192.990 99.040 193.535 ;
        RECT 75.295 190.985 80.640 191.420 ;
        RECT 80.815 190.985 86.160 191.420 ;
        RECT 86.330 190.985 86.620 192.150 ;
        RECT 86.790 192.075 87.310 192.615 ;
        RECT 87.480 192.245 88.000 192.785 ;
        RECT 86.790 190.985 88.000 192.075 ;
        RECT 89.765 191.420 90.115 192.670 ;
        RECT 91.595 192.160 91.935 192.990 ;
        RECT 95.285 191.420 95.635 192.670 ;
        RECT 97.115 192.160 97.455 192.990 ;
        RECT 99.210 192.810 99.500 193.535 ;
        RECT 100.135 192.990 105.480 193.535 ;
        RECT 105.655 192.990 111.000 193.535 ;
        RECT 88.175 190.985 93.520 191.420 ;
        RECT 93.695 190.985 99.040 191.420 ;
        RECT 99.210 190.985 99.500 192.150 ;
        RECT 101.725 191.420 102.075 192.670 ;
        RECT 103.555 192.160 103.895 192.990 ;
        RECT 107.245 191.420 107.595 192.670 ;
        RECT 109.075 192.160 109.415 192.990 ;
        RECT 111.170 192.785 112.380 193.535 ;
        RECT 111.170 192.075 111.690 192.615 ;
        RECT 111.860 192.245 112.380 192.785 ;
        RECT 100.135 190.985 105.480 191.420 ;
        RECT 105.655 190.985 111.000 191.420 ;
        RECT 111.170 190.985 112.380 192.075 ;
        RECT 18.165 190.815 112.465 190.985 ;
        RECT 18.250 189.725 19.460 190.815 ;
        RECT 18.250 189.015 18.770 189.555 ;
        RECT 18.940 189.185 19.460 189.725 ;
        RECT 20.090 189.725 23.600 190.815 ;
        RECT 23.775 190.380 29.120 190.815 ;
        RECT 29.295 190.380 34.640 190.815 ;
        RECT 20.090 189.205 21.780 189.725 ;
        RECT 21.950 189.035 23.600 189.555 ;
        RECT 25.365 189.130 25.715 190.380 ;
        RECT 18.250 188.265 19.460 189.015 ;
        RECT 20.090 188.265 23.600 189.035 ;
        RECT 27.195 188.810 27.535 189.640 ;
        RECT 30.885 189.130 31.235 190.380 ;
        RECT 34.810 189.650 35.100 190.815 ;
        RECT 35.730 189.725 38.320 190.815 ;
        RECT 38.495 190.380 43.840 190.815 ;
        RECT 44.015 190.380 49.360 190.815 ;
        RECT 49.535 190.380 54.880 190.815 ;
        RECT 55.055 190.380 60.400 190.815 ;
        RECT 32.715 188.810 33.055 189.640 ;
        RECT 35.730 189.205 36.940 189.725 ;
        RECT 37.110 189.035 38.320 189.555 ;
        RECT 40.085 189.130 40.435 190.380 ;
        RECT 23.775 188.265 29.120 188.810 ;
        RECT 29.295 188.265 34.640 188.810 ;
        RECT 34.810 188.265 35.100 188.990 ;
        RECT 35.730 188.265 38.320 189.035 ;
        RECT 41.915 188.810 42.255 189.640 ;
        RECT 45.605 189.130 45.955 190.380 ;
        RECT 47.435 188.810 47.775 189.640 ;
        RECT 51.125 189.130 51.475 190.380 ;
        RECT 52.955 188.810 53.295 189.640 ;
        RECT 56.645 189.130 56.995 190.380 ;
        RECT 60.570 189.650 60.860 190.815 ;
        RECT 61.030 189.725 62.700 190.815 ;
        RECT 62.875 190.380 68.220 190.815 ;
        RECT 58.475 188.810 58.815 189.640 ;
        RECT 61.030 189.205 61.780 189.725 ;
        RECT 61.950 189.035 62.700 189.555 ;
        RECT 64.465 189.130 64.815 190.380 ;
        RECT 68.450 189.675 68.660 190.815 ;
        RECT 68.830 189.665 69.160 190.645 ;
        RECT 69.330 189.675 69.560 190.815 ;
        RECT 69.775 190.380 75.120 190.815 ;
        RECT 75.295 190.380 80.640 190.815 ;
        RECT 80.815 190.380 86.160 190.815 ;
        RECT 38.495 188.265 43.840 188.810 ;
        RECT 44.015 188.265 49.360 188.810 ;
        RECT 49.535 188.265 54.880 188.810 ;
        RECT 55.055 188.265 60.400 188.810 ;
        RECT 60.570 188.265 60.860 188.990 ;
        RECT 61.030 188.265 62.700 189.035 ;
        RECT 66.295 188.810 66.635 189.640 ;
        RECT 62.875 188.265 68.220 188.810 ;
        RECT 68.450 188.265 68.660 189.085 ;
        RECT 68.830 189.065 69.080 189.665 ;
        RECT 69.250 189.255 69.580 189.505 ;
        RECT 71.365 189.130 71.715 190.380 ;
        RECT 68.830 188.435 69.160 189.065 ;
        RECT 69.330 188.265 69.560 189.085 ;
        RECT 73.195 188.810 73.535 189.640 ;
        RECT 76.885 189.130 77.235 190.380 ;
        RECT 78.715 188.810 79.055 189.640 ;
        RECT 82.405 189.130 82.755 190.380 ;
        RECT 86.330 189.650 86.620 190.815 ;
        RECT 87.250 189.725 88.920 190.815 ;
        RECT 89.095 190.380 94.440 190.815 ;
        RECT 94.615 190.380 99.960 190.815 ;
        RECT 100.135 190.380 105.480 190.815 ;
        RECT 105.655 190.380 111.000 190.815 ;
        RECT 84.235 188.810 84.575 189.640 ;
        RECT 87.250 189.205 88.000 189.725 ;
        RECT 88.170 189.035 88.920 189.555 ;
        RECT 90.685 189.130 91.035 190.380 ;
        RECT 69.775 188.265 75.120 188.810 ;
        RECT 75.295 188.265 80.640 188.810 ;
        RECT 80.815 188.265 86.160 188.810 ;
        RECT 86.330 188.265 86.620 188.990 ;
        RECT 87.250 188.265 88.920 189.035 ;
        RECT 92.515 188.810 92.855 189.640 ;
        RECT 96.205 189.130 96.555 190.380 ;
        RECT 98.035 188.810 98.375 189.640 ;
        RECT 101.725 189.130 102.075 190.380 ;
        RECT 103.555 188.810 103.895 189.640 ;
        RECT 107.245 189.130 107.595 190.380 ;
        RECT 111.170 189.725 112.380 190.815 ;
        RECT 109.075 188.810 109.415 189.640 ;
        RECT 111.170 189.185 111.690 189.725 ;
        RECT 111.860 189.015 112.380 189.555 ;
        RECT 89.095 188.265 94.440 188.810 ;
        RECT 94.615 188.265 99.960 188.810 ;
        RECT 100.135 188.265 105.480 188.810 ;
        RECT 105.655 188.265 111.000 188.810 ;
        RECT 111.170 188.265 112.380 189.015 ;
        RECT 18.165 188.095 112.465 188.265 ;
        RECT 18.250 187.345 19.460 188.095 ;
        RECT 18.250 186.805 18.770 187.345 ;
        RECT 20.090 187.325 21.760 188.095 ;
        RECT 21.930 187.370 22.220 188.095 ;
        RECT 22.850 187.325 25.440 188.095 ;
        RECT 25.615 187.550 30.960 188.095 ;
        RECT 31.135 187.550 36.480 188.095 ;
        RECT 36.655 187.550 42.000 188.095 ;
        RECT 42.175 187.550 47.520 188.095 ;
        RECT 18.940 186.635 19.460 187.175 ;
        RECT 18.250 185.545 19.460 186.635 ;
        RECT 20.090 186.635 20.840 187.155 ;
        RECT 21.010 186.805 21.760 187.325 ;
        RECT 20.090 185.545 21.760 186.635 ;
        RECT 21.930 185.545 22.220 186.710 ;
        RECT 22.850 186.635 24.060 187.155 ;
        RECT 24.230 186.805 25.440 187.325 ;
        RECT 22.850 185.545 25.440 186.635 ;
        RECT 27.205 185.980 27.555 187.230 ;
        RECT 29.035 186.720 29.375 187.550 ;
        RECT 32.725 185.980 33.075 187.230 ;
        RECT 34.555 186.720 34.895 187.550 ;
        RECT 38.245 185.980 38.595 187.230 ;
        RECT 40.075 186.720 40.415 187.550 ;
        RECT 43.765 185.980 44.115 187.230 ;
        RECT 45.595 186.720 45.935 187.550 ;
        RECT 47.690 187.370 47.980 188.095 ;
        RECT 48.150 187.325 50.740 188.095 ;
        RECT 50.915 187.550 56.260 188.095 ;
        RECT 25.615 185.545 30.960 185.980 ;
        RECT 31.135 185.545 36.480 185.980 ;
        RECT 36.655 185.545 42.000 185.980 ;
        RECT 42.175 185.545 47.520 185.980 ;
        RECT 47.690 185.545 47.980 186.710 ;
        RECT 48.150 186.635 49.360 187.155 ;
        RECT 49.530 186.805 50.740 187.325 ;
        RECT 48.150 185.545 50.740 186.635 ;
        RECT 52.505 185.980 52.855 187.230 ;
        RECT 54.335 186.720 54.675 187.550 ;
        RECT 56.490 187.275 56.700 188.095 ;
        RECT 56.870 187.295 57.200 187.925 ;
        RECT 56.870 186.695 57.120 187.295 ;
        RECT 57.370 187.275 57.600 188.095 ;
        RECT 57.850 187.275 58.080 188.095 ;
        RECT 58.250 187.295 58.580 187.925 ;
        RECT 57.290 186.855 57.620 187.105 ;
        RECT 57.830 186.855 58.160 187.105 ;
        RECT 58.330 186.695 58.580 187.295 ;
        RECT 58.750 187.275 58.960 188.095 ;
        RECT 59.195 187.385 59.450 187.915 ;
        RECT 59.620 187.635 59.925 188.095 ;
        RECT 60.170 187.715 61.240 187.885 ;
        RECT 50.915 185.545 56.260 185.980 ;
        RECT 56.490 185.545 56.700 186.685 ;
        RECT 56.870 185.715 57.200 186.695 ;
        RECT 57.370 185.545 57.600 186.685 ;
        RECT 57.850 185.545 58.080 186.685 ;
        RECT 58.250 185.715 58.580 186.695 ;
        RECT 59.195 186.735 59.405 187.385 ;
        RECT 60.170 187.360 60.490 187.715 ;
        RECT 60.165 187.185 60.490 187.360 ;
        RECT 59.575 186.885 60.490 187.185 ;
        RECT 60.660 187.145 60.900 187.545 ;
        RECT 61.070 187.485 61.240 187.715 ;
        RECT 61.410 187.655 61.600 188.095 ;
        RECT 61.770 187.645 62.720 187.925 ;
        RECT 62.940 187.735 63.290 187.905 ;
        RECT 61.070 187.315 61.600 187.485 ;
        RECT 59.575 186.855 60.315 186.885 ;
        RECT 58.750 185.545 58.960 186.685 ;
        RECT 59.195 185.855 59.450 186.735 ;
        RECT 59.620 185.545 59.925 186.685 ;
        RECT 60.145 186.265 60.315 186.855 ;
        RECT 60.660 186.775 61.200 187.145 ;
        RECT 61.380 187.035 61.600 187.315 ;
        RECT 61.770 186.865 61.940 187.645 ;
        RECT 61.535 186.695 61.940 186.865 ;
        RECT 62.110 186.855 62.460 187.475 ;
        RECT 61.535 186.605 61.705 186.695 ;
        RECT 62.630 186.685 62.840 187.475 ;
        RECT 60.485 186.435 61.705 186.605 ;
        RECT 62.165 186.525 62.840 186.685 ;
        RECT 60.145 186.095 60.945 186.265 ;
        RECT 60.265 185.545 60.595 185.925 ;
        RECT 60.775 185.805 60.945 186.095 ;
        RECT 61.535 186.055 61.705 186.435 ;
        RECT 61.875 186.515 62.840 186.525 ;
        RECT 63.030 187.345 63.290 187.735 ;
        RECT 63.500 187.635 63.830 188.095 ;
        RECT 64.705 187.705 65.560 187.875 ;
        RECT 65.765 187.705 66.260 187.875 ;
        RECT 66.430 187.735 66.760 188.095 ;
        RECT 63.030 186.655 63.200 187.345 ;
        RECT 63.370 186.995 63.540 187.175 ;
        RECT 63.710 187.165 64.500 187.415 ;
        RECT 64.705 186.995 64.875 187.705 ;
        RECT 65.045 187.195 65.400 187.415 ;
        RECT 63.370 186.825 65.060 186.995 ;
        RECT 61.875 186.225 62.335 186.515 ;
        RECT 63.030 186.485 64.530 186.655 ;
        RECT 63.030 186.345 63.200 186.485 ;
        RECT 62.640 186.175 63.200 186.345 ;
        RECT 61.115 185.545 61.365 186.005 ;
        RECT 61.535 185.715 62.405 186.055 ;
        RECT 62.640 185.715 62.810 186.175 ;
        RECT 63.645 186.145 64.720 186.315 ;
        RECT 62.980 185.545 63.350 186.005 ;
        RECT 63.645 185.805 63.815 186.145 ;
        RECT 63.985 185.545 64.315 185.975 ;
        RECT 64.550 185.805 64.720 186.145 ;
        RECT 64.890 186.045 65.060 186.825 ;
        RECT 65.230 186.605 65.400 187.195 ;
        RECT 65.570 186.795 65.920 187.415 ;
        RECT 65.230 186.215 65.695 186.605 ;
        RECT 66.090 186.345 66.260 187.705 ;
        RECT 66.430 186.515 66.890 187.565 ;
        RECT 65.865 186.175 66.260 186.345 ;
        RECT 65.865 186.045 66.035 186.175 ;
        RECT 64.890 185.715 65.570 186.045 ;
        RECT 65.785 185.715 66.035 186.045 ;
        RECT 66.205 185.545 66.455 186.005 ;
        RECT 66.625 185.730 66.950 186.515 ;
        RECT 67.120 185.715 67.290 187.835 ;
        RECT 67.460 187.715 67.790 188.095 ;
        RECT 67.960 187.545 68.215 187.835 ;
        RECT 67.465 187.375 68.215 187.545 ;
        RECT 67.465 186.385 67.695 187.375 ;
        RECT 68.390 187.355 68.710 187.835 ;
        RECT 68.880 187.525 69.110 187.925 ;
        RECT 69.280 187.705 69.630 188.095 ;
        RECT 68.880 187.445 69.390 187.525 ;
        RECT 69.800 187.445 70.130 187.925 ;
        RECT 68.880 187.355 70.130 187.445 ;
        RECT 67.865 186.555 68.215 187.205 ;
        RECT 68.390 186.425 68.560 187.355 ;
        RECT 69.220 187.275 70.130 187.355 ;
        RECT 70.300 187.275 70.470 188.095 ;
        RECT 70.975 187.355 71.440 187.900 ;
        RECT 68.730 186.765 68.900 187.185 ;
        RECT 69.130 186.935 69.730 187.105 ;
        RECT 68.730 186.595 69.390 186.765 ;
        RECT 67.465 186.215 68.215 186.385 ;
        RECT 68.390 186.225 69.050 186.425 ;
        RECT 69.220 186.395 69.390 186.595 ;
        RECT 69.560 186.735 69.730 186.935 ;
        RECT 69.900 186.905 70.595 187.105 ;
        RECT 70.855 186.735 71.100 187.185 ;
        RECT 69.560 186.565 71.100 186.735 ;
        RECT 71.270 186.395 71.440 187.355 ;
        RECT 71.610 187.325 73.280 188.095 ;
        RECT 73.450 187.370 73.740 188.095 ;
        RECT 74.830 187.325 78.340 188.095 ;
        RECT 78.515 187.550 83.860 188.095 ;
        RECT 84.035 187.550 89.380 188.095 ;
        RECT 89.555 187.550 94.900 188.095 ;
        RECT 69.220 186.225 71.440 186.395 ;
        RECT 71.610 186.635 72.360 187.155 ;
        RECT 72.530 186.805 73.280 187.325 ;
        RECT 67.460 185.545 67.790 186.045 ;
        RECT 67.960 185.715 68.215 186.215 ;
        RECT 68.880 186.055 69.050 186.225 ;
        RECT 68.410 185.545 68.710 186.055 ;
        RECT 68.880 185.885 69.260 186.055 ;
        RECT 69.840 185.545 70.470 186.055 ;
        RECT 70.640 185.715 70.970 186.225 ;
        RECT 71.140 185.545 71.440 186.055 ;
        RECT 71.610 185.545 73.280 186.635 ;
        RECT 73.450 185.545 73.740 186.710 ;
        RECT 74.830 186.635 76.520 187.155 ;
        RECT 76.690 186.805 78.340 187.325 ;
        RECT 74.830 185.545 78.340 186.635 ;
        RECT 80.105 185.980 80.455 187.230 ;
        RECT 81.935 186.720 82.275 187.550 ;
        RECT 85.625 185.980 85.975 187.230 ;
        RECT 87.455 186.720 87.795 187.550 ;
        RECT 91.145 185.980 91.495 187.230 ;
        RECT 92.975 186.720 93.315 187.550 ;
        RECT 95.110 187.275 95.340 188.095 ;
        RECT 95.510 187.295 95.840 187.925 ;
        RECT 95.090 186.855 95.420 187.105 ;
        RECT 95.590 186.695 95.840 187.295 ;
        RECT 96.010 187.275 96.220 188.095 ;
        RECT 96.450 187.325 99.040 188.095 ;
        RECT 99.210 187.370 99.500 188.095 ;
        RECT 100.135 187.550 105.480 188.095 ;
        RECT 105.655 187.550 111.000 188.095 ;
        RECT 78.515 185.545 83.860 185.980 ;
        RECT 84.035 185.545 89.380 185.980 ;
        RECT 89.555 185.545 94.900 185.980 ;
        RECT 95.110 185.545 95.340 186.685 ;
        RECT 95.510 185.715 95.840 186.695 ;
        RECT 96.010 185.545 96.220 186.685 ;
        RECT 96.450 186.635 97.660 187.155 ;
        RECT 97.830 186.805 99.040 187.325 ;
        RECT 96.450 185.545 99.040 186.635 ;
        RECT 99.210 185.545 99.500 186.710 ;
        RECT 101.725 185.980 102.075 187.230 ;
        RECT 103.555 186.720 103.895 187.550 ;
        RECT 107.245 185.980 107.595 187.230 ;
        RECT 109.075 186.720 109.415 187.550 ;
        RECT 111.170 187.345 112.380 188.095 ;
        RECT 111.170 186.635 111.690 187.175 ;
        RECT 111.860 186.805 112.380 187.345 ;
        RECT 100.135 185.545 105.480 185.980 ;
        RECT 105.655 185.545 111.000 185.980 ;
        RECT 111.170 185.545 112.380 186.635 ;
        RECT 18.165 185.375 112.465 185.545 ;
        RECT 18.250 184.285 19.460 185.375 ;
        RECT 18.250 183.575 18.770 184.115 ;
        RECT 18.940 183.745 19.460 184.285 ;
        RECT 20.090 184.285 23.600 185.375 ;
        RECT 23.775 184.940 29.120 185.375 ;
        RECT 29.295 184.940 34.640 185.375 ;
        RECT 20.090 183.765 21.780 184.285 ;
        RECT 21.950 183.595 23.600 184.115 ;
        RECT 25.365 183.690 25.715 184.940 ;
        RECT 18.250 182.825 19.460 183.575 ;
        RECT 20.090 182.825 23.600 183.595 ;
        RECT 27.195 183.370 27.535 184.200 ;
        RECT 30.885 183.690 31.235 184.940 ;
        RECT 34.810 184.210 35.100 185.375 ;
        RECT 35.270 184.285 36.480 185.375 ;
        RECT 36.650 184.285 40.160 185.375 ;
        RECT 40.335 184.940 45.680 185.375 ;
        RECT 45.855 184.940 51.200 185.375 ;
        RECT 32.715 183.370 33.055 184.200 ;
        RECT 35.270 183.745 35.790 184.285 ;
        RECT 35.960 183.575 36.480 184.115 ;
        RECT 36.650 183.765 38.340 184.285 ;
        RECT 38.510 183.595 40.160 184.115 ;
        RECT 41.925 183.690 42.275 184.940 ;
        RECT 23.775 182.825 29.120 183.370 ;
        RECT 29.295 182.825 34.640 183.370 ;
        RECT 34.810 182.825 35.100 183.550 ;
        RECT 35.270 182.825 36.480 183.575 ;
        RECT 36.650 182.825 40.160 183.595 ;
        RECT 43.755 183.370 44.095 184.200 ;
        RECT 47.445 183.690 47.795 184.940 ;
        RECT 51.375 184.705 51.630 185.205 ;
        RECT 51.800 184.875 52.130 185.375 ;
        RECT 51.375 184.535 52.125 184.705 ;
        RECT 49.275 183.370 49.615 184.200 ;
        RECT 51.375 183.715 51.725 184.365 ;
        RECT 51.895 183.545 52.125 184.535 ;
        RECT 51.375 183.375 52.125 183.545 ;
        RECT 40.335 182.825 45.680 183.370 ;
        RECT 45.855 182.825 51.200 183.370 ;
        RECT 51.375 183.085 51.630 183.375 ;
        RECT 51.800 182.825 52.130 183.205 ;
        RECT 52.300 183.085 52.470 185.205 ;
        RECT 52.640 184.405 52.965 185.190 ;
        RECT 53.135 184.915 53.385 185.375 ;
        RECT 53.555 184.875 53.805 185.205 ;
        RECT 54.020 184.875 54.700 185.205 ;
        RECT 53.555 184.745 53.725 184.875 ;
        RECT 53.330 184.575 53.725 184.745 ;
        RECT 52.700 183.355 53.160 184.405 ;
        RECT 53.330 183.215 53.500 184.575 ;
        RECT 53.895 184.315 54.360 184.705 ;
        RECT 53.670 183.505 54.020 184.125 ;
        RECT 54.190 183.725 54.360 184.315 ;
        RECT 54.530 184.095 54.700 184.875 ;
        RECT 54.870 184.775 55.040 185.115 ;
        RECT 55.275 184.945 55.605 185.375 ;
        RECT 55.775 184.775 55.945 185.115 ;
        RECT 56.240 184.915 56.610 185.375 ;
        RECT 54.870 184.605 55.945 184.775 ;
        RECT 56.780 184.745 56.950 185.205 ;
        RECT 57.185 184.865 58.055 185.205 ;
        RECT 58.225 184.915 58.475 185.375 ;
        RECT 56.390 184.575 56.950 184.745 ;
        RECT 56.390 184.435 56.560 184.575 ;
        RECT 55.060 184.265 56.560 184.435 ;
        RECT 57.255 184.405 57.715 184.695 ;
        RECT 54.530 183.925 56.220 184.095 ;
        RECT 54.190 183.505 54.545 183.725 ;
        RECT 54.715 183.215 54.885 183.925 ;
        RECT 55.090 183.505 55.880 183.755 ;
        RECT 56.050 183.745 56.220 183.925 ;
        RECT 56.390 183.575 56.560 184.265 ;
        RECT 52.830 182.825 53.160 183.185 ;
        RECT 53.330 183.045 53.825 183.215 ;
        RECT 54.030 183.045 54.885 183.215 ;
        RECT 55.760 182.825 56.090 183.285 ;
        RECT 56.300 183.185 56.560 183.575 ;
        RECT 56.750 184.395 57.715 184.405 ;
        RECT 57.885 184.485 58.055 184.865 ;
        RECT 58.645 184.825 58.815 185.115 ;
        RECT 58.995 184.995 59.325 185.375 ;
        RECT 58.645 184.655 59.445 184.825 ;
        RECT 56.750 184.235 57.425 184.395 ;
        RECT 57.885 184.315 59.105 184.485 ;
        RECT 56.750 183.445 56.960 184.235 ;
        RECT 57.885 184.225 58.055 184.315 ;
        RECT 57.130 183.445 57.480 184.065 ;
        RECT 57.650 184.055 58.055 184.225 ;
        RECT 57.650 183.275 57.820 184.055 ;
        RECT 57.990 183.605 58.210 183.885 ;
        RECT 58.390 183.775 58.930 184.145 ;
        RECT 59.275 184.065 59.445 184.655 ;
        RECT 59.665 184.235 59.970 185.375 ;
        RECT 60.140 184.185 60.395 185.065 ;
        RECT 60.570 184.210 60.860 185.375 ;
        RECT 61.120 184.445 61.290 185.205 ;
        RECT 61.505 184.615 61.835 185.375 ;
        RECT 61.120 184.275 61.835 184.445 ;
        RECT 62.005 184.300 62.260 185.205 ;
        RECT 59.275 184.035 60.015 184.065 ;
        RECT 57.990 183.435 58.520 183.605 ;
        RECT 56.300 183.015 56.650 183.185 ;
        RECT 56.870 182.995 57.820 183.275 ;
        RECT 57.990 182.825 58.180 183.265 ;
        RECT 58.350 183.205 58.520 183.435 ;
        RECT 58.690 183.375 58.930 183.775 ;
        RECT 59.100 183.735 60.015 184.035 ;
        RECT 59.100 183.560 59.425 183.735 ;
        RECT 59.100 183.205 59.420 183.560 ;
        RECT 60.185 183.535 60.395 184.185 ;
        RECT 61.030 183.725 61.385 184.095 ;
        RECT 61.665 184.065 61.835 184.275 ;
        RECT 61.665 183.735 61.920 184.065 ;
        RECT 58.350 183.035 59.420 183.205 ;
        RECT 59.665 182.825 59.970 183.285 ;
        RECT 60.140 183.005 60.395 183.535 ;
        RECT 60.570 182.825 60.860 183.550 ;
        RECT 61.665 183.545 61.835 183.735 ;
        RECT 62.090 183.570 62.260 184.300 ;
        RECT 62.435 184.225 62.695 185.375 ;
        RECT 63.790 184.300 64.060 185.205 ;
        RECT 64.230 184.615 64.560 185.375 ;
        RECT 64.740 184.445 64.910 185.205 ;
        RECT 61.120 183.375 61.835 183.545 ;
        RECT 61.120 182.995 61.290 183.375 ;
        RECT 61.505 182.825 61.835 183.205 ;
        RECT 62.005 182.995 62.260 183.570 ;
        RECT 62.435 182.825 62.695 183.665 ;
        RECT 63.790 183.500 63.960 184.300 ;
        RECT 64.245 184.275 64.910 184.445 ;
        RECT 64.245 184.130 64.415 184.275 ;
        RECT 64.130 183.800 64.415 184.130 ;
        RECT 65.175 184.185 65.430 185.065 ;
        RECT 65.600 184.235 65.905 185.375 ;
        RECT 66.245 184.995 66.575 185.375 ;
        RECT 66.755 184.825 66.925 185.115 ;
        RECT 67.095 184.915 67.345 185.375 ;
        RECT 66.125 184.655 66.925 184.825 ;
        RECT 67.515 184.865 68.385 185.205 ;
        RECT 64.245 183.545 64.415 183.800 ;
        RECT 64.650 183.725 64.980 184.095 ;
        RECT 63.790 182.995 64.050 183.500 ;
        RECT 64.245 183.375 64.910 183.545 ;
        RECT 64.230 182.825 64.560 183.205 ;
        RECT 64.740 182.995 64.910 183.375 ;
        RECT 65.175 183.535 65.385 184.185 ;
        RECT 66.125 184.065 66.295 184.655 ;
        RECT 67.515 184.485 67.685 184.865 ;
        RECT 68.620 184.745 68.790 185.205 ;
        RECT 68.960 184.915 69.330 185.375 ;
        RECT 69.625 184.775 69.795 185.115 ;
        RECT 69.965 184.945 70.295 185.375 ;
        RECT 70.530 184.775 70.700 185.115 ;
        RECT 66.465 184.315 67.685 184.485 ;
        RECT 67.855 184.405 68.315 184.695 ;
        RECT 68.620 184.575 69.180 184.745 ;
        RECT 69.625 184.605 70.700 184.775 ;
        RECT 70.870 184.875 71.550 185.205 ;
        RECT 71.765 184.875 72.015 185.205 ;
        RECT 72.185 184.915 72.435 185.375 ;
        RECT 69.010 184.435 69.180 184.575 ;
        RECT 67.855 184.395 68.820 184.405 ;
        RECT 67.515 184.225 67.685 184.315 ;
        RECT 68.145 184.235 68.820 184.395 ;
        RECT 65.555 184.035 66.295 184.065 ;
        RECT 65.555 183.735 66.470 184.035 ;
        RECT 66.145 183.560 66.470 183.735 ;
        RECT 65.175 183.005 65.430 183.535 ;
        RECT 65.600 182.825 65.905 183.285 ;
        RECT 66.150 183.205 66.470 183.560 ;
        RECT 66.640 183.775 67.180 184.145 ;
        RECT 67.515 184.055 67.920 184.225 ;
        RECT 66.640 183.375 66.880 183.775 ;
        RECT 67.360 183.605 67.580 183.885 ;
        RECT 67.050 183.435 67.580 183.605 ;
        RECT 67.050 183.205 67.220 183.435 ;
        RECT 67.750 183.275 67.920 184.055 ;
        RECT 68.090 183.445 68.440 184.065 ;
        RECT 68.610 183.445 68.820 184.235 ;
        RECT 69.010 184.265 70.510 184.435 ;
        RECT 69.010 183.575 69.180 184.265 ;
        RECT 70.870 184.095 71.040 184.875 ;
        RECT 71.845 184.745 72.015 184.875 ;
        RECT 69.350 183.925 71.040 184.095 ;
        RECT 71.210 184.315 71.675 184.705 ;
        RECT 71.845 184.575 72.240 184.745 ;
        RECT 69.350 183.745 69.520 183.925 ;
        RECT 66.150 183.035 67.220 183.205 ;
        RECT 67.390 182.825 67.580 183.265 ;
        RECT 67.750 182.995 68.700 183.275 ;
        RECT 69.010 183.185 69.270 183.575 ;
        RECT 69.690 183.505 70.480 183.755 ;
        RECT 68.920 183.015 69.270 183.185 ;
        RECT 69.480 182.825 69.810 183.285 ;
        RECT 70.685 183.215 70.855 183.925 ;
        RECT 71.210 183.725 71.380 184.315 ;
        RECT 71.025 183.505 71.380 183.725 ;
        RECT 71.550 183.505 71.900 184.125 ;
        RECT 72.070 183.215 72.240 184.575 ;
        RECT 72.605 184.405 72.930 185.190 ;
        RECT 72.410 183.355 72.870 184.405 ;
        RECT 70.685 183.045 71.540 183.215 ;
        RECT 71.745 183.045 72.240 183.215 ;
        RECT 72.410 182.825 72.740 183.185 ;
        RECT 73.100 183.085 73.270 185.205 ;
        RECT 73.440 184.875 73.770 185.375 ;
        RECT 73.940 184.705 74.195 185.205 ;
        RECT 73.445 184.535 74.195 184.705 ;
        RECT 73.445 183.545 73.675 184.535 ;
        RECT 73.845 183.715 74.195 184.365 ;
        RECT 74.410 184.235 74.640 185.375 ;
        RECT 74.810 184.225 75.140 185.205 ;
        RECT 75.310 184.235 75.520 185.375 ;
        RECT 75.750 184.285 78.340 185.375 ;
        RECT 74.390 183.815 74.720 184.065 ;
        RECT 73.445 183.375 74.195 183.545 ;
        RECT 73.440 182.825 73.770 183.205 ;
        RECT 73.940 183.085 74.195 183.375 ;
        RECT 74.410 182.825 74.640 183.645 ;
        RECT 74.890 183.625 75.140 184.225 ;
        RECT 75.750 183.765 76.960 184.285 ;
        RECT 78.550 184.235 78.780 185.375 ;
        RECT 78.950 184.225 79.280 185.205 ;
        RECT 79.450 184.235 79.660 185.375 ;
        RECT 79.890 184.615 80.405 185.025 ;
        RECT 80.640 184.615 80.810 185.375 ;
        RECT 80.980 185.035 83.010 185.205 ;
        RECT 74.810 182.995 75.140 183.625 ;
        RECT 75.310 182.825 75.520 183.645 ;
        RECT 77.130 183.595 78.340 184.115 ;
        RECT 78.530 183.815 78.860 184.065 ;
        RECT 75.750 182.825 78.340 183.595 ;
        RECT 78.550 182.825 78.780 183.645 ;
        RECT 79.030 183.625 79.280 184.225 ;
        RECT 79.890 183.805 80.230 184.615 ;
        RECT 80.980 184.370 81.150 185.035 ;
        RECT 81.545 184.695 82.670 184.865 ;
        RECT 80.400 184.180 81.150 184.370 ;
        RECT 81.320 184.355 82.330 184.525 ;
        RECT 78.950 182.995 79.280 183.625 ;
        RECT 79.450 182.825 79.660 183.645 ;
        RECT 79.890 183.635 81.120 183.805 ;
        RECT 80.165 183.030 80.410 183.635 ;
        RECT 80.630 182.825 81.140 183.360 ;
        RECT 81.320 182.995 81.510 184.355 ;
        RECT 81.680 183.335 81.955 184.155 ;
        RECT 82.160 183.555 82.330 184.355 ;
        RECT 82.500 183.565 82.670 184.695 ;
        RECT 82.840 184.065 83.010 185.035 ;
        RECT 83.180 184.235 83.350 185.375 ;
        RECT 83.520 184.235 83.855 185.205 ;
        RECT 84.120 184.445 84.290 185.205 ;
        RECT 84.470 184.615 84.800 185.375 ;
        RECT 84.120 184.275 84.785 184.445 ;
        RECT 84.970 184.300 85.240 185.205 ;
        RECT 82.840 183.735 83.035 184.065 ;
        RECT 83.260 183.735 83.515 184.065 ;
        RECT 83.260 183.565 83.430 183.735 ;
        RECT 83.685 183.565 83.855 184.235 ;
        RECT 84.615 184.130 84.785 184.275 ;
        RECT 84.050 183.725 84.380 184.095 ;
        RECT 84.615 183.800 84.900 184.130 ;
        RECT 82.500 183.395 83.430 183.565 ;
        RECT 82.500 183.360 82.675 183.395 ;
        RECT 81.680 183.165 81.960 183.335 ;
        RECT 81.680 182.995 81.955 183.165 ;
        RECT 82.145 182.995 82.675 183.360 ;
        RECT 83.100 182.825 83.430 183.225 ;
        RECT 83.600 182.995 83.855 183.565 ;
        RECT 84.615 183.545 84.785 183.800 ;
        RECT 84.120 183.375 84.785 183.545 ;
        RECT 85.070 183.500 85.240 184.300 ;
        RECT 86.330 184.210 86.620 185.375 ;
        RECT 86.830 184.235 87.060 185.375 ;
        RECT 87.230 184.225 87.560 185.205 ;
        RECT 87.730 184.235 87.940 185.375 ;
        RECT 88.175 184.705 88.430 185.205 ;
        RECT 88.600 184.875 88.930 185.375 ;
        RECT 88.175 184.535 88.925 184.705 ;
        RECT 86.810 183.815 87.140 184.065 ;
        RECT 84.120 182.995 84.290 183.375 ;
        RECT 84.470 182.825 84.800 183.205 ;
        RECT 84.980 182.995 85.240 183.500 ;
        RECT 86.330 182.825 86.620 183.550 ;
        RECT 86.830 182.825 87.060 183.645 ;
        RECT 87.310 183.625 87.560 184.225 ;
        RECT 88.175 183.715 88.525 184.365 ;
        RECT 87.230 182.995 87.560 183.625 ;
        RECT 87.730 182.825 87.940 183.645 ;
        RECT 88.695 183.545 88.925 184.535 ;
        RECT 88.175 183.375 88.925 183.545 ;
        RECT 88.175 183.085 88.430 183.375 ;
        RECT 88.600 182.825 88.930 183.205 ;
        RECT 89.100 183.085 89.270 185.205 ;
        RECT 89.440 184.405 89.765 185.190 ;
        RECT 89.935 184.915 90.185 185.375 ;
        RECT 90.355 184.875 90.605 185.205 ;
        RECT 90.820 184.875 91.500 185.205 ;
        RECT 90.355 184.745 90.525 184.875 ;
        RECT 90.130 184.575 90.525 184.745 ;
        RECT 89.500 183.355 89.960 184.405 ;
        RECT 90.130 183.215 90.300 184.575 ;
        RECT 90.695 184.315 91.160 184.705 ;
        RECT 90.470 183.505 90.820 184.125 ;
        RECT 90.990 183.725 91.160 184.315 ;
        RECT 91.330 184.095 91.500 184.875 ;
        RECT 91.670 184.775 91.840 185.115 ;
        RECT 92.075 184.945 92.405 185.375 ;
        RECT 92.575 184.775 92.745 185.115 ;
        RECT 93.040 184.915 93.410 185.375 ;
        RECT 91.670 184.605 92.745 184.775 ;
        RECT 93.580 184.745 93.750 185.205 ;
        RECT 93.985 184.865 94.855 185.205 ;
        RECT 95.025 184.915 95.275 185.375 ;
        RECT 93.190 184.575 93.750 184.745 ;
        RECT 93.190 184.435 93.360 184.575 ;
        RECT 91.860 184.265 93.360 184.435 ;
        RECT 94.055 184.405 94.515 184.695 ;
        RECT 91.330 183.925 93.020 184.095 ;
        RECT 90.990 183.505 91.345 183.725 ;
        RECT 91.515 183.215 91.685 183.925 ;
        RECT 91.890 183.505 92.680 183.755 ;
        RECT 92.850 183.745 93.020 183.925 ;
        RECT 93.190 183.575 93.360 184.265 ;
        RECT 89.630 182.825 89.960 183.185 ;
        RECT 90.130 183.045 90.625 183.215 ;
        RECT 90.830 183.045 91.685 183.215 ;
        RECT 92.560 182.825 92.890 183.285 ;
        RECT 93.100 183.185 93.360 183.575 ;
        RECT 93.550 184.395 94.515 184.405 ;
        RECT 94.685 184.485 94.855 184.865 ;
        RECT 95.445 184.825 95.615 185.115 ;
        RECT 95.795 184.995 96.125 185.375 ;
        RECT 95.445 184.655 96.245 184.825 ;
        RECT 93.550 184.235 94.225 184.395 ;
        RECT 94.685 184.315 95.905 184.485 ;
        RECT 93.550 183.445 93.760 184.235 ;
        RECT 94.685 184.225 94.855 184.315 ;
        RECT 93.930 183.445 94.280 184.065 ;
        RECT 94.450 184.055 94.855 184.225 ;
        RECT 94.450 183.275 94.620 184.055 ;
        RECT 94.790 183.605 95.010 183.885 ;
        RECT 95.190 183.775 95.730 184.145 ;
        RECT 96.075 184.065 96.245 184.655 ;
        RECT 96.465 184.235 96.770 185.375 ;
        RECT 96.940 184.185 97.195 185.065 ;
        RECT 96.075 184.035 96.815 184.065 ;
        RECT 94.790 183.435 95.320 183.605 ;
        RECT 93.100 183.015 93.450 183.185 ;
        RECT 93.670 182.995 94.620 183.275 ;
        RECT 94.790 182.825 94.980 183.265 ;
        RECT 95.150 183.205 95.320 183.435 ;
        RECT 95.490 183.375 95.730 183.775 ;
        RECT 95.900 183.735 96.815 184.035 ;
        RECT 95.900 183.560 96.225 183.735 ;
        RECT 95.900 183.205 96.220 183.560 ;
        RECT 96.985 183.535 97.195 184.185 ;
        RECT 95.150 183.035 96.220 183.205 ;
        RECT 96.465 182.825 96.770 183.285 ;
        RECT 96.940 183.005 97.195 183.535 ;
        RECT 97.375 184.185 97.630 185.065 ;
        RECT 97.800 184.235 98.105 185.375 ;
        RECT 98.445 184.995 98.775 185.375 ;
        RECT 98.955 184.825 99.125 185.115 ;
        RECT 99.295 184.915 99.545 185.375 ;
        RECT 98.325 184.655 99.125 184.825 ;
        RECT 99.715 184.865 100.585 185.205 ;
        RECT 97.375 183.535 97.585 184.185 ;
        RECT 98.325 184.065 98.495 184.655 ;
        RECT 99.715 184.485 99.885 184.865 ;
        RECT 100.820 184.745 100.990 185.205 ;
        RECT 101.160 184.915 101.530 185.375 ;
        RECT 101.825 184.775 101.995 185.115 ;
        RECT 102.165 184.945 102.495 185.375 ;
        RECT 102.730 184.775 102.900 185.115 ;
        RECT 98.665 184.315 99.885 184.485 ;
        RECT 100.055 184.405 100.515 184.695 ;
        RECT 100.820 184.575 101.380 184.745 ;
        RECT 101.825 184.605 102.900 184.775 ;
        RECT 103.070 184.875 103.750 185.205 ;
        RECT 103.965 184.875 104.215 185.205 ;
        RECT 104.385 184.915 104.635 185.375 ;
        RECT 101.210 184.435 101.380 184.575 ;
        RECT 100.055 184.395 101.020 184.405 ;
        RECT 99.715 184.225 99.885 184.315 ;
        RECT 100.345 184.235 101.020 184.395 ;
        RECT 97.755 184.035 98.495 184.065 ;
        RECT 97.755 183.735 98.670 184.035 ;
        RECT 98.345 183.560 98.670 183.735 ;
        RECT 97.375 183.005 97.630 183.535 ;
        RECT 97.800 182.825 98.105 183.285 ;
        RECT 98.350 183.205 98.670 183.560 ;
        RECT 98.840 183.775 99.380 184.145 ;
        RECT 99.715 184.055 100.120 184.225 ;
        RECT 98.840 183.375 99.080 183.775 ;
        RECT 99.560 183.605 99.780 183.885 ;
        RECT 99.250 183.435 99.780 183.605 ;
        RECT 99.250 183.205 99.420 183.435 ;
        RECT 99.950 183.275 100.120 184.055 ;
        RECT 100.290 183.445 100.640 184.065 ;
        RECT 100.810 183.445 101.020 184.235 ;
        RECT 101.210 184.265 102.710 184.435 ;
        RECT 101.210 183.575 101.380 184.265 ;
        RECT 103.070 184.095 103.240 184.875 ;
        RECT 104.045 184.745 104.215 184.875 ;
        RECT 101.550 183.925 103.240 184.095 ;
        RECT 103.410 184.315 103.875 184.705 ;
        RECT 104.045 184.575 104.440 184.745 ;
        RECT 101.550 183.745 101.720 183.925 ;
        RECT 98.350 183.035 99.420 183.205 ;
        RECT 99.590 182.825 99.780 183.265 ;
        RECT 99.950 182.995 100.900 183.275 ;
        RECT 101.210 183.185 101.470 183.575 ;
        RECT 101.890 183.505 102.680 183.755 ;
        RECT 101.120 183.015 101.470 183.185 ;
        RECT 101.680 182.825 102.010 183.285 ;
        RECT 102.885 183.215 103.055 183.925 ;
        RECT 103.410 183.725 103.580 184.315 ;
        RECT 103.225 183.505 103.580 183.725 ;
        RECT 103.750 183.505 104.100 184.125 ;
        RECT 104.270 183.215 104.440 184.575 ;
        RECT 104.805 184.405 105.130 185.190 ;
        RECT 104.610 183.355 105.070 184.405 ;
        RECT 102.885 183.045 103.740 183.215 ;
        RECT 103.945 183.045 104.440 183.215 ;
        RECT 104.610 182.825 104.940 183.185 ;
        RECT 105.300 183.085 105.470 185.205 ;
        RECT 105.640 184.875 105.970 185.375 ;
        RECT 106.140 184.705 106.395 185.205 ;
        RECT 105.645 184.535 106.395 184.705 ;
        RECT 105.645 183.545 105.875 184.535 ;
        RECT 106.045 183.715 106.395 184.365 ;
        RECT 107.490 184.285 111.000 185.375 ;
        RECT 111.170 184.285 112.380 185.375 ;
        RECT 107.490 183.765 109.180 184.285 ;
        RECT 109.350 183.595 111.000 184.115 ;
        RECT 111.170 183.745 111.690 184.285 ;
        RECT 105.645 183.375 106.395 183.545 ;
        RECT 105.640 182.825 105.970 183.205 ;
        RECT 106.140 183.085 106.395 183.375 ;
        RECT 107.490 182.825 111.000 183.595 ;
        RECT 111.860 183.575 112.380 184.115 ;
        RECT 111.170 182.825 112.380 183.575 ;
        RECT 18.165 182.655 112.465 182.825 ;
        RECT 18.250 181.905 19.460 182.655 ;
        RECT 18.250 181.365 18.770 181.905 ;
        RECT 20.090 181.885 21.760 182.655 ;
        RECT 21.930 181.930 22.220 182.655 ;
        RECT 22.850 181.885 25.440 182.655 ;
        RECT 25.615 182.110 30.960 182.655 ;
        RECT 31.135 182.110 36.480 182.655 ;
        RECT 36.655 182.110 42.000 182.655 ;
        RECT 42.175 182.110 47.520 182.655 ;
        RECT 18.940 181.195 19.460 181.735 ;
        RECT 18.250 180.105 19.460 181.195 ;
        RECT 20.090 181.195 20.840 181.715 ;
        RECT 21.010 181.365 21.760 181.885 ;
        RECT 20.090 180.105 21.760 181.195 ;
        RECT 21.930 180.105 22.220 181.270 ;
        RECT 22.850 181.195 24.060 181.715 ;
        RECT 24.230 181.365 25.440 181.885 ;
        RECT 22.850 180.105 25.440 181.195 ;
        RECT 27.205 180.540 27.555 181.790 ;
        RECT 29.035 181.280 29.375 182.110 ;
        RECT 32.725 180.540 33.075 181.790 ;
        RECT 34.555 181.280 34.895 182.110 ;
        RECT 38.245 180.540 38.595 181.790 ;
        RECT 40.075 181.280 40.415 182.110 ;
        RECT 43.765 180.540 44.115 181.790 ;
        RECT 45.595 181.280 45.935 182.110 ;
        RECT 47.690 181.930 47.980 182.655 ;
        RECT 48.150 181.885 51.660 182.655 ;
        RECT 51.835 182.110 57.180 182.655 ;
        RECT 25.615 180.105 30.960 180.540 ;
        RECT 31.135 180.105 36.480 180.540 ;
        RECT 36.655 180.105 42.000 180.540 ;
        RECT 42.175 180.105 47.520 180.540 ;
        RECT 47.690 180.105 47.980 181.270 ;
        RECT 48.150 181.195 49.840 181.715 ;
        RECT 50.010 181.365 51.660 181.885 ;
        RECT 48.150 180.105 51.660 181.195 ;
        RECT 53.425 180.540 53.775 181.790 ;
        RECT 55.255 181.280 55.595 182.110 ;
        RECT 57.435 182.085 57.610 182.485 ;
        RECT 57.780 182.275 58.110 182.655 ;
        RECT 58.355 182.155 58.585 182.485 ;
        RECT 57.435 181.915 58.065 182.085 ;
        RECT 57.895 181.745 58.065 181.915 ;
        RECT 57.350 181.065 57.715 181.745 ;
        RECT 57.895 181.415 58.245 181.745 ;
        RECT 57.895 180.895 58.065 181.415 ;
        RECT 57.435 180.725 58.065 180.895 ;
        RECT 58.415 180.865 58.585 182.155 ;
        RECT 58.785 181.045 59.065 182.320 ;
        RECT 59.290 182.315 59.560 182.320 ;
        RECT 59.250 182.145 59.560 182.315 ;
        RECT 60.020 182.275 60.350 182.655 ;
        RECT 60.520 182.400 60.855 182.445 ;
        RECT 59.290 181.045 59.560 182.145 ;
        RECT 59.750 181.045 60.090 182.075 ;
        RECT 60.520 181.935 60.860 182.400 ;
        RECT 60.260 181.415 60.520 181.745 ;
        RECT 60.260 180.865 60.430 181.415 ;
        RECT 60.690 181.245 60.860 181.935 ;
        RECT 51.835 180.105 57.180 180.540 ;
        RECT 57.435 180.275 57.610 180.725 ;
        RECT 58.415 180.695 60.430 180.865 ;
        RECT 57.780 180.105 58.110 180.545 ;
        RECT 58.415 180.275 58.585 180.695 ;
        RECT 58.820 180.105 59.490 180.515 ;
        RECT 59.705 180.275 59.875 180.695 ;
        RECT 60.075 180.105 60.405 180.515 ;
        RECT 60.600 180.275 60.860 181.245 ;
        RECT 61.030 182.155 61.290 182.485 ;
        RECT 61.600 182.275 61.930 182.655 ;
        RECT 62.110 182.315 63.590 182.485 ;
        RECT 61.030 181.455 61.200 182.155 ;
        RECT 62.110 181.985 62.510 182.315 ;
        RECT 61.550 181.795 61.760 181.975 ;
        RECT 61.550 181.625 62.170 181.795 ;
        RECT 62.340 181.505 62.510 181.985 ;
        RECT 62.700 181.815 63.250 182.145 ;
        RECT 61.030 181.285 62.160 181.455 ;
        RECT 62.340 181.335 62.910 181.505 ;
        RECT 61.030 180.605 61.200 181.285 ;
        RECT 61.990 181.165 62.160 181.285 ;
        RECT 61.370 180.785 61.720 181.115 ;
        RECT 61.990 180.995 62.570 181.165 ;
        RECT 62.740 180.825 62.910 181.335 ;
        RECT 62.170 180.655 62.910 180.825 ;
        RECT 63.080 180.825 63.250 181.815 ;
        RECT 63.420 181.415 63.590 182.315 ;
        RECT 63.840 181.745 64.025 182.325 ;
        RECT 64.295 181.745 64.490 182.320 ;
        RECT 64.700 182.275 65.030 182.655 ;
        RECT 63.840 181.415 64.070 181.745 ;
        RECT 64.295 181.415 64.550 181.745 ;
        RECT 63.840 181.105 64.025 181.415 ;
        RECT 64.295 181.105 64.490 181.415 ;
        RECT 64.860 180.825 65.030 181.745 ;
        RECT 63.080 180.655 65.030 180.825 ;
        RECT 61.030 180.275 61.290 180.605 ;
        RECT 61.600 180.105 61.930 180.485 ;
        RECT 62.170 180.275 62.360 180.655 ;
        RECT 62.610 180.105 62.940 180.485 ;
        RECT 63.150 180.275 63.320 180.655 ;
        RECT 63.515 180.105 63.845 180.485 ;
        RECT 64.105 180.275 64.275 180.655 ;
        RECT 64.700 180.105 65.030 180.485 ;
        RECT 65.200 180.275 65.460 182.485 ;
        RECT 65.630 182.155 65.890 182.485 ;
        RECT 66.100 182.175 66.375 182.655 ;
        RECT 65.630 181.245 65.800 182.155 ;
        RECT 66.585 182.085 66.790 182.485 ;
        RECT 66.960 182.255 67.295 182.655 ;
        RECT 67.635 182.145 67.875 182.655 ;
        RECT 68.055 182.145 68.335 182.475 ;
        RECT 68.565 182.145 68.780 182.655 ;
        RECT 65.970 181.415 66.330 181.995 ;
        RECT 66.585 181.915 67.270 182.085 ;
        RECT 66.510 181.245 66.760 181.745 ;
        RECT 65.630 181.075 66.760 181.245 ;
        RECT 65.630 180.305 65.900 181.075 ;
        RECT 66.930 180.885 67.270 181.915 ;
        RECT 67.530 181.415 67.885 181.975 ;
        RECT 68.055 181.245 68.225 182.145 ;
        RECT 68.395 181.415 68.660 181.975 ;
        RECT 68.950 181.915 69.565 182.485 ;
        RECT 68.910 181.245 69.080 181.745 ;
        RECT 67.655 181.075 69.080 181.245 ;
        RECT 67.655 180.900 68.045 181.075 ;
        RECT 66.070 180.105 66.400 180.885 ;
        RECT 66.605 180.710 67.270 180.885 ;
        RECT 66.605 180.305 66.790 180.710 ;
        RECT 66.960 180.105 67.295 180.530 ;
        RECT 68.530 180.105 68.860 180.905 ;
        RECT 69.250 180.895 69.565 181.915 ;
        RECT 69.030 180.275 69.565 180.895 ;
        RECT 69.770 182.005 70.030 182.485 ;
        RECT 70.200 182.115 70.450 182.655 ;
        RECT 69.770 180.975 69.940 182.005 ;
        RECT 70.620 181.950 70.840 182.435 ;
        RECT 70.110 181.355 70.340 181.750 ;
        RECT 70.510 181.525 70.840 181.950 ;
        RECT 71.010 182.275 71.900 182.445 ;
        RECT 71.010 181.550 71.180 182.275 ;
        RECT 71.350 181.720 71.900 182.105 ;
        RECT 72.070 181.905 73.280 182.655 ;
        RECT 73.450 181.930 73.740 182.655 ;
        RECT 71.010 181.480 71.900 181.550 ;
        RECT 71.005 181.455 71.900 181.480 ;
        RECT 70.995 181.440 71.900 181.455 ;
        RECT 70.990 181.425 71.900 181.440 ;
        RECT 70.980 181.420 71.900 181.425 ;
        RECT 70.975 181.410 71.900 181.420 ;
        RECT 70.970 181.400 71.900 181.410 ;
        RECT 70.960 181.395 71.900 181.400 ;
        RECT 70.950 181.385 71.900 181.395 ;
        RECT 70.940 181.380 71.900 181.385 ;
        RECT 70.940 181.375 71.275 181.380 ;
        RECT 70.925 181.370 71.275 181.375 ;
        RECT 70.910 181.360 71.275 181.370 ;
        RECT 70.885 181.355 71.275 181.360 ;
        RECT 70.110 181.350 71.275 181.355 ;
        RECT 70.110 181.315 71.245 181.350 ;
        RECT 70.110 181.290 71.210 181.315 ;
        RECT 70.110 181.260 71.180 181.290 ;
        RECT 70.110 181.230 71.160 181.260 ;
        RECT 70.110 181.200 71.140 181.230 ;
        RECT 70.110 181.190 71.070 181.200 ;
        RECT 70.110 181.180 71.045 181.190 ;
        RECT 70.110 181.165 71.025 181.180 ;
        RECT 70.110 181.150 71.005 181.165 ;
        RECT 70.215 181.140 71.000 181.150 ;
        RECT 70.215 181.105 70.985 181.140 ;
        RECT 69.770 180.275 70.045 180.975 ;
        RECT 70.215 180.855 70.970 181.105 ;
        RECT 71.140 180.785 71.470 181.030 ;
        RECT 71.640 180.930 71.900 181.380 ;
        RECT 72.070 181.195 72.590 181.735 ;
        RECT 72.760 181.365 73.280 181.905 ;
        RECT 73.910 181.885 76.500 182.655 ;
        RECT 71.285 180.760 71.470 180.785 ;
        RECT 71.285 180.660 71.900 180.760 ;
        RECT 70.215 180.105 70.470 180.650 ;
        RECT 70.640 180.275 71.120 180.615 ;
        RECT 71.295 180.105 71.900 180.660 ;
        RECT 72.070 180.105 73.280 181.195 ;
        RECT 73.450 180.105 73.740 181.270 ;
        RECT 73.910 181.195 75.120 181.715 ;
        RECT 75.290 181.365 76.500 181.885 ;
        RECT 76.710 181.835 76.940 182.655 ;
        RECT 77.110 181.855 77.440 182.485 ;
        RECT 76.690 181.415 77.020 181.665 ;
        RECT 77.190 181.255 77.440 181.855 ;
        RECT 77.610 181.835 77.820 182.655 ;
        RECT 78.055 181.945 78.310 182.475 ;
        RECT 78.480 182.195 78.785 182.655 ;
        RECT 79.030 182.275 80.100 182.445 ;
        RECT 73.910 180.105 76.500 181.195 ;
        RECT 76.710 180.105 76.940 181.245 ;
        RECT 77.110 180.275 77.440 181.255 ;
        RECT 78.055 181.295 78.265 181.945 ;
        RECT 79.030 181.920 79.350 182.275 ;
        RECT 79.025 181.745 79.350 181.920 ;
        RECT 78.435 181.445 79.350 181.745 ;
        RECT 79.520 181.705 79.760 182.105 ;
        RECT 79.930 182.045 80.100 182.275 ;
        RECT 80.270 182.215 80.460 182.655 ;
        RECT 80.630 182.205 81.580 182.485 ;
        RECT 81.800 182.295 82.150 182.465 ;
        RECT 79.930 181.875 80.460 182.045 ;
        RECT 78.435 181.415 79.175 181.445 ;
        RECT 77.610 180.105 77.820 181.245 ;
        RECT 78.055 180.415 78.310 181.295 ;
        RECT 78.480 180.105 78.785 181.245 ;
        RECT 79.005 180.825 79.175 181.415 ;
        RECT 79.520 181.335 80.060 181.705 ;
        RECT 80.240 181.595 80.460 181.875 ;
        RECT 80.630 181.425 80.800 182.205 ;
        RECT 80.395 181.255 80.800 181.425 ;
        RECT 80.970 181.415 81.320 182.035 ;
        RECT 80.395 181.165 80.565 181.255 ;
        RECT 81.490 181.245 81.700 182.035 ;
        RECT 79.345 180.995 80.565 181.165 ;
        RECT 81.025 181.085 81.700 181.245 ;
        RECT 79.005 180.655 79.805 180.825 ;
        RECT 79.125 180.105 79.455 180.485 ;
        RECT 79.635 180.365 79.805 180.655 ;
        RECT 80.395 180.615 80.565 180.995 ;
        RECT 80.735 181.075 81.700 181.085 ;
        RECT 81.890 181.905 82.150 182.295 ;
        RECT 82.360 182.195 82.690 182.655 ;
        RECT 83.565 182.265 84.420 182.435 ;
        RECT 84.625 182.265 85.120 182.435 ;
        RECT 85.290 182.295 85.620 182.655 ;
        RECT 81.890 181.215 82.060 181.905 ;
        RECT 82.230 181.555 82.400 181.735 ;
        RECT 82.570 181.725 83.360 181.975 ;
        RECT 83.565 181.555 83.735 182.265 ;
        RECT 83.905 181.755 84.260 181.975 ;
        RECT 82.230 181.385 83.920 181.555 ;
        RECT 80.735 180.785 81.195 181.075 ;
        RECT 81.890 181.045 83.390 181.215 ;
        RECT 81.890 180.905 82.060 181.045 ;
        RECT 81.500 180.735 82.060 180.905 ;
        RECT 79.975 180.105 80.225 180.565 ;
        RECT 80.395 180.275 81.265 180.615 ;
        RECT 81.500 180.275 81.670 180.735 ;
        RECT 82.505 180.705 83.580 180.875 ;
        RECT 81.840 180.105 82.210 180.565 ;
        RECT 82.505 180.365 82.675 180.705 ;
        RECT 82.845 180.105 83.175 180.535 ;
        RECT 83.410 180.365 83.580 180.705 ;
        RECT 83.750 180.605 83.920 181.385 ;
        RECT 84.090 181.165 84.260 181.755 ;
        RECT 84.430 181.355 84.780 181.975 ;
        RECT 84.090 180.775 84.555 181.165 ;
        RECT 84.950 180.905 85.120 182.265 ;
        RECT 85.290 181.075 85.750 182.125 ;
        RECT 84.725 180.735 85.120 180.905 ;
        RECT 84.725 180.605 84.895 180.735 ;
        RECT 83.750 180.275 84.430 180.605 ;
        RECT 84.645 180.275 84.895 180.605 ;
        RECT 85.065 180.105 85.315 180.565 ;
        RECT 85.485 180.290 85.810 181.075 ;
        RECT 85.980 180.275 86.150 182.395 ;
        RECT 86.320 182.275 86.650 182.655 ;
        RECT 86.820 182.105 87.075 182.395 ;
        RECT 86.325 181.935 87.075 182.105 ;
        RECT 86.325 180.945 86.555 181.935 ;
        RECT 87.710 181.885 89.380 182.655 ;
        RECT 86.725 181.115 87.075 181.765 ;
        RECT 87.710 181.195 88.460 181.715 ;
        RECT 88.630 181.365 89.380 181.885 ;
        RECT 89.550 181.980 89.810 182.485 ;
        RECT 89.990 182.275 90.320 182.655 ;
        RECT 90.500 182.105 90.670 182.485 ;
        RECT 86.325 180.775 87.075 180.945 ;
        RECT 86.320 180.105 86.650 180.605 ;
        RECT 86.820 180.275 87.075 180.775 ;
        RECT 87.710 180.105 89.380 181.195 ;
        RECT 89.550 181.180 89.720 181.980 ;
        RECT 90.005 181.935 90.670 182.105 ;
        RECT 90.005 181.680 90.175 181.935 ;
        RECT 90.935 181.915 91.190 182.485 ;
        RECT 91.360 182.255 91.690 182.655 ;
        RECT 92.115 182.120 92.645 182.485 ;
        RECT 92.115 182.085 92.290 182.120 ;
        RECT 91.360 181.915 92.290 182.085 ;
        RECT 89.890 181.350 90.175 181.680 ;
        RECT 90.410 181.385 90.740 181.755 ;
        RECT 90.005 181.205 90.175 181.350 ;
        RECT 90.935 181.245 91.105 181.915 ;
        RECT 91.360 181.745 91.530 181.915 ;
        RECT 91.275 181.415 91.530 181.745 ;
        RECT 91.755 181.415 91.950 181.745 ;
        RECT 89.550 180.275 89.820 181.180 ;
        RECT 90.005 181.035 90.670 181.205 ;
        RECT 89.990 180.105 90.320 180.865 ;
        RECT 90.500 180.275 90.670 181.035 ;
        RECT 90.935 180.275 91.270 181.245 ;
        RECT 91.440 180.105 91.610 181.245 ;
        RECT 91.780 180.445 91.950 181.415 ;
        RECT 92.120 180.785 92.290 181.915 ;
        RECT 92.460 181.125 92.630 181.925 ;
        RECT 92.835 181.635 93.110 182.485 ;
        RECT 92.830 181.465 93.110 181.635 ;
        RECT 92.835 181.325 93.110 181.465 ;
        RECT 93.280 181.125 93.470 182.485 ;
        RECT 93.650 182.120 94.160 182.655 ;
        RECT 94.380 181.845 94.625 182.450 ;
        RECT 95.345 181.845 95.590 182.450 ;
        RECT 95.810 182.120 96.320 182.655 ;
        RECT 93.670 181.675 94.900 181.845 ;
        RECT 92.460 180.955 93.470 181.125 ;
        RECT 93.640 181.110 94.390 181.300 ;
        RECT 92.120 180.615 93.245 180.785 ;
        RECT 93.640 180.445 93.810 181.110 ;
        RECT 94.560 180.865 94.900 181.675 ;
        RECT 91.780 180.275 93.810 180.445 ;
        RECT 93.980 180.105 94.150 180.865 ;
        RECT 94.385 180.455 94.900 180.865 ;
        RECT 95.070 181.675 96.300 181.845 ;
        RECT 95.070 180.865 95.410 181.675 ;
        RECT 95.580 181.110 96.330 181.300 ;
        RECT 95.070 180.455 95.585 180.865 ;
        RECT 95.820 180.105 95.990 180.865 ;
        RECT 96.160 180.445 96.330 181.110 ;
        RECT 96.500 181.125 96.690 182.485 ;
        RECT 96.860 181.975 97.135 182.485 ;
        RECT 97.325 182.120 97.855 182.485 ;
        RECT 98.280 182.255 98.610 182.655 ;
        RECT 97.680 182.085 97.855 182.120 ;
        RECT 96.860 181.805 97.140 181.975 ;
        RECT 96.860 181.325 97.135 181.805 ;
        RECT 97.340 181.125 97.510 181.925 ;
        RECT 96.500 180.955 97.510 181.125 ;
        RECT 97.680 181.915 98.610 182.085 ;
        RECT 98.780 181.915 99.035 182.485 ;
        RECT 99.210 181.930 99.500 182.655 ;
        RECT 99.760 182.105 99.930 182.485 ;
        RECT 100.110 182.275 100.440 182.655 ;
        RECT 99.760 181.935 100.425 182.105 ;
        RECT 100.620 181.980 100.880 182.485 ;
        RECT 97.680 180.785 97.850 181.915 ;
        RECT 98.440 181.745 98.610 181.915 ;
        RECT 96.725 180.615 97.850 180.785 ;
        RECT 98.020 181.415 98.215 181.745 ;
        RECT 98.440 181.415 98.695 181.745 ;
        RECT 98.020 180.445 98.190 181.415 ;
        RECT 98.865 181.245 99.035 181.915 ;
        RECT 99.690 181.385 100.020 181.755 ;
        RECT 100.255 181.680 100.425 181.935 ;
        RECT 100.255 181.350 100.540 181.680 ;
        RECT 96.160 180.275 98.190 180.445 ;
        RECT 98.360 180.105 98.530 181.245 ;
        RECT 98.700 180.275 99.035 181.245 ;
        RECT 99.210 180.105 99.500 181.270 ;
        RECT 100.255 181.205 100.425 181.350 ;
        RECT 99.760 181.035 100.425 181.205 ;
        RECT 100.710 181.180 100.880 181.980 ;
        RECT 101.970 181.885 105.480 182.655 ;
        RECT 105.655 182.110 111.000 182.655 ;
        RECT 99.760 180.275 99.930 181.035 ;
        RECT 100.110 180.105 100.440 180.865 ;
        RECT 100.610 180.275 100.880 181.180 ;
        RECT 101.970 181.195 103.660 181.715 ;
        RECT 103.830 181.365 105.480 181.885 ;
        RECT 101.970 180.105 105.480 181.195 ;
        RECT 107.245 180.540 107.595 181.790 ;
        RECT 109.075 181.280 109.415 182.110 ;
        RECT 111.170 181.905 112.380 182.655 ;
        RECT 111.170 181.195 111.690 181.735 ;
        RECT 111.860 181.365 112.380 181.905 ;
        RECT 105.655 180.105 111.000 180.540 ;
        RECT 111.170 180.105 112.380 181.195 ;
        RECT 18.165 179.935 112.465 180.105 ;
        RECT 18.250 178.845 19.460 179.935 ;
        RECT 18.250 178.135 18.770 178.675 ;
        RECT 18.940 178.305 19.460 178.845 ;
        RECT 20.090 178.845 23.600 179.935 ;
        RECT 23.775 179.500 29.120 179.935 ;
        RECT 29.295 179.500 34.640 179.935 ;
        RECT 20.090 178.325 21.780 178.845 ;
        RECT 21.950 178.155 23.600 178.675 ;
        RECT 25.365 178.250 25.715 179.500 ;
        RECT 18.250 177.385 19.460 178.135 ;
        RECT 20.090 177.385 23.600 178.155 ;
        RECT 27.195 177.930 27.535 178.760 ;
        RECT 30.885 178.250 31.235 179.500 ;
        RECT 34.810 178.770 35.100 179.935 ;
        RECT 35.270 178.845 36.940 179.935 ;
        RECT 37.115 179.500 42.460 179.935 ;
        RECT 32.715 177.930 33.055 178.760 ;
        RECT 35.270 178.325 36.020 178.845 ;
        RECT 36.190 178.155 36.940 178.675 ;
        RECT 38.705 178.250 39.055 179.500 ;
        RECT 42.690 178.795 42.900 179.935 ;
        RECT 43.070 178.785 43.400 179.765 ;
        RECT 43.570 178.795 43.800 179.935 ;
        RECT 44.385 178.955 44.640 179.625 ;
        RECT 44.820 179.135 45.105 179.935 ;
        RECT 45.285 179.215 45.615 179.725 ;
        RECT 23.775 177.385 29.120 177.930 ;
        RECT 29.295 177.385 34.640 177.930 ;
        RECT 34.810 177.385 35.100 178.110 ;
        RECT 35.270 177.385 36.940 178.155 ;
        RECT 40.535 177.930 40.875 178.760 ;
        RECT 37.115 177.385 42.460 177.930 ;
        RECT 42.690 177.385 42.900 178.205 ;
        RECT 43.070 178.185 43.320 178.785 ;
        RECT 43.490 178.375 43.820 178.625 ;
        RECT 43.070 177.555 43.400 178.185 ;
        RECT 43.570 177.385 43.800 178.205 ;
        RECT 44.385 178.095 44.565 178.955 ;
        RECT 45.285 178.625 45.535 179.215 ;
        RECT 45.885 179.065 46.055 179.675 ;
        RECT 46.225 179.245 46.555 179.935 ;
        RECT 46.785 179.385 47.025 179.675 ;
        RECT 47.225 179.555 47.645 179.935 ;
        RECT 47.825 179.465 48.455 179.715 ;
        RECT 48.925 179.555 49.255 179.935 ;
        RECT 47.825 179.385 47.995 179.465 ;
        RECT 49.425 179.385 49.595 179.675 ;
        RECT 49.775 179.555 50.155 179.935 ;
        RECT 50.395 179.550 51.225 179.720 ;
        RECT 46.785 179.215 47.995 179.385 ;
        RECT 44.735 178.295 45.535 178.625 ;
        RECT 44.385 177.895 44.640 178.095 ;
        RECT 44.300 177.725 44.640 177.895 ;
        RECT 44.385 177.565 44.640 177.725 ;
        RECT 44.820 177.385 45.105 177.845 ;
        RECT 45.285 177.645 45.535 178.295 ;
        RECT 45.735 179.045 46.055 179.065 ;
        RECT 45.735 178.875 47.655 179.045 ;
        RECT 45.735 177.980 45.925 178.875 ;
        RECT 47.825 178.705 47.995 179.215 ;
        RECT 48.165 178.955 48.685 179.265 ;
        RECT 46.095 178.535 47.995 178.705 ;
        RECT 46.095 178.475 46.425 178.535 ;
        RECT 46.575 178.305 46.905 178.365 ;
        RECT 46.245 178.035 46.905 178.305 ;
        RECT 45.735 177.650 46.055 177.980 ;
        RECT 46.235 177.385 46.895 177.865 ;
        RECT 47.095 177.775 47.265 178.535 ;
        RECT 48.165 178.365 48.345 178.775 ;
        RECT 47.435 178.195 47.765 178.315 ;
        RECT 48.515 178.195 48.685 178.955 ;
        RECT 47.435 178.025 48.685 178.195 ;
        RECT 48.855 179.135 50.225 179.385 ;
        RECT 48.855 178.365 49.045 179.135 ;
        RECT 49.975 178.875 50.225 179.135 ;
        RECT 49.215 178.705 49.465 178.865 ;
        RECT 50.395 178.705 50.565 179.550 ;
        RECT 51.460 179.265 51.630 179.765 ;
        RECT 51.800 179.435 52.130 179.935 ;
        RECT 50.735 178.875 51.235 179.255 ;
        RECT 51.460 179.095 52.155 179.265 ;
        RECT 49.215 178.535 50.565 178.705 ;
        RECT 50.145 178.495 50.565 178.535 ;
        RECT 48.855 178.025 49.275 178.365 ;
        RECT 49.565 178.035 49.975 178.365 ;
        RECT 47.095 177.605 47.945 177.775 ;
        RECT 48.505 177.385 48.825 177.845 ;
        RECT 49.025 177.595 49.275 178.025 ;
        RECT 49.565 177.385 49.975 177.825 ;
        RECT 50.145 177.765 50.315 178.495 ;
        RECT 50.485 177.945 50.835 178.315 ;
        RECT 51.015 178.005 51.235 178.875 ;
        RECT 51.405 178.305 51.815 178.925 ;
        RECT 51.985 178.125 52.155 179.095 ;
        RECT 51.460 177.935 52.155 178.125 ;
        RECT 50.145 177.565 51.160 177.765 ;
        RECT 51.460 177.605 51.630 177.935 ;
        RECT 51.800 177.385 52.130 177.765 ;
        RECT 52.345 177.645 52.570 179.765 ;
        RECT 52.740 179.435 53.070 179.935 ;
        RECT 53.240 179.265 53.410 179.765 ;
        RECT 52.745 179.095 53.410 179.265 ;
        RECT 52.745 178.105 52.975 179.095 ;
        RECT 53.145 178.275 53.495 178.925 ;
        RECT 53.670 178.845 54.880 179.935 ;
        RECT 55.050 178.845 58.560 179.935 ;
        RECT 58.730 178.965 59.000 179.735 ;
        RECT 59.170 179.155 59.500 179.935 ;
        RECT 59.705 179.330 59.890 179.735 ;
        RECT 60.060 179.510 60.395 179.935 ;
        RECT 59.705 179.155 60.370 179.330 ;
        RECT 53.670 178.305 54.190 178.845 ;
        RECT 54.360 178.135 54.880 178.675 ;
        RECT 55.050 178.325 56.740 178.845 ;
        RECT 58.730 178.795 59.860 178.965 ;
        RECT 56.910 178.155 58.560 178.675 ;
        RECT 52.745 177.935 53.410 178.105 ;
        RECT 52.740 177.385 53.070 177.765 ;
        RECT 53.240 177.645 53.410 177.935 ;
        RECT 53.670 177.385 54.880 178.135 ;
        RECT 55.050 177.385 58.560 178.155 ;
        RECT 58.730 177.885 58.900 178.795 ;
        RECT 59.070 178.045 59.430 178.625 ;
        RECT 59.610 178.295 59.860 178.795 ;
        RECT 60.030 178.125 60.370 179.155 ;
        RECT 60.570 178.770 60.860 179.935 ;
        RECT 61.950 179.380 62.555 179.935 ;
        RECT 62.730 179.425 63.210 179.765 ;
        RECT 63.380 179.390 63.635 179.935 ;
        RECT 61.950 179.280 62.565 179.380 ;
        RECT 62.380 179.255 62.565 179.280 ;
        RECT 61.950 178.660 62.210 179.110 ;
        RECT 62.380 179.010 62.710 179.255 ;
        RECT 62.880 178.935 63.635 179.185 ;
        RECT 63.805 179.065 64.080 179.765 ;
        RECT 62.865 178.900 63.635 178.935 ;
        RECT 62.850 178.890 63.635 178.900 ;
        RECT 62.845 178.875 63.740 178.890 ;
        RECT 62.825 178.860 63.740 178.875 ;
        RECT 62.805 178.850 63.740 178.860 ;
        RECT 62.780 178.840 63.740 178.850 ;
        RECT 62.710 178.810 63.740 178.840 ;
        RECT 62.690 178.780 63.740 178.810 ;
        RECT 62.670 178.750 63.740 178.780 ;
        RECT 62.640 178.725 63.740 178.750 ;
        RECT 62.605 178.690 63.740 178.725 ;
        RECT 62.575 178.685 63.740 178.690 ;
        RECT 62.575 178.680 62.965 178.685 ;
        RECT 62.575 178.670 62.940 178.680 ;
        RECT 62.575 178.665 62.925 178.670 ;
        RECT 62.575 178.660 62.910 178.665 ;
        RECT 61.950 178.655 62.910 178.660 ;
        RECT 61.950 178.645 62.900 178.655 ;
        RECT 61.950 178.640 62.890 178.645 ;
        RECT 61.950 178.630 62.880 178.640 ;
        RECT 61.950 178.620 62.875 178.630 ;
        RECT 61.950 178.615 62.870 178.620 ;
        RECT 61.950 178.600 62.860 178.615 ;
        RECT 61.950 178.585 62.855 178.600 ;
        RECT 61.950 178.560 62.845 178.585 ;
        RECT 61.950 178.490 62.840 178.560 ;
        RECT 59.685 177.955 60.370 178.125 ;
        RECT 58.730 177.555 58.990 177.885 ;
        RECT 59.200 177.385 59.475 177.865 ;
        RECT 59.685 177.555 59.890 177.955 ;
        RECT 60.060 177.385 60.395 177.785 ;
        RECT 60.570 177.385 60.860 178.110 ;
        RECT 61.950 177.935 62.500 178.320 ;
        RECT 62.670 177.765 62.840 178.490 ;
        RECT 61.950 177.595 62.840 177.765 ;
        RECT 63.010 178.090 63.340 178.515 ;
        RECT 63.510 178.290 63.740 178.685 ;
        RECT 63.010 177.605 63.230 178.090 ;
        RECT 63.910 178.035 64.080 179.065 ;
        RECT 63.400 177.385 63.650 177.925 ;
        RECT 63.820 177.555 64.080 178.035 ;
        RECT 64.260 178.875 64.590 179.725 ;
        RECT 64.260 178.110 64.450 178.875 ;
        RECT 64.760 178.795 65.010 179.935 ;
        RECT 65.200 179.295 65.450 179.715 ;
        RECT 65.680 179.465 66.010 179.935 ;
        RECT 66.240 179.295 66.490 179.715 ;
        RECT 65.200 179.125 66.490 179.295 ;
        RECT 66.670 179.295 67.000 179.725 ;
        RECT 66.670 179.125 67.125 179.295 ;
        RECT 65.190 178.625 65.405 178.955 ;
        RECT 64.620 178.295 64.930 178.625 ;
        RECT 65.100 178.295 65.405 178.625 ;
        RECT 65.580 178.295 65.865 178.955 ;
        RECT 66.060 178.295 66.325 178.955 ;
        RECT 66.540 178.295 66.785 178.955 ;
        RECT 64.760 178.125 64.930 178.295 ;
        RECT 66.955 178.125 67.125 179.125 ;
        RECT 64.260 177.600 64.590 178.110 ;
        RECT 64.760 177.955 67.125 178.125 ;
        RECT 67.470 178.860 67.740 179.765 ;
        RECT 67.910 179.175 68.240 179.935 ;
        RECT 68.420 179.005 68.590 179.765 ;
        RECT 67.470 178.060 67.640 178.860 ;
        RECT 67.925 178.835 68.590 179.005 ;
        RECT 67.925 178.690 68.095 178.835 ;
        RECT 68.850 178.795 69.130 179.935 ;
        RECT 69.300 178.785 69.630 179.765 ;
        RECT 69.800 178.795 70.060 179.935 ;
        RECT 71.150 178.845 74.660 179.935 ;
        RECT 75.205 178.955 75.460 179.625 ;
        RECT 75.640 179.135 75.925 179.935 ;
        RECT 76.105 179.215 76.435 179.725 ;
        RECT 67.810 178.360 68.095 178.690 ;
        RECT 67.925 178.105 68.095 178.360 ;
        RECT 68.330 178.285 68.660 178.655 ;
        RECT 68.860 178.355 69.195 178.625 ;
        RECT 69.365 178.185 69.535 178.785 ;
        RECT 69.705 178.375 70.040 178.625 ;
        RECT 71.150 178.325 72.840 178.845 ;
        RECT 64.760 177.385 65.090 177.785 ;
        RECT 66.140 177.615 66.470 177.955 ;
        RECT 66.640 177.385 66.970 177.785 ;
        RECT 67.470 177.555 67.730 178.060 ;
        RECT 67.925 177.935 68.590 178.105 ;
        RECT 67.910 177.385 68.240 177.765 ;
        RECT 68.420 177.555 68.590 177.935 ;
        RECT 68.850 177.385 69.160 178.185 ;
        RECT 69.365 177.555 70.060 178.185 ;
        RECT 73.010 178.155 74.660 178.675 ;
        RECT 75.205 178.235 75.385 178.955 ;
        RECT 76.105 178.625 76.355 179.215 ;
        RECT 76.705 179.065 76.875 179.675 ;
        RECT 77.045 179.245 77.375 179.935 ;
        RECT 77.605 179.385 77.845 179.675 ;
        RECT 78.045 179.555 78.465 179.935 ;
        RECT 78.645 179.465 79.275 179.715 ;
        RECT 79.745 179.555 80.075 179.935 ;
        RECT 78.645 179.385 78.815 179.465 ;
        RECT 80.245 179.385 80.415 179.675 ;
        RECT 80.595 179.555 80.975 179.935 ;
        RECT 81.215 179.550 82.045 179.720 ;
        RECT 77.605 179.215 78.815 179.385 ;
        RECT 75.555 178.295 76.355 178.625 ;
        RECT 71.150 177.385 74.660 178.155 ;
        RECT 75.120 178.095 75.385 178.235 ;
        RECT 75.120 178.065 75.460 178.095 ;
        RECT 75.205 177.565 75.460 178.065 ;
        RECT 75.640 177.385 75.925 177.845 ;
        RECT 76.105 177.645 76.355 178.295 ;
        RECT 76.555 179.045 76.875 179.065 ;
        RECT 76.555 178.875 78.475 179.045 ;
        RECT 76.555 177.980 76.745 178.875 ;
        RECT 78.645 178.705 78.815 179.215 ;
        RECT 78.985 178.955 79.505 179.265 ;
        RECT 76.915 178.535 78.815 178.705 ;
        RECT 76.915 178.475 77.245 178.535 ;
        RECT 77.395 178.305 77.725 178.365 ;
        RECT 77.065 178.035 77.725 178.305 ;
        RECT 76.555 177.650 76.875 177.980 ;
        RECT 77.055 177.385 77.715 177.865 ;
        RECT 77.915 177.775 78.085 178.535 ;
        RECT 78.985 178.365 79.165 178.775 ;
        RECT 78.255 178.195 78.585 178.315 ;
        RECT 79.335 178.195 79.505 178.955 ;
        RECT 78.255 178.025 79.505 178.195 ;
        RECT 79.675 179.135 81.045 179.385 ;
        RECT 79.675 178.365 79.865 179.135 ;
        RECT 80.795 178.875 81.045 179.135 ;
        RECT 80.035 178.705 80.285 178.865 ;
        RECT 81.215 178.705 81.385 179.550 ;
        RECT 82.280 179.265 82.450 179.765 ;
        RECT 82.620 179.435 82.950 179.935 ;
        RECT 81.555 178.875 82.055 179.255 ;
        RECT 82.280 179.095 82.975 179.265 ;
        RECT 80.035 178.535 81.385 178.705 ;
        RECT 80.965 178.495 81.385 178.535 ;
        RECT 79.675 178.025 80.095 178.365 ;
        RECT 80.385 178.035 80.795 178.365 ;
        RECT 77.915 177.605 78.765 177.775 ;
        RECT 79.325 177.385 79.645 177.845 ;
        RECT 79.845 177.595 80.095 178.025 ;
        RECT 80.385 177.385 80.795 177.825 ;
        RECT 80.965 177.765 81.135 178.495 ;
        RECT 81.305 177.945 81.655 178.315 ;
        RECT 81.835 178.005 82.055 178.875 ;
        RECT 82.225 178.305 82.635 178.925 ;
        RECT 82.805 178.125 82.975 179.095 ;
        RECT 82.280 177.935 82.975 178.125 ;
        RECT 80.965 177.565 81.980 177.765 ;
        RECT 82.280 177.605 82.450 177.935 ;
        RECT 82.620 177.385 82.950 177.765 ;
        RECT 83.165 177.645 83.390 179.765 ;
        RECT 83.560 179.435 83.890 179.935 ;
        RECT 84.060 179.265 84.230 179.765 ;
        RECT 83.565 179.095 84.230 179.265 ;
        RECT 83.565 178.105 83.795 179.095 ;
        RECT 83.965 178.275 84.315 178.925 ;
        RECT 84.490 178.860 84.760 179.765 ;
        RECT 84.930 179.175 85.260 179.935 ;
        RECT 85.440 179.005 85.610 179.765 ;
        RECT 83.565 177.935 84.230 178.105 ;
        RECT 83.560 177.385 83.890 177.765 ;
        RECT 84.060 177.645 84.230 177.935 ;
        RECT 84.490 178.060 84.660 178.860 ;
        RECT 84.945 178.835 85.610 179.005 ;
        RECT 84.945 178.690 85.115 178.835 ;
        RECT 86.330 178.770 86.620 179.935 ;
        RECT 86.795 179.500 92.140 179.935 ;
        RECT 84.830 178.360 85.115 178.690 ;
        RECT 84.945 178.105 85.115 178.360 ;
        RECT 85.350 178.285 85.680 178.655 ;
        RECT 88.385 178.250 88.735 179.500 ;
        RECT 92.350 178.795 92.580 179.935 ;
        RECT 92.750 178.785 93.080 179.765 ;
        RECT 93.250 178.795 93.460 179.935 ;
        RECT 84.490 177.555 84.750 178.060 ;
        RECT 84.945 177.935 85.610 178.105 ;
        RECT 84.930 177.385 85.260 177.765 ;
        RECT 85.440 177.555 85.610 177.935 ;
        RECT 86.330 177.385 86.620 178.110 ;
        RECT 90.215 177.930 90.555 178.760 ;
        RECT 92.330 178.375 92.660 178.625 ;
        RECT 86.795 177.385 92.140 177.930 ;
        RECT 92.350 177.385 92.580 178.205 ;
        RECT 92.830 178.185 93.080 178.785 ;
        RECT 93.695 178.745 93.950 179.625 ;
        RECT 94.120 178.795 94.425 179.935 ;
        RECT 94.765 179.555 95.095 179.935 ;
        RECT 95.275 179.385 95.445 179.675 ;
        RECT 95.615 179.475 95.865 179.935 ;
        RECT 94.645 179.215 95.445 179.385 ;
        RECT 96.035 179.425 96.905 179.765 ;
        RECT 92.750 177.555 93.080 178.185 ;
        RECT 93.250 177.385 93.460 178.205 ;
        RECT 93.695 178.095 93.905 178.745 ;
        RECT 94.645 178.625 94.815 179.215 ;
        RECT 96.035 179.045 96.205 179.425 ;
        RECT 97.140 179.305 97.310 179.765 ;
        RECT 97.480 179.475 97.850 179.935 ;
        RECT 98.145 179.335 98.315 179.675 ;
        RECT 98.485 179.505 98.815 179.935 ;
        RECT 99.050 179.335 99.220 179.675 ;
        RECT 94.985 178.875 96.205 179.045 ;
        RECT 96.375 178.965 96.835 179.255 ;
        RECT 97.140 179.135 97.700 179.305 ;
        RECT 98.145 179.165 99.220 179.335 ;
        RECT 99.390 179.435 100.070 179.765 ;
        RECT 100.285 179.435 100.535 179.765 ;
        RECT 100.705 179.475 100.955 179.935 ;
        RECT 97.530 178.995 97.700 179.135 ;
        RECT 96.375 178.955 97.340 178.965 ;
        RECT 96.035 178.785 96.205 178.875 ;
        RECT 96.665 178.795 97.340 178.955 ;
        RECT 94.075 178.595 94.815 178.625 ;
        RECT 94.075 178.295 94.990 178.595 ;
        RECT 94.665 178.120 94.990 178.295 ;
        RECT 93.695 177.565 93.950 178.095 ;
        RECT 94.120 177.385 94.425 177.845 ;
        RECT 94.670 177.765 94.990 178.120 ;
        RECT 95.160 178.335 95.700 178.705 ;
        RECT 96.035 178.615 96.440 178.785 ;
        RECT 95.160 177.935 95.400 178.335 ;
        RECT 95.880 178.165 96.100 178.445 ;
        RECT 95.570 177.995 96.100 178.165 ;
        RECT 95.570 177.765 95.740 177.995 ;
        RECT 96.270 177.835 96.440 178.615 ;
        RECT 96.610 178.005 96.960 178.625 ;
        RECT 97.130 178.005 97.340 178.795 ;
        RECT 97.530 178.825 99.030 178.995 ;
        RECT 97.530 178.135 97.700 178.825 ;
        RECT 99.390 178.655 99.560 179.435 ;
        RECT 100.365 179.305 100.535 179.435 ;
        RECT 97.870 178.485 99.560 178.655 ;
        RECT 99.730 178.875 100.195 179.265 ;
        RECT 100.365 179.135 100.760 179.305 ;
        RECT 97.870 178.305 98.040 178.485 ;
        RECT 94.670 177.595 95.740 177.765 ;
        RECT 95.910 177.385 96.100 177.825 ;
        RECT 96.270 177.555 97.220 177.835 ;
        RECT 97.530 177.745 97.790 178.135 ;
        RECT 98.210 178.065 99.000 178.315 ;
        RECT 97.440 177.575 97.790 177.745 ;
        RECT 98.000 177.385 98.330 177.845 ;
        RECT 99.205 177.775 99.375 178.485 ;
        RECT 99.730 178.285 99.900 178.875 ;
        RECT 99.545 178.065 99.900 178.285 ;
        RECT 100.070 178.065 100.420 178.685 ;
        RECT 100.590 177.775 100.760 179.135 ;
        RECT 101.125 178.965 101.450 179.750 ;
        RECT 100.930 177.915 101.390 178.965 ;
        RECT 99.205 177.605 100.060 177.775 ;
        RECT 100.265 177.605 100.760 177.775 ;
        RECT 100.930 177.385 101.260 177.745 ;
        RECT 101.620 177.645 101.790 179.765 ;
        RECT 101.960 179.435 102.290 179.935 ;
        RECT 102.460 179.265 102.715 179.765 ;
        RECT 101.965 179.095 102.715 179.265 ;
        RECT 101.965 178.105 102.195 179.095 ;
        RECT 102.365 178.275 102.715 178.925 ;
        RECT 102.890 178.860 103.160 179.765 ;
        RECT 103.330 179.175 103.660 179.935 ;
        RECT 103.840 179.005 104.010 179.765 ;
        RECT 101.965 177.935 102.715 178.105 ;
        RECT 101.960 177.385 102.290 177.765 ;
        RECT 102.460 177.645 102.715 177.935 ;
        RECT 102.890 178.060 103.060 178.860 ;
        RECT 103.345 178.835 104.010 179.005 ;
        RECT 104.270 178.845 105.480 179.935 ;
        RECT 105.655 179.500 111.000 179.935 ;
        RECT 103.345 178.690 103.515 178.835 ;
        RECT 103.230 178.360 103.515 178.690 ;
        RECT 103.345 178.105 103.515 178.360 ;
        RECT 103.750 178.285 104.080 178.655 ;
        RECT 104.270 178.305 104.790 178.845 ;
        RECT 104.960 178.135 105.480 178.675 ;
        RECT 107.245 178.250 107.595 179.500 ;
        RECT 111.170 178.845 112.380 179.935 ;
        RECT 102.890 177.555 103.150 178.060 ;
        RECT 103.345 177.935 104.010 178.105 ;
        RECT 103.330 177.385 103.660 177.765 ;
        RECT 103.840 177.555 104.010 177.935 ;
        RECT 104.270 177.385 105.480 178.135 ;
        RECT 109.075 177.930 109.415 178.760 ;
        RECT 111.170 178.305 111.690 178.845 ;
        RECT 111.860 178.135 112.380 178.675 ;
        RECT 105.655 177.385 111.000 177.930 ;
        RECT 111.170 177.385 112.380 178.135 ;
        RECT 18.165 177.215 112.465 177.385 ;
        RECT 18.250 176.465 19.460 177.215 ;
        RECT 18.250 175.925 18.770 176.465 ;
        RECT 20.090 176.445 21.760 177.215 ;
        RECT 21.930 176.490 22.220 177.215 ;
        RECT 23.310 176.445 26.820 177.215 ;
        RECT 26.995 176.670 32.340 177.215 ;
        RECT 32.515 176.670 37.860 177.215 ;
        RECT 18.940 175.755 19.460 176.295 ;
        RECT 18.250 174.665 19.460 175.755 ;
        RECT 20.090 175.755 20.840 176.275 ;
        RECT 21.010 175.925 21.760 176.445 ;
        RECT 20.090 174.665 21.760 175.755 ;
        RECT 21.930 174.665 22.220 175.830 ;
        RECT 23.310 175.755 25.000 176.275 ;
        RECT 25.170 175.925 26.820 176.445 ;
        RECT 23.310 174.665 26.820 175.755 ;
        RECT 28.585 175.100 28.935 176.350 ;
        RECT 30.415 175.840 30.755 176.670 ;
        RECT 34.105 175.100 34.455 176.350 ;
        RECT 35.935 175.840 36.275 176.670 ;
        RECT 38.405 176.505 38.660 177.035 ;
        RECT 38.840 176.755 39.125 177.215 ;
        RECT 38.405 175.855 38.585 176.505 ;
        RECT 39.305 176.305 39.555 176.955 ;
        RECT 38.755 175.975 39.555 176.305 ;
        RECT 38.320 175.685 38.585 175.855 ;
        RECT 38.405 175.645 38.585 175.685 ;
        RECT 26.995 174.665 32.340 175.100 ;
        RECT 32.515 174.665 37.860 175.100 ;
        RECT 38.405 174.975 38.660 175.645 ;
        RECT 38.840 174.665 39.125 175.465 ;
        RECT 39.305 175.385 39.555 175.975 ;
        RECT 39.755 176.620 40.075 176.950 ;
        RECT 40.255 176.735 40.915 177.215 ;
        RECT 41.115 176.825 41.965 176.995 ;
        RECT 39.755 175.725 39.945 176.620 ;
        RECT 40.265 176.295 40.925 176.565 ;
        RECT 40.595 176.235 40.925 176.295 ;
        RECT 40.115 176.065 40.445 176.125 ;
        RECT 41.115 176.065 41.285 176.825 ;
        RECT 42.525 176.755 42.845 177.215 ;
        RECT 43.045 176.575 43.295 177.005 ;
        RECT 43.585 176.775 43.995 177.215 ;
        RECT 44.165 176.835 45.180 177.035 ;
        RECT 41.455 176.405 42.705 176.575 ;
        RECT 41.455 176.285 41.785 176.405 ;
        RECT 40.115 175.895 42.015 176.065 ;
        RECT 39.755 175.555 41.675 175.725 ;
        RECT 39.755 175.535 40.075 175.555 ;
        RECT 39.305 174.875 39.635 175.385 ;
        RECT 39.905 174.925 40.075 175.535 ;
        RECT 41.845 175.385 42.015 175.895 ;
        RECT 42.185 175.825 42.365 176.235 ;
        RECT 42.535 175.645 42.705 176.405 ;
        RECT 40.245 174.665 40.575 175.355 ;
        RECT 40.805 175.215 42.015 175.385 ;
        RECT 42.185 175.335 42.705 175.645 ;
        RECT 42.875 176.235 43.295 176.575 ;
        RECT 43.585 176.235 43.995 176.565 ;
        RECT 42.875 175.465 43.065 176.235 ;
        RECT 44.165 176.105 44.335 176.835 ;
        RECT 45.480 176.665 45.650 176.995 ;
        RECT 45.820 176.835 46.150 177.215 ;
        RECT 44.505 176.285 44.855 176.655 ;
        RECT 44.165 176.065 44.585 176.105 ;
        RECT 43.235 175.895 44.585 176.065 ;
        RECT 43.235 175.735 43.485 175.895 ;
        RECT 43.995 175.465 44.245 175.725 ;
        RECT 42.875 175.215 44.245 175.465 ;
        RECT 40.805 174.925 41.045 175.215 ;
        RECT 41.845 175.135 42.015 175.215 ;
        RECT 41.245 174.665 41.665 175.045 ;
        RECT 41.845 174.885 42.475 175.135 ;
        RECT 42.945 174.665 43.275 175.045 ;
        RECT 43.445 174.925 43.615 175.215 ;
        RECT 44.415 175.050 44.585 175.895 ;
        RECT 45.035 175.725 45.255 176.595 ;
        RECT 45.480 176.475 46.175 176.665 ;
        RECT 44.755 175.345 45.255 175.725 ;
        RECT 45.425 175.675 45.835 176.295 ;
        RECT 46.005 175.505 46.175 176.475 ;
        RECT 45.480 175.335 46.175 175.505 ;
        RECT 43.795 174.665 44.175 175.045 ;
        RECT 44.415 174.880 45.245 175.050 ;
        RECT 45.480 174.835 45.650 175.335 ;
        RECT 45.820 174.665 46.150 175.165 ;
        RECT 46.365 174.835 46.590 176.955 ;
        RECT 46.760 176.835 47.090 177.215 ;
        RECT 47.260 176.665 47.430 176.955 ;
        RECT 46.765 176.495 47.430 176.665 ;
        RECT 46.765 175.505 46.995 176.495 ;
        RECT 47.690 176.490 47.980 177.215 ;
        RECT 48.210 176.395 48.420 177.215 ;
        RECT 48.590 176.415 48.920 177.045 ;
        RECT 47.165 175.675 47.515 176.325 ;
        RECT 46.765 175.335 47.430 175.505 ;
        RECT 46.760 174.665 47.090 175.165 ;
        RECT 47.260 174.835 47.430 175.335 ;
        RECT 47.690 174.665 47.980 175.830 ;
        RECT 48.590 175.815 48.840 176.415 ;
        RECT 49.090 176.395 49.320 177.215 ;
        RECT 50.540 176.665 50.710 177.045 ;
        RECT 50.890 176.835 51.220 177.215 ;
        RECT 50.540 176.495 51.205 176.665 ;
        RECT 51.400 176.540 51.660 177.045 ;
        RECT 49.010 175.975 49.340 176.225 ;
        RECT 50.470 175.945 50.800 176.315 ;
        RECT 51.035 176.240 51.205 176.495 ;
        RECT 51.035 175.910 51.320 176.240 ;
        RECT 48.210 174.665 48.420 175.805 ;
        RECT 48.590 174.835 48.920 175.815 ;
        RECT 49.090 174.665 49.320 175.805 ;
        RECT 51.035 175.765 51.205 175.910 ;
        RECT 50.540 175.595 51.205 175.765 ;
        RECT 51.490 175.740 51.660 176.540 ;
        RECT 51.890 176.395 52.100 177.215 ;
        RECT 52.270 176.415 52.600 177.045 ;
        RECT 52.270 175.815 52.520 176.415 ;
        RECT 52.770 176.395 53.000 177.215 ;
        RECT 53.210 176.540 53.470 177.045 ;
        RECT 53.650 176.835 53.980 177.215 ;
        RECT 54.160 176.665 54.330 177.045 ;
        RECT 55.360 176.745 55.530 177.215 ;
        RECT 52.690 175.975 53.020 176.225 ;
        RECT 50.540 174.835 50.710 175.595 ;
        RECT 50.890 174.665 51.220 175.425 ;
        RECT 51.390 174.835 51.660 175.740 ;
        RECT 51.890 174.665 52.100 175.805 ;
        RECT 52.270 174.835 52.600 175.815 ;
        RECT 52.770 174.665 53.000 175.805 ;
        RECT 53.210 175.740 53.380 176.540 ;
        RECT 53.665 176.495 54.330 176.665 ;
        RECT 55.700 176.565 56.030 177.045 ;
        RECT 56.200 176.745 56.370 177.215 ;
        RECT 56.540 176.565 56.870 177.045 ;
        RECT 53.665 176.240 53.835 176.495 ;
        RECT 55.105 176.395 56.870 176.565 ;
        RECT 57.040 176.405 57.210 177.215 ;
        RECT 57.410 176.835 58.480 177.005 ;
        RECT 57.410 176.480 57.730 176.835 ;
        RECT 53.550 175.910 53.835 176.240 ;
        RECT 54.070 175.945 54.400 176.315 ;
        RECT 53.665 175.765 53.835 175.910 ;
        RECT 55.105 175.845 55.515 176.395 ;
        RECT 57.405 176.225 57.730 176.480 ;
        RECT 55.700 176.015 57.730 176.225 ;
        RECT 57.385 176.005 57.730 176.015 ;
        RECT 57.900 176.265 58.140 176.665 ;
        RECT 58.310 176.605 58.480 176.835 ;
        RECT 58.650 176.775 58.840 177.215 ;
        RECT 59.010 176.765 59.960 177.045 ;
        RECT 60.180 176.855 60.530 177.025 ;
        RECT 58.310 176.435 58.840 176.605 ;
        RECT 53.210 174.835 53.480 175.740 ;
        RECT 53.665 175.595 54.330 175.765 ;
        RECT 55.105 175.675 56.830 175.845 ;
        RECT 53.650 174.665 53.980 175.425 ;
        RECT 54.160 174.835 54.330 175.595 ;
        RECT 55.360 174.665 55.530 175.505 ;
        RECT 55.740 174.835 55.990 175.675 ;
        RECT 56.200 174.665 56.370 175.505 ;
        RECT 56.540 174.835 56.830 175.675 ;
        RECT 57.040 174.665 57.210 175.725 ;
        RECT 57.385 175.385 57.555 176.005 ;
        RECT 57.900 175.895 58.440 176.265 ;
        RECT 58.620 176.155 58.840 176.435 ;
        RECT 59.010 175.985 59.180 176.765 ;
        RECT 58.775 175.815 59.180 175.985 ;
        RECT 59.350 175.975 59.700 176.595 ;
        RECT 58.775 175.725 58.945 175.815 ;
        RECT 59.870 175.805 60.080 176.595 ;
        RECT 57.725 175.555 58.945 175.725 ;
        RECT 59.405 175.645 60.080 175.805 ;
        RECT 57.385 175.215 58.185 175.385 ;
        RECT 57.505 174.665 57.835 175.045 ;
        RECT 58.015 174.925 58.185 175.215 ;
        RECT 58.775 175.175 58.945 175.555 ;
        RECT 59.115 175.635 60.080 175.645 ;
        RECT 60.270 176.465 60.530 176.855 ;
        RECT 60.740 176.755 61.070 177.215 ;
        RECT 61.945 176.825 62.800 176.995 ;
        RECT 63.005 176.825 63.500 176.995 ;
        RECT 63.670 176.855 64.000 177.215 ;
        RECT 60.270 175.775 60.440 176.465 ;
        RECT 60.610 176.115 60.780 176.295 ;
        RECT 60.950 176.285 61.740 176.535 ;
        RECT 61.945 176.115 62.115 176.825 ;
        RECT 62.285 176.315 62.640 176.535 ;
        RECT 60.610 175.945 62.300 176.115 ;
        RECT 59.115 175.345 59.575 175.635 ;
        RECT 60.270 175.605 61.770 175.775 ;
        RECT 60.270 175.465 60.440 175.605 ;
        RECT 59.880 175.295 60.440 175.465 ;
        RECT 58.355 174.665 58.605 175.125 ;
        RECT 58.775 174.835 59.645 175.175 ;
        RECT 59.880 174.835 60.050 175.295 ;
        RECT 60.885 175.265 61.960 175.435 ;
        RECT 60.220 174.665 60.590 175.125 ;
        RECT 60.885 174.925 61.055 175.265 ;
        RECT 61.225 174.665 61.555 175.095 ;
        RECT 61.790 174.925 61.960 175.265 ;
        RECT 62.130 175.165 62.300 175.945 ;
        RECT 62.470 175.725 62.640 176.315 ;
        RECT 62.810 175.915 63.160 176.535 ;
        RECT 62.470 175.335 62.935 175.725 ;
        RECT 63.330 175.465 63.500 176.825 ;
        RECT 63.670 175.635 64.130 176.685 ;
        RECT 63.105 175.295 63.500 175.465 ;
        RECT 63.105 175.165 63.275 175.295 ;
        RECT 62.130 174.835 62.810 175.165 ;
        RECT 63.025 174.835 63.275 175.165 ;
        RECT 63.445 174.665 63.695 175.125 ;
        RECT 63.865 174.850 64.190 175.635 ;
        RECT 64.360 174.835 64.530 176.955 ;
        RECT 64.700 176.835 65.030 177.215 ;
        RECT 65.200 176.665 65.455 176.955 ;
        RECT 64.705 176.495 65.455 176.665 ;
        RECT 64.705 175.505 64.935 176.495 ;
        RECT 65.630 176.395 65.890 177.215 ;
        RECT 66.060 176.395 66.390 176.815 ;
        RECT 66.570 176.645 66.830 177.045 ;
        RECT 67.000 176.815 67.330 177.215 ;
        RECT 67.500 176.645 67.670 176.995 ;
        RECT 67.840 176.815 68.215 177.215 ;
        RECT 66.570 176.475 68.235 176.645 ;
        RECT 68.405 176.540 68.680 176.885 ;
        RECT 65.105 175.675 65.455 176.325 ;
        RECT 66.140 176.305 66.390 176.395 ;
        RECT 68.065 176.305 68.235 176.475 ;
        RECT 65.635 175.975 65.970 176.225 ;
        RECT 66.140 175.975 66.855 176.305 ;
        RECT 67.070 175.975 67.895 176.305 ;
        RECT 68.065 175.975 68.340 176.305 ;
        RECT 64.705 175.335 65.455 175.505 ;
        RECT 64.700 174.665 65.030 175.165 ;
        RECT 65.200 174.835 65.455 175.335 ;
        RECT 65.630 174.665 65.890 175.805 ;
        RECT 66.140 175.415 66.310 175.975 ;
        RECT 66.570 175.515 66.900 175.805 ;
        RECT 67.070 175.685 67.315 175.975 ;
        RECT 68.065 175.805 68.235 175.975 ;
        RECT 68.510 175.805 68.680 176.540 ;
        RECT 69.585 176.405 69.830 177.010 ;
        RECT 70.050 176.680 70.560 177.215 ;
        RECT 67.575 175.635 68.235 175.805 ;
        RECT 67.575 175.515 67.745 175.635 ;
        RECT 66.570 175.345 67.745 175.515 ;
        RECT 66.130 174.845 67.745 175.175 ;
        RECT 67.915 174.665 68.195 175.465 ;
        RECT 68.405 174.835 68.680 175.805 ;
        RECT 69.310 176.235 70.540 176.405 ;
        RECT 69.310 175.425 69.650 176.235 ;
        RECT 69.820 175.670 70.570 175.860 ;
        RECT 69.310 175.015 69.825 175.425 ;
        RECT 70.060 174.665 70.230 175.425 ;
        RECT 70.400 175.005 70.570 175.670 ;
        RECT 70.740 175.685 70.930 177.045 ;
        RECT 71.100 176.195 71.375 177.045 ;
        RECT 71.565 176.680 72.095 177.045 ;
        RECT 72.520 176.815 72.850 177.215 ;
        RECT 71.920 176.645 72.095 176.680 ;
        RECT 71.100 176.025 71.380 176.195 ;
        RECT 71.100 175.885 71.375 176.025 ;
        RECT 71.580 175.685 71.750 176.485 ;
        RECT 70.740 175.515 71.750 175.685 ;
        RECT 71.920 176.475 72.850 176.645 ;
        RECT 73.020 176.475 73.275 177.045 ;
        RECT 73.450 176.490 73.740 177.215 ;
        RECT 74.285 176.505 74.540 177.035 ;
        RECT 74.720 176.755 75.005 177.215 ;
        RECT 71.920 175.345 72.090 176.475 ;
        RECT 72.680 176.305 72.850 176.475 ;
        RECT 70.965 175.175 72.090 175.345 ;
        RECT 72.260 175.975 72.455 176.305 ;
        RECT 72.680 175.975 72.935 176.305 ;
        RECT 72.260 175.005 72.430 175.975 ;
        RECT 73.105 175.805 73.275 176.475 ;
        RECT 70.400 174.835 72.430 175.005 ;
        RECT 72.600 174.665 72.770 175.805 ;
        RECT 72.940 174.835 73.275 175.805 ;
        RECT 73.450 174.665 73.740 175.830 ;
        RECT 74.285 175.645 74.465 176.505 ;
        RECT 75.185 176.305 75.435 176.955 ;
        RECT 74.635 175.975 75.435 176.305 ;
        RECT 74.285 175.175 74.540 175.645 ;
        RECT 74.200 175.005 74.540 175.175 ;
        RECT 74.285 174.975 74.540 175.005 ;
        RECT 74.720 174.665 75.005 175.465 ;
        RECT 75.185 175.385 75.435 175.975 ;
        RECT 75.635 176.620 75.955 176.950 ;
        RECT 76.135 176.735 76.795 177.215 ;
        RECT 76.995 176.825 77.845 176.995 ;
        RECT 75.635 175.725 75.825 176.620 ;
        RECT 76.145 176.295 76.805 176.565 ;
        RECT 76.475 176.235 76.805 176.295 ;
        RECT 75.995 176.065 76.325 176.125 ;
        RECT 76.995 176.065 77.165 176.825 ;
        RECT 78.405 176.755 78.725 177.215 ;
        RECT 78.925 176.575 79.175 177.005 ;
        RECT 79.465 176.775 79.875 177.215 ;
        RECT 80.045 176.835 81.060 177.035 ;
        RECT 77.335 176.405 78.585 176.575 ;
        RECT 77.335 176.285 77.665 176.405 ;
        RECT 75.995 175.895 77.895 176.065 ;
        RECT 75.635 175.555 77.555 175.725 ;
        RECT 75.635 175.535 75.955 175.555 ;
        RECT 75.185 174.875 75.515 175.385 ;
        RECT 75.785 174.925 75.955 175.535 ;
        RECT 77.725 175.385 77.895 175.895 ;
        RECT 78.065 175.825 78.245 176.235 ;
        RECT 78.415 175.645 78.585 176.405 ;
        RECT 76.125 174.665 76.455 175.355 ;
        RECT 76.685 175.215 77.895 175.385 ;
        RECT 78.065 175.335 78.585 175.645 ;
        RECT 78.755 176.235 79.175 176.575 ;
        RECT 79.465 176.235 79.875 176.565 ;
        RECT 78.755 175.465 78.945 176.235 ;
        RECT 80.045 176.105 80.215 176.835 ;
        RECT 81.360 176.665 81.530 176.995 ;
        RECT 81.700 176.835 82.030 177.215 ;
        RECT 80.385 176.285 80.735 176.655 ;
        RECT 80.045 176.065 80.465 176.105 ;
        RECT 79.115 175.895 80.465 176.065 ;
        RECT 79.115 175.735 79.365 175.895 ;
        RECT 79.875 175.465 80.125 175.725 ;
        RECT 78.755 175.215 80.125 175.465 ;
        RECT 76.685 174.925 76.925 175.215 ;
        RECT 77.725 175.135 77.895 175.215 ;
        RECT 77.125 174.665 77.545 175.045 ;
        RECT 77.725 174.885 78.355 175.135 ;
        RECT 78.825 174.665 79.155 175.045 ;
        RECT 79.325 174.925 79.495 175.215 ;
        RECT 80.295 175.050 80.465 175.895 ;
        RECT 80.915 175.725 81.135 176.595 ;
        RECT 81.360 176.475 82.055 176.665 ;
        RECT 80.635 175.345 81.135 175.725 ;
        RECT 81.305 175.675 81.715 176.295 ;
        RECT 81.885 175.505 82.055 176.475 ;
        RECT 81.360 175.335 82.055 175.505 ;
        RECT 79.675 174.665 80.055 175.045 ;
        RECT 80.295 174.880 81.125 175.050 ;
        RECT 81.360 174.835 81.530 175.335 ;
        RECT 81.700 174.665 82.030 175.165 ;
        RECT 82.245 174.835 82.470 176.955 ;
        RECT 82.640 176.835 82.970 177.215 ;
        RECT 83.140 176.665 83.310 176.955 ;
        RECT 82.645 176.495 83.310 176.665 ;
        RECT 82.645 175.505 82.875 176.495 ;
        RECT 84.030 176.445 85.700 177.215 ;
        RECT 83.045 175.675 83.395 176.325 ;
        RECT 84.030 175.755 84.780 176.275 ;
        RECT 84.950 175.925 85.700 176.445 ;
        RECT 85.910 176.395 86.140 177.215 ;
        RECT 86.310 176.415 86.640 177.045 ;
        RECT 85.890 175.975 86.220 176.225 ;
        RECT 86.390 175.815 86.640 176.415 ;
        RECT 86.810 176.395 87.020 177.215 ;
        RECT 87.800 176.665 87.970 177.045 ;
        RECT 88.150 176.835 88.480 177.215 ;
        RECT 87.800 176.495 88.465 176.665 ;
        RECT 88.660 176.540 88.920 177.045 ;
        RECT 87.730 175.945 88.060 176.315 ;
        RECT 88.295 176.240 88.465 176.495 ;
        RECT 82.645 175.335 83.310 175.505 ;
        RECT 82.640 174.665 82.970 175.165 ;
        RECT 83.140 174.835 83.310 175.335 ;
        RECT 84.030 174.665 85.700 175.755 ;
        RECT 85.910 174.665 86.140 175.805 ;
        RECT 86.310 174.835 86.640 175.815 ;
        RECT 88.295 175.910 88.580 176.240 ;
        RECT 86.810 174.665 87.020 175.805 ;
        RECT 88.295 175.765 88.465 175.910 ;
        RECT 87.800 175.595 88.465 175.765 ;
        RECT 88.750 175.740 88.920 176.540 ;
        RECT 87.800 174.835 87.970 175.595 ;
        RECT 88.150 174.665 88.480 175.425 ;
        RECT 88.650 174.835 88.920 175.740 ;
        RECT 89.095 176.505 89.350 177.035 ;
        RECT 89.520 176.755 89.825 177.215 ;
        RECT 90.070 176.835 91.140 177.005 ;
        RECT 89.095 175.855 89.305 176.505 ;
        RECT 90.070 176.480 90.390 176.835 ;
        RECT 90.065 176.305 90.390 176.480 ;
        RECT 89.475 176.005 90.390 176.305 ;
        RECT 90.560 176.265 90.800 176.665 ;
        RECT 90.970 176.605 91.140 176.835 ;
        RECT 91.310 176.775 91.500 177.215 ;
        RECT 91.670 176.765 92.620 177.045 ;
        RECT 92.840 176.855 93.190 177.025 ;
        RECT 90.970 176.435 91.500 176.605 ;
        RECT 89.475 175.975 90.215 176.005 ;
        RECT 89.095 174.975 89.350 175.855 ;
        RECT 89.520 174.665 89.825 175.805 ;
        RECT 90.045 175.385 90.215 175.975 ;
        RECT 90.560 175.895 91.100 176.265 ;
        RECT 91.280 176.155 91.500 176.435 ;
        RECT 91.670 175.985 91.840 176.765 ;
        RECT 91.435 175.815 91.840 175.985 ;
        RECT 92.010 175.975 92.360 176.595 ;
        RECT 91.435 175.725 91.605 175.815 ;
        RECT 92.530 175.805 92.740 176.595 ;
        RECT 90.385 175.555 91.605 175.725 ;
        RECT 92.065 175.645 92.740 175.805 ;
        RECT 90.045 175.215 90.845 175.385 ;
        RECT 90.165 174.665 90.495 175.045 ;
        RECT 90.675 174.925 90.845 175.215 ;
        RECT 91.435 175.175 91.605 175.555 ;
        RECT 91.775 175.635 92.740 175.645 ;
        RECT 92.930 176.465 93.190 176.855 ;
        RECT 93.400 176.755 93.730 177.215 ;
        RECT 94.605 176.825 95.460 176.995 ;
        RECT 95.665 176.825 96.160 176.995 ;
        RECT 96.330 176.855 96.660 177.215 ;
        RECT 92.930 175.775 93.100 176.465 ;
        RECT 93.270 176.115 93.440 176.295 ;
        RECT 93.610 176.285 94.400 176.535 ;
        RECT 94.605 176.115 94.775 176.825 ;
        RECT 94.945 176.315 95.300 176.535 ;
        RECT 93.270 175.945 94.960 176.115 ;
        RECT 91.775 175.345 92.235 175.635 ;
        RECT 92.930 175.605 94.430 175.775 ;
        RECT 92.930 175.465 93.100 175.605 ;
        RECT 92.540 175.295 93.100 175.465 ;
        RECT 91.015 174.665 91.265 175.125 ;
        RECT 91.435 174.835 92.305 175.175 ;
        RECT 92.540 174.835 92.710 175.295 ;
        RECT 93.545 175.265 94.620 175.435 ;
        RECT 92.880 174.665 93.250 175.125 ;
        RECT 93.545 174.925 93.715 175.265 ;
        RECT 93.885 174.665 94.215 175.095 ;
        RECT 94.450 174.925 94.620 175.265 ;
        RECT 94.790 175.165 94.960 175.945 ;
        RECT 95.130 175.725 95.300 176.315 ;
        RECT 95.470 175.915 95.820 176.535 ;
        RECT 95.130 175.335 95.595 175.725 ;
        RECT 95.990 175.465 96.160 176.825 ;
        RECT 96.330 175.635 96.790 176.685 ;
        RECT 95.765 175.295 96.160 175.465 ;
        RECT 95.765 175.165 95.935 175.295 ;
        RECT 94.790 174.835 95.470 175.165 ;
        RECT 95.685 174.835 95.935 175.165 ;
        RECT 96.105 174.665 96.355 175.125 ;
        RECT 96.525 174.850 96.850 175.635 ;
        RECT 97.020 174.835 97.190 176.955 ;
        RECT 97.360 176.835 97.690 177.215 ;
        RECT 97.860 176.665 98.115 176.955 ;
        RECT 97.365 176.495 98.115 176.665 ;
        RECT 97.365 175.505 97.595 176.495 ;
        RECT 99.210 176.490 99.500 177.215 ;
        RECT 100.130 176.445 101.800 177.215 ;
        RECT 97.765 175.675 98.115 176.325 ;
        RECT 97.365 175.335 98.115 175.505 ;
        RECT 97.360 174.665 97.690 175.165 ;
        RECT 97.860 174.835 98.115 175.335 ;
        RECT 99.210 174.665 99.500 175.830 ;
        RECT 100.130 175.755 100.880 176.275 ;
        RECT 101.050 175.925 101.800 176.445 ;
        RECT 102.010 176.395 102.240 177.215 ;
        RECT 102.410 176.415 102.740 177.045 ;
        RECT 101.990 175.975 102.320 176.225 ;
        RECT 102.490 175.815 102.740 176.415 ;
        RECT 102.910 176.395 103.120 177.215 ;
        RECT 103.410 176.395 103.620 177.215 ;
        RECT 103.790 176.415 104.120 177.045 ;
        RECT 100.130 174.665 101.800 175.755 ;
        RECT 102.010 174.665 102.240 175.805 ;
        RECT 102.410 174.835 102.740 175.815 ;
        RECT 103.790 175.815 104.040 176.415 ;
        RECT 104.290 176.395 104.520 177.215 ;
        RECT 105.655 176.670 111.000 177.215 ;
        RECT 104.210 175.975 104.540 176.225 ;
        RECT 102.910 174.665 103.120 175.805 ;
        RECT 103.410 174.665 103.620 175.805 ;
        RECT 103.790 174.835 104.120 175.815 ;
        RECT 104.290 174.665 104.520 175.805 ;
        RECT 107.245 175.100 107.595 176.350 ;
        RECT 109.075 175.840 109.415 176.670 ;
        RECT 111.170 176.465 112.380 177.215 ;
        RECT 111.170 175.755 111.690 176.295 ;
        RECT 111.860 175.925 112.380 176.465 ;
        RECT 105.655 174.665 111.000 175.100 ;
        RECT 111.170 174.665 112.380 175.755 ;
        RECT 18.165 174.495 112.465 174.665 ;
        RECT 18.250 173.405 19.460 174.495 ;
        RECT 18.250 172.695 18.770 173.235 ;
        RECT 18.940 172.865 19.460 173.405 ;
        RECT 20.090 173.405 23.600 174.495 ;
        RECT 23.775 174.060 29.120 174.495 ;
        RECT 29.295 174.060 34.640 174.495 ;
        RECT 20.090 172.885 21.780 173.405 ;
        RECT 21.950 172.715 23.600 173.235 ;
        RECT 25.365 172.810 25.715 174.060 ;
        RECT 18.250 171.945 19.460 172.695 ;
        RECT 20.090 171.945 23.600 172.715 ;
        RECT 27.195 172.490 27.535 173.320 ;
        RECT 30.885 172.810 31.235 174.060 ;
        RECT 34.810 173.330 35.100 174.495 ;
        RECT 35.730 173.405 38.320 174.495 ;
        RECT 32.715 172.490 33.055 173.320 ;
        RECT 35.730 172.885 36.940 173.405 ;
        RECT 38.530 173.355 38.760 174.495 ;
        RECT 38.930 173.345 39.260 174.325 ;
        RECT 39.430 173.355 39.640 174.495 ;
        RECT 39.870 173.735 40.385 174.145 ;
        RECT 40.620 173.735 40.790 174.495 ;
        RECT 40.960 174.155 42.990 174.325 ;
        RECT 37.110 172.715 38.320 173.235 ;
        RECT 38.510 172.935 38.840 173.185 ;
        RECT 23.775 171.945 29.120 172.490 ;
        RECT 29.295 171.945 34.640 172.490 ;
        RECT 34.810 171.945 35.100 172.670 ;
        RECT 35.730 171.945 38.320 172.715 ;
        RECT 38.530 171.945 38.760 172.765 ;
        RECT 39.010 172.745 39.260 173.345 ;
        RECT 39.870 172.925 40.210 173.735 ;
        RECT 40.960 173.490 41.130 174.155 ;
        RECT 41.525 173.815 42.650 173.985 ;
        RECT 40.380 173.300 41.130 173.490 ;
        RECT 41.300 173.475 42.310 173.645 ;
        RECT 38.930 172.115 39.260 172.745 ;
        RECT 39.430 171.945 39.640 172.765 ;
        RECT 39.870 172.755 41.100 172.925 ;
        RECT 40.145 172.150 40.390 172.755 ;
        RECT 40.610 171.945 41.120 172.480 ;
        RECT 41.300 172.115 41.490 173.475 ;
        RECT 41.660 172.795 41.935 173.275 ;
        RECT 41.660 172.625 41.940 172.795 ;
        RECT 42.140 172.675 42.310 173.475 ;
        RECT 42.480 172.685 42.650 173.815 ;
        RECT 42.820 173.185 42.990 174.155 ;
        RECT 43.160 173.355 43.330 174.495 ;
        RECT 43.500 173.355 43.835 174.325 ;
        RECT 42.820 172.855 43.015 173.185 ;
        RECT 43.240 172.855 43.495 173.185 ;
        RECT 43.240 172.685 43.410 172.855 ;
        RECT 43.665 172.685 43.835 173.355 ;
        RECT 44.010 173.735 44.525 174.145 ;
        RECT 44.760 173.735 44.930 174.495 ;
        RECT 45.100 174.155 47.130 174.325 ;
        RECT 44.010 172.925 44.350 173.735 ;
        RECT 45.100 173.490 45.270 174.155 ;
        RECT 45.665 173.815 46.790 173.985 ;
        RECT 44.520 173.300 45.270 173.490 ;
        RECT 45.440 173.475 46.450 173.645 ;
        RECT 44.010 172.755 45.240 172.925 ;
        RECT 41.660 172.115 41.935 172.625 ;
        RECT 42.480 172.515 43.410 172.685 ;
        RECT 42.480 172.480 42.655 172.515 ;
        RECT 42.125 172.115 42.655 172.480 ;
        RECT 43.080 171.945 43.410 172.345 ;
        RECT 43.580 172.115 43.835 172.685 ;
        RECT 44.285 172.150 44.530 172.755 ;
        RECT 44.750 171.945 45.260 172.480 ;
        RECT 45.440 172.115 45.630 173.475 ;
        RECT 45.800 172.455 46.075 173.275 ;
        RECT 46.280 172.675 46.450 173.475 ;
        RECT 46.620 172.685 46.790 173.815 ;
        RECT 46.960 173.185 47.130 174.155 ;
        RECT 47.300 173.355 47.470 174.495 ;
        RECT 47.640 173.355 47.975 174.325 ;
        RECT 46.960 172.855 47.155 173.185 ;
        RECT 47.380 172.855 47.635 173.185 ;
        RECT 47.380 172.685 47.550 172.855 ;
        RECT 47.805 172.685 47.975 173.355 ;
        RECT 46.620 172.515 47.550 172.685 ;
        RECT 46.620 172.480 46.795 172.515 ;
        RECT 45.800 172.285 46.080 172.455 ;
        RECT 45.800 172.115 46.075 172.285 ;
        RECT 46.265 172.115 46.795 172.480 ;
        RECT 47.220 171.945 47.550 172.345 ;
        RECT 47.720 172.115 47.975 172.685 ;
        RECT 48.525 173.515 48.780 174.185 ;
        RECT 48.960 173.695 49.245 174.495 ;
        RECT 49.425 173.775 49.755 174.285 ;
        RECT 48.525 172.655 48.705 173.515 ;
        RECT 49.425 173.185 49.675 173.775 ;
        RECT 50.025 173.625 50.195 174.235 ;
        RECT 50.365 173.805 50.695 174.495 ;
        RECT 50.925 173.945 51.165 174.235 ;
        RECT 51.365 174.115 51.785 174.495 ;
        RECT 51.965 174.025 52.595 174.275 ;
        RECT 53.065 174.115 53.395 174.495 ;
        RECT 51.965 173.945 52.135 174.025 ;
        RECT 53.565 173.945 53.735 174.235 ;
        RECT 53.915 174.115 54.295 174.495 ;
        RECT 54.535 174.110 55.365 174.280 ;
        RECT 50.925 173.775 52.135 173.945 ;
        RECT 48.875 172.855 49.675 173.185 ;
        RECT 48.525 172.455 48.780 172.655 ;
        RECT 48.440 172.285 48.780 172.455 ;
        RECT 48.525 172.125 48.780 172.285 ;
        RECT 48.960 171.945 49.245 172.405 ;
        RECT 49.425 172.205 49.675 172.855 ;
        RECT 49.875 173.605 50.195 173.625 ;
        RECT 49.875 173.435 51.795 173.605 ;
        RECT 49.875 172.540 50.065 173.435 ;
        RECT 51.965 173.265 52.135 173.775 ;
        RECT 52.305 173.515 52.825 173.825 ;
        RECT 50.235 173.095 52.135 173.265 ;
        RECT 50.235 173.035 50.565 173.095 ;
        RECT 50.715 172.865 51.045 172.925 ;
        RECT 50.385 172.595 51.045 172.865 ;
        RECT 49.875 172.210 50.195 172.540 ;
        RECT 50.375 171.945 51.035 172.425 ;
        RECT 51.235 172.335 51.405 173.095 ;
        RECT 52.305 172.925 52.485 173.335 ;
        RECT 51.575 172.755 51.905 172.875 ;
        RECT 52.655 172.755 52.825 173.515 ;
        RECT 51.575 172.585 52.825 172.755 ;
        RECT 52.995 173.695 54.365 173.945 ;
        RECT 52.995 172.925 53.185 173.695 ;
        RECT 54.115 173.435 54.365 173.695 ;
        RECT 53.355 173.265 53.605 173.425 ;
        RECT 54.535 173.265 54.705 174.110 ;
        RECT 55.600 173.825 55.770 174.325 ;
        RECT 55.940 173.995 56.270 174.495 ;
        RECT 54.875 173.435 55.375 173.815 ;
        RECT 55.600 173.655 56.295 173.825 ;
        RECT 53.355 173.095 54.705 173.265 ;
        RECT 54.285 173.055 54.705 173.095 ;
        RECT 52.995 172.585 53.415 172.925 ;
        RECT 53.705 172.595 54.115 172.925 ;
        RECT 51.235 172.165 52.085 172.335 ;
        RECT 52.645 171.945 52.965 172.405 ;
        RECT 53.165 172.155 53.415 172.585 ;
        RECT 53.705 171.945 54.115 172.385 ;
        RECT 54.285 172.325 54.455 173.055 ;
        RECT 54.625 172.505 54.975 172.875 ;
        RECT 55.155 172.565 55.375 173.435 ;
        RECT 55.545 172.865 55.955 173.485 ;
        RECT 56.125 172.685 56.295 173.655 ;
        RECT 55.600 172.495 56.295 172.685 ;
        RECT 54.285 172.125 55.300 172.325 ;
        RECT 55.600 172.165 55.770 172.495 ;
        RECT 55.940 171.945 56.270 172.325 ;
        RECT 56.485 172.205 56.710 174.325 ;
        RECT 56.880 173.995 57.210 174.495 ;
        RECT 57.380 173.825 57.550 174.325 ;
        RECT 56.885 173.655 57.550 173.825 ;
        RECT 56.885 172.665 57.115 173.655 ;
        RECT 57.285 172.835 57.635 173.485 ;
        RECT 57.810 173.405 59.020 174.495 ;
        RECT 57.810 172.865 58.330 173.405 ;
        RECT 59.250 173.355 59.460 174.495 ;
        RECT 59.630 173.345 59.960 174.325 ;
        RECT 60.130 173.355 60.360 174.495 ;
        RECT 58.500 172.695 59.020 173.235 ;
        RECT 56.885 172.495 57.550 172.665 ;
        RECT 56.880 171.945 57.210 172.325 ;
        RECT 57.380 172.205 57.550 172.495 ;
        RECT 57.810 171.945 59.020 172.695 ;
        RECT 59.250 171.945 59.460 172.765 ;
        RECT 59.630 172.745 59.880 173.345 ;
        RECT 60.570 173.330 60.860 174.495 ;
        RECT 62.010 173.355 62.220 174.495 ;
        RECT 62.390 173.345 62.720 174.325 ;
        RECT 62.890 173.355 63.120 174.495 ;
        RECT 64.250 173.355 64.510 174.495 ;
        RECT 64.750 173.985 66.365 174.315 ;
        RECT 60.050 172.935 60.380 173.185 ;
        RECT 59.630 172.115 59.960 172.745 ;
        RECT 60.130 171.945 60.360 172.765 ;
        RECT 60.570 171.945 60.860 172.670 ;
        RECT 62.010 171.945 62.220 172.765 ;
        RECT 62.390 172.745 62.640 173.345 ;
        RECT 64.760 173.185 64.930 173.745 ;
        RECT 65.190 173.645 66.365 173.815 ;
        RECT 66.535 173.695 66.815 174.495 ;
        RECT 65.190 173.355 65.520 173.645 ;
        RECT 66.195 173.525 66.365 173.645 ;
        RECT 65.690 173.185 65.935 173.475 ;
        RECT 66.195 173.355 66.855 173.525 ;
        RECT 67.025 173.355 67.300 174.325 ;
        RECT 67.490 173.985 67.790 174.495 ;
        RECT 67.960 173.985 68.340 174.155 ;
        RECT 68.920 173.985 69.550 174.495 ;
        RECT 67.960 173.815 68.130 173.985 ;
        RECT 69.720 173.815 70.050 174.325 ;
        RECT 70.220 173.985 70.520 174.495 ;
        RECT 66.685 173.185 66.855 173.355 ;
        RECT 62.810 172.935 63.140 173.185 ;
        RECT 64.255 172.935 64.590 173.185 ;
        RECT 64.760 172.855 65.475 173.185 ;
        RECT 65.690 172.855 66.515 173.185 ;
        RECT 66.685 172.855 66.960 173.185 ;
        RECT 64.760 172.765 65.010 172.855 ;
        RECT 62.390 172.115 62.720 172.745 ;
        RECT 62.890 171.945 63.120 172.765 ;
        RECT 64.250 171.945 64.510 172.765 ;
        RECT 64.680 172.345 65.010 172.765 ;
        RECT 66.685 172.685 66.855 172.855 ;
        RECT 65.190 172.515 66.855 172.685 ;
        RECT 67.130 172.620 67.300 173.355 ;
        RECT 65.190 172.115 65.450 172.515 ;
        RECT 65.620 171.945 65.950 172.345 ;
        RECT 66.120 172.165 66.290 172.515 ;
        RECT 66.460 171.945 66.835 172.345 ;
        RECT 67.025 172.275 67.300 172.620 ;
        RECT 67.470 173.615 68.130 173.815 ;
        RECT 68.300 173.645 70.520 173.815 ;
        RECT 67.470 172.685 67.640 173.615 ;
        RECT 68.300 173.445 68.470 173.645 ;
        RECT 67.810 173.275 68.470 173.445 ;
        RECT 68.640 173.305 70.180 173.475 ;
        RECT 67.810 172.855 67.980 173.275 ;
        RECT 68.640 173.105 68.810 173.305 ;
        RECT 68.210 172.935 68.810 173.105 ;
        RECT 68.980 172.935 69.675 173.135 ;
        RECT 69.935 172.855 70.180 173.305 ;
        RECT 68.300 172.685 69.210 172.765 ;
        RECT 67.470 172.205 67.790 172.685 ;
        RECT 67.960 172.595 69.210 172.685 ;
        RECT 67.960 172.515 68.470 172.595 ;
        RECT 67.960 172.115 68.190 172.515 ;
        RECT 68.360 171.945 68.710 172.335 ;
        RECT 68.880 172.115 69.210 172.595 ;
        RECT 69.380 171.945 69.550 172.765 ;
        RECT 70.350 172.685 70.520 173.645 ;
        RECT 70.690 173.355 70.950 174.495 ;
        RECT 71.120 173.525 71.450 174.325 ;
        RECT 71.620 173.695 71.790 174.495 ;
        RECT 71.990 173.525 72.320 174.325 ;
        RECT 72.520 173.695 72.800 174.495 ;
        RECT 71.120 173.355 72.400 173.525 ;
        RECT 70.715 172.855 71.000 173.185 ;
        RECT 71.200 172.855 71.580 173.185 ;
        RECT 71.750 172.855 72.060 173.185 ;
        RECT 70.055 172.140 70.520 172.685 ;
        RECT 70.695 171.945 71.030 172.685 ;
        RECT 71.200 172.160 71.415 172.855 ;
        RECT 71.750 172.685 71.955 172.855 ;
        RECT 72.230 172.685 72.400 173.355 ;
        RECT 72.580 172.855 72.820 173.525 ;
        RECT 73.950 173.355 74.180 174.495 ;
        RECT 74.350 173.345 74.680 174.325 ;
        RECT 74.850 173.355 75.060 174.495 ;
        RECT 75.290 173.735 75.805 174.145 ;
        RECT 76.040 173.735 76.210 174.495 ;
        RECT 76.380 174.155 78.410 174.325 ;
        RECT 73.930 172.935 74.260 173.185 ;
        RECT 71.605 172.160 71.955 172.685 ;
        RECT 72.125 172.115 72.820 172.685 ;
        RECT 73.950 171.945 74.180 172.765 ;
        RECT 74.430 172.745 74.680 173.345 ;
        RECT 75.290 172.925 75.630 173.735 ;
        RECT 76.380 173.490 76.550 174.155 ;
        RECT 76.945 173.815 78.070 173.985 ;
        RECT 75.800 173.300 76.550 173.490 ;
        RECT 76.720 173.475 77.730 173.645 ;
        RECT 74.350 172.115 74.680 172.745 ;
        RECT 74.850 171.945 75.060 172.765 ;
        RECT 75.290 172.755 76.520 172.925 ;
        RECT 75.565 172.150 75.810 172.755 ;
        RECT 76.030 171.945 76.540 172.480 ;
        RECT 76.720 172.115 76.910 173.475 ;
        RECT 77.080 172.455 77.355 173.275 ;
        RECT 77.560 172.675 77.730 173.475 ;
        RECT 77.900 172.685 78.070 173.815 ;
        RECT 78.240 173.185 78.410 174.155 ;
        RECT 78.580 173.355 78.750 174.495 ;
        RECT 78.920 173.355 79.255 174.325 ;
        RECT 78.240 172.855 78.435 173.185 ;
        RECT 78.660 172.855 78.915 173.185 ;
        RECT 78.660 172.685 78.830 172.855 ;
        RECT 79.085 172.685 79.255 173.355 ;
        RECT 77.900 172.515 78.830 172.685 ;
        RECT 77.900 172.480 78.075 172.515 ;
        RECT 77.080 172.285 77.360 172.455 ;
        RECT 77.080 172.115 77.355 172.285 ;
        RECT 77.545 172.115 78.075 172.480 ;
        RECT 78.500 171.945 78.830 172.345 ;
        RECT 79.000 172.115 79.255 172.685 ;
        RECT 80.350 173.420 80.620 174.325 ;
        RECT 80.790 173.735 81.120 174.495 ;
        RECT 81.300 173.565 81.470 174.325 ;
        RECT 80.350 172.620 80.520 173.420 ;
        RECT 80.805 173.395 81.470 173.565 ;
        RECT 81.730 173.420 82.000 174.325 ;
        RECT 82.170 173.735 82.500 174.495 ;
        RECT 82.680 173.565 82.850 174.325 ;
        RECT 80.805 173.250 80.975 173.395 ;
        RECT 80.690 172.920 80.975 173.250 ;
        RECT 80.805 172.665 80.975 172.920 ;
        RECT 81.210 172.845 81.540 173.215 ;
        RECT 80.350 172.115 80.610 172.620 ;
        RECT 80.805 172.495 81.470 172.665 ;
        RECT 80.790 171.945 81.120 172.325 ;
        RECT 81.300 172.115 81.470 172.495 ;
        RECT 81.730 172.620 81.900 173.420 ;
        RECT 82.185 173.395 82.850 173.565 ;
        RECT 83.110 173.405 84.780 174.495 ;
        RECT 82.185 173.250 82.355 173.395 ;
        RECT 82.070 172.920 82.355 173.250 ;
        RECT 82.185 172.665 82.355 172.920 ;
        RECT 82.590 172.845 82.920 173.215 ;
        RECT 83.110 172.885 83.860 173.405 ;
        RECT 84.990 173.355 85.220 174.495 ;
        RECT 85.390 173.345 85.720 174.325 ;
        RECT 85.890 173.355 86.100 174.495 ;
        RECT 84.030 172.715 84.780 173.235 ;
        RECT 84.970 172.935 85.300 173.185 ;
        RECT 81.730 172.115 81.990 172.620 ;
        RECT 82.185 172.495 82.850 172.665 ;
        RECT 82.170 171.945 82.500 172.325 ;
        RECT 82.680 172.115 82.850 172.495 ;
        RECT 83.110 171.945 84.780 172.715 ;
        RECT 84.990 171.945 85.220 172.765 ;
        RECT 85.470 172.745 85.720 173.345 ;
        RECT 86.330 173.330 86.620 174.495 ;
        RECT 86.795 173.305 87.050 174.185 ;
        RECT 87.220 173.355 87.525 174.495 ;
        RECT 87.865 174.115 88.195 174.495 ;
        RECT 88.375 173.945 88.545 174.235 ;
        RECT 88.715 174.035 88.965 174.495 ;
        RECT 87.745 173.775 88.545 173.945 ;
        RECT 89.135 173.985 90.005 174.325 ;
        RECT 85.390 172.115 85.720 172.745 ;
        RECT 85.890 171.945 86.100 172.765 ;
        RECT 86.330 171.945 86.620 172.670 ;
        RECT 86.795 172.655 87.005 173.305 ;
        RECT 87.745 173.185 87.915 173.775 ;
        RECT 89.135 173.605 89.305 173.985 ;
        RECT 90.240 173.865 90.410 174.325 ;
        RECT 90.580 174.035 90.950 174.495 ;
        RECT 91.245 173.895 91.415 174.235 ;
        RECT 91.585 174.065 91.915 174.495 ;
        RECT 92.150 173.895 92.320 174.235 ;
        RECT 88.085 173.435 89.305 173.605 ;
        RECT 89.475 173.525 89.935 173.815 ;
        RECT 90.240 173.695 90.800 173.865 ;
        RECT 91.245 173.725 92.320 173.895 ;
        RECT 92.490 173.995 93.170 174.325 ;
        RECT 93.385 173.995 93.635 174.325 ;
        RECT 93.805 174.035 94.055 174.495 ;
        RECT 90.630 173.555 90.800 173.695 ;
        RECT 89.475 173.515 90.440 173.525 ;
        RECT 89.135 173.345 89.305 173.435 ;
        RECT 89.765 173.355 90.440 173.515 ;
        RECT 87.175 173.155 87.915 173.185 ;
        RECT 87.175 172.855 88.090 173.155 ;
        RECT 87.765 172.680 88.090 172.855 ;
        RECT 86.795 172.125 87.050 172.655 ;
        RECT 87.220 171.945 87.525 172.405 ;
        RECT 87.770 172.325 88.090 172.680 ;
        RECT 88.260 172.895 88.800 173.265 ;
        RECT 89.135 173.175 89.540 173.345 ;
        RECT 88.260 172.495 88.500 172.895 ;
        RECT 88.980 172.725 89.200 173.005 ;
        RECT 88.670 172.555 89.200 172.725 ;
        RECT 88.670 172.325 88.840 172.555 ;
        RECT 89.370 172.395 89.540 173.175 ;
        RECT 89.710 172.565 90.060 173.185 ;
        RECT 90.230 172.565 90.440 173.355 ;
        RECT 90.630 173.385 92.130 173.555 ;
        RECT 90.630 172.695 90.800 173.385 ;
        RECT 92.490 173.215 92.660 173.995 ;
        RECT 93.465 173.865 93.635 173.995 ;
        RECT 90.970 173.045 92.660 173.215 ;
        RECT 92.830 173.435 93.295 173.825 ;
        RECT 93.465 173.695 93.860 173.865 ;
        RECT 90.970 172.865 91.140 173.045 ;
        RECT 87.770 172.155 88.840 172.325 ;
        RECT 89.010 171.945 89.200 172.385 ;
        RECT 89.370 172.115 90.320 172.395 ;
        RECT 90.630 172.305 90.890 172.695 ;
        RECT 91.310 172.625 92.100 172.875 ;
        RECT 90.540 172.135 90.890 172.305 ;
        RECT 91.100 171.945 91.430 172.405 ;
        RECT 92.305 172.335 92.475 173.045 ;
        RECT 92.830 172.845 93.000 173.435 ;
        RECT 92.645 172.625 93.000 172.845 ;
        RECT 93.170 172.625 93.520 173.245 ;
        RECT 93.690 172.335 93.860 173.695 ;
        RECT 94.225 173.525 94.550 174.310 ;
        RECT 94.030 172.475 94.490 173.525 ;
        RECT 92.305 172.165 93.160 172.335 ;
        RECT 93.365 172.165 93.860 172.335 ;
        RECT 94.030 171.945 94.360 172.305 ;
        RECT 94.720 172.205 94.890 174.325 ;
        RECT 95.060 173.995 95.390 174.495 ;
        RECT 95.560 173.825 95.815 174.325 ;
        RECT 95.065 173.655 95.815 173.825 ;
        RECT 95.990 173.735 96.505 174.145 ;
        RECT 96.740 173.735 96.910 174.495 ;
        RECT 97.080 174.155 99.110 174.325 ;
        RECT 95.065 172.665 95.295 173.655 ;
        RECT 95.465 172.835 95.815 173.485 ;
        RECT 95.990 172.925 96.330 173.735 ;
        RECT 97.080 173.490 97.250 174.155 ;
        RECT 97.645 173.815 98.770 173.985 ;
        RECT 96.500 173.300 97.250 173.490 ;
        RECT 97.420 173.475 98.430 173.645 ;
        RECT 95.990 172.755 97.220 172.925 ;
        RECT 95.065 172.495 95.815 172.665 ;
        RECT 95.060 171.945 95.390 172.325 ;
        RECT 95.560 172.205 95.815 172.495 ;
        RECT 96.265 172.150 96.510 172.755 ;
        RECT 96.730 171.945 97.240 172.480 ;
        RECT 97.420 172.115 97.610 173.475 ;
        RECT 97.780 172.795 98.055 173.275 ;
        RECT 97.780 172.625 98.060 172.795 ;
        RECT 98.260 172.675 98.430 173.475 ;
        RECT 98.600 172.685 98.770 173.815 ;
        RECT 98.940 173.185 99.110 174.155 ;
        RECT 99.280 173.355 99.450 174.495 ;
        RECT 99.620 173.355 99.955 174.325 ;
        RECT 98.940 172.855 99.135 173.185 ;
        RECT 99.360 172.855 99.615 173.185 ;
        RECT 99.360 172.685 99.530 172.855 ;
        RECT 99.785 172.685 99.955 173.355 ;
        RECT 97.780 172.115 98.055 172.625 ;
        RECT 98.600 172.515 99.530 172.685 ;
        RECT 98.600 172.480 98.775 172.515 ;
        RECT 98.245 172.115 98.775 172.480 ;
        RECT 99.200 171.945 99.530 172.345 ;
        RECT 99.700 172.115 99.955 172.685 ;
        RECT 101.055 173.305 101.310 174.185 ;
        RECT 101.480 173.355 101.785 174.495 ;
        RECT 102.125 174.115 102.455 174.495 ;
        RECT 102.635 173.945 102.805 174.235 ;
        RECT 102.975 174.035 103.225 174.495 ;
        RECT 102.005 173.775 102.805 173.945 ;
        RECT 103.395 173.985 104.265 174.325 ;
        RECT 101.055 172.655 101.265 173.305 ;
        RECT 102.005 173.185 102.175 173.775 ;
        RECT 103.395 173.605 103.565 173.985 ;
        RECT 104.500 173.865 104.670 174.325 ;
        RECT 104.840 174.035 105.210 174.495 ;
        RECT 105.505 173.895 105.675 174.235 ;
        RECT 105.845 174.065 106.175 174.495 ;
        RECT 106.410 173.895 106.580 174.235 ;
        RECT 102.345 173.435 103.565 173.605 ;
        RECT 103.735 173.525 104.195 173.815 ;
        RECT 104.500 173.695 105.060 173.865 ;
        RECT 105.505 173.725 106.580 173.895 ;
        RECT 106.750 173.995 107.430 174.325 ;
        RECT 107.645 173.995 107.895 174.325 ;
        RECT 108.065 174.035 108.315 174.495 ;
        RECT 104.890 173.555 105.060 173.695 ;
        RECT 103.735 173.515 104.700 173.525 ;
        RECT 103.395 173.345 103.565 173.435 ;
        RECT 104.025 173.355 104.700 173.515 ;
        RECT 101.435 173.155 102.175 173.185 ;
        RECT 101.435 172.855 102.350 173.155 ;
        RECT 102.025 172.680 102.350 172.855 ;
        RECT 101.055 172.125 101.310 172.655 ;
        RECT 101.480 171.945 101.785 172.405 ;
        RECT 102.030 172.325 102.350 172.680 ;
        RECT 102.520 172.895 103.060 173.265 ;
        RECT 103.395 173.175 103.800 173.345 ;
        RECT 102.520 172.495 102.760 172.895 ;
        RECT 103.240 172.725 103.460 173.005 ;
        RECT 102.930 172.555 103.460 172.725 ;
        RECT 102.930 172.325 103.100 172.555 ;
        RECT 103.630 172.395 103.800 173.175 ;
        RECT 103.970 172.565 104.320 173.185 ;
        RECT 104.490 172.565 104.700 173.355 ;
        RECT 104.890 173.385 106.390 173.555 ;
        RECT 104.890 172.695 105.060 173.385 ;
        RECT 106.750 173.215 106.920 173.995 ;
        RECT 107.725 173.865 107.895 173.995 ;
        RECT 105.230 173.045 106.920 173.215 ;
        RECT 107.090 173.435 107.555 173.825 ;
        RECT 107.725 173.695 108.120 173.865 ;
        RECT 105.230 172.865 105.400 173.045 ;
        RECT 102.030 172.155 103.100 172.325 ;
        RECT 103.270 171.945 103.460 172.385 ;
        RECT 103.630 172.115 104.580 172.395 ;
        RECT 104.890 172.305 105.150 172.695 ;
        RECT 105.570 172.625 106.360 172.875 ;
        RECT 104.800 172.135 105.150 172.305 ;
        RECT 105.360 171.945 105.690 172.405 ;
        RECT 106.565 172.335 106.735 173.045 ;
        RECT 107.090 172.845 107.260 173.435 ;
        RECT 106.905 172.625 107.260 172.845 ;
        RECT 107.430 172.625 107.780 173.245 ;
        RECT 107.950 172.335 108.120 173.695 ;
        RECT 108.485 173.525 108.810 174.310 ;
        RECT 108.290 172.475 108.750 173.525 ;
        RECT 106.565 172.165 107.420 172.335 ;
        RECT 107.625 172.165 108.120 172.335 ;
        RECT 108.290 171.945 108.620 172.305 ;
        RECT 108.980 172.205 109.150 174.325 ;
        RECT 109.320 173.995 109.650 174.495 ;
        RECT 109.820 173.825 110.075 174.325 ;
        RECT 109.325 173.655 110.075 173.825 ;
        RECT 109.325 172.665 109.555 173.655 ;
        RECT 109.725 172.835 110.075 173.485 ;
        RECT 111.170 173.405 112.380 174.495 ;
        RECT 111.170 172.865 111.690 173.405 ;
        RECT 111.860 172.695 112.380 173.235 ;
        RECT 109.325 172.495 110.075 172.665 ;
        RECT 109.320 171.945 109.650 172.325 ;
        RECT 109.820 172.205 110.075 172.495 ;
        RECT 111.170 171.945 112.380 172.695 ;
        RECT 18.165 171.775 112.465 171.945 ;
        RECT 18.250 171.025 19.460 171.775 ;
        RECT 18.250 170.485 18.770 171.025 ;
        RECT 20.090 171.005 21.760 171.775 ;
        RECT 21.930 171.050 22.220 171.775 ;
        RECT 22.850 171.005 25.440 171.775 ;
        RECT 18.940 170.315 19.460 170.855 ;
        RECT 18.250 169.225 19.460 170.315 ;
        RECT 20.090 170.315 20.840 170.835 ;
        RECT 21.010 170.485 21.760 171.005 ;
        RECT 20.090 169.225 21.760 170.315 ;
        RECT 21.930 169.225 22.220 170.390 ;
        RECT 22.850 170.315 24.060 170.835 ;
        RECT 24.230 170.485 25.440 171.005 ;
        RECT 25.650 170.955 25.880 171.775 ;
        RECT 26.050 170.975 26.380 171.605 ;
        RECT 25.630 170.535 25.960 170.785 ;
        RECT 26.130 170.375 26.380 170.975 ;
        RECT 26.550 170.955 26.760 171.775 ;
        RECT 27.030 170.955 27.260 171.775 ;
        RECT 27.430 170.975 27.760 171.605 ;
        RECT 27.010 170.535 27.340 170.785 ;
        RECT 27.510 170.375 27.760 170.975 ;
        RECT 27.930 170.955 28.140 171.775 ;
        RECT 28.460 171.225 28.630 171.605 ;
        RECT 28.810 171.395 29.140 171.775 ;
        RECT 28.460 171.055 29.125 171.225 ;
        RECT 29.320 171.100 29.580 171.605 ;
        RECT 28.390 170.505 28.720 170.875 ;
        RECT 28.955 170.800 29.125 171.055 ;
        RECT 22.850 169.225 25.440 170.315 ;
        RECT 25.650 169.225 25.880 170.365 ;
        RECT 26.050 169.395 26.380 170.375 ;
        RECT 26.550 169.225 26.760 170.365 ;
        RECT 27.030 169.225 27.260 170.365 ;
        RECT 27.430 169.395 27.760 170.375 ;
        RECT 28.955 170.470 29.240 170.800 ;
        RECT 27.930 169.225 28.140 170.365 ;
        RECT 28.955 170.325 29.125 170.470 ;
        RECT 28.460 170.155 29.125 170.325 ;
        RECT 29.410 170.300 29.580 171.100 ;
        RECT 28.460 169.395 28.630 170.155 ;
        RECT 28.810 169.225 29.140 169.985 ;
        RECT 29.310 169.395 29.580 170.300 ;
        RECT 29.750 170.975 30.090 171.605 ;
        RECT 30.260 170.975 30.510 171.775 ;
        RECT 30.700 171.125 31.030 171.605 ;
        RECT 31.200 171.315 31.425 171.775 ;
        RECT 31.595 171.125 31.925 171.605 ;
        RECT 29.750 170.415 29.925 170.975 ;
        RECT 30.700 170.955 31.925 171.125 ;
        RECT 32.555 170.995 33.055 171.605 ;
        RECT 33.435 171.225 33.690 171.515 ;
        RECT 33.860 171.395 34.190 171.775 ;
        RECT 33.435 171.055 34.185 171.225 ;
        RECT 30.095 170.615 30.790 170.785 ;
        RECT 29.750 170.365 29.980 170.415 ;
        RECT 30.620 170.365 30.790 170.615 ;
        RECT 30.965 170.585 31.385 170.785 ;
        RECT 31.555 170.585 31.885 170.785 ;
        RECT 32.055 170.585 32.385 170.785 ;
        RECT 32.555 170.365 32.725 170.995 ;
        RECT 32.910 170.535 33.260 170.785 ;
        RECT 29.750 169.395 30.090 170.365 ;
        RECT 30.260 169.225 30.430 170.365 ;
        RECT 30.620 170.195 33.055 170.365 ;
        RECT 33.435 170.235 33.785 170.885 ;
        RECT 30.700 169.225 30.950 170.025 ;
        RECT 31.595 169.395 31.925 170.195 ;
        RECT 32.225 169.225 32.555 170.025 ;
        RECT 32.725 169.395 33.055 170.195 ;
        RECT 33.955 170.065 34.185 171.055 ;
        RECT 33.435 169.895 34.185 170.065 ;
        RECT 33.435 169.395 33.690 169.895 ;
        RECT 33.860 169.225 34.190 169.725 ;
        RECT 34.360 169.395 34.530 171.515 ;
        RECT 34.890 171.415 35.220 171.775 ;
        RECT 35.390 171.385 35.885 171.555 ;
        RECT 36.090 171.385 36.945 171.555 ;
        RECT 34.760 170.195 35.220 171.245 ;
        RECT 34.700 169.410 35.025 170.195 ;
        RECT 35.390 170.025 35.560 171.385 ;
        RECT 35.730 170.475 36.080 171.095 ;
        RECT 36.250 170.875 36.605 171.095 ;
        RECT 36.250 170.285 36.420 170.875 ;
        RECT 36.775 170.675 36.945 171.385 ;
        RECT 37.820 171.315 38.150 171.775 ;
        RECT 38.360 171.415 38.710 171.585 ;
        RECT 37.150 170.845 37.940 171.095 ;
        RECT 38.360 171.025 38.620 171.415 ;
        RECT 38.930 171.325 39.880 171.605 ;
        RECT 40.050 171.335 40.240 171.775 ;
        RECT 40.410 171.395 41.480 171.565 ;
        RECT 38.110 170.675 38.280 170.855 ;
        RECT 35.390 169.855 35.785 170.025 ;
        RECT 35.955 169.895 36.420 170.285 ;
        RECT 36.590 170.505 38.280 170.675 ;
        RECT 35.615 169.725 35.785 169.855 ;
        RECT 36.590 169.725 36.760 170.505 ;
        RECT 38.450 170.335 38.620 171.025 ;
        RECT 37.120 170.165 38.620 170.335 ;
        RECT 38.810 170.365 39.020 171.155 ;
        RECT 39.190 170.535 39.540 171.155 ;
        RECT 39.710 170.545 39.880 171.325 ;
        RECT 40.410 171.165 40.580 171.395 ;
        RECT 40.050 170.995 40.580 171.165 ;
        RECT 40.050 170.715 40.270 170.995 ;
        RECT 40.750 170.825 40.990 171.225 ;
        RECT 39.710 170.375 40.115 170.545 ;
        RECT 40.450 170.455 40.990 170.825 ;
        RECT 41.160 171.040 41.480 171.395 ;
        RECT 41.725 171.315 42.030 171.775 ;
        RECT 42.200 171.065 42.455 171.595 ;
        RECT 41.160 170.865 41.485 171.040 ;
        RECT 41.160 170.565 42.075 170.865 ;
        RECT 41.335 170.535 42.075 170.565 ;
        RECT 38.810 170.205 39.485 170.365 ;
        RECT 39.945 170.285 40.115 170.375 ;
        RECT 38.810 170.195 39.775 170.205 ;
        RECT 38.450 170.025 38.620 170.165 ;
        RECT 35.195 169.225 35.445 169.685 ;
        RECT 35.615 169.395 35.865 169.725 ;
        RECT 36.080 169.395 36.760 169.725 ;
        RECT 36.930 169.825 38.005 169.995 ;
        RECT 38.450 169.855 39.010 170.025 ;
        RECT 39.315 169.905 39.775 170.195 ;
        RECT 39.945 170.115 41.165 170.285 ;
        RECT 36.930 169.485 37.100 169.825 ;
        RECT 37.335 169.225 37.665 169.655 ;
        RECT 37.835 169.485 38.005 169.825 ;
        RECT 38.300 169.225 38.670 169.685 ;
        RECT 38.840 169.395 39.010 169.855 ;
        RECT 39.945 169.735 40.115 170.115 ;
        RECT 41.335 169.945 41.505 170.535 ;
        RECT 42.245 170.415 42.455 171.065 ;
        RECT 43.090 171.005 45.680 171.775 ;
        RECT 39.245 169.395 40.115 169.735 ;
        RECT 40.705 169.775 41.505 169.945 ;
        RECT 40.285 169.225 40.535 169.685 ;
        RECT 40.705 169.485 40.875 169.775 ;
        RECT 41.055 169.225 41.385 169.605 ;
        RECT 41.725 169.225 42.030 170.365 ;
        RECT 42.200 169.535 42.455 170.415 ;
        RECT 43.090 170.315 44.300 170.835 ;
        RECT 44.470 170.485 45.680 171.005 ;
        RECT 45.850 171.100 46.110 171.605 ;
        RECT 46.290 171.395 46.620 171.775 ;
        RECT 46.800 171.225 46.970 171.605 ;
        RECT 43.090 169.225 45.680 170.315 ;
        RECT 45.850 170.300 46.020 171.100 ;
        RECT 46.305 171.055 46.970 171.225 ;
        RECT 46.305 170.800 46.475 171.055 ;
        RECT 47.690 171.050 47.980 171.775 ;
        RECT 48.650 170.955 48.880 171.775 ;
        RECT 49.050 170.975 49.380 171.605 ;
        RECT 46.190 170.470 46.475 170.800 ;
        RECT 46.710 170.505 47.040 170.875 ;
        RECT 48.630 170.535 48.960 170.785 ;
        RECT 46.305 170.325 46.475 170.470 ;
        RECT 45.850 169.395 46.120 170.300 ;
        RECT 46.305 170.155 46.970 170.325 ;
        RECT 46.290 169.225 46.620 169.985 ;
        RECT 46.800 169.395 46.970 170.155 ;
        RECT 47.690 169.225 47.980 170.390 ;
        RECT 49.130 170.375 49.380 170.975 ;
        RECT 49.550 170.955 49.760 171.775 ;
        RECT 50.265 170.965 50.510 171.570 ;
        RECT 50.730 171.240 51.240 171.775 ;
        RECT 48.650 169.225 48.880 170.365 ;
        RECT 49.050 169.395 49.380 170.375 ;
        RECT 49.990 170.795 51.220 170.965 ;
        RECT 49.550 169.225 49.760 170.365 ;
        RECT 49.990 169.985 50.330 170.795 ;
        RECT 50.500 170.230 51.250 170.420 ;
        RECT 49.990 169.575 50.505 169.985 ;
        RECT 50.740 169.225 50.910 169.985 ;
        RECT 51.080 169.565 51.250 170.230 ;
        RECT 51.420 170.245 51.610 171.605 ;
        RECT 51.780 170.755 52.055 171.605 ;
        RECT 52.245 171.240 52.775 171.605 ;
        RECT 53.200 171.375 53.530 171.775 ;
        RECT 52.600 171.205 52.775 171.240 ;
        RECT 51.780 170.585 52.060 170.755 ;
        RECT 51.780 170.445 52.055 170.585 ;
        RECT 52.260 170.245 52.430 171.045 ;
        RECT 51.420 170.075 52.430 170.245 ;
        RECT 52.600 171.035 53.530 171.205 ;
        RECT 53.700 171.035 53.955 171.605 ;
        RECT 54.220 171.225 54.390 171.605 ;
        RECT 54.570 171.395 54.900 171.775 ;
        RECT 54.220 171.055 54.885 171.225 ;
        RECT 55.080 171.100 55.340 171.605 ;
        RECT 52.600 169.905 52.770 171.035 ;
        RECT 53.360 170.865 53.530 171.035 ;
        RECT 51.645 169.735 52.770 169.905 ;
        RECT 52.940 170.535 53.135 170.865 ;
        RECT 53.360 170.535 53.615 170.865 ;
        RECT 52.940 169.565 53.110 170.535 ;
        RECT 53.785 170.365 53.955 171.035 ;
        RECT 54.150 170.505 54.480 170.875 ;
        RECT 54.715 170.800 54.885 171.055 ;
        RECT 51.080 169.395 53.110 169.565 ;
        RECT 53.280 169.225 53.450 170.365 ;
        RECT 53.620 169.395 53.955 170.365 ;
        RECT 54.715 170.470 55.000 170.800 ;
        RECT 54.715 170.325 54.885 170.470 ;
        RECT 54.220 170.155 54.885 170.325 ;
        RECT 55.170 170.300 55.340 171.100 ;
        RECT 55.625 171.145 55.910 171.605 ;
        RECT 56.080 171.315 56.350 171.775 ;
        RECT 55.625 170.975 56.580 171.145 ;
        RECT 54.220 169.395 54.390 170.155 ;
        RECT 54.570 169.225 54.900 169.985 ;
        RECT 55.070 169.395 55.340 170.300 ;
        RECT 55.510 170.245 56.200 170.805 ;
        RECT 56.370 170.075 56.580 170.975 ;
        RECT 55.625 169.855 56.580 170.075 ;
        RECT 56.750 170.805 57.150 171.605 ;
        RECT 57.340 171.145 57.620 171.605 ;
        RECT 58.140 171.315 58.465 171.775 ;
        RECT 57.340 170.975 58.465 171.145 ;
        RECT 58.635 171.035 59.020 171.605 ;
        RECT 58.015 170.865 58.465 170.975 ;
        RECT 56.750 170.245 57.845 170.805 ;
        RECT 58.015 170.535 58.570 170.865 ;
        RECT 55.625 169.395 55.910 169.855 ;
        RECT 56.080 169.225 56.350 169.685 ;
        RECT 56.750 169.395 57.150 170.245 ;
        RECT 58.015 170.075 58.465 170.535 ;
        RECT 58.740 170.365 59.020 171.035 ;
        RECT 57.340 169.855 58.465 170.075 ;
        RECT 57.340 169.395 57.620 169.855 ;
        RECT 58.140 169.225 58.465 169.685 ;
        RECT 58.635 169.395 59.020 170.365 ;
        RECT 59.195 171.065 59.450 171.595 ;
        RECT 59.620 171.315 59.925 171.775 ;
        RECT 60.170 171.395 61.240 171.565 ;
        RECT 59.195 170.415 59.405 171.065 ;
        RECT 60.170 171.040 60.490 171.395 ;
        RECT 60.165 170.865 60.490 171.040 ;
        RECT 59.575 170.565 60.490 170.865 ;
        RECT 60.660 170.825 60.900 171.225 ;
        RECT 61.070 171.165 61.240 171.395 ;
        RECT 61.410 171.335 61.600 171.775 ;
        RECT 61.770 171.325 62.720 171.605 ;
        RECT 62.940 171.415 63.290 171.585 ;
        RECT 61.070 170.995 61.600 171.165 ;
        RECT 59.575 170.535 60.315 170.565 ;
        RECT 59.195 169.535 59.450 170.415 ;
        RECT 59.620 169.225 59.925 170.365 ;
        RECT 60.145 169.945 60.315 170.535 ;
        RECT 60.660 170.455 61.200 170.825 ;
        RECT 61.380 170.715 61.600 170.995 ;
        RECT 61.770 170.545 61.940 171.325 ;
        RECT 61.535 170.375 61.940 170.545 ;
        RECT 62.110 170.535 62.460 171.155 ;
        RECT 61.535 170.285 61.705 170.375 ;
        RECT 62.630 170.365 62.840 171.155 ;
        RECT 60.485 170.115 61.705 170.285 ;
        RECT 62.165 170.205 62.840 170.365 ;
        RECT 60.145 169.775 60.945 169.945 ;
        RECT 60.265 169.225 60.595 169.605 ;
        RECT 60.775 169.485 60.945 169.775 ;
        RECT 61.535 169.735 61.705 170.115 ;
        RECT 61.875 170.195 62.840 170.205 ;
        RECT 63.030 171.025 63.290 171.415 ;
        RECT 63.500 171.315 63.830 171.775 ;
        RECT 64.705 171.385 65.560 171.555 ;
        RECT 65.765 171.385 66.260 171.555 ;
        RECT 66.430 171.415 66.760 171.775 ;
        RECT 63.030 170.335 63.200 171.025 ;
        RECT 63.370 170.675 63.540 170.855 ;
        RECT 63.710 170.845 64.500 171.095 ;
        RECT 64.705 170.675 64.875 171.385 ;
        RECT 65.045 170.875 65.400 171.095 ;
        RECT 63.370 170.505 65.060 170.675 ;
        RECT 61.875 169.905 62.335 170.195 ;
        RECT 63.030 170.165 64.530 170.335 ;
        RECT 63.030 170.025 63.200 170.165 ;
        RECT 62.640 169.855 63.200 170.025 ;
        RECT 61.115 169.225 61.365 169.685 ;
        RECT 61.535 169.395 62.405 169.735 ;
        RECT 62.640 169.395 62.810 169.855 ;
        RECT 63.645 169.825 64.720 169.995 ;
        RECT 62.980 169.225 63.350 169.685 ;
        RECT 63.645 169.485 63.815 169.825 ;
        RECT 63.985 169.225 64.315 169.655 ;
        RECT 64.550 169.485 64.720 169.825 ;
        RECT 64.890 169.725 65.060 170.505 ;
        RECT 65.230 170.285 65.400 170.875 ;
        RECT 65.570 170.475 65.920 171.095 ;
        RECT 65.230 169.895 65.695 170.285 ;
        RECT 66.090 170.025 66.260 171.385 ;
        RECT 66.430 170.195 66.890 171.245 ;
        RECT 65.865 169.855 66.260 170.025 ;
        RECT 65.865 169.725 66.035 169.855 ;
        RECT 64.890 169.395 65.570 169.725 ;
        RECT 65.785 169.395 66.035 169.725 ;
        RECT 66.205 169.225 66.455 169.685 ;
        RECT 66.625 169.410 66.950 170.195 ;
        RECT 67.120 169.395 67.290 171.515 ;
        RECT 67.460 171.395 67.790 171.775 ;
        RECT 67.960 171.225 68.215 171.515 ;
        RECT 67.465 171.055 68.215 171.225 ;
        RECT 68.480 171.125 68.650 171.605 ;
        RECT 68.830 171.295 69.070 171.775 ;
        RECT 69.320 171.125 69.490 171.605 ;
        RECT 69.660 171.295 69.990 171.775 ;
        RECT 70.160 171.125 70.330 171.605 ;
        RECT 67.465 170.065 67.695 171.055 ;
        RECT 68.480 170.955 69.115 171.125 ;
        RECT 69.320 170.955 70.330 171.125 ;
        RECT 70.500 170.975 70.830 171.775 ;
        RECT 71.610 171.005 73.280 171.775 ;
        RECT 73.450 171.050 73.740 171.775 ;
        RECT 67.865 170.235 68.215 170.885 ;
        RECT 68.945 170.785 69.115 170.955 ;
        RECT 69.830 170.925 70.330 170.955 ;
        RECT 68.395 170.545 68.775 170.785 ;
        RECT 68.945 170.615 69.445 170.785 ;
        RECT 68.945 170.375 69.115 170.615 ;
        RECT 69.835 170.415 70.330 170.925 ;
        RECT 68.400 170.205 69.115 170.375 ;
        RECT 69.320 170.245 70.330 170.415 ;
        RECT 67.465 169.895 68.215 170.065 ;
        RECT 67.460 169.225 67.790 169.725 ;
        RECT 67.960 169.395 68.215 169.895 ;
        RECT 68.400 169.395 68.730 170.205 ;
        RECT 68.900 169.225 69.140 170.025 ;
        RECT 69.320 169.395 69.490 170.245 ;
        RECT 69.660 169.225 69.990 170.025 ;
        RECT 70.160 169.395 70.330 170.245 ;
        RECT 70.500 169.225 70.830 170.375 ;
        RECT 71.610 170.315 72.360 170.835 ;
        RECT 72.530 170.485 73.280 171.005 ;
        RECT 74.870 170.955 75.100 171.775 ;
        RECT 75.270 170.975 75.600 171.605 ;
        RECT 74.850 170.535 75.180 170.785 ;
        RECT 71.610 169.225 73.280 170.315 ;
        RECT 73.450 169.225 73.740 170.390 ;
        RECT 75.350 170.375 75.600 170.975 ;
        RECT 75.770 170.955 75.980 171.775 ;
        RECT 76.215 171.065 76.470 171.595 ;
        RECT 76.640 171.315 76.945 171.775 ;
        RECT 77.190 171.395 78.260 171.565 ;
        RECT 74.870 169.225 75.100 170.365 ;
        RECT 75.270 169.395 75.600 170.375 ;
        RECT 76.215 170.415 76.425 171.065 ;
        RECT 77.190 171.040 77.510 171.395 ;
        RECT 77.185 170.865 77.510 171.040 ;
        RECT 76.595 170.565 77.510 170.865 ;
        RECT 77.680 170.825 77.920 171.225 ;
        RECT 78.090 171.165 78.260 171.395 ;
        RECT 78.430 171.335 78.620 171.775 ;
        RECT 78.790 171.325 79.740 171.605 ;
        RECT 79.960 171.415 80.310 171.585 ;
        RECT 78.090 170.995 78.620 171.165 ;
        RECT 76.595 170.535 77.335 170.565 ;
        RECT 75.770 169.225 75.980 170.365 ;
        RECT 76.215 169.535 76.470 170.415 ;
        RECT 76.640 169.225 76.945 170.365 ;
        RECT 77.165 169.945 77.335 170.535 ;
        RECT 77.680 170.455 78.220 170.825 ;
        RECT 78.400 170.715 78.620 170.995 ;
        RECT 78.790 170.545 78.960 171.325 ;
        RECT 78.555 170.375 78.960 170.545 ;
        RECT 79.130 170.535 79.480 171.155 ;
        RECT 78.555 170.285 78.725 170.375 ;
        RECT 79.650 170.365 79.860 171.155 ;
        RECT 77.505 170.115 78.725 170.285 ;
        RECT 79.185 170.205 79.860 170.365 ;
        RECT 77.165 169.775 77.965 169.945 ;
        RECT 77.285 169.225 77.615 169.605 ;
        RECT 77.795 169.485 77.965 169.775 ;
        RECT 78.555 169.735 78.725 170.115 ;
        RECT 78.895 170.195 79.860 170.205 ;
        RECT 80.050 171.025 80.310 171.415 ;
        RECT 80.520 171.315 80.850 171.775 ;
        RECT 81.725 171.385 82.580 171.555 ;
        RECT 82.785 171.385 83.280 171.555 ;
        RECT 83.450 171.415 83.780 171.775 ;
        RECT 80.050 170.335 80.220 171.025 ;
        RECT 80.390 170.675 80.560 170.855 ;
        RECT 80.730 170.845 81.520 171.095 ;
        RECT 81.725 170.675 81.895 171.385 ;
        RECT 82.065 170.875 82.420 171.095 ;
        RECT 80.390 170.505 82.080 170.675 ;
        RECT 78.895 169.905 79.355 170.195 ;
        RECT 80.050 170.165 81.550 170.335 ;
        RECT 80.050 170.025 80.220 170.165 ;
        RECT 79.660 169.855 80.220 170.025 ;
        RECT 78.135 169.225 78.385 169.685 ;
        RECT 78.555 169.395 79.425 169.735 ;
        RECT 79.660 169.395 79.830 169.855 ;
        RECT 80.665 169.825 81.740 169.995 ;
        RECT 80.000 169.225 80.370 169.685 ;
        RECT 80.665 169.485 80.835 169.825 ;
        RECT 81.005 169.225 81.335 169.655 ;
        RECT 81.570 169.485 81.740 169.825 ;
        RECT 81.910 169.725 82.080 170.505 ;
        RECT 82.250 170.285 82.420 170.875 ;
        RECT 82.590 170.475 82.940 171.095 ;
        RECT 82.250 169.895 82.715 170.285 ;
        RECT 83.110 170.025 83.280 171.385 ;
        RECT 83.450 170.195 83.910 171.245 ;
        RECT 82.885 169.855 83.280 170.025 ;
        RECT 82.885 169.725 83.055 169.855 ;
        RECT 81.910 169.395 82.590 169.725 ;
        RECT 82.805 169.395 83.055 169.725 ;
        RECT 83.225 169.225 83.475 169.685 ;
        RECT 83.645 169.410 83.970 170.195 ;
        RECT 84.140 169.395 84.310 171.515 ;
        RECT 84.480 171.395 84.810 171.775 ;
        RECT 84.980 171.225 85.235 171.515 ;
        RECT 84.485 171.055 85.235 171.225 ;
        RECT 84.485 170.065 84.715 171.055 ;
        RECT 85.870 171.005 87.540 171.775 ;
        RECT 84.885 170.235 85.235 170.885 ;
        RECT 85.870 170.315 86.620 170.835 ;
        RECT 86.790 170.485 87.540 171.005 ;
        RECT 87.715 171.035 87.970 171.605 ;
        RECT 88.140 171.375 88.470 171.775 ;
        RECT 88.895 171.240 89.425 171.605 ;
        RECT 88.895 171.205 89.070 171.240 ;
        RECT 88.140 171.035 89.070 171.205 ;
        RECT 89.615 171.095 89.890 171.605 ;
        RECT 87.715 170.365 87.885 171.035 ;
        RECT 88.140 170.865 88.310 171.035 ;
        RECT 88.055 170.535 88.310 170.865 ;
        RECT 88.535 170.535 88.730 170.865 ;
        RECT 84.485 169.895 85.235 170.065 ;
        RECT 84.480 169.225 84.810 169.725 ;
        RECT 84.980 169.395 85.235 169.895 ;
        RECT 85.870 169.225 87.540 170.315 ;
        RECT 87.715 169.395 88.050 170.365 ;
        RECT 88.220 169.225 88.390 170.365 ;
        RECT 88.560 169.565 88.730 170.535 ;
        RECT 88.900 169.905 89.070 171.035 ;
        RECT 89.240 170.245 89.410 171.045 ;
        RECT 89.610 170.925 89.890 171.095 ;
        RECT 89.615 170.445 89.890 170.925 ;
        RECT 90.060 170.245 90.250 171.605 ;
        RECT 90.430 171.240 90.940 171.775 ;
        RECT 91.160 170.965 91.405 171.570 ;
        RECT 93.045 170.965 93.290 171.570 ;
        RECT 93.510 171.240 94.020 171.775 ;
        RECT 90.450 170.795 91.680 170.965 ;
        RECT 89.240 170.075 90.250 170.245 ;
        RECT 90.420 170.230 91.170 170.420 ;
        RECT 88.900 169.735 90.025 169.905 ;
        RECT 90.420 169.565 90.590 170.230 ;
        RECT 91.340 169.985 91.680 170.795 ;
        RECT 88.560 169.395 90.590 169.565 ;
        RECT 90.760 169.225 90.930 169.985 ;
        RECT 91.165 169.575 91.680 169.985 ;
        RECT 92.770 170.795 94.000 170.965 ;
        RECT 92.770 169.985 93.110 170.795 ;
        RECT 93.280 170.230 94.030 170.420 ;
        RECT 92.770 169.575 93.285 169.985 ;
        RECT 93.520 169.225 93.690 169.985 ;
        RECT 93.860 169.565 94.030 170.230 ;
        RECT 94.200 170.245 94.390 171.605 ;
        RECT 94.560 170.755 94.835 171.605 ;
        RECT 95.025 171.240 95.555 171.605 ;
        RECT 95.980 171.375 96.310 171.775 ;
        RECT 95.380 171.205 95.555 171.240 ;
        RECT 94.560 170.585 94.840 170.755 ;
        RECT 94.560 170.445 94.835 170.585 ;
        RECT 95.040 170.245 95.210 171.045 ;
        RECT 94.200 170.075 95.210 170.245 ;
        RECT 95.380 171.035 96.310 171.205 ;
        RECT 96.480 171.035 96.735 171.605 ;
        RECT 95.380 169.905 95.550 171.035 ;
        RECT 96.140 170.865 96.310 171.035 ;
        RECT 94.425 169.735 95.550 169.905 ;
        RECT 95.720 170.535 95.915 170.865 ;
        RECT 96.140 170.535 96.395 170.865 ;
        RECT 95.720 169.565 95.890 170.535 ;
        RECT 96.565 170.365 96.735 171.035 ;
        RECT 93.860 169.395 95.890 169.565 ;
        RECT 96.060 169.225 96.230 170.365 ;
        RECT 96.400 169.395 96.735 170.365 ;
        RECT 96.910 171.100 97.170 171.605 ;
        RECT 97.350 171.395 97.680 171.775 ;
        RECT 97.860 171.225 98.030 171.605 ;
        RECT 96.910 170.300 97.080 171.100 ;
        RECT 97.365 171.055 98.030 171.225 ;
        RECT 97.365 170.800 97.535 171.055 ;
        RECT 99.210 171.050 99.500 171.775 ;
        RECT 100.595 171.065 100.850 171.595 ;
        RECT 101.020 171.315 101.325 171.775 ;
        RECT 101.570 171.395 102.640 171.565 ;
        RECT 97.250 170.470 97.535 170.800 ;
        RECT 97.770 170.505 98.100 170.875 ;
        RECT 97.365 170.325 97.535 170.470 ;
        RECT 100.595 170.415 100.805 171.065 ;
        RECT 101.570 171.040 101.890 171.395 ;
        RECT 101.565 170.865 101.890 171.040 ;
        RECT 100.975 170.565 101.890 170.865 ;
        RECT 102.060 170.825 102.300 171.225 ;
        RECT 102.470 171.165 102.640 171.395 ;
        RECT 102.810 171.335 103.000 171.775 ;
        RECT 103.170 171.325 104.120 171.605 ;
        RECT 104.340 171.415 104.690 171.585 ;
        RECT 102.470 170.995 103.000 171.165 ;
        RECT 100.975 170.535 101.715 170.565 ;
        RECT 96.910 169.395 97.180 170.300 ;
        RECT 97.365 170.155 98.030 170.325 ;
        RECT 97.350 169.225 97.680 169.985 ;
        RECT 97.860 169.395 98.030 170.155 ;
        RECT 99.210 169.225 99.500 170.390 ;
        RECT 100.595 169.535 100.850 170.415 ;
        RECT 101.020 169.225 101.325 170.365 ;
        RECT 101.545 169.945 101.715 170.535 ;
        RECT 102.060 170.455 102.600 170.825 ;
        RECT 102.780 170.715 103.000 170.995 ;
        RECT 103.170 170.545 103.340 171.325 ;
        RECT 102.935 170.375 103.340 170.545 ;
        RECT 103.510 170.535 103.860 171.155 ;
        RECT 102.935 170.285 103.105 170.375 ;
        RECT 104.030 170.365 104.240 171.155 ;
        RECT 101.885 170.115 103.105 170.285 ;
        RECT 103.565 170.205 104.240 170.365 ;
        RECT 101.545 169.775 102.345 169.945 ;
        RECT 101.665 169.225 101.995 169.605 ;
        RECT 102.175 169.485 102.345 169.775 ;
        RECT 102.935 169.735 103.105 170.115 ;
        RECT 103.275 170.195 104.240 170.205 ;
        RECT 104.430 171.025 104.690 171.415 ;
        RECT 104.900 171.315 105.230 171.775 ;
        RECT 106.105 171.385 106.960 171.555 ;
        RECT 107.165 171.385 107.660 171.555 ;
        RECT 107.830 171.415 108.160 171.775 ;
        RECT 104.430 170.335 104.600 171.025 ;
        RECT 104.770 170.675 104.940 170.855 ;
        RECT 105.110 170.845 105.900 171.095 ;
        RECT 106.105 170.675 106.275 171.385 ;
        RECT 106.445 170.875 106.800 171.095 ;
        RECT 104.770 170.505 106.460 170.675 ;
        RECT 103.275 169.905 103.735 170.195 ;
        RECT 104.430 170.165 105.930 170.335 ;
        RECT 104.430 170.025 104.600 170.165 ;
        RECT 104.040 169.855 104.600 170.025 ;
        RECT 102.515 169.225 102.765 169.685 ;
        RECT 102.935 169.395 103.805 169.735 ;
        RECT 104.040 169.395 104.210 169.855 ;
        RECT 105.045 169.825 106.120 169.995 ;
        RECT 104.380 169.225 104.750 169.685 ;
        RECT 105.045 169.485 105.215 169.825 ;
        RECT 105.385 169.225 105.715 169.655 ;
        RECT 105.950 169.485 106.120 169.825 ;
        RECT 106.290 169.725 106.460 170.505 ;
        RECT 106.630 170.285 106.800 170.875 ;
        RECT 106.970 170.475 107.320 171.095 ;
        RECT 106.630 169.895 107.095 170.285 ;
        RECT 107.490 170.025 107.660 171.385 ;
        RECT 107.830 170.195 108.290 171.245 ;
        RECT 107.265 169.855 107.660 170.025 ;
        RECT 107.265 169.725 107.435 169.855 ;
        RECT 106.290 169.395 106.970 169.725 ;
        RECT 107.185 169.395 107.435 169.725 ;
        RECT 107.605 169.225 107.855 169.685 ;
        RECT 108.025 169.410 108.350 170.195 ;
        RECT 108.520 169.395 108.690 171.515 ;
        RECT 108.860 171.395 109.190 171.775 ;
        RECT 109.360 171.225 109.615 171.515 ;
        RECT 108.865 171.055 109.615 171.225 ;
        RECT 109.790 171.100 110.050 171.605 ;
        RECT 110.230 171.395 110.560 171.775 ;
        RECT 110.740 171.225 110.910 171.605 ;
        RECT 108.865 170.065 109.095 171.055 ;
        RECT 109.265 170.235 109.615 170.885 ;
        RECT 109.790 170.300 109.960 171.100 ;
        RECT 110.245 171.055 110.910 171.225 ;
        RECT 110.245 170.800 110.415 171.055 ;
        RECT 111.170 171.025 112.380 171.775 ;
        RECT 110.130 170.470 110.415 170.800 ;
        RECT 110.650 170.505 110.980 170.875 ;
        RECT 110.245 170.325 110.415 170.470 ;
        RECT 108.865 169.895 109.615 170.065 ;
        RECT 108.860 169.225 109.190 169.725 ;
        RECT 109.360 169.395 109.615 169.895 ;
        RECT 109.790 169.395 110.060 170.300 ;
        RECT 110.245 170.155 110.910 170.325 ;
        RECT 110.230 169.225 110.560 169.985 ;
        RECT 110.740 169.395 110.910 170.155 ;
        RECT 111.170 170.315 111.690 170.855 ;
        RECT 111.860 170.485 112.380 171.025 ;
        RECT 111.170 169.225 112.380 170.315 ;
        RECT 18.165 169.055 112.465 169.225 ;
        RECT 18.250 167.965 19.460 169.055 ;
        RECT 20.095 168.620 25.440 169.055 ;
        RECT 18.250 167.255 18.770 167.795 ;
        RECT 18.940 167.425 19.460 167.965 ;
        RECT 21.685 167.370 22.035 168.620 ;
        RECT 25.615 168.385 25.870 168.885 ;
        RECT 26.040 168.555 26.370 169.055 ;
        RECT 25.615 168.215 26.365 168.385 ;
        RECT 18.250 166.505 19.460 167.255 ;
        RECT 23.515 167.050 23.855 167.880 ;
        RECT 25.615 167.395 25.965 168.045 ;
        RECT 26.135 167.225 26.365 168.215 ;
        RECT 25.615 167.055 26.365 167.225 ;
        RECT 20.095 166.505 25.440 167.050 ;
        RECT 25.615 166.765 25.870 167.055 ;
        RECT 26.040 166.505 26.370 166.885 ;
        RECT 26.540 166.765 26.710 168.885 ;
        RECT 26.880 168.085 27.205 168.870 ;
        RECT 27.375 168.595 27.625 169.055 ;
        RECT 27.795 168.555 28.045 168.885 ;
        RECT 28.260 168.555 28.940 168.885 ;
        RECT 27.795 168.425 27.965 168.555 ;
        RECT 27.570 168.255 27.965 168.425 ;
        RECT 26.940 167.035 27.400 168.085 ;
        RECT 27.570 166.895 27.740 168.255 ;
        RECT 28.135 167.995 28.600 168.385 ;
        RECT 27.910 167.185 28.260 167.805 ;
        RECT 28.430 167.405 28.600 167.995 ;
        RECT 28.770 167.775 28.940 168.555 ;
        RECT 29.110 168.455 29.280 168.795 ;
        RECT 29.515 168.625 29.845 169.055 ;
        RECT 30.015 168.455 30.185 168.795 ;
        RECT 30.480 168.595 30.850 169.055 ;
        RECT 29.110 168.285 30.185 168.455 ;
        RECT 31.020 168.425 31.190 168.885 ;
        RECT 31.425 168.545 32.295 168.885 ;
        RECT 32.465 168.595 32.715 169.055 ;
        RECT 30.630 168.255 31.190 168.425 ;
        RECT 30.630 168.115 30.800 168.255 ;
        RECT 29.300 167.945 30.800 168.115 ;
        RECT 31.495 168.085 31.955 168.375 ;
        RECT 28.770 167.605 30.460 167.775 ;
        RECT 28.430 167.185 28.785 167.405 ;
        RECT 28.955 166.895 29.125 167.605 ;
        RECT 29.330 167.185 30.120 167.435 ;
        RECT 30.290 167.425 30.460 167.605 ;
        RECT 30.630 167.255 30.800 167.945 ;
        RECT 27.070 166.505 27.400 166.865 ;
        RECT 27.570 166.725 28.065 166.895 ;
        RECT 28.270 166.725 29.125 166.895 ;
        RECT 30.000 166.505 30.330 166.965 ;
        RECT 30.540 166.865 30.800 167.255 ;
        RECT 30.990 168.075 31.955 168.085 ;
        RECT 32.125 168.165 32.295 168.545 ;
        RECT 32.885 168.505 33.055 168.795 ;
        RECT 33.235 168.675 33.565 169.055 ;
        RECT 32.885 168.335 33.685 168.505 ;
        RECT 30.990 167.915 31.665 168.075 ;
        RECT 32.125 167.995 33.345 168.165 ;
        RECT 30.990 167.125 31.200 167.915 ;
        RECT 32.125 167.905 32.295 167.995 ;
        RECT 31.370 167.125 31.720 167.745 ;
        RECT 31.890 167.735 32.295 167.905 ;
        RECT 31.890 166.955 32.060 167.735 ;
        RECT 32.230 167.285 32.450 167.565 ;
        RECT 32.630 167.455 33.170 167.825 ;
        RECT 33.515 167.745 33.685 168.335 ;
        RECT 33.905 167.915 34.210 169.055 ;
        RECT 34.380 167.865 34.635 168.745 ;
        RECT 34.810 167.890 35.100 169.055 ;
        RECT 35.270 167.980 35.540 168.885 ;
        RECT 35.710 168.295 36.040 169.055 ;
        RECT 36.220 168.125 36.390 168.885 ;
        RECT 33.515 167.715 34.255 167.745 ;
        RECT 32.230 167.115 32.760 167.285 ;
        RECT 30.540 166.695 30.890 166.865 ;
        RECT 31.110 166.675 32.060 166.955 ;
        RECT 32.230 166.505 32.420 166.945 ;
        RECT 32.590 166.885 32.760 167.115 ;
        RECT 32.930 167.055 33.170 167.455 ;
        RECT 33.340 167.415 34.255 167.715 ;
        RECT 33.340 167.240 33.665 167.415 ;
        RECT 33.340 166.885 33.660 167.240 ;
        RECT 34.425 167.215 34.635 167.865 ;
        RECT 32.590 166.715 33.660 166.885 ;
        RECT 33.905 166.505 34.210 166.965 ;
        RECT 34.380 166.685 34.635 167.215 ;
        RECT 34.810 166.505 35.100 167.230 ;
        RECT 35.270 167.180 35.440 167.980 ;
        RECT 35.725 167.955 36.390 168.125 ;
        RECT 35.725 167.810 35.895 167.955 ;
        RECT 35.610 167.480 35.895 167.810 ;
        RECT 36.655 167.865 36.910 168.745 ;
        RECT 37.080 167.915 37.385 169.055 ;
        RECT 37.725 168.675 38.055 169.055 ;
        RECT 38.235 168.505 38.405 168.795 ;
        RECT 38.575 168.595 38.825 169.055 ;
        RECT 37.605 168.335 38.405 168.505 ;
        RECT 38.995 168.545 39.865 168.885 ;
        RECT 35.725 167.225 35.895 167.480 ;
        RECT 36.130 167.405 36.460 167.775 ;
        RECT 35.270 166.675 35.530 167.180 ;
        RECT 35.725 167.055 36.390 167.225 ;
        RECT 35.710 166.505 36.040 166.885 ;
        RECT 36.220 166.675 36.390 167.055 ;
        RECT 36.655 167.215 36.865 167.865 ;
        RECT 37.605 167.745 37.775 168.335 ;
        RECT 38.995 168.165 39.165 168.545 ;
        RECT 40.100 168.425 40.270 168.885 ;
        RECT 40.440 168.595 40.810 169.055 ;
        RECT 41.105 168.455 41.275 168.795 ;
        RECT 41.445 168.625 41.775 169.055 ;
        RECT 42.010 168.455 42.180 168.795 ;
        RECT 37.945 167.995 39.165 168.165 ;
        RECT 39.335 168.085 39.795 168.375 ;
        RECT 40.100 168.255 40.660 168.425 ;
        RECT 41.105 168.285 42.180 168.455 ;
        RECT 42.350 168.555 43.030 168.885 ;
        RECT 43.245 168.555 43.495 168.885 ;
        RECT 43.665 168.595 43.915 169.055 ;
        RECT 40.490 168.115 40.660 168.255 ;
        RECT 39.335 168.075 40.300 168.085 ;
        RECT 38.995 167.905 39.165 167.995 ;
        RECT 39.625 167.915 40.300 168.075 ;
        RECT 37.035 167.715 37.775 167.745 ;
        RECT 37.035 167.415 37.950 167.715 ;
        RECT 37.625 167.240 37.950 167.415 ;
        RECT 36.655 166.685 36.910 167.215 ;
        RECT 37.080 166.505 37.385 166.965 ;
        RECT 37.630 166.885 37.950 167.240 ;
        RECT 38.120 167.455 38.660 167.825 ;
        RECT 38.995 167.735 39.400 167.905 ;
        RECT 38.120 167.055 38.360 167.455 ;
        RECT 38.840 167.285 39.060 167.565 ;
        RECT 38.530 167.115 39.060 167.285 ;
        RECT 38.530 166.885 38.700 167.115 ;
        RECT 39.230 166.955 39.400 167.735 ;
        RECT 39.570 167.125 39.920 167.745 ;
        RECT 40.090 167.125 40.300 167.915 ;
        RECT 40.490 167.945 41.990 168.115 ;
        RECT 40.490 167.255 40.660 167.945 ;
        RECT 42.350 167.775 42.520 168.555 ;
        RECT 43.325 168.425 43.495 168.555 ;
        RECT 40.830 167.605 42.520 167.775 ;
        RECT 42.690 167.995 43.155 168.385 ;
        RECT 43.325 168.255 43.720 168.425 ;
        RECT 40.830 167.425 41.000 167.605 ;
        RECT 37.630 166.715 38.700 166.885 ;
        RECT 38.870 166.505 39.060 166.945 ;
        RECT 39.230 166.675 40.180 166.955 ;
        RECT 40.490 166.865 40.750 167.255 ;
        RECT 41.170 167.185 41.960 167.435 ;
        RECT 40.400 166.695 40.750 166.865 ;
        RECT 40.960 166.505 41.290 166.965 ;
        RECT 42.165 166.895 42.335 167.605 ;
        RECT 42.690 167.405 42.860 167.995 ;
        RECT 42.505 167.185 42.860 167.405 ;
        RECT 43.030 167.185 43.380 167.805 ;
        RECT 43.550 166.895 43.720 168.255 ;
        RECT 44.085 168.085 44.410 168.870 ;
        RECT 43.890 167.035 44.350 168.085 ;
        RECT 42.165 166.725 43.020 166.895 ;
        RECT 43.225 166.725 43.720 166.895 ;
        RECT 43.890 166.505 44.220 166.865 ;
        RECT 44.580 166.765 44.750 168.885 ;
        RECT 44.920 168.555 45.250 169.055 ;
        RECT 45.420 168.385 45.675 168.885 ;
        RECT 44.925 168.215 45.675 168.385 ;
        RECT 44.925 167.225 45.155 168.215 ;
        RECT 45.325 167.395 45.675 168.045 ;
        RECT 45.850 167.915 46.190 168.885 ;
        RECT 46.360 167.915 46.530 169.055 ;
        RECT 46.800 168.255 47.050 169.055 ;
        RECT 47.695 168.085 48.025 168.885 ;
        RECT 48.325 168.255 48.655 169.055 ;
        RECT 48.825 168.085 49.155 168.885 ;
        RECT 46.720 167.915 49.155 168.085 ;
        RECT 50.450 168.295 50.965 168.705 ;
        RECT 51.200 168.295 51.370 169.055 ;
        RECT 51.540 168.715 53.570 168.885 ;
        RECT 45.850 167.305 46.025 167.915 ;
        RECT 46.720 167.665 46.890 167.915 ;
        RECT 46.195 167.495 46.890 167.665 ;
        RECT 47.065 167.495 47.485 167.695 ;
        RECT 47.655 167.495 47.985 167.695 ;
        RECT 48.155 167.495 48.485 167.695 ;
        RECT 44.925 167.055 45.675 167.225 ;
        RECT 44.920 166.505 45.250 166.885 ;
        RECT 45.420 166.765 45.675 167.055 ;
        RECT 45.850 166.675 46.190 167.305 ;
        RECT 46.360 166.505 46.610 167.305 ;
        RECT 46.800 167.155 48.025 167.325 ;
        RECT 46.800 166.675 47.130 167.155 ;
        RECT 47.300 166.505 47.525 166.965 ;
        RECT 47.695 166.675 48.025 167.155 ;
        RECT 48.655 167.285 48.825 167.915 ;
        RECT 49.010 167.495 49.360 167.745 ;
        RECT 50.450 167.485 50.790 168.295 ;
        RECT 51.540 168.050 51.710 168.715 ;
        RECT 52.105 168.375 53.230 168.545 ;
        RECT 50.960 167.860 51.710 168.050 ;
        RECT 51.880 168.035 52.890 168.205 ;
        RECT 50.450 167.315 51.680 167.485 ;
        RECT 48.655 166.675 49.155 167.285 ;
        RECT 50.725 166.710 50.970 167.315 ;
        RECT 51.190 166.505 51.700 167.040 ;
        RECT 51.880 166.675 52.070 168.035 ;
        RECT 52.240 167.355 52.515 167.835 ;
        RECT 52.240 167.185 52.520 167.355 ;
        RECT 52.720 167.235 52.890 168.035 ;
        RECT 53.060 167.245 53.230 168.375 ;
        RECT 53.400 167.745 53.570 168.715 ;
        RECT 53.740 167.915 53.910 169.055 ;
        RECT 54.080 167.915 54.415 168.885 ;
        RECT 55.140 168.125 55.310 168.885 ;
        RECT 55.490 168.295 55.820 169.055 ;
        RECT 55.140 167.955 55.805 168.125 ;
        RECT 55.990 167.980 56.260 168.885 ;
        RECT 53.400 167.415 53.595 167.745 ;
        RECT 53.820 167.415 54.075 167.745 ;
        RECT 53.820 167.245 53.990 167.415 ;
        RECT 54.245 167.245 54.415 167.915 ;
        RECT 55.635 167.810 55.805 167.955 ;
        RECT 55.070 167.405 55.400 167.775 ;
        RECT 55.635 167.480 55.920 167.810 ;
        RECT 52.240 166.675 52.515 167.185 ;
        RECT 53.060 167.075 53.990 167.245 ;
        RECT 53.060 167.040 53.235 167.075 ;
        RECT 52.705 166.675 53.235 167.040 ;
        RECT 53.660 166.505 53.990 166.905 ;
        RECT 54.160 166.675 54.415 167.245 ;
        RECT 55.635 167.225 55.805 167.480 ;
        RECT 55.140 167.055 55.805 167.225 ;
        RECT 56.090 167.180 56.260 167.980 ;
        RECT 56.890 167.965 60.400 169.055 ;
        RECT 56.890 167.445 58.580 167.965 ;
        RECT 60.570 167.890 60.860 169.055 ;
        RECT 61.030 167.965 64.540 169.055 ;
        RECT 64.715 168.620 70.060 169.055 ;
        RECT 58.750 167.275 60.400 167.795 ;
        RECT 61.030 167.445 62.720 167.965 ;
        RECT 62.890 167.275 64.540 167.795 ;
        RECT 66.305 167.370 66.655 168.620 ;
        RECT 70.240 168.075 70.570 168.885 ;
        RECT 70.740 168.255 70.980 169.055 ;
        RECT 70.240 167.905 70.955 168.075 ;
        RECT 55.140 166.675 55.310 167.055 ;
        RECT 55.490 166.505 55.820 166.885 ;
        RECT 56.000 166.675 56.260 167.180 ;
        RECT 56.890 166.505 60.400 167.275 ;
        RECT 60.570 166.505 60.860 167.230 ;
        RECT 61.030 166.505 64.540 167.275 ;
        RECT 68.135 167.050 68.475 167.880 ;
        RECT 70.235 167.495 70.615 167.735 ;
        RECT 70.785 167.665 70.955 167.905 ;
        RECT 71.160 168.035 71.330 168.885 ;
        RECT 71.500 168.255 71.830 169.055 ;
        RECT 72.000 168.035 72.170 168.885 ;
        RECT 71.160 167.865 72.170 168.035 ;
        RECT 72.340 167.905 72.670 169.055 ;
        RECT 70.785 167.495 71.285 167.665 ;
        RECT 70.785 167.325 70.955 167.495 ;
        RECT 71.675 167.325 72.170 167.865 ;
        RECT 70.320 167.155 70.955 167.325 ;
        RECT 71.160 167.155 72.170 167.325 ;
        RECT 72.995 167.865 73.250 168.745 ;
        RECT 73.420 167.915 73.725 169.055 ;
        RECT 74.065 168.675 74.395 169.055 ;
        RECT 74.575 168.505 74.745 168.795 ;
        RECT 74.915 168.595 75.165 169.055 ;
        RECT 73.945 168.335 74.745 168.505 ;
        RECT 75.335 168.545 76.205 168.885 ;
        RECT 64.715 166.505 70.060 167.050 ;
        RECT 70.320 166.675 70.490 167.155 ;
        RECT 70.670 166.505 70.910 166.985 ;
        RECT 71.160 166.675 71.330 167.155 ;
        RECT 71.500 166.505 71.830 166.985 ;
        RECT 72.000 166.675 72.170 167.155 ;
        RECT 72.340 166.505 72.670 167.305 ;
        RECT 72.995 167.215 73.205 167.865 ;
        RECT 73.945 167.745 74.115 168.335 ;
        RECT 75.335 168.165 75.505 168.545 ;
        RECT 76.440 168.425 76.610 168.885 ;
        RECT 76.780 168.595 77.150 169.055 ;
        RECT 77.445 168.455 77.615 168.795 ;
        RECT 77.785 168.625 78.115 169.055 ;
        RECT 78.350 168.455 78.520 168.795 ;
        RECT 74.285 167.995 75.505 168.165 ;
        RECT 75.675 168.085 76.135 168.375 ;
        RECT 76.440 168.255 77.000 168.425 ;
        RECT 77.445 168.285 78.520 168.455 ;
        RECT 78.690 168.555 79.370 168.885 ;
        RECT 79.585 168.555 79.835 168.885 ;
        RECT 80.005 168.595 80.255 169.055 ;
        RECT 76.830 168.115 77.000 168.255 ;
        RECT 75.675 168.075 76.640 168.085 ;
        RECT 75.335 167.905 75.505 167.995 ;
        RECT 75.965 167.915 76.640 168.075 ;
        RECT 73.375 167.715 74.115 167.745 ;
        RECT 73.375 167.415 74.290 167.715 ;
        RECT 73.965 167.240 74.290 167.415 ;
        RECT 72.995 166.685 73.250 167.215 ;
        RECT 73.420 166.505 73.725 166.965 ;
        RECT 73.970 166.885 74.290 167.240 ;
        RECT 74.460 167.455 75.000 167.825 ;
        RECT 75.335 167.735 75.740 167.905 ;
        RECT 74.460 167.055 74.700 167.455 ;
        RECT 75.180 167.285 75.400 167.565 ;
        RECT 74.870 167.115 75.400 167.285 ;
        RECT 74.870 166.885 75.040 167.115 ;
        RECT 75.570 166.955 75.740 167.735 ;
        RECT 75.910 167.125 76.260 167.745 ;
        RECT 76.430 167.125 76.640 167.915 ;
        RECT 76.830 167.945 78.330 168.115 ;
        RECT 76.830 167.255 77.000 167.945 ;
        RECT 78.690 167.775 78.860 168.555 ;
        RECT 79.665 168.425 79.835 168.555 ;
        RECT 77.170 167.605 78.860 167.775 ;
        RECT 79.030 167.995 79.495 168.385 ;
        RECT 79.665 168.255 80.060 168.425 ;
        RECT 77.170 167.425 77.340 167.605 ;
        RECT 73.970 166.715 75.040 166.885 ;
        RECT 75.210 166.505 75.400 166.945 ;
        RECT 75.570 166.675 76.520 166.955 ;
        RECT 76.830 166.865 77.090 167.255 ;
        RECT 77.510 167.185 78.300 167.435 ;
        RECT 76.740 166.695 77.090 166.865 ;
        RECT 77.300 166.505 77.630 166.965 ;
        RECT 78.505 166.895 78.675 167.605 ;
        RECT 79.030 167.405 79.200 167.995 ;
        RECT 78.845 167.185 79.200 167.405 ;
        RECT 79.370 167.185 79.720 167.805 ;
        RECT 79.890 166.895 80.060 168.255 ;
        RECT 80.425 168.085 80.750 168.870 ;
        RECT 80.230 167.035 80.690 168.085 ;
        RECT 78.505 166.725 79.360 166.895 ;
        RECT 79.565 166.725 80.060 166.895 ;
        RECT 80.230 166.505 80.560 166.865 ;
        RECT 80.920 166.765 81.090 168.885 ;
        RECT 81.260 168.555 81.590 169.055 ;
        RECT 81.760 168.385 82.015 168.885 ;
        RECT 81.265 168.215 82.015 168.385 ;
        RECT 82.190 168.295 82.705 168.705 ;
        RECT 82.940 168.295 83.110 169.055 ;
        RECT 83.280 168.715 85.310 168.885 ;
        RECT 81.265 167.225 81.495 168.215 ;
        RECT 81.665 167.395 82.015 168.045 ;
        RECT 82.190 167.485 82.530 168.295 ;
        RECT 83.280 168.050 83.450 168.715 ;
        RECT 83.845 168.375 84.970 168.545 ;
        RECT 82.700 167.860 83.450 168.050 ;
        RECT 83.620 168.035 84.630 168.205 ;
        RECT 82.190 167.315 83.420 167.485 ;
        RECT 81.265 167.055 82.015 167.225 ;
        RECT 81.260 166.505 81.590 166.885 ;
        RECT 81.760 166.765 82.015 167.055 ;
        RECT 82.465 166.710 82.710 167.315 ;
        RECT 82.930 166.505 83.440 167.040 ;
        RECT 83.620 166.675 83.810 168.035 ;
        RECT 83.980 167.015 84.255 167.835 ;
        RECT 84.460 167.235 84.630 168.035 ;
        RECT 84.800 167.245 84.970 168.375 ;
        RECT 85.140 167.745 85.310 168.715 ;
        RECT 85.480 167.915 85.650 169.055 ;
        RECT 85.820 167.915 86.155 168.885 ;
        RECT 85.140 167.415 85.335 167.745 ;
        RECT 85.560 167.415 85.815 167.745 ;
        RECT 85.560 167.245 85.730 167.415 ;
        RECT 85.985 167.245 86.155 167.915 ;
        RECT 86.330 167.890 86.620 169.055 ;
        RECT 86.790 167.980 87.060 168.885 ;
        RECT 87.230 168.295 87.560 169.055 ;
        RECT 87.740 168.125 87.910 168.885 ;
        RECT 84.800 167.075 85.730 167.245 ;
        RECT 84.800 167.040 84.975 167.075 ;
        RECT 83.980 166.845 84.260 167.015 ;
        RECT 83.980 166.675 84.255 166.845 ;
        RECT 84.445 166.675 84.975 167.040 ;
        RECT 85.400 166.505 85.730 166.905 ;
        RECT 85.900 166.675 86.155 167.245 ;
        RECT 86.330 166.505 86.620 167.230 ;
        RECT 86.790 167.180 86.960 167.980 ;
        RECT 87.245 167.955 87.910 168.125 ;
        RECT 87.245 167.810 87.415 167.955 ;
        RECT 88.230 167.915 88.440 169.055 ;
        RECT 87.130 167.480 87.415 167.810 ;
        RECT 88.610 167.905 88.940 168.885 ;
        RECT 89.110 167.915 89.340 169.055 ;
        RECT 90.510 167.915 90.740 169.055 ;
        RECT 90.910 167.905 91.240 168.885 ;
        RECT 91.410 167.915 91.620 169.055 ;
        RECT 91.855 168.385 92.110 168.885 ;
        RECT 92.280 168.555 92.610 169.055 ;
        RECT 91.855 168.215 92.605 168.385 ;
        RECT 87.245 167.225 87.415 167.480 ;
        RECT 87.650 167.405 87.980 167.775 ;
        RECT 86.790 166.675 87.050 167.180 ;
        RECT 87.245 167.055 87.910 167.225 ;
        RECT 87.230 166.505 87.560 166.885 ;
        RECT 87.740 166.675 87.910 167.055 ;
        RECT 88.230 166.505 88.440 167.325 ;
        RECT 88.610 167.305 88.860 167.905 ;
        RECT 89.030 167.495 89.360 167.745 ;
        RECT 90.490 167.495 90.820 167.745 ;
        RECT 88.610 166.675 88.940 167.305 ;
        RECT 89.110 166.505 89.340 167.325 ;
        RECT 90.510 166.505 90.740 167.325 ;
        RECT 90.990 167.305 91.240 167.905 ;
        RECT 91.855 167.395 92.205 168.045 ;
        RECT 90.910 166.675 91.240 167.305 ;
        RECT 91.410 166.505 91.620 167.325 ;
        RECT 92.375 167.225 92.605 168.215 ;
        RECT 91.855 167.055 92.605 167.225 ;
        RECT 91.855 166.765 92.110 167.055 ;
        RECT 92.280 166.505 92.610 166.885 ;
        RECT 92.780 166.765 92.950 168.885 ;
        RECT 93.120 168.085 93.445 168.870 ;
        RECT 93.615 168.595 93.865 169.055 ;
        RECT 94.035 168.555 94.285 168.885 ;
        RECT 94.500 168.555 95.180 168.885 ;
        RECT 94.035 168.425 94.205 168.555 ;
        RECT 93.810 168.255 94.205 168.425 ;
        RECT 93.180 167.035 93.640 168.085 ;
        RECT 93.810 166.895 93.980 168.255 ;
        RECT 94.375 167.995 94.840 168.385 ;
        RECT 94.150 167.185 94.500 167.805 ;
        RECT 94.670 167.405 94.840 167.995 ;
        RECT 95.010 167.775 95.180 168.555 ;
        RECT 95.350 168.455 95.520 168.795 ;
        RECT 95.755 168.625 96.085 169.055 ;
        RECT 96.255 168.455 96.425 168.795 ;
        RECT 96.720 168.595 97.090 169.055 ;
        RECT 95.350 168.285 96.425 168.455 ;
        RECT 97.260 168.425 97.430 168.885 ;
        RECT 97.665 168.545 98.535 168.885 ;
        RECT 98.705 168.595 98.955 169.055 ;
        RECT 96.870 168.255 97.430 168.425 ;
        RECT 96.870 168.115 97.040 168.255 ;
        RECT 95.540 167.945 97.040 168.115 ;
        RECT 97.735 168.085 98.195 168.375 ;
        RECT 95.010 167.605 96.700 167.775 ;
        RECT 94.670 167.185 95.025 167.405 ;
        RECT 95.195 166.895 95.365 167.605 ;
        RECT 95.570 167.185 96.360 167.435 ;
        RECT 96.530 167.425 96.700 167.605 ;
        RECT 96.870 167.255 97.040 167.945 ;
        RECT 93.310 166.505 93.640 166.865 ;
        RECT 93.810 166.725 94.305 166.895 ;
        RECT 94.510 166.725 95.365 166.895 ;
        RECT 96.240 166.505 96.570 166.965 ;
        RECT 96.780 166.865 97.040 167.255 ;
        RECT 97.230 168.075 98.195 168.085 ;
        RECT 98.365 168.165 98.535 168.545 ;
        RECT 99.125 168.505 99.295 168.795 ;
        RECT 99.475 168.675 99.805 169.055 ;
        RECT 99.125 168.335 99.925 168.505 ;
        RECT 97.230 167.915 97.905 168.075 ;
        RECT 98.365 167.995 99.585 168.165 ;
        RECT 97.230 167.125 97.440 167.915 ;
        RECT 98.365 167.905 98.535 167.995 ;
        RECT 97.610 167.125 97.960 167.745 ;
        RECT 98.130 167.735 98.535 167.905 ;
        RECT 98.130 166.955 98.300 167.735 ;
        RECT 98.470 167.285 98.690 167.565 ;
        RECT 98.870 167.455 99.410 167.825 ;
        RECT 99.755 167.745 99.925 168.335 ;
        RECT 100.145 167.915 100.450 169.055 ;
        RECT 100.620 167.865 100.875 168.745 ;
        RECT 99.755 167.715 100.495 167.745 ;
        RECT 98.470 167.115 99.000 167.285 ;
        RECT 96.780 166.695 97.130 166.865 ;
        RECT 97.350 166.675 98.300 166.955 ;
        RECT 98.470 166.505 98.660 166.945 ;
        RECT 98.830 166.885 99.000 167.115 ;
        RECT 99.170 167.055 99.410 167.455 ;
        RECT 99.580 167.415 100.495 167.715 ;
        RECT 99.580 167.240 99.905 167.415 ;
        RECT 99.580 166.885 99.900 167.240 ;
        RECT 100.665 167.215 100.875 167.865 ;
        RECT 101.050 168.295 101.565 168.705 ;
        RECT 101.800 168.295 101.970 169.055 ;
        RECT 102.140 168.715 104.170 168.885 ;
        RECT 101.050 167.485 101.390 168.295 ;
        RECT 102.140 168.050 102.310 168.715 ;
        RECT 102.705 168.375 103.830 168.545 ;
        RECT 101.560 167.860 102.310 168.050 ;
        RECT 102.480 168.035 103.490 168.205 ;
        RECT 101.050 167.315 102.280 167.485 ;
        RECT 98.830 166.715 99.900 166.885 ;
        RECT 100.145 166.505 100.450 166.965 ;
        RECT 100.620 166.685 100.875 167.215 ;
        RECT 101.325 166.710 101.570 167.315 ;
        RECT 101.790 166.505 102.300 167.040 ;
        RECT 102.480 166.675 102.670 168.035 ;
        RECT 102.840 167.355 103.115 167.835 ;
        RECT 102.840 167.185 103.120 167.355 ;
        RECT 103.320 167.235 103.490 168.035 ;
        RECT 103.660 167.245 103.830 168.375 ;
        RECT 104.000 167.745 104.170 168.715 ;
        RECT 104.340 167.915 104.510 169.055 ;
        RECT 104.680 167.915 105.015 168.885 ;
        RECT 105.740 168.125 105.910 168.885 ;
        RECT 106.090 168.295 106.420 169.055 ;
        RECT 105.740 167.955 106.405 168.125 ;
        RECT 106.590 167.980 106.860 168.885 ;
        RECT 104.000 167.415 104.195 167.745 ;
        RECT 104.420 167.415 104.675 167.745 ;
        RECT 104.420 167.245 104.590 167.415 ;
        RECT 104.845 167.245 105.015 167.915 ;
        RECT 106.235 167.810 106.405 167.955 ;
        RECT 105.670 167.405 106.000 167.775 ;
        RECT 106.235 167.480 106.520 167.810 ;
        RECT 102.840 166.675 103.115 167.185 ;
        RECT 103.660 167.075 104.590 167.245 ;
        RECT 103.660 167.040 103.835 167.075 ;
        RECT 103.305 166.675 103.835 167.040 ;
        RECT 104.260 166.505 104.590 166.905 ;
        RECT 104.760 166.675 105.015 167.245 ;
        RECT 106.235 167.225 106.405 167.480 ;
        RECT 105.740 167.055 106.405 167.225 ;
        RECT 106.690 167.180 106.860 167.980 ;
        RECT 107.490 167.965 111.000 169.055 ;
        RECT 111.170 167.965 112.380 169.055 ;
        RECT 107.490 167.445 109.180 167.965 ;
        RECT 109.350 167.275 111.000 167.795 ;
        RECT 111.170 167.425 111.690 167.965 ;
        RECT 105.740 166.675 105.910 167.055 ;
        RECT 106.090 166.505 106.420 166.885 ;
        RECT 106.600 166.675 106.860 167.180 ;
        RECT 107.490 166.505 111.000 167.275 ;
        RECT 111.860 167.255 112.380 167.795 ;
        RECT 111.170 166.505 112.380 167.255 ;
        RECT 18.165 166.335 112.465 166.505 ;
        RECT 18.250 165.585 19.460 166.335 ;
        RECT 18.250 165.045 18.770 165.585 ;
        RECT 20.090 165.565 21.760 166.335 ;
        RECT 21.930 165.610 22.220 166.335 ;
        RECT 22.480 165.785 22.650 166.165 ;
        RECT 22.830 165.955 23.160 166.335 ;
        RECT 22.480 165.615 23.145 165.785 ;
        RECT 23.340 165.660 23.600 166.165 ;
        RECT 18.940 164.875 19.460 165.415 ;
        RECT 18.250 163.785 19.460 164.875 ;
        RECT 20.090 164.875 20.840 165.395 ;
        RECT 21.010 165.045 21.760 165.565 ;
        RECT 22.410 165.065 22.740 165.435 ;
        RECT 22.975 165.360 23.145 165.615 ;
        RECT 22.975 165.030 23.260 165.360 ;
        RECT 20.090 163.785 21.760 164.875 ;
        RECT 21.930 163.785 22.220 164.950 ;
        RECT 22.975 164.885 23.145 165.030 ;
        RECT 22.480 164.715 23.145 164.885 ;
        RECT 23.430 164.860 23.600 165.660 ;
        RECT 23.775 165.785 24.030 166.075 ;
        RECT 24.200 165.955 24.530 166.335 ;
        RECT 23.775 165.615 24.525 165.785 ;
        RECT 22.480 163.955 22.650 164.715 ;
        RECT 22.830 163.785 23.160 164.545 ;
        RECT 23.330 163.955 23.600 164.860 ;
        RECT 23.775 164.795 24.125 165.445 ;
        RECT 24.295 164.625 24.525 165.615 ;
        RECT 23.775 164.455 24.525 164.625 ;
        RECT 23.775 163.955 24.030 164.455 ;
        RECT 24.200 163.785 24.530 164.285 ;
        RECT 24.700 163.955 24.870 166.075 ;
        RECT 25.230 165.975 25.560 166.335 ;
        RECT 25.730 165.945 26.225 166.115 ;
        RECT 26.430 165.945 27.285 166.115 ;
        RECT 25.100 164.755 25.560 165.805 ;
        RECT 25.040 163.970 25.365 164.755 ;
        RECT 25.730 164.585 25.900 165.945 ;
        RECT 26.070 165.035 26.420 165.655 ;
        RECT 26.590 165.435 26.945 165.655 ;
        RECT 26.590 164.845 26.760 165.435 ;
        RECT 27.115 165.235 27.285 165.945 ;
        RECT 28.160 165.875 28.490 166.335 ;
        RECT 28.700 165.975 29.050 166.145 ;
        RECT 27.490 165.405 28.280 165.655 ;
        RECT 28.700 165.585 28.960 165.975 ;
        RECT 29.270 165.885 30.220 166.165 ;
        RECT 30.390 165.895 30.580 166.335 ;
        RECT 30.750 165.955 31.820 166.125 ;
        RECT 28.450 165.235 28.620 165.415 ;
        RECT 25.730 164.415 26.125 164.585 ;
        RECT 26.295 164.455 26.760 164.845 ;
        RECT 26.930 165.065 28.620 165.235 ;
        RECT 25.955 164.285 26.125 164.415 ;
        RECT 26.930 164.285 27.100 165.065 ;
        RECT 28.790 164.895 28.960 165.585 ;
        RECT 27.460 164.725 28.960 164.895 ;
        RECT 29.150 164.925 29.360 165.715 ;
        RECT 29.530 165.095 29.880 165.715 ;
        RECT 30.050 165.105 30.220 165.885 ;
        RECT 30.750 165.725 30.920 165.955 ;
        RECT 30.390 165.555 30.920 165.725 ;
        RECT 30.390 165.275 30.610 165.555 ;
        RECT 31.090 165.385 31.330 165.785 ;
        RECT 30.050 164.935 30.455 165.105 ;
        RECT 30.790 165.015 31.330 165.385 ;
        RECT 31.500 165.600 31.820 165.955 ;
        RECT 32.065 165.875 32.370 166.335 ;
        RECT 32.540 165.625 32.795 166.155 ;
        RECT 31.500 165.425 31.825 165.600 ;
        RECT 31.500 165.125 32.415 165.425 ;
        RECT 31.675 165.095 32.415 165.125 ;
        RECT 29.150 164.765 29.825 164.925 ;
        RECT 30.285 164.845 30.455 164.935 ;
        RECT 29.150 164.755 30.115 164.765 ;
        RECT 28.790 164.585 28.960 164.725 ;
        RECT 25.535 163.785 25.785 164.245 ;
        RECT 25.955 163.955 26.205 164.285 ;
        RECT 26.420 163.955 27.100 164.285 ;
        RECT 27.270 164.385 28.345 164.555 ;
        RECT 28.790 164.415 29.350 164.585 ;
        RECT 29.655 164.465 30.115 164.755 ;
        RECT 30.285 164.675 31.505 164.845 ;
        RECT 27.270 164.045 27.440 164.385 ;
        RECT 27.675 163.785 28.005 164.215 ;
        RECT 28.175 164.045 28.345 164.385 ;
        RECT 28.640 163.785 29.010 164.245 ;
        RECT 29.180 163.955 29.350 164.415 ;
        RECT 30.285 164.295 30.455 164.675 ;
        RECT 31.675 164.505 31.845 165.095 ;
        RECT 32.585 164.975 32.795 165.625 ;
        RECT 33.085 165.705 33.370 166.165 ;
        RECT 33.540 165.875 33.810 166.335 ;
        RECT 33.085 165.535 34.040 165.705 ;
        RECT 29.585 163.955 30.455 164.295 ;
        RECT 31.045 164.335 31.845 164.505 ;
        RECT 30.625 163.785 30.875 164.245 ;
        RECT 31.045 164.045 31.215 164.335 ;
        RECT 31.395 163.785 31.725 164.165 ;
        RECT 32.065 163.785 32.370 164.925 ;
        RECT 32.540 164.095 32.795 164.975 ;
        RECT 32.970 164.805 33.660 165.365 ;
        RECT 33.830 164.635 34.040 165.535 ;
        RECT 33.085 164.415 34.040 164.635 ;
        RECT 34.210 165.365 34.610 166.165 ;
        RECT 34.800 165.705 35.080 166.165 ;
        RECT 35.600 165.875 35.925 166.335 ;
        RECT 34.800 165.535 35.925 165.705 ;
        RECT 36.095 165.595 36.480 166.165 ;
        RECT 35.475 165.425 35.925 165.535 ;
        RECT 34.210 164.805 35.305 165.365 ;
        RECT 35.475 165.095 36.030 165.425 ;
        RECT 33.085 163.955 33.370 164.415 ;
        RECT 33.540 163.785 33.810 164.245 ;
        RECT 34.210 163.955 34.610 164.805 ;
        RECT 35.475 164.635 35.925 165.095 ;
        RECT 36.200 164.925 36.480 165.595 ;
        RECT 34.800 164.415 35.925 164.635 ;
        RECT 34.800 163.955 35.080 164.415 ;
        RECT 35.600 163.785 35.925 164.245 ;
        RECT 36.095 163.955 36.480 164.925 ;
        RECT 36.655 165.595 36.910 166.165 ;
        RECT 37.080 165.935 37.410 166.335 ;
        RECT 37.835 165.800 38.365 166.165 ;
        RECT 37.835 165.765 38.010 165.800 ;
        RECT 37.080 165.595 38.010 165.765 ;
        RECT 38.555 165.655 38.830 166.165 ;
        RECT 36.655 164.925 36.825 165.595 ;
        RECT 37.080 165.425 37.250 165.595 ;
        RECT 36.995 165.095 37.250 165.425 ;
        RECT 37.475 165.095 37.670 165.425 ;
        RECT 36.655 163.955 36.990 164.925 ;
        RECT 37.160 163.785 37.330 164.925 ;
        RECT 37.500 164.125 37.670 165.095 ;
        RECT 37.840 164.465 38.010 165.595 ;
        RECT 38.180 164.805 38.350 165.605 ;
        RECT 38.550 165.485 38.830 165.655 ;
        RECT 38.555 165.005 38.830 165.485 ;
        RECT 39.000 164.805 39.190 166.165 ;
        RECT 39.370 165.800 39.880 166.335 ;
        RECT 40.100 165.525 40.345 166.130 ;
        RECT 41.065 165.525 41.310 166.130 ;
        RECT 41.530 165.800 42.040 166.335 ;
        RECT 39.390 165.355 40.620 165.525 ;
        RECT 38.180 164.635 39.190 164.805 ;
        RECT 39.360 164.790 40.110 164.980 ;
        RECT 37.840 164.295 38.965 164.465 ;
        RECT 39.360 164.125 39.530 164.790 ;
        RECT 40.280 164.545 40.620 165.355 ;
        RECT 37.500 163.955 39.530 164.125 ;
        RECT 39.700 163.785 39.870 164.545 ;
        RECT 40.105 164.135 40.620 164.545 ;
        RECT 40.790 165.355 42.020 165.525 ;
        RECT 40.790 164.545 41.130 165.355 ;
        RECT 41.300 164.790 42.050 164.980 ;
        RECT 40.790 164.135 41.305 164.545 ;
        RECT 41.540 163.785 41.710 164.545 ;
        RECT 41.880 164.125 42.050 164.790 ;
        RECT 42.220 164.805 42.410 166.165 ;
        RECT 42.580 165.315 42.855 166.165 ;
        RECT 43.045 165.800 43.575 166.165 ;
        RECT 44.000 165.935 44.330 166.335 ;
        RECT 43.400 165.765 43.575 165.800 ;
        RECT 42.580 165.145 42.860 165.315 ;
        RECT 42.580 165.005 42.855 165.145 ;
        RECT 43.060 164.805 43.230 165.605 ;
        RECT 42.220 164.635 43.230 164.805 ;
        RECT 43.400 165.595 44.330 165.765 ;
        RECT 44.500 165.595 44.755 166.165 ;
        RECT 43.400 164.465 43.570 165.595 ;
        RECT 44.160 165.425 44.330 165.595 ;
        RECT 42.445 164.295 43.570 164.465 ;
        RECT 43.740 165.095 43.935 165.425 ;
        RECT 44.160 165.095 44.415 165.425 ;
        RECT 43.740 164.125 43.910 165.095 ;
        RECT 44.585 164.925 44.755 165.595 ;
        RECT 44.930 165.585 46.140 166.335 ;
        RECT 41.880 163.955 43.910 164.125 ;
        RECT 44.080 163.785 44.250 164.925 ;
        RECT 44.420 163.955 44.755 164.925 ;
        RECT 44.930 164.875 45.450 165.415 ;
        RECT 45.620 165.045 46.140 165.585 ;
        RECT 46.350 165.515 46.580 166.335 ;
        RECT 46.750 165.535 47.080 166.165 ;
        RECT 46.330 165.095 46.660 165.345 ;
        RECT 46.830 164.935 47.080 165.535 ;
        RECT 47.250 165.515 47.460 166.335 ;
        RECT 47.690 165.610 47.980 166.335 ;
        RECT 48.150 165.565 49.820 166.335 ;
        RECT 44.930 163.785 46.140 164.875 ;
        RECT 46.350 163.785 46.580 164.925 ;
        RECT 46.750 163.955 47.080 164.935 ;
        RECT 47.250 163.785 47.460 164.925 ;
        RECT 47.690 163.785 47.980 164.950 ;
        RECT 48.150 164.875 48.900 165.395 ;
        RECT 49.070 165.045 49.820 165.565 ;
        RECT 50.365 165.625 50.620 166.155 ;
        RECT 50.800 165.875 51.085 166.335 ;
        RECT 50.365 164.975 50.545 165.625 ;
        RECT 51.265 165.425 51.515 166.075 ;
        RECT 50.715 165.095 51.515 165.425 ;
        RECT 48.150 163.785 49.820 164.875 ;
        RECT 50.280 164.805 50.545 164.975 ;
        RECT 50.365 164.765 50.545 164.805 ;
        RECT 50.365 164.095 50.620 164.765 ;
        RECT 50.800 163.785 51.085 164.585 ;
        RECT 51.265 164.505 51.515 165.095 ;
        RECT 51.715 165.740 52.035 166.070 ;
        RECT 52.215 165.855 52.875 166.335 ;
        RECT 53.075 165.945 53.925 166.115 ;
        RECT 51.715 164.845 51.905 165.740 ;
        RECT 52.225 165.415 52.885 165.685 ;
        RECT 52.555 165.355 52.885 165.415 ;
        RECT 52.075 165.185 52.405 165.245 ;
        RECT 53.075 165.185 53.245 165.945 ;
        RECT 54.485 165.875 54.805 166.335 ;
        RECT 55.005 165.695 55.255 166.125 ;
        RECT 55.545 165.895 55.955 166.335 ;
        RECT 56.125 165.955 57.140 166.155 ;
        RECT 53.415 165.525 54.665 165.695 ;
        RECT 53.415 165.405 53.745 165.525 ;
        RECT 52.075 165.015 53.975 165.185 ;
        RECT 51.715 164.675 53.635 164.845 ;
        RECT 51.715 164.655 52.035 164.675 ;
        RECT 51.265 163.995 51.595 164.505 ;
        RECT 51.865 164.045 52.035 164.655 ;
        RECT 53.805 164.505 53.975 165.015 ;
        RECT 54.145 164.945 54.325 165.355 ;
        RECT 54.495 164.765 54.665 165.525 ;
        RECT 52.205 163.785 52.535 164.475 ;
        RECT 52.765 164.335 53.975 164.505 ;
        RECT 54.145 164.455 54.665 164.765 ;
        RECT 54.835 165.355 55.255 165.695 ;
        RECT 55.545 165.355 55.955 165.685 ;
        RECT 54.835 164.585 55.025 165.355 ;
        RECT 56.125 165.225 56.295 165.955 ;
        RECT 57.440 165.785 57.610 166.115 ;
        RECT 57.780 165.955 58.110 166.335 ;
        RECT 56.465 165.405 56.815 165.775 ;
        RECT 56.125 165.185 56.545 165.225 ;
        RECT 55.195 165.015 56.545 165.185 ;
        RECT 55.195 164.855 55.445 165.015 ;
        RECT 55.955 164.585 56.205 164.845 ;
        RECT 54.835 164.335 56.205 164.585 ;
        RECT 52.765 164.045 53.005 164.335 ;
        RECT 53.805 164.255 53.975 164.335 ;
        RECT 53.205 163.785 53.625 164.165 ;
        RECT 53.805 164.005 54.435 164.255 ;
        RECT 54.905 163.785 55.235 164.165 ;
        RECT 55.405 164.045 55.575 164.335 ;
        RECT 56.375 164.170 56.545 165.015 ;
        RECT 56.995 164.845 57.215 165.715 ;
        RECT 57.440 165.595 58.135 165.785 ;
        RECT 56.715 164.465 57.215 164.845 ;
        RECT 57.385 164.795 57.795 165.415 ;
        RECT 57.965 164.625 58.135 165.595 ;
        RECT 57.440 164.455 58.135 164.625 ;
        RECT 55.755 163.785 56.135 164.165 ;
        RECT 56.375 164.000 57.205 164.170 ;
        RECT 57.440 163.955 57.610 164.455 ;
        RECT 57.780 163.785 58.110 164.285 ;
        RECT 58.325 163.955 58.550 166.075 ;
        RECT 58.720 165.955 59.050 166.335 ;
        RECT 59.220 165.785 59.390 166.075 ;
        RECT 58.725 165.615 59.390 165.785 ;
        RECT 58.725 164.625 58.955 165.615 ;
        RECT 59.710 165.515 59.920 166.335 ;
        RECT 60.090 165.535 60.420 166.165 ;
        RECT 59.125 164.795 59.475 165.445 ;
        RECT 60.090 164.935 60.340 165.535 ;
        RECT 60.590 165.515 60.820 166.335 ;
        RECT 61.030 165.565 64.540 166.335 ;
        RECT 60.510 165.095 60.840 165.345 ;
        RECT 58.725 164.455 59.390 164.625 ;
        RECT 58.720 163.785 59.050 164.285 ;
        RECT 59.220 163.955 59.390 164.455 ;
        RECT 59.710 163.785 59.920 164.925 ;
        RECT 60.090 163.955 60.420 164.935 ;
        RECT 60.590 163.785 60.820 164.925 ;
        RECT 61.030 164.875 62.720 165.395 ;
        RECT 62.890 165.045 64.540 165.565 ;
        RECT 64.750 165.515 64.980 166.335 ;
        RECT 65.150 165.535 65.480 166.165 ;
        RECT 64.730 165.095 65.060 165.345 ;
        RECT 65.230 164.935 65.480 165.535 ;
        RECT 65.650 165.515 65.860 166.335 ;
        RECT 66.360 165.940 66.690 166.335 ;
        RECT 66.860 165.765 67.060 166.120 ;
        RECT 67.230 165.935 67.560 166.335 ;
        RECT 67.730 165.765 67.930 166.110 ;
        RECT 66.090 165.595 67.930 165.765 ;
        RECT 68.100 165.595 68.430 166.335 ;
        RECT 68.665 165.765 68.835 166.015 ;
        RECT 69.615 165.765 69.785 166.015 ;
        RECT 68.665 165.595 69.140 165.765 ;
        RECT 61.030 163.785 64.540 164.875 ;
        RECT 64.750 163.785 64.980 164.925 ;
        RECT 65.150 163.955 65.480 164.935 ;
        RECT 65.650 163.785 65.860 164.925 ;
        RECT 66.090 163.970 66.350 165.595 ;
        RECT 66.530 164.625 66.750 165.425 ;
        RECT 66.990 164.805 67.290 165.425 ;
        RECT 67.460 164.805 67.790 165.425 ;
        RECT 67.960 164.805 68.280 165.425 ;
        RECT 68.450 164.805 68.800 165.425 ;
        RECT 68.970 164.625 69.140 165.595 ;
        RECT 66.530 164.415 69.140 164.625 ;
        RECT 69.310 165.595 69.785 165.765 ;
        RECT 70.020 165.595 70.350 166.335 ;
        RECT 70.520 165.765 70.720 166.110 ;
        RECT 70.890 165.935 71.220 166.335 ;
        RECT 71.390 165.765 71.590 166.120 ;
        RECT 71.760 165.940 72.090 166.335 ;
        RECT 70.520 165.595 72.360 165.765 ;
        RECT 73.450 165.610 73.740 166.335 ;
        RECT 69.310 164.625 69.480 165.595 ;
        RECT 69.650 164.805 70.000 165.425 ;
        RECT 70.170 164.805 70.490 165.425 ;
        RECT 70.660 164.805 70.990 165.425 ;
        RECT 71.160 164.805 71.460 165.425 ;
        RECT 71.700 164.625 71.920 165.425 ;
        RECT 69.310 164.415 71.920 164.625 ;
        RECT 68.100 163.785 68.430 164.235 ;
        RECT 70.020 163.785 70.350 164.235 ;
        RECT 72.100 163.970 72.360 165.595 ;
        RECT 74.870 165.515 75.100 166.335 ;
        RECT 75.270 165.535 75.600 166.165 ;
        RECT 74.850 165.095 75.180 165.345 ;
        RECT 73.450 163.785 73.740 164.950 ;
        RECT 75.350 164.935 75.600 165.535 ;
        RECT 75.770 165.515 75.980 166.335 ;
        RECT 76.485 165.525 76.730 166.130 ;
        RECT 76.950 165.800 77.460 166.335 ;
        RECT 74.870 163.785 75.100 164.925 ;
        RECT 75.270 163.955 75.600 164.935 ;
        RECT 76.210 165.355 77.440 165.525 ;
        RECT 75.770 163.785 75.980 164.925 ;
        RECT 76.210 164.545 76.550 165.355 ;
        RECT 76.720 164.790 77.470 164.980 ;
        RECT 76.210 164.135 76.725 164.545 ;
        RECT 76.960 163.785 77.130 164.545 ;
        RECT 77.300 164.125 77.470 164.790 ;
        RECT 77.640 164.805 77.830 166.165 ;
        RECT 78.000 165.655 78.275 166.165 ;
        RECT 78.465 165.800 78.995 166.165 ;
        RECT 79.420 165.935 79.750 166.335 ;
        RECT 78.820 165.765 78.995 165.800 ;
        RECT 78.000 165.485 78.280 165.655 ;
        RECT 78.000 165.005 78.275 165.485 ;
        RECT 78.480 164.805 78.650 165.605 ;
        RECT 77.640 164.635 78.650 164.805 ;
        RECT 78.820 165.595 79.750 165.765 ;
        RECT 79.920 165.595 80.175 166.165 ;
        RECT 80.870 165.865 81.170 166.335 ;
        RECT 81.340 165.695 81.595 166.140 ;
        RECT 81.765 165.865 82.025 166.335 ;
        RECT 82.195 165.695 82.455 166.140 ;
        RECT 82.625 165.865 82.920 166.335 ;
        RECT 78.820 164.465 78.990 165.595 ;
        RECT 79.580 165.425 79.750 165.595 ;
        RECT 77.865 164.295 78.990 164.465 ;
        RECT 79.160 165.095 79.355 165.425 ;
        RECT 79.580 165.095 79.835 165.425 ;
        RECT 79.160 164.125 79.330 165.095 ;
        RECT 80.005 164.925 80.175 165.595 ;
        RECT 77.300 163.955 79.330 164.125 ;
        RECT 79.500 163.785 79.670 164.925 ;
        RECT 79.840 163.955 80.175 164.925 ;
        RECT 80.350 165.525 83.380 165.695 ;
        RECT 80.350 164.960 80.650 165.525 ;
        RECT 80.825 165.130 83.040 165.355 ;
        RECT 83.210 164.960 83.380 165.525 ;
        RECT 83.630 165.515 83.840 166.335 ;
        RECT 84.010 165.535 84.340 166.165 ;
        RECT 80.350 164.790 83.380 164.960 ;
        RECT 84.010 164.935 84.260 165.535 ;
        RECT 84.510 165.515 84.740 166.335 ;
        RECT 85.415 165.625 85.670 166.155 ;
        RECT 85.840 165.875 86.145 166.335 ;
        RECT 86.390 165.955 87.460 166.125 ;
        RECT 84.430 165.095 84.760 165.345 ;
        RECT 85.415 164.975 85.625 165.625 ;
        RECT 86.390 165.600 86.710 165.955 ;
        RECT 86.385 165.425 86.710 165.600 ;
        RECT 85.795 165.125 86.710 165.425 ;
        RECT 86.880 165.385 87.120 165.785 ;
        RECT 87.290 165.725 87.460 165.955 ;
        RECT 87.630 165.895 87.820 166.335 ;
        RECT 87.990 165.885 88.940 166.165 ;
        RECT 89.160 165.975 89.510 166.145 ;
        RECT 87.290 165.555 87.820 165.725 ;
        RECT 85.795 165.095 86.535 165.125 ;
        RECT 80.350 163.785 80.735 164.620 ;
        RECT 80.905 163.985 81.165 164.790 ;
        RECT 81.335 163.785 81.595 164.620 ;
        RECT 81.765 163.985 82.020 164.790 ;
        RECT 82.195 163.785 82.455 164.620 ;
        RECT 82.625 163.985 82.880 164.790 ;
        RECT 83.055 163.785 83.400 164.620 ;
        RECT 83.630 163.785 83.840 164.925 ;
        RECT 84.010 163.955 84.340 164.935 ;
        RECT 84.510 163.785 84.740 164.925 ;
        RECT 85.415 164.095 85.670 164.975 ;
        RECT 85.840 163.785 86.145 164.925 ;
        RECT 86.365 164.505 86.535 165.095 ;
        RECT 86.880 165.015 87.420 165.385 ;
        RECT 87.600 165.275 87.820 165.555 ;
        RECT 87.990 165.105 88.160 165.885 ;
        RECT 87.755 164.935 88.160 165.105 ;
        RECT 88.330 165.095 88.680 165.715 ;
        RECT 87.755 164.845 87.925 164.935 ;
        RECT 88.850 164.925 89.060 165.715 ;
        RECT 86.705 164.675 87.925 164.845 ;
        RECT 88.385 164.765 89.060 164.925 ;
        RECT 86.365 164.335 87.165 164.505 ;
        RECT 86.485 163.785 86.815 164.165 ;
        RECT 86.995 164.045 87.165 164.335 ;
        RECT 87.755 164.295 87.925 164.675 ;
        RECT 88.095 164.755 89.060 164.765 ;
        RECT 89.250 165.585 89.510 165.975 ;
        RECT 89.720 165.875 90.050 166.335 ;
        RECT 90.925 165.945 91.780 166.115 ;
        RECT 91.985 165.945 92.480 166.115 ;
        RECT 92.650 165.975 92.980 166.335 ;
        RECT 89.250 164.895 89.420 165.585 ;
        RECT 89.590 165.235 89.760 165.415 ;
        RECT 89.930 165.405 90.720 165.655 ;
        RECT 90.925 165.235 91.095 165.945 ;
        RECT 91.265 165.435 91.620 165.655 ;
        RECT 89.590 165.065 91.280 165.235 ;
        RECT 88.095 164.465 88.555 164.755 ;
        RECT 89.250 164.725 90.750 164.895 ;
        RECT 89.250 164.585 89.420 164.725 ;
        RECT 88.860 164.415 89.420 164.585 ;
        RECT 87.335 163.785 87.585 164.245 ;
        RECT 87.755 163.955 88.625 164.295 ;
        RECT 88.860 163.955 89.030 164.415 ;
        RECT 89.865 164.385 90.940 164.555 ;
        RECT 89.200 163.785 89.570 164.245 ;
        RECT 89.865 164.045 90.035 164.385 ;
        RECT 90.205 163.785 90.535 164.215 ;
        RECT 90.770 164.045 90.940 164.385 ;
        RECT 91.110 164.285 91.280 165.065 ;
        RECT 91.450 164.845 91.620 165.435 ;
        RECT 91.790 165.035 92.140 165.655 ;
        RECT 91.450 164.455 91.915 164.845 ;
        RECT 92.310 164.585 92.480 165.945 ;
        RECT 92.650 164.755 93.110 165.805 ;
        RECT 92.085 164.415 92.480 164.585 ;
        RECT 92.085 164.285 92.255 164.415 ;
        RECT 91.110 163.955 91.790 164.285 ;
        RECT 92.005 163.955 92.255 164.285 ;
        RECT 92.425 163.785 92.675 164.245 ;
        RECT 92.845 163.970 93.170 164.755 ;
        RECT 93.340 163.955 93.510 166.075 ;
        RECT 93.680 165.955 94.010 166.335 ;
        RECT 94.180 165.785 94.435 166.075 ;
        RECT 93.685 165.615 94.435 165.785 ;
        RECT 93.685 164.625 93.915 165.615 ;
        RECT 94.615 165.595 94.870 166.165 ;
        RECT 95.040 165.935 95.370 166.335 ;
        RECT 95.795 165.800 96.325 166.165 ;
        RECT 96.515 165.995 96.790 166.165 ;
        RECT 96.510 165.825 96.790 165.995 ;
        RECT 95.795 165.765 95.970 165.800 ;
        RECT 95.040 165.595 95.970 165.765 ;
        RECT 94.085 164.795 94.435 165.445 ;
        RECT 94.615 164.925 94.785 165.595 ;
        RECT 95.040 165.425 95.210 165.595 ;
        RECT 94.955 165.095 95.210 165.425 ;
        RECT 95.435 165.095 95.630 165.425 ;
        RECT 93.685 164.455 94.435 164.625 ;
        RECT 93.680 163.785 94.010 164.285 ;
        RECT 94.180 163.955 94.435 164.455 ;
        RECT 94.615 163.955 94.950 164.925 ;
        RECT 95.120 163.785 95.290 164.925 ;
        RECT 95.460 164.125 95.630 165.095 ;
        RECT 95.800 164.465 95.970 165.595 ;
        RECT 96.140 164.805 96.310 165.605 ;
        RECT 96.515 165.005 96.790 165.825 ;
        RECT 96.960 164.805 97.150 166.165 ;
        RECT 97.330 165.800 97.840 166.335 ;
        RECT 98.060 165.525 98.305 166.130 ;
        RECT 99.210 165.610 99.500 166.335 ;
        RECT 100.405 165.525 100.650 166.130 ;
        RECT 100.870 165.800 101.380 166.335 ;
        RECT 97.350 165.355 98.580 165.525 ;
        RECT 96.140 164.635 97.150 164.805 ;
        RECT 97.320 164.790 98.070 164.980 ;
        RECT 95.800 164.295 96.925 164.465 ;
        RECT 97.320 164.125 97.490 164.790 ;
        RECT 98.240 164.545 98.580 165.355 ;
        RECT 100.130 165.355 101.360 165.525 ;
        RECT 95.460 163.955 97.490 164.125 ;
        RECT 97.660 163.785 97.830 164.545 ;
        RECT 98.065 164.135 98.580 164.545 ;
        RECT 99.210 163.785 99.500 164.950 ;
        RECT 100.130 164.545 100.470 165.355 ;
        RECT 100.640 164.790 101.390 164.980 ;
        RECT 100.130 164.135 100.645 164.545 ;
        RECT 100.880 163.785 101.050 164.545 ;
        RECT 101.220 164.125 101.390 164.790 ;
        RECT 101.560 164.805 101.750 166.165 ;
        RECT 101.920 165.655 102.195 166.165 ;
        RECT 102.385 165.800 102.915 166.165 ;
        RECT 103.340 165.935 103.670 166.335 ;
        RECT 102.740 165.765 102.915 165.800 ;
        RECT 101.920 165.485 102.200 165.655 ;
        RECT 101.920 165.005 102.195 165.485 ;
        RECT 102.400 164.805 102.570 165.605 ;
        RECT 101.560 164.635 102.570 164.805 ;
        RECT 102.740 165.595 103.670 165.765 ;
        RECT 103.840 165.595 104.095 166.165 ;
        RECT 102.740 164.465 102.910 165.595 ;
        RECT 103.500 165.425 103.670 165.595 ;
        RECT 101.785 164.295 102.910 164.465 ;
        RECT 103.080 165.095 103.275 165.425 ;
        RECT 103.500 165.095 103.755 165.425 ;
        RECT 103.080 164.125 103.250 165.095 ;
        RECT 103.925 164.925 104.095 165.595 ;
        RECT 104.310 165.515 104.540 166.335 ;
        RECT 104.710 165.535 105.040 166.165 ;
        RECT 104.290 165.095 104.620 165.345 ;
        RECT 104.790 164.935 105.040 165.535 ;
        RECT 105.210 165.515 105.420 166.335 ;
        RECT 106.660 165.785 106.830 166.165 ;
        RECT 107.010 165.955 107.340 166.335 ;
        RECT 106.660 165.615 107.325 165.785 ;
        RECT 107.520 165.660 107.780 166.165 ;
        RECT 106.590 165.065 106.920 165.435 ;
        RECT 107.155 165.360 107.325 165.615 ;
        RECT 101.220 163.955 103.250 164.125 ;
        RECT 103.420 163.785 103.590 164.925 ;
        RECT 103.760 163.955 104.095 164.925 ;
        RECT 104.310 163.785 104.540 164.925 ;
        RECT 104.710 163.955 105.040 164.935 ;
        RECT 107.155 165.030 107.440 165.360 ;
        RECT 105.210 163.785 105.420 164.925 ;
        RECT 107.155 164.885 107.325 165.030 ;
        RECT 106.660 164.715 107.325 164.885 ;
        RECT 107.610 164.860 107.780 165.660 ;
        RECT 108.410 165.565 111.000 166.335 ;
        RECT 111.170 165.585 112.380 166.335 ;
        RECT 106.660 163.955 106.830 164.715 ;
        RECT 107.010 163.785 107.340 164.545 ;
        RECT 107.510 163.955 107.780 164.860 ;
        RECT 108.410 164.875 109.620 165.395 ;
        RECT 109.790 165.045 111.000 165.565 ;
        RECT 111.170 164.875 111.690 165.415 ;
        RECT 111.860 165.045 112.380 165.585 ;
        RECT 108.410 163.785 111.000 164.875 ;
        RECT 111.170 163.785 112.380 164.875 ;
        RECT 18.165 163.615 112.465 163.785 ;
        RECT 18.250 162.525 19.460 163.615 ;
        RECT 18.250 161.815 18.770 162.355 ;
        RECT 18.940 161.985 19.460 162.525 ;
        RECT 19.630 162.525 21.300 163.615 ;
        RECT 19.630 162.005 20.380 162.525 ;
        RECT 21.510 162.475 21.740 163.615 ;
        RECT 21.910 162.465 22.240 163.445 ;
        RECT 22.410 162.475 22.620 163.615 ;
        RECT 22.910 162.475 23.120 163.615 ;
        RECT 20.550 161.835 21.300 162.355 ;
        RECT 21.490 162.055 21.820 162.305 ;
        RECT 18.250 161.065 19.460 161.815 ;
        RECT 19.630 161.065 21.300 161.835 ;
        RECT 21.510 161.065 21.740 161.885 ;
        RECT 21.990 161.865 22.240 162.465 ;
        RECT 23.290 162.465 23.620 163.445 ;
        RECT 23.790 162.475 24.020 163.615 ;
        RECT 24.230 162.525 25.440 163.615 ;
        RECT 21.910 161.235 22.240 161.865 ;
        RECT 22.410 161.065 22.620 161.885 ;
        RECT 22.910 161.065 23.120 161.885 ;
        RECT 23.290 161.865 23.540 162.465 ;
        RECT 23.710 162.055 24.040 162.305 ;
        RECT 24.230 161.985 24.750 162.525 ;
        RECT 25.615 162.425 25.870 163.305 ;
        RECT 26.040 162.475 26.345 163.615 ;
        RECT 26.685 163.235 27.015 163.615 ;
        RECT 27.195 163.065 27.365 163.355 ;
        RECT 27.535 163.155 27.785 163.615 ;
        RECT 26.565 162.895 27.365 163.065 ;
        RECT 27.955 163.105 28.825 163.445 ;
        RECT 23.290 161.235 23.620 161.865 ;
        RECT 23.790 161.065 24.020 161.885 ;
        RECT 24.920 161.815 25.440 162.355 ;
        RECT 24.230 161.065 25.440 161.815 ;
        RECT 25.615 161.775 25.825 162.425 ;
        RECT 26.565 162.305 26.735 162.895 ;
        RECT 27.955 162.725 28.125 163.105 ;
        RECT 29.060 162.985 29.230 163.445 ;
        RECT 29.400 163.155 29.770 163.615 ;
        RECT 30.065 163.015 30.235 163.355 ;
        RECT 30.405 163.185 30.735 163.615 ;
        RECT 30.970 163.015 31.140 163.355 ;
        RECT 26.905 162.555 28.125 162.725 ;
        RECT 28.295 162.645 28.755 162.935 ;
        RECT 29.060 162.815 29.620 162.985 ;
        RECT 30.065 162.845 31.140 163.015 ;
        RECT 31.310 163.115 31.990 163.445 ;
        RECT 32.205 163.115 32.455 163.445 ;
        RECT 32.625 163.155 32.875 163.615 ;
        RECT 29.450 162.675 29.620 162.815 ;
        RECT 28.295 162.635 29.260 162.645 ;
        RECT 27.955 162.465 28.125 162.555 ;
        RECT 28.585 162.475 29.260 162.635 ;
        RECT 25.995 162.275 26.735 162.305 ;
        RECT 25.995 161.975 26.910 162.275 ;
        RECT 26.585 161.800 26.910 161.975 ;
        RECT 25.615 161.245 25.870 161.775 ;
        RECT 26.040 161.065 26.345 161.525 ;
        RECT 26.590 161.445 26.910 161.800 ;
        RECT 27.080 162.015 27.620 162.385 ;
        RECT 27.955 162.295 28.360 162.465 ;
        RECT 27.080 161.615 27.320 162.015 ;
        RECT 27.800 161.845 28.020 162.125 ;
        RECT 27.490 161.675 28.020 161.845 ;
        RECT 27.490 161.445 27.660 161.675 ;
        RECT 28.190 161.515 28.360 162.295 ;
        RECT 28.530 161.685 28.880 162.305 ;
        RECT 29.050 161.685 29.260 162.475 ;
        RECT 29.450 162.505 30.950 162.675 ;
        RECT 29.450 161.815 29.620 162.505 ;
        RECT 31.310 162.335 31.480 163.115 ;
        RECT 32.285 162.985 32.455 163.115 ;
        RECT 29.790 162.165 31.480 162.335 ;
        RECT 31.650 162.555 32.115 162.945 ;
        RECT 32.285 162.815 32.680 162.985 ;
        RECT 29.790 161.985 29.960 162.165 ;
        RECT 26.590 161.275 27.660 161.445 ;
        RECT 27.830 161.065 28.020 161.505 ;
        RECT 28.190 161.235 29.140 161.515 ;
        RECT 29.450 161.425 29.710 161.815 ;
        RECT 30.130 161.745 30.920 161.995 ;
        RECT 29.360 161.255 29.710 161.425 ;
        RECT 29.920 161.065 30.250 161.525 ;
        RECT 31.125 161.455 31.295 162.165 ;
        RECT 31.650 161.965 31.820 162.555 ;
        RECT 31.465 161.745 31.820 161.965 ;
        RECT 31.990 161.745 32.340 162.365 ;
        RECT 32.510 161.455 32.680 162.815 ;
        RECT 33.045 162.645 33.370 163.430 ;
        RECT 32.850 161.595 33.310 162.645 ;
        RECT 31.125 161.285 31.980 161.455 ;
        RECT 32.185 161.285 32.680 161.455 ;
        RECT 32.850 161.065 33.180 161.425 ;
        RECT 33.540 161.325 33.710 163.445 ;
        RECT 33.880 163.115 34.210 163.615 ;
        RECT 34.380 162.945 34.635 163.445 ;
        RECT 33.885 162.775 34.635 162.945 ;
        RECT 33.885 161.785 34.115 162.775 ;
        RECT 34.285 161.955 34.635 162.605 ;
        RECT 34.810 162.450 35.100 163.615 ;
        RECT 35.275 162.475 35.610 163.445 ;
        RECT 35.780 162.475 35.950 163.615 ;
        RECT 36.120 163.275 38.150 163.445 ;
        RECT 35.275 161.805 35.445 162.475 ;
        RECT 36.120 162.305 36.290 163.275 ;
        RECT 35.615 161.975 35.870 162.305 ;
        RECT 36.095 161.975 36.290 162.305 ;
        RECT 36.460 162.935 37.585 163.105 ;
        RECT 35.700 161.805 35.870 161.975 ;
        RECT 36.460 161.805 36.630 162.935 ;
        RECT 33.885 161.615 34.635 161.785 ;
        RECT 33.880 161.065 34.210 161.445 ;
        RECT 34.380 161.325 34.635 161.615 ;
        RECT 34.810 161.065 35.100 161.790 ;
        RECT 35.275 161.235 35.530 161.805 ;
        RECT 35.700 161.635 36.630 161.805 ;
        RECT 36.800 162.595 37.810 162.765 ;
        RECT 36.800 161.795 36.970 162.595 ;
        RECT 37.175 162.255 37.450 162.395 ;
        RECT 37.170 162.085 37.450 162.255 ;
        RECT 36.455 161.600 36.630 161.635 ;
        RECT 35.700 161.065 36.030 161.465 ;
        RECT 36.455 161.235 36.985 161.600 ;
        RECT 37.175 161.235 37.450 162.085 ;
        RECT 37.620 161.235 37.810 162.595 ;
        RECT 37.980 162.610 38.150 163.275 ;
        RECT 38.320 162.855 38.490 163.615 ;
        RECT 38.725 162.855 39.240 163.265 ;
        RECT 37.980 162.420 38.730 162.610 ;
        RECT 38.900 162.045 39.240 162.855 ;
        RECT 40.535 162.645 40.865 163.445 ;
        RECT 41.035 162.815 41.365 163.615 ;
        RECT 41.665 162.645 41.995 163.445 ;
        RECT 42.640 162.815 42.890 163.615 ;
        RECT 40.535 162.475 42.970 162.645 ;
        RECT 43.160 162.475 43.330 163.615 ;
        RECT 43.500 162.475 43.840 163.445 ;
        RECT 40.330 162.055 40.680 162.305 ;
        RECT 38.010 161.875 39.240 162.045 ;
        RECT 37.990 161.065 38.500 161.600 ;
        RECT 38.720 161.270 38.965 161.875 ;
        RECT 40.865 161.845 41.035 162.475 ;
        RECT 41.205 162.055 41.535 162.255 ;
        RECT 41.705 162.055 42.035 162.255 ;
        RECT 42.205 162.055 42.625 162.255 ;
        RECT 42.800 162.225 42.970 162.475 ;
        RECT 43.610 162.425 43.840 162.475 ;
        RECT 42.800 162.055 43.495 162.225 ;
        RECT 40.535 161.235 41.035 161.845 ;
        RECT 41.665 161.715 42.890 161.885 ;
        RECT 43.665 161.865 43.840 162.425 ;
        RECT 41.665 161.235 41.995 161.715 ;
        RECT 42.165 161.065 42.390 161.525 ;
        RECT 42.560 161.235 42.890 161.715 ;
        RECT 43.080 161.065 43.330 161.865 ;
        RECT 43.500 161.235 43.840 161.865 ;
        RECT 44.010 162.475 44.350 163.445 ;
        RECT 44.520 162.475 44.690 163.615 ;
        RECT 44.960 162.815 45.210 163.615 ;
        RECT 45.855 162.645 46.185 163.445 ;
        RECT 46.485 162.815 46.815 163.615 ;
        RECT 46.985 162.645 47.315 163.445 ;
        RECT 44.880 162.475 47.315 162.645 ;
        RECT 48.065 162.635 48.320 163.305 ;
        RECT 48.500 162.815 48.785 163.615 ;
        RECT 48.965 162.895 49.295 163.405 ;
        RECT 44.010 162.425 44.240 162.475 ;
        RECT 44.010 161.865 44.185 162.425 ;
        RECT 44.880 162.225 45.050 162.475 ;
        RECT 44.355 162.055 45.050 162.225 ;
        RECT 45.225 162.055 45.645 162.255 ;
        RECT 45.815 162.055 46.145 162.255 ;
        RECT 46.315 162.055 46.645 162.255 ;
        RECT 44.010 161.235 44.350 161.865 ;
        RECT 44.520 161.065 44.770 161.865 ;
        RECT 44.960 161.715 46.185 161.885 ;
        RECT 44.960 161.235 45.290 161.715 ;
        RECT 45.460 161.065 45.685 161.525 ;
        RECT 45.855 161.235 46.185 161.715 ;
        RECT 46.815 161.845 46.985 162.475 ;
        RECT 47.170 162.055 47.520 162.305 ;
        RECT 46.815 161.235 47.315 161.845 ;
        RECT 48.065 161.775 48.245 162.635 ;
        RECT 48.965 162.305 49.215 162.895 ;
        RECT 49.565 162.745 49.735 163.355 ;
        RECT 49.905 162.925 50.235 163.615 ;
        RECT 50.465 163.065 50.705 163.355 ;
        RECT 50.905 163.235 51.325 163.615 ;
        RECT 51.505 163.145 52.135 163.395 ;
        RECT 52.605 163.235 52.935 163.615 ;
        RECT 51.505 163.065 51.675 163.145 ;
        RECT 53.105 163.065 53.275 163.355 ;
        RECT 53.455 163.235 53.835 163.615 ;
        RECT 54.075 163.230 54.905 163.400 ;
        RECT 50.465 162.895 51.675 163.065 ;
        RECT 48.415 161.975 49.215 162.305 ;
        RECT 48.065 161.575 48.320 161.775 ;
        RECT 47.980 161.405 48.320 161.575 ;
        RECT 48.065 161.245 48.320 161.405 ;
        RECT 48.500 161.065 48.785 161.525 ;
        RECT 48.965 161.325 49.215 161.975 ;
        RECT 49.415 162.725 49.735 162.745 ;
        RECT 49.415 162.555 51.335 162.725 ;
        RECT 49.415 161.660 49.605 162.555 ;
        RECT 51.505 162.385 51.675 162.895 ;
        RECT 51.845 162.635 52.365 162.945 ;
        RECT 49.775 162.215 51.675 162.385 ;
        RECT 49.775 162.155 50.105 162.215 ;
        RECT 50.255 161.985 50.585 162.045 ;
        RECT 49.925 161.715 50.585 161.985 ;
        RECT 49.415 161.330 49.735 161.660 ;
        RECT 49.915 161.065 50.575 161.545 ;
        RECT 50.775 161.455 50.945 162.215 ;
        RECT 51.845 162.045 52.025 162.455 ;
        RECT 51.115 161.875 51.445 161.995 ;
        RECT 52.195 161.875 52.365 162.635 ;
        RECT 51.115 161.705 52.365 161.875 ;
        RECT 52.535 162.815 53.905 163.065 ;
        RECT 52.535 162.045 52.725 162.815 ;
        RECT 53.655 162.555 53.905 162.815 ;
        RECT 52.895 162.385 53.145 162.545 ;
        RECT 54.075 162.385 54.245 163.230 ;
        RECT 55.140 162.945 55.310 163.445 ;
        RECT 55.480 163.115 55.810 163.615 ;
        RECT 54.415 162.555 54.915 162.935 ;
        RECT 55.140 162.775 55.835 162.945 ;
        RECT 52.895 162.215 54.245 162.385 ;
        RECT 53.825 162.175 54.245 162.215 ;
        RECT 52.535 161.705 52.955 162.045 ;
        RECT 53.245 161.715 53.655 162.045 ;
        RECT 50.775 161.285 51.625 161.455 ;
        RECT 52.185 161.065 52.505 161.525 ;
        RECT 52.705 161.275 52.955 161.705 ;
        RECT 53.245 161.065 53.655 161.505 ;
        RECT 53.825 161.445 53.995 162.175 ;
        RECT 54.165 161.625 54.515 161.995 ;
        RECT 54.695 161.685 54.915 162.555 ;
        RECT 55.085 161.985 55.495 162.605 ;
        RECT 55.665 161.805 55.835 162.775 ;
        RECT 55.140 161.615 55.835 161.805 ;
        RECT 53.825 161.245 54.840 161.445 ;
        RECT 55.140 161.285 55.310 161.615 ;
        RECT 55.480 161.065 55.810 161.445 ;
        RECT 56.025 161.325 56.250 163.445 ;
        RECT 56.420 163.115 56.750 163.615 ;
        RECT 56.920 162.945 57.090 163.445 ;
        RECT 56.425 162.775 57.090 162.945 ;
        RECT 56.425 161.785 56.655 162.775 ;
        RECT 56.825 161.955 57.175 162.605 ;
        RECT 57.810 162.540 58.080 163.445 ;
        RECT 58.250 162.855 58.580 163.615 ;
        RECT 58.760 162.685 58.930 163.445 ;
        RECT 56.425 161.615 57.090 161.785 ;
        RECT 56.420 161.065 56.750 161.445 ;
        RECT 56.920 161.325 57.090 161.615 ;
        RECT 57.810 161.740 57.980 162.540 ;
        RECT 58.265 162.515 58.930 162.685 ;
        RECT 59.280 162.685 59.450 163.445 ;
        RECT 59.630 162.855 59.960 163.615 ;
        RECT 59.280 162.515 59.945 162.685 ;
        RECT 60.130 162.540 60.400 163.445 ;
        RECT 58.265 162.370 58.435 162.515 ;
        RECT 58.150 162.040 58.435 162.370 ;
        RECT 59.775 162.370 59.945 162.515 ;
        RECT 58.265 161.785 58.435 162.040 ;
        RECT 58.670 161.965 59.000 162.335 ;
        RECT 59.210 161.965 59.540 162.335 ;
        RECT 59.775 162.040 60.060 162.370 ;
        RECT 59.775 161.785 59.945 162.040 ;
        RECT 57.810 161.235 58.070 161.740 ;
        RECT 58.265 161.615 58.930 161.785 ;
        RECT 58.250 161.065 58.580 161.445 ;
        RECT 58.760 161.235 58.930 161.615 ;
        RECT 59.280 161.615 59.945 161.785 ;
        RECT 60.230 161.740 60.400 162.540 ;
        RECT 60.570 162.450 60.860 163.615 ;
        RECT 61.490 161.805 61.750 163.430 ;
        RECT 63.500 163.165 63.830 163.615 ;
        RECT 64.710 163.115 64.970 163.445 ;
        RECT 65.280 163.235 65.610 163.615 ;
        RECT 61.930 162.775 64.540 162.985 ;
        RECT 61.930 161.975 62.150 162.775 ;
        RECT 62.390 161.975 62.690 162.595 ;
        RECT 62.860 161.975 63.190 162.595 ;
        RECT 63.360 161.975 63.680 162.595 ;
        RECT 63.850 161.975 64.200 162.595 ;
        RECT 64.370 161.805 64.540 162.775 ;
        RECT 59.280 161.235 59.450 161.615 ;
        RECT 59.630 161.065 59.960 161.445 ;
        RECT 60.140 161.235 60.400 161.740 ;
        RECT 60.570 161.065 60.860 161.790 ;
        RECT 61.490 161.635 63.330 161.805 ;
        RECT 61.760 161.065 62.090 161.460 ;
        RECT 62.260 161.280 62.460 161.635 ;
        RECT 62.630 161.065 62.960 161.465 ;
        RECT 63.130 161.290 63.330 161.635 ;
        RECT 63.500 161.065 63.830 161.805 ;
        RECT 64.065 161.635 64.540 161.805 ;
        RECT 64.710 162.435 64.880 163.115 ;
        RECT 65.850 163.065 66.040 163.445 ;
        RECT 66.290 163.235 66.620 163.615 ;
        RECT 66.830 163.065 67.000 163.445 ;
        RECT 67.195 163.235 67.525 163.615 ;
        RECT 67.785 163.065 67.955 163.445 ;
        RECT 68.380 163.235 68.710 163.615 ;
        RECT 65.050 162.605 65.400 162.935 ;
        RECT 65.850 162.895 66.590 163.065 ;
        RECT 65.670 162.555 66.250 162.725 ;
        RECT 65.670 162.435 65.840 162.555 ;
        RECT 64.710 162.265 65.840 162.435 ;
        RECT 66.420 162.385 66.590 162.895 ;
        RECT 64.065 161.385 64.235 161.635 ;
        RECT 64.710 161.565 64.880 162.265 ;
        RECT 66.020 162.215 66.590 162.385 ;
        RECT 66.760 162.895 68.710 163.065 ;
        RECT 65.230 161.925 65.850 162.095 ;
        RECT 65.230 161.745 65.440 161.925 ;
        RECT 66.020 161.735 66.190 162.215 ;
        RECT 66.760 161.905 66.930 162.895 ;
        RECT 67.520 162.305 67.705 162.615 ;
        RECT 67.975 162.305 68.170 162.615 ;
        RECT 64.710 161.235 64.970 161.565 ;
        RECT 65.280 161.065 65.610 161.445 ;
        RECT 65.790 161.405 66.190 161.735 ;
        RECT 66.380 161.575 66.930 161.905 ;
        RECT 67.100 161.405 67.270 162.305 ;
        RECT 65.790 161.235 67.270 161.405 ;
        RECT 67.520 161.975 67.750 162.305 ;
        RECT 67.975 161.975 68.230 162.305 ;
        RECT 68.540 161.975 68.710 162.895 ;
        RECT 67.520 161.395 67.705 161.975 ;
        RECT 67.975 161.400 68.170 161.975 ;
        RECT 68.380 161.065 68.710 161.445 ;
        RECT 68.880 161.235 69.140 163.445 ;
        RECT 69.310 162.645 69.620 163.445 ;
        RECT 69.790 162.815 70.100 163.615 ;
        RECT 70.270 162.985 70.530 163.445 ;
        RECT 70.700 163.155 70.955 163.615 ;
        RECT 71.130 162.985 71.390 163.445 ;
        RECT 70.270 162.815 71.390 162.985 ;
        RECT 69.310 162.475 70.340 162.645 ;
        RECT 69.310 161.565 69.480 162.475 ;
        RECT 69.650 161.735 70.000 162.305 ;
        RECT 70.170 162.225 70.340 162.475 ;
        RECT 71.130 162.565 71.390 162.815 ;
        RECT 71.560 162.745 71.845 163.615 ;
        RECT 72.080 162.805 72.375 163.615 ;
        RECT 71.130 162.395 71.885 162.565 ;
        RECT 70.170 162.055 71.310 162.225 ;
        RECT 71.480 161.885 71.885 162.395 ;
        RECT 72.555 162.305 72.800 163.445 ;
        RECT 72.975 162.805 73.235 163.615 ;
        RECT 73.835 163.610 80.110 163.615 ;
        RECT 73.415 162.305 73.665 163.440 ;
        RECT 73.835 162.815 74.095 163.610 ;
        RECT 74.265 162.715 74.525 163.440 ;
        RECT 74.695 162.885 74.955 163.610 ;
        RECT 75.125 162.715 75.385 163.440 ;
        RECT 75.555 162.885 75.815 163.610 ;
        RECT 75.985 162.715 76.245 163.440 ;
        RECT 76.415 162.885 76.675 163.610 ;
        RECT 76.845 162.715 77.105 163.440 ;
        RECT 77.275 162.885 77.520 163.610 ;
        RECT 77.690 162.715 77.950 163.440 ;
        RECT 78.135 162.885 78.380 163.610 ;
        RECT 78.550 162.715 78.810 163.440 ;
        RECT 78.995 162.885 79.240 163.610 ;
        RECT 79.410 162.715 79.670 163.440 ;
        RECT 79.855 162.885 80.110 163.610 ;
        RECT 74.265 162.700 79.670 162.715 ;
        RECT 80.280 162.700 80.570 163.440 ;
        RECT 80.740 162.870 81.010 163.615 ;
        RECT 82.190 162.855 82.705 163.265 ;
        RECT 82.940 162.855 83.110 163.615 ;
        RECT 83.280 163.275 85.310 163.445 ;
        RECT 74.265 162.475 81.010 162.700 ;
        RECT 70.235 161.715 71.885 161.885 ;
        RECT 72.070 161.745 72.385 162.305 ;
        RECT 72.555 162.055 79.675 162.305 ;
        RECT 69.310 161.235 69.610 161.565 ;
        RECT 69.780 161.065 70.055 161.545 ;
        RECT 70.235 161.325 70.530 161.715 ;
        RECT 70.700 161.065 70.955 161.545 ;
        RECT 71.130 161.325 71.390 161.715 ;
        RECT 71.560 161.065 71.840 161.545 ;
        RECT 72.070 161.065 72.375 161.575 ;
        RECT 72.555 161.245 72.805 162.055 ;
        RECT 72.975 161.065 73.235 161.590 ;
        RECT 73.415 161.245 73.665 162.055 ;
        RECT 79.845 161.885 81.010 162.475 ;
        RECT 74.265 161.715 81.010 161.885 ;
        RECT 82.190 162.045 82.530 162.855 ;
        RECT 83.280 162.610 83.450 163.275 ;
        RECT 83.845 162.935 84.970 163.105 ;
        RECT 82.700 162.420 83.450 162.610 ;
        RECT 83.620 162.595 84.630 162.765 ;
        RECT 82.190 161.875 83.420 162.045 ;
        RECT 73.835 161.065 74.095 161.625 ;
        RECT 74.265 161.260 74.525 161.715 ;
        RECT 74.695 161.065 74.955 161.545 ;
        RECT 75.125 161.260 75.385 161.715 ;
        RECT 75.555 161.065 75.815 161.545 ;
        RECT 75.985 161.260 76.245 161.715 ;
        RECT 76.415 161.065 76.660 161.545 ;
        RECT 76.830 161.260 77.105 161.715 ;
        RECT 77.275 161.065 77.520 161.545 ;
        RECT 77.690 161.260 77.950 161.715 ;
        RECT 78.130 161.065 78.380 161.545 ;
        RECT 78.550 161.260 78.810 161.715 ;
        RECT 78.990 161.065 79.240 161.545 ;
        RECT 79.410 161.260 79.670 161.715 ;
        RECT 79.850 161.065 80.110 161.545 ;
        RECT 80.280 161.260 80.540 161.715 ;
        RECT 80.710 161.065 81.010 161.545 ;
        RECT 82.465 161.270 82.710 161.875 ;
        RECT 82.930 161.065 83.440 161.600 ;
        RECT 83.620 161.235 83.810 162.595 ;
        RECT 83.980 161.575 84.255 162.395 ;
        RECT 84.460 161.795 84.630 162.595 ;
        RECT 84.800 161.805 84.970 162.935 ;
        RECT 85.140 162.305 85.310 163.275 ;
        RECT 85.480 162.475 85.650 163.615 ;
        RECT 85.820 162.475 86.155 163.445 ;
        RECT 85.140 161.975 85.335 162.305 ;
        RECT 85.560 161.975 85.815 162.305 ;
        RECT 85.560 161.805 85.730 161.975 ;
        RECT 85.985 161.805 86.155 162.475 ;
        RECT 86.330 162.450 86.620 163.615 ;
        RECT 86.850 162.475 87.060 163.615 ;
        RECT 87.230 162.465 87.560 163.445 ;
        RECT 87.730 162.475 87.960 163.615 ;
        RECT 89.150 162.780 89.405 163.615 ;
        RECT 89.575 162.610 89.835 163.415 ;
        RECT 90.005 162.780 90.265 163.615 ;
        RECT 90.435 162.610 90.690 163.415 ;
        RECT 84.800 161.635 85.730 161.805 ;
        RECT 84.800 161.600 84.975 161.635 ;
        RECT 83.980 161.405 84.260 161.575 ;
        RECT 83.980 161.235 84.255 161.405 ;
        RECT 84.445 161.235 84.975 161.600 ;
        RECT 85.400 161.065 85.730 161.465 ;
        RECT 85.900 161.235 86.155 161.805 ;
        RECT 86.330 161.065 86.620 161.790 ;
        RECT 86.850 161.065 87.060 161.885 ;
        RECT 87.230 161.865 87.480 162.465 ;
        RECT 89.090 162.440 90.690 162.610 ;
        RECT 91.020 162.685 91.190 163.445 ;
        RECT 91.370 162.855 91.700 163.615 ;
        RECT 91.020 162.515 91.685 162.685 ;
        RECT 91.870 162.540 92.140 163.445 ;
        RECT 87.650 162.055 87.980 162.305 ;
        RECT 87.230 161.235 87.560 161.865 ;
        RECT 87.730 161.065 87.960 161.885 ;
        RECT 89.090 161.875 89.370 162.440 ;
        RECT 91.515 162.370 91.685 162.515 ;
        RECT 89.540 162.045 90.760 162.270 ;
        RECT 90.950 161.965 91.280 162.335 ;
        RECT 91.515 162.040 91.800 162.370 ;
        RECT 89.090 161.705 89.820 161.875 ;
        RECT 91.515 161.785 91.685 162.040 ;
        RECT 89.095 161.065 89.425 161.535 ;
        RECT 89.595 161.260 89.820 161.705 ;
        RECT 91.020 161.615 91.685 161.785 ;
        RECT 91.970 161.740 92.140 162.540 ;
        RECT 92.770 162.525 95.360 163.615 ;
        RECT 95.530 162.540 95.800 163.445 ;
        RECT 95.970 162.855 96.300 163.615 ;
        RECT 96.480 162.685 96.650 163.445 ;
        RECT 92.770 162.005 93.980 162.525 ;
        RECT 94.150 161.835 95.360 162.355 ;
        RECT 89.990 161.065 90.285 161.590 ;
        RECT 91.020 161.235 91.190 161.615 ;
        RECT 91.370 161.065 91.700 161.445 ;
        RECT 91.880 161.235 92.140 161.740 ;
        RECT 92.770 161.065 95.360 161.835 ;
        RECT 95.530 161.740 95.700 162.540 ;
        RECT 95.985 162.515 96.650 162.685 ;
        RECT 96.910 162.855 97.425 163.265 ;
        RECT 97.660 162.855 97.830 163.615 ;
        RECT 98.000 163.275 100.030 163.445 ;
        RECT 95.985 162.370 96.155 162.515 ;
        RECT 95.870 162.040 96.155 162.370 ;
        RECT 95.985 161.785 96.155 162.040 ;
        RECT 96.390 161.965 96.720 162.335 ;
        RECT 96.910 162.045 97.250 162.855 ;
        RECT 98.000 162.610 98.170 163.275 ;
        RECT 98.565 162.935 99.690 163.105 ;
        RECT 97.420 162.420 98.170 162.610 ;
        RECT 98.340 162.595 99.350 162.765 ;
        RECT 96.910 161.875 98.140 162.045 ;
        RECT 95.530 161.235 95.790 161.740 ;
        RECT 95.985 161.615 96.650 161.785 ;
        RECT 95.970 161.065 96.300 161.445 ;
        RECT 96.480 161.235 96.650 161.615 ;
        RECT 97.185 161.270 97.430 161.875 ;
        RECT 97.650 161.065 98.160 161.600 ;
        RECT 98.340 161.235 98.530 162.595 ;
        RECT 98.700 161.915 98.975 162.395 ;
        RECT 98.700 161.745 98.980 161.915 ;
        RECT 99.180 161.795 99.350 162.595 ;
        RECT 99.520 161.805 99.690 162.935 ;
        RECT 99.860 162.305 100.030 163.275 ;
        RECT 100.200 162.475 100.370 163.615 ;
        RECT 100.540 162.475 100.875 163.445 ;
        RECT 99.860 161.975 100.055 162.305 ;
        RECT 100.280 161.975 100.535 162.305 ;
        RECT 100.280 161.805 100.450 161.975 ;
        RECT 100.705 161.805 100.875 162.475 ;
        RECT 98.700 161.235 98.975 161.745 ;
        RECT 99.520 161.635 100.450 161.805 ;
        RECT 99.520 161.600 99.695 161.635 ;
        RECT 99.165 161.235 99.695 161.600 ;
        RECT 100.120 161.065 100.450 161.465 ;
        RECT 100.620 161.235 100.875 161.805 ;
        RECT 101.055 162.425 101.310 163.305 ;
        RECT 101.480 162.475 101.785 163.615 ;
        RECT 102.125 163.235 102.455 163.615 ;
        RECT 102.635 163.065 102.805 163.355 ;
        RECT 102.975 163.155 103.225 163.615 ;
        RECT 102.005 162.895 102.805 163.065 ;
        RECT 103.395 163.105 104.265 163.445 ;
        RECT 101.055 161.775 101.265 162.425 ;
        RECT 102.005 162.305 102.175 162.895 ;
        RECT 103.395 162.725 103.565 163.105 ;
        RECT 104.500 162.985 104.670 163.445 ;
        RECT 104.840 163.155 105.210 163.615 ;
        RECT 105.505 163.015 105.675 163.355 ;
        RECT 105.845 163.185 106.175 163.615 ;
        RECT 106.410 163.015 106.580 163.355 ;
        RECT 102.345 162.555 103.565 162.725 ;
        RECT 103.735 162.645 104.195 162.935 ;
        RECT 104.500 162.815 105.060 162.985 ;
        RECT 105.505 162.845 106.580 163.015 ;
        RECT 106.750 163.115 107.430 163.445 ;
        RECT 107.645 163.115 107.895 163.445 ;
        RECT 108.065 163.155 108.315 163.615 ;
        RECT 104.890 162.675 105.060 162.815 ;
        RECT 103.735 162.635 104.700 162.645 ;
        RECT 103.395 162.465 103.565 162.555 ;
        RECT 104.025 162.475 104.700 162.635 ;
        RECT 101.435 162.275 102.175 162.305 ;
        RECT 101.435 161.975 102.350 162.275 ;
        RECT 102.025 161.800 102.350 161.975 ;
        RECT 101.055 161.245 101.310 161.775 ;
        RECT 101.480 161.065 101.785 161.525 ;
        RECT 102.030 161.445 102.350 161.800 ;
        RECT 102.520 162.015 103.060 162.385 ;
        RECT 103.395 162.295 103.800 162.465 ;
        RECT 102.520 161.615 102.760 162.015 ;
        RECT 103.240 161.845 103.460 162.125 ;
        RECT 102.930 161.675 103.460 161.845 ;
        RECT 102.930 161.445 103.100 161.675 ;
        RECT 103.630 161.515 103.800 162.295 ;
        RECT 103.970 161.685 104.320 162.305 ;
        RECT 104.490 161.685 104.700 162.475 ;
        RECT 104.890 162.505 106.390 162.675 ;
        RECT 104.890 161.815 105.060 162.505 ;
        RECT 106.750 162.335 106.920 163.115 ;
        RECT 107.725 162.985 107.895 163.115 ;
        RECT 105.230 162.165 106.920 162.335 ;
        RECT 107.090 162.555 107.555 162.945 ;
        RECT 107.725 162.815 108.120 162.985 ;
        RECT 105.230 161.985 105.400 162.165 ;
        RECT 102.030 161.275 103.100 161.445 ;
        RECT 103.270 161.065 103.460 161.505 ;
        RECT 103.630 161.235 104.580 161.515 ;
        RECT 104.890 161.425 105.150 161.815 ;
        RECT 105.570 161.745 106.360 161.995 ;
        RECT 104.800 161.255 105.150 161.425 ;
        RECT 105.360 161.065 105.690 161.525 ;
        RECT 106.565 161.455 106.735 162.165 ;
        RECT 107.090 161.965 107.260 162.555 ;
        RECT 106.905 161.745 107.260 161.965 ;
        RECT 107.430 161.745 107.780 162.365 ;
        RECT 107.950 161.455 108.120 162.815 ;
        RECT 108.485 162.645 108.810 163.430 ;
        RECT 108.290 161.595 108.750 162.645 ;
        RECT 106.565 161.285 107.420 161.455 ;
        RECT 107.625 161.285 108.120 161.455 ;
        RECT 108.290 161.065 108.620 161.425 ;
        RECT 108.980 161.325 109.150 163.445 ;
        RECT 109.320 163.115 109.650 163.615 ;
        RECT 109.820 162.945 110.075 163.445 ;
        RECT 109.325 162.775 110.075 162.945 ;
        RECT 109.325 161.785 109.555 162.775 ;
        RECT 109.725 161.955 110.075 162.605 ;
        RECT 111.170 162.525 112.380 163.615 ;
        RECT 111.170 161.985 111.690 162.525 ;
        RECT 111.860 161.815 112.380 162.355 ;
        RECT 109.325 161.615 110.075 161.785 ;
        RECT 109.320 161.065 109.650 161.445 ;
        RECT 109.820 161.325 110.075 161.615 ;
        RECT 111.170 161.065 112.380 161.815 ;
        RECT 18.165 160.895 112.465 161.065 ;
        RECT 18.250 160.145 19.460 160.895 ;
        RECT 20.640 160.345 20.810 160.725 ;
        RECT 20.990 160.515 21.320 160.895 ;
        RECT 20.640 160.175 21.305 160.345 ;
        RECT 21.500 160.220 21.760 160.725 ;
        RECT 18.250 159.605 18.770 160.145 ;
        RECT 18.940 159.435 19.460 159.975 ;
        RECT 20.570 159.625 20.900 159.995 ;
        RECT 21.135 159.920 21.305 160.175 ;
        RECT 21.135 159.590 21.420 159.920 ;
        RECT 21.135 159.445 21.305 159.590 ;
        RECT 18.250 158.345 19.460 159.435 ;
        RECT 20.640 159.275 21.305 159.445 ;
        RECT 21.590 159.420 21.760 160.220 ;
        RECT 21.930 160.170 22.220 160.895 ;
        RECT 23.000 160.095 23.330 160.895 ;
        RECT 23.500 160.245 23.670 160.725 ;
        RECT 23.840 160.415 24.170 160.895 ;
        RECT 24.340 160.245 24.510 160.725 ;
        RECT 24.760 160.415 25.000 160.895 ;
        RECT 25.180 160.245 25.350 160.725 ;
        RECT 23.500 160.075 24.510 160.245 ;
        RECT 24.715 160.075 25.350 160.245 ;
        RECT 25.615 160.155 25.870 160.725 ;
        RECT 26.040 160.495 26.370 160.895 ;
        RECT 26.795 160.360 27.325 160.725 ;
        RECT 26.795 160.325 26.970 160.360 ;
        RECT 26.040 160.155 26.970 160.325 ;
        RECT 23.500 160.045 24.000 160.075 ;
        RECT 23.500 159.535 23.995 160.045 ;
        RECT 24.715 159.905 24.885 160.075 ;
        RECT 24.385 159.735 24.885 159.905 ;
        RECT 20.640 158.515 20.810 159.275 ;
        RECT 20.990 158.345 21.320 159.105 ;
        RECT 21.490 158.515 21.760 159.420 ;
        RECT 21.930 158.345 22.220 159.510 ;
        RECT 23.000 158.345 23.330 159.495 ;
        RECT 23.500 159.365 24.510 159.535 ;
        RECT 23.500 158.515 23.670 159.365 ;
        RECT 23.840 158.345 24.170 159.145 ;
        RECT 24.340 158.515 24.510 159.365 ;
        RECT 24.715 159.495 24.885 159.735 ;
        RECT 25.055 159.665 25.435 159.905 ;
        RECT 24.715 159.325 25.430 159.495 ;
        RECT 24.690 158.345 24.930 159.145 ;
        RECT 25.100 158.515 25.430 159.325 ;
        RECT 25.615 159.485 25.785 160.155 ;
        RECT 26.040 159.985 26.210 160.155 ;
        RECT 25.955 159.655 26.210 159.985 ;
        RECT 26.435 159.655 26.630 159.985 ;
        RECT 25.615 158.515 25.950 159.485 ;
        RECT 26.120 158.345 26.290 159.485 ;
        RECT 26.460 158.685 26.630 159.655 ;
        RECT 26.800 159.025 26.970 160.155 ;
        RECT 27.140 159.365 27.310 160.165 ;
        RECT 27.515 159.875 27.790 160.725 ;
        RECT 27.510 159.705 27.790 159.875 ;
        RECT 27.515 159.565 27.790 159.705 ;
        RECT 27.960 159.365 28.150 160.725 ;
        RECT 28.330 160.360 28.840 160.895 ;
        RECT 29.060 160.085 29.305 160.690 ;
        RECT 30.210 160.125 31.880 160.895 ;
        RECT 28.350 159.915 29.580 160.085 ;
        RECT 27.140 159.195 28.150 159.365 ;
        RECT 28.320 159.350 29.070 159.540 ;
        RECT 26.800 158.855 27.925 159.025 ;
        RECT 28.320 158.685 28.490 159.350 ;
        RECT 29.240 159.105 29.580 159.915 ;
        RECT 26.460 158.515 28.490 158.685 ;
        RECT 28.660 158.345 28.830 159.105 ;
        RECT 29.065 158.695 29.580 159.105 ;
        RECT 30.210 159.435 30.960 159.955 ;
        RECT 31.130 159.605 31.880 160.125 ;
        RECT 32.055 160.185 32.310 160.715 ;
        RECT 32.480 160.435 32.785 160.895 ;
        RECT 33.030 160.515 34.100 160.685 ;
        RECT 32.055 159.535 32.265 160.185 ;
        RECT 33.030 160.160 33.350 160.515 ;
        RECT 33.025 159.985 33.350 160.160 ;
        RECT 32.435 159.685 33.350 159.985 ;
        RECT 33.520 159.945 33.760 160.345 ;
        RECT 33.930 160.285 34.100 160.515 ;
        RECT 34.270 160.455 34.460 160.895 ;
        RECT 34.630 160.445 35.580 160.725 ;
        RECT 35.800 160.535 36.150 160.705 ;
        RECT 33.930 160.115 34.460 160.285 ;
        RECT 32.435 159.655 33.175 159.685 ;
        RECT 30.210 158.345 31.880 159.435 ;
        RECT 32.055 158.655 32.310 159.535 ;
        RECT 32.480 158.345 32.785 159.485 ;
        RECT 33.005 159.065 33.175 159.655 ;
        RECT 33.520 159.575 34.060 159.945 ;
        RECT 34.240 159.835 34.460 160.115 ;
        RECT 34.630 159.665 34.800 160.445 ;
        RECT 34.395 159.495 34.800 159.665 ;
        RECT 34.970 159.655 35.320 160.275 ;
        RECT 34.395 159.405 34.565 159.495 ;
        RECT 35.490 159.485 35.700 160.275 ;
        RECT 33.345 159.235 34.565 159.405 ;
        RECT 35.025 159.325 35.700 159.485 ;
        RECT 33.005 158.895 33.805 159.065 ;
        RECT 33.125 158.345 33.455 158.725 ;
        RECT 33.635 158.605 33.805 158.895 ;
        RECT 34.395 158.855 34.565 159.235 ;
        RECT 34.735 159.315 35.700 159.325 ;
        RECT 35.890 160.145 36.150 160.535 ;
        RECT 36.360 160.435 36.690 160.895 ;
        RECT 37.565 160.505 38.420 160.675 ;
        RECT 38.625 160.505 39.120 160.675 ;
        RECT 39.290 160.535 39.620 160.895 ;
        RECT 35.890 159.455 36.060 160.145 ;
        RECT 36.230 159.795 36.400 159.975 ;
        RECT 36.570 159.965 37.360 160.215 ;
        RECT 37.565 159.795 37.735 160.505 ;
        RECT 37.905 159.995 38.260 160.215 ;
        RECT 36.230 159.625 37.920 159.795 ;
        RECT 34.735 159.025 35.195 159.315 ;
        RECT 35.890 159.285 37.390 159.455 ;
        RECT 35.890 159.145 36.060 159.285 ;
        RECT 35.500 158.975 36.060 159.145 ;
        RECT 33.975 158.345 34.225 158.805 ;
        RECT 34.395 158.515 35.265 158.855 ;
        RECT 35.500 158.515 35.670 158.975 ;
        RECT 36.505 158.945 37.580 159.115 ;
        RECT 35.840 158.345 36.210 158.805 ;
        RECT 36.505 158.605 36.675 158.945 ;
        RECT 36.845 158.345 37.175 158.775 ;
        RECT 37.410 158.605 37.580 158.945 ;
        RECT 37.750 158.845 37.920 159.625 ;
        RECT 38.090 159.405 38.260 159.995 ;
        RECT 38.430 159.595 38.780 160.215 ;
        RECT 38.090 159.015 38.555 159.405 ;
        RECT 38.950 159.145 39.120 160.505 ;
        RECT 39.290 159.315 39.750 160.365 ;
        RECT 38.725 158.975 39.120 159.145 ;
        RECT 38.725 158.845 38.895 158.975 ;
        RECT 37.750 158.515 38.430 158.845 ;
        RECT 38.645 158.515 38.895 158.845 ;
        RECT 39.065 158.345 39.315 158.805 ;
        RECT 39.485 158.530 39.810 159.315 ;
        RECT 39.980 158.515 40.150 160.635 ;
        RECT 40.320 160.515 40.650 160.895 ;
        RECT 40.820 160.345 41.075 160.635 ;
        RECT 41.310 160.415 41.590 160.895 ;
        RECT 40.325 160.175 41.075 160.345 ;
        RECT 41.760 160.245 42.020 160.635 ;
        RECT 42.195 160.415 42.450 160.895 ;
        RECT 42.620 160.245 42.915 160.635 ;
        RECT 43.095 160.415 43.370 160.895 ;
        RECT 43.540 160.395 43.840 160.725 ;
        RECT 40.325 159.185 40.555 160.175 ;
        RECT 41.265 160.075 42.915 160.245 ;
        RECT 40.725 159.355 41.075 160.005 ;
        RECT 41.265 159.565 41.670 160.075 ;
        RECT 41.840 159.735 42.980 159.905 ;
        RECT 41.265 159.395 42.020 159.565 ;
        RECT 40.325 159.015 41.075 159.185 ;
        RECT 40.320 158.345 40.650 158.845 ;
        RECT 40.820 158.515 41.075 159.015 ;
        RECT 41.305 158.345 41.590 159.215 ;
        RECT 41.760 159.145 42.020 159.395 ;
        RECT 42.810 159.485 42.980 159.735 ;
        RECT 43.150 159.655 43.500 160.225 ;
        RECT 43.670 159.485 43.840 160.395 ;
        RECT 42.810 159.315 43.840 159.485 ;
        RECT 41.760 158.975 42.880 159.145 ;
        RECT 41.760 158.515 42.020 158.975 ;
        RECT 42.195 158.345 42.450 158.805 ;
        RECT 42.620 158.515 42.880 158.975 ;
        RECT 43.050 158.345 43.360 159.145 ;
        RECT 43.530 158.515 43.840 159.315 ;
        RECT 44.010 160.095 44.350 160.725 ;
        RECT 44.520 160.095 44.770 160.895 ;
        RECT 44.960 160.245 45.290 160.725 ;
        RECT 45.460 160.435 45.685 160.895 ;
        RECT 45.855 160.245 46.185 160.725 ;
        RECT 44.010 159.485 44.185 160.095 ;
        RECT 44.960 160.075 46.185 160.245 ;
        RECT 46.815 160.115 47.315 160.725 ;
        RECT 47.690 160.170 47.980 160.895 ;
        RECT 44.355 159.735 45.050 159.905 ;
        RECT 44.880 159.485 45.050 159.735 ;
        RECT 45.225 159.705 45.645 159.905 ;
        RECT 45.815 159.705 46.145 159.905 ;
        RECT 46.315 159.705 46.645 159.905 ;
        RECT 46.815 159.485 46.985 160.115 ;
        RECT 48.425 160.085 48.670 160.690 ;
        RECT 48.890 160.360 49.400 160.895 ;
        RECT 48.150 159.915 49.380 160.085 ;
        RECT 47.170 159.655 47.520 159.905 ;
        RECT 44.010 158.515 44.350 159.485 ;
        RECT 44.520 158.345 44.690 159.485 ;
        RECT 44.880 159.315 47.315 159.485 ;
        RECT 44.960 158.345 45.210 159.145 ;
        RECT 45.855 158.515 46.185 159.315 ;
        RECT 46.485 158.345 46.815 159.145 ;
        RECT 46.985 158.515 47.315 159.315 ;
        RECT 47.690 158.345 47.980 159.510 ;
        RECT 48.150 159.105 48.490 159.915 ;
        RECT 48.660 159.350 49.410 159.540 ;
        RECT 48.150 158.695 48.665 159.105 ;
        RECT 48.900 158.345 49.070 159.105 ;
        RECT 49.240 158.685 49.410 159.350 ;
        RECT 49.580 159.365 49.770 160.725 ;
        RECT 49.940 160.555 50.215 160.725 ;
        RECT 49.940 160.385 50.220 160.555 ;
        RECT 49.940 159.565 50.215 160.385 ;
        RECT 50.405 160.360 50.935 160.725 ;
        RECT 51.360 160.495 51.690 160.895 ;
        RECT 50.760 160.325 50.935 160.360 ;
        RECT 50.420 159.365 50.590 160.165 ;
        RECT 49.580 159.195 50.590 159.365 ;
        RECT 50.760 160.155 51.690 160.325 ;
        RECT 51.860 160.155 52.115 160.725 ;
        RECT 50.760 159.025 50.930 160.155 ;
        RECT 51.520 159.985 51.690 160.155 ;
        RECT 49.805 158.855 50.930 159.025 ;
        RECT 51.100 159.655 51.295 159.985 ;
        RECT 51.520 159.655 51.775 159.985 ;
        RECT 51.100 158.685 51.270 159.655 ;
        RECT 51.945 159.485 52.115 160.155 ;
        RECT 52.380 160.245 52.550 160.725 ;
        RECT 52.730 160.415 52.970 160.895 ;
        RECT 53.220 160.245 53.390 160.725 ;
        RECT 53.560 160.415 53.890 160.895 ;
        RECT 54.060 160.245 54.230 160.725 ;
        RECT 52.380 160.075 53.015 160.245 ;
        RECT 53.220 160.075 54.230 160.245 ;
        RECT 54.400 160.095 54.730 160.895 ;
        RECT 55.110 160.415 55.390 160.895 ;
        RECT 55.560 160.245 55.820 160.635 ;
        RECT 55.995 160.415 56.250 160.895 ;
        RECT 56.420 160.245 56.715 160.635 ;
        RECT 56.895 160.415 57.170 160.895 ;
        RECT 57.340 160.395 57.640 160.725 ;
        RECT 52.845 159.905 53.015 160.075 ;
        RECT 52.295 159.665 52.675 159.905 ;
        RECT 52.845 159.735 53.345 159.905 ;
        RECT 53.735 159.875 54.230 160.075 ;
        RECT 52.845 159.495 53.015 159.735 ;
        RECT 53.730 159.705 54.230 159.875 ;
        RECT 53.735 159.535 54.230 159.705 ;
        RECT 49.240 158.515 51.270 158.685 ;
        RECT 51.440 158.345 51.610 159.485 ;
        RECT 51.780 158.515 52.115 159.485 ;
        RECT 52.300 159.325 53.015 159.495 ;
        RECT 53.220 159.365 54.230 159.535 ;
        RECT 55.065 160.075 56.715 160.245 ;
        RECT 55.065 159.565 55.470 160.075 ;
        RECT 55.640 159.735 56.780 159.905 ;
        RECT 52.300 158.515 52.630 159.325 ;
        RECT 52.800 158.345 53.040 159.145 ;
        RECT 53.220 158.515 53.390 159.365 ;
        RECT 53.560 158.345 53.890 159.145 ;
        RECT 54.060 158.515 54.230 159.365 ;
        RECT 54.400 158.345 54.730 159.495 ;
        RECT 55.065 159.395 55.820 159.565 ;
        RECT 55.105 158.345 55.390 159.215 ;
        RECT 55.560 159.145 55.820 159.395 ;
        RECT 56.610 159.485 56.780 159.735 ;
        RECT 56.950 159.655 57.300 160.225 ;
        RECT 57.470 159.485 57.640 160.395 ;
        RECT 58.275 160.055 58.535 160.895 ;
        RECT 58.710 160.150 58.965 160.725 ;
        RECT 59.135 160.515 59.465 160.895 ;
        RECT 59.680 160.345 59.850 160.725 ;
        RECT 59.135 160.175 59.850 160.345 ;
        RECT 56.610 159.315 57.640 159.485 ;
        RECT 55.560 158.975 56.680 159.145 ;
        RECT 55.560 158.515 55.820 158.975 ;
        RECT 55.995 158.345 56.250 158.805 ;
        RECT 56.420 158.515 56.680 158.975 ;
        RECT 56.850 158.345 57.160 159.145 ;
        RECT 57.330 158.515 57.640 159.315 ;
        RECT 58.275 158.345 58.535 159.495 ;
        RECT 58.710 159.420 58.880 160.150 ;
        RECT 59.135 159.985 59.305 160.175 ;
        RECT 60.115 160.055 60.375 160.895 ;
        RECT 60.550 160.150 60.805 160.725 ;
        RECT 60.975 160.515 61.305 160.895 ;
        RECT 61.520 160.345 61.690 160.725 ;
        RECT 60.975 160.175 61.690 160.345 ;
        RECT 62.040 160.345 62.210 160.725 ;
        RECT 62.390 160.515 62.720 160.895 ;
        RECT 62.040 160.175 62.705 160.345 ;
        RECT 62.900 160.220 63.160 160.725 ;
        RECT 59.050 159.655 59.305 159.985 ;
        RECT 59.135 159.445 59.305 159.655 ;
        RECT 59.585 159.625 59.940 159.995 ;
        RECT 58.710 158.515 58.965 159.420 ;
        RECT 59.135 159.275 59.850 159.445 ;
        RECT 59.135 158.345 59.465 159.105 ;
        RECT 59.680 158.515 59.850 159.275 ;
        RECT 60.115 158.345 60.375 159.495 ;
        RECT 60.550 159.420 60.720 160.150 ;
        RECT 60.975 159.985 61.145 160.175 ;
        RECT 60.890 159.655 61.145 159.985 ;
        RECT 60.975 159.445 61.145 159.655 ;
        RECT 61.425 159.625 61.780 159.995 ;
        RECT 61.970 159.625 62.300 159.995 ;
        RECT 62.535 159.920 62.705 160.175 ;
        RECT 62.535 159.590 62.820 159.920 ;
        RECT 62.535 159.445 62.705 159.590 ;
        RECT 60.550 158.515 60.805 159.420 ;
        RECT 60.975 159.275 61.690 159.445 ;
        RECT 60.975 158.345 61.305 159.105 ;
        RECT 61.520 158.515 61.690 159.275 ;
        RECT 62.040 159.275 62.705 159.445 ;
        RECT 62.990 159.420 63.160 160.220 ;
        RECT 63.340 160.365 63.670 160.725 ;
        RECT 63.840 160.535 64.170 160.895 ;
        RECT 64.370 160.365 64.700 160.725 ;
        RECT 63.340 160.155 64.700 160.365 ;
        RECT 65.210 160.135 65.920 160.725 ;
        RECT 66.360 160.500 66.690 160.895 ;
        RECT 66.860 160.325 67.060 160.680 ;
        RECT 67.230 160.495 67.560 160.895 ;
        RECT 67.730 160.325 67.930 160.670 ;
        RECT 65.690 160.045 65.920 160.135 ;
        RECT 63.330 159.655 63.640 159.985 ;
        RECT 63.850 159.655 64.225 159.985 ;
        RECT 64.545 159.655 65.040 159.985 ;
        RECT 62.040 158.515 62.210 159.275 ;
        RECT 62.390 158.345 62.720 159.105 ;
        RECT 62.890 158.515 63.160 159.420 ;
        RECT 63.340 158.345 63.670 159.405 ;
        RECT 63.850 158.730 64.020 159.655 ;
        RECT 64.190 159.165 64.520 159.385 ;
        RECT 64.715 159.365 65.040 159.655 ;
        RECT 65.215 159.365 65.545 159.905 ;
        RECT 65.715 159.165 65.920 160.045 ;
        RECT 64.190 158.935 65.920 159.165 ;
        RECT 64.190 158.535 64.520 158.935 ;
        RECT 64.690 158.345 65.020 158.705 ;
        RECT 65.220 158.515 65.920 158.935 ;
        RECT 66.090 160.155 67.930 160.325 ;
        RECT 68.100 160.155 68.430 160.895 ;
        RECT 68.665 160.325 68.835 160.575 ;
        RECT 68.665 160.155 69.140 160.325 ;
        RECT 66.090 158.530 66.350 160.155 ;
        RECT 66.530 159.185 66.750 159.985 ;
        RECT 66.990 159.365 67.290 159.985 ;
        RECT 67.460 159.365 67.790 159.985 ;
        RECT 67.960 159.365 68.280 159.985 ;
        RECT 68.450 159.365 68.800 159.985 ;
        RECT 68.970 159.185 69.140 160.155 ;
        RECT 69.310 160.145 70.520 160.895 ;
        RECT 66.530 158.975 69.140 159.185 ;
        RECT 69.310 159.435 69.830 159.975 ;
        RECT 70.000 159.605 70.520 160.145 ;
        RECT 70.690 160.395 70.990 160.725 ;
        RECT 71.160 160.415 71.435 160.895 ;
        RECT 70.690 159.485 70.860 160.395 ;
        RECT 71.615 160.245 71.910 160.635 ;
        RECT 72.080 160.415 72.335 160.895 ;
        RECT 72.510 160.245 72.770 160.635 ;
        RECT 72.940 160.415 73.220 160.895 ;
        RECT 71.030 159.655 71.380 160.225 ;
        RECT 71.615 160.075 73.265 160.245 ;
        RECT 73.450 160.170 73.740 160.895 ;
        RECT 75.205 160.555 75.460 160.715 ;
        RECT 75.120 160.385 75.460 160.555 ;
        RECT 75.640 160.435 75.925 160.895 ;
        RECT 75.205 160.185 75.460 160.385 ;
        RECT 71.550 159.735 72.690 159.905 ;
        RECT 71.550 159.485 71.720 159.735 ;
        RECT 72.860 159.565 73.265 160.075 ;
        RECT 68.100 158.345 68.430 158.795 ;
        RECT 69.310 158.345 70.520 159.435 ;
        RECT 70.690 159.315 71.720 159.485 ;
        RECT 72.510 159.395 73.265 159.565 ;
        RECT 70.690 158.515 71.000 159.315 ;
        RECT 72.510 159.145 72.770 159.395 ;
        RECT 71.170 158.345 71.480 159.145 ;
        RECT 71.650 158.975 72.770 159.145 ;
        RECT 71.650 158.515 71.910 158.975 ;
        RECT 72.080 158.345 72.335 158.805 ;
        RECT 72.510 158.515 72.770 158.975 ;
        RECT 72.940 158.345 73.225 159.215 ;
        RECT 73.450 158.345 73.740 159.510 ;
        RECT 75.205 159.325 75.385 160.185 ;
        RECT 76.105 159.985 76.355 160.635 ;
        RECT 75.555 159.655 76.355 159.985 ;
        RECT 75.205 158.655 75.460 159.325 ;
        RECT 75.640 158.345 75.925 159.145 ;
        RECT 76.105 159.065 76.355 159.655 ;
        RECT 76.555 160.300 76.875 160.630 ;
        RECT 77.055 160.415 77.715 160.895 ;
        RECT 77.915 160.505 78.765 160.675 ;
        RECT 76.555 159.405 76.745 160.300 ;
        RECT 77.065 159.975 77.725 160.245 ;
        RECT 77.395 159.915 77.725 159.975 ;
        RECT 76.915 159.745 77.245 159.805 ;
        RECT 77.915 159.745 78.085 160.505 ;
        RECT 79.325 160.435 79.645 160.895 ;
        RECT 79.845 160.255 80.095 160.685 ;
        RECT 80.385 160.455 80.795 160.895 ;
        RECT 80.965 160.515 81.980 160.715 ;
        RECT 78.255 160.085 79.505 160.255 ;
        RECT 78.255 159.965 78.585 160.085 ;
        RECT 76.915 159.575 78.815 159.745 ;
        RECT 76.555 159.235 78.475 159.405 ;
        RECT 76.555 159.215 76.875 159.235 ;
        RECT 76.105 158.555 76.435 159.065 ;
        RECT 76.705 158.605 76.875 159.215 ;
        RECT 78.645 159.065 78.815 159.575 ;
        RECT 78.985 159.505 79.165 159.915 ;
        RECT 79.335 159.325 79.505 160.085 ;
        RECT 77.045 158.345 77.375 159.035 ;
        RECT 77.605 158.895 78.815 159.065 ;
        RECT 78.985 159.015 79.505 159.325 ;
        RECT 79.675 159.915 80.095 160.255 ;
        RECT 80.385 159.915 80.795 160.245 ;
        RECT 79.675 159.145 79.865 159.915 ;
        RECT 80.965 159.785 81.135 160.515 ;
        RECT 82.280 160.345 82.450 160.675 ;
        RECT 82.620 160.515 82.950 160.895 ;
        RECT 81.305 159.965 81.655 160.335 ;
        RECT 80.965 159.745 81.385 159.785 ;
        RECT 80.035 159.575 81.385 159.745 ;
        RECT 80.035 159.415 80.285 159.575 ;
        RECT 80.795 159.145 81.045 159.405 ;
        RECT 79.675 158.895 81.045 159.145 ;
        RECT 77.605 158.605 77.845 158.895 ;
        RECT 78.645 158.815 78.815 158.895 ;
        RECT 78.045 158.345 78.465 158.725 ;
        RECT 78.645 158.565 79.275 158.815 ;
        RECT 79.745 158.345 80.075 158.725 ;
        RECT 80.245 158.605 80.415 158.895 ;
        RECT 81.215 158.730 81.385 159.575 ;
        RECT 81.835 159.405 82.055 160.275 ;
        RECT 82.280 160.155 82.975 160.345 ;
        RECT 81.555 159.025 82.055 159.405 ;
        RECT 82.225 159.355 82.635 159.975 ;
        RECT 82.805 159.185 82.975 160.155 ;
        RECT 82.280 159.015 82.975 159.185 ;
        RECT 80.595 158.345 80.975 158.725 ;
        RECT 81.215 158.560 82.045 158.730 ;
        RECT 82.280 158.515 82.450 159.015 ;
        RECT 82.620 158.345 82.950 158.845 ;
        RECT 83.165 158.515 83.390 160.635 ;
        RECT 83.560 160.515 83.890 160.895 ;
        RECT 84.060 160.345 84.230 160.635 ;
        RECT 83.565 160.175 84.230 160.345 ;
        RECT 84.490 160.220 84.750 160.725 ;
        RECT 84.930 160.515 85.260 160.895 ;
        RECT 85.440 160.345 85.610 160.725 ;
        RECT 83.565 159.185 83.795 160.175 ;
        RECT 83.965 159.355 84.315 160.005 ;
        RECT 84.490 159.420 84.660 160.220 ;
        RECT 84.945 160.175 85.610 160.345 ;
        RECT 84.945 159.920 85.115 160.175 ;
        RECT 86.075 160.115 86.575 160.725 ;
        RECT 84.830 159.590 85.115 159.920 ;
        RECT 85.350 159.625 85.680 159.995 ;
        RECT 85.870 159.655 86.220 159.905 ;
        RECT 84.945 159.445 85.115 159.590 ;
        RECT 86.405 159.485 86.575 160.115 ;
        RECT 87.205 160.245 87.535 160.725 ;
        RECT 87.705 160.435 87.930 160.895 ;
        RECT 88.100 160.245 88.430 160.725 ;
        RECT 87.205 160.075 88.430 160.245 ;
        RECT 88.620 160.095 88.870 160.895 ;
        RECT 89.040 160.095 89.380 160.725 ;
        RECT 86.745 159.705 87.075 159.905 ;
        RECT 87.245 159.705 87.575 159.905 ;
        RECT 87.745 159.705 88.165 159.905 ;
        RECT 88.340 159.735 89.035 159.905 ;
        RECT 88.340 159.485 88.510 159.735 ;
        RECT 89.205 159.485 89.380 160.095 ;
        RECT 89.825 160.085 90.070 160.690 ;
        RECT 90.290 160.360 90.800 160.895 ;
        RECT 83.565 159.015 84.230 159.185 ;
        RECT 83.560 158.345 83.890 158.845 ;
        RECT 84.060 158.515 84.230 159.015 ;
        RECT 84.490 158.515 84.760 159.420 ;
        RECT 84.945 159.275 85.610 159.445 ;
        RECT 84.930 158.345 85.260 159.105 ;
        RECT 85.440 158.515 85.610 159.275 ;
        RECT 86.075 159.315 88.510 159.485 ;
        RECT 86.075 158.515 86.405 159.315 ;
        RECT 86.575 158.345 86.905 159.145 ;
        RECT 87.205 158.515 87.535 159.315 ;
        RECT 88.180 158.345 88.430 159.145 ;
        RECT 88.700 158.345 88.870 159.485 ;
        RECT 89.040 158.515 89.380 159.485 ;
        RECT 89.550 159.915 90.780 160.085 ;
        RECT 89.550 159.105 89.890 159.915 ;
        RECT 90.060 159.350 90.810 159.540 ;
        RECT 89.550 158.695 90.065 159.105 ;
        RECT 90.300 158.345 90.470 159.105 ;
        RECT 90.640 158.685 90.810 159.350 ;
        RECT 90.980 159.365 91.170 160.725 ;
        RECT 91.340 160.215 91.615 160.725 ;
        RECT 91.805 160.360 92.335 160.725 ;
        RECT 92.760 160.495 93.090 160.895 ;
        RECT 92.160 160.325 92.335 160.360 ;
        RECT 91.340 160.045 91.620 160.215 ;
        RECT 91.340 159.565 91.615 160.045 ;
        RECT 91.820 159.365 91.990 160.165 ;
        RECT 90.980 159.195 91.990 159.365 ;
        RECT 92.160 160.155 93.090 160.325 ;
        RECT 93.260 160.155 93.515 160.725 ;
        RECT 93.780 160.345 93.950 160.725 ;
        RECT 94.130 160.515 94.460 160.895 ;
        RECT 93.780 160.175 94.445 160.345 ;
        RECT 94.640 160.220 94.900 160.725 ;
        RECT 92.160 159.025 92.330 160.155 ;
        RECT 92.920 159.985 93.090 160.155 ;
        RECT 91.205 158.855 92.330 159.025 ;
        RECT 92.500 159.655 92.695 159.985 ;
        RECT 92.920 159.655 93.175 159.985 ;
        RECT 92.500 158.685 92.670 159.655 ;
        RECT 93.345 159.485 93.515 160.155 ;
        RECT 93.710 159.625 94.040 159.995 ;
        RECT 94.275 159.920 94.445 160.175 ;
        RECT 90.640 158.515 92.670 158.685 ;
        RECT 92.840 158.345 93.010 159.485 ;
        RECT 93.180 158.515 93.515 159.485 ;
        RECT 94.275 159.590 94.560 159.920 ;
        RECT 94.275 159.445 94.445 159.590 ;
        RECT 93.780 159.275 94.445 159.445 ;
        RECT 94.730 159.420 94.900 160.220 ;
        RECT 93.780 158.515 93.950 159.275 ;
        RECT 94.130 158.345 94.460 159.105 ;
        RECT 94.630 158.515 94.900 159.420 ;
        RECT 95.530 160.095 95.870 160.725 ;
        RECT 96.040 160.095 96.290 160.895 ;
        RECT 96.480 160.245 96.810 160.725 ;
        RECT 96.980 160.435 97.205 160.895 ;
        RECT 97.375 160.245 97.705 160.725 ;
        RECT 95.530 159.485 95.705 160.095 ;
        RECT 96.480 160.075 97.705 160.245 ;
        RECT 98.335 160.115 98.835 160.725 ;
        RECT 99.210 160.170 99.500 160.895 ;
        RECT 99.875 160.115 100.375 160.725 ;
        RECT 95.875 159.735 96.570 159.905 ;
        RECT 96.400 159.485 96.570 159.735 ;
        RECT 96.745 159.705 97.165 159.905 ;
        RECT 97.335 159.705 97.665 159.905 ;
        RECT 97.835 159.705 98.165 159.905 ;
        RECT 98.335 159.485 98.505 160.115 ;
        RECT 98.690 159.655 99.040 159.905 ;
        RECT 99.670 159.655 100.020 159.905 ;
        RECT 95.530 158.515 95.870 159.485 ;
        RECT 96.040 158.345 96.210 159.485 ;
        RECT 96.400 159.315 98.835 159.485 ;
        RECT 96.480 158.345 96.730 159.145 ;
        RECT 97.375 158.515 97.705 159.315 ;
        RECT 98.005 158.345 98.335 159.145 ;
        RECT 98.505 158.515 98.835 159.315 ;
        RECT 99.210 158.345 99.500 159.510 ;
        RECT 100.205 159.485 100.375 160.115 ;
        RECT 101.005 160.245 101.335 160.725 ;
        RECT 101.505 160.435 101.730 160.895 ;
        RECT 101.900 160.245 102.230 160.725 ;
        RECT 101.005 160.075 102.230 160.245 ;
        RECT 102.420 160.095 102.670 160.895 ;
        RECT 102.840 160.095 103.180 160.725 ;
        RECT 100.545 159.705 100.875 159.905 ;
        RECT 101.045 159.705 101.375 159.905 ;
        RECT 101.545 159.705 101.965 159.905 ;
        RECT 102.140 159.735 102.835 159.905 ;
        RECT 102.140 159.485 102.310 159.735 ;
        RECT 103.005 159.485 103.180 160.095 ;
        RECT 104.310 160.075 104.540 160.895 ;
        RECT 104.710 160.095 105.040 160.725 ;
        RECT 104.290 159.655 104.620 159.905 ;
        RECT 104.790 159.495 105.040 160.095 ;
        RECT 105.210 160.075 105.420 160.895 ;
        RECT 105.650 160.145 106.860 160.895 ;
        RECT 107.035 160.495 107.370 160.895 ;
        RECT 107.540 160.325 107.745 160.725 ;
        RECT 107.955 160.415 108.230 160.895 ;
        RECT 108.440 160.395 108.700 160.725 ;
        RECT 99.875 159.315 102.310 159.485 ;
        RECT 99.875 158.515 100.205 159.315 ;
        RECT 100.375 158.345 100.705 159.145 ;
        RECT 101.005 158.515 101.335 159.315 ;
        RECT 101.980 158.345 102.230 159.145 ;
        RECT 102.500 158.345 102.670 159.485 ;
        RECT 102.840 158.515 103.180 159.485 ;
        RECT 104.310 158.345 104.540 159.485 ;
        RECT 104.710 158.515 105.040 159.495 ;
        RECT 105.210 158.345 105.420 159.485 ;
        RECT 105.650 159.435 106.170 159.975 ;
        RECT 106.340 159.605 106.860 160.145 ;
        RECT 107.060 160.155 107.745 160.325 ;
        RECT 105.650 158.345 106.860 159.435 ;
        RECT 107.060 159.125 107.400 160.155 ;
        RECT 107.570 159.485 107.820 159.985 ;
        RECT 108.000 159.655 108.360 160.235 ;
        RECT 108.530 159.485 108.700 160.395 ;
        RECT 109.330 160.125 111.000 160.895 ;
        RECT 111.170 160.145 112.380 160.895 ;
        RECT 107.570 159.315 108.700 159.485 ;
        RECT 107.060 158.950 107.725 159.125 ;
        RECT 107.035 158.345 107.370 158.770 ;
        RECT 107.540 158.545 107.725 158.950 ;
        RECT 107.930 158.345 108.260 159.125 ;
        RECT 108.430 158.545 108.700 159.315 ;
        RECT 109.330 159.435 110.080 159.955 ;
        RECT 110.250 159.605 111.000 160.125 ;
        RECT 111.170 159.435 111.690 159.975 ;
        RECT 111.860 159.605 112.380 160.145 ;
        RECT 109.330 158.345 111.000 159.435 ;
        RECT 111.170 158.345 112.380 159.435 ;
        RECT 18.165 158.175 112.465 158.345 ;
        RECT 18.250 157.085 19.460 158.175 ;
        RECT 18.250 156.375 18.770 156.915 ;
        RECT 18.940 156.545 19.460 157.085 ;
        RECT 19.635 156.985 19.890 157.865 ;
        RECT 20.060 157.035 20.365 158.175 ;
        RECT 20.705 157.795 21.035 158.175 ;
        RECT 21.215 157.625 21.385 157.915 ;
        RECT 21.555 157.715 21.805 158.175 ;
        RECT 20.585 157.455 21.385 157.625 ;
        RECT 21.975 157.665 22.845 158.005 ;
        RECT 18.250 155.625 19.460 156.375 ;
        RECT 19.635 156.335 19.845 156.985 ;
        RECT 20.585 156.865 20.755 157.455 ;
        RECT 21.975 157.285 22.145 157.665 ;
        RECT 23.080 157.545 23.250 158.005 ;
        RECT 23.420 157.715 23.790 158.175 ;
        RECT 24.085 157.575 24.255 157.915 ;
        RECT 24.425 157.745 24.755 158.175 ;
        RECT 24.990 157.575 25.160 157.915 ;
        RECT 20.925 157.115 22.145 157.285 ;
        RECT 22.315 157.205 22.775 157.495 ;
        RECT 23.080 157.375 23.640 157.545 ;
        RECT 24.085 157.405 25.160 157.575 ;
        RECT 25.330 157.675 26.010 158.005 ;
        RECT 26.225 157.675 26.475 158.005 ;
        RECT 26.645 157.715 26.895 158.175 ;
        RECT 23.470 157.235 23.640 157.375 ;
        RECT 22.315 157.195 23.280 157.205 ;
        RECT 21.975 157.025 22.145 157.115 ;
        RECT 22.605 157.035 23.280 157.195 ;
        RECT 20.015 156.835 20.755 156.865 ;
        RECT 20.015 156.535 20.930 156.835 ;
        RECT 20.605 156.360 20.930 156.535 ;
        RECT 19.635 155.805 19.890 156.335 ;
        RECT 20.060 155.625 20.365 156.085 ;
        RECT 20.610 156.005 20.930 156.360 ;
        RECT 21.100 156.575 21.640 156.945 ;
        RECT 21.975 156.855 22.380 157.025 ;
        RECT 21.100 156.175 21.340 156.575 ;
        RECT 21.820 156.405 22.040 156.685 ;
        RECT 21.510 156.235 22.040 156.405 ;
        RECT 21.510 156.005 21.680 156.235 ;
        RECT 22.210 156.075 22.380 156.855 ;
        RECT 22.550 156.245 22.900 156.865 ;
        RECT 23.070 156.245 23.280 157.035 ;
        RECT 23.470 157.065 24.970 157.235 ;
        RECT 23.470 156.375 23.640 157.065 ;
        RECT 25.330 156.895 25.500 157.675 ;
        RECT 26.305 157.545 26.475 157.675 ;
        RECT 23.810 156.725 25.500 156.895 ;
        RECT 25.670 157.115 26.135 157.505 ;
        RECT 26.305 157.375 26.700 157.545 ;
        RECT 23.810 156.545 23.980 156.725 ;
        RECT 20.610 155.835 21.680 156.005 ;
        RECT 21.850 155.625 22.040 156.065 ;
        RECT 22.210 155.795 23.160 156.075 ;
        RECT 23.470 155.985 23.730 156.375 ;
        RECT 24.150 156.305 24.940 156.555 ;
        RECT 23.380 155.815 23.730 155.985 ;
        RECT 23.940 155.625 24.270 156.085 ;
        RECT 25.145 156.015 25.315 156.725 ;
        RECT 25.670 156.525 25.840 157.115 ;
        RECT 25.485 156.305 25.840 156.525 ;
        RECT 26.010 156.305 26.360 156.925 ;
        RECT 26.530 156.015 26.700 157.375 ;
        RECT 27.065 157.205 27.390 157.990 ;
        RECT 26.870 156.155 27.330 157.205 ;
        RECT 25.145 155.845 26.000 156.015 ;
        RECT 26.205 155.845 26.700 156.015 ;
        RECT 26.870 155.625 27.200 155.985 ;
        RECT 27.560 155.885 27.730 158.005 ;
        RECT 27.900 157.675 28.230 158.175 ;
        RECT 28.400 157.505 28.655 158.005 ;
        RECT 27.905 157.335 28.655 157.505 ;
        RECT 27.905 156.345 28.135 157.335 ;
        RECT 28.305 156.515 28.655 157.165 ;
        RECT 29.350 157.035 29.560 158.175 ;
        RECT 29.730 157.025 30.060 158.005 ;
        RECT 30.230 157.035 30.460 158.175 ;
        RECT 30.670 157.415 31.185 157.825 ;
        RECT 31.420 157.415 31.590 158.175 ;
        RECT 31.760 157.835 33.790 158.005 ;
        RECT 27.905 156.175 28.655 156.345 ;
        RECT 27.900 155.625 28.230 156.005 ;
        RECT 28.400 155.885 28.655 156.175 ;
        RECT 29.350 155.625 29.560 156.445 ;
        RECT 29.730 156.425 29.980 157.025 ;
        RECT 30.150 156.615 30.480 156.865 ;
        RECT 30.670 156.605 31.010 157.415 ;
        RECT 31.760 157.170 31.930 157.835 ;
        RECT 32.325 157.495 33.450 157.665 ;
        RECT 31.180 156.980 31.930 157.170 ;
        RECT 32.100 157.155 33.110 157.325 ;
        RECT 29.730 155.795 30.060 156.425 ;
        RECT 30.230 155.625 30.460 156.445 ;
        RECT 30.670 156.435 31.900 156.605 ;
        RECT 30.945 155.830 31.190 156.435 ;
        RECT 31.410 155.625 31.920 156.160 ;
        RECT 32.100 155.795 32.290 157.155 ;
        RECT 32.460 156.815 32.735 156.955 ;
        RECT 32.460 156.645 32.740 156.815 ;
        RECT 32.460 155.795 32.735 156.645 ;
        RECT 32.940 156.355 33.110 157.155 ;
        RECT 33.280 156.365 33.450 157.495 ;
        RECT 33.620 156.865 33.790 157.835 ;
        RECT 33.960 157.035 34.130 158.175 ;
        RECT 34.300 157.035 34.635 158.005 ;
        RECT 33.620 156.535 33.815 156.865 ;
        RECT 34.040 156.535 34.295 156.865 ;
        RECT 34.040 156.365 34.210 156.535 ;
        RECT 34.465 156.365 34.635 157.035 ;
        RECT 34.810 157.010 35.100 158.175 ;
        RECT 35.270 157.085 36.480 158.175 ;
        RECT 36.855 157.205 37.185 158.005 ;
        RECT 37.355 157.375 37.685 158.175 ;
        RECT 37.985 157.205 38.315 158.005 ;
        RECT 38.960 157.375 39.210 158.175 ;
        RECT 35.270 156.545 35.790 157.085 ;
        RECT 36.855 157.035 39.290 157.205 ;
        RECT 39.480 157.035 39.650 158.175 ;
        RECT 39.820 157.035 40.160 158.005 ;
        RECT 40.535 157.205 40.865 158.005 ;
        RECT 41.035 157.375 41.365 158.175 ;
        RECT 41.665 157.205 41.995 158.005 ;
        RECT 42.640 157.375 42.890 158.175 ;
        RECT 40.535 157.035 42.970 157.205 ;
        RECT 43.160 157.035 43.330 158.175 ;
        RECT 43.500 157.035 43.840 158.005 ;
        RECT 44.100 157.430 44.370 158.175 ;
        RECT 45.000 158.170 51.275 158.175 ;
        RECT 44.540 157.260 44.830 158.000 ;
        RECT 45.000 157.445 45.255 158.170 ;
        RECT 45.440 157.275 45.700 158.000 ;
        RECT 45.870 157.445 46.115 158.170 ;
        RECT 46.300 157.275 46.560 158.000 ;
        RECT 46.730 157.445 46.975 158.170 ;
        RECT 47.160 157.275 47.420 158.000 ;
        RECT 47.590 157.445 47.835 158.170 ;
        RECT 48.005 157.275 48.265 158.000 ;
        RECT 48.435 157.445 48.695 158.170 ;
        RECT 48.865 157.275 49.125 158.000 ;
        RECT 49.295 157.445 49.555 158.170 ;
        RECT 49.725 157.275 49.985 158.000 ;
        RECT 50.155 157.445 50.415 158.170 ;
        RECT 50.585 157.275 50.845 158.000 ;
        RECT 51.015 157.375 51.275 158.170 ;
        RECT 45.440 157.260 50.845 157.275 ;
        RECT 35.960 156.375 36.480 156.915 ;
        RECT 36.650 156.615 37.000 156.865 ;
        RECT 37.185 156.405 37.355 157.035 ;
        RECT 37.525 156.615 37.855 156.815 ;
        RECT 38.025 156.615 38.355 156.815 ;
        RECT 38.525 156.615 38.945 156.815 ;
        RECT 39.120 156.785 39.290 157.035 ;
        RECT 39.120 156.615 39.815 156.785 ;
        RECT 39.985 156.475 40.160 157.035 ;
        RECT 40.330 156.615 40.680 156.865 ;
        RECT 33.280 156.195 34.210 156.365 ;
        RECT 33.280 156.160 33.455 156.195 ;
        RECT 32.925 155.795 33.455 156.160 ;
        RECT 33.880 155.625 34.210 156.025 ;
        RECT 34.380 155.795 34.635 156.365 ;
        RECT 34.810 155.625 35.100 156.350 ;
        RECT 35.270 155.625 36.480 156.375 ;
        RECT 36.855 155.795 37.355 156.405 ;
        RECT 37.985 156.275 39.210 156.445 ;
        RECT 39.930 156.425 40.160 156.475 ;
        RECT 37.985 155.795 38.315 156.275 ;
        RECT 38.485 155.625 38.710 156.085 ;
        RECT 38.880 155.795 39.210 156.275 ;
        RECT 39.400 155.625 39.650 156.425 ;
        RECT 39.820 155.795 40.160 156.425 ;
        RECT 40.865 156.405 41.035 157.035 ;
        RECT 41.205 156.615 41.535 156.815 ;
        RECT 41.705 156.615 42.035 156.815 ;
        RECT 42.205 156.615 42.625 156.815 ;
        RECT 42.800 156.785 42.970 157.035 ;
        RECT 42.800 156.615 43.495 156.785 ;
        RECT 40.535 155.795 41.035 156.405 ;
        RECT 41.665 156.275 42.890 156.445 ;
        RECT 43.665 156.425 43.840 157.035 ;
        RECT 41.665 155.795 41.995 156.275 ;
        RECT 42.165 155.625 42.390 156.085 ;
        RECT 42.560 155.795 42.890 156.275 ;
        RECT 43.080 155.625 43.330 156.425 ;
        RECT 43.500 155.795 43.840 156.425 ;
        RECT 44.100 157.035 50.845 157.260 ;
        RECT 44.100 156.445 45.265 157.035 ;
        RECT 51.445 156.865 51.695 158.000 ;
        RECT 51.875 157.365 52.135 158.175 ;
        RECT 52.310 156.865 52.555 158.005 ;
        RECT 52.735 157.365 53.030 158.175 ;
        RECT 53.310 157.715 53.480 158.175 ;
        RECT 53.650 157.225 53.980 158.005 ;
        RECT 54.150 157.375 54.320 158.175 ;
        RECT 53.210 157.205 53.980 157.225 ;
        RECT 54.490 157.205 54.820 158.005 ;
        RECT 54.990 157.375 55.160 158.175 ;
        RECT 55.330 157.205 55.660 158.005 ;
        RECT 53.210 157.035 55.660 157.205 ;
        RECT 55.920 157.035 56.215 158.175 ;
        RECT 45.435 156.615 52.555 156.865 ;
        RECT 44.100 156.275 50.845 156.445 ;
        RECT 44.100 155.625 44.400 156.105 ;
        RECT 44.570 155.820 44.830 156.275 ;
        RECT 45.000 155.625 45.260 156.105 ;
        RECT 45.440 155.820 45.700 156.275 ;
        RECT 45.870 155.625 46.120 156.105 ;
        RECT 46.300 155.820 46.560 156.275 ;
        RECT 46.730 155.625 46.980 156.105 ;
        RECT 47.160 155.820 47.420 156.275 ;
        RECT 47.590 155.625 47.835 156.105 ;
        RECT 48.005 155.820 48.280 156.275 ;
        RECT 48.450 155.625 48.695 156.105 ;
        RECT 48.865 155.820 49.125 156.275 ;
        RECT 49.295 155.625 49.555 156.105 ;
        RECT 49.725 155.820 49.985 156.275 ;
        RECT 50.155 155.625 50.415 156.105 ;
        RECT 50.585 155.820 50.845 156.275 ;
        RECT 51.015 155.625 51.275 156.185 ;
        RECT 51.445 155.805 51.695 156.615 ;
        RECT 51.875 155.625 52.135 156.150 ;
        RECT 52.305 155.805 52.555 156.615 ;
        RECT 52.725 156.305 53.040 156.865 ;
        RECT 53.210 156.445 53.560 157.035 ;
        RECT 56.435 157.025 56.695 158.175 ;
        RECT 56.870 157.100 57.125 158.005 ;
        RECT 57.295 157.415 57.625 158.175 ;
        RECT 57.840 157.245 58.010 158.005 ;
        RECT 53.730 156.615 56.240 156.865 ;
        RECT 53.210 156.265 55.580 156.445 ;
        RECT 52.735 155.625 53.040 156.135 ;
        RECT 53.310 155.625 53.560 156.090 ;
        RECT 53.730 155.795 53.900 156.265 ;
        RECT 54.150 155.625 54.320 156.085 ;
        RECT 54.570 155.795 54.740 156.265 ;
        RECT 54.990 155.625 55.160 156.085 ;
        RECT 55.410 155.795 55.580 156.265 ;
        RECT 55.950 155.625 56.215 156.085 ;
        RECT 56.435 155.625 56.695 156.465 ;
        RECT 56.870 156.370 57.040 157.100 ;
        RECT 57.295 157.075 58.010 157.245 ;
        RECT 59.280 157.245 59.450 158.005 ;
        RECT 59.630 157.415 59.960 158.175 ;
        RECT 59.280 157.075 59.945 157.245 ;
        RECT 60.130 157.100 60.400 158.005 ;
        RECT 57.295 156.865 57.465 157.075 ;
        RECT 59.775 156.930 59.945 157.075 ;
        RECT 57.210 156.535 57.465 156.865 ;
        RECT 56.870 155.795 57.125 156.370 ;
        RECT 57.295 156.345 57.465 156.535 ;
        RECT 57.745 156.525 58.100 156.895 ;
        RECT 59.210 156.525 59.540 156.895 ;
        RECT 59.775 156.600 60.060 156.930 ;
        RECT 59.775 156.345 59.945 156.600 ;
        RECT 57.295 156.175 58.010 156.345 ;
        RECT 57.295 155.625 57.625 156.005 ;
        RECT 57.840 155.795 58.010 156.175 ;
        RECT 59.280 156.175 59.945 156.345 ;
        RECT 60.230 156.300 60.400 157.100 ;
        RECT 60.570 157.010 60.860 158.175 ;
        RECT 62.040 157.245 62.210 158.005 ;
        RECT 62.425 157.415 62.755 158.175 ;
        RECT 62.040 157.075 62.755 157.245 ;
        RECT 62.925 157.100 63.180 158.005 ;
        RECT 61.950 156.525 62.305 156.895 ;
        RECT 62.585 156.865 62.755 157.075 ;
        RECT 62.585 156.535 62.840 156.865 ;
        RECT 59.280 155.795 59.450 156.175 ;
        RECT 59.630 155.625 59.960 156.005 ;
        RECT 60.140 155.795 60.400 156.300 ;
        RECT 60.570 155.625 60.860 156.350 ;
        RECT 62.585 156.345 62.755 156.535 ;
        RECT 63.010 156.370 63.180 157.100 ;
        RECT 63.355 157.025 63.615 158.175 ;
        RECT 64.715 157.025 64.975 158.175 ;
        RECT 65.150 157.100 65.405 158.005 ;
        RECT 65.575 157.415 65.905 158.175 ;
        RECT 66.120 157.245 66.290 158.005 ;
        RECT 62.040 156.175 62.755 156.345 ;
        RECT 62.040 155.795 62.210 156.175 ;
        RECT 62.425 155.625 62.755 156.005 ;
        RECT 62.925 155.795 63.180 156.370 ;
        RECT 63.355 155.625 63.615 156.465 ;
        RECT 64.715 155.625 64.975 156.465 ;
        RECT 65.150 156.370 65.320 157.100 ;
        RECT 65.575 157.075 66.290 157.245 ;
        RECT 66.620 157.235 66.880 158.005 ;
        RECT 67.050 157.405 67.380 158.175 ;
        RECT 67.550 157.835 68.670 158.005 ;
        RECT 67.550 157.235 67.740 157.835 ;
        RECT 65.575 156.865 65.745 157.075 ;
        RECT 66.620 157.065 67.740 157.235 ;
        RECT 67.910 157.250 68.240 157.665 ;
        RECT 68.410 157.640 68.670 157.835 ;
        RECT 68.900 157.455 69.230 158.175 ;
        RECT 69.400 157.250 69.590 158.005 ;
        RECT 69.760 157.455 70.090 158.175 ;
        RECT 70.260 157.250 70.520 158.005 ;
        RECT 70.690 157.715 70.950 158.175 ;
        RECT 67.910 157.080 70.520 157.250 ;
        RECT 65.490 156.535 65.745 156.865 ;
        RECT 65.150 155.795 65.405 156.370 ;
        RECT 65.575 156.345 65.745 156.535 ;
        RECT 66.025 156.525 66.380 156.895 ;
        RECT 66.610 156.785 67.505 156.835 ;
        RECT 66.610 156.615 67.560 156.785 ;
        RECT 67.730 156.615 68.700 156.895 ;
        RECT 69.160 156.615 70.020 156.905 ;
        RECT 65.575 156.175 66.290 156.345 ;
        RECT 66.610 156.305 66.950 156.615 ;
        RECT 65.575 155.625 65.905 156.005 ;
        RECT 66.120 155.795 66.290 156.175 ;
        RECT 67.120 156.175 69.660 156.385 ;
        RECT 67.120 156.055 67.310 156.175 ;
        RECT 69.830 156.005 70.020 156.430 ;
        RECT 70.190 156.210 70.520 157.080 ;
        RECT 70.690 156.535 70.980 157.510 ;
        RECT 71.150 157.415 71.665 157.825 ;
        RECT 71.900 157.415 72.070 158.175 ;
        RECT 72.240 157.835 74.270 158.005 ;
        RECT 71.150 156.605 71.490 157.415 ;
        RECT 72.240 157.170 72.410 157.835 ;
        RECT 72.805 157.495 73.930 157.665 ;
        RECT 71.660 156.980 72.410 157.170 ;
        RECT 72.580 157.155 73.590 157.325 ;
        RECT 71.150 156.435 72.380 156.605 ;
        RECT 68.900 155.985 70.020 156.005 ;
        RECT 66.620 155.625 66.950 155.985 ;
        RECT 67.480 155.625 67.810 155.985 ;
        RECT 68.340 155.625 68.670 155.985 ;
        RECT 68.900 155.795 70.970 155.985 ;
        RECT 71.425 155.830 71.670 156.435 ;
        RECT 71.890 155.625 72.400 156.160 ;
        RECT 72.580 155.795 72.770 157.155 ;
        RECT 72.940 156.135 73.215 156.955 ;
        RECT 73.420 156.355 73.590 157.155 ;
        RECT 73.760 156.365 73.930 157.495 ;
        RECT 74.100 156.865 74.270 157.835 ;
        RECT 74.440 157.035 74.610 158.175 ;
        RECT 74.780 157.035 75.115 158.005 ;
        RECT 74.100 156.535 74.295 156.865 ;
        RECT 74.520 156.535 74.775 156.865 ;
        RECT 74.520 156.365 74.690 156.535 ;
        RECT 74.945 156.365 75.115 157.035 ;
        RECT 73.760 156.195 74.690 156.365 ;
        RECT 73.760 156.160 73.935 156.195 ;
        RECT 72.940 155.965 73.220 156.135 ;
        RECT 72.940 155.795 73.215 155.965 ;
        RECT 73.405 155.795 73.935 156.160 ;
        RECT 74.360 155.625 74.690 156.025 ;
        RECT 74.860 155.795 75.115 156.365 ;
        RECT 75.665 157.195 75.920 157.865 ;
        RECT 76.100 157.375 76.385 158.175 ;
        RECT 76.565 157.455 76.895 157.965 ;
        RECT 75.665 156.335 75.845 157.195 ;
        RECT 76.565 156.865 76.815 157.455 ;
        RECT 77.165 157.305 77.335 157.915 ;
        RECT 77.505 157.485 77.835 158.175 ;
        RECT 78.065 157.625 78.305 157.915 ;
        RECT 78.505 157.795 78.925 158.175 ;
        RECT 79.105 157.705 79.735 157.955 ;
        RECT 80.205 157.795 80.535 158.175 ;
        RECT 79.105 157.625 79.275 157.705 ;
        RECT 80.705 157.625 80.875 157.915 ;
        RECT 81.055 157.795 81.435 158.175 ;
        RECT 81.675 157.790 82.505 157.960 ;
        RECT 78.065 157.455 79.275 157.625 ;
        RECT 76.015 156.535 76.815 156.865 ;
        RECT 75.665 156.135 75.920 156.335 ;
        RECT 75.580 155.965 75.920 156.135 ;
        RECT 75.665 155.805 75.920 155.965 ;
        RECT 76.100 155.625 76.385 156.085 ;
        RECT 76.565 155.885 76.815 156.535 ;
        RECT 77.015 157.285 77.335 157.305 ;
        RECT 77.015 157.115 78.935 157.285 ;
        RECT 77.015 156.220 77.205 157.115 ;
        RECT 79.105 156.945 79.275 157.455 ;
        RECT 79.445 157.195 79.965 157.505 ;
        RECT 77.375 156.775 79.275 156.945 ;
        RECT 77.375 156.715 77.705 156.775 ;
        RECT 77.855 156.545 78.185 156.605 ;
        RECT 77.525 156.275 78.185 156.545 ;
        RECT 77.015 155.890 77.335 156.220 ;
        RECT 77.515 155.625 78.175 156.105 ;
        RECT 78.375 156.015 78.545 156.775 ;
        RECT 79.445 156.605 79.625 157.015 ;
        RECT 78.715 156.435 79.045 156.555 ;
        RECT 79.795 156.435 79.965 157.195 ;
        RECT 78.715 156.265 79.965 156.435 ;
        RECT 80.135 157.375 81.505 157.625 ;
        RECT 80.135 156.605 80.325 157.375 ;
        RECT 81.255 157.115 81.505 157.375 ;
        RECT 80.495 156.945 80.745 157.105 ;
        RECT 81.675 156.945 81.845 157.790 ;
        RECT 82.740 157.505 82.910 158.005 ;
        RECT 83.080 157.675 83.410 158.175 ;
        RECT 82.015 157.115 82.515 157.495 ;
        RECT 82.740 157.335 83.435 157.505 ;
        RECT 80.495 156.775 81.845 156.945 ;
        RECT 81.425 156.735 81.845 156.775 ;
        RECT 80.135 156.265 80.555 156.605 ;
        RECT 80.845 156.275 81.255 156.605 ;
        RECT 78.375 155.845 79.225 156.015 ;
        RECT 79.785 155.625 80.105 156.085 ;
        RECT 80.305 155.835 80.555 156.265 ;
        RECT 80.845 155.625 81.255 156.065 ;
        RECT 81.425 156.005 81.595 156.735 ;
        RECT 81.765 156.185 82.115 156.555 ;
        RECT 82.295 156.245 82.515 157.115 ;
        RECT 82.685 156.545 83.095 157.165 ;
        RECT 83.265 156.365 83.435 157.335 ;
        RECT 82.740 156.175 83.435 156.365 ;
        RECT 81.425 155.805 82.440 156.005 ;
        RECT 82.740 155.845 82.910 156.175 ;
        RECT 83.080 155.625 83.410 156.005 ;
        RECT 83.625 155.885 83.850 158.005 ;
        RECT 84.020 157.675 84.350 158.175 ;
        RECT 84.520 157.505 84.690 158.005 ;
        RECT 84.025 157.335 84.690 157.505 ;
        RECT 84.025 156.345 84.255 157.335 ;
        RECT 84.425 156.515 84.775 157.165 ;
        RECT 84.950 157.100 85.220 158.005 ;
        RECT 85.390 157.415 85.720 158.175 ;
        RECT 85.900 157.245 86.070 158.005 ;
        RECT 84.025 156.175 84.690 156.345 ;
        RECT 84.020 155.625 84.350 156.005 ;
        RECT 84.520 155.885 84.690 156.175 ;
        RECT 84.950 156.300 85.120 157.100 ;
        RECT 85.405 157.075 86.070 157.245 ;
        RECT 85.405 156.930 85.575 157.075 ;
        RECT 86.330 157.010 86.620 158.175 ;
        RECT 87.165 157.195 87.420 157.865 ;
        RECT 87.600 157.375 87.885 158.175 ;
        RECT 88.065 157.455 88.395 157.965 ;
        RECT 87.165 157.155 87.345 157.195 ;
        RECT 87.080 156.985 87.345 157.155 ;
        RECT 85.290 156.600 85.575 156.930 ;
        RECT 85.405 156.345 85.575 156.600 ;
        RECT 85.810 156.525 86.140 156.895 ;
        RECT 84.950 155.795 85.210 156.300 ;
        RECT 85.405 156.175 86.070 156.345 ;
        RECT 85.390 155.625 85.720 156.005 ;
        RECT 85.900 155.795 86.070 156.175 ;
        RECT 86.330 155.625 86.620 156.350 ;
        RECT 87.165 156.335 87.345 156.985 ;
        RECT 88.065 156.865 88.315 157.455 ;
        RECT 88.665 157.305 88.835 157.915 ;
        RECT 89.005 157.485 89.335 158.175 ;
        RECT 89.565 157.625 89.805 157.915 ;
        RECT 90.005 157.795 90.425 158.175 ;
        RECT 90.605 157.705 91.235 157.955 ;
        RECT 91.705 157.795 92.035 158.175 ;
        RECT 90.605 157.625 90.775 157.705 ;
        RECT 92.205 157.625 92.375 157.915 ;
        RECT 92.555 157.795 92.935 158.175 ;
        RECT 93.175 157.790 94.005 157.960 ;
        RECT 89.565 157.455 90.775 157.625 ;
        RECT 87.515 156.535 88.315 156.865 ;
        RECT 87.165 155.805 87.420 156.335 ;
        RECT 87.600 155.625 87.885 156.085 ;
        RECT 88.065 155.885 88.315 156.535 ;
        RECT 88.515 157.285 88.835 157.305 ;
        RECT 88.515 157.115 90.435 157.285 ;
        RECT 88.515 156.220 88.705 157.115 ;
        RECT 90.605 156.945 90.775 157.455 ;
        RECT 90.945 157.195 91.465 157.505 ;
        RECT 88.875 156.775 90.775 156.945 ;
        RECT 88.875 156.715 89.205 156.775 ;
        RECT 89.355 156.545 89.685 156.605 ;
        RECT 89.025 156.275 89.685 156.545 ;
        RECT 88.515 155.890 88.835 156.220 ;
        RECT 89.015 155.625 89.675 156.105 ;
        RECT 89.875 156.015 90.045 156.775 ;
        RECT 90.945 156.605 91.125 157.015 ;
        RECT 90.215 156.435 90.545 156.555 ;
        RECT 91.295 156.435 91.465 157.195 ;
        RECT 90.215 156.265 91.465 156.435 ;
        RECT 91.635 157.375 93.005 157.625 ;
        RECT 91.635 156.605 91.825 157.375 ;
        RECT 92.755 157.115 93.005 157.375 ;
        RECT 91.995 156.945 92.245 157.105 ;
        RECT 93.175 156.945 93.345 157.790 ;
        RECT 94.240 157.505 94.410 158.005 ;
        RECT 94.580 157.675 94.910 158.175 ;
        RECT 93.515 157.115 94.015 157.495 ;
        RECT 94.240 157.335 94.935 157.505 ;
        RECT 91.995 156.775 93.345 156.945 ;
        RECT 92.925 156.735 93.345 156.775 ;
        RECT 91.635 156.265 92.055 156.605 ;
        RECT 92.345 156.275 92.755 156.605 ;
        RECT 89.875 155.845 90.725 156.015 ;
        RECT 91.285 155.625 91.605 156.085 ;
        RECT 91.805 155.835 92.055 156.265 ;
        RECT 92.345 155.625 92.755 156.065 ;
        RECT 92.925 156.005 93.095 156.735 ;
        RECT 93.265 156.185 93.615 156.555 ;
        RECT 93.795 156.245 94.015 157.115 ;
        RECT 94.185 156.545 94.595 157.165 ;
        RECT 94.765 156.365 94.935 157.335 ;
        RECT 94.240 156.175 94.935 156.365 ;
        RECT 92.925 155.805 93.940 156.005 ;
        RECT 94.240 155.845 94.410 156.175 ;
        RECT 94.580 155.625 94.910 156.005 ;
        RECT 95.125 155.885 95.350 158.005 ;
        RECT 95.520 157.675 95.850 158.175 ;
        RECT 96.020 157.505 96.190 158.005 ;
        RECT 95.525 157.335 96.190 157.505 ;
        RECT 96.910 157.415 97.425 157.825 ;
        RECT 97.660 157.415 97.830 158.175 ;
        RECT 98.000 157.835 100.030 158.005 ;
        RECT 95.525 156.345 95.755 157.335 ;
        RECT 95.925 156.515 96.275 157.165 ;
        RECT 96.910 156.605 97.250 157.415 ;
        RECT 98.000 157.170 98.170 157.835 ;
        RECT 98.565 157.495 99.690 157.665 ;
        RECT 97.420 156.980 98.170 157.170 ;
        RECT 98.340 157.155 99.350 157.325 ;
        RECT 96.910 156.435 98.140 156.605 ;
        RECT 95.525 156.175 96.190 156.345 ;
        RECT 95.520 155.625 95.850 156.005 ;
        RECT 96.020 155.885 96.190 156.175 ;
        RECT 97.185 155.830 97.430 156.435 ;
        RECT 97.650 155.625 98.160 156.160 ;
        RECT 98.340 155.795 98.530 157.155 ;
        RECT 98.700 156.475 98.975 156.955 ;
        RECT 98.700 156.305 98.980 156.475 ;
        RECT 99.180 156.355 99.350 157.155 ;
        RECT 99.520 156.365 99.690 157.495 ;
        RECT 99.860 156.865 100.030 157.835 ;
        RECT 100.200 157.035 100.370 158.175 ;
        RECT 100.540 157.035 100.875 158.005 ;
        RECT 99.860 156.535 100.055 156.865 ;
        RECT 100.280 156.535 100.535 156.865 ;
        RECT 100.280 156.365 100.450 156.535 ;
        RECT 100.705 156.365 100.875 157.035 ;
        RECT 101.425 157.195 101.680 157.865 ;
        RECT 101.860 157.375 102.145 158.175 ;
        RECT 102.325 157.455 102.655 157.965 ;
        RECT 101.425 156.815 101.605 157.195 ;
        RECT 102.325 156.865 102.575 157.455 ;
        RECT 102.925 157.305 103.095 157.915 ;
        RECT 103.265 157.485 103.595 158.175 ;
        RECT 103.825 157.625 104.065 157.915 ;
        RECT 104.265 157.795 104.685 158.175 ;
        RECT 104.865 157.705 105.495 157.955 ;
        RECT 105.965 157.795 106.295 158.175 ;
        RECT 104.865 157.625 105.035 157.705 ;
        RECT 106.465 157.625 106.635 157.915 ;
        RECT 106.815 157.795 107.195 158.175 ;
        RECT 107.435 157.790 108.265 157.960 ;
        RECT 103.825 157.455 105.035 157.625 ;
        RECT 101.340 156.645 101.605 156.815 ;
        RECT 98.700 155.795 98.975 156.305 ;
        RECT 99.520 156.195 100.450 156.365 ;
        RECT 99.520 156.160 99.695 156.195 ;
        RECT 99.165 155.795 99.695 156.160 ;
        RECT 100.120 155.625 100.450 156.025 ;
        RECT 100.620 155.795 100.875 156.365 ;
        RECT 101.425 156.335 101.605 156.645 ;
        RECT 101.775 156.535 102.575 156.865 ;
        RECT 101.425 155.805 101.680 156.335 ;
        RECT 101.860 155.625 102.145 156.085 ;
        RECT 102.325 155.885 102.575 156.535 ;
        RECT 102.775 157.285 103.095 157.305 ;
        RECT 102.775 157.115 104.695 157.285 ;
        RECT 102.775 156.220 102.965 157.115 ;
        RECT 104.865 156.945 105.035 157.455 ;
        RECT 105.205 157.195 105.725 157.505 ;
        RECT 103.135 156.775 105.035 156.945 ;
        RECT 103.135 156.715 103.465 156.775 ;
        RECT 103.615 156.545 103.945 156.605 ;
        RECT 103.285 156.275 103.945 156.545 ;
        RECT 102.775 155.890 103.095 156.220 ;
        RECT 103.275 155.625 103.935 156.105 ;
        RECT 104.135 156.015 104.305 156.775 ;
        RECT 105.205 156.605 105.385 157.015 ;
        RECT 104.475 156.435 104.805 156.555 ;
        RECT 105.555 156.435 105.725 157.195 ;
        RECT 104.475 156.265 105.725 156.435 ;
        RECT 105.895 157.375 107.265 157.625 ;
        RECT 105.895 156.605 106.085 157.375 ;
        RECT 107.015 157.115 107.265 157.375 ;
        RECT 106.255 156.945 106.505 157.105 ;
        RECT 107.435 156.945 107.605 157.790 ;
        RECT 108.500 157.505 108.670 158.005 ;
        RECT 108.840 157.675 109.170 158.175 ;
        RECT 107.775 157.115 108.275 157.495 ;
        RECT 108.500 157.335 109.195 157.505 ;
        RECT 106.255 156.775 107.605 156.945 ;
        RECT 107.185 156.735 107.605 156.775 ;
        RECT 105.895 156.265 106.315 156.605 ;
        RECT 106.605 156.275 107.015 156.605 ;
        RECT 104.135 155.845 104.985 156.015 ;
        RECT 105.545 155.625 105.865 156.085 ;
        RECT 106.065 155.835 106.315 156.265 ;
        RECT 106.605 155.625 107.015 156.065 ;
        RECT 107.185 156.005 107.355 156.735 ;
        RECT 107.525 156.185 107.875 156.555 ;
        RECT 108.055 156.245 108.275 157.115 ;
        RECT 108.445 156.545 108.855 157.165 ;
        RECT 109.025 156.365 109.195 157.335 ;
        RECT 108.500 156.175 109.195 156.365 ;
        RECT 107.185 155.805 108.200 156.005 ;
        RECT 108.500 155.845 108.670 156.175 ;
        RECT 108.840 155.625 109.170 156.005 ;
        RECT 109.385 155.885 109.610 158.005 ;
        RECT 109.780 157.675 110.110 158.175 ;
        RECT 110.280 157.505 110.450 158.005 ;
        RECT 109.785 157.335 110.450 157.505 ;
        RECT 109.785 156.345 110.015 157.335 ;
        RECT 110.185 156.515 110.535 157.165 ;
        RECT 111.170 157.085 112.380 158.175 ;
        RECT 111.170 156.545 111.690 157.085 ;
        RECT 111.860 156.375 112.380 156.915 ;
        RECT 109.785 156.175 110.450 156.345 ;
        RECT 109.780 155.625 110.110 156.005 ;
        RECT 110.280 155.885 110.450 156.175 ;
        RECT 111.170 155.625 112.380 156.375 ;
        RECT 18.165 155.455 112.465 155.625 ;
        RECT 18.250 154.705 19.460 155.455 ;
        RECT 18.250 154.165 18.770 154.705 ;
        RECT 20.090 154.685 21.760 155.455 ;
        RECT 21.930 154.730 22.220 155.455 ;
        RECT 22.940 154.905 23.110 155.285 ;
        RECT 23.290 155.075 23.620 155.455 ;
        RECT 22.940 154.735 23.605 154.905 ;
        RECT 23.800 154.780 24.060 155.285 ;
        RECT 18.940 153.995 19.460 154.535 ;
        RECT 18.250 152.905 19.460 153.995 ;
        RECT 20.090 153.995 20.840 154.515 ;
        RECT 21.010 154.165 21.760 154.685 ;
        RECT 22.870 154.185 23.200 154.555 ;
        RECT 23.435 154.480 23.605 154.735 ;
        RECT 23.435 154.150 23.720 154.480 ;
        RECT 20.090 152.905 21.760 153.995 ;
        RECT 21.930 152.905 22.220 154.070 ;
        RECT 23.435 154.005 23.605 154.150 ;
        RECT 22.940 153.835 23.605 154.005 ;
        RECT 23.890 153.980 24.060 154.780 ;
        RECT 22.940 153.075 23.110 153.835 ;
        RECT 23.290 152.905 23.620 153.665 ;
        RECT 23.790 153.075 24.060 153.980 ;
        RECT 24.235 154.715 24.490 155.285 ;
        RECT 24.660 155.055 24.990 155.455 ;
        RECT 25.415 154.920 25.945 155.285 ;
        RECT 25.415 154.885 25.590 154.920 ;
        RECT 24.660 154.715 25.590 154.885 ;
        RECT 26.135 154.775 26.410 155.285 ;
        RECT 24.235 154.045 24.405 154.715 ;
        RECT 24.660 154.545 24.830 154.715 ;
        RECT 24.575 154.215 24.830 154.545 ;
        RECT 25.055 154.215 25.250 154.545 ;
        RECT 24.235 153.075 24.570 154.045 ;
        RECT 24.740 152.905 24.910 154.045 ;
        RECT 25.080 153.245 25.250 154.215 ;
        RECT 25.420 153.585 25.590 154.715 ;
        RECT 25.760 153.925 25.930 154.725 ;
        RECT 26.130 154.605 26.410 154.775 ;
        RECT 26.135 154.125 26.410 154.605 ;
        RECT 26.580 153.925 26.770 155.285 ;
        RECT 26.950 154.920 27.460 155.455 ;
        RECT 27.680 154.645 27.925 155.250 ;
        RECT 28.370 154.685 30.040 155.455 ;
        RECT 30.300 154.975 30.600 155.455 ;
        RECT 30.770 154.805 31.030 155.260 ;
        RECT 31.200 154.975 31.460 155.455 ;
        RECT 31.640 154.805 31.900 155.260 ;
        RECT 32.070 154.975 32.320 155.455 ;
        RECT 32.500 154.805 32.760 155.260 ;
        RECT 32.930 154.975 33.180 155.455 ;
        RECT 33.360 154.805 33.620 155.260 ;
        RECT 33.790 154.975 34.035 155.455 ;
        RECT 34.205 154.805 34.480 155.260 ;
        RECT 34.650 154.975 34.895 155.455 ;
        RECT 35.065 154.805 35.325 155.260 ;
        RECT 35.495 154.975 35.755 155.455 ;
        RECT 35.925 154.805 36.185 155.260 ;
        RECT 36.355 154.975 36.615 155.455 ;
        RECT 36.785 154.805 37.045 155.260 ;
        RECT 37.215 154.895 37.475 155.455 ;
        RECT 26.970 154.475 28.200 154.645 ;
        RECT 25.760 153.755 26.770 153.925 ;
        RECT 26.940 153.910 27.690 154.100 ;
        RECT 25.420 153.415 26.545 153.585 ;
        RECT 26.940 153.245 27.110 153.910 ;
        RECT 27.860 153.665 28.200 154.475 ;
        RECT 25.080 153.075 27.110 153.245 ;
        RECT 27.280 152.905 27.450 153.665 ;
        RECT 27.685 153.255 28.200 153.665 ;
        RECT 28.370 153.995 29.120 154.515 ;
        RECT 29.290 154.165 30.040 154.685 ;
        RECT 30.300 154.635 37.045 154.805 ;
        RECT 30.300 154.045 31.465 154.635 ;
        RECT 37.645 154.465 37.895 155.275 ;
        RECT 38.075 154.930 38.335 155.455 ;
        RECT 38.505 154.465 38.755 155.275 ;
        RECT 38.935 154.945 39.240 155.455 ;
        RECT 31.635 154.215 38.755 154.465 ;
        RECT 38.925 154.215 39.240 154.775 ;
        RECT 39.870 154.685 41.540 155.455 ;
        RECT 28.370 152.905 30.040 153.995 ;
        RECT 30.300 153.820 37.045 154.045 ;
        RECT 30.300 152.905 30.570 153.650 ;
        RECT 30.740 153.080 31.030 153.820 ;
        RECT 31.640 153.805 37.045 153.820 ;
        RECT 31.200 152.910 31.455 153.635 ;
        RECT 31.640 153.080 31.900 153.805 ;
        RECT 32.070 152.910 32.315 153.635 ;
        RECT 32.500 153.080 32.760 153.805 ;
        RECT 32.930 152.910 33.175 153.635 ;
        RECT 33.360 153.080 33.620 153.805 ;
        RECT 33.790 152.910 34.035 153.635 ;
        RECT 34.205 153.080 34.465 153.805 ;
        RECT 34.635 152.910 34.895 153.635 ;
        RECT 35.065 153.080 35.325 153.805 ;
        RECT 35.495 152.910 35.755 153.635 ;
        RECT 35.925 153.080 36.185 153.805 ;
        RECT 36.355 152.910 36.615 153.635 ;
        RECT 36.785 153.080 37.045 153.805 ;
        RECT 37.215 152.910 37.475 153.705 ;
        RECT 37.645 153.080 37.895 154.215 ;
        RECT 31.200 152.905 37.475 152.910 ;
        RECT 38.075 152.905 38.335 153.715 ;
        RECT 38.510 153.075 38.755 154.215 ;
        RECT 39.870 153.995 40.620 154.515 ;
        RECT 40.790 154.165 41.540 154.685 ;
        RECT 41.710 154.655 42.050 155.285 ;
        RECT 42.220 154.655 42.470 155.455 ;
        RECT 42.660 154.805 42.990 155.285 ;
        RECT 43.160 154.995 43.385 155.455 ;
        RECT 43.555 154.805 43.885 155.285 ;
        RECT 41.710 154.045 41.885 154.655 ;
        RECT 42.660 154.635 43.885 154.805 ;
        RECT 44.515 154.675 45.015 155.285 ;
        RECT 45.850 154.685 47.520 155.455 ;
        RECT 47.690 154.730 47.980 155.455 ;
        RECT 42.055 154.295 42.750 154.465 ;
        RECT 42.580 154.045 42.750 154.295 ;
        RECT 42.925 154.265 43.345 154.465 ;
        RECT 43.515 154.265 43.845 154.465 ;
        RECT 44.015 154.265 44.345 154.465 ;
        RECT 44.515 154.045 44.685 154.675 ;
        RECT 44.870 154.215 45.220 154.465 ;
        RECT 38.935 152.905 39.230 153.715 ;
        RECT 39.870 152.905 41.540 153.995 ;
        RECT 41.710 153.075 42.050 154.045 ;
        RECT 42.220 152.905 42.390 154.045 ;
        RECT 42.580 153.875 45.015 154.045 ;
        RECT 42.660 152.905 42.910 153.705 ;
        RECT 43.555 153.075 43.885 153.875 ;
        RECT 44.185 152.905 44.515 153.705 ;
        RECT 44.685 153.075 45.015 153.875 ;
        RECT 45.850 153.995 46.600 154.515 ;
        RECT 46.770 154.165 47.520 154.685 ;
        RECT 48.150 154.655 48.490 155.285 ;
        RECT 48.660 154.655 48.910 155.455 ;
        RECT 49.100 154.805 49.430 155.285 ;
        RECT 49.600 154.995 49.825 155.455 ;
        RECT 49.995 154.805 50.325 155.285 ;
        RECT 45.850 152.905 47.520 153.995 ;
        RECT 47.690 152.905 47.980 154.070 ;
        RECT 48.150 154.045 48.325 154.655 ;
        RECT 49.100 154.635 50.325 154.805 ;
        RECT 50.955 154.675 51.455 155.285 ;
        RECT 51.830 154.705 53.040 155.455 ;
        RECT 48.495 154.295 49.190 154.465 ;
        RECT 49.020 154.045 49.190 154.295 ;
        RECT 49.365 154.265 49.785 154.465 ;
        RECT 49.955 154.265 50.285 154.465 ;
        RECT 50.455 154.265 50.785 154.465 ;
        RECT 50.955 154.045 51.125 154.675 ;
        RECT 51.310 154.215 51.660 154.465 ;
        RECT 48.150 153.075 48.490 154.045 ;
        RECT 48.660 152.905 48.830 154.045 ;
        RECT 49.020 153.875 51.455 154.045 ;
        RECT 49.100 152.905 49.350 153.705 ;
        RECT 49.995 153.075 50.325 153.875 ;
        RECT 50.625 152.905 50.955 153.705 ;
        RECT 51.125 153.075 51.455 153.875 ;
        RECT 51.830 153.995 52.350 154.535 ;
        RECT 52.520 154.165 53.040 154.705 ;
        RECT 53.585 154.745 53.840 155.275 ;
        RECT 54.020 154.995 54.305 155.455 ;
        RECT 51.830 152.905 53.040 153.995 ;
        RECT 53.585 153.885 53.765 154.745 ;
        RECT 54.485 154.545 54.735 155.195 ;
        RECT 53.935 154.215 54.735 154.545 ;
        RECT 53.585 153.415 53.840 153.885 ;
        RECT 53.500 153.245 53.840 153.415 ;
        RECT 53.585 153.215 53.840 153.245 ;
        RECT 54.020 152.905 54.305 153.705 ;
        RECT 54.485 153.625 54.735 154.215 ;
        RECT 54.935 154.860 55.255 155.190 ;
        RECT 55.435 154.975 56.095 155.455 ;
        RECT 56.295 155.065 57.145 155.235 ;
        RECT 54.935 153.965 55.125 154.860 ;
        RECT 55.445 154.535 56.105 154.805 ;
        RECT 55.775 154.475 56.105 154.535 ;
        RECT 55.295 154.305 55.625 154.365 ;
        RECT 56.295 154.305 56.465 155.065 ;
        RECT 57.705 154.995 58.025 155.455 ;
        RECT 58.225 154.815 58.475 155.245 ;
        RECT 58.765 155.015 59.175 155.455 ;
        RECT 59.345 155.075 60.360 155.275 ;
        RECT 56.635 154.645 57.885 154.815 ;
        RECT 56.635 154.525 56.965 154.645 ;
        RECT 55.295 154.135 57.195 154.305 ;
        RECT 54.935 153.795 56.855 153.965 ;
        RECT 54.935 153.775 55.255 153.795 ;
        RECT 54.485 153.115 54.815 153.625 ;
        RECT 55.085 153.165 55.255 153.775 ;
        RECT 57.025 153.625 57.195 154.135 ;
        RECT 57.365 154.065 57.545 154.475 ;
        RECT 57.715 153.885 57.885 154.645 ;
        RECT 55.425 152.905 55.755 153.595 ;
        RECT 55.985 153.455 57.195 153.625 ;
        RECT 57.365 153.575 57.885 153.885 ;
        RECT 58.055 154.475 58.475 154.815 ;
        RECT 58.765 154.475 59.175 154.805 ;
        RECT 58.055 153.705 58.245 154.475 ;
        RECT 59.345 154.345 59.515 155.075 ;
        RECT 60.660 154.905 60.830 155.235 ;
        RECT 61.000 155.075 61.330 155.455 ;
        RECT 59.685 154.525 60.035 154.895 ;
        RECT 59.345 154.305 59.765 154.345 ;
        RECT 58.415 154.135 59.765 154.305 ;
        RECT 58.415 153.975 58.665 154.135 ;
        RECT 59.175 153.705 59.425 153.965 ;
        RECT 58.055 153.455 59.425 153.705 ;
        RECT 55.985 153.165 56.225 153.455 ;
        RECT 57.025 153.375 57.195 153.455 ;
        RECT 56.425 152.905 56.845 153.285 ;
        RECT 57.025 153.125 57.655 153.375 ;
        RECT 58.125 152.905 58.455 153.285 ;
        RECT 58.625 153.165 58.795 153.455 ;
        RECT 59.595 153.290 59.765 154.135 ;
        RECT 60.215 153.965 60.435 154.835 ;
        RECT 60.660 154.715 61.355 154.905 ;
        RECT 59.935 153.585 60.435 153.965 ;
        RECT 60.605 153.915 61.015 154.535 ;
        RECT 61.185 153.745 61.355 154.715 ;
        RECT 60.660 153.575 61.355 153.745 ;
        RECT 58.975 152.905 59.355 153.285 ;
        RECT 59.595 153.120 60.425 153.290 ;
        RECT 60.660 153.075 60.830 153.575 ;
        RECT 61.000 152.905 61.330 153.405 ;
        RECT 61.545 153.075 61.770 155.195 ;
        RECT 61.940 155.075 62.270 155.455 ;
        RECT 62.440 154.905 62.610 155.195 ;
        RECT 61.945 154.735 62.610 154.905 ;
        RECT 62.960 154.905 63.130 155.285 ;
        RECT 63.310 155.075 63.640 155.455 ;
        RECT 62.960 154.735 63.625 154.905 ;
        RECT 63.820 154.780 64.080 155.285 ;
        RECT 61.945 153.745 62.175 154.735 ;
        RECT 62.345 153.915 62.695 154.565 ;
        RECT 62.890 154.185 63.220 154.555 ;
        RECT 63.455 154.480 63.625 154.735 ;
        RECT 63.455 154.150 63.740 154.480 ;
        RECT 63.455 154.005 63.625 154.150 ;
        RECT 62.960 153.835 63.625 154.005 ;
        RECT 63.910 153.980 64.080 154.780 ;
        RECT 64.255 154.615 64.515 155.455 ;
        RECT 64.690 154.710 64.945 155.285 ;
        RECT 65.115 155.075 65.445 155.455 ;
        RECT 65.660 154.905 65.830 155.285 ;
        RECT 65.115 154.735 65.830 154.905 ;
        RECT 61.945 153.575 62.610 153.745 ;
        RECT 61.940 152.905 62.270 153.405 ;
        RECT 62.440 153.075 62.610 153.575 ;
        RECT 62.960 153.075 63.130 153.835 ;
        RECT 63.310 152.905 63.640 153.665 ;
        RECT 63.810 153.075 64.080 153.980 ;
        RECT 64.255 152.905 64.515 154.055 ;
        RECT 64.690 153.980 64.860 154.710 ;
        RECT 65.115 154.545 65.285 154.735 ;
        RECT 66.295 154.675 66.795 155.285 ;
        RECT 65.030 154.215 65.285 154.545 ;
        RECT 65.115 154.005 65.285 154.215 ;
        RECT 65.565 154.185 65.920 154.555 ;
        RECT 66.090 154.215 66.440 154.465 ;
        RECT 66.625 154.045 66.795 154.675 ;
        RECT 67.425 154.805 67.755 155.285 ;
        RECT 67.925 154.995 68.150 155.455 ;
        RECT 68.320 154.805 68.650 155.285 ;
        RECT 67.425 154.635 68.650 154.805 ;
        RECT 68.840 154.655 69.090 155.455 ;
        RECT 69.260 154.655 69.600 155.285 ;
        RECT 69.975 154.675 70.475 155.285 ;
        RECT 66.965 154.265 67.295 154.465 ;
        RECT 67.465 154.265 67.795 154.465 ;
        RECT 67.965 154.265 68.385 154.465 ;
        RECT 68.560 154.295 69.255 154.465 ;
        RECT 68.560 154.045 68.730 154.295 ;
        RECT 69.425 154.045 69.600 154.655 ;
        RECT 69.770 154.215 70.120 154.465 ;
        RECT 70.305 154.045 70.475 154.675 ;
        RECT 71.105 154.805 71.435 155.285 ;
        RECT 71.605 154.995 71.830 155.455 ;
        RECT 72.000 154.805 72.330 155.285 ;
        RECT 71.105 154.635 72.330 154.805 ;
        RECT 72.520 154.655 72.770 155.455 ;
        RECT 72.940 154.655 73.280 155.285 ;
        RECT 73.450 154.730 73.740 155.455 ;
        RECT 73.970 154.975 74.250 155.455 ;
        RECT 74.420 154.805 74.680 155.195 ;
        RECT 74.855 154.975 75.110 155.455 ;
        RECT 75.280 154.805 75.575 155.195 ;
        RECT 75.755 154.975 76.030 155.455 ;
        RECT 76.200 154.955 76.500 155.285 ;
        RECT 70.645 154.265 70.975 154.465 ;
        RECT 71.145 154.265 71.475 154.465 ;
        RECT 71.645 154.265 72.065 154.465 ;
        RECT 72.240 154.295 72.935 154.465 ;
        RECT 72.240 154.045 72.410 154.295 ;
        RECT 73.105 154.045 73.280 154.655 ;
        RECT 73.925 154.635 75.575 154.805 ;
        RECT 73.925 154.125 74.330 154.635 ;
        RECT 74.500 154.295 75.640 154.465 ;
        RECT 64.690 153.075 64.945 153.980 ;
        RECT 65.115 153.835 65.830 154.005 ;
        RECT 65.115 152.905 65.445 153.665 ;
        RECT 65.660 153.075 65.830 153.835 ;
        RECT 66.295 153.875 68.730 154.045 ;
        RECT 66.295 153.075 66.625 153.875 ;
        RECT 66.795 152.905 67.125 153.705 ;
        RECT 67.425 153.075 67.755 153.875 ;
        RECT 68.400 152.905 68.650 153.705 ;
        RECT 68.920 152.905 69.090 154.045 ;
        RECT 69.260 153.075 69.600 154.045 ;
        RECT 69.975 153.875 72.410 154.045 ;
        RECT 69.975 153.075 70.305 153.875 ;
        RECT 70.475 152.905 70.805 153.705 ;
        RECT 71.105 153.075 71.435 153.875 ;
        RECT 72.080 152.905 72.330 153.705 ;
        RECT 72.600 152.905 72.770 154.045 ;
        RECT 72.940 153.075 73.280 154.045 ;
        RECT 73.450 152.905 73.740 154.070 ;
        RECT 73.925 153.955 74.680 154.125 ;
        RECT 73.965 152.905 74.250 153.775 ;
        RECT 74.420 153.705 74.680 153.955 ;
        RECT 75.470 154.045 75.640 154.295 ;
        RECT 75.810 154.215 76.160 154.785 ;
        RECT 76.330 154.045 76.500 154.955 ;
        RECT 76.945 154.645 77.190 155.250 ;
        RECT 77.410 154.920 77.920 155.455 ;
        RECT 75.470 153.875 76.500 154.045 ;
        RECT 74.420 153.535 75.540 153.705 ;
        RECT 74.420 153.075 74.680 153.535 ;
        RECT 74.855 152.905 75.110 153.365 ;
        RECT 75.280 153.075 75.540 153.535 ;
        RECT 75.710 152.905 76.020 153.705 ;
        RECT 76.190 153.075 76.500 153.875 ;
        RECT 76.670 154.475 77.900 154.645 ;
        RECT 76.670 153.665 77.010 154.475 ;
        RECT 77.180 153.910 77.930 154.100 ;
        RECT 76.670 153.255 77.185 153.665 ;
        RECT 77.420 152.905 77.590 153.665 ;
        RECT 77.760 153.245 77.930 153.910 ;
        RECT 78.100 153.925 78.290 155.285 ;
        RECT 78.460 154.435 78.735 155.285 ;
        RECT 78.925 154.920 79.455 155.285 ;
        RECT 79.880 155.055 80.210 155.455 ;
        RECT 79.280 154.885 79.455 154.920 ;
        RECT 78.460 154.265 78.740 154.435 ;
        RECT 78.460 154.125 78.735 154.265 ;
        RECT 78.940 153.925 79.110 154.725 ;
        RECT 78.100 153.755 79.110 153.925 ;
        RECT 79.280 154.715 80.210 154.885 ;
        RECT 80.380 154.715 80.635 155.285 ;
        RECT 81.730 154.945 82.035 155.455 ;
        RECT 79.280 153.585 79.450 154.715 ;
        RECT 80.040 154.545 80.210 154.715 ;
        RECT 78.325 153.415 79.450 153.585 ;
        RECT 79.620 154.215 79.815 154.545 ;
        RECT 80.040 154.215 80.295 154.545 ;
        RECT 79.620 153.245 79.790 154.215 ;
        RECT 80.465 154.045 80.635 154.715 ;
        RECT 81.730 154.215 82.045 154.775 ;
        RECT 82.215 154.465 82.465 155.275 ;
        RECT 82.635 154.930 82.895 155.455 ;
        RECT 83.075 154.465 83.325 155.275 ;
        RECT 83.495 154.895 83.755 155.455 ;
        RECT 83.925 154.805 84.185 155.260 ;
        RECT 84.355 154.975 84.615 155.455 ;
        RECT 84.785 154.805 85.045 155.260 ;
        RECT 85.215 154.975 85.475 155.455 ;
        RECT 85.645 154.805 85.905 155.260 ;
        RECT 86.075 154.975 86.320 155.455 ;
        RECT 86.490 154.805 86.765 155.260 ;
        RECT 86.935 154.975 87.180 155.455 ;
        RECT 87.350 154.805 87.610 155.260 ;
        RECT 87.790 154.975 88.040 155.455 ;
        RECT 88.210 154.805 88.470 155.260 ;
        RECT 88.650 154.975 88.900 155.455 ;
        RECT 89.070 154.805 89.330 155.260 ;
        RECT 89.510 154.975 89.770 155.455 ;
        RECT 89.940 154.805 90.200 155.260 ;
        RECT 90.370 154.975 90.670 155.455 ;
        RECT 83.925 154.635 90.670 154.805 ;
        RECT 82.215 154.215 89.335 154.465 ;
        RECT 77.760 153.075 79.790 153.245 ;
        RECT 79.960 152.905 80.130 154.045 ;
        RECT 80.300 153.075 80.635 154.045 ;
        RECT 81.740 152.905 82.035 153.715 ;
        RECT 82.215 153.075 82.460 154.215 ;
        RECT 82.635 152.905 82.895 153.715 ;
        RECT 83.075 153.080 83.325 154.215 ;
        RECT 89.505 154.045 90.670 154.635 ;
        RECT 83.925 153.820 90.670 154.045 ;
        RECT 90.930 154.655 91.270 155.285 ;
        RECT 91.440 154.655 91.690 155.455 ;
        RECT 91.880 154.805 92.210 155.285 ;
        RECT 92.380 154.995 92.605 155.455 ;
        RECT 92.775 154.805 93.105 155.285 ;
        RECT 90.930 154.045 91.105 154.655 ;
        RECT 91.880 154.635 93.105 154.805 ;
        RECT 93.735 154.675 94.235 155.285 ;
        RECT 95.735 154.675 96.235 155.285 ;
        RECT 91.275 154.295 91.970 154.465 ;
        RECT 91.800 154.045 91.970 154.295 ;
        RECT 92.145 154.265 92.565 154.465 ;
        RECT 92.735 154.265 93.065 154.465 ;
        RECT 93.235 154.265 93.565 154.465 ;
        RECT 93.735 154.045 93.905 154.675 ;
        RECT 94.090 154.215 94.440 154.465 ;
        RECT 95.530 154.215 95.880 154.465 ;
        RECT 96.065 154.045 96.235 154.675 ;
        RECT 96.865 154.805 97.195 155.285 ;
        RECT 97.365 154.995 97.590 155.455 ;
        RECT 97.760 154.805 98.090 155.285 ;
        RECT 96.865 154.635 98.090 154.805 ;
        RECT 98.280 154.655 98.530 155.455 ;
        RECT 98.700 154.655 99.040 155.285 ;
        RECT 99.210 154.730 99.500 155.455 ;
        RECT 99.875 154.675 100.375 155.285 ;
        RECT 98.810 154.605 99.040 154.655 ;
        RECT 96.405 154.265 96.735 154.465 ;
        RECT 96.905 154.265 97.235 154.465 ;
        RECT 97.405 154.265 97.825 154.465 ;
        RECT 98.000 154.295 98.695 154.465 ;
        RECT 98.000 154.045 98.170 154.295 ;
        RECT 98.865 154.045 99.040 154.605 ;
        RECT 99.670 154.215 100.020 154.465 ;
        RECT 83.925 153.805 89.330 153.820 ;
        RECT 83.495 152.910 83.755 153.705 ;
        RECT 83.925 153.080 84.185 153.805 ;
        RECT 84.355 152.910 84.615 153.635 ;
        RECT 84.785 153.080 85.045 153.805 ;
        RECT 85.215 152.910 85.475 153.635 ;
        RECT 85.645 153.080 85.905 153.805 ;
        RECT 86.075 152.910 86.335 153.635 ;
        RECT 86.505 153.080 86.765 153.805 ;
        RECT 86.935 152.910 87.180 153.635 ;
        RECT 87.350 153.080 87.610 153.805 ;
        RECT 87.795 152.910 88.040 153.635 ;
        RECT 88.210 153.080 88.470 153.805 ;
        RECT 88.655 152.910 88.900 153.635 ;
        RECT 89.070 153.080 89.330 153.805 ;
        RECT 89.515 152.910 89.770 153.635 ;
        RECT 89.940 153.080 90.230 153.820 ;
        RECT 83.495 152.905 89.770 152.910 ;
        RECT 90.400 152.905 90.670 153.650 ;
        RECT 90.930 153.075 91.270 154.045 ;
        RECT 91.440 152.905 91.610 154.045 ;
        RECT 91.800 153.875 94.235 154.045 ;
        RECT 91.880 152.905 92.130 153.705 ;
        RECT 92.775 153.075 93.105 153.875 ;
        RECT 93.405 152.905 93.735 153.705 ;
        RECT 93.905 153.075 94.235 153.875 ;
        RECT 95.735 153.875 98.170 154.045 ;
        RECT 95.735 153.075 96.065 153.875 ;
        RECT 96.235 152.905 96.565 153.705 ;
        RECT 96.865 153.075 97.195 153.875 ;
        RECT 97.840 152.905 98.090 153.705 ;
        RECT 98.360 152.905 98.530 154.045 ;
        RECT 98.700 153.075 99.040 154.045 ;
        RECT 99.210 152.905 99.500 154.070 ;
        RECT 100.205 154.045 100.375 154.675 ;
        RECT 101.005 154.805 101.335 155.285 ;
        RECT 101.505 154.995 101.730 155.455 ;
        RECT 101.900 154.805 102.230 155.285 ;
        RECT 101.005 154.635 102.230 154.805 ;
        RECT 102.420 154.655 102.670 155.455 ;
        RECT 102.840 154.655 103.180 155.285 ;
        RECT 103.500 154.655 103.830 155.455 ;
        RECT 104.000 154.805 104.170 155.285 ;
        RECT 104.340 154.975 104.670 155.455 ;
        RECT 104.840 154.805 105.010 155.285 ;
        RECT 105.260 154.975 105.500 155.455 ;
        RECT 105.680 154.805 105.850 155.285 ;
        RECT 100.545 154.265 100.875 154.465 ;
        RECT 101.045 154.265 101.375 154.465 ;
        RECT 101.545 154.265 101.965 154.465 ;
        RECT 102.140 154.295 102.835 154.465 ;
        RECT 102.140 154.045 102.310 154.295 ;
        RECT 103.005 154.045 103.180 154.655 ;
        RECT 104.000 154.635 105.010 154.805 ;
        RECT 105.215 154.635 105.850 154.805 ;
        RECT 106.200 154.905 106.370 155.285 ;
        RECT 106.550 155.075 106.880 155.455 ;
        RECT 106.200 154.735 106.865 154.905 ;
        RECT 107.060 154.780 107.320 155.285 ;
        RECT 104.000 154.605 104.500 154.635 ;
        RECT 104.000 154.095 104.495 154.605 ;
        RECT 105.215 154.465 105.385 154.635 ;
        RECT 104.885 154.295 105.385 154.465 ;
        RECT 99.875 153.875 102.310 154.045 ;
        RECT 99.875 153.075 100.205 153.875 ;
        RECT 100.375 152.905 100.705 153.705 ;
        RECT 101.005 153.075 101.335 153.875 ;
        RECT 101.980 152.905 102.230 153.705 ;
        RECT 102.500 152.905 102.670 154.045 ;
        RECT 102.840 153.075 103.180 154.045 ;
        RECT 103.500 152.905 103.830 154.055 ;
        RECT 104.000 153.925 105.010 154.095 ;
        RECT 104.000 153.075 104.170 153.925 ;
        RECT 104.340 152.905 104.670 153.705 ;
        RECT 104.840 153.075 105.010 153.925 ;
        RECT 105.215 154.055 105.385 154.295 ;
        RECT 105.555 154.225 105.935 154.465 ;
        RECT 106.130 154.185 106.460 154.555 ;
        RECT 106.695 154.480 106.865 154.735 ;
        RECT 106.695 154.150 106.980 154.480 ;
        RECT 105.215 153.885 105.930 154.055 ;
        RECT 106.695 154.005 106.865 154.150 ;
        RECT 105.190 152.905 105.430 153.705 ;
        RECT 105.600 153.075 105.930 153.885 ;
        RECT 106.200 153.835 106.865 154.005 ;
        RECT 107.150 153.980 107.320 154.780 ;
        RECT 107.490 154.685 111.000 155.455 ;
        RECT 111.170 154.705 112.380 155.455 ;
        RECT 106.200 153.075 106.370 153.835 ;
        RECT 106.550 152.905 106.880 153.665 ;
        RECT 107.050 153.075 107.320 153.980 ;
        RECT 107.490 153.995 109.180 154.515 ;
        RECT 109.350 154.165 111.000 154.685 ;
        RECT 111.170 153.995 111.690 154.535 ;
        RECT 111.860 154.165 112.380 154.705 ;
        RECT 107.490 152.905 111.000 153.995 ;
        RECT 111.170 152.905 112.380 153.995 ;
        RECT 18.165 152.735 112.465 152.905 ;
        RECT 18.250 151.645 19.460 152.735 ;
        RECT 18.250 150.935 18.770 151.475 ;
        RECT 18.940 151.105 19.460 151.645 ;
        RECT 19.690 151.595 19.900 152.735 ;
        RECT 20.070 151.585 20.400 152.565 ;
        RECT 20.570 151.595 20.800 152.735 ;
        RECT 21.015 152.065 21.270 152.565 ;
        RECT 21.440 152.235 21.770 152.735 ;
        RECT 21.015 151.895 21.765 152.065 ;
        RECT 18.250 150.185 19.460 150.935 ;
        RECT 19.690 150.185 19.900 151.005 ;
        RECT 20.070 150.985 20.320 151.585 ;
        RECT 20.490 151.175 20.820 151.425 ;
        RECT 21.015 151.075 21.365 151.725 ;
        RECT 20.070 150.355 20.400 150.985 ;
        RECT 20.570 150.185 20.800 151.005 ;
        RECT 21.535 150.905 21.765 151.895 ;
        RECT 21.015 150.735 21.765 150.905 ;
        RECT 21.015 150.445 21.270 150.735 ;
        RECT 21.440 150.185 21.770 150.565 ;
        RECT 21.940 150.445 22.110 152.565 ;
        RECT 22.280 151.765 22.605 152.550 ;
        RECT 22.775 152.275 23.025 152.735 ;
        RECT 23.195 152.235 23.445 152.565 ;
        RECT 23.660 152.235 24.340 152.565 ;
        RECT 23.195 152.105 23.365 152.235 ;
        RECT 22.970 151.935 23.365 152.105 ;
        RECT 22.340 150.715 22.800 151.765 ;
        RECT 22.970 150.575 23.140 151.935 ;
        RECT 23.535 151.675 24.000 152.065 ;
        RECT 23.310 150.865 23.660 151.485 ;
        RECT 23.830 151.085 24.000 151.675 ;
        RECT 24.170 151.455 24.340 152.235 ;
        RECT 24.510 152.135 24.680 152.475 ;
        RECT 24.915 152.305 25.245 152.735 ;
        RECT 25.415 152.135 25.585 152.475 ;
        RECT 25.880 152.275 26.250 152.735 ;
        RECT 24.510 151.965 25.585 152.135 ;
        RECT 26.420 152.105 26.590 152.565 ;
        RECT 26.825 152.225 27.695 152.565 ;
        RECT 27.865 152.275 28.115 152.735 ;
        RECT 26.030 151.935 26.590 152.105 ;
        RECT 26.030 151.795 26.200 151.935 ;
        RECT 24.700 151.625 26.200 151.795 ;
        RECT 26.895 151.765 27.355 152.055 ;
        RECT 24.170 151.285 25.860 151.455 ;
        RECT 23.830 150.865 24.185 151.085 ;
        RECT 24.355 150.575 24.525 151.285 ;
        RECT 24.730 150.865 25.520 151.115 ;
        RECT 25.690 151.105 25.860 151.285 ;
        RECT 26.030 150.935 26.200 151.625 ;
        RECT 22.470 150.185 22.800 150.545 ;
        RECT 22.970 150.405 23.465 150.575 ;
        RECT 23.670 150.405 24.525 150.575 ;
        RECT 25.400 150.185 25.730 150.645 ;
        RECT 25.940 150.545 26.200 150.935 ;
        RECT 26.390 151.755 27.355 151.765 ;
        RECT 27.525 151.845 27.695 152.225 ;
        RECT 28.285 152.185 28.455 152.475 ;
        RECT 28.635 152.355 28.965 152.735 ;
        RECT 28.285 152.015 29.085 152.185 ;
        RECT 26.390 151.595 27.065 151.755 ;
        RECT 27.525 151.675 28.745 151.845 ;
        RECT 26.390 150.805 26.600 151.595 ;
        RECT 27.525 151.585 27.695 151.675 ;
        RECT 26.770 150.805 27.120 151.425 ;
        RECT 27.290 151.415 27.695 151.585 ;
        RECT 27.290 150.635 27.460 151.415 ;
        RECT 27.630 150.965 27.850 151.245 ;
        RECT 28.030 151.135 28.570 151.505 ;
        RECT 28.915 151.425 29.085 152.015 ;
        RECT 29.305 151.595 29.610 152.735 ;
        RECT 29.780 151.545 30.035 152.425 ;
        RECT 28.915 151.395 29.655 151.425 ;
        RECT 27.630 150.795 28.160 150.965 ;
        RECT 25.940 150.375 26.290 150.545 ;
        RECT 26.510 150.355 27.460 150.635 ;
        RECT 27.630 150.185 27.820 150.625 ;
        RECT 27.990 150.565 28.160 150.795 ;
        RECT 28.330 150.735 28.570 151.135 ;
        RECT 28.740 151.095 29.655 151.395 ;
        RECT 28.740 150.920 29.065 151.095 ;
        RECT 28.740 150.565 29.060 150.920 ;
        RECT 29.825 150.895 30.035 151.545 ;
        RECT 30.670 151.975 31.185 152.385 ;
        RECT 31.420 151.975 31.590 152.735 ;
        RECT 31.760 152.395 33.790 152.565 ;
        RECT 30.670 151.165 31.010 151.975 ;
        RECT 31.760 151.730 31.930 152.395 ;
        RECT 32.325 152.055 33.450 152.225 ;
        RECT 31.180 151.540 31.930 151.730 ;
        RECT 32.100 151.715 33.110 151.885 ;
        RECT 30.670 150.995 31.900 151.165 ;
        RECT 27.990 150.395 29.060 150.565 ;
        RECT 29.305 150.185 29.610 150.645 ;
        RECT 29.780 150.365 30.035 150.895 ;
        RECT 30.945 150.390 31.190 150.995 ;
        RECT 31.410 150.185 31.920 150.720 ;
        RECT 32.100 150.355 32.290 151.715 ;
        RECT 32.460 151.375 32.735 151.515 ;
        RECT 32.460 151.205 32.740 151.375 ;
        RECT 32.460 150.355 32.735 151.205 ;
        RECT 32.940 150.915 33.110 151.715 ;
        RECT 33.280 150.925 33.450 152.055 ;
        RECT 33.620 151.425 33.790 152.395 ;
        RECT 33.960 151.595 34.130 152.735 ;
        RECT 34.300 151.595 34.635 152.565 ;
        RECT 33.620 151.095 33.815 151.425 ;
        RECT 34.040 151.095 34.295 151.425 ;
        RECT 34.040 150.925 34.210 151.095 ;
        RECT 34.465 150.925 34.635 151.595 ;
        RECT 34.810 151.570 35.100 152.735 ;
        RECT 35.730 151.975 36.245 152.385 ;
        RECT 36.480 151.975 36.650 152.735 ;
        RECT 36.820 152.395 38.850 152.565 ;
        RECT 35.730 151.165 36.070 151.975 ;
        RECT 36.820 151.730 36.990 152.395 ;
        RECT 37.385 152.055 38.510 152.225 ;
        RECT 36.240 151.540 36.990 151.730 ;
        RECT 37.160 151.715 38.170 151.885 ;
        RECT 35.730 150.995 36.960 151.165 ;
        RECT 33.280 150.755 34.210 150.925 ;
        RECT 33.280 150.720 33.455 150.755 ;
        RECT 32.925 150.355 33.455 150.720 ;
        RECT 33.880 150.185 34.210 150.585 ;
        RECT 34.380 150.355 34.635 150.925 ;
        RECT 34.810 150.185 35.100 150.910 ;
        RECT 36.005 150.390 36.250 150.995 ;
        RECT 36.470 150.185 36.980 150.720 ;
        RECT 37.160 150.355 37.350 151.715 ;
        RECT 37.520 151.375 37.795 151.515 ;
        RECT 37.520 151.205 37.800 151.375 ;
        RECT 37.520 150.355 37.795 151.205 ;
        RECT 38.000 150.915 38.170 151.715 ;
        RECT 38.340 150.925 38.510 152.055 ;
        RECT 38.680 151.425 38.850 152.395 ;
        RECT 39.020 151.595 39.190 152.735 ;
        RECT 39.360 151.595 39.695 152.565 ;
        RECT 38.680 151.095 38.875 151.425 ;
        RECT 39.100 151.095 39.355 151.425 ;
        RECT 39.100 150.925 39.270 151.095 ;
        RECT 39.525 150.925 39.695 151.595 ;
        RECT 38.340 150.755 39.270 150.925 ;
        RECT 38.340 150.720 38.515 150.755 ;
        RECT 37.985 150.355 38.515 150.720 ;
        RECT 38.940 150.185 39.270 150.585 ;
        RECT 39.440 150.355 39.695 150.925 ;
        RECT 39.870 151.660 40.140 152.565 ;
        RECT 40.310 151.975 40.640 152.735 ;
        RECT 40.820 151.805 40.990 152.565 ;
        RECT 39.870 150.860 40.040 151.660 ;
        RECT 40.325 151.635 40.990 151.805 ;
        RECT 40.325 151.490 40.495 151.635 ;
        RECT 40.210 151.160 40.495 151.490 ;
        RECT 41.710 151.595 42.050 152.565 ;
        RECT 42.220 151.595 42.390 152.735 ;
        RECT 42.660 151.935 42.910 152.735 ;
        RECT 43.555 151.765 43.885 152.565 ;
        RECT 44.185 151.935 44.515 152.735 ;
        RECT 44.685 151.765 45.015 152.565 ;
        RECT 42.580 151.595 45.015 151.765 ;
        RECT 45.595 151.765 45.925 152.565 ;
        RECT 46.095 151.935 46.425 152.735 ;
        RECT 46.725 151.765 47.055 152.565 ;
        RECT 47.700 151.935 47.950 152.735 ;
        RECT 45.595 151.595 48.030 151.765 ;
        RECT 48.220 151.595 48.390 152.735 ;
        RECT 48.560 151.595 48.900 152.565 ;
        RECT 40.325 150.905 40.495 151.160 ;
        RECT 40.730 151.085 41.060 151.455 ;
        RECT 41.710 150.985 41.885 151.595 ;
        RECT 42.580 151.345 42.750 151.595 ;
        RECT 42.055 151.175 42.750 151.345 ;
        RECT 42.925 151.175 43.345 151.375 ;
        RECT 43.515 151.175 43.845 151.375 ;
        RECT 44.015 151.175 44.345 151.375 ;
        RECT 39.870 150.355 40.130 150.860 ;
        RECT 40.325 150.735 40.990 150.905 ;
        RECT 40.310 150.185 40.640 150.565 ;
        RECT 40.820 150.355 40.990 150.735 ;
        RECT 41.710 150.355 42.050 150.985 ;
        RECT 42.220 150.185 42.470 150.985 ;
        RECT 42.660 150.835 43.885 151.005 ;
        RECT 42.660 150.355 42.990 150.835 ;
        RECT 43.160 150.185 43.385 150.645 ;
        RECT 43.555 150.355 43.885 150.835 ;
        RECT 44.515 150.965 44.685 151.595 ;
        RECT 44.870 151.175 45.220 151.425 ;
        RECT 45.390 151.175 45.740 151.425 ;
        RECT 45.925 150.965 46.095 151.595 ;
        RECT 46.265 151.175 46.595 151.375 ;
        RECT 46.765 151.175 47.095 151.375 ;
        RECT 47.265 151.175 47.685 151.375 ;
        RECT 47.860 151.345 48.030 151.595 ;
        RECT 47.860 151.175 48.555 151.345 ;
        RECT 44.515 150.355 45.015 150.965 ;
        RECT 45.595 150.355 46.095 150.965 ;
        RECT 46.725 150.835 47.950 151.005 ;
        RECT 48.725 150.985 48.900 151.595 ;
        RECT 49.070 151.645 50.740 152.735 ;
        RECT 51.285 151.755 51.540 152.425 ;
        RECT 51.720 151.935 52.005 152.735 ;
        RECT 52.185 152.015 52.515 152.525 ;
        RECT 49.070 151.125 49.820 151.645 ;
        RECT 46.725 150.355 47.055 150.835 ;
        RECT 47.225 150.185 47.450 150.645 ;
        RECT 47.620 150.355 47.950 150.835 ;
        RECT 48.140 150.185 48.390 150.985 ;
        RECT 48.560 150.355 48.900 150.985 ;
        RECT 49.990 150.955 50.740 151.475 ;
        RECT 49.070 150.185 50.740 150.955 ;
        RECT 51.285 150.895 51.465 151.755 ;
        RECT 52.185 151.425 52.435 152.015 ;
        RECT 52.785 151.865 52.955 152.475 ;
        RECT 53.125 152.045 53.455 152.735 ;
        RECT 53.685 152.185 53.925 152.475 ;
        RECT 54.125 152.355 54.545 152.735 ;
        RECT 54.725 152.265 55.355 152.515 ;
        RECT 55.825 152.355 56.155 152.735 ;
        RECT 54.725 152.185 54.895 152.265 ;
        RECT 56.325 152.185 56.495 152.475 ;
        RECT 56.675 152.355 57.055 152.735 ;
        RECT 57.295 152.350 58.125 152.520 ;
        RECT 53.685 152.015 54.895 152.185 ;
        RECT 51.635 151.095 52.435 151.425 ;
        RECT 51.285 150.695 51.540 150.895 ;
        RECT 51.200 150.525 51.540 150.695 ;
        RECT 51.285 150.365 51.540 150.525 ;
        RECT 51.720 150.185 52.005 150.645 ;
        RECT 52.185 150.445 52.435 151.095 ;
        RECT 52.635 151.845 52.955 151.865 ;
        RECT 52.635 151.675 54.555 151.845 ;
        RECT 52.635 150.780 52.825 151.675 ;
        RECT 54.725 151.505 54.895 152.015 ;
        RECT 55.065 151.755 55.585 152.065 ;
        RECT 52.995 151.335 54.895 151.505 ;
        RECT 52.995 151.275 53.325 151.335 ;
        RECT 53.475 151.105 53.805 151.165 ;
        RECT 53.145 150.835 53.805 151.105 ;
        RECT 52.635 150.450 52.955 150.780 ;
        RECT 53.135 150.185 53.795 150.665 ;
        RECT 53.995 150.575 54.165 151.335 ;
        RECT 55.065 151.165 55.245 151.575 ;
        RECT 54.335 150.995 54.665 151.115 ;
        RECT 55.415 150.995 55.585 151.755 ;
        RECT 54.335 150.825 55.585 150.995 ;
        RECT 55.755 151.935 57.125 152.185 ;
        RECT 55.755 151.165 55.945 151.935 ;
        RECT 56.875 151.675 57.125 151.935 ;
        RECT 56.115 151.505 56.365 151.665 ;
        RECT 57.295 151.505 57.465 152.350 ;
        RECT 58.360 152.065 58.530 152.565 ;
        RECT 58.700 152.235 59.030 152.735 ;
        RECT 57.635 151.675 58.135 152.055 ;
        RECT 58.360 151.895 59.055 152.065 ;
        RECT 56.115 151.335 57.465 151.505 ;
        RECT 57.045 151.295 57.465 151.335 ;
        RECT 55.755 150.825 56.175 151.165 ;
        RECT 56.465 150.835 56.875 151.165 ;
        RECT 53.995 150.405 54.845 150.575 ;
        RECT 55.405 150.185 55.725 150.645 ;
        RECT 55.925 150.395 56.175 150.825 ;
        RECT 56.465 150.185 56.875 150.625 ;
        RECT 57.045 150.565 57.215 151.295 ;
        RECT 57.385 150.745 57.735 151.115 ;
        RECT 57.915 150.805 58.135 151.675 ;
        RECT 58.305 151.105 58.715 151.725 ;
        RECT 58.885 150.925 59.055 151.895 ;
        RECT 58.360 150.735 59.055 150.925 ;
        RECT 57.045 150.365 58.060 150.565 ;
        RECT 58.360 150.405 58.530 150.735 ;
        RECT 58.700 150.185 59.030 150.565 ;
        RECT 59.245 150.445 59.470 152.565 ;
        RECT 59.640 152.235 59.970 152.735 ;
        RECT 60.140 152.065 60.310 152.565 ;
        RECT 59.645 151.895 60.310 152.065 ;
        RECT 59.645 150.905 59.875 151.895 ;
        RECT 60.045 151.075 60.395 151.725 ;
        RECT 60.570 151.570 60.860 152.735 ;
        RECT 61.030 151.660 61.300 152.565 ;
        RECT 61.470 151.975 61.800 152.735 ;
        RECT 61.980 151.805 62.150 152.565 ;
        RECT 59.645 150.735 60.310 150.905 ;
        RECT 59.640 150.185 59.970 150.565 ;
        RECT 60.140 150.445 60.310 150.735 ;
        RECT 60.570 150.185 60.860 150.910 ;
        RECT 61.030 150.860 61.200 151.660 ;
        RECT 61.485 151.635 62.150 151.805 ;
        RECT 61.485 151.490 61.655 151.635 ;
        RECT 62.470 151.595 62.680 152.735 ;
        RECT 61.370 151.160 61.655 151.490 ;
        RECT 62.850 151.585 63.180 152.565 ;
        RECT 63.350 151.595 63.580 152.735 ;
        RECT 64.340 151.805 64.510 152.565 ;
        RECT 64.725 151.975 65.055 152.735 ;
        RECT 64.340 151.635 65.055 151.805 ;
        RECT 65.225 151.660 65.480 152.565 ;
        RECT 61.485 150.905 61.655 151.160 ;
        RECT 61.890 151.085 62.220 151.455 ;
        RECT 61.030 150.355 61.290 150.860 ;
        RECT 61.485 150.735 62.150 150.905 ;
        RECT 61.470 150.185 61.800 150.565 ;
        RECT 61.980 150.355 62.150 150.735 ;
        RECT 62.470 150.185 62.680 151.005 ;
        RECT 62.850 150.985 63.100 151.585 ;
        RECT 63.270 151.175 63.600 151.425 ;
        RECT 64.250 151.085 64.605 151.455 ;
        RECT 64.885 151.425 65.055 151.635 ;
        RECT 64.885 151.095 65.140 151.425 ;
        RECT 62.850 150.355 63.180 150.985 ;
        RECT 63.350 150.185 63.580 151.005 ;
        RECT 64.885 150.905 65.055 151.095 ;
        RECT 65.310 150.930 65.480 151.660 ;
        RECT 65.655 151.585 65.915 152.735 ;
        RECT 66.180 151.805 66.350 152.565 ;
        RECT 66.565 151.975 66.895 152.735 ;
        RECT 66.180 151.635 66.895 151.805 ;
        RECT 67.065 151.660 67.320 152.565 ;
        RECT 66.090 151.085 66.445 151.455 ;
        RECT 66.725 151.425 66.895 151.635 ;
        RECT 66.725 151.095 66.980 151.425 ;
        RECT 64.340 150.735 65.055 150.905 ;
        RECT 64.340 150.355 64.510 150.735 ;
        RECT 64.725 150.185 65.055 150.565 ;
        RECT 65.225 150.355 65.480 150.930 ;
        RECT 65.655 150.185 65.915 151.025 ;
        RECT 66.725 150.905 66.895 151.095 ;
        RECT 67.150 150.930 67.320 151.660 ;
        RECT 67.495 151.585 67.755 152.735 ;
        RECT 68.850 151.595 69.190 152.565 ;
        RECT 69.360 151.595 69.530 152.735 ;
        RECT 69.800 151.935 70.050 152.735 ;
        RECT 70.695 151.765 71.025 152.565 ;
        RECT 71.325 151.935 71.655 152.735 ;
        RECT 71.825 151.765 72.155 152.565 ;
        RECT 69.720 151.595 72.155 151.765 ;
        RECT 72.530 151.595 72.870 152.565 ;
        RECT 73.040 151.595 73.210 152.735 ;
        RECT 73.480 151.935 73.730 152.735 ;
        RECT 74.375 151.765 74.705 152.565 ;
        RECT 75.005 151.935 75.335 152.735 ;
        RECT 75.505 151.765 75.835 152.565 ;
        RECT 73.400 151.595 75.835 151.765 ;
        RECT 76.585 151.755 76.840 152.425 ;
        RECT 77.020 151.935 77.305 152.735 ;
        RECT 77.485 152.015 77.815 152.525 ;
        RECT 66.180 150.735 66.895 150.905 ;
        RECT 66.180 150.355 66.350 150.735 ;
        RECT 66.565 150.185 66.895 150.565 ;
        RECT 67.065 150.355 67.320 150.930 ;
        RECT 67.495 150.185 67.755 151.025 ;
        RECT 68.850 150.985 69.025 151.595 ;
        RECT 69.720 151.345 69.890 151.595 ;
        RECT 69.195 151.175 69.890 151.345 ;
        RECT 70.065 151.175 70.485 151.375 ;
        RECT 70.655 151.175 70.985 151.375 ;
        RECT 71.155 151.175 71.485 151.375 ;
        RECT 68.850 150.355 69.190 150.985 ;
        RECT 69.360 150.185 69.610 150.985 ;
        RECT 69.800 150.835 71.025 151.005 ;
        RECT 69.800 150.355 70.130 150.835 ;
        RECT 70.300 150.185 70.525 150.645 ;
        RECT 70.695 150.355 71.025 150.835 ;
        RECT 71.655 150.965 71.825 151.595 ;
        RECT 72.010 151.175 72.360 151.425 ;
        RECT 72.530 150.985 72.705 151.595 ;
        RECT 73.400 151.345 73.570 151.595 ;
        RECT 72.875 151.175 73.570 151.345 ;
        RECT 73.745 151.175 74.165 151.375 ;
        RECT 74.335 151.175 74.665 151.375 ;
        RECT 74.835 151.175 75.165 151.375 ;
        RECT 71.655 150.355 72.155 150.965 ;
        RECT 72.530 150.355 72.870 150.985 ;
        RECT 73.040 150.185 73.290 150.985 ;
        RECT 73.480 150.835 74.705 151.005 ;
        RECT 73.480 150.355 73.810 150.835 ;
        RECT 73.980 150.185 74.205 150.645 ;
        RECT 74.375 150.355 74.705 150.835 ;
        RECT 75.335 150.965 75.505 151.595 ;
        RECT 75.690 151.175 76.040 151.425 ;
        RECT 75.335 150.355 75.835 150.965 ;
        RECT 76.585 150.895 76.765 151.755 ;
        RECT 77.485 151.425 77.735 152.015 ;
        RECT 78.085 151.865 78.255 152.475 ;
        RECT 78.425 152.045 78.755 152.735 ;
        RECT 78.985 152.185 79.225 152.475 ;
        RECT 79.425 152.355 79.845 152.735 ;
        RECT 80.025 152.265 80.655 152.515 ;
        RECT 81.125 152.355 81.455 152.735 ;
        RECT 80.025 152.185 80.195 152.265 ;
        RECT 81.625 152.185 81.795 152.475 ;
        RECT 81.975 152.355 82.355 152.735 ;
        RECT 82.595 152.350 83.425 152.520 ;
        RECT 78.985 152.015 80.195 152.185 ;
        RECT 76.935 151.095 77.735 151.425 ;
        RECT 76.585 150.695 76.840 150.895 ;
        RECT 76.500 150.525 76.840 150.695 ;
        RECT 76.585 150.365 76.840 150.525 ;
        RECT 77.020 150.185 77.305 150.645 ;
        RECT 77.485 150.445 77.735 151.095 ;
        RECT 77.935 151.845 78.255 151.865 ;
        RECT 77.935 151.675 79.855 151.845 ;
        RECT 77.935 150.780 78.125 151.675 ;
        RECT 80.025 151.505 80.195 152.015 ;
        RECT 80.365 151.755 80.885 152.065 ;
        RECT 78.295 151.335 80.195 151.505 ;
        RECT 78.295 151.275 78.625 151.335 ;
        RECT 78.775 151.105 79.105 151.165 ;
        RECT 78.445 150.835 79.105 151.105 ;
        RECT 77.935 150.450 78.255 150.780 ;
        RECT 78.435 150.185 79.095 150.665 ;
        RECT 79.295 150.575 79.465 151.335 ;
        RECT 80.365 151.165 80.545 151.575 ;
        RECT 79.635 150.995 79.965 151.115 ;
        RECT 80.715 150.995 80.885 151.755 ;
        RECT 79.635 150.825 80.885 150.995 ;
        RECT 81.055 151.935 82.425 152.185 ;
        RECT 81.055 151.165 81.245 151.935 ;
        RECT 82.175 151.675 82.425 151.935 ;
        RECT 81.415 151.505 81.665 151.665 ;
        RECT 82.595 151.505 82.765 152.350 ;
        RECT 83.660 152.065 83.830 152.565 ;
        RECT 84.000 152.235 84.330 152.735 ;
        RECT 82.935 151.675 83.435 152.055 ;
        RECT 83.660 151.895 84.355 152.065 ;
        RECT 81.415 151.335 82.765 151.505 ;
        RECT 82.345 151.295 82.765 151.335 ;
        RECT 81.055 150.825 81.475 151.165 ;
        RECT 81.765 150.835 82.175 151.165 ;
        RECT 79.295 150.405 80.145 150.575 ;
        RECT 80.705 150.185 81.025 150.645 ;
        RECT 81.225 150.395 81.475 150.825 ;
        RECT 81.765 150.185 82.175 150.625 ;
        RECT 82.345 150.565 82.515 151.295 ;
        RECT 82.685 150.745 83.035 151.115 ;
        RECT 83.215 150.805 83.435 151.675 ;
        RECT 83.605 151.105 84.015 151.725 ;
        RECT 84.185 150.925 84.355 151.895 ;
        RECT 83.660 150.735 84.355 150.925 ;
        RECT 82.345 150.365 83.360 150.565 ;
        RECT 83.660 150.405 83.830 150.735 ;
        RECT 84.000 150.185 84.330 150.565 ;
        RECT 84.545 150.445 84.770 152.565 ;
        RECT 84.940 152.235 85.270 152.735 ;
        RECT 85.440 152.065 85.610 152.565 ;
        RECT 84.945 151.895 85.610 152.065 ;
        RECT 84.945 150.905 85.175 151.895 ;
        RECT 85.345 151.075 85.695 151.725 ;
        RECT 86.330 151.570 86.620 152.735 ;
        RECT 87.750 151.595 87.980 152.735 ;
        RECT 88.150 151.585 88.480 152.565 ;
        RECT 88.650 151.595 88.860 152.735 ;
        RECT 89.295 151.765 89.625 152.565 ;
        RECT 89.795 151.935 90.125 152.735 ;
        RECT 90.425 151.765 90.755 152.565 ;
        RECT 91.400 151.935 91.650 152.735 ;
        RECT 89.295 151.595 91.730 151.765 ;
        RECT 91.920 151.595 92.090 152.735 ;
        RECT 92.260 151.595 92.600 152.565 ;
        RECT 92.975 151.765 93.305 152.565 ;
        RECT 93.475 151.935 93.805 152.735 ;
        RECT 94.105 151.765 94.435 152.565 ;
        RECT 95.080 151.935 95.330 152.735 ;
        RECT 92.975 151.595 95.410 151.765 ;
        RECT 95.600 151.595 95.770 152.735 ;
        RECT 95.940 151.595 96.280 152.565 ;
        RECT 97.575 151.765 97.905 152.565 ;
        RECT 98.075 151.935 98.405 152.735 ;
        RECT 98.705 151.765 99.035 152.565 ;
        RECT 99.680 151.935 99.930 152.735 ;
        RECT 97.575 151.595 100.010 151.765 ;
        RECT 100.200 151.595 100.370 152.735 ;
        RECT 100.540 151.595 100.880 152.565 ;
        RECT 87.730 151.175 88.060 151.425 ;
        RECT 84.945 150.735 85.610 150.905 ;
        RECT 84.940 150.185 85.270 150.565 ;
        RECT 85.440 150.445 85.610 150.735 ;
        RECT 86.330 150.185 86.620 150.910 ;
        RECT 87.750 150.185 87.980 151.005 ;
        RECT 88.230 150.985 88.480 151.585 ;
        RECT 89.090 151.175 89.440 151.425 ;
        RECT 88.150 150.355 88.480 150.985 ;
        RECT 88.650 150.185 88.860 151.005 ;
        RECT 89.625 150.965 89.795 151.595 ;
        RECT 89.965 151.175 90.295 151.375 ;
        RECT 90.465 151.175 90.795 151.375 ;
        RECT 90.965 151.175 91.385 151.375 ;
        RECT 91.560 151.345 91.730 151.595 ;
        RECT 91.560 151.175 92.255 151.345 ;
        RECT 89.295 150.355 89.795 150.965 ;
        RECT 90.425 150.835 91.650 151.005 ;
        RECT 92.425 150.985 92.600 151.595 ;
        RECT 92.770 151.175 93.120 151.425 ;
        RECT 90.425 150.355 90.755 150.835 ;
        RECT 90.925 150.185 91.150 150.645 ;
        RECT 91.320 150.355 91.650 150.835 ;
        RECT 91.840 150.185 92.090 150.985 ;
        RECT 92.260 150.355 92.600 150.985 ;
        RECT 93.305 150.965 93.475 151.595 ;
        RECT 93.645 151.175 93.975 151.375 ;
        RECT 94.145 151.175 94.475 151.375 ;
        RECT 94.645 151.175 95.065 151.375 ;
        RECT 95.240 151.345 95.410 151.595 ;
        RECT 95.240 151.175 95.935 151.345 ;
        RECT 92.975 150.355 93.475 150.965 ;
        RECT 94.105 150.835 95.330 151.005 ;
        RECT 96.105 150.985 96.280 151.595 ;
        RECT 97.370 151.175 97.720 151.425 ;
        RECT 94.105 150.355 94.435 150.835 ;
        RECT 94.605 150.185 94.830 150.645 ;
        RECT 95.000 150.355 95.330 150.835 ;
        RECT 95.520 150.185 95.770 150.985 ;
        RECT 95.940 150.355 96.280 150.985 ;
        RECT 97.905 150.965 98.075 151.595 ;
        RECT 98.245 151.175 98.575 151.375 ;
        RECT 98.745 151.175 99.075 151.375 ;
        RECT 99.245 151.175 99.665 151.375 ;
        RECT 99.840 151.345 100.010 151.595 ;
        RECT 99.840 151.175 100.535 151.345 ;
        RECT 97.575 150.355 98.075 150.965 ;
        RECT 98.705 150.835 99.930 151.005 ;
        RECT 100.705 150.985 100.880 151.595 ;
        RECT 98.705 150.355 99.035 150.835 ;
        RECT 99.205 150.185 99.430 150.645 ;
        RECT 99.600 150.355 99.930 150.835 ;
        RECT 100.120 150.185 100.370 150.985 ;
        RECT 100.540 150.355 100.880 150.985 ;
        RECT 101.515 151.545 101.770 152.425 ;
        RECT 101.940 151.595 102.245 152.735 ;
        RECT 102.585 152.355 102.915 152.735 ;
        RECT 103.095 152.185 103.265 152.475 ;
        RECT 103.435 152.275 103.685 152.735 ;
        RECT 102.465 152.015 103.265 152.185 ;
        RECT 103.855 152.225 104.725 152.565 ;
        RECT 101.515 150.895 101.725 151.545 ;
        RECT 102.465 151.425 102.635 152.015 ;
        RECT 103.855 151.845 104.025 152.225 ;
        RECT 104.960 152.105 105.130 152.565 ;
        RECT 105.300 152.275 105.670 152.735 ;
        RECT 105.965 152.135 106.135 152.475 ;
        RECT 106.305 152.305 106.635 152.735 ;
        RECT 106.870 152.135 107.040 152.475 ;
        RECT 102.805 151.675 104.025 151.845 ;
        RECT 104.195 151.765 104.655 152.055 ;
        RECT 104.960 151.935 105.520 152.105 ;
        RECT 105.965 151.965 107.040 152.135 ;
        RECT 107.210 152.235 107.890 152.565 ;
        RECT 108.105 152.235 108.355 152.565 ;
        RECT 108.525 152.275 108.775 152.735 ;
        RECT 105.350 151.795 105.520 151.935 ;
        RECT 104.195 151.755 105.160 151.765 ;
        RECT 103.855 151.585 104.025 151.675 ;
        RECT 104.485 151.595 105.160 151.755 ;
        RECT 101.895 151.395 102.635 151.425 ;
        RECT 101.895 151.095 102.810 151.395 ;
        RECT 102.485 150.920 102.810 151.095 ;
        RECT 101.515 150.365 101.770 150.895 ;
        RECT 101.940 150.185 102.245 150.645 ;
        RECT 102.490 150.565 102.810 150.920 ;
        RECT 102.980 151.135 103.520 151.505 ;
        RECT 103.855 151.415 104.260 151.585 ;
        RECT 102.980 150.735 103.220 151.135 ;
        RECT 103.700 150.965 103.920 151.245 ;
        RECT 103.390 150.795 103.920 150.965 ;
        RECT 103.390 150.565 103.560 150.795 ;
        RECT 104.090 150.635 104.260 151.415 ;
        RECT 104.430 150.805 104.780 151.425 ;
        RECT 104.950 150.805 105.160 151.595 ;
        RECT 105.350 151.625 106.850 151.795 ;
        RECT 105.350 150.935 105.520 151.625 ;
        RECT 107.210 151.455 107.380 152.235 ;
        RECT 108.185 152.105 108.355 152.235 ;
        RECT 105.690 151.285 107.380 151.455 ;
        RECT 107.550 151.675 108.015 152.065 ;
        RECT 108.185 151.935 108.580 152.105 ;
        RECT 105.690 151.105 105.860 151.285 ;
        RECT 102.490 150.395 103.560 150.565 ;
        RECT 103.730 150.185 103.920 150.625 ;
        RECT 104.090 150.355 105.040 150.635 ;
        RECT 105.350 150.545 105.610 150.935 ;
        RECT 106.030 150.865 106.820 151.115 ;
        RECT 105.260 150.375 105.610 150.545 ;
        RECT 105.820 150.185 106.150 150.645 ;
        RECT 107.025 150.575 107.195 151.285 ;
        RECT 107.550 151.085 107.720 151.675 ;
        RECT 107.365 150.865 107.720 151.085 ;
        RECT 107.890 150.865 108.240 151.485 ;
        RECT 108.410 150.575 108.580 151.935 ;
        RECT 108.945 151.765 109.270 152.550 ;
        RECT 108.750 150.715 109.210 151.765 ;
        RECT 107.025 150.405 107.880 150.575 ;
        RECT 108.085 150.405 108.580 150.575 ;
        RECT 108.750 150.185 109.080 150.545 ;
        RECT 109.440 150.445 109.610 152.565 ;
        RECT 109.780 152.235 110.110 152.735 ;
        RECT 110.280 152.065 110.535 152.565 ;
        RECT 109.785 151.895 110.535 152.065 ;
        RECT 109.785 150.905 110.015 151.895 ;
        RECT 110.185 151.075 110.535 151.725 ;
        RECT 111.170 151.645 112.380 152.735 ;
        RECT 111.170 151.105 111.690 151.645 ;
        RECT 111.860 150.935 112.380 151.475 ;
        RECT 109.785 150.735 110.535 150.905 ;
        RECT 109.780 150.185 110.110 150.565 ;
        RECT 110.280 150.445 110.535 150.735 ;
        RECT 111.170 150.185 112.380 150.935 ;
        RECT 18.165 150.015 112.465 150.185 ;
        RECT 18.250 149.265 19.460 150.015 ;
        RECT 18.250 148.725 18.770 149.265 ;
        RECT 20.090 149.245 21.760 150.015 ;
        RECT 21.930 149.290 22.220 150.015 ;
        RECT 18.940 148.555 19.460 149.095 ;
        RECT 18.250 147.465 19.460 148.555 ;
        RECT 20.090 148.555 20.840 149.075 ;
        RECT 21.010 148.725 21.760 149.245 ;
        RECT 22.430 149.195 22.660 150.015 ;
        RECT 22.830 149.215 23.160 149.845 ;
        RECT 22.410 148.775 22.740 149.025 ;
        RECT 20.090 147.465 21.760 148.555 ;
        RECT 21.930 147.465 22.220 148.630 ;
        RECT 22.910 148.615 23.160 149.215 ;
        RECT 23.330 149.195 23.540 150.015 ;
        RECT 23.770 149.340 24.030 149.845 ;
        RECT 24.210 149.635 24.540 150.015 ;
        RECT 24.720 149.465 24.890 149.845 ;
        RECT 22.430 147.465 22.660 148.605 ;
        RECT 22.830 147.635 23.160 148.615 ;
        RECT 23.330 147.465 23.540 148.605 ;
        RECT 23.770 148.540 23.940 149.340 ;
        RECT 24.225 149.295 24.890 149.465 ;
        RECT 24.225 149.040 24.395 149.295 ;
        RECT 25.155 149.275 25.410 149.845 ;
        RECT 25.580 149.615 25.910 150.015 ;
        RECT 26.335 149.480 26.865 149.845 ;
        RECT 26.335 149.445 26.510 149.480 ;
        RECT 25.580 149.275 26.510 149.445 ;
        RECT 24.110 148.710 24.395 149.040 ;
        RECT 24.630 148.745 24.960 149.115 ;
        RECT 24.225 148.565 24.395 148.710 ;
        RECT 25.155 148.605 25.325 149.275 ;
        RECT 25.580 149.105 25.750 149.275 ;
        RECT 25.495 148.775 25.750 149.105 ;
        RECT 25.975 148.775 26.170 149.105 ;
        RECT 23.770 147.635 24.040 148.540 ;
        RECT 24.225 148.395 24.890 148.565 ;
        RECT 24.210 147.465 24.540 148.225 ;
        RECT 24.720 147.635 24.890 148.395 ;
        RECT 25.155 147.635 25.490 148.605 ;
        RECT 25.660 147.465 25.830 148.605 ;
        RECT 26.000 147.805 26.170 148.775 ;
        RECT 26.340 148.145 26.510 149.275 ;
        RECT 26.680 148.485 26.850 149.285 ;
        RECT 27.055 148.995 27.330 149.845 ;
        RECT 27.050 148.825 27.330 148.995 ;
        RECT 27.055 148.685 27.330 148.825 ;
        RECT 27.500 148.485 27.690 149.845 ;
        RECT 27.870 149.480 28.380 150.015 ;
        RECT 28.600 149.205 28.845 149.810 ;
        RECT 27.890 149.035 29.120 149.205 ;
        RECT 29.330 149.195 29.560 150.015 ;
        RECT 29.730 149.215 30.060 149.845 ;
        RECT 26.680 148.315 27.690 148.485 ;
        RECT 27.860 148.470 28.610 148.660 ;
        RECT 26.340 147.975 27.465 148.145 ;
        RECT 27.860 147.805 28.030 148.470 ;
        RECT 28.780 148.225 29.120 149.035 ;
        RECT 29.310 148.775 29.640 149.025 ;
        RECT 29.810 148.615 30.060 149.215 ;
        RECT 30.230 149.195 30.440 150.015 ;
        RECT 30.760 149.465 30.930 149.755 ;
        RECT 31.100 149.635 31.430 150.015 ;
        RECT 30.760 149.295 31.425 149.465 ;
        RECT 26.000 147.635 28.030 147.805 ;
        RECT 28.200 147.465 28.370 148.225 ;
        RECT 28.605 147.815 29.120 148.225 ;
        RECT 29.330 147.465 29.560 148.605 ;
        RECT 29.730 147.635 30.060 148.615 ;
        RECT 30.230 147.465 30.440 148.605 ;
        RECT 30.675 148.475 31.025 149.125 ;
        RECT 31.195 148.305 31.425 149.295 ;
        RECT 30.760 148.135 31.425 148.305 ;
        RECT 30.760 147.635 30.930 148.135 ;
        RECT 31.100 147.465 31.430 147.965 ;
        RECT 31.600 147.635 31.825 149.755 ;
        RECT 32.040 149.635 32.370 150.015 ;
        RECT 32.540 149.465 32.710 149.795 ;
        RECT 33.010 149.635 34.025 149.835 ;
        RECT 32.015 149.275 32.710 149.465 ;
        RECT 32.015 148.305 32.185 149.275 ;
        RECT 32.355 148.475 32.765 149.095 ;
        RECT 32.935 148.525 33.155 149.395 ;
        RECT 33.335 149.085 33.685 149.455 ;
        RECT 33.855 148.905 34.025 149.635 ;
        RECT 34.195 149.575 34.605 150.015 ;
        RECT 34.895 149.375 35.145 149.805 ;
        RECT 35.345 149.555 35.665 150.015 ;
        RECT 36.225 149.625 37.075 149.795 ;
        RECT 34.195 149.035 34.605 149.365 ;
        RECT 34.895 149.035 35.315 149.375 ;
        RECT 33.605 148.865 34.025 148.905 ;
        RECT 33.605 148.695 34.955 148.865 ;
        RECT 32.015 148.135 32.710 148.305 ;
        RECT 32.935 148.145 33.435 148.525 ;
        RECT 32.040 147.465 32.370 147.965 ;
        RECT 32.540 147.635 32.710 148.135 ;
        RECT 33.605 147.850 33.775 148.695 ;
        RECT 34.705 148.535 34.955 148.695 ;
        RECT 33.945 148.265 34.195 148.525 ;
        RECT 35.125 148.265 35.315 149.035 ;
        RECT 33.945 148.015 35.315 148.265 ;
        RECT 35.485 149.205 36.735 149.375 ;
        RECT 35.485 148.445 35.655 149.205 ;
        RECT 36.405 149.085 36.735 149.205 ;
        RECT 35.825 148.625 36.005 149.035 ;
        RECT 36.905 148.865 37.075 149.625 ;
        RECT 37.275 149.535 37.935 150.015 ;
        RECT 38.115 149.420 38.435 149.750 ;
        RECT 37.265 149.095 37.925 149.365 ;
        RECT 37.265 149.035 37.595 149.095 ;
        RECT 37.745 148.865 38.075 148.925 ;
        RECT 36.175 148.695 38.075 148.865 ;
        RECT 35.485 148.135 36.005 148.445 ;
        RECT 36.175 148.185 36.345 148.695 ;
        RECT 38.245 148.525 38.435 149.420 ;
        RECT 36.515 148.355 38.435 148.525 ;
        RECT 38.115 148.335 38.435 148.355 ;
        RECT 38.635 149.105 38.885 149.755 ;
        RECT 39.065 149.555 39.350 150.015 ;
        RECT 39.530 149.305 39.785 149.835 ;
        RECT 40.430 149.550 40.680 150.015 ;
        RECT 40.850 149.375 41.020 149.845 ;
        RECT 41.270 149.555 41.440 150.015 ;
        RECT 41.690 149.375 41.860 149.845 ;
        RECT 42.110 149.555 42.280 150.015 ;
        RECT 42.530 149.375 42.700 149.845 ;
        RECT 43.070 149.555 43.335 150.015 ;
        RECT 38.635 148.775 39.435 149.105 ;
        RECT 36.175 148.015 37.385 148.185 ;
        RECT 32.945 147.680 33.775 147.850 ;
        RECT 34.015 147.465 34.395 147.845 ;
        RECT 34.575 147.725 34.745 148.015 ;
        RECT 36.175 147.935 36.345 148.015 ;
        RECT 34.915 147.465 35.245 147.845 ;
        RECT 35.715 147.685 36.345 147.935 ;
        RECT 36.525 147.465 36.945 147.845 ;
        RECT 37.145 147.725 37.385 148.015 ;
        RECT 37.615 147.465 37.945 148.155 ;
        RECT 38.115 147.725 38.285 148.335 ;
        RECT 38.635 148.185 38.885 148.775 ;
        RECT 39.605 148.445 39.785 149.305 ;
        RECT 39.530 148.315 39.785 148.445 ;
        RECT 40.330 149.195 42.700 149.375 ;
        RECT 44.010 149.215 44.350 149.845 ;
        RECT 44.520 149.215 44.770 150.015 ;
        RECT 44.960 149.365 45.290 149.845 ;
        RECT 45.460 149.555 45.685 150.015 ;
        RECT 45.855 149.365 46.185 149.845 ;
        RECT 40.330 148.605 40.680 149.195 ;
        RECT 40.850 148.775 43.360 149.025 ;
        RECT 44.010 148.605 44.185 149.215 ;
        RECT 44.960 149.195 46.185 149.365 ;
        RECT 46.815 149.235 47.315 149.845 ;
        RECT 47.690 149.290 47.980 150.015 ;
        RECT 44.355 148.855 45.050 149.025 ;
        RECT 44.880 148.605 45.050 148.855 ;
        RECT 45.225 148.825 45.645 149.025 ;
        RECT 45.815 148.825 46.145 149.025 ;
        RECT 46.315 148.825 46.645 149.025 ;
        RECT 46.815 148.605 46.985 149.235 ;
        RECT 48.610 149.215 48.950 149.845 ;
        RECT 49.120 149.215 49.370 150.015 ;
        RECT 49.560 149.365 49.890 149.845 ;
        RECT 50.060 149.555 50.285 150.015 ;
        RECT 50.455 149.365 50.785 149.845 ;
        RECT 47.170 148.775 47.520 149.025 ;
        RECT 40.330 148.435 42.780 148.605 ;
        RECT 40.330 148.415 41.100 148.435 ;
        RECT 38.555 147.675 38.885 148.185 ;
        RECT 39.065 147.465 39.350 148.265 ;
        RECT 39.530 148.145 39.870 148.315 ;
        RECT 39.530 147.775 39.785 148.145 ;
        RECT 40.430 147.465 40.600 147.925 ;
        RECT 40.770 147.635 41.100 148.415 ;
        RECT 41.270 147.465 41.440 148.265 ;
        RECT 41.610 147.635 41.940 148.435 ;
        RECT 42.110 147.465 42.280 148.265 ;
        RECT 42.450 147.635 42.780 148.435 ;
        RECT 43.040 147.465 43.335 148.605 ;
        RECT 44.010 147.635 44.350 148.605 ;
        RECT 44.520 147.465 44.690 148.605 ;
        RECT 44.880 148.435 47.315 148.605 ;
        RECT 44.960 147.465 45.210 148.265 ;
        RECT 45.855 147.635 46.185 148.435 ;
        RECT 46.485 147.465 46.815 148.265 ;
        RECT 46.985 147.635 47.315 148.435 ;
        RECT 47.690 147.465 47.980 148.630 ;
        RECT 48.610 148.605 48.785 149.215 ;
        RECT 49.560 149.195 50.785 149.365 ;
        RECT 51.415 149.235 51.915 149.845 ;
        RECT 48.955 148.855 49.650 149.025 ;
        RECT 49.480 148.605 49.650 148.855 ;
        RECT 49.825 148.825 50.245 149.025 ;
        RECT 50.415 148.825 50.745 149.025 ;
        RECT 50.915 148.825 51.245 149.025 ;
        RECT 51.415 148.605 51.585 149.235 ;
        RECT 52.565 149.205 52.810 149.810 ;
        RECT 53.030 149.480 53.540 150.015 ;
        RECT 52.290 149.035 53.520 149.205 ;
        RECT 51.770 148.775 52.120 149.025 ;
        RECT 48.610 147.635 48.950 148.605 ;
        RECT 49.120 147.465 49.290 148.605 ;
        RECT 49.480 148.435 51.915 148.605 ;
        RECT 49.560 147.465 49.810 148.265 ;
        RECT 50.455 147.635 50.785 148.435 ;
        RECT 51.085 147.465 51.415 148.265 ;
        RECT 51.585 147.635 51.915 148.435 ;
        RECT 52.290 148.225 52.630 149.035 ;
        RECT 52.800 148.470 53.550 148.660 ;
        RECT 52.290 147.815 52.805 148.225 ;
        RECT 53.040 147.465 53.210 148.225 ;
        RECT 53.380 147.805 53.550 148.470 ;
        RECT 53.720 148.485 53.910 149.845 ;
        RECT 54.080 149.335 54.355 149.845 ;
        RECT 54.545 149.480 55.075 149.845 ;
        RECT 55.500 149.615 55.830 150.015 ;
        RECT 54.900 149.445 55.075 149.480 ;
        RECT 54.080 149.165 54.360 149.335 ;
        RECT 54.080 148.685 54.355 149.165 ;
        RECT 54.560 148.485 54.730 149.285 ;
        RECT 53.720 148.315 54.730 148.485 ;
        RECT 54.900 149.275 55.830 149.445 ;
        RECT 56.000 149.275 56.255 149.845 ;
        RECT 54.900 148.145 55.070 149.275 ;
        RECT 55.660 149.105 55.830 149.275 ;
        RECT 53.945 147.975 55.070 148.145 ;
        RECT 55.240 148.775 55.435 149.105 ;
        RECT 55.660 148.775 55.915 149.105 ;
        RECT 55.240 147.805 55.410 148.775 ;
        RECT 56.085 148.605 56.255 149.275 ;
        RECT 56.705 149.205 56.950 149.810 ;
        RECT 57.170 149.480 57.680 150.015 ;
        RECT 53.380 147.635 55.410 147.805 ;
        RECT 55.580 147.465 55.750 148.605 ;
        RECT 55.920 147.635 56.255 148.605 ;
        RECT 56.430 149.035 57.660 149.205 ;
        RECT 56.430 148.225 56.770 149.035 ;
        RECT 56.940 148.470 57.690 148.660 ;
        RECT 56.430 147.815 56.945 148.225 ;
        RECT 57.180 147.465 57.350 148.225 ;
        RECT 57.520 147.805 57.690 148.470 ;
        RECT 57.860 148.485 58.050 149.845 ;
        RECT 58.220 148.995 58.495 149.845 ;
        RECT 58.685 149.480 59.215 149.845 ;
        RECT 59.640 149.615 59.970 150.015 ;
        RECT 59.040 149.445 59.215 149.480 ;
        RECT 58.220 148.825 58.500 148.995 ;
        RECT 58.220 148.685 58.495 148.825 ;
        RECT 58.700 148.485 58.870 149.285 ;
        RECT 57.860 148.315 58.870 148.485 ;
        RECT 59.040 149.275 59.970 149.445 ;
        RECT 60.140 149.275 60.395 149.845 ;
        RECT 59.040 148.145 59.210 149.275 ;
        RECT 59.800 149.105 59.970 149.275 ;
        RECT 58.085 147.975 59.210 148.145 ;
        RECT 59.380 148.775 59.575 149.105 ;
        RECT 59.800 148.775 60.055 149.105 ;
        RECT 59.380 147.805 59.550 148.775 ;
        RECT 60.225 148.605 60.395 149.275 ;
        RECT 57.520 147.635 59.550 147.805 ;
        RECT 59.720 147.465 59.890 148.605 ;
        RECT 60.060 147.635 60.395 148.605 ;
        RECT 60.570 149.340 60.830 149.845 ;
        RECT 61.010 149.635 61.340 150.015 ;
        RECT 61.520 149.465 61.690 149.845 ;
        RECT 60.570 148.540 60.740 149.340 ;
        RECT 61.025 149.295 61.690 149.465 ;
        RECT 61.025 149.040 61.195 149.295 ;
        RECT 61.990 149.195 62.220 150.015 ;
        RECT 62.390 149.215 62.720 149.845 ;
        RECT 60.910 148.710 61.195 149.040 ;
        RECT 61.430 148.745 61.760 149.115 ;
        RECT 61.970 148.775 62.300 149.025 ;
        RECT 61.025 148.565 61.195 148.710 ;
        RECT 62.470 148.615 62.720 149.215 ;
        RECT 62.890 149.195 63.100 150.015 ;
        RECT 63.420 149.465 63.590 149.845 ;
        RECT 63.805 149.635 64.135 150.015 ;
        RECT 63.420 149.295 64.135 149.465 ;
        RECT 63.330 148.745 63.685 149.115 ;
        RECT 63.965 149.105 64.135 149.295 ;
        RECT 64.305 149.270 64.560 149.845 ;
        RECT 63.965 148.775 64.220 149.105 ;
        RECT 60.570 147.635 60.840 148.540 ;
        RECT 61.025 148.395 61.690 148.565 ;
        RECT 61.010 147.465 61.340 148.225 ;
        RECT 61.520 147.635 61.690 148.395 ;
        RECT 61.990 147.465 62.220 148.605 ;
        RECT 62.390 147.635 62.720 148.615 ;
        RECT 62.890 147.465 63.100 148.605 ;
        RECT 63.965 148.565 64.135 148.775 ;
        RECT 63.420 148.395 64.135 148.565 ;
        RECT 64.390 148.540 64.560 149.270 ;
        RECT 64.735 149.175 64.995 150.015 ;
        RECT 65.175 149.250 65.630 150.015 ;
        RECT 65.905 149.635 67.205 149.845 ;
        RECT 67.460 149.655 67.790 150.015 ;
        RECT 67.035 149.485 67.205 149.635 ;
        RECT 67.960 149.515 68.220 149.845 ;
        RECT 66.105 149.025 66.325 149.425 ;
        RECT 65.170 148.825 65.660 149.025 ;
        RECT 65.850 148.815 66.325 149.025 ;
        RECT 66.570 149.025 66.780 149.425 ;
        RECT 67.035 149.360 67.790 149.485 ;
        RECT 67.035 149.315 67.880 149.360 ;
        RECT 67.610 149.195 67.880 149.315 ;
        RECT 66.570 148.815 66.900 149.025 ;
        RECT 67.070 148.755 67.480 149.060 ;
        RECT 63.420 147.635 63.590 148.395 ;
        RECT 63.805 147.465 64.135 148.225 ;
        RECT 64.305 147.635 64.560 148.540 ;
        RECT 64.735 147.465 64.995 148.615 ;
        RECT 65.175 148.585 66.350 148.645 ;
        RECT 67.710 148.620 67.880 149.195 ;
        RECT 67.680 148.585 67.880 148.620 ;
        RECT 65.175 148.475 67.880 148.585 ;
        RECT 65.175 147.855 65.430 148.475 ;
        RECT 66.020 148.415 67.820 148.475 ;
        RECT 66.020 148.385 66.350 148.415 ;
        RECT 68.050 148.315 68.220 149.515 ;
        RECT 68.395 149.175 68.655 150.015 ;
        RECT 68.830 149.270 69.085 149.845 ;
        RECT 69.255 149.635 69.585 150.015 ;
        RECT 69.800 149.465 69.970 149.845 ;
        RECT 69.255 149.295 69.970 149.465 ;
        RECT 70.320 149.465 70.490 149.845 ;
        RECT 70.705 149.635 71.035 150.015 ;
        RECT 70.320 149.295 71.035 149.465 ;
        RECT 65.680 148.215 65.865 148.305 ;
        RECT 66.455 148.215 67.290 148.225 ;
        RECT 65.680 148.015 67.290 148.215 ;
        RECT 65.680 147.975 65.910 148.015 ;
        RECT 65.175 147.635 65.510 147.855 ;
        RECT 66.515 147.465 66.870 147.845 ;
        RECT 67.040 147.635 67.290 148.015 ;
        RECT 67.540 147.465 67.790 148.245 ;
        RECT 67.960 147.635 68.220 148.315 ;
        RECT 68.395 147.465 68.655 148.615 ;
        RECT 68.830 148.540 69.000 149.270 ;
        RECT 69.255 149.105 69.425 149.295 ;
        RECT 69.170 148.775 69.425 149.105 ;
        RECT 69.255 148.565 69.425 148.775 ;
        RECT 69.705 148.745 70.060 149.115 ;
        RECT 70.230 148.745 70.585 149.115 ;
        RECT 70.865 149.105 71.035 149.295 ;
        RECT 71.205 149.270 71.460 149.845 ;
        RECT 70.865 148.775 71.120 149.105 ;
        RECT 70.865 148.565 71.035 148.775 ;
        RECT 68.830 147.635 69.085 148.540 ;
        RECT 69.255 148.395 69.970 148.565 ;
        RECT 69.255 147.465 69.585 148.225 ;
        RECT 69.800 147.635 69.970 148.395 ;
        RECT 70.320 148.395 71.035 148.565 ;
        RECT 71.290 148.540 71.460 149.270 ;
        RECT 71.635 149.175 71.895 150.015 ;
        RECT 72.070 149.340 72.330 149.845 ;
        RECT 72.510 149.635 72.840 150.015 ;
        RECT 73.020 149.465 73.190 149.845 ;
        RECT 70.320 147.635 70.490 148.395 ;
        RECT 70.705 147.465 71.035 148.225 ;
        RECT 71.205 147.635 71.460 148.540 ;
        RECT 71.635 147.465 71.895 148.615 ;
        RECT 72.070 148.540 72.240 149.340 ;
        RECT 72.525 149.295 73.190 149.465 ;
        RECT 72.525 149.040 72.695 149.295 ;
        RECT 73.450 149.290 73.740 150.015 ;
        RECT 74.370 149.245 77.880 150.015 ;
        RECT 72.410 148.710 72.695 149.040 ;
        RECT 72.930 148.745 73.260 149.115 ;
        RECT 72.525 148.565 72.695 148.710 ;
        RECT 72.070 147.635 72.340 148.540 ;
        RECT 72.525 148.395 73.190 148.565 ;
        RECT 72.510 147.465 72.840 148.225 ;
        RECT 73.020 147.635 73.190 148.395 ;
        RECT 73.450 147.465 73.740 148.630 ;
        RECT 74.370 148.555 76.060 149.075 ;
        RECT 76.230 148.725 77.880 149.245 ;
        RECT 78.110 149.195 78.320 150.015 ;
        RECT 78.490 149.215 78.820 149.845 ;
        RECT 78.490 148.615 78.740 149.215 ;
        RECT 78.990 149.195 79.220 150.015 ;
        RECT 79.470 149.195 79.700 150.015 ;
        RECT 79.870 149.215 80.200 149.845 ;
        RECT 78.910 148.775 79.240 149.025 ;
        RECT 79.450 148.775 79.780 149.025 ;
        RECT 79.950 148.615 80.200 149.215 ;
        RECT 80.370 149.195 80.580 150.015 ;
        RECT 81.085 149.205 81.330 149.810 ;
        RECT 81.550 149.480 82.060 150.015 ;
        RECT 74.370 147.465 77.880 148.555 ;
        RECT 78.110 147.465 78.320 148.605 ;
        RECT 78.490 147.635 78.820 148.615 ;
        RECT 78.990 147.465 79.220 148.605 ;
        RECT 79.470 147.465 79.700 148.605 ;
        RECT 79.870 147.635 80.200 148.615 ;
        RECT 80.810 149.035 82.040 149.205 ;
        RECT 80.370 147.465 80.580 148.605 ;
        RECT 80.810 148.225 81.150 149.035 ;
        RECT 81.320 148.470 82.070 148.660 ;
        RECT 80.810 147.815 81.325 148.225 ;
        RECT 81.560 147.465 81.730 148.225 ;
        RECT 81.900 147.805 82.070 148.470 ;
        RECT 82.240 148.485 82.430 149.845 ;
        RECT 82.600 149.335 82.875 149.845 ;
        RECT 83.065 149.480 83.595 149.845 ;
        RECT 84.020 149.615 84.350 150.015 ;
        RECT 83.420 149.445 83.595 149.480 ;
        RECT 82.600 149.165 82.880 149.335 ;
        RECT 82.600 148.685 82.875 149.165 ;
        RECT 83.080 148.485 83.250 149.285 ;
        RECT 82.240 148.315 83.250 148.485 ;
        RECT 83.420 149.275 84.350 149.445 ;
        RECT 84.520 149.275 84.775 149.845 ;
        RECT 83.420 148.145 83.590 149.275 ;
        RECT 84.180 149.105 84.350 149.275 ;
        RECT 82.465 147.975 83.590 148.145 ;
        RECT 83.760 148.775 83.955 149.105 ;
        RECT 84.180 148.775 84.435 149.105 ;
        RECT 83.760 147.805 83.930 148.775 ;
        RECT 84.605 148.605 84.775 149.275 ;
        RECT 81.900 147.635 83.930 147.805 ;
        RECT 84.100 147.465 84.270 148.605 ;
        RECT 84.440 147.635 84.775 148.605 ;
        RECT 84.950 149.340 85.210 149.845 ;
        RECT 85.390 149.635 85.720 150.015 ;
        RECT 85.900 149.465 86.070 149.845 ;
        RECT 84.950 148.540 85.120 149.340 ;
        RECT 85.405 149.295 86.070 149.465 ;
        RECT 85.405 149.040 85.575 149.295 ;
        RECT 86.330 149.245 88.920 150.015 ;
        RECT 85.290 148.710 85.575 149.040 ;
        RECT 85.810 148.745 86.140 149.115 ;
        RECT 85.405 148.565 85.575 148.710 ;
        RECT 84.950 147.635 85.220 148.540 ;
        RECT 85.405 148.395 86.070 148.565 ;
        RECT 85.390 147.465 85.720 148.225 ;
        RECT 85.900 147.635 86.070 148.395 ;
        RECT 86.330 148.555 87.540 149.075 ;
        RECT 87.710 148.725 88.920 149.245 ;
        RECT 89.090 149.215 89.430 149.845 ;
        RECT 89.600 149.215 89.850 150.015 ;
        RECT 90.040 149.365 90.370 149.845 ;
        RECT 90.540 149.555 90.765 150.015 ;
        RECT 90.935 149.365 91.265 149.845 ;
        RECT 89.090 148.605 89.265 149.215 ;
        RECT 90.040 149.195 91.265 149.365 ;
        RECT 91.895 149.235 92.395 149.845 ;
        RECT 92.975 149.235 93.475 149.845 ;
        RECT 89.435 148.855 90.130 149.025 ;
        RECT 89.960 148.605 90.130 148.855 ;
        RECT 90.305 148.825 90.725 149.025 ;
        RECT 90.895 148.825 91.225 149.025 ;
        RECT 91.395 148.825 91.725 149.025 ;
        RECT 91.895 148.605 92.065 149.235 ;
        RECT 92.250 148.775 92.600 149.025 ;
        RECT 92.770 148.775 93.120 149.025 ;
        RECT 93.305 148.605 93.475 149.235 ;
        RECT 94.105 149.365 94.435 149.845 ;
        RECT 94.605 149.555 94.830 150.015 ;
        RECT 95.000 149.365 95.330 149.845 ;
        RECT 94.105 149.195 95.330 149.365 ;
        RECT 95.520 149.215 95.770 150.015 ;
        RECT 95.940 149.215 96.280 149.845 ;
        RECT 96.460 149.515 96.790 150.015 ;
        RECT 96.990 149.445 97.160 149.795 ;
        RECT 97.360 149.615 97.690 150.015 ;
        RECT 97.860 149.445 98.030 149.795 ;
        RECT 98.200 149.615 98.580 150.015 ;
        RECT 93.645 148.825 93.975 149.025 ;
        RECT 94.145 148.825 94.475 149.025 ;
        RECT 94.645 148.825 95.065 149.025 ;
        RECT 95.240 148.855 95.935 149.025 ;
        RECT 95.240 148.605 95.410 148.855 ;
        RECT 96.105 148.605 96.280 149.215 ;
        RECT 96.455 148.775 96.805 149.345 ;
        RECT 96.990 149.275 98.600 149.445 ;
        RECT 98.770 149.340 99.040 149.685 ;
        RECT 98.430 149.105 98.600 149.275 ;
        RECT 96.975 148.655 97.685 149.105 ;
        RECT 97.855 148.775 98.260 149.105 ;
        RECT 98.430 148.775 98.700 149.105 ;
        RECT 86.330 147.465 88.920 148.555 ;
        RECT 89.090 147.635 89.430 148.605 ;
        RECT 89.600 147.465 89.770 148.605 ;
        RECT 89.960 148.435 92.395 148.605 ;
        RECT 90.040 147.465 90.290 148.265 ;
        RECT 90.935 147.635 91.265 148.435 ;
        RECT 91.565 147.465 91.895 148.265 ;
        RECT 92.065 147.635 92.395 148.435 ;
        RECT 92.975 148.435 95.410 148.605 ;
        RECT 92.975 147.635 93.305 148.435 ;
        RECT 93.475 147.465 93.805 148.265 ;
        RECT 94.105 147.635 94.435 148.435 ;
        RECT 95.080 147.465 95.330 148.265 ;
        RECT 95.600 147.465 95.770 148.605 ;
        RECT 95.940 147.635 96.280 148.605 ;
        RECT 96.455 148.315 96.775 148.605 ;
        RECT 96.970 148.485 97.685 148.655 ;
        RECT 98.430 148.605 98.600 148.775 ;
        RECT 98.870 148.605 99.040 149.340 ;
        RECT 99.210 149.290 99.500 150.015 ;
        RECT 100.170 149.195 100.400 150.015 ;
        RECT 100.570 149.215 100.900 149.845 ;
        RECT 100.150 148.775 100.480 149.025 ;
        RECT 97.875 148.435 98.600 148.605 ;
        RECT 97.875 148.315 98.045 148.435 ;
        RECT 96.455 148.145 98.045 148.315 ;
        RECT 96.455 147.685 98.110 147.975 ;
        RECT 98.280 147.465 98.560 148.265 ;
        RECT 98.770 147.635 99.040 148.605 ;
        RECT 99.210 147.465 99.500 148.630 ;
        RECT 100.650 148.615 100.900 149.215 ;
        RECT 101.070 149.195 101.280 150.015 ;
        RECT 101.885 149.305 102.140 149.835 ;
        RECT 102.320 149.555 102.605 150.015 ;
        RECT 100.170 147.465 100.400 148.605 ;
        RECT 100.570 147.635 100.900 148.615 ;
        RECT 101.070 147.465 101.280 148.605 ;
        RECT 101.885 148.445 102.065 149.305 ;
        RECT 102.785 149.105 103.035 149.755 ;
        RECT 102.235 148.775 103.035 149.105 ;
        RECT 101.885 147.975 102.140 148.445 ;
        RECT 101.800 147.805 102.140 147.975 ;
        RECT 101.885 147.775 102.140 147.805 ;
        RECT 102.320 147.465 102.605 148.265 ;
        RECT 102.785 148.185 103.035 148.775 ;
        RECT 103.235 149.420 103.555 149.750 ;
        RECT 103.735 149.535 104.395 150.015 ;
        RECT 104.595 149.625 105.445 149.795 ;
        RECT 103.235 148.525 103.425 149.420 ;
        RECT 103.745 149.095 104.405 149.365 ;
        RECT 104.075 149.035 104.405 149.095 ;
        RECT 103.595 148.865 103.925 148.925 ;
        RECT 104.595 148.865 104.765 149.625 ;
        RECT 106.005 149.555 106.325 150.015 ;
        RECT 106.525 149.375 106.775 149.805 ;
        RECT 107.065 149.575 107.475 150.015 ;
        RECT 107.645 149.635 108.660 149.835 ;
        RECT 104.935 149.205 106.185 149.375 ;
        RECT 104.935 149.085 105.265 149.205 ;
        RECT 103.595 148.695 105.495 148.865 ;
        RECT 103.235 148.355 105.155 148.525 ;
        RECT 103.235 148.335 103.555 148.355 ;
        RECT 102.785 147.675 103.115 148.185 ;
        RECT 103.385 147.725 103.555 148.335 ;
        RECT 105.325 148.185 105.495 148.695 ;
        RECT 105.665 148.625 105.845 149.035 ;
        RECT 106.015 148.445 106.185 149.205 ;
        RECT 103.725 147.465 104.055 148.155 ;
        RECT 104.285 148.015 105.495 148.185 ;
        RECT 105.665 148.135 106.185 148.445 ;
        RECT 106.355 149.035 106.775 149.375 ;
        RECT 107.065 149.035 107.475 149.365 ;
        RECT 106.355 148.265 106.545 149.035 ;
        RECT 107.645 148.905 107.815 149.635 ;
        RECT 108.960 149.465 109.130 149.795 ;
        RECT 109.300 149.635 109.630 150.015 ;
        RECT 107.985 149.085 108.335 149.455 ;
        RECT 107.645 148.865 108.065 148.905 ;
        RECT 106.715 148.695 108.065 148.865 ;
        RECT 106.715 148.535 106.965 148.695 ;
        RECT 107.475 148.265 107.725 148.525 ;
        RECT 106.355 148.015 107.725 148.265 ;
        RECT 104.285 147.725 104.525 148.015 ;
        RECT 105.325 147.935 105.495 148.015 ;
        RECT 104.725 147.465 105.145 147.845 ;
        RECT 105.325 147.685 105.955 147.935 ;
        RECT 106.425 147.465 106.755 147.845 ;
        RECT 106.925 147.725 107.095 148.015 ;
        RECT 107.895 147.850 108.065 148.695 ;
        RECT 108.515 148.525 108.735 149.395 ;
        RECT 108.960 149.275 109.655 149.465 ;
        RECT 108.235 148.145 108.735 148.525 ;
        RECT 108.905 148.475 109.315 149.095 ;
        RECT 109.485 148.305 109.655 149.275 ;
        RECT 108.960 148.135 109.655 148.305 ;
        RECT 107.275 147.465 107.655 147.845 ;
        RECT 107.895 147.680 108.725 147.850 ;
        RECT 108.960 147.635 109.130 148.135 ;
        RECT 109.300 147.465 109.630 147.965 ;
        RECT 109.845 147.635 110.070 149.755 ;
        RECT 110.240 149.635 110.570 150.015 ;
        RECT 110.740 149.465 110.910 149.755 ;
        RECT 110.245 149.295 110.910 149.465 ;
        RECT 110.245 148.305 110.475 149.295 ;
        RECT 111.170 149.265 112.380 150.015 ;
        RECT 110.645 148.475 110.995 149.125 ;
        RECT 111.170 148.555 111.690 149.095 ;
        RECT 111.860 148.725 112.380 149.265 ;
        RECT 110.245 148.135 110.910 148.305 ;
        RECT 110.240 147.465 110.570 147.965 ;
        RECT 110.740 147.635 110.910 148.135 ;
        RECT 111.170 147.465 112.380 148.555 ;
        RECT 18.165 147.295 112.465 147.465 ;
        RECT 18.250 146.205 19.460 147.295 ;
        RECT 18.250 145.495 18.770 146.035 ;
        RECT 18.940 145.665 19.460 146.205 ;
        RECT 19.630 146.205 20.840 147.295 ;
        RECT 19.630 145.665 20.150 146.205 ;
        RECT 21.015 146.105 21.270 146.985 ;
        RECT 21.440 146.155 21.745 147.295 ;
        RECT 22.085 146.915 22.415 147.295 ;
        RECT 22.595 146.745 22.765 147.035 ;
        RECT 22.935 146.835 23.185 147.295 ;
        RECT 21.965 146.575 22.765 146.745 ;
        RECT 23.355 146.785 24.225 147.125 ;
        RECT 20.320 145.495 20.840 146.035 ;
        RECT 18.250 144.745 19.460 145.495 ;
        RECT 19.630 144.745 20.840 145.495 ;
        RECT 21.015 145.455 21.225 146.105 ;
        RECT 21.965 145.985 22.135 146.575 ;
        RECT 23.355 146.405 23.525 146.785 ;
        RECT 24.460 146.665 24.630 147.125 ;
        RECT 24.800 146.835 25.170 147.295 ;
        RECT 25.465 146.695 25.635 147.035 ;
        RECT 25.805 146.865 26.135 147.295 ;
        RECT 26.370 146.695 26.540 147.035 ;
        RECT 22.305 146.235 23.525 146.405 ;
        RECT 23.695 146.325 24.155 146.615 ;
        RECT 24.460 146.495 25.020 146.665 ;
        RECT 25.465 146.525 26.540 146.695 ;
        RECT 26.710 146.795 27.390 147.125 ;
        RECT 27.605 146.795 27.855 147.125 ;
        RECT 28.025 146.835 28.275 147.295 ;
        RECT 24.850 146.355 25.020 146.495 ;
        RECT 23.695 146.315 24.660 146.325 ;
        RECT 23.355 146.145 23.525 146.235 ;
        RECT 23.985 146.155 24.660 146.315 ;
        RECT 21.395 145.955 22.135 145.985 ;
        RECT 21.395 145.655 22.310 145.955 ;
        RECT 21.985 145.480 22.310 145.655 ;
        RECT 21.015 144.925 21.270 145.455 ;
        RECT 21.440 144.745 21.745 145.205 ;
        RECT 21.990 145.125 22.310 145.480 ;
        RECT 22.480 145.695 23.020 146.065 ;
        RECT 23.355 145.975 23.760 146.145 ;
        RECT 22.480 145.295 22.720 145.695 ;
        RECT 23.200 145.525 23.420 145.805 ;
        RECT 22.890 145.355 23.420 145.525 ;
        RECT 22.890 145.125 23.060 145.355 ;
        RECT 23.590 145.195 23.760 145.975 ;
        RECT 23.930 145.365 24.280 145.985 ;
        RECT 24.450 145.365 24.660 146.155 ;
        RECT 24.850 146.185 26.350 146.355 ;
        RECT 24.850 145.495 25.020 146.185 ;
        RECT 26.710 146.015 26.880 146.795 ;
        RECT 27.685 146.665 27.855 146.795 ;
        RECT 25.190 145.845 26.880 146.015 ;
        RECT 27.050 146.235 27.515 146.625 ;
        RECT 27.685 146.495 28.080 146.665 ;
        RECT 25.190 145.665 25.360 145.845 ;
        RECT 21.990 144.955 23.060 145.125 ;
        RECT 23.230 144.745 23.420 145.185 ;
        RECT 23.590 144.915 24.540 145.195 ;
        RECT 24.850 145.105 25.110 145.495 ;
        RECT 25.530 145.425 26.320 145.675 ;
        RECT 24.760 144.935 25.110 145.105 ;
        RECT 25.320 144.745 25.650 145.205 ;
        RECT 26.525 145.135 26.695 145.845 ;
        RECT 27.050 145.645 27.220 146.235 ;
        RECT 26.865 145.425 27.220 145.645 ;
        RECT 27.390 145.425 27.740 146.045 ;
        RECT 27.910 145.135 28.080 146.495 ;
        RECT 28.445 146.325 28.770 147.110 ;
        RECT 28.250 145.275 28.710 146.325 ;
        RECT 26.525 144.965 27.380 145.135 ;
        RECT 27.585 144.965 28.080 145.135 ;
        RECT 28.250 144.745 28.580 145.105 ;
        RECT 28.940 145.005 29.110 147.125 ;
        RECT 29.280 146.795 29.610 147.295 ;
        RECT 29.780 146.625 30.035 147.125 ;
        RECT 29.285 146.455 30.035 146.625 ;
        RECT 29.285 145.465 29.515 146.455 ;
        RECT 29.685 145.635 30.035 146.285 ;
        RECT 30.210 146.220 30.480 147.125 ;
        RECT 30.650 146.535 30.980 147.295 ;
        RECT 31.160 146.365 31.330 147.125 ;
        RECT 29.285 145.295 30.035 145.465 ;
        RECT 29.280 144.745 29.610 145.125 ;
        RECT 29.780 145.005 30.035 145.295 ;
        RECT 30.210 145.420 30.380 146.220 ;
        RECT 30.665 146.195 31.330 146.365 ;
        RECT 30.665 146.050 30.835 146.195 ;
        RECT 32.090 146.155 32.320 147.295 ;
        RECT 32.490 146.145 32.820 147.125 ;
        RECT 32.990 146.155 33.200 147.295 ;
        RECT 33.430 146.220 33.700 147.125 ;
        RECT 33.870 146.535 34.200 147.295 ;
        RECT 34.380 146.365 34.550 147.125 ;
        RECT 30.550 145.720 30.835 146.050 ;
        RECT 30.665 145.465 30.835 145.720 ;
        RECT 31.070 145.645 31.400 146.015 ;
        RECT 32.070 145.735 32.400 145.985 ;
        RECT 30.210 144.915 30.470 145.420 ;
        RECT 30.665 145.295 31.330 145.465 ;
        RECT 30.650 144.745 30.980 145.125 ;
        RECT 31.160 144.915 31.330 145.295 ;
        RECT 32.090 144.745 32.320 145.565 ;
        RECT 32.570 145.545 32.820 146.145 ;
        RECT 32.490 144.915 32.820 145.545 ;
        RECT 32.990 144.745 33.200 145.565 ;
        RECT 33.430 145.420 33.600 146.220 ;
        RECT 33.885 146.195 34.550 146.365 ;
        RECT 33.885 146.050 34.055 146.195 ;
        RECT 34.810 146.130 35.100 147.295 ;
        RECT 35.275 146.155 35.610 147.125 ;
        RECT 35.780 146.155 35.950 147.295 ;
        RECT 36.120 146.955 38.150 147.125 ;
        RECT 33.770 145.720 34.055 146.050 ;
        RECT 33.885 145.465 34.055 145.720 ;
        RECT 34.290 145.645 34.620 146.015 ;
        RECT 35.275 145.485 35.445 146.155 ;
        RECT 36.120 145.985 36.290 146.955 ;
        RECT 35.615 145.655 35.870 145.985 ;
        RECT 36.095 145.655 36.290 145.985 ;
        RECT 36.460 146.615 37.585 146.785 ;
        RECT 35.700 145.485 35.870 145.655 ;
        RECT 36.460 145.485 36.630 146.615 ;
        RECT 33.430 144.915 33.690 145.420 ;
        RECT 33.885 145.295 34.550 145.465 ;
        RECT 33.870 144.745 34.200 145.125 ;
        RECT 34.380 144.915 34.550 145.295 ;
        RECT 34.810 144.745 35.100 145.470 ;
        RECT 35.275 144.915 35.530 145.485 ;
        RECT 35.700 145.315 36.630 145.485 ;
        RECT 36.800 146.275 37.810 146.445 ;
        RECT 36.800 145.475 36.970 146.275 ;
        RECT 37.175 145.935 37.450 146.075 ;
        RECT 37.170 145.765 37.450 145.935 ;
        RECT 36.455 145.280 36.630 145.315 ;
        RECT 35.700 144.745 36.030 145.145 ;
        RECT 36.455 144.915 36.985 145.280 ;
        RECT 37.175 144.915 37.450 145.765 ;
        RECT 37.620 144.915 37.810 146.275 ;
        RECT 37.980 146.290 38.150 146.955 ;
        RECT 38.320 146.535 38.490 147.295 ;
        RECT 38.725 146.535 39.240 146.945 ;
        RECT 37.980 146.100 38.730 146.290 ;
        RECT 38.900 145.725 39.240 146.535 ;
        RECT 38.010 145.555 39.240 145.725 ;
        RECT 39.410 146.205 41.080 147.295 ;
        RECT 39.410 145.685 40.160 146.205 ;
        RECT 41.250 146.155 41.590 147.125 ;
        RECT 41.760 146.155 41.930 147.295 ;
        RECT 42.200 146.495 42.450 147.295 ;
        RECT 43.095 146.325 43.425 147.125 ;
        RECT 43.725 146.495 44.055 147.295 ;
        RECT 44.225 146.325 44.555 147.125 ;
        RECT 42.120 146.155 44.555 146.325 ;
        RECT 44.930 146.155 45.270 147.125 ;
        RECT 45.440 146.155 45.610 147.295 ;
        RECT 45.880 146.495 46.130 147.295 ;
        RECT 46.775 146.325 47.105 147.125 ;
        RECT 47.405 146.495 47.735 147.295 ;
        RECT 47.905 146.325 48.235 147.125 ;
        RECT 45.800 146.155 48.235 146.325 ;
        RECT 49.070 146.155 49.410 147.125 ;
        RECT 49.580 146.155 49.750 147.295 ;
        RECT 50.020 146.495 50.270 147.295 ;
        RECT 50.915 146.325 51.245 147.125 ;
        RECT 51.545 146.495 51.875 147.295 ;
        RECT 52.045 146.325 52.375 147.125 ;
        RECT 52.865 146.665 53.150 147.125 ;
        RECT 53.320 146.835 53.590 147.295 ;
        RECT 52.865 146.445 53.820 146.665 ;
        RECT 49.940 146.155 52.375 146.325 ;
        RECT 37.990 144.745 38.500 145.280 ;
        RECT 38.720 144.950 38.965 145.555 ;
        RECT 40.330 145.515 41.080 146.035 ;
        RECT 39.410 144.745 41.080 145.515 ;
        RECT 41.250 145.595 41.425 146.155 ;
        RECT 42.120 145.905 42.290 146.155 ;
        RECT 41.595 145.735 42.290 145.905 ;
        RECT 42.465 145.735 42.885 145.935 ;
        RECT 43.055 145.735 43.385 145.935 ;
        RECT 43.555 145.735 43.885 145.935 ;
        RECT 41.250 145.545 41.480 145.595 ;
        RECT 41.250 144.915 41.590 145.545 ;
        RECT 41.760 144.745 42.010 145.545 ;
        RECT 42.200 145.395 43.425 145.565 ;
        RECT 42.200 144.915 42.530 145.395 ;
        RECT 42.700 144.745 42.925 145.205 ;
        RECT 43.095 144.915 43.425 145.395 ;
        RECT 44.055 145.525 44.225 146.155 ;
        RECT 44.410 145.735 44.760 145.985 ;
        RECT 44.930 145.545 45.105 146.155 ;
        RECT 45.800 145.905 45.970 146.155 ;
        RECT 45.275 145.735 45.970 145.905 ;
        RECT 46.145 145.735 46.565 145.935 ;
        RECT 46.735 145.735 47.065 145.935 ;
        RECT 47.235 145.735 47.565 145.935 ;
        RECT 44.055 144.915 44.555 145.525 ;
        RECT 44.930 144.915 45.270 145.545 ;
        RECT 45.440 144.745 45.690 145.545 ;
        RECT 45.880 145.395 47.105 145.565 ;
        RECT 45.880 144.915 46.210 145.395 ;
        RECT 46.380 144.745 46.605 145.205 ;
        RECT 46.775 144.915 47.105 145.395 ;
        RECT 47.735 145.525 47.905 146.155 ;
        RECT 49.070 146.105 49.300 146.155 ;
        RECT 48.090 145.735 48.440 145.985 ;
        RECT 49.070 145.545 49.245 146.105 ;
        RECT 49.940 145.905 50.110 146.155 ;
        RECT 49.415 145.735 50.110 145.905 ;
        RECT 50.285 145.735 50.705 145.935 ;
        RECT 50.875 145.735 51.205 145.935 ;
        RECT 51.375 145.735 51.705 145.935 ;
        RECT 47.735 144.915 48.235 145.525 ;
        RECT 49.070 144.915 49.410 145.545 ;
        RECT 49.580 144.745 49.830 145.545 ;
        RECT 50.020 145.395 51.245 145.565 ;
        RECT 50.020 144.915 50.350 145.395 ;
        RECT 50.520 144.745 50.745 145.205 ;
        RECT 50.915 144.915 51.245 145.395 ;
        RECT 51.875 145.525 52.045 146.155 ;
        RECT 52.230 145.735 52.580 145.985 ;
        RECT 52.750 145.715 53.440 146.275 ;
        RECT 53.610 145.545 53.820 146.445 ;
        RECT 51.875 144.915 52.375 145.525 ;
        RECT 52.865 145.375 53.820 145.545 ;
        RECT 53.990 146.275 54.390 147.125 ;
        RECT 54.580 146.665 54.860 147.125 ;
        RECT 55.380 146.835 55.705 147.295 ;
        RECT 54.580 146.445 55.705 146.665 ;
        RECT 53.990 145.715 55.085 146.275 ;
        RECT 55.255 145.985 55.705 146.445 ;
        RECT 55.875 146.155 56.260 147.125 ;
        RECT 52.865 144.915 53.150 145.375 ;
        RECT 53.320 144.745 53.590 145.205 ;
        RECT 53.990 144.915 54.390 145.715 ;
        RECT 55.255 145.655 55.810 145.985 ;
        RECT 55.255 145.545 55.705 145.655 ;
        RECT 54.580 145.375 55.705 145.545 ;
        RECT 55.980 145.485 56.260 146.155 ;
        RECT 56.430 146.535 56.945 146.945 ;
        RECT 57.180 146.535 57.350 147.295 ;
        RECT 57.520 146.955 59.550 147.125 ;
        RECT 56.430 145.725 56.770 146.535 ;
        RECT 57.520 146.290 57.690 146.955 ;
        RECT 58.085 146.615 59.210 146.785 ;
        RECT 56.940 146.100 57.690 146.290 ;
        RECT 57.860 146.275 58.870 146.445 ;
        RECT 56.430 145.555 57.660 145.725 ;
        RECT 54.580 144.915 54.860 145.375 ;
        RECT 55.380 144.745 55.705 145.205 ;
        RECT 55.875 144.915 56.260 145.485 ;
        RECT 56.705 144.950 56.950 145.555 ;
        RECT 57.170 144.745 57.680 145.280 ;
        RECT 57.860 144.915 58.050 146.275 ;
        RECT 58.220 145.935 58.495 146.075 ;
        RECT 58.220 145.765 58.500 145.935 ;
        RECT 58.220 144.915 58.495 145.765 ;
        RECT 58.700 145.475 58.870 146.275 ;
        RECT 59.040 145.485 59.210 146.615 ;
        RECT 59.380 145.985 59.550 146.955 ;
        RECT 59.720 146.155 59.890 147.295 ;
        RECT 60.060 146.155 60.395 147.125 ;
        RECT 59.380 145.655 59.575 145.985 ;
        RECT 59.800 145.655 60.055 145.985 ;
        RECT 59.800 145.485 59.970 145.655 ;
        RECT 60.225 145.485 60.395 146.155 ;
        RECT 60.570 146.130 60.860 147.295 ;
        RECT 61.405 146.315 61.660 146.985 ;
        RECT 61.840 146.495 62.125 147.295 ;
        RECT 62.305 146.575 62.635 147.085 ;
        RECT 61.405 145.935 61.585 146.315 ;
        RECT 62.305 145.985 62.555 146.575 ;
        RECT 62.905 146.425 63.075 147.035 ;
        RECT 63.245 146.605 63.575 147.295 ;
        RECT 63.805 146.745 64.045 147.035 ;
        RECT 64.245 146.915 64.665 147.295 ;
        RECT 64.845 146.825 65.475 147.075 ;
        RECT 65.945 146.915 66.275 147.295 ;
        RECT 64.845 146.745 65.015 146.825 ;
        RECT 66.445 146.745 66.615 147.035 ;
        RECT 66.795 146.915 67.175 147.295 ;
        RECT 67.415 146.910 68.245 147.080 ;
        RECT 63.805 146.575 65.015 146.745 ;
        RECT 61.320 145.765 61.585 145.935 ;
        RECT 59.040 145.315 59.970 145.485 ;
        RECT 59.040 145.280 59.215 145.315 ;
        RECT 58.685 144.915 59.215 145.280 ;
        RECT 59.640 144.745 59.970 145.145 ;
        RECT 60.140 144.915 60.395 145.485 ;
        RECT 60.570 144.745 60.860 145.470 ;
        RECT 61.405 145.455 61.585 145.765 ;
        RECT 61.755 145.655 62.555 145.985 ;
        RECT 61.405 144.925 61.660 145.455 ;
        RECT 61.840 144.745 62.125 145.205 ;
        RECT 62.305 145.005 62.555 145.655 ;
        RECT 62.755 146.405 63.075 146.425 ;
        RECT 62.755 146.235 64.675 146.405 ;
        RECT 62.755 145.340 62.945 146.235 ;
        RECT 64.845 146.065 65.015 146.575 ;
        RECT 65.185 146.315 65.705 146.625 ;
        RECT 63.115 145.895 65.015 146.065 ;
        RECT 63.115 145.835 63.445 145.895 ;
        RECT 63.595 145.665 63.925 145.725 ;
        RECT 63.265 145.395 63.925 145.665 ;
        RECT 62.755 145.010 63.075 145.340 ;
        RECT 63.255 144.745 63.915 145.225 ;
        RECT 64.115 145.135 64.285 145.895 ;
        RECT 65.185 145.725 65.365 146.135 ;
        RECT 64.455 145.555 64.785 145.675 ;
        RECT 65.535 145.555 65.705 146.315 ;
        RECT 64.455 145.385 65.705 145.555 ;
        RECT 65.875 146.495 67.245 146.745 ;
        RECT 65.875 145.725 66.065 146.495 ;
        RECT 66.995 146.235 67.245 146.495 ;
        RECT 66.235 146.065 66.485 146.225 ;
        RECT 67.415 146.065 67.585 146.910 ;
        RECT 68.480 146.625 68.650 147.125 ;
        RECT 68.820 146.795 69.150 147.295 ;
        RECT 67.755 146.235 68.255 146.615 ;
        RECT 68.480 146.455 69.175 146.625 ;
        RECT 66.235 145.895 67.585 146.065 ;
        RECT 67.165 145.855 67.585 145.895 ;
        RECT 65.875 145.385 66.295 145.725 ;
        RECT 66.585 145.395 66.995 145.725 ;
        RECT 64.115 144.965 64.965 145.135 ;
        RECT 65.525 144.745 65.845 145.205 ;
        RECT 66.045 144.955 66.295 145.385 ;
        RECT 66.585 144.745 66.995 145.185 ;
        RECT 67.165 145.125 67.335 145.855 ;
        RECT 67.505 145.305 67.855 145.675 ;
        RECT 68.035 145.365 68.255 146.235 ;
        RECT 68.425 145.665 68.835 146.285 ;
        RECT 69.005 145.485 69.175 146.455 ;
        RECT 68.480 145.295 69.175 145.485 ;
        RECT 67.165 144.925 68.180 145.125 ;
        RECT 68.480 144.965 68.650 145.295 ;
        RECT 68.820 144.745 69.150 145.125 ;
        RECT 69.365 145.005 69.590 147.125 ;
        RECT 69.760 146.795 70.090 147.295 ;
        RECT 70.260 146.625 70.430 147.125 ;
        RECT 71.615 146.860 76.960 147.295 ;
        RECT 69.765 146.455 70.430 146.625 ;
        RECT 69.765 145.465 69.995 146.455 ;
        RECT 70.165 145.635 70.515 146.285 ;
        RECT 73.205 145.610 73.555 146.860 ;
        RECT 69.765 145.295 70.430 145.465 ;
        RECT 69.760 144.745 70.090 145.125 ;
        RECT 70.260 145.005 70.430 145.295 ;
        RECT 75.035 145.290 75.375 146.120 ;
        RECT 77.135 146.105 77.390 146.985 ;
        RECT 77.560 146.155 77.865 147.295 ;
        RECT 78.205 146.915 78.535 147.295 ;
        RECT 78.715 146.745 78.885 147.035 ;
        RECT 79.055 146.835 79.305 147.295 ;
        RECT 78.085 146.575 78.885 146.745 ;
        RECT 79.475 146.785 80.345 147.125 ;
        RECT 77.135 145.455 77.345 146.105 ;
        RECT 78.085 145.985 78.255 146.575 ;
        RECT 79.475 146.405 79.645 146.785 ;
        RECT 80.580 146.665 80.750 147.125 ;
        RECT 80.920 146.835 81.290 147.295 ;
        RECT 81.585 146.695 81.755 147.035 ;
        RECT 81.925 146.865 82.255 147.295 ;
        RECT 82.490 146.695 82.660 147.035 ;
        RECT 78.425 146.235 79.645 146.405 ;
        RECT 79.815 146.325 80.275 146.615 ;
        RECT 80.580 146.495 81.140 146.665 ;
        RECT 81.585 146.525 82.660 146.695 ;
        RECT 82.830 146.795 83.510 147.125 ;
        RECT 83.725 146.795 83.975 147.125 ;
        RECT 84.145 146.835 84.395 147.295 ;
        RECT 80.970 146.355 81.140 146.495 ;
        RECT 79.815 146.315 80.780 146.325 ;
        RECT 79.475 146.145 79.645 146.235 ;
        RECT 80.105 146.155 80.780 146.315 ;
        RECT 77.515 145.955 78.255 145.985 ;
        RECT 77.515 145.655 78.430 145.955 ;
        RECT 78.105 145.480 78.430 145.655 ;
        RECT 71.615 144.745 76.960 145.290 ;
        RECT 77.135 144.925 77.390 145.455 ;
        RECT 77.560 144.745 77.865 145.205 ;
        RECT 78.110 145.125 78.430 145.480 ;
        RECT 78.600 145.695 79.140 146.065 ;
        RECT 79.475 145.975 79.880 146.145 ;
        RECT 78.600 145.295 78.840 145.695 ;
        RECT 79.320 145.525 79.540 145.805 ;
        RECT 79.010 145.355 79.540 145.525 ;
        RECT 79.010 145.125 79.180 145.355 ;
        RECT 79.710 145.195 79.880 145.975 ;
        RECT 80.050 145.365 80.400 145.985 ;
        RECT 80.570 145.365 80.780 146.155 ;
        RECT 80.970 146.185 82.470 146.355 ;
        RECT 80.970 145.495 81.140 146.185 ;
        RECT 82.830 146.015 83.000 146.795 ;
        RECT 83.805 146.665 83.975 146.795 ;
        RECT 81.310 145.845 83.000 146.015 ;
        RECT 83.170 146.235 83.635 146.625 ;
        RECT 83.805 146.495 84.200 146.665 ;
        RECT 81.310 145.665 81.480 145.845 ;
        RECT 78.110 144.955 79.180 145.125 ;
        RECT 79.350 144.745 79.540 145.185 ;
        RECT 79.710 144.915 80.660 145.195 ;
        RECT 80.970 145.105 81.230 145.495 ;
        RECT 81.650 145.425 82.440 145.675 ;
        RECT 80.880 144.935 81.230 145.105 ;
        RECT 81.440 144.745 81.770 145.205 ;
        RECT 82.645 145.135 82.815 145.845 ;
        RECT 83.170 145.645 83.340 146.235 ;
        RECT 82.985 145.425 83.340 145.645 ;
        RECT 83.510 145.425 83.860 146.045 ;
        RECT 84.030 145.135 84.200 146.495 ;
        RECT 84.565 146.325 84.890 147.110 ;
        RECT 84.370 145.275 84.830 146.325 ;
        RECT 82.645 144.965 83.500 145.135 ;
        RECT 83.705 144.965 84.200 145.135 ;
        RECT 84.370 144.745 84.700 145.105 ;
        RECT 85.060 145.005 85.230 147.125 ;
        RECT 85.400 146.795 85.730 147.295 ;
        RECT 85.900 146.625 86.155 147.125 ;
        RECT 85.405 146.455 86.155 146.625 ;
        RECT 85.405 145.465 85.635 146.455 ;
        RECT 85.805 145.635 86.155 146.285 ;
        RECT 86.330 146.130 86.620 147.295 ;
        RECT 87.455 146.325 87.785 147.125 ;
        RECT 87.955 146.495 88.285 147.295 ;
        RECT 88.585 146.325 88.915 147.125 ;
        RECT 89.560 146.495 89.810 147.295 ;
        RECT 87.455 146.155 89.890 146.325 ;
        RECT 90.080 146.155 90.250 147.295 ;
        RECT 90.420 146.155 90.760 147.125 ;
        RECT 87.250 145.735 87.600 145.985 ;
        RECT 87.785 145.525 87.955 146.155 ;
        RECT 88.125 145.735 88.455 145.935 ;
        RECT 88.625 145.735 88.955 145.935 ;
        RECT 89.125 145.735 89.545 145.935 ;
        RECT 89.720 145.905 89.890 146.155 ;
        RECT 89.720 145.735 90.415 145.905 ;
        RECT 85.405 145.295 86.155 145.465 ;
        RECT 85.400 144.745 85.730 145.125 ;
        RECT 85.900 145.005 86.155 145.295 ;
        RECT 86.330 144.745 86.620 145.470 ;
        RECT 87.455 144.915 87.955 145.525 ;
        RECT 88.585 145.395 89.810 145.565 ;
        RECT 90.585 145.545 90.760 146.155 ;
        RECT 90.930 146.205 92.600 147.295 ;
        RECT 92.975 146.325 93.305 147.125 ;
        RECT 93.475 146.495 93.805 147.295 ;
        RECT 94.105 146.325 94.435 147.125 ;
        RECT 95.080 146.495 95.330 147.295 ;
        RECT 90.930 145.685 91.680 146.205 ;
        RECT 92.975 146.155 95.410 146.325 ;
        RECT 95.600 146.155 95.770 147.295 ;
        RECT 95.940 146.155 96.280 147.125 ;
        RECT 88.585 144.915 88.915 145.395 ;
        RECT 89.085 144.745 89.310 145.205 ;
        RECT 89.480 144.915 89.810 145.395 ;
        RECT 90.000 144.745 90.250 145.545 ;
        RECT 90.420 144.915 90.760 145.545 ;
        RECT 91.850 145.515 92.600 146.035 ;
        RECT 92.770 145.735 93.120 145.985 ;
        RECT 93.305 145.525 93.475 146.155 ;
        RECT 93.645 145.735 93.975 145.935 ;
        RECT 94.145 145.735 94.475 145.935 ;
        RECT 94.645 145.735 95.065 145.935 ;
        RECT 95.240 145.905 95.410 146.155 ;
        RECT 95.240 145.735 95.935 145.905 ;
        RECT 90.930 144.745 92.600 145.515 ;
        RECT 92.975 144.915 93.475 145.525 ;
        RECT 94.105 145.395 95.330 145.565 ;
        RECT 96.105 145.545 96.280 146.155 ;
        RECT 96.450 146.205 97.660 147.295 ;
        RECT 96.450 145.665 96.970 146.205 ;
        RECT 97.830 146.155 98.170 147.125 ;
        RECT 98.340 146.155 98.510 147.295 ;
        RECT 98.780 146.495 99.030 147.295 ;
        RECT 99.675 146.325 100.005 147.125 ;
        RECT 100.305 146.495 100.635 147.295 ;
        RECT 100.805 146.325 101.135 147.125 ;
        RECT 98.700 146.155 101.135 146.325 ;
        RECT 101.510 146.535 102.025 146.945 ;
        RECT 102.260 146.535 102.430 147.295 ;
        RECT 102.600 146.955 104.630 147.125 ;
        RECT 94.105 144.915 94.435 145.395 ;
        RECT 94.605 144.745 94.830 145.205 ;
        RECT 95.000 144.915 95.330 145.395 ;
        RECT 95.520 144.745 95.770 145.545 ;
        RECT 95.940 144.915 96.280 145.545 ;
        RECT 97.140 145.495 97.660 146.035 ;
        RECT 96.450 144.745 97.660 145.495 ;
        RECT 97.830 145.545 98.005 146.155 ;
        RECT 98.700 145.905 98.870 146.155 ;
        RECT 98.175 145.735 98.870 145.905 ;
        RECT 99.045 145.735 99.465 145.935 ;
        RECT 99.635 145.735 99.965 145.935 ;
        RECT 100.135 145.735 100.465 145.935 ;
        RECT 97.830 144.915 98.170 145.545 ;
        RECT 98.340 144.745 98.590 145.545 ;
        RECT 98.780 145.395 100.005 145.565 ;
        RECT 98.780 144.915 99.110 145.395 ;
        RECT 99.280 144.745 99.505 145.205 ;
        RECT 99.675 144.915 100.005 145.395 ;
        RECT 100.635 145.525 100.805 146.155 ;
        RECT 100.990 145.735 101.340 145.985 ;
        RECT 101.510 145.725 101.850 146.535 ;
        RECT 102.600 146.290 102.770 146.955 ;
        RECT 103.165 146.615 104.290 146.785 ;
        RECT 102.020 146.100 102.770 146.290 ;
        RECT 102.940 146.275 103.950 146.445 ;
        RECT 101.510 145.555 102.740 145.725 ;
        RECT 100.635 144.915 101.135 145.525 ;
        RECT 101.785 144.950 102.030 145.555 ;
        RECT 102.250 144.745 102.760 145.280 ;
        RECT 102.940 144.915 103.130 146.275 ;
        RECT 103.300 145.935 103.575 146.075 ;
        RECT 103.300 145.765 103.580 145.935 ;
        RECT 103.300 144.915 103.575 145.765 ;
        RECT 103.780 145.475 103.950 146.275 ;
        RECT 104.120 145.485 104.290 146.615 ;
        RECT 104.460 145.985 104.630 146.955 ;
        RECT 104.800 146.155 104.970 147.295 ;
        RECT 105.140 146.155 105.475 147.125 ;
        RECT 105.710 146.155 105.920 147.295 ;
        RECT 104.460 145.655 104.655 145.985 ;
        RECT 104.880 145.655 105.135 145.985 ;
        RECT 104.880 145.485 105.050 145.655 ;
        RECT 105.305 145.485 105.475 146.155 ;
        RECT 106.090 146.145 106.420 147.125 ;
        RECT 106.590 146.155 106.820 147.295 ;
        RECT 107.120 146.365 107.290 147.125 ;
        RECT 107.470 146.535 107.800 147.295 ;
        RECT 107.120 146.195 107.785 146.365 ;
        RECT 107.970 146.220 108.240 147.125 ;
        RECT 104.120 145.315 105.050 145.485 ;
        RECT 104.120 145.280 104.295 145.315 ;
        RECT 103.765 144.915 104.295 145.280 ;
        RECT 104.720 144.745 105.050 145.145 ;
        RECT 105.220 144.915 105.475 145.485 ;
        RECT 105.710 144.745 105.920 145.565 ;
        RECT 106.090 145.545 106.340 146.145 ;
        RECT 107.615 146.050 107.785 146.195 ;
        RECT 106.510 145.735 106.840 145.985 ;
        RECT 107.050 145.645 107.380 146.015 ;
        RECT 107.615 145.720 107.900 146.050 ;
        RECT 106.090 144.915 106.420 145.545 ;
        RECT 106.590 144.745 106.820 145.565 ;
        RECT 107.615 145.465 107.785 145.720 ;
        RECT 107.120 145.295 107.785 145.465 ;
        RECT 108.070 145.420 108.240 146.220 ;
        RECT 108.500 146.365 108.670 147.125 ;
        RECT 108.850 146.535 109.180 147.295 ;
        RECT 108.500 146.195 109.165 146.365 ;
        RECT 109.350 146.220 109.620 147.125 ;
        RECT 108.995 146.050 109.165 146.195 ;
        RECT 108.430 145.645 108.760 146.015 ;
        RECT 108.995 145.720 109.280 146.050 ;
        RECT 108.995 145.465 109.165 145.720 ;
        RECT 107.120 144.915 107.290 145.295 ;
        RECT 107.470 144.745 107.800 145.125 ;
        RECT 107.980 144.915 108.240 145.420 ;
        RECT 108.500 145.295 109.165 145.465 ;
        RECT 109.450 145.420 109.620 146.220 ;
        RECT 109.790 146.205 111.000 147.295 ;
        RECT 111.170 146.205 112.380 147.295 ;
        RECT 109.790 145.665 110.310 146.205 ;
        RECT 110.480 145.495 111.000 146.035 ;
        RECT 111.170 145.665 111.690 146.205 ;
        RECT 111.860 145.495 112.380 146.035 ;
        RECT 108.500 144.915 108.670 145.295 ;
        RECT 108.850 144.745 109.180 145.125 ;
        RECT 109.360 144.915 109.620 145.420 ;
        RECT 109.790 144.745 111.000 145.495 ;
        RECT 111.170 144.745 112.380 145.495 ;
        RECT 18.165 144.575 112.465 144.745 ;
        RECT 18.250 143.825 19.460 144.575 ;
        RECT 18.250 143.285 18.770 143.825 ;
        RECT 20.090 143.805 21.760 144.575 ;
        RECT 21.930 143.850 22.220 144.575 ;
        RECT 22.390 143.805 24.980 144.575 ;
        RECT 18.940 143.115 19.460 143.655 ;
        RECT 18.250 142.025 19.460 143.115 ;
        RECT 20.090 143.115 20.840 143.635 ;
        RECT 21.010 143.285 21.760 143.805 ;
        RECT 20.090 142.025 21.760 143.115 ;
        RECT 21.930 142.025 22.220 143.190 ;
        RECT 22.390 143.115 23.600 143.635 ;
        RECT 23.770 143.285 24.980 143.805 ;
        RECT 25.425 143.765 25.670 144.370 ;
        RECT 25.890 144.040 26.400 144.575 ;
        RECT 25.150 143.595 26.380 143.765 ;
        RECT 22.390 142.025 24.980 143.115 ;
        RECT 25.150 142.785 25.490 143.595 ;
        RECT 25.660 143.030 26.410 143.220 ;
        RECT 25.150 142.375 25.665 142.785 ;
        RECT 25.900 142.025 26.070 142.785 ;
        RECT 26.240 142.365 26.410 143.030 ;
        RECT 26.580 143.045 26.770 144.405 ;
        RECT 26.940 143.895 27.215 144.405 ;
        RECT 27.405 144.040 27.935 144.405 ;
        RECT 28.360 144.175 28.690 144.575 ;
        RECT 27.760 144.005 27.935 144.040 ;
        RECT 26.940 143.725 27.220 143.895 ;
        RECT 26.940 143.245 27.215 143.725 ;
        RECT 27.420 143.045 27.590 143.845 ;
        RECT 26.580 142.875 27.590 143.045 ;
        RECT 27.760 143.835 28.690 144.005 ;
        RECT 28.860 143.835 29.115 144.405 ;
        RECT 27.760 142.705 27.930 143.835 ;
        RECT 28.520 143.665 28.690 143.835 ;
        RECT 26.805 142.535 27.930 142.705 ;
        RECT 28.100 143.335 28.295 143.665 ;
        RECT 28.520 143.335 28.775 143.665 ;
        RECT 28.100 142.365 28.270 143.335 ;
        RECT 28.945 143.165 29.115 143.835 ;
        RECT 30.250 143.755 30.480 144.575 ;
        RECT 30.650 143.775 30.980 144.405 ;
        RECT 30.230 143.335 30.560 143.585 ;
        RECT 30.730 143.175 30.980 143.775 ;
        RECT 31.150 143.755 31.360 144.575 ;
        RECT 31.595 143.865 31.850 144.395 ;
        RECT 32.020 144.115 32.325 144.575 ;
        RECT 32.570 144.195 33.640 144.365 ;
        RECT 26.240 142.195 28.270 142.365 ;
        RECT 28.440 142.025 28.610 143.165 ;
        RECT 28.780 142.195 29.115 143.165 ;
        RECT 30.250 142.025 30.480 143.165 ;
        RECT 30.650 142.195 30.980 143.175 ;
        RECT 31.595 143.215 31.805 143.865 ;
        RECT 32.570 143.840 32.890 144.195 ;
        RECT 32.565 143.665 32.890 143.840 ;
        RECT 31.975 143.365 32.890 143.665 ;
        RECT 33.060 143.625 33.300 144.025 ;
        RECT 33.470 143.965 33.640 144.195 ;
        RECT 33.810 144.135 34.000 144.575 ;
        RECT 34.170 144.125 35.120 144.405 ;
        RECT 35.340 144.215 35.690 144.385 ;
        RECT 33.470 143.795 34.000 143.965 ;
        RECT 31.975 143.335 32.715 143.365 ;
        RECT 31.150 142.025 31.360 143.165 ;
        RECT 31.595 142.335 31.850 143.215 ;
        RECT 32.020 142.025 32.325 143.165 ;
        RECT 32.545 142.745 32.715 143.335 ;
        RECT 33.060 143.255 33.600 143.625 ;
        RECT 33.780 143.515 34.000 143.795 ;
        RECT 34.170 143.345 34.340 144.125 ;
        RECT 33.935 143.175 34.340 143.345 ;
        RECT 34.510 143.335 34.860 143.955 ;
        RECT 33.935 143.085 34.105 143.175 ;
        RECT 35.030 143.165 35.240 143.955 ;
        RECT 32.885 142.915 34.105 143.085 ;
        RECT 34.565 143.005 35.240 143.165 ;
        RECT 32.545 142.575 33.345 142.745 ;
        RECT 32.665 142.025 32.995 142.405 ;
        RECT 33.175 142.285 33.345 142.575 ;
        RECT 33.935 142.535 34.105 142.915 ;
        RECT 34.275 142.995 35.240 143.005 ;
        RECT 35.430 143.825 35.690 144.215 ;
        RECT 35.900 144.115 36.230 144.575 ;
        RECT 37.105 144.185 37.960 144.355 ;
        RECT 38.165 144.185 38.660 144.355 ;
        RECT 38.830 144.215 39.160 144.575 ;
        RECT 35.430 143.135 35.600 143.825 ;
        RECT 35.770 143.475 35.940 143.655 ;
        RECT 36.110 143.645 36.900 143.895 ;
        RECT 37.105 143.475 37.275 144.185 ;
        RECT 37.445 143.675 37.800 143.895 ;
        RECT 35.770 143.305 37.460 143.475 ;
        RECT 34.275 142.705 34.735 142.995 ;
        RECT 35.430 142.965 36.930 143.135 ;
        RECT 35.430 142.825 35.600 142.965 ;
        RECT 35.040 142.655 35.600 142.825 ;
        RECT 33.515 142.025 33.765 142.485 ;
        RECT 33.935 142.195 34.805 142.535 ;
        RECT 35.040 142.195 35.210 142.655 ;
        RECT 36.045 142.625 37.120 142.795 ;
        RECT 35.380 142.025 35.750 142.485 ;
        RECT 36.045 142.285 36.215 142.625 ;
        RECT 36.385 142.025 36.715 142.455 ;
        RECT 36.950 142.285 37.120 142.625 ;
        RECT 37.290 142.525 37.460 143.305 ;
        RECT 37.630 143.085 37.800 143.675 ;
        RECT 37.970 143.275 38.320 143.895 ;
        RECT 37.630 142.695 38.095 143.085 ;
        RECT 38.490 142.825 38.660 144.185 ;
        RECT 38.830 142.995 39.290 144.045 ;
        RECT 38.265 142.655 38.660 142.825 ;
        RECT 38.265 142.525 38.435 142.655 ;
        RECT 37.290 142.195 37.970 142.525 ;
        RECT 38.185 142.195 38.435 142.525 ;
        RECT 38.605 142.025 38.855 142.485 ;
        RECT 39.025 142.210 39.350 142.995 ;
        RECT 39.520 142.195 39.690 144.315 ;
        RECT 39.860 144.195 40.190 144.575 ;
        RECT 40.360 144.025 40.615 144.315 ;
        RECT 39.865 143.855 40.615 144.025 ;
        RECT 41.250 143.900 41.520 144.245 ;
        RECT 41.710 144.175 42.090 144.575 ;
        RECT 42.260 144.005 42.430 144.355 ;
        RECT 42.600 144.175 42.930 144.575 ;
        RECT 43.130 144.005 43.300 144.355 ;
        RECT 43.500 144.075 43.830 144.575 ;
        RECT 39.865 142.865 40.095 143.855 ;
        RECT 40.265 143.035 40.615 143.685 ;
        RECT 41.250 143.165 41.420 143.900 ;
        RECT 41.690 143.835 43.300 144.005 ;
        RECT 41.690 143.665 41.860 143.835 ;
        RECT 41.590 143.335 41.860 143.665 ;
        RECT 42.030 143.335 42.435 143.665 ;
        RECT 41.690 143.165 41.860 143.335 ;
        RECT 39.865 142.695 40.615 142.865 ;
        RECT 39.860 142.025 40.190 142.525 ;
        RECT 40.360 142.195 40.615 142.695 ;
        RECT 41.250 142.195 41.520 143.165 ;
        RECT 41.690 142.995 42.415 143.165 ;
        RECT 42.605 143.045 43.315 143.665 ;
        RECT 43.485 143.335 43.835 143.905 ;
        RECT 44.215 143.795 44.715 144.405 ;
        RECT 44.010 143.335 44.360 143.585 ;
        RECT 44.545 143.165 44.715 143.795 ;
        RECT 45.345 143.925 45.675 144.405 ;
        RECT 45.845 144.115 46.070 144.575 ;
        RECT 46.240 143.925 46.570 144.405 ;
        RECT 45.345 143.755 46.570 143.925 ;
        RECT 46.760 143.775 47.010 144.575 ;
        RECT 47.180 143.775 47.520 144.405 ;
        RECT 47.690 143.850 47.980 144.575 ;
        RECT 44.885 143.385 45.215 143.585 ;
        RECT 45.385 143.385 45.715 143.585 ;
        RECT 45.885 143.385 46.305 143.585 ;
        RECT 46.480 143.415 47.175 143.585 ;
        RECT 46.480 143.165 46.650 143.415 ;
        RECT 47.345 143.165 47.520 143.775 ;
        RECT 48.610 143.775 48.950 144.405 ;
        RECT 49.120 143.775 49.370 144.575 ;
        RECT 49.560 143.925 49.890 144.405 ;
        RECT 50.060 144.115 50.285 144.575 ;
        RECT 50.455 143.925 50.785 144.405 ;
        RECT 48.610 143.725 48.840 143.775 ;
        RECT 49.560 143.755 50.785 143.925 ;
        RECT 51.415 143.795 51.915 144.405 ;
        RECT 42.245 142.875 42.415 142.995 ;
        RECT 43.515 142.875 43.835 143.165 ;
        RECT 41.730 142.025 42.010 142.825 ;
        RECT 42.245 142.705 43.835 142.875 ;
        RECT 44.215 142.995 46.650 143.165 ;
        RECT 42.180 142.245 43.835 142.535 ;
        RECT 44.215 142.195 44.545 142.995 ;
        RECT 44.715 142.025 45.045 142.825 ;
        RECT 45.345 142.195 45.675 142.995 ;
        RECT 46.320 142.025 46.570 142.825 ;
        RECT 46.840 142.025 47.010 143.165 ;
        RECT 47.180 142.195 47.520 143.165 ;
        RECT 47.690 142.025 47.980 143.190 ;
        RECT 48.610 143.165 48.785 143.725 ;
        RECT 48.955 143.415 49.650 143.585 ;
        RECT 49.480 143.165 49.650 143.415 ;
        RECT 49.825 143.385 50.245 143.585 ;
        RECT 50.415 143.385 50.745 143.585 ;
        RECT 50.915 143.385 51.245 143.585 ;
        RECT 51.415 143.165 51.585 143.795 ;
        RECT 52.290 143.775 52.630 144.405 ;
        RECT 52.800 143.775 53.050 144.575 ;
        RECT 53.240 143.925 53.570 144.405 ;
        RECT 53.740 144.115 53.965 144.575 ;
        RECT 54.135 143.925 54.465 144.405 ;
        RECT 51.770 143.335 52.120 143.585 ;
        RECT 52.290 143.165 52.465 143.775 ;
        RECT 53.240 143.755 54.465 143.925 ;
        RECT 55.095 143.795 55.595 144.405 ;
        RECT 56.520 144.095 56.820 144.575 ;
        RECT 56.990 143.925 57.250 144.380 ;
        RECT 57.420 144.095 57.680 144.575 ;
        RECT 57.860 143.925 58.120 144.380 ;
        RECT 58.290 144.095 58.540 144.575 ;
        RECT 58.720 143.925 58.980 144.380 ;
        RECT 59.150 144.095 59.400 144.575 ;
        RECT 59.580 143.925 59.840 144.380 ;
        RECT 60.010 144.095 60.255 144.575 ;
        RECT 60.425 143.925 60.700 144.380 ;
        RECT 60.870 144.095 61.115 144.575 ;
        RECT 61.285 143.925 61.545 144.380 ;
        RECT 61.715 144.095 61.975 144.575 ;
        RECT 62.145 143.925 62.405 144.380 ;
        RECT 62.575 144.095 62.835 144.575 ;
        RECT 63.005 143.925 63.265 144.380 ;
        RECT 63.435 144.015 63.695 144.575 ;
        RECT 52.635 143.415 53.330 143.585 ;
        RECT 53.160 143.165 53.330 143.415 ;
        RECT 53.505 143.385 53.925 143.585 ;
        RECT 54.095 143.385 54.425 143.585 ;
        RECT 54.595 143.385 54.925 143.585 ;
        RECT 55.095 143.165 55.265 143.795 ;
        RECT 56.520 143.755 63.265 143.925 ;
        RECT 55.450 143.335 55.800 143.585 ;
        RECT 56.520 143.555 57.685 143.755 ;
        RECT 63.865 143.585 64.115 144.395 ;
        RECT 64.295 144.050 64.555 144.575 ;
        RECT 64.725 143.585 64.975 144.395 ;
        RECT 65.155 144.065 65.460 144.575 ;
        RECT 56.490 143.385 57.685 143.555 ;
        RECT 56.520 143.165 57.685 143.385 ;
        RECT 57.855 143.335 64.975 143.585 ;
        RECT 65.145 143.335 65.460 143.895 ;
        RECT 65.630 143.825 66.840 144.575 ;
        RECT 67.070 144.095 67.350 144.575 ;
        RECT 67.520 143.925 67.780 144.315 ;
        RECT 67.955 144.095 68.210 144.575 ;
        RECT 68.380 143.925 68.675 144.315 ;
        RECT 68.855 144.095 69.130 144.575 ;
        RECT 69.300 144.075 69.600 144.405 ;
        RECT 48.610 142.195 48.950 143.165 ;
        RECT 49.120 142.025 49.290 143.165 ;
        RECT 49.480 142.995 51.915 143.165 ;
        RECT 49.560 142.025 49.810 142.825 ;
        RECT 50.455 142.195 50.785 142.995 ;
        RECT 51.085 142.025 51.415 142.825 ;
        RECT 51.585 142.195 51.915 142.995 ;
        RECT 52.290 142.195 52.630 143.165 ;
        RECT 52.800 142.025 52.970 143.165 ;
        RECT 53.160 142.995 55.595 143.165 ;
        RECT 53.240 142.025 53.490 142.825 ;
        RECT 54.135 142.195 54.465 142.995 ;
        RECT 54.765 142.025 55.095 142.825 ;
        RECT 55.265 142.195 55.595 142.995 ;
        RECT 56.520 142.940 63.265 143.165 ;
        RECT 56.520 142.025 56.790 142.770 ;
        RECT 56.960 142.200 57.250 142.940 ;
        RECT 57.860 142.925 63.265 142.940 ;
        RECT 57.420 142.030 57.675 142.755 ;
        RECT 57.860 142.200 58.120 142.925 ;
        RECT 58.290 142.030 58.535 142.755 ;
        RECT 58.720 142.200 58.980 142.925 ;
        RECT 59.150 142.030 59.395 142.755 ;
        RECT 59.580 142.200 59.840 142.925 ;
        RECT 60.010 142.030 60.255 142.755 ;
        RECT 60.425 142.200 60.685 142.925 ;
        RECT 60.855 142.030 61.115 142.755 ;
        RECT 61.285 142.200 61.545 142.925 ;
        RECT 61.715 142.030 61.975 142.755 ;
        RECT 62.145 142.200 62.405 142.925 ;
        RECT 62.575 142.030 62.835 142.755 ;
        RECT 63.005 142.200 63.265 142.925 ;
        RECT 63.435 142.030 63.695 142.825 ;
        RECT 63.865 142.200 64.115 143.335 ;
        RECT 57.420 142.025 63.695 142.030 ;
        RECT 64.295 142.025 64.555 142.835 ;
        RECT 64.730 142.195 64.975 143.335 ;
        RECT 65.630 143.115 66.150 143.655 ;
        RECT 66.320 143.285 66.840 143.825 ;
        RECT 67.025 143.755 68.675 143.925 ;
        RECT 67.025 143.245 67.430 143.755 ;
        RECT 67.600 143.415 68.740 143.585 ;
        RECT 65.155 142.025 65.450 142.835 ;
        RECT 65.630 142.025 66.840 143.115 ;
        RECT 67.025 143.075 67.780 143.245 ;
        RECT 67.065 142.025 67.350 142.895 ;
        RECT 67.520 142.825 67.780 143.075 ;
        RECT 68.570 143.165 68.740 143.415 ;
        RECT 68.910 143.335 69.260 143.905 ;
        RECT 69.430 143.165 69.600 144.075 ;
        RECT 69.780 144.045 70.110 144.405 ;
        RECT 70.280 144.215 70.610 144.575 ;
        RECT 70.810 144.045 71.140 144.405 ;
        RECT 69.780 143.835 71.140 144.045 ;
        RECT 71.650 143.815 72.360 144.405 ;
        RECT 73.450 143.850 73.740 144.575 ;
        RECT 73.910 144.075 74.210 144.405 ;
        RECT 74.380 144.095 74.655 144.575 ;
        RECT 72.130 143.725 72.360 143.815 ;
        RECT 69.770 143.335 70.080 143.665 ;
        RECT 70.290 143.335 70.665 143.665 ;
        RECT 70.985 143.335 71.480 143.665 ;
        RECT 68.570 142.995 69.600 143.165 ;
        RECT 67.520 142.655 68.640 142.825 ;
        RECT 67.520 142.195 67.780 142.655 ;
        RECT 67.955 142.025 68.210 142.485 ;
        RECT 68.380 142.195 68.640 142.655 ;
        RECT 68.810 142.025 69.120 142.825 ;
        RECT 69.290 142.195 69.600 142.995 ;
        RECT 69.780 142.025 70.110 143.085 ;
        RECT 70.290 142.410 70.460 143.335 ;
        RECT 70.630 142.845 70.960 143.065 ;
        RECT 71.155 143.045 71.480 143.335 ;
        RECT 71.655 143.045 71.985 143.585 ;
        RECT 72.155 142.845 72.360 143.725 ;
        RECT 70.630 142.615 72.360 142.845 ;
        RECT 70.630 142.215 70.960 142.615 ;
        RECT 71.130 142.025 71.460 142.385 ;
        RECT 71.660 142.195 72.360 142.615 ;
        RECT 73.450 142.025 73.740 143.190 ;
        RECT 73.910 143.165 74.080 144.075 ;
        RECT 74.835 143.925 75.130 144.315 ;
        RECT 75.300 144.095 75.555 144.575 ;
        RECT 75.730 143.925 75.990 144.315 ;
        RECT 76.160 144.095 76.440 144.575 ;
        RECT 74.250 143.335 74.600 143.905 ;
        RECT 74.835 143.755 76.485 143.925 ;
        RECT 76.670 143.805 79.260 144.575 ;
        RECT 74.770 143.415 75.910 143.585 ;
        RECT 74.770 143.165 74.940 143.415 ;
        RECT 76.080 143.245 76.485 143.755 ;
        RECT 73.910 142.995 74.940 143.165 ;
        RECT 75.730 143.075 76.485 143.245 ;
        RECT 76.670 143.115 77.880 143.635 ;
        RECT 78.050 143.285 79.260 143.805 ;
        RECT 79.705 143.765 79.950 144.370 ;
        RECT 80.170 144.040 80.680 144.575 ;
        RECT 79.430 143.595 80.660 143.765 ;
        RECT 73.910 142.195 74.220 142.995 ;
        RECT 75.730 142.825 75.990 143.075 ;
        RECT 74.390 142.025 74.700 142.825 ;
        RECT 74.870 142.655 75.990 142.825 ;
        RECT 74.870 142.195 75.130 142.655 ;
        RECT 75.300 142.025 75.555 142.485 ;
        RECT 75.730 142.195 75.990 142.655 ;
        RECT 76.160 142.025 76.445 142.895 ;
        RECT 76.670 142.025 79.260 143.115 ;
        RECT 79.430 142.785 79.770 143.595 ;
        RECT 79.940 143.030 80.690 143.220 ;
        RECT 79.430 142.375 79.945 142.785 ;
        RECT 80.180 142.025 80.350 142.785 ;
        RECT 80.520 142.365 80.690 143.030 ;
        RECT 80.860 143.045 81.050 144.405 ;
        RECT 81.220 143.555 81.495 144.405 ;
        RECT 81.685 144.040 82.215 144.405 ;
        RECT 82.640 144.175 82.970 144.575 ;
        RECT 82.040 144.005 82.215 144.040 ;
        RECT 81.220 143.385 81.500 143.555 ;
        RECT 81.220 143.245 81.495 143.385 ;
        RECT 81.700 143.045 81.870 143.845 ;
        RECT 80.860 142.875 81.870 143.045 ;
        RECT 82.040 143.835 82.970 144.005 ;
        RECT 83.140 143.835 83.395 144.405 ;
        RECT 83.660 144.025 83.830 144.405 ;
        RECT 84.010 144.195 84.340 144.575 ;
        RECT 83.660 143.855 84.325 144.025 ;
        RECT 84.520 143.900 84.780 144.405 ;
        RECT 82.040 142.705 82.210 143.835 ;
        RECT 82.800 143.665 82.970 143.835 ;
        RECT 81.085 142.535 82.210 142.705 ;
        RECT 82.380 143.335 82.575 143.665 ;
        RECT 82.800 143.335 83.055 143.665 ;
        RECT 82.380 142.365 82.550 143.335 ;
        RECT 83.225 143.165 83.395 143.835 ;
        RECT 83.590 143.305 83.920 143.675 ;
        RECT 84.155 143.600 84.325 143.855 ;
        RECT 80.520 142.195 82.550 142.365 ;
        RECT 82.720 142.025 82.890 143.165 ;
        RECT 83.060 142.195 83.395 143.165 ;
        RECT 84.155 143.270 84.440 143.600 ;
        RECT 84.155 143.125 84.325 143.270 ;
        RECT 83.660 142.955 84.325 143.125 ;
        RECT 84.610 143.100 84.780 143.900 ;
        RECT 85.410 143.805 88.000 144.575 ;
        RECT 88.180 144.075 88.510 144.575 ;
        RECT 88.710 144.005 88.880 144.355 ;
        RECT 89.080 144.175 89.410 144.575 ;
        RECT 89.580 144.005 89.750 144.355 ;
        RECT 89.920 144.175 90.300 144.575 ;
        RECT 83.660 142.195 83.830 142.955 ;
        RECT 84.010 142.025 84.340 142.785 ;
        RECT 84.510 142.195 84.780 143.100 ;
        RECT 85.410 143.115 86.620 143.635 ;
        RECT 86.790 143.285 88.000 143.805 ;
        RECT 88.175 143.335 88.525 143.905 ;
        RECT 88.710 143.835 90.320 144.005 ;
        RECT 90.490 143.900 90.760 144.245 ;
        RECT 90.150 143.665 90.320 143.835 ;
        RECT 85.410 142.025 88.000 143.115 ;
        RECT 88.175 142.875 88.495 143.165 ;
        RECT 88.695 143.045 89.405 143.665 ;
        RECT 89.575 143.335 89.980 143.665 ;
        RECT 90.150 143.335 90.420 143.665 ;
        RECT 90.150 143.165 90.320 143.335 ;
        RECT 90.590 143.165 90.760 143.900 ;
        RECT 89.595 142.995 90.320 143.165 ;
        RECT 89.595 142.875 89.765 142.995 ;
        RECT 88.175 142.705 89.765 142.875 ;
        RECT 88.175 142.245 89.830 142.535 ;
        RECT 90.000 142.025 90.280 142.825 ;
        RECT 90.490 142.195 90.760 143.165 ;
        RECT 90.930 143.775 91.270 144.405 ;
        RECT 91.440 143.775 91.690 144.575 ;
        RECT 91.880 143.925 92.210 144.405 ;
        RECT 92.380 144.115 92.605 144.575 ;
        RECT 92.775 143.925 93.105 144.405 ;
        RECT 90.930 143.725 91.160 143.775 ;
        RECT 91.880 143.755 93.105 143.925 ;
        RECT 93.735 143.795 94.235 144.405 ;
        RECT 95.735 143.795 96.235 144.405 ;
        RECT 90.930 143.165 91.105 143.725 ;
        RECT 91.275 143.415 91.970 143.585 ;
        RECT 91.800 143.165 91.970 143.415 ;
        RECT 92.145 143.385 92.565 143.585 ;
        RECT 92.735 143.385 93.065 143.585 ;
        RECT 93.235 143.385 93.565 143.585 ;
        RECT 93.735 143.165 93.905 143.795 ;
        RECT 94.090 143.335 94.440 143.585 ;
        RECT 95.530 143.335 95.880 143.585 ;
        RECT 96.065 143.165 96.235 143.795 ;
        RECT 96.865 143.925 97.195 144.405 ;
        RECT 97.365 144.115 97.590 144.575 ;
        RECT 97.760 143.925 98.090 144.405 ;
        RECT 96.865 143.755 98.090 143.925 ;
        RECT 98.280 143.775 98.530 144.575 ;
        RECT 98.700 143.775 99.040 144.405 ;
        RECT 99.210 143.850 99.500 144.575 ;
        RECT 99.680 144.075 100.010 144.575 ;
        RECT 100.210 144.005 100.380 144.355 ;
        RECT 100.580 144.175 100.910 144.575 ;
        RECT 101.080 144.005 101.250 144.355 ;
        RECT 101.420 144.175 101.800 144.575 ;
        RECT 96.405 143.385 96.735 143.585 ;
        RECT 96.905 143.385 97.235 143.585 ;
        RECT 97.405 143.385 97.825 143.585 ;
        RECT 98.000 143.415 98.695 143.585 ;
        RECT 98.000 143.165 98.170 143.415 ;
        RECT 98.865 143.165 99.040 143.775 ;
        RECT 99.675 143.335 100.025 143.905 ;
        RECT 100.210 143.835 101.820 144.005 ;
        RECT 101.990 143.900 102.260 144.245 ;
        RECT 101.650 143.665 101.820 143.835 ;
        RECT 90.930 142.195 91.270 143.165 ;
        RECT 91.440 142.025 91.610 143.165 ;
        RECT 91.800 142.995 94.235 143.165 ;
        RECT 91.880 142.025 92.130 142.825 ;
        RECT 92.775 142.195 93.105 142.995 ;
        RECT 93.405 142.025 93.735 142.825 ;
        RECT 93.905 142.195 94.235 142.995 ;
        RECT 95.735 142.995 98.170 143.165 ;
        RECT 95.735 142.195 96.065 142.995 ;
        RECT 96.235 142.025 96.565 142.825 ;
        RECT 96.865 142.195 97.195 142.995 ;
        RECT 97.840 142.025 98.090 142.825 ;
        RECT 98.360 142.025 98.530 143.165 ;
        RECT 98.700 142.195 99.040 143.165 ;
        RECT 99.210 142.025 99.500 143.190 ;
        RECT 99.675 142.875 99.995 143.165 ;
        RECT 100.195 143.045 100.905 143.665 ;
        RECT 101.075 143.335 101.480 143.665 ;
        RECT 101.650 143.335 101.920 143.665 ;
        RECT 101.650 143.165 101.820 143.335 ;
        RECT 102.090 143.165 102.260 143.900 ;
        RECT 102.705 143.765 102.950 144.370 ;
        RECT 103.170 144.040 103.680 144.575 ;
        RECT 101.095 142.995 101.820 143.165 ;
        RECT 101.095 142.875 101.265 142.995 ;
        RECT 99.675 142.705 101.265 142.875 ;
        RECT 99.675 142.245 101.330 142.535 ;
        RECT 101.500 142.025 101.780 142.825 ;
        RECT 101.990 142.195 102.260 143.165 ;
        RECT 102.430 143.595 103.660 143.765 ;
        RECT 102.430 142.785 102.770 143.595 ;
        RECT 102.940 143.030 103.690 143.220 ;
        RECT 102.430 142.375 102.945 142.785 ;
        RECT 103.180 142.025 103.350 142.785 ;
        RECT 103.520 142.365 103.690 143.030 ;
        RECT 103.860 143.045 104.050 144.405 ;
        RECT 104.220 144.235 104.495 144.405 ;
        RECT 104.220 144.065 104.500 144.235 ;
        RECT 104.220 143.245 104.495 144.065 ;
        RECT 104.685 144.040 105.215 144.405 ;
        RECT 105.640 144.175 105.970 144.575 ;
        RECT 105.040 144.005 105.215 144.040 ;
        RECT 104.700 143.045 104.870 143.845 ;
        RECT 103.860 142.875 104.870 143.045 ;
        RECT 105.040 143.835 105.970 144.005 ;
        RECT 106.140 143.835 106.395 144.405 ;
        RECT 105.040 142.705 105.210 143.835 ;
        RECT 105.800 143.665 105.970 143.835 ;
        RECT 104.085 142.535 105.210 142.705 ;
        RECT 105.380 143.335 105.575 143.665 ;
        RECT 105.800 143.335 106.055 143.665 ;
        RECT 105.380 142.365 105.550 143.335 ;
        RECT 106.225 143.165 106.395 143.835 ;
        RECT 107.490 143.805 111.000 144.575 ;
        RECT 111.170 143.825 112.380 144.575 ;
        RECT 103.520 142.195 105.550 142.365 ;
        RECT 105.720 142.025 105.890 143.165 ;
        RECT 106.060 142.195 106.395 143.165 ;
        RECT 107.490 143.115 109.180 143.635 ;
        RECT 109.350 143.285 111.000 143.805 ;
        RECT 111.170 143.115 111.690 143.655 ;
        RECT 111.860 143.285 112.380 143.825 ;
        RECT 107.490 142.025 111.000 143.115 ;
        RECT 111.170 142.025 112.380 143.115 ;
        RECT 18.165 141.855 112.465 142.025 ;
        RECT 18.250 140.765 19.460 141.855 ;
        RECT 18.250 140.055 18.770 140.595 ;
        RECT 18.940 140.225 19.460 140.765 ;
        RECT 19.635 140.665 19.890 141.545 ;
        RECT 20.060 140.715 20.365 141.855 ;
        RECT 20.705 141.475 21.035 141.855 ;
        RECT 21.215 141.305 21.385 141.595 ;
        RECT 21.555 141.395 21.805 141.855 ;
        RECT 20.585 141.135 21.385 141.305 ;
        RECT 21.975 141.345 22.845 141.685 ;
        RECT 18.250 139.305 19.460 140.055 ;
        RECT 19.635 140.015 19.845 140.665 ;
        RECT 20.585 140.545 20.755 141.135 ;
        RECT 21.975 140.965 22.145 141.345 ;
        RECT 23.080 141.225 23.250 141.685 ;
        RECT 23.420 141.395 23.790 141.855 ;
        RECT 24.085 141.255 24.255 141.595 ;
        RECT 24.425 141.425 24.755 141.855 ;
        RECT 24.990 141.255 25.160 141.595 ;
        RECT 20.925 140.795 22.145 140.965 ;
        RECT 22.315 140.885 22.775 141.175 ;
        RECT 23.080 141.055 23.640 141.225 ;
        RECT 24.085 141.085 25.160 141.255 ;
        RECT 25.330 141.355 26.010 141.685 ;
        RECT 26.225 141.355 26.475 141.685 ;
        RECT 26.645 141.395 26.895 141.855 ;
        RECT 23.470 140.915 23.640 141.055 ;
        RECT 22.315 140.875 23.280 140.885 ;
        RECT 21.975 140.705 22.145 140.795 ;
        RECT 22.605 140.715 23.280 140.875 ;
        RECT 20.015 140.515 20.755 140.545 ;
        RECT 20.015 140.215 20.930 140.515 ;
        RECT 20.605 140.040 20.930 140.215 ;
        RECT 19.635 139.485 19.890 140.015 ;
        RECT 20.060 139.305 20.365 139.765 ;
        RECT 20.610 139.685 20.930 140.040 ;
        RECT 21.100 140.255 21.640 140.625 ;
        RECT 21.975 140.535 22.380 140.705 ;
        RECT 21.100 139.855 21.340 140.255 ;
        RECT 21.820 140.085 22.040 140.365 ;
        RECT 21.510 139.915 22.040 140.085 ;
        RECT 21.510 139.685 21.680 139.915 ;
        RECT 22.210 139.755 22.380 140.535 ;
        RECT 22.550 139.925 22.900 140.545 ;
        RECT 23.070 139.925 23.280 140.715 ;
        RECT 23.470 140.745 24.970 140.915 ;
        RECT 23.470 140.055 23.640 140.745 ;
        RECT 25.330 140.575 25.500 141.355 ;
        RECT 26.305 141.225 26.475 141.355 ;
        RECT 23.810 140.405 25.500 140.575 ;
        RECT 25.670 140.795 26.135 141.185 ;
        RECT 26.305 141.055 26.700 141.225 ;
        RECT 23.810 140.225 23.980 140.405 ;
        RECT 20.610 139.515 21.680 139.685 ;
        RECT 21.850 139.305 22.040 139.745 ;
        RECT 22.210 139.475 23.160 139.755 ;
        RECT 23.470 139.665 23.730 140.055 ;
        RECT 24.150 139.985 24.940 140.235 ;
        RECT 23.380 139.495 23.730 139.665 ;
        RECT 23.940 139.305 24.270 139.765 ;
        RECT 25.145 139.695 25.315 140.405 ;
        RECT 25.670 140.205 25.840 140.795 ;
        RECT 25.485 139.985 25.840 140.205 ;
        RECT 26.010 139.985 26.360 140.605 ;
        RECT 26.530 139.695 26.700 141.055 ;
        RECT 27.065 140.885 27.390 141.670 ;
        RECT 26.870 139.835 27.330 140.885 ;
        RECT 25.145 139.525 26.000 139.695 ;
        RECT 26.205 139.525 26.700 139.695 ;
        RECT 26.870 139.305 27.200 139.665 ;
        RECT 27.560 139.565 27.730 141.685 ;
        RECT 27.900 141.355 28.230 141.855 ;
        RECT 28.400 141.185 28.655 141.685 ;
        RECT 27.905 141.015 28.655 141.185 ;
        RECT 28.945 141.225 29.230 141.685 ;
        RECT 29.400 141.395 29.670 141.855 ;
        RECT 27.905 140.025 28.135 141.015 ;
        RECT 28.945 141.005 29.900 141.225 ;
        RECT 28.305 140.195 28.655 140.845 ;
        RECT 28.830 140.275 29.520 140.835 ;
        RECT 29.690 140.105 29.900 141.005 ;
        RECT 27.905 139.855 28.655 140.025 ;
        RECT 27.900 139.305 28.230 139.685 ;
        RECT 28.400 139.565 28.655 139.855 ;
        RECT 28.945 139.935 29.900 140.105 ;
        RECT 30.070 140.835 30.470 141.685 ;
        RECT 30.660 141.225 30.940 141.685 ;
        RECT 31.460 141.395 31.785 141.855 ;
        RECT 30.660 141.005 31.785 141.225 ;
        RECT 30.070 140.275 31.165 140.835 ;
        RECT 31.335 140.545 31.785 141.005 ;
        RECT 31.955 140.715 32.340 141.685 ;
        RECT 28.945 139.475 29.230 139.935 ;
        RECT 29.400 139.305 29.670 139.765 ;
        RECT 30.070 139.475 30.470 140.275 ;
        RECT 31.335 140.215 31.890 140.545 ;
        RECT 31.335 140.105 31.785 140.215 ;
        RECT 30.660 139.935 31.785 140.105 ;
        RECT 32.060 140.045 32.340 140.715 ;
        RECT 30.660 139.475 30.940 139.935 ;
        RECT 31.460 139.305 31.785 139.765 ;
        RECT 31.955 139.475 32.340 140.045 ;
        RECT 33.430 140.780 33.700 141.685 ;
        RECT 33.870 141.095 34.200 141.855 ;
        RECT 34.380 140.925 34.550 141.685 ;
        RECT 33.430 139.980 33.600 140.780 ;
        RECT 33.885 140.755 34.550 140.925 ;
        RECT 33.885 140.610 34.055 140.755 ;
        RECT 34.810 140.690 35.100 141.855 ;
        RECT 36.280 140.925 36.450 141.685 ;
        RECT 36.630 141.095 36.960 141.855 ;
        RECT 36.280 140.755 36.945 140.925 ;
        RECT 37.130 140.780 37.400 141.685 ;
        RECT 33.770 140.280 34.055 140.610 ;
        RECT 36.775 140.610 36.945 140.755 ;
        RECT 33.885 140.025 34.055 140.280 ;
        RECT 34.290 140.205 34.620 140.575 ;
        RECT 36.210 140.205 36.540 140.575 ;
        RECT 36.775 140.280 37.060 140.610 ;
        RECT 33.430 139.475 33.690 139.980 ;
        RECT 33.885 139.855 34.550 140.025 ;
        RECT 33.870 139.305 34.200 139.685 ;
        RECT 34.380 139.475 34.550 139.855 ;
        RECT 34.810 139.305 35.100 140.030 ;
        RECT 36.775 140.025 36.945 140.280 ;
        RECT 36.280 139.855 36.945 140.025 ;
        RECT 37.230 139.980 37.400 140.780 ;
        RECT 37.720 140.705 38.050 141.855 ;
        RECT 38.220 140.835 38.390 141.685 ;
        RECT 38.560 141.055 38.890 141.855 ;
        RECT 39.060 140.835 39.230 141.685 ;
        RECT 39.410 141.055 39.650 141.855 ;
        RECT 39.820 140.875 40.150 141.685 ;
        RECT 40.335 141.345 41.990 141.635 ;
        RECT 38.220 140.665 39.230 140.835 ;
        RECT 39.435 140.705 40.150 140.875 ;
        RECT 40.335 141.005 41.925 141.175 ;
        RECT 42.160 141.055 42.440 141.855 ;
        RECT 40.335 140.715 40.655 141.005 ;
        RECT 41.755 140.885 41.925 141.005 ;
        RECT 38.220 140.125 38.715 140.665 ;
        RECT 39.435 140.465 39.605 140.705 ;
        RECT 39.105 140.295 39.605 140.465 ;
        RECT 39.775 140.295 40.155 140.535 ;
        RECT 39.435 140.125 39.605 140.295 ;
        RECT 36.280 139.475 36.450 139.855 ;
        RECT 36.630 139.305 36.960 139.685 ;
        RECT 37.140 139.475 37.400 139.980 ;
        RECT 37.720 139.305 38.050 140.105 ;
        RECT 38.220 139.955 39.230 140.125 ;
        RECT 39.435 139.955 40.070 140.125 ;
        RECT 40.335 139.975 40.685 140.545 ;
        RECT 40.855 140.215 41.565 140.835 ;
        RECT 41.755 140.715 42.480 140.885 ;
        RECT 42.650 140.715 42.920 141.685 ;
        RECT 42.310 140.545 42.480 140.715 ;
        RECT 41.735 140.215 42.140 140.545 ;
        RECT 42.310 140.215 42.580 140.545 ;
        RECT 42.310 140.045 42.480 140.215 ;
        RECT 38.220 139.475 38.390 139.955 ;
        RECT 38.560 139.305 38.890 139.785 ;
        RECT 39.060 139.475 39.230 139.955 ;
        RECT 39.480 139.305 39.720 139.785 ;
        RECT 39.900 139.475 40.070 139.955 ;
        RECT 40.870 139.875 42.480 140.045 ;
        RECT 42.750 139.980 42.920 140.715 ;
        RECT 40.340 139.305 40.670 139.805 ;
        RECT 40.870 139.525 41.040 139.875 ;
        RECT 41.240 139.305 41.570 139.705 ;
        RECT 41.740 139.525 41.910 139.875 ;
        RECT 42.080 139.305 42.460 139.705 ;
        RECT 42.650 139.635 42.920 139.980 ;
        RECT 43.090 140.715 43.430 141.685 ;
        RECT 43.600 140.715 43.770 141.855 ;
        RECT 44.040 141.055 44.290 141.855 ;
        RECT 44.935 140.885 45.265 141.685 ;
        RECT 45.565 141.055 45.895 141.855 ;
        RECT 46.065 140.885 46.395 141.685 ;
        RECT 43.960 140.715 46.395 140.885 ;
        RECT 47.270 140.715 47.500 141.855 ;
        RECT 43.090 140.105 43.265 140.715 ;
        RECT 43.960 140.465 44.130 140.715 ;
        RECT 43.435 140.295 44.130 140.465 ;
        RECT 44.305 140.295 44.725 140.495 ;
        RECT 44.895 140.295 45.225 140.495 ;
        RECT 45.395 140.295 45.725 140.495 ;
        RECT 43.090 139.475 43.430 140.105 ;
        RECT 43.600 139.305 43.850 140.105 ;
        RECT 44.040 139.955 45.265 140.125 ;
        RECT 44.040 139.475 44.370 139.955 ;
        RECT 44.540 139.305 44.765 139.765 ;
        RECT 44.935 139.475 45.265 139.955 ;
        RECT 45.895 140.085 46.065 140.715 ;
        RECT 47.670 140.705 48.000 141.685 ;
        RECT 48.170 140.715 48.380 141.855 ;
        RECT 48.615 141.345 50.270 141.635 ;
        RECT 48.615 141.005 50.205 141.175 ;
        RECT 50.440 141.055 50.720 141.855 ;
        RECT 48.615 140.715 48.935 141.005 ;
        RECT 50.035 140.885 50.205 141.005 ;
        RECT 46.250 140.295 46.600 140.545 ;
        RECT 47.250 140.295 47.580 140.545 ;
        RECT 45.895 139.475 46.395 140.085 ;
        RECT 47.270 139.305 47.500 140.125 ;
        RECT 47.750 140.105 48.000 140.705 ;
        RECT 49.130 140.665 49.845 140.835 ;
        RECT 50.035 140.715 50.760 140.885 ;
        RECT 50.930 140.715 51.200 141.685 ;
        RECT 47.670 139.475 48.000 140.105 ;
        RECT 48.170 139.305 48.380 140.125 ;
        RECT 48.615 139.975 48.965 140.545 ;
        RECT 49.135 140.215 49.845 140.665 ;
        RECT 50.590 140.545 50.760 140.715 ;
        RECT 50.015 140.215 50.420 140.545 ;
        RECT 50.590 140.215 50.860 140.545 ;
        RECT 50.590 140.045 50.760 140.215 ;
        RECT 49.150 139.875 50.760 140.045 ;
        RECT 51.030 139.980 51.200 140.715 ;
        RECT 48.620 139.305 48.950 139.805 ;
        RECT 49.150 139.525 49.320 139.875 ;
        RECT 49.520 139.305 49.850 139.705 ;
        RECT 50.020 139.525 50.190 139.875 ;
        RECT 50.360 139.305 50.740 139.705 ;
        RECT 50.930 139.635 51.200 139.980 ;
        RECT 51.375 140.665 51.630 141.545 ;
        RECT 51.800 140.715 52.105 141.855 ;
        RECT 52.445 141.475 52.775 141.855 ;
        RECT 52.955 141.305 53.125 141.595 ;
        RECT 53.295 141.395 53.545 141.855 ;
        RECT 52.325 141.135 53.125 141.305 ;
        RECT 53.715 141.345 54.585 141.685 ;
        RECT 51.375 140.015 51.585 140.665 ;
        RECT 52.325 140.545 52.495 141.135 ;
        RECT 53.715 140.965 53.885 141.345 ;
        RECT 54.820 141.225 54.990 141.685 ;
        RECT 55.160 141.395 55.530 141.855 ;
        RECT 55.825 141.255 55.995 141.595 ;
        RECT 56.165 141.425 56.495 141.855 ;
        RECT 56.730 141.255 56.900 141.595 ;
        RECT 52.665 140.795 53.885 140.965 ;
        RECT 54.055 140.885 54.515 141.175 ;
        RECT 54.820 141.055 55.380 141.225 ;
        RECT 55.825 141.085 56.900 141.255 ;
        RECT 57.070 141.355 57.750 141.685 ;
        RECT 57.965 141.355 58.215 141.685 ;
        RECT 58.385 141.395 58.635 141.855 ;
        RECT 55.210 140.915 55.380 141.055 ;
        RECT 54.055 140.875 55.020 140.885 ;
        RECT 53.715 140.705 53.885 140.795 ;
        RECT 54.345 140.715 55.020 140.875 ;
        RECT 51.755 140.515 52.495 140.545 ;
        RECT 51.755 140.215 52.670 140.515 ;
        RECT 52.345 140.040 52.670 140.215 ;
        RECT 51.375 139.485 51.630 140.015 ;
        RECT 51.800 139.305 52.105 139.765 ;
        RECT 52.350 139.685 52.670 140.040 ;
        RECT 52.840 140.255 53.380 140.625 ;
        RECT 53.715 140.535 54.120 140.705 ;
        RECT 52.840 139.855 53.080 140.255 ;
        RECT 53.560 140.085 53.780 140.365 ;
        RECT 53.250 139.915 53.780 140.085 ;
        RECT 53.250 139.685 53.420 139.915 ;
        RECT 53.950 139.755 54.120 140.535 ;
        RECT 54.290 139.925 54.640 140.545 ;
        RECT 54.810 139.925 55.020 140.715 ;
        RECT 55.210 140.745 56.710 140.915 ;
        RECT 55.210 140.055 55.380 140.745 ;
        RECT 57.070 140.575 57.240 141.355 ;
        RECT 58.045 141.225 58.215 141.355 ;
        RECT 55.550 140.405 57.240 140.575 ;
        RECT 57.410 140.795 57.875 141.185 ;
        RECT 58.045 141.055 58.440 141.225 ;
        RECT 55.550 140.225 55.720 140.405 ;
        RECT 52.350 139.515 53.420 139.685 ;
        RECT 53.590 139.305 53.780 139.745 ;
        RECT 53.950 139.475 54.900 139.755 ;
        RECT 55.210 139.665 55.470 140.055 ;
        RECT 55.890 139.985 56.680 140.235 ;
        RECT 55.120 139.495 55.470 139.665 ;
        RECT 55.680 139.305 56.010 139.765 ;
        RECT 56.885 139.695 57.055 140.405 ;
        RECT 57.410 140.205 57.580 140.795 ;
        RECT 57.225 139.985 57.580 140.205 ;
        RECT 57.750 139.985 58.100 140.605 ;
        RECT 58.270 139.695 58.440 141.055 ;
        RECT 58.805 140.885 59.130 141.670 ;
        RECT 58.610 139.835 59.070 140.885 ;
        RECT 56.885 139.525 57.740 139.695 ;
        RECT 57.945 139.525 58.440 139.695 ;
        RECT 58.610 139.305 58.940 139.665 ;
        RECT 59.300 139.565 59.470 141.685 ;
        RECT 59.640 141.355 59.970 141.855 ;
        RECT 60.140 141.185 60.395 141.685 ;
        RECT 59.645 141.015 60.395 141.185 ;
        RECT 59.645 140.025 59.875 141.015 ;
        RECT 60.045 140.195 60.395 140.845 ;
        RECT 60.570 140.690 60.860 141.855 ;
        RECT 61.495 140.705 61.755 141.855 ;
        RECT 61.930 140.780 62.185 141.685 ;
        RECT 62.355 141.095 62.685 141.855 ;
        RECT 62.900 140.925 63.070 141.685 ;
        RECT 59.645 139.855 60.395 140.025 ;
        RECT 59.640 139.305 59.970 139.685 ;
        RECT 60.140 139.565 60.395 139.855 ;
        RECT 60.570 139.305 60.860 140.030 ;
        RECT 61.495 139.305 61.755 140.145 ;
        RECT 61.930 140.050 62.100 140.780 ;
        RECT 62.355 140.755 63.070 140.925 ;
        RECT 62.355 140.545 62.525 140.755 ;
        RECT 63.335 140.705 63.595 141.855 ;
        RECT 63.770 140.780 64.025 141.685 ;
        RECT 64.195 141.095 64.525 141.855 ;
        RECT 64.740 140.925 64.910 141.685 ;
        RECT 62.270 140.215 62.525 140.545 ;
        RECT 61.930 139.475 62.185 140.050 ;
        RECT 62.355 140.025 62.525 140.215 ;
        RECT 62.805 140.205 63.160 140.575 ;
        RECT 62.355 139.855 63.070 140.025 ;
        RECT 62.355 139.305 62.685 139.685 ;
        RECT 62.900 139.475 63.070 139.855 ;
        RECT 63.335 139.305 63.595 140.145 ;
        RECT 63.770 140.050 63.940 140.780 ;
        RECT 64.195 140.755 64.910 140.925 ;
        RECT 65.260 140.925 65.430 141.685 ;
        RECT 65.645 141.095 65.975 141.855 ;
        RECT 65.260 140.755 65.975 140.925 ;
        RECT 66.145 140.780 66.400 141.685 ;
        RECT 64.195 140.545 64.365 140.755 ;
        RECT 64.110 140.215 64.365 140.545 ;
        RECT 63.770 139.475 64.025 140.050 ;
        RECT 64.195 140.025 64.365 140.215 ;
        RECT 64.645 140.205 65.000 140.575 ;
        RECT 65.170 140.205 65.525 140.575 ;
        RECT 65.805 140.545 65.975 140.755 ;
        RECT 65.805 140.215 66.060 140.545 ;
        RECT 65.805 140.025 65.975 140.215 ;
        RECT 66.230 140.050 66.400 140.780 ;
        RECT 66.575 140.705 66.835 141.855 ;
        RECT 67.100 140.925 67.270 141.685 ;
        RECT 67.485 141.095 67.815 141.855 ;
        RECT 67.100 140.755 67.815 140.925 ;
        RECT 67.985 140.780 68.240 141.685 ;
        RECT 67.010 140.205 67.365 140.575 ;
        RECT 67.645 140.545 67.815 140.755 ;
        RECT 67.645 140.215 67.900 140.545 ;
        RECT 64.195 139.855 64.910 140.025 ;
        RECT 64.195 139.305 64.525 139.685 ;
        RECT 64.740 139.475 64.910 139.855 ;
        RECT 65.260 139.855 65.975 140.025 ;
        RECT 65.260 139.475 65.430 139.855 ;
        RECT 65.645 139.305 65.975 139.685 ;
        RECT 66.145 139.475 66.400 140.050 ;
        RECT 66.575 139.305 66.835 140.145 ;
        RECT 67.645 140.025 67.815 140.215 ;
        RECT 68.070 140.050 68.240 140.780 ;
        RECT 68.415 140.705 68.675 141.855 ;
        RECT 68.850 140.715 69.190 141.685 ;
        RECT 69.360 140.715 69.530 141.855 ;
        RECT 69.800 141.055 70.050 141.855 ;
        RECT 70.695 140.885 71.025 141.685 ;
        RECT 71.325 141.055 71.655 141.855 ;
        RECT 71.825 140.885 72.155 141.685 ;
        RECT 69.720 140.715 72.155 140.885 ;
        RECT 72.530 140.715 72.870 141.685 ;
        RECT 73.040 140.715 73.210 141.855 ;
        RECT 73.480 141.055 73.730 141.855 ;
        RECT 74.375 140.885 74.705 141.685 ;
        RECT 75.005 141.055 75.335 141.855 ;
        RECT 75.505 140.885 75.835 141.685 ;
        RECT 73.400 140.715 75.835 140.885 ;
        RECT 77.045 140.875 77.300 141.545 ;
        RECT 77.480 141.055 77.765 141.855 ;
        RECT 77.945 141.135 78.275 141.645 ;
        RECT 68.850 140.665 69.080 140.715 ;
        RECT 67.100 139.855 67.815 140.025 ;
        RECT 67.100 139.475 67.270 139.855 ;
        RECT 67.485 139.305 67.815 139.685 ;
        RECT 67.985 139.475 68.240 140.050 ;
        RECT 68.415 139.305 68.675 140.145 ;
        RECT 68.850 140.105 69.025 140.665 ;
        RECT 69.720 140.465 69.890 140.715 ;
        RECT 69.195 140.295 69.890 140.465 ;
        RECT 70.065 140.295 70.485 140.495 ;
        RECT 70.655 140.295 70.985 140.495 ;
        RECT 71.155 140.295 71.485 140.495 ;
        RECT 68.850 139.475 69.190 140.105 ;
        RECT 69.360 139.305 69.610 140.105 ;
        RECT 69.800 139.955 71.025 140.125 ;
        RECT 69.800 139.475 70.130 139.955 ;
        RECT 70.300 139.305 70.525 139.765 ;
        RECT 70.695 139.475 71.025 139.955 ;
        RECT 71.655 140.085 71.825 140.715 ;
        RECT 72.010 140.295 72.360 140.545 ;
        RECT 72.530 140.105 72.705 140.715 ;
        RECT 73.400 140.465 73.570 140.715 ;
        RECT 72.875 140.295 73.570 140.465 ;
        RECT 73.745 140.295 74.165 140.495 ;
        RECT 74.335 140.295 74.665 140.495 ;
        RECT 74.835 140.295 75.165 140.495 ;
        RECT 71.655 139.475 72.155 140.085 ;
        RECT 72.530 139.475 72.870 140.105 ;
        RECT 73.040 139.305 73.290 140.105 ;
        RECT 73.480 139.955 74.705 140.125 ;
        RECT 73.480 139.475 73.810 139.955 ;
        RECT 73.980 139.305 74.205 139.765 ;
        RECT 74.375 139.475 74.705 139.955 ;
        RECT 75.335 140.085 75.505 140.715 ;
        RECT 75.690 140.295 76.040 140.545 ;
        RECT 75.335 139.475 75.835 140.085 ;
        RECT 77.045 140.015 77.225 140.875 ;
        RECT 77.945 140.545 78.195 141.135 ;
        RECT 78.545 140.985 78.715 141.595 ;
        RECT 78.885 141.165 79.215 141.855 ;
        RECT 79.445 141.305 79.685 141.595 ;
        RECT 79.885 141.475 80.305 141.855 ;
        RECT 80.485 141.385 81.115 141.635 ;
        RECT 81.585 141.475 81.915 141.855 ;
        RECT 80.485 141.305 80.655 141.385 ;
        RECT 82.085 141.305 82.255 141.595 ;
        RECT 82.435 141.475 82.815 141.855 ;
        RECT 83.055 141.470 83.885 141.640 ;
        RECT 79.445 141.135 80.655 141.305 ;
        RECT 77.395 140.215 78.195 140.545 ;
        RECT 77.045 139.815 77.300 140.015 ;
        RECT 76.960 139.645 77.300 139.815 ;
        RECT 77.045 139.485 77.300 139.645 ;
        RECT 77.480 139.305 77.765 139.765 ;
        RECT 77.945 139.565 78.195 140.215 ;
        RECT 78.395 140.965 78.715 140.985 ;
        RECT 78.395 140.795 80.315 140.965 ;
        RECT 78.395 139.900 78.585 140.795 ;
        RECT 80.485 140.625 80.655 141.135 ;
        RECT 80.825 140.875 81.345 141.185 ;
        RECT 78.755 140.455 80.655 140.625 ;
        RECT 78.755 140.395 79.085 140.455 ;
        RECT 79.235 140.225 79.565 140.285 ;
        RECT 78.905 139.955 79.565 140.225 ;
        RECT 78.395 139.570 78.715 139.900 ;
        RECT 78.895 139.305 79.555 139.785 ;
        RECT 79.755 139.695 79.925 140.455 ;
        RECT 80.825 140.285 81.005 140.695 ;
        RECT 80.095 140.115 80.425 140.235 ;
        RECT 81.175 140.115 81.345 140.875 ;
        RECT 80.095 139.945 81.345 140.115 ;
        RECT 81.515 141.055 82.885 141.305 ;
        RECT 81.515 140.285 81.705 141.055 ;
        RECT 82.635 140.795 82.885 141.055 ;
        RECT 81.875 140.625 82.125 140.785 ;
        RECT 83.055 140.625 83.225 141.470 ;
        RECT 84.120 141.185 84.290 141.685 ;
        RECT 84.460 141.355 84.790 141.855 ;
        RECT 83.395 140.795 83.895 141.175 ;
        RECT 84.120 141.015 84.815 141.185 ;
        RECT 81.875 140.455 83.225 140.625 ;
        RECT 82.805 140.415 83.225 140.455 ;
        RECT 81.515 139.945 81.935 140.285 ;
        RECT 82.225 139.955 82.635 140.285 ;
        RECT 79.755 139.525 80.605 139.695 ;
        RECT 81.165 139.305 81.485 139.765 ;
        RECT 81.685 139.515 81.935 139.945 ;
        RECT 82.225 139.305 82.635 139.745 ;
        RECT 82.805 139.685 82.975 140.415 ;
        RECT 83.145 139.865 83.495 140.235 ;
        RECT 83.675 139.925 83.895 140.795 ;
        RECT 84.065 140.225 84.475 140.845 ;
        RECT 84.645 140.045 84.815 141.015 ;
        RECT 84.120 139.855 84.815 140.045 ;
        RECT 82.805 139.485 83.820 139.685 ;
        RECT 84.120 139.525 84.290 139.855 ;
        RECT 84.460 139.305 84.790 139.685 ;
        RECT 85.005 139.565 85.230 141.685 ;
        RECT 85.400 141.355 85.730 141.855 ;
        RECT 85.900 141.185 86.070 141.685 ;
        RECT 85.405 141.015 86.070 141.185 ;
        RECT 85.405 140.025 85.635 141.015 ;
        RECT 85.805 140.195 86.155 140.845 ;
        RECT 86.330 140.690 86.620 141.855 ;
        RECT 86.790 140.765 88.000 141.855 ;
        RECT 86.790 140.225 87.310 140.765 ;
        RECT 88.170 140.715 88.440 141.685 ;
        RECT 88.650 141.055 88.930 141.855 ;
        RECT 89.100 141.345 90.755 141.635 ;
        RECT 89.165 141.005 90.755 141.175 ;
        RECT 89.165 140.885 89.335 141.005 ;
        RECT 88.610 140.715 89.335 140.885 ;
        RECT 87.480 140.055 88.000 140.595 ;
        RECT 85.405 139.855 86.070 140.025 ;
        RECT 85.400 139.305 85.730 139.685 ;
        RECT 85.900 139.565 86.070 139.855 ;
        RECT 86.330 139.305 86.620 140.030 ;
        RECT 86.790 139.305 88.000 140.055 ;
        RECT 88.170 139.980 88.340 140.715 ;
        RECT 88.610 140.545 88.780 140.715 ;
        RECT 89.525 140.665 90.240 140.835 ;
        RECT 90.435 140.715 90.755 141.005 ;
        RECT 90.930 140.715 91.270 141.685 ;
        RECT 91.440 140.715 91.610 141.855 ;
        RECT 91.880 141.055 92.130 141.855 ;
        RECT 92.775 140.885 93.105 141.685 ;
        RECT 93.405 141.055 93.735 141.855 ;
        RECT 93.905 140.885 94.235 141.685 ;
        RECT 91.800 140.715 94.235 140.885 ;
        RECT 94.610 140.765 95.820 141.855 ;
        RECT 88.510 140.215 88.780 140.545 ;
        RECT 88.950 140.215 89.355 140.545 ;
        RECT 89.525 140.215 90.235 140.665 ;
        RECT 88.610 140.045 88.780 140.215 ;
        RECT 88.170 139.635 88.440 139.980 ;
        RECT 88.610 139.875 90.220 140.045 ;
        RECT 90.405 139.975 90.755 140.545 ;
        RECT 90.930 140.155 91.105 140.715 ;
        RECT 91.800 140.465 91.970 140.715 ;
        RECT 91.275 140.295 91.970 140.465 ;
        RECT 92.145 140.295 92.565 140.495 ;
        RECT 92.735 140.295 93.065 140.495 ;
        RECT 93.235 140.295 93.565 140.495 ;
        RECT 90.930 140.105 91.160 140.155 ;
        RECT 88.630 139.305 89.010 139.705 ;
        RECT 89.180 139.525 89.350 139.875 ;
        RECT 89.520 139.305 89.850 139.705 ;
        RECT 90.050 139.525 90.220 139.875 ;
        RECT 90.420 139.305 90.750 139.805 ;
        RECT 90.930 139.475 91.270 140.105 ;
        RECT 91.440 139.305 91.690 140.105 ;
        RECT 91.880 139.955 93.105 140.125 ;
        RECT 91.880 139.475 92.210 139.955 ;
        RECT 92.380 139.305 92.605 139.765 ;
        RECT 92.775 139.475 93.105 139.955 ;
        RECT 93.735 140.085 93.905 140.715 ;
        RECT 94.090 140.295 94.440 140.545 ;
        RECT 94.610 140.225 95.130 140.765 ;
        RECT 95.990 140.715 96.330 141.685 ;
        RECT 96.500 140.715 96.670 141.855 ;
        RECT 96.940 141.055 97.190 141.855 ;
        RECT 97.835 140.885 98.165 141.685 ;
        RECT 98.465 141.055 98.795 141.855 ;
        RECT 98.965 140.885 99.295 141.685 ;
        RECT 99.675 141.345 101.330 141.635 ;
        RECT 96.860 140.715 99.295 140.885 ;
        RECT 99.675 141.005 101.265 141.175 ;
        RECT 101.500 141.055 101.780 141.855 ;
        RECT 99.675 140.715 99.995 141.005 ;
        RECT 101.095 140.885 101.265 141.005 ;
        RECT 93.735 139.475 94.235 140.085 ;
        RECT 95.300 140.055 95.820 140.595 ;
        RECT 94.610 139.305 95.820 140.055 ;
        RECT 95.990 140.105 96.165 140.715 ;
        RECT 96.860 140.465 97.030 140.715 ;
        RECT 96.335 140.295 97.030 140.465 ;
        RECT 97.205 140.295 97.625 140.495 ;
        RECT 97.795 140.295 98.125 140.495 ;
        RECT 98.295 140.295 98.625 140.495 ;
        RECT 95.990 139.475 96.330 140.105 ;
        RECT 96.500 139.305 96.750 140.105 ;
        RECT 96.940 139.955 98.165 140.125 ;
        RECT 96.940 139.475 97.270 139.955 ;
        RECT 97.440 139.305 97.665 139.765 ;
        RECT 97.835 139.475 98.165 139.955 ;
        RECT 98.795 140.085 98.965 140.715 ;
        RECT 100.190 140.665 100.905 140.835 ;
        RECT 101.095 140.715 101.820 140.885 ;
        RECT 101.990 140.715 102.260 141.685 ;
        RECT 99.150 140.295 99.500 140.545 ;
        RECT 98.795 139.475 99.295 140.085 ;
        RECT 99.675 139.975 100.025 140.545 ;
        RECT 100.195 140.215 100.905 140.665 ;
        RECT 101.650 140.545 101.820 140.715 ;
        RECT 101.075 140.215 101.480 140.545 ;
        RECT 101.650 140.215 101.920 140.545 ;
        RECT 101.650 140.045 101.820 140.215 ;
        RECT 100.210 139.875 101.820 140.045 ;
        RECT 102.090 139.980 102.260 140.715 ;
        RECT 102.430 141.095 102.945 141.505 ;
        RECT 103.180 141.095 103.350 141.855 ;
        RECT 103.520 141.515 105.550 141.685 ;
        RECT 102.430 140.285 102.770 141.095 ;
        RECT 103.520 140.850 103.690 141.515 ;
        RECT 104.085 141.175 105.210 141.345 ;
        RECT 102.940 140.660 103.690 140.850 ;
        RECT 103.860 140.835 104.870 141.005 ;
        RECT 102.430 140.115 103.660 140.285 ;
        RECT 99.680 139.305 100.010 139.805 ;
        RECT 100.210 139.525 100.380 139.875 ;
        RECT 100.580 139.305 100.910 139.705 ;
        RECT 101.080 139.525 101.250 139.875 ;
        RECT 101.420 139.305 101.800 139.705 ;
        RECT 101.990 139.635 102.260 139.980 ;
        RECT 102.705 139.510 102.950 140.115 ;
        RECT 103.170 139.305 103.680 139.840 ;
        RECT 103.860 139.475 104.050 140.835 ;
        RECT 104.220 140.495 104.495 140.635 ;
        RECT 104.220 140.325 104.500 140.495 ;
        RECT 104.220 139.475 104.495 140.325 ;
        RECT 104.700 140.035 104.870 140.835 ;
        RECT 105.040 140.045 105.210 141.175 ;
        RECT 105.380 140.545 105.550 141.515 ;
        RECT 105.720 140.715 105.890 141.855 ;
        RECT 106.060 140.715 106.395 141.685 ;
        RECT 106.610 140.715 106.840 141.855 ;
        RECT 105.380 140.215 105.575 140.545 ;
        RECT 105.800 140.215 106.055 140.545 ;
        RECT 105.800 140.045 105.970 140.215 ;
        RECT 106.225 140.045 106.395 140.715 ;
        RECT 107.010 140.705 107.340 141.685 ;
        RECT 107.510 140.715 107.720 141.855 ;
        RECT 108.040 140.925 108.210 141.685 ;
        RECT 108.390 141.095 108.720 141.855 ;
        RECT 108.040 140.755 108.705 140.925 ;
        RECT 108.890 140.780 109.160 141.685 ;
        RECT 106.590 140.295 106.920 140.545 ;
        RECT 105.040 139.875 105.970 140.045 ;
        RECT 105.040 139.840 105.215 139.875 ;
        RECT 104.685 139.475 105.215 139.840 ;
        RECT 105.640 139.305 105.970 139.705 ;
        RECT 106.140 139.475 106.395 140.045 ;
        RECT 106.610 139.305 106.840 140.125 ;
        RECT 107.090 140.105 107.340 140.705 ;
        RECT 108.535 140.610 108.705 140.755 ;
        RECT 107.970 140.205 108.300 140.575 ;
        RECT 108.535 140.280 108.820 140.610 ;
        RECT 107.010 139.475 107.340 140.105 ;
        RECT 107.510 139.305 107.720 140.125 ;
        RECT 108.535 140.025 108.705 140.280 ;
        RECT 108.040 139.855 108.705 140.025 ;
        RECT 108.990 139.980 109.160 140.780 ;
        RECT 109.330 140.765 111.000 141.855 ;
        RECT 111.170 140.765 112.380 141.855 ;
        RECT 109.330 140.245 110.080 140.765 ;
        RECT 110.250 140.075 111.000 140.595 ;
        RECT 111.170 140.225 111.690 140.765 ;
        RECT 108.040 139.475 108.210 139.855 ;
        RECT 108.390 139.305 108.720 139.685 ;
        RECT 108.900 139.475 109.160 139.980 ;
        RECT 109.330 139.305 111.000 140.075 ;
        RECT 111.860 140.055 112.380 140.595 ;
        RECT 111.170 139.305 112.380 140.055 ;
        RECT 18.165 139.135 112.465 139.305 ;
        RECT 18.250 138.385 19.460 139.135 ;
        RECT 18.250 137.845 18.770 138.385 ;
        RECT 20.610 138.315 20.820 139.135 ;
        RECT 20.990 138.335 21.320 138.965 ;
        RECT 18.940 137.675 19.460 138.215 ;
        RECT 20.990 137.735 21.240 138.335 ;
        RECT 21.490 138.315 21.720 139.135 ;
        RECT 21.930 138.410 22.220 139.135 ;
        RECT 22.450 138.315 22.660 139.135 ;
        RECT 22.830 138.335 23.160 138.965 ;
        RECT 21.410 137.895 21.740 138.145 ;
        RECT 18.250 136.585 19.460 137.675 ;
        RECT 20.610 136.585 20.820 137.725 ;
        RECT 20.990 136.755 21.320 137.735 ;
        RECT 21.490 136.585 21.720 137.725 ;
        RECT 21.930 136.585 22.220 137.750 ;
        RECT 22.830 137.735 23.080 138.335 ;
        RECT 23.330 138.315 23.560 139.135 ;
        RECT 24.045 138.325 24.290 138.930 ;
        RECT 24.510 138.600 25.020 139.135 ;
        RECT 23.770 138.155 25.000 138.325 ;
        RECT 23.250 137.895 23.580 138.145 ;
        RECT 22.450 136.585 22.660 137.725 ;
        RECT 22.830 136.755 23.160 137.735 ;
        RECT 23.330 136.585 23.560 137.725 ;
        RECT 23.770 137.345 24.110 138.155 ;
        RECT 24.280 137.590 25.030 137.780 ;
        RECT 23.770 136.935 24.285 137.345 ;
        RECT 24.520 136.585 24.690 137.345 ;
        RECT 24.860 136.925 25.030 137.590 ;
        RECT 25.200 137.605 25.390 138.965 ;
        RECT 25.560 138.115 25.835 138.965 ;
        RECT 26.025 138.600 26.555 138.965 ;
        RECT 26.980 138.735 27.310 139.135 ;
        RECT 26.380 138.565 26.555 138.600 ;
        RECT 25.560 137.945 25.840 138.115 ;
        RECT 25.560 137.805 25.835 137.945 ;
        RECT 26.040 137.605 26.210 138.405 ;
        RECT 25.200 137.435 26.210 137.605 ;
        RECT 26.380 138.395 27.310 138.565 ;
        RECT 27.480 138.395 27.735 138.965 ;
        RECT 26.380 137.265 26.550 138.395 ;
        RECT 27.140 138.225 27.310 138.395 ;
        RECT 25.425 137.095 26.550 137.265 ;
        RECT 26.720 137.895 26.915 138.225 ;
        RECT 27.140 137.895 27.395 138.225 ;
        RECT 26.720 136.925 26.890 137.895 ;
        RECT 27.565 137.725 27.735 138.395 ;
        RECT 24.860 136.755 26.890 136.925 ;
        RECT 27.060 136.585 27.230 137.725 ;
        RECT 27.400 136.755 27.735 137.725 ;
        RECT 27.910 138.460 28.170 138.965 ;
        RECT 28.350 138.755 28.680 139.135 ;
        RECT 28.860 138.585 29.030 138.965 ;
        RECT 27.910 137.660 28.080 138.460 ;
        RECT 28.365 138.415 29.030 138.585 ;
        RECT 28.365 138.160 28.535 138.415 ;
        RECT 29.290 138.365 30.960 139.135 ;
        RECT 31.135 138.585 31.390 138.875 ;
        RECT 31.560 138.755 31.890 139.135 ;
        RECT 31.135 138.415 31.885 138.585 ;
        RECT 28.250 137.830 28.535 138.160 ;
        RECT 28.770 137.865 29.100 138.235 ;
        RECT 28.365 137.685 28.535 137.830 ;
        RECT 27.910 136.755 28.180 137.660 ;
        RECT 28.365 137.515 29.030 137.685 ;
        RECT 28.350 136.585 28.680 137.345 ;
        RECT 28.860 136.755 29.030 137.515 ;
        RECT 29.290 137.675 30.040 138.195 ;
        RECT 30.210 137.845 30.960 138.365 ;
        RECT 29.290 136.585 30.960 137.675 ;
        RECT 31.135 137.595 31.485 138.245 ;
        RECT 31.655 137.425 31.885 138.415 ;
        RECT 31.135 137.255 31.885 137.425 ;
        RECT 31.135 136.755 31.390 137.255 ;
        RECT 31.560 136.585 31.890 137.085 ;
        RECT 32.060 136.755 32.230 138.875 ;
        RECT 32.590 138.775 32.920 139.135 ;
        RECT 33.090 138.745 33.585 138.915 ;
        RECT 33.790 138.745 34.645 138.915 ;
        RECT 32.460 137.555 32.920 138.605 ;
        RECT 32.400 136.770 32.725 137.555 ;
        RECT 33.090 137.385 33.260 138.745 ;
        RECT 33.430 137.835 33.780 138.455 ;
        RECT 33.950 138.235 34.305 138.455 ;
        RECT 33.950 137.645 34.120 138.235 ;
        RECT 34.475 138.035 34.645 138.745 ;
        RECT 35.520 138.675 35.850 139.135 ;
        RECT 36.060 138.775 36.410 138.945 ;
        RECT 34.850 138.205 35.640 138.455 ;
        RECT 36.060 138.385 36.320 138.775 ;
        RECT 36.630 138.685 37.580 138.965 ;
        RECT 37.750 138.695 37.940 139.135 ;
        RECT 38.110 138.755 39.180 138.925 ;
        RECT 35.810 138.035 35.980 138.215 ;
        RECT 33.090 137.215 33.485 137.385 ;
        RECT 33.655 137.255 34.120 137.645 ;
        RECT 34.290 137.865 35.980 138.035 ;
        RECT 33.315 137.085 33.485 137.215 ;
        RECT 34.290 137.085 34.460 137.865 ;
        RECT 36.150 137.695 36.320 138.385 ;
        RECT 34.820 137.525 36.320 137.695 ;
        RECT 36.510 137.725 36.720 138.515 ;
        RECT 36.890 137.895 37.240 138.515 ;
        RECT 37.410 137.905 37.580 138.685 ;
        RECT 38.110 138.525 38.280 138.755 ;
        RECT 37.750 138.355 38.280 138.525 ;
        RECT 37.750 138.075 37.970 138.355 ;
        RECT 38.450 138.185 38.690 138.585 ;
        RECT 37.410 137.735 37.815 137.905 ;
        RECT 38.150 137.815 38.690 138.185 ;
        RECT 38.860 138.400 39.180 138.755 ;
        RECT 39.425 138.675 39.730 139.135 ;
        RECT 39.900 138.425 40.155 138.955 ;
        RECT 38.860 138.225 39.185 138.400 ;
        RECT 38.860 137.925 39.775 138.225 ;
        RECT 39.035 137.895 39.775 137.925 ;
        RECT 36.510 137.565 37.185 137.725 ;
        RECT 37.645 137.645 37.815 137.735 ;
        RECT 36.510 137.555 37.475 137.565 ;
        RECT 36.150 137.385 36.320 137.525 ;
        RECT 32.895 136.585 33.145 137.045 ;
        RECT 33.315 136.755 33.565 137.085 ;
        RECT 33.780 136.755 34.460 137.085 ;
        RECT 34.630 137.185 35.705 137.355 ;
        RECT 36.150 137.215 36.710 137.385 ;
        RECT 37.015 137.265 37.475 137.555 ;
        RECT 37.645 137.475 38.865 137.645 ;
        RECT 34.630 136.845 34.800 137.185 ;
        RECT 35.035 136.585 35.365 137.015 ;
        RECT 35.535 136.845 35.705 137.185 ;
        RECT 36.000 136.585 36.370 137.045 ;
        RECT 36.540 136.755 36.710 137.215 ;
        RECT 37.645 137.095 37.815 137.475 ;
        RECT 39.035 137.305 39.205 137.895 ;
        RECT 39.945 137.775 40.155 138.425 ;
        RECT 36.945 136.755 37.815 137.095 ;
        RECT 38.405 137.135 39.205 137.305 ;
        RECT 37.985 136.585 38.235 137.045 ;
        RECT 38.405 136.845 38.575 137.135 ;
        RECT 38.755 136.585 39.085 136.965 ;
        RECT 39.425 136.585 39.730 137.725 ;
        RECT 39.900 136.895 40.155 137.775 ;
        RECT 40.330 138.460 40.600 138.805 ;
        RECT 40.790 138.735 41.170 139.135 ;
        RECT 41.340 138.565 41.510 138.915 ;
        RECT 41.680 138.735 42.010 139.135 ;
        RECT 42.210 138.565 42.380 138.915 ;
        RECT 42.580 138.635 42.910 139.135 ;
        RECT 40.330 137.725 40.500 138.460 ;
        RECT 40.770 138.395 42.380 138.565 ;
        RECT 40.770 138.225 40.940 138.395 ;
        RECT 40.670 137.895 40.940 138.225 ;
        RECT 41.110 137.895 41.515 138.225 ;
        RECT 40.770 137.725 40.940 137.895 ;
        RECT 41.685 137.775 42.395 138.225 ;
        RECT 42.565 137.895 42.915 138.465 ;
        RECT 43.755 138.355 44.255 138.965 ;
        RECT 43.550 137.895 43.900 138.145 ;
        RECT 40.330 136.755 40.600 137.725 ;
        RECT 40.770 137.555 41.495 137.725 ;
        RECT 41.685 137.605 42.400 137.775 ;
        RECT 44.085 137.725 44.255 138.355 ;
        RECT 44.885 138.485 45.215 138.965 ;
        RECT 45.385 138.675 45.610 139.135 ;
        RECT 45.780 138.485 46.110 138.965 ;
        RECT 44.885 138.315 46.110 138.485 ;
        RECT 46.300 138.335 46.550 139.135 ;
        RECT 46.720 138.335 47.060 138.965 ;
        RECT 47.690 138.410 47.980 139.135 ;
        RECT 44.425 137.945 44.755 138.145 ;
        RECT 44.925 137.945 45.255 138.145 ;
        RECT 45.425 137.945 45.845 138.145 ;
        RECT 46.020 137.975 46.715 138.145 ;
        RECT 46.020 137.725 46.190 137.975 ;
        RECT 46.885 137.725 47.060 138.335 ;
        RECT 48.610 138.335 48.950 138.965 ;
        RECT 49.120 138.335 49.370 139.135 ;
        RECT 49.560 138.485 49.890 138.965 ;
        RECT 50.060 138.675 50.285 139.135 ;
        RECT 50.455 138.485 50.785 138.965 ;
        RECT 41.325 137.435 41.495 137.555 ;
        RECT 42.595 137.435 42.915 137.725 ;
        RECT 40.810 136.585 41.090 137.385 ;
        RECT 41.325 137.265 42.915 137.435 ;
        RECT 43.755 137.555 46.190 137.725 ;
        RECT 41.260 136.805 42.915 137.095 ;
        RECT 43.755 136.755 44.085 137.555 ;
        RECT 44.255 136.585 44.585 137.385 ;
        RECT 44.885 136.755 45.215 137.555 ;
        RECT 45.860 136.585 46.110 137.385 ;
        RECT 46.380 136.585 46.550 137.725 ;
        RECT 46.720 136.755 47.060 137.725 ;
        RECT 47.690 136.585 47.980 137.750 ;
        RECT 48.610 137.725 48.785 138.335 ;
        RECT 49.560 138.315 50.785 138.485 ;
        RECT 51.415 138.355 51.915 138.965 ;
        RECT 52.665 138.425 52.920 138.955 ;
        RECT 53.100 138.675 53.385 139.135 ;
        RECT 48.955 137.975 49.650 138.145 ;
        RECT 49.480 137.725 49.650 137.975 ;
        RECT 49.825 137.945 50.245 138.145 ;
        RECT 50.415 137.945 50.745 138.145 ;
        RECT 50.915 137.945 51.245 138.145 ;
        RECT 51.415 137.725 51.585 138.355 ;
        RECT 51.770 137.895 52.120 138.145 ;
        RECT 48.610 136.755 48.950 137.725 ;
        RECT 49.120 136.585 49.290 137.725 ;
        RECT 49.480 137.555 51.915 137.725 ;
        RECT 49.560 136.585 49.810 137.385 ;
        RECT 50.455 136.755 50.785 137.555 ;
        RECT 51.085 136.585 51.415 137.385 ;
        RECT 51.585 136.755 51.915 137.555 ;
        RECT 52.665 137.565 52.845 138.425 ;
        RECT 53.565 138.225 53.815 138.875 ;
        RECT 53.015 137.895 53.815 138.225 ;
        RECT 52.665 137.095 52.920 137.565 ;
        RECT 52.580 136.925 52.920 137.095 ;
        RECT 52.665 136.895 52.920 136.925 ;
        RECT 53.100 136.585 53.385 137.385 ;
        RECT 53.565 137.305 53.815 137.895 ;
        RECT 54.015 138.540 54.335 138.870 ;
        RECT 54.515 138.655 55.175 139.135 ;
        RECT 55.375 138.745 56.225 138.915 ;
        RECT 54.015 137.645 54.205 138.540 ;
        RECT 54.525 138.215 55.185 138.485 ;
        RECT 54.855 138.155 55.185 138.215 ;
        RECT 54.375 137.985 54.705 138.045 ;
        RECT 55.375 137.985 55.545 138.745 ;
        RECT 56.785 138.675 57.105 139.135 ;
        RECT 57.305 138.495 57.555 138.925 ;
        RECT 57.845 138.695 58.255 139.135 ;
        RECT 58.425 138.755 59.440 138.955 ;
        RECT 55.715 138.325 56.965 138.495 ;
        RECT 55.715 138.205 56.045 138.325 ;
        RECT 54.375 137.815 56.275 137.985 ;
        RECT 54.015 137.475 55.935 137.645 ;
        RECT 54.015 137.455 54.335 137.475 ;
        RECT 53.565 136.795 53.895 137.305 ;
        RECT 54.165 136.845 54.335 137.455 ;
        RECT 56.105 137.305 56.275 137.815 ;
        RECT 56.445 137.745 56.625 138.155 ;
        RECT 56.795 137.565 56.965 138.325 ;
        RECT 54.505 136.585 54.835 137.275 ;
        RECT 55.065 137.135 56.275 137.305 ;
        RECT 56.445 137.255 56.965 137.565 ;
        RECT 57.135 138.155 57.555 138.495 ;
        RECT 57.845 138.155 58.255 138.485 ;
        RECT 57.135 137.385 57.325 138.155 ;
        RECT 58.425 138.025 58.595 138.755 ;
        RECT 59.740 138.585 59.910 138.915 ;
        RECT 60.080 138.755 60.410 139.135 ;
        RECT 58.765 138.205 59.115 138.575 ;
        RECT 58.425 137.985 58.845 138.025 ;
        RECT 57.495 137.815 58.845 137.985 ;
        RECT 57.495 137.655 57.745 137.815 ;
        RECT 58.255 137.385 58.505 137.645 ;
        RECT 57.135 137.135 58.505 137.385 ;
        RECT 55.065 136.845 55.305 137.135 ;
        RECT 56.105 137.055 56.275 137.135 ;
        RECT 55.505 136.585 55.925 136.965 ;
        RECT 56.105 136.805 56.735 137.055 ;
        RECT 57.205 136.585 57.535 136.965 ;
        RECT 57.705 136.845 57.875 137.135 ;
        RECT 58.675 136.970 58.845 137.815 ;
        RECT 59.295 137.645 59.515 138.515 ;
        RECT 59.740 138.395 60.435 138.585 ;
        RECT 59.015 137.265 59.515 137.645 ;
        RECT 59.685 137.595 60.095 138.215 ;
        RECT 60.265 137.425 60.435 138.395 ;
        RECT 59.740 137.255 60.435 137.425 ;
        RECT 58.055 136.585 58.435 136.965 ;
        RECT 58.675 136.800 59.505 136.970 ;
        RECT 59.740 136.755 59.910 137.255 ;
        RECT 60.080 136.585 60.410 137.085 ;
        RECT 60.625 136.755 60.850 138.875 ;
        RECT 61.020 138.755 61.350 139.135 ;
        RECT 61.520 138.585 61.690 138.875 ;
        RECT 61.025 138.415 61.690 138.585 ;
        RECT 61.950 138.460 62.210 138.965 ;
        RECT 62.390 138.755 62.720 139.135 ;
        RECT 62.900 138.585 63.070 138.965 ;
        RECT 61.025 137.425 61.255 138.415 ;
        RECT 61.425 137.595 61.775 138.245 ;
        RECT 61.950 137.660 62.120 138.460 ;
        RECT 62.405 138.415 63.070 138.585 ;
        RECT 62.405 138.160 62.575 138.415 ;
        RECT 63.335 138.295 63.595 139.135 ;
        RECT 63.770 138.390 64.025 138.965 ;
        RECT 64.195 138.755 64.525 139.135 ;
        RECT 64.740 138.585 64.910 138.965 ;
        RECT 64.195 138.415 64.910 138.585 ;
        RECT 65.260 138.585 65.430 138.965 ;
        RECT 65.645 138.755 65.975 139.135 ;
        RECT 65.260 138.415 65.975 138.585 ;
        RECT 62.290 137.830 62.575 138.160 ;
        RECT 62.810 137.865 63.140 138.235 ;
        RECT 62.405 137.685 62.575 137.830 ;
        RECT 61.025 137.255 61.690 137.425 ;
        RECT 61.020 136.585 61.350 137.085 ;
        RECT 61.520 136.755 61.690 137.255 ;
        RECT 61.950 136.755 62.220 137.660 ;
        RECT 62.405 137.515 63.070 137.685 ;
        RECT 62.390 136.585 62.720 137.345 ;
        RECT 62.900 136.755 63.070 137.515 ;
        RECT 63.335 136.585 63.595 137.735 ;
        RECT 63.770 137.660 63.940 138.390 ;
        RECT 64.195 138.225 64.365 138.415 ;
        RECT 64.110 137.895 64.365 138.225 ;
        RECT 64.195 137.685 64.365 137.895 ;
        RECT 64.645 137.865 65.000 138.235 ;
        RECT 65.170 137.865 65.525 138.235 ;
        RECT 65.805 138.225 65.975 138.415 ;
        RECT 66.145 138.390 66.400 138.965 ;
        RECT 65.805 137.895 66.060 138.225 ;
        RECT 65.805 137.685 65.975 137.895 ;
        RECT 63.770 136.755 64.025 137.660 ;
        RECT 64.195 137.515 64.910 137.685 ;
        RECT 64.195 136.585 64.525 137.345 ;
        RECT 64.740 136.755 64.910 137.515 ;
        RECT 65.260 137.515 65.975 137.685 ;
        RECT 66.230 137.660 66.400 138.390 ;
        RECT 66.575 138.295 66.835 139.135 ;
        RECT 67.100 138.585 67.270 138.965 ;
        RECT 67.485 138.755 67.815 139.135 ;
        RECT 67.100 138.415 67.815 138.585 ;
        RECT 67.010 137.865 67.365 138.235 ;
        RECT 67.645 138.225 67.815 138.415 ;
        RECT 67.985 138.390 68.240 138.965 ;
        RECT 67.645 137.895 67.900 138.225 ;
        RECT 65.260 136.755 65.430 137.515 ;
        RECT 65.645 136.585 65.975 137.345 ;
        RECT 66.145 136.755 66.400 137.660 ;
        RECT 66.575 136.585 66.835 137.735 ;
        RECT 67.645 137.685 67.815 137.895 ;
        RECT 67.100 137.515 67.815 137.685 ;
        RECT 68.070 137.660 68.240 138.390 ;
        RECT 68.415 138.295 68.675 139.135 ;
        RECT 69.770 138.335 70.110 138.965 ;
        RECT 70.280 138.335 70.530 139.135 ;
        RECT 70.720 138.485 71.050 138.965 ;
        RECT 71.220 138.675 71.445 139.135 ;
        RECT 71.615 138.485 71.945 138.965 ;
        RECT 67.100 136.755 67.270 137.515 ;
        RECT 67.485 136.585 67.815 137.345 ;
        RECT 67.985 136.755 68.240 137.660 ;
        RECT 68.415 136.585 68.675 137.735 ;
        RECT 69.770 137.725 69.945 138.335 ;
        RECT 70.720 138.315 71.945 138.485 ;
        RECT 72.575 138.355 73.075 138.965 ;
        RECT 73.450 138.410 73.740 139.135 ;
        RECT 70.115 137.975 70.810 138.145 ;
        RECT 70.640 137.725 70.810 137.975 ;
        RECT 70.985 137.945 71.405 138.145 ;
        RECT 71.575 137.945 71.905 138.145 ;
        RECT 72.075 137.945 72.405 138.145 ;
        RECT 72.575 137.725 72.745 138.355 ;
        RECT 73.910 138.335 74.250 138.965 ;
        RECT 74.420 138.335 74.670 139.135 ;
        RECT 74.860 138.485 75.190 138.965 ;
        RECT 75.360 138.675 75.585 139.135 ;
        RECT 75.755 138.485 76.085 138.965 ;
        RECT 72.930 137.895 73.280 138.145 ;
        RECT 69.770 136.755 70.110 137.725 ;
        RECT 70.280 136.585 70.450 137.725 ;
        RECT 70.640 137.555 73.075 137.725 ;
        RECT 70.720 136.585 70.970 137.385 ;
        RECT 71.615 136.755 71.945 137.555 ;
        RECT 72.245 136.585 72.575 137.385 ;
        RECT 72.745 136.755 73.075 137.555 ;
        RECT 73.450 136.585 73.740 137.750 ;
        RECT 73.910 137.725 74.085 138.335 ;
        RECT 74.860 138.315 76.085 138.485 ;
        RECT 76.715 138.355 77.215 138.965 ;
        RECT 78.050 138.365 79.720 139.135 ;
        RECT 74.255 137.975 74.950 138.145 ;
        RECT 74.780 137.725 74.950 137.975 ;
        RECT 75.125 137.945 75.545 138.145 ;
        RECT 75.715 137.945 76.045 138.145 ;
        RECT 76.215 137.945 76.545 138.145 ;
        RECT 76.715 137.725 76.885 138.355 ;
        RECT 77.070 137.895 77.420 138.145 ;
        RECT 73.910 136.755 74.250 137.725 ;
        RECT 74.420 136.585 74.590 137.725 ;
        RECT 74.780 137.555 77.215 137.725 ;
        RECT 74.860 136.585 75.110 137.385 ;
        RECT 75.755 136.755 76.085 137.555 ;
        RECT 76.385 136.585 76.715 137.385 ;
        RECT 76.885 136.755 77.215 137.555 ;
        RECT 78.050 137.675 78.800 138.195 ;
        RECT 78.970 137.845 79.720 138.365 ;
        RECT 80.165 138.325 80.410 138.930 ;
        RECT 80.630 138.600 81.140 139.135 ;
        RECT 79.890 138.155 81.120 138.325 ;
        RECT 78.050 136.585 79.720 137.675 ;
        RECT 79.890 137.345 80.230 138.155 ;
        RECT 80.400 137.590 81.150 137.780 ;
        RECT 79.890 136.935 80.405 137.345 ;
        RECT 80.640 136.585 80.810 137.345 ;
        RECT 80.980 136.925 81.150 137.590 ;
        RECT 81.320 137.605 81.510 138.965 ;
        RECT 81.680 138.115 81.955 138.965 ;
        RECT 82.145 138.600 82.675 138.965 ;
        RECT 83.100 138.735 83.430 139.135 ;
        RECT 82.500 138.565 82.675 138.600 ;
        RECT 81.680 137.945 81.960 138.115 ;
        RECT 81.680 137.805 81.955 137.945 ;
        RECT 82.160 137.605 82.330 138.405 ;
        RECT 81.320 137.435 82.330 137.605 ;
        RECT 82.500 138.395 83.430 138.565 ;
        RECT 83.600 138.395 83.855 138.965 ;
        RECT 82.500 137.265 82.670 138.395 ;
        RECT 83.260 138.225 83.430 138.395 ;
        RECT 81.545 137.095 82.670 137.265 ;
        RECT 82.840 137.895 83.035 138.225 ;
        RECT 83.260 137.895 83.515 138.225 ;
        RECT 82.840 136.925 83.010 137.895 ;
        RECT 83.685 137.725 83.855 138.395 ;
        RECT 84.090 138.315 84.300 139.135 ;
        RECT 84.470 138.335 84.800 138.965 ;
        RECT 84.470 137.735 84.720 138.335 ;
        RECT 84.970 138.315 85.200 139.135 ;
        RECT 85.410 138.460 85.670 138.965 ;
        RECT 85.850 138.755 86.180 139.135 ;
        RECT 86.360 138.585 86.530 138.965 ;
        RECT 84.890 137.895 85.220 138.145 ;
        RECT 80.980 136.755 83.010 136.925 ;
        RECT 83.180 136.585 83.350 137.725 ;
        RECT 83.520 136.755 83.855 137.725 ;
        RECT 84.090 136.585 84.300 137.725 ;
        RECT 84.470 136.755 84.800 137.735 ;
        RECT 84.970 136.585 85.200 137.725 ;
        RECT 85.410 137.660 85.580 138.460 ;
        RECT 85.865 138.415 86.530 138.585 ;
        RECT 85.865 138.160 86.035 138.415 ;
        RECT 86.790 138.385 88.000 139.135 ;
        RECT 88.175 138.590 93.520 139.135 ;
        RECT 93.700 138.635 94.030 139.135 ;
        RECT 85.750 137.830 86.035 138.160 ;
        RECT 86.270 137.865 86.600 138.235 ;
        RECT 85.865 137.685 86.035 137.830 ;
        RECT 85.410 136.755 85.680 137.660 ;
        RECT 85.865 137.515 86.530 137.685 ;
        RECT 85.850 136.585 86.180 137.345 ;
        RECT 86.360 136.755 86.530 137.515 ;
        RECT 86.790 137.675 87.310 138.215 ;
        RECT 87.480 137.845 88.000 138.385 ;
        RECT 86.790 136.585 88.000 137.675 ;
        RECT 89.765 137.020 90.115 138.270 ;
        RECT 91.595 137.760 91.935 138.590 ;
        RECT 94.230 138.565 94.400 138.915 ;
        RECT 94.600 138.735 94.930 139.135 ;
        RECT 95.100 138.565 95.270 138.915 ;
        RECT 95.440 138.735 95.820 139.135 ;
        RECT 93.695 137.895 94.045 138.465 ;
        RECT 94.230 138.395 95.840 138.565 ;
        RECT 96.010 138.460 96.280 138.805 ;
        RECT 95.670 138.225 95.840 138.395 ;
        RECT 93.695 137.435 94.015 137.725 ;
        RECT 94.215 137.605 94.925 138.225 ;
        RECT 95.095 137.895 95.500 138.225 ;
        RECT 95.670 137.895 95.940 138.225 ;
        RECT 95.670 137.725 95.840 137.895 ;
        RECT 96.110 137.725 96.280 138.460 ;
        RECT 96.540 138.485 96.710 138.965 ;
        RECT 96.890 138.655 97.130 139.135 ;
        RECT 97.380 138.485 97.550 138.965 ;
        RECT 97.720 138.655 98.050 139.135 ;
        RECT 98.220 138.485 98.390 138.965 ;
        RECT 96.540 138.315 97.175 138.485 ;
        RECT 97.380 138.315 98.390 138.485 ;
        RECT 98.560 138.335 98.890 139.135 ;
        RECT 99.210 138.410 99.500 139.135 ;
        RECT 100.170 138.315 100.400 139.135 ;
        RECT 100.570 138.335 100.900 138.965 ;
        RECT 97.005 138.145 97.175 138.315 ;
        RECT 96.455 137.905 96.835 138.145 ;
        RECT 97.005 137.975 97.505 138.145 ;
        RECT 97.005 137.735 97.175 137.975 ;
        RECT 97.895 137.775 98.390 138.315 ;
        RECT 100.150 137.895 100.480 138.145 ;
        RECT 95.115 137.555 95.840 137.725 ;
        RECT 95.115 137.435 95.285 137.555 ;
        RECT 93.695 137.265 95.285 137.435 ;
        RECT 88.175 136.585 93.520 137.020 ;
        RECT 93.695 136.805 95.350 137.095 ;
        RECT 95.520 136.585 95.800 137.385 ;
        RECT 96.010 136.755 96.280 137.725 ;
        RECT 96.460 137.565 97.175 137.735 ;
        RECT 97.380 137.605 98.390 137.775 ;
        RECT 96.460 136.755 96.790 137.565 ;
        RECT 96.960 136.585 97.200 137.385 ;
        RECT 97.380 136.755 97.550 137.605 ;
        RECT 97.720 136.585 98.050 137.385 ;
        RECT 98.220 136.755 98.390 137.605 ;
        RECT 98.560 136.585 98.890 137.735 ;
        RECT 99.210 136.585 99.500 137.750 ;
        RECT 100.650 137.735 100.900 138.335 ;
        RECT 101.070 138.315 101.280 139.135 ;
        RECT 101.885 138.795 102.140 138.955 ;
        RECT 101.800 138.625 102.140 138.795 ;
        RECT 102.320 138.675 102.605 139.135 ;
        RECT 101.885 138.425 102.140 138.625 ;
        RECT 100.170 136.585 100.400 137.725 ;
        RECT 100.570 136.755 100.900 137.735 ;
        RECT 101.070 136.585 101.280 137.725 ;
        RECT 101.885 137.565 102.065 138.425 ;
        RECT 102.785 138.225 103.035 138.875 ;
        RECT 102.235 137.895 103.035 138.225 ;
        RECT 101.885 136.895 102.140 137.565 ;
        RECT 102.320 136.585 102.605 137.385 ;
        RECT 102.785 137.305 103.035 137.895 ;
        RECT 103.235 138.540 103.555 138.870 ;
        RECT 103.735 138.655 104.395 139.135 ;
        RECT 104.595 138.745 105.445 138.915 ;
        RECT 103.235 137.645 103.425 138.540 ;
        RECT 103.745 138.215 104.405 138.485 ;
        RECT 104.075 138.155 104.405 138.215 ;
        RECT 103.595 137.985 103.925 138.045 ;
        RECT 104.595 137.985 104.765 138.745 ;
        RECT 106.005 138.675 106.325 139.135 ;
        RECT 106.525 138.495 106.775 138.925 ;
        RECT 107.065 138.695 107.475 139.135 ;
        RECT 107.645 138.755 108.660 138.955 ;
        RECT 104.935 138.325 106.185 138.495 ;
        RECT 104.935 138.205 105.265 138.325 ;
        RECT 103.595 137.815 105.495 137.985 ;
        RECT 103.235 137.475 105.155 137.645 ;
        RECT 103.235 137.455 103.555 137.475 ;
        RECT 102.785 136.795 103.115 137.305 ;
        RECT 103.385 136.845 103.555 137.455 ;
        RECT 105.325 137.305 105.495 137.815 ;
        RECT 105.665 137.745 105.845 138.155 ;
        RECT 106.015 137.565 106.185 138.325 ;
        RECT 103.725 136.585 104.055 137.275 ;
        RECT 104.285 137.135 105.495 137.305 ;
        RECT 105.665 137.255 106.185 137.565 ;
        RECT 106.355 138.155 106.775 138.495 ;
        RECT 107.065 138.155 107.475 138.485 ;
        RECT 106.355 137.385 106.545 138.155 ;
        RECT 107.645 138.025 107.815 138.755 ;
        RECT 108.960 138.585 109.130 138.915 ;
        RECT 109.300 138.755 109.630 139.135 ;
        RECT 107.985 138.205 108.335 138.575 ;
        RECT 107.645 137.985 108.065 138.025 ;
        RECT 106.715 137.815 108.065 137.985 ;
        RECT 106.715 137.655 106.965 137.815 ;
        RECT 107.475 137.385 107.725 137.645 ;
        RECT 106.355 137.135 107.725 137.385 ;
        RECT 104.285 136.845 104.525 137.135 ;
        RECT 105.325 137.055 105.495 137.135 ;
        RECT 104.725 136.585 105.145 136.965 ;
        RECT 105.325 136.805 105.955 137.055 ;
        RECT 106.425 136.585 106.755 136.965 ;
        RECT 106.925 136.845 107.095 137.135 ;
        RECT 107.895 136.970 108.065 137.815 ;
        RECT 108.515 137.645 108.735 138.515 ;
        RECT 108.960 138.395 109.655 138.585 ;
        RECT 108.235 137.265 108.735 137.645 ;
        RECT 108.905 137.595 109.315 138.215 ;
        RECT 109.485 137.425 109.655 138.395 ;
        RECT 108.960 137.255 109.655 137.425 ;
        RECT 107.275 136.585 107.655 136.965 ;
        RECT 107.895 136.800 108.725 136.970 ;
        RECT 108.960 136.755 109.130 137.255 ;
        RECT 109.300 136.585 109.630 137.085 ;
        RECT 109.845 136.755 110.070 138.875 ;
        RECT 110.240 138.755 110.570 139.135 ;
        RECT 110.740 138.585 110.910 138.875 ;
        RECT 110.245 138.415 110.910 138.585 ;
        RECT 110.245 137.425 110.475 138.415 ;
        RECT 111.170 138.385 112.380 139.135 ;
        RECT 110.645 137.595 110.995 138.245 ;
        RECT 111.170 137.675 111.690 138.215 ;
        RECT 111.860 137.845 112.380 138.385 ;
        RECT 110.245 137.255 110.910 137.425 ;
        RECT 110.240 136.585 110.570 137.085 ;
        RECT 110.740 136.755 110.910 137.255 ;
        RECT 111.170 136.585 112.380 137.675 ;
        RECT 18.165 136.415 112.465 136.585 ;
        RECT 18.250 135.325 19.460 136.415 ;
        RECT 18.250 134.615 18.770 135.155 ;
        RECT 18.940 134.785 19.460 135.325 ;
        RECT 20.095 135.225 20.350 136.105 ;
        RECT 20.520 135.275 20.825 136.415 ;
        RECT 21.165 136.035 21.495 136.415 ;
        RECT 21.675 135.865 21.845 136.155 ;
        RECT 22.015 135.955 22.265 136.415 ;
        RECT 21.045 135.695 21.845 135.865 ;
        RECT 22.435 135.905 23.305 136.245 ;
        RECT 18.250 133.865 19.460 134.615 ;
        RECT 20.095 134.575 20.305 135.225 ;
        RECT 21.045 135.105 21.215 135.695 ;
        RECT 22.435 135.525 22.605 135.905 ;
        RECT 23.540 135.785 23.710 136.245 ;
        RECT 23.880 135.955 24.250 136.415 ;
        RECT 24.545 135.815 24.715 136.155 ;
        RECT 24.885 135.985 25.215 136.415 ;
        RECT 25.450 135.815 25.620 136.155 ;
        RECT 21.385 135.355 22.605 135.525 ;
        RECT 22.775 135.445 23.235 135.735 ;
        RECT 23.540 135.615 24.100 135.785 ;
        RECT 24.545 135.645 25.620 135.815 ;
        RECT 25.790 135.915 26.470 136.245 ;
        RECT 26.685 135.915 26.935 136.245 ;
        RECT 27.105 135.955 27.355 136.415 ;
        RECT 23.930 135.475 24.100 135.615 ;
        RECT 22.775 135.435 23.740 135.445 ;
        RECT 22.435 135.265 22.605 135.355 ;
        RECT 23.065 135.275 23.740 135.435 ;
        RECT 20.475 135.075 21.215 135.105 ;
        RECT 20.475 134.775 21.390 135.075 ;
        RECT 21.065 134.600 21.390 134.775 ;
        RECT 20.095 134.045 20.350 134.575 ;
        RECT 20.520 133.865 20.825 134.325 ;
        RECT 21.070 134.245 21.390 134.600 ;
        RECT 21.560 134.815 22.100 135.185 ;
        RECT 22.435 135.095 22.840 135.265 ;
        RECT 21.560 134.415 21.800 134.815 ;
        RECT 22.280 134.645 22.500 134.925 ;
        RECT 21.970 134.475 22.500 134.645 ;
        RECT 21.970 134.245 22.140 134.475 ;
        RECT 22.670 134.315 22.840 135.095 ;
        RECT 23.010 134.485 23.360 135.105 ;
        RECT 23.530 134.485 23.740 135.275 ;
        RECT 23.930 135.305 25.430 135.475 ;
        RECT 23.930 134.615 24.100 135.305 ;
        RECT 25.790 135.135 25.960 135.915 ;
        RECT 26.765 135.785 26.935 135.915 ;
        RECT 24.270 134.965 25.960 135.135 ;
        RECT 26.130 135.355 26.595 135.745 ;
        RECT 26.765 135.615 27.160 135.785 ;
        RECT 24.270 134.785 24.440 134.965 ;
        RECT 21.070 134.075 22.140 134.245 ;
        RECT 22.310 133.865 22.500 134.305 ;
        RECT 22.670 134.035 23.620 134.315 ;
        RECT 23.930 134.225 24.190 134.615 ;
        RECT 24.610 134.545 25.400 134.795 ;
        RECT 23.840 134.055 24.190 134.225 ;
        RECT 24.400 133.865 24.730 134.325 ;
        RECT 25.605 134.255 25.775 134.965 ;
        RECT 26.130 134.765 26.300 135.355 ;
        RECT 25.945 134.545 26.300 134.765 ;
        RECT 26.470 134.545 26.820 135.165 ;
        RECT 26.990 134.255 27.160 135.615 ;
        RECT 27.525 135.445 27.850 136.230 ;
        RECT 27.330 134.395 27.790 135.445 ;
        RECT 25.605 134.085 26.460 134.255 ;
        RECT 26.665 134.085 27.160 134.255 ;
        RECT 27.330 133.865 27.660 134.225 ;
        RECT 28.020 134.125 28.190 136.245 ;
        RECT 28.360 135.915 28.690 136.415 ;
        RECT 28.860 135.745 29.115 136.245 ;
        RECT 28.365 135.575 29.115 135.745 ;
        RECT 28.365 134.585 28.595 135.575 ;
        RECT 28.765 134.755 29.115 135.405 ;
        RECT 29.330 135.275 29.560 136.415 ;
        RECT 29.730 135.265 30.060 136.245 ;
        RECT 30.230 135.275 30.440 136.415 ;
        RECT 30.670 135.655 31.185 136.065 ;
        RECT 31.420 135.655 31.590 136.415 ;
        RECT 31.760 136.075 33.790 136.245 ;
        RECT 29.310 134.855 29.640 135.105 ;
        RECT 28.365 134.415 29.115 134.585 ;
        RECT 28.360 133.865 28.690 134.245 ;
        RECT 28.860 134.125 29.115 134.415 ;
        RECT 29.330 133.865 29.560 134.685 ;
        RECT 29.810 134.665 30.060 135.265 ;
        RECT 30.670 134.845 31.010 135.655 ;
        RECT 31.760 135.410 31.930 136.075 ;
        RECT 32.325 135.735 33.450 135.905 ;
        RECT 31.180 135.220 31.930 135.410 ;
        RECT 32.100 135.395 33.110 135.565 ;
        RECT 29.730 134.035 30.060 134.665 ;
        RECT 30.230 133.865 30.440 134.685 ;
        RECT 30.670 134.675 31.900 134.845 ;
        RECT 30.945 134.070 31.190 134.675 ;
        RECT 31.410 133.865 31.920 134.400 ;
        RECT 32.100 134.035 32.290 135.395 ;
        RECT 32.460 135.055 32.735 135.195 ;
        RECT 32.460 134.885 32.740 135.055 ;
        RECT 32.460 134.035 32.735 134.885 ;
        RECT 32.940 134.595 33.110 135.395 ;
        RECT 33.280 134.605 33.450 135.735 ;
        RECT 33.620 135.105 33.790 136.075 ;
        RECT 33.960 135.275 34.130 136.415 ;
        RECT 34.300 135.275 34.635 136.245 ;
        RECT 33.620 134.775 33.815 135.105 ;
        RECT 34.040 134.775 34.295 135.105 ;
        RECT 34.040 134.605 34.210 134.775 ;
        RECT 34.465 134.605 34.635 135.275 ;
        RECT 34.810 135.250 35.100 136.415 ;
        RECT 35.275 135.275 35.610 136.245 ;
        RECT 35.780 135.275 35.950 136.415 ;
        RECT 36.120 136.075 38.150 136.245 ;
        RECT 33.280 134.435 34.210 134.605 ;
        RECT 33.280 134.400 33.455 134.435 ;
        RECT 32.925 134.035 33.455 134.400 ;
        RECT 33.880 133.865 34.210 134.265 ;
        RECT 34.380 134.035 34.635 134.605 ;
        RECT 35.275 134.605 35.445 135.275 ;
        RECT 36.120 135.105 36.290 136.075 ;
        RECT 35.615 134.775 35.870 135.105 ;
        RECT 36.095 134.775 36.290 135.105 ;
        RECT 36.460 135.735 37.585 135.905 ;
        RECT 35.700 134.605 35.870 134.775 ;
        RECT 36.460 134.605 36.630 135.735 ;
        RECT 34.810 133.865 35.100 134.590 ;
        RECT 35.275 134.035 35.530 134.605 ;
        RECT 35.700 134.435 36.630 134.605 ;
        RECT 36.800 135.395 37.810 135.565 ;
        RECT 36.800 134.595 36.970 135.395 ;
        RECT 37.175 134.715 37.450 135.195 ;
        RECT 37.170 134.545 37.450 134.715 ;
        RECT 36.455 134.400 36.630 134.435 ;
        RECT 35.700 133.865 36.030 134.265 ;
        RECT 36.455 134.035 36.985 134.400 ;
        RECT 37.175 134.035 37.450 134.545 ;
        RECT 37.620 134.035 37.810 135.395 ;
        RECT 37.980 135.410 38.150 136.075 ;
        RECT 38.320 135.655 38.490 136.415 ;
        RECT 38.725 135.655 39.240 136.065 ;
        RECT 37.980 135.220 38.730 135.410 ;
        RECT 38.900 134.845 39.240 135.655 ;
        RECT 38.010 134.675 39.240 134.845 ;
        RECT 39.870 135.275 40.140 136.245 ;
        RECT 40.350 135.615 40.630 136.415 ;
        RECT 40.800 135.905 42.455 136.195 ;
        RECT 40.865 135.565 42.455 135.735 ;
        RECT 40.865 135.445 41.035 135.565 ;
        RECT 40.310 135.275 41.035 135.445 ;
        RECT 37.990 133.865 38.500 134.400 ;
        RECT 38.720 134.070 38.965 134.675 ;
        RECT 39.870 134.540 40.040 135.275 ;
        RECT 40.310 135.105 40.480 135.275 ;
        RECT 41.225 135.225 41.940 135.395 ;
        RECT 42.135 135.275 42.455 135.565 ;
        RECT 42.630 135.275 42.970 136.245 ;
        RECT 43.140 135.275 43.310 136.415 ;
        RECT 43.580 135.615 43.830 136.415 ;
        RECT 44.475 135.445 44.805 136.245 ;
        RECT 45.105 135.615 45.435 136.415 ;
        RECT 45.605 135.445 45.935 136.245 ;
        RECT 43.500 135.275 45.935 135.445 ;
        RECT 46.310 135.275 46.650 136.245 ;
        RECT 46.820 135.275 46.990 136.415 ;
        RECT 47.260 135.615 47.510 136.415 ;
        RECT 48.155 135.445 48.485 136.245 ;
        RECT 48.785 135.615 49.115 136.415 ;
        RECT 49.285 135.445 49.615 136.245 ;
        RECT 47.180 135.275 49.615 135.445 ;
        RECT 50.450 135.275 50.790 136.245 ;
        RECT 50.960 135.275 51.130 136.415 ;
        RECT 51.400 135.615 51.650 136.415 ;
        RECT 52.295 135.445 52.625 136.245 ;
        RECT 52.925 135.615 53.255 136.415 ;
        RECT 53.425 135.445 53.755 136.245 ;
        RECT 51.320 135.275 53.755 135.445 ;
        RECT 55.090 135.275 55.320 136.415 ;
        RECT 40.210 134.775 40.480 135.105 ;
        RECT 40.650 134.775 41.055 135.105 ;
        RECT 41.225 134.775 41.935 135.225 ;
        RECT 40.310 134.605 40.480 134.775 ;
        RECT 39.870 134.195 40.140 134.540 ;
        RECT 40.310 134.435 41.920 134.605 ;
        RECT 42.105 134.535 42.455 135.105 ;
        RECT 42.630 134.665 42.805 135.275 ;
        RECT 43.500 135.025 43.670 135.275 ;
        RECT 42.975 134.855 43.670 135.025 ;
        RECT 43.840 134.885 44.265 135.055 ;
        RECT 43.845 134.855 44.265 134.885 ;
        RECT 44.435 134.855 44.765 135.055 ;
        RECT 44.935 134.855 45.265 135.055 ;
        RECT 40.330 133.865 40.710 134.265 ;
        RECT 40.880 134.085 41.050 134.435 ;
        RECT 41.220 133.865 41.550 134.265 ;
        RECT 41.750 134.085 41.920 134.435 ;
        RECT 42.120 133.865 42.450 134.365 ;
        RECT 42.630 134.035 42.970 134.665 ;
        RECT 43.140 133.865 43.390 134.665 ;
        RECT 43.580 134.515 44.805 134.685 ;
        RECT 43.580 134.035 43.910 134.515 ;
        RECT 44.080 133.865 44.305 134.325 ;
        RECT 44.475 134.035 44.805 134.515 ;
        RECT 45.435 134.645 45.605 135.275 ;
        RECT 45.790 134.855 46.140 135.105 ;
        RECT 46.310 134.665 46.485 135.275 ;
        RECT 47.180 135.025 47.350 135.275 ;
        RECT 46.655 134.855 47.350 135.025 ;
        RECT 47.525 134.855 47.945 135.055 ;
        RECT 48.115 134.855 48.445 135.055 ;
        RECT 48.615 134.855 48.945 135.055 ;
        RECT 45.435 134.035 45.935 134.645 ;
        RECT 46.310 134.035 46.650 134.665 ;
        RECT 46.820 133.865 47.070 134.665 ;
        RECT 47.260 134.515 48.485 134.685 ;
        RECT 47.260 134.035 47.590 134.515 ;
        RECT 47.760 133.865 47.985 134.325 ;
        RECT 48.155 134.035 48.485 134.515 ;
        RECT 49.115 134.645 49.285 135.275 ;
        RECT 49.470 134.855 49.820 135.105 ;
        RECT 50.450 134.665 50.625 135.275 ;
        RECT 51.320 135.025 51.490 135.275 ;
        RECT 50.795 134.855 51.490 135.025 ;
        RECT 51.665 134.855 52.085 135.055 ;
        RECT 52.255 134.855 52.585 135.055 ;
        RECT 52.755 134.855 53.085 135.055 ;
        RECT 49.115 134.035 49.615 134.645 ;
        RECT 50.450 134.035 50.790 134.665 ;
        RECT 50.960 133.865 51.210 134.665 ;
        RECT 51.400 134.515 52.625 134.685 ;
        RECT 51.400 134.035 51.730 134.515 ;
        RECT 51.900 133.865 52.125 134.325 ;
        RECT 52.295 134.035 52.625 134.515 ;
        RECT 53.255 134.645 53.425 135.275 ;
        RECT 55.490 135.265 55.820 136.245 ;
        RECT 55.990 135.275 56.200 136.415 ;
        RECT 56.430 135.655 56.945 136.065 ;
        RECT 57.180 135.655 57.350 136.415 ;
        RECT 57.520 136.075 59.550 136.245 ;
        RECT 53.610 134.855 53.960 135.105 ;
        RECT 55.070 134.855 55.400 135.105 ;
        RECT 53.255 134.035 53.755 134.645 ;
        RECT 55.090 133.865 55.320 134.685 ;
        RECT 55.570 134.665 55.820 135.265 ;
        RECT 56.430 134.845 56.770 135.655 ;
        RECT 57.520 135.410 57.690 136.075 ;
        RECT 58.085 135.735 59.210 135.905 ;
        RECT 56.940 135.220 57.690 135.410 ;
        RECT 57.860 135.395 58.870 135.565 ;
        RECT 55.490 134.035 55.820 134.665 ;
        RECT 55.990 133.865 56.200 134.685 ;
        RECT 56.430 134.675 57.660 134.845 ;
        RECT 56.705 134.070 56.950 134.675 ;
        RECT 57.170 133.865 57.680 134.400 ;
        RECT 57.860 134.035 58.050 135.395 ;
        RECT 58.220 135.055 58.495 135.195 ;
        RECT 58.220 134.885 58.500 135.055 ;
        RECT 58.220 134.035 58.495 134.885 ;
        RECT 58.700 134.595 58.870 135.395 ;
        RECT 59.040 134.605 59.210 135.735 ;
        RECT 59.380 135.105 59.550 136.075 ;
        RECT 59.720 135.275 59.890 136.415 ;
        RECT 60.060 135.275 60.395 136.245 ;
        RECT 59.380 134.775 59.575 135.105 ;
        RECT 59.800 134.775 60.055 135.105 ;
        RECT 59.800 134.605 59.970 134.775 ;
        RECT 60.225 134.605 60.395 135.275 ;
        RECT 60.570 135.250 60.860 136.415 ;
        RECT 61.950 135.340 62.220 136.245 ;
        RECT 62.390 135.655 62.720 136.415 ;
        RECT 62.900 135.485 63.070 136.245 ;
        RECT 59.040 134.435 59.970 134.605 ;
        RECT 59.040 134.400 59.215 134.435 ;
        RECT 58.685 134.035 59.215 134.400 ;
        RECT 59.640 133.865 59.970 134.265 ;
        RECT 60.140 134.035 60.395 134.605 ;
        RECT 60.570 133.865 60.860 134.590 ;
        RECT 61.950 134.540 62.120 135.340 ;
        RECT 62.405 135.315 63.070 135.485 ;
        RECT 62.405 135.170 62.575 135.315 ;
        RECT 63.390 135.275 63.600 136.415 ;
        RECT 62.290 134.840 62.575 135.170 ;
        RECT 63.770 135.265 64.100 136.245 ;
        RECT 64.270 135.275 64.500 136.415 ;
        RECT 64.800 135.485 64.970 136.245 ;
        RECT 65.150 135.655 65.480 136.415 ;
        RECT 64.800 135.315 65.465 135.485 ;
        RECT 65.650 135.340 65.920 136.245 ;
        RECT 62.405 134.585 62.575 134.840 ;
        RECT 62.810 134.765 63.140 135.135 ;
        RECT 61.950 134.035 62.210 134.540 ;
        RECT 62.405 134.415 63.070 134.585 ;
        RECT 62.390 133.865 62.720 134.245 ;
        RECT 62.900 134.035 63.070 134.415 ;
        RECT 63.390 133.865 63.600 134.685 ;
        RECT 63.770 134.665 64.020 135.265 ;
        RECT 65.295 135.170 65.465 135.315 ;
        RECT 64.190 134.855 64.520 135.105 ;
        RECT 64.730 134.765 65.060 135.135 ;
        RECT 65.295 134.840 65.580 135.170 ;
        RECT 63.770 134.035 64.100 134.665 ;
        RECT 64.270 133.865 64.500 134.685 ;
        RECT 65.295 134.585 65.465 134.840 ;
        RECT 64.800 134.415 65.465 134.585 ;
        RECT 65.750 134.540 65.920 135.340 ;
        RECT 66.640 135.485 66.810 136.245 ;
        RECT 66.990 135.655 67.320 136.415 ;
        RECT 66.640 135.315 67.305 135.485 ;
        RECT 67.490 135.340 67.760 136.245 ;
        RECT 67.135 135.170 67.305 135.315 ;
        RECT 66.570 134.765 66.900 135.135 ;
        RECT 67.135 134.840 67.420 135.170 ;
        RECT 67.135 134.585 67.305 134.840 ;
        RECT 64.800 134.035 64.970 134.415 ;
        RECT 65.150 133.865 65.480 134.245 ;
        RECT 65.660 134.035 65.920 134.540 ;
        RECT 66.640 134.415 67.305 134.585 ;
        RECT 67.590 134.540 67.760 135.340 ;
        RECT 67.930 135.325 71.440 136.415 ;
        RECT 67.930 134.805 69.620 135.325 ;
        RECT 71.610 135.275 71.880 136.245 ;
        RECT 72.090 135.615 72.370 136.415 ;
        RECT 72.540 135.905 74.195 136.195 ;
        RECT 72.605 135.565 74.195 135.735 ;
        RECT 72.605 135.445 72.775 135.565 ;
        RECT 72.050 135.275 72.775 135.445 ;
        RECT 69.790 134.635 71.440 135.155 ;
        RECT 66.640 134.035 66.810 134.415 ;
        RECT 66.990 133.865 67.320 134.245 ;
        RECT 67.500 134.035 67.760 134.540 ;
        RECT 67.930 133.865 71.440 134.635 ;
        RECT 71.610 134.540 71.780 135.275 ;
        RECT 72.050 135.105 72.220 135.275 ;
        RECT 72.965 135.225 73.680 135.395 ;
        RECT 73.875 135.275 74.195 135.565 ;
        RECT 74.370 135.275 74.710 136.245 ;
        RECT 74.880 135.275 75.050 136.415 ;
        RECT 75.320 135.615 75.570 136.415 ;
        RECT 76.215 135.445 76.545 136.245 ;
        RECT 76.845 135.615 77.175 136.415 ;
        RECT 77.345 135.445 77.675 136.245 ;
        RECT 75.240 135.275 77.675 135.445 ;
        RECT 78.510 135.325 80.180 136.415 ;
        RECT 80.350 135.655 80.865 136.065 ;
        RECT 81.100 135.655 81.270 136.415 ;
        RECT 81.440 136.075 83.470 136.245 ;
        RECT 71.950 134.775 72.220 135.105 ;
        RECT 72.390 134.775 72.795 135.105 ;
        RECT 72.965 134.775 73.675 135.225 ;
        RECT 72.050 134.605 72.220 134.775 ;
        RECT 71.610 134.195 71.880 134.540 ;
        RECT 72.050 134.435 73.660 134.605 ;
        RECT 73.845 134.535 74.195 135.105 ;
        RECT 74.370 134.715 74.545 135.275 ;
        RECT 75.240 135.025 75.410 135.275 ;
        RECT 74.715 134.855 75.410 135.025 ;
        RECT 75.585 134.855 76.005 135.055 ;
        RECT 76.175 134.855 76.505 135.055 ;
        RECT 76.675 134.855 77.005 135.055 ;
        RECT 74.370 134.665 74.600 134.715 ;
        RECT 72.070 133.865 72.450 134.265 ;
        RECT 72.620 134.085 72.790 134.435 ;
        RECT 72.960 133.865 73.290 134.265 ;
        RECT 73.490 134.085 73.660 134.435 ;
        RECT 73.860 133.865 74.190 134.365 ;
        RECT 74.370 134.035 74.710 134.665 ;
        RECT 74.880 133.865 75.130 134.665 ;
        RECT 75.320 134.515 76.545 134.685 ;
        RECT 75.320 134.035 75.650 134.515 ;
        RECT 75.820 133.865 76.045 134.325 ;
        RECT 76.215 134.035 76.545 134.515 ;
        RECT 77.175 134.645 77.345 135.275 ;
        RECT 77.530 134.855 77.880 135.105 ;
        RECT 78.510 134.805 79.260 135.325 ;
        RECT 77.175 134.035 77.675 134.645 ;
        RECT 79.430 134.635 80.180 135.155 ;
        RECT 80.350 134.845 80.690 135.655 ;
        RECT 81.440 135.410 81.610 136.075 ;
        RECT 82.005 135.735 83.130 135.905 ;
        RECT 80.860 135.220 81.610 135.410 ;
        RECT 81.780 135.395 82.790 135.565 ;
        RECT 80.350 134.675 81.580 134.845 ;
        RECT 78.510 133.865 80.180 134.635 ;
        RECT 80.625 134.070 80.870 134.675 ;
        RECT 81.090 133.865 81.600 134.400 ;
        RECT 81.780 134.035 81.970 135.395 ;
        RECT 82.140 134.715 82.415 135.195 ;
        RECT 82.140 134.545 82.420 134.715 ;
        RECT 82.620 134.595 82.790 135.395 ;
        RECT 82.960 134.605 83.130 135.735 ;
        RECT 83.300 135.105 83.470 136.075 ;
        RECT 83.640 135.275 83.810 136.415 ;
        RECT 83.980 135.275 84.315 136.245 ;
        RECT 85.040 135.485 85.210 136.245 ;
        RECT 85.390 135.655 85.720 136.415 ;
        RECT 85.040 135.315 85.705 135.485 ;
        RECT 85.890 135.340 86.160 136.245 ;
        RECT 83.300 134.775 83.495 135.105 ;
        RECT 83.720 134.775 83.975 135.105 ;
        RECT 83.720 134.605 83.890 134.775 ;
        RECT 84.145 134.605 84.315 135.275 ;
        RECT 85.535 135.170 85.705 135.315 ;
        RECT 84.970 134.765 85.300 135.135 ;
        RECT 85.535 134.840 85.820 135.170 ;
        RECT 82.140 134.035 82.415 134.545 ;
        RECT 82.960 134.435 83.890 134.605 ;
        RECT 82.960 134.400 83.135 134.435 ;
        RECT 82.605 134.035 83.135 134.400 ;
        RECT 83.560 133.865 83.890 134.265 ;
        RECT 84.060 134.035 84.315 134.605 ;
        RECT 85.535 134.585 85.705 134.840 ;
        RECT 85.040 134.415 85.705 134.585 ;
        RECT 85.990 134.540 86.160 135.340 ;
        RECT 86.330 135.250 86.620 136.415 ;
        RECT 87.250 135.325 89.840 136.415 ;
        RECT 87.250 134.805 88.460 135.325 ;
        RECT 90.050 135.275 90.280 136.415 ;
        RECT 90.450 135.265 90.780 136.245 ;
        RECT 90.950 135.275 91.160 136.415 ;
        RECT 91.390 135.655 91.905 136.065 ;
        RECT 92.140 135.655 92.310 136.415 ;
        RECT 92.480 136.075 94.510 136.245 ;
        RECT 88.630 134.635 89.840 135.155 ;
        RECT 90.030 134.855 90.360 135.105 ;
        RECT 85.040 134.035 85.210 134.415 ;
        RECT 85.390 133.865 85.720 134.245 ;
        RECT 85.900 134.035 86.160 134.540 ;
        RECT 86.330 133.865 86.620 134.590 ;
        RECT 87.250 133.865 89.840 134.635 ;
        RECT 90.050 133.865 90.280 134.685 ;
        RECT 90.530 134.665 90.780 135.265 ;
        RECT 91.390 134.845 91.730 135.655 ;
        RECT 92.480 135.410 92.650 136.075 ;
        RECT 93.045 135.735 94.170 135.905 ;
        RECT 91.900 135.220 92.650 135.410 ;
        RECT 92.820 135.395 93.830 135.565 ;
        RECT 90.450 134.035 90.780 134.665 ;
        RECT 90.950 133.865 91.160 134.685 ;
        RECT 91.390 134.675 92.620 134.845 ;
        RECT 91.665 134.070 91.910 134.675 ;
        RECT 92.130 133.865 92.640 134.400 ;
        RECT 92.820 134.035 93.010 135.395 ;
        RECT 93.180 135.055 93.455 135.195 ;
        RECT 93.180 134.885 93.460 135.055 ;
        RECT 93.180 134.035 93.455 134.885 ;
        RECT 93.660 134.595 93.830 135.395 ;
        RECT 94.000 134.605 94.170 135.735 ;
        RECT 94.340 135.105 94.510 136.075 ;
        RECT 94.680 135.275 94.850 136.415 ;
        RECT 95.020 135.275 95.355 136.245 ;
        RECT 94.340 134.775 94.535 135.105 ;
        RECT 94.760 134.775 95.015 135.105 ;
        RECT 94.760 134.605 94.930 134.775 ;
        RECT 95.185 134.605 95.355 135.275 ;
        RECT 95.990 135.655 96.505 136.065 ;
        RECT 96.740 135.655 96.910 136.415 ;
        RECT 97.080 136.075 99.110 136.245 ;
        RECT 95.990 134.845 96.330 135.655 ;
        RECT 97.080 135.410 97.250 136.075 ;
        RECT 97.645 135.735 98.770 135.905 ;
        RECT 96.500 135.220 97.250 135.410 ;
        RECT 97.420 135.395 98.430 135.565 ;
        RECT 95.990 134.675 97.220 134.845 ;
        RECT 94.000 134.435 94.930 134.605 ;
        RECT 94.000 134.400 94.175 134.435 ;
        RECT 93.645 134.035 94.175 134.400 ;
        RECT 94.600 133.865 94.930 134.265 ;
        RECT 95.100 134.035 95.355 134.605 ;
        RECT 96.265 134.070 96.510 134.675 ;
        RECT 96.730 133.865 97.240 134.400 ;
        RECT 97.420 134.035 97.610 135.395 ;
        RECT 97.780 135.055 98.055 135.195 ;
        RECT 97.780 134.885 98.060 135.055 ;
        RECT 97.780 134.035 98.055 134.885 ;
        RECT 98.260 134.595 98.430 135.395 ;
        RECT 98.600 134.605 98.770 135.735 ;
        RECT 98.940 135.105 99.110 136.075 ;
        RECT 99.280 135.275 99.450 136.415 ;
        RECT 99.620 135.275 99.955 136.245 ;
        RECT 101.425 135.435 101.680 136.105 ;
        RECT 101.860 135.615 102.145 136.415 ;
        RECT 102.325 135.695 102.655 136.205 ;
        RECT 101.425 135.395 101.605 135.435 ;
        RECT 98.940 134.775 99.135 135.105 ;
        RECT 99.360 134.775 99.615 135.105 ;
        RECT 99.360 134.605 99.530 134.775 ;
        RECT 99.785 134.605 99.955 135.275 ;
        RECT 101.340 135.225 101.605 135.395 ;
        RECT 98.600 134.435 99.530 134.605 ;
        RECT 98.600 134.400 98.775 134.435 ;
        RECT 98.245 134.035 98.775 134.400 ;
        RECT 99.200 133.865 99.530 134.265 ;
        RECT 99.700 134.035 99.955 134.605 ;
        RECT 101.425 134.575 101.605 135.225 ;
        RECT 102.325 135.105 102.575 135.695 ;
        RECT 102.925 135.545 103.095 136.155 ;
        RECT 103.265 135.725 103.595 136.415 ;
        RECT 103.825 135.865 104.065 136.155 ;
        RECT 104.265 136.035 104.685 136.415 ;
        RECT 104.865 135.945 105.495 136.195 ;
        RECT 105.965 136.035 106.295 136.415 ;
        RECT 104.865 135.865 105.035 135.945 ;
        RECT 106.465 135.865 106.635 136.155 ;
        RECT 106.815 136.035 107.195 136.415 ;
        RECT 107.435 136.030 108.265 136.200 ;
        RECT 103.825 135.695 105.035 135.865 ;
        RECT 101.775 134.775 102.575 135.105 ;
        RECT 101.425 134.045 101.680 134.575 ;
        RECT 101.860 133.865 102.145 134.325 ;
        RECT 102.325 134.125 102.575 134.775 ;
        RECT 102.775 135.525 103.095 135.545 ;
        RECT 102.775 135.355 104.695 135.525 ;
        RECT 102.775 134.460 102.965 135.355 ;
        RECT 104.865 135.185 105.035 135.695 ;
        RECT 105.205 135.435 105.725 135.745 ;
        RECT 103.135 135.015 105.035 135.185 ;
        RECT 103.135 134.955 103.465 135.015 ;
        RECT 103.615 134.785 103.945 134.845 ;
        RECT 103.285 134.515 103.945 134.785 ;
        RECT 102.775 134.130 103.095 134.460 ;
        RECT 103.275 133.865 103.935 134.345 ;
        RECT 104.135 134.255 104.305 135.015 ;
        RECT 105.205 134.845 105.385 135.255 ;
        RECT 104.475 134.675 104.805 134.795 ;
        RECT 105.555 134.675 105.725 135.435 ;
        RECT 104.475 134.505 105.725 134.675 ;
        RECT 105.895 135.615 107.265 135.865 ;
        RECT 105.895 134.845 106.085 135.615 ;
        RECT 107.015 135.355 107.265 135.615 ;
        RECT 106.255 135.185 106.505 135.345 ;
        RECT 107.435 135.185 107.605 136.030 ;
        RECT 108.500 135.745 108.670 136.245 ;
        RECT 108.840 135.915 109.170 136.415 ;
        RECT 107.775 135.355 108.275 135.735 ;
        RECT 108.500 135.575 109.195 135.745 ;
        RECT 106.255 135.015 107.605 135.185 ;
        RECT 107.185 134.975 107.605 135.015 ;
        RECT 105.895 134.505 106.315 134.845 ;
        RECT 106.605 134.515 107.015 134.845 ;
        RECT 104.135 134.085 104.985 134.255 ;
        RECT 105.545 133.865 105.865 134.325 ;
        RECT 106.065 134.075 106.315 134.505 ;
        RECT 106.605 133.865 107.015 134.305 ;
        RECT 107.185 134.245 107.355 134.975 ;
        RECT 107.525 134.425 107.875 134.795 ;
        RECT 108.055 134.485 108.275 135.355 ;
        RECT 108.445 134.785 108.855 135.405 ;
        RECT 109.025 134.605 109.195 135.575 ;
        RECT 108.500 134.415 109.195 134.605 ;
        RECT 107.185 134.045 108.200 134.245 ;
        RECT 108.500 134.085 108.670 134.415 ;
        RECT 108.840 133.865 109.170 134.245 ;
        RECT 109.385 134.125 109.610 136.245 ;
        RECT 109.780 135.915 110.110 136.415 ;
        RECT 110.280 135.745 110.450 136.245 ;
        RECT 109.785 135.575 110.450 135.745 ;
        RECT 109.785 134.585 110.015 135.575 ;
        RECT 110.185 134.755 110.535 135.405 ;
        RECT 111.170 135.325 112.380 136.415 ;
        RECT 111.170 134.785 111.690 135.325 ;
        RECT 111.860 134.615 112.380 135.155 ;
        RECT 109.785 134.415 110.450 134.585 ;
        RECT 109.780 133.865 110.110 134.245 ;
        RECT 110.280 134.125 110.450 134.415 ;
        RECT 111.170 133.865 112.380 134.615 ;
        RECT 18.165 133.695 112.465 133.865 ;
        RECT 18.250 132.945 19.460 133.695 ;
        RECT 18.250 132.405 18.770 132.945 ;
        RECT 20.090 132.925 21.760 133.695 ;
        RECT 21.930 132.970 22.220 133.695 ;
        RECT 18.940 132.235 19.460 132.775 ;
        RECT 18.250 131.145 19.460 132.235 ;
        RECT 20.090 132.235 20.840 132.755 ;
        RECT 21.010 132.405 21.760 132.925 ;
        RECT 22.890 132.875 23.120 133.695 ;
        RECT 23.290 132.895 23.620 133.525 ;
        RECT 22.870 132.455 23.200 132.705 ;
        RECT 20.090 131.145 21.760 132.235 ;
        RECT 21.930 131.145 22.220 132.310 ;
        RECT 23.370 132.295 23.620 132.895 ;
        RECT 23.790 132.875 24.000 133.695 ;
        RECT 24.320 133.145 24.490 133.525 ;
        RECT 24.670 133.315 25.000 133.695 ;
        RECT 24.320 132.975 24.985 133.145 ;
        RECT 25.180 133.020 25.440 133.525 ;
        RECT 24.250 132.425 24.580 132.795 ;
        RECT 24.815 132.720 24.985 132.975 ;
        RECT 22.890 131.145 23.120 132.285 ;
        RECT 23.290 131.315 23.620 132.295 ;
        RECT 24.815 132.390 25.100 132.720 ;
        RECT 23.790 131.145 24.000 132.285 ;
        RECT 24.815 132.245 24.985 132.390 ;
        RECT 24.320 132.075 24.985 132.245 ;
        RECT 25.270 132.220 25.440 133.020 ;
        RECT 24.320 131.315 24.490 132.075 ;
        RECT 24.670 131.145 25.000 131.905 ;
        RECT 25.170 131.315 25.440 132.220 ;
        RECT 25.615 132.985 25.870 133.515 ;
        RECT 26.040 133.235 26.345 133.695 ;
        RECT 26.590 133.315 27.660 133.485 ;
        RECT 25.615 132.335 25.825 132.985 ;
        RECT 26.590 132.960 26.910 133.315 ;
        RECT 26.585 132.785 26.910 132.960 ;
        RECT 25.995 132.485 26.910 132.785 ;
        RECT 27.080 132.745 27.320 133.145 ;
        RECT 27.490 133.085 27.660 133.315 ;
        RECT 27.830 133.255 28.020 133.695 ;
        RECT 28.190 133.245 29.140 133.525 ;
        RECT 29.360 133.335 29.710 133.505 ;
        RECT 27.490 132.915 28.020 133.085 ;
        RECT 25.995 132.455 26.735 132.485 ;
        RECT 25.615 131.455 25.870 132.335 ;
        RECT 26.040 131.145 26.345 132.285 ;
        RECT 26.565 131.865 26.735 132.455 ;
        RECT 27.080 132.375 27.620 132.745 ;
        RECT 27.800 132.635 28.020 132.915 ;
        RECT 28.190 132.465 28.360 133.245 ;
        RECT 27.955 132.295 28.360 132.465 ;
        RECT 28.530 132.455 28.880 133.075 ;
        RECT 27.955 132.205 28.125 132.295 ;
        RECT 29.050 132.285 29.260 133.075 ;
        RECT 26.905 132.035 28.125 132.205 ;
        RECT 28.585 132.125 29.260 132.285 ;
        RECT 26.565 131.695 27.365 131.865 ;
        RECT 26.685 131.145 27.015 131.525 ;
        RECT 27.195 131.405 27.365 131.695 ;
        RECT 27.955 131.655 28.125 132.035 ;
        RECT 28.295 132.115 29.260 132.125 ;
        RECT 29.450 132.945 29.710 133.335 ;
        RECT 29.920 133.235 30.250 133.695 ;
        RECT 31.125 133.305 31.980 133.475 ;
        RECT 32.185 133.305 32.680 133.475 ;
        RECT 32.850 133.335 33.180 133.695 ;
        RECT 29.450 132.255 29.620 132.945 ;
        RECT 29.790 132.595 29.960 132.775 ;
        RECT 30.130 132.765 30.920 133.015 ;
        RECT 31.125 132.595 31.295 133.305 ;
        RECT 31.465 132.795 31.820 133.015 ;
        RECT 29.790 132.425 31.480 132.595 ;
        RECT 28.295 131.825 28.755 132.115 ;
        RECT 29.450 132.085 30.950 132.255 ;
        RECT 29.450 131.945 29.620 132.085 ;
        RECT 29.060 131.775 29.620 131.945 ;
        RECT 27.535 131.145 27.785 131.605 ;
        RECT 27.955 131.315 28.825 131.655 ;
        RECT 29.060 131.315 29.230 131.775 ;
        RECT 30.065 131.745 31.140 131.915 ;
        RECT 29.400 131.145 29.770 131.605 ;
        RECT 30.065 131.405 30.235 131.745 ;
        RECT 30.405 131.145 30.735 131.575 ;
        RECT 30.970 131.405 31.140 131.745 ;
        RECT 31.310 131.645 31.480 132.425 ;
        RECT 31.650 132.205 31.820 132.795 ;
        RECT 31.990 132.395 32.340 133.015 ;
        RECT 31.650 131.815 32.115 132.205 ;
        RECT 32.510 131.945 32.680 133.305 ;
        RECT 32.850 132.115 33.310 133.165 ;
        RECT 32.285 131.775 32.680 131.945 ;
        RECT 32.285 131.645 32.455 131.775 ;
        RECT 31.310 131.315 31.990 131.645 ;
        RECT 32.205 131.315 32.455 131.645 ;
        RECT 32.625 131.145 32.875 131.605 ;
        RECT 33.045 131.330 33.370 132.115 ;
        RECT 33.540 131.315 33.710 133.435 ;
        RECT 33.880 133.315 34.210 133.695 ;
        RECT 34.380 133.145 34.635 133.435 ;
        RECT 33.885 132.975 34.635 133.145 ;
        RECT 34.810 133.020 35.070 133.525 ;
        RECT 35.250 133.315 35.580 133.695 ;
        RECT 35.760 133.145 35.930 133.525 ;
        RECT 33.885 131.985 34.115 132.975 ;
        RECT 34.285 132.155 34.635 132.805 ;
        RECT 34.810 132.220 34.980 133.020 ;
        RECT 35.265 132.975 35.930 133.145 ;
        RECT 35.265 132.720 35.435 132.975 ;
        RECT 36.190 132.925 37.860 133.695 ;
        RECT 35.150 132.390 35.435 132.720 ;
        RECT 35.670 132.425 36.000 132.795 ;
        RECT 35.265 132.245 35.435 132.390 ;
        RECT 33.885 131.815 34.635 131.985 ;
        RECT 33.880 131.145 34.210 131.645 ;
        RECT 34.380 131.315 34.635 131.815 ;
        RECT 34.810 131.315 35.080 132.220 ;
        RECT 35.265 132.075 35.930 132.245 ;
        RECT 35.250 131.145 35.580 131.905 ;
        RECT 35.760 131.315 35.930 132.075 ;
        RECT 36.190 132.235 36.940 132.755 ;
        RECT 37.110 132.405 37.860 132.925 ;
        RECT 38.230 133.065 38.560 133.425 ;
        RECT 39.180 133.235 39.430 133.695 ;
        RECT 39.600 133.235 40.160 133.525 ;
        RECT 38.230 132.875 39.620 133.065 ;
        RECT 39.450 132.785 39.620 132.875 ;
        RECT 38.045 132.455 38.720 132.705 ;
        RECT 38.940 132.455 39.280 132.705 ;
        RECT 39.450 132.455 39.740 132.785 ;
        RECT 36.190 131.145 37.860 132.235 ;
        RECT 38.045 132.095 38.310 132.455 ;
        RECT 39.450 132.205 39.620 132.455 ;
        RECT 38.680 132.035 39.620 132.205 ;
        RECT 38.230 131.145 38.510 131.815 ;
        RECT 38.680 131.485 38.980 132.035 ;
        RECT 39.910 131.865 40.160 133.235 ;
        RECT 40.340 133.195 40.670 133.695 ;
        RECT 40.870 133.125 41.040 133.475 ;
        RECT 41.240 133.295 41.570 133.695 ;
        RECT 41.740 133.125 41.910 133.475 ;
        RECT 42.080 133.295 42.460 133.695 ;
        RECT 40.335 132.455 40.685 133.025 ;
        RECT 40.870 132.955 42.480 133.125 ;
        RECT 42.650 133.020 42.920 133.365 ;
        RECT 42.310 132.785 42.480 132.955 ;
        RECT 39.180 131.145 39.510 131.865 ;
        RECT 39.700 131.315 40.160 131.865 ;
        RECT 40.335 131.995 40.655 132.285 ;
        RECT 40.855 132.165 41.565 132.785 ;
        RECT 41.735 132.455 42.140 132.785 ;
        RECT 42.310 132.455 42.580 132.785 ;
        RECT 42.310 132.285 42.480 132.455 ;
        RECT 42.750 132.285 42.920 133.020 ;
        RECT 41.755 132.115 42.480 132.285 ;
        RECT 41.755 131.995 41.925 132.115 ;
        RECT 40.335 131.825 41.925 131.995 ;
        RECT 40.335 131.365 41.990 131.655 ;
        RECT 42.160 131.145 42.440 131.945 ;
        RECT 42.650 131.315 42.920 132.285 ;
        RECT 43.090 132.895 43.430 133.525 ;
        RECT 43.600 132.895 43.850 133.695 ;
        RECT 44.040 133.045 44.370 133.525 ;
        RECT 44.540 133.235 44.765 133.695 ;
        RECT 44.935 133.045 45.265 133.525 ;
        RECT 43.090 132.285 43.265 132.895 ;
        RECT 44.040 132.875 45.265 133.045 ;
        RECT 45.895 132.915 46.395 133.525 ;
        RECT 47.690 132.970 47.980 133.695 ;
        RECT 48.150 132.925 51.660 133.695 ;
        RECT 43.435 132.535 44.130 132.705 ;
        RECT 43.960 132.285 44.130 132.535 ;
        RECT 44.305 132.505 44.725 132.705 ;
        RECT 44.895 132.505 45.225 132.705 ;
        RECT 45.395 132.505 45.725 132.705 ;
        RECT 45.895 132.285 46.065 132.915 ;
        RECT 46.250 132.455 46.600 132.705 ;
        RECT 43.090 131.315 43.430 132.285 ;
        RECT 43.600 131.145 43.770 132.285 ;
        RECT 43.960 132.115 46.395 132.285 ;
        RECT 44.040 131.145 44.290 131.945 ;
        RECT 44.935 131.315 45.265 132.115 ;
        RECT 45.565 131.145 45.895 131.945 ;
        RECT 46.065 131.315 46.395 132.115 ;
        RECT 47.690 131.145 47.980 132.310 ;
        RECT 48.150 132.235 49.840 132.755 ;
        RECT 50.010 132.405 51.660 132.925 ;
        RECT 51.830 132.895 52.170 133.525 ;
        RECT 52.340 132.895 52.590 133.695 ;
        RECT 52.780 133.045 53.110 133.525 ;
        RECT 53.280 133.235 53.505 133.695 ;
        RECT 53.675 133.045 54.005 133.525 ;
        RECT 51.830 132.285 52.005 132.895 ;
        RECT 52.780 132.875 54.005 133.045 ;
        RECT 54.635 132.915 55.135 133.525 ;
        RECT 52.175 132.535 52.870 132.705 ;
        RECT 52.700 132.285 52.870 132.535 ;
        RECT 53.045 132.505 53.465 132.705 ;
        RECT 53.635 132.505 53.965 132.705 ;
        RECT 54.135 132.505 54.465 132.705 ;
        RECT 54.635 132.285 54.805 132.915 ;
        RECT 55.785 132.885 56.030 133.490 ;
        RECT 56.250 133.160 56.760 133.695 ;
        RECT 55.510 132.715 56.740 132.885 ;
        RECT 54.990 132.455 55.340 132.705 ;
        RECT 48.150 131.145 51.660 132.235 ;
        RECT 51.830 131.315 52.170 132.285 ;
        RECT 52.340 131.145 52.510 132.285 ;
        RECT 52.700 132.115 55.135 132.285 ;
        RECT 52.780 131.145 53.030 131.945 ;
        RECT 53.675 131.315 54.005 132.115 ;
        RECT 54.305 131.145 54.635 131.945 ;
        RECT 54.805 131.315 55.135 132.115 ;
        RECT 55.510 131.905 55.850 132.715 ;
        RECT 56.020 132.150 56.770 132.340 ;
        RECT 55.510 131.495 56.025 131.905 ;
        RECT 56.260 131.145 56.430 131.905 ;
        RECT 56.600 131.485 56.770 132.150 ;
        RECT 56.940 132.165 57.130 133.525 ;
        RECT 57.300 133.355 57.575 133.525 ;
        RECT 57.300 133.185 57.580 133.355 ;
        RECT 57.300 132.365 57.575 133.185 ;
        RECT 57.765 133.160 58.295 133.525 ;
        RECT 58.720 133.295 59.050 133.695 ;
        RECT 58.120 133.125 58.295 133.160 ;
        RECT 57.780 132.165 57.950 132.965 ;
        RECT 56.940 131.995 57.950 132.165 ;
        RECT 58.120 132.955 59.050 133.125 ;
        RECT 59.220 132.955 59.475 133.525 ;
        RECT 58.120 131.825 58.290 132.955 ;
        RECT 58.880 132.785 59.050 132.955 ;
        RECT 57.165 131.655 58.290 131.825 ;
        RECT 58.460 132.455 58.655 132.785 ;
        RECT 58.880 132.455 59.135 132.785 ;
        RECT 58.460 131.485 58.630 132.455 ;
        RECT 59.305 132.285 59.475 132.955 ;
        RECT 56.600 131.315 58.630 131.485 ;
        RECT 58.800 131.145 58.970 132.285 ;
        RECT 59.140 131.315 59.475 132.285 ;
        RECT 60.025 132.985 60.280 133.515 ;
        RECT 60.460 133.235 60.745 133.695 ;
        RECT 60.025 132.125 60.205 132.985 ;
        RECT 60.925 132.785 61.175 133.435 ;
        RECT 60.375 132.455 61.175 132.785 ;
        RECT 60.025 131.655 60.280 132.125 ;
        RECT 59.940 131.485 60.280 131.655 ;
        RECT 60.025 131.455 60.280 131.485 ;
        RECT 60.460 131.145 60.745 131.945 ;
        RECT 60.925 131.865 61.175 132.455 ;
        RECT 61.375 133.100 61.695 133.430 ;
        RECT 61.875 133.215 62.535 133.695 ;
        RECT 62.735 133.305 63.585 133.475 ;
        RECT 61.375 132.205 61.565 133.100 ;
        RECT 61.885 132.775 62.545 133.045 ;
        RECT 62.215 132.715 62.545 132.775 ;
        RECT 61.735 132.545 62.065 132.605 ;
        RECT 62.735 132.545 62.905 133.305 ;
        RECT 64.145 133.235 64.465 133.695 ;
        RECT 64.665 133.055 64.915 133.485 ;
        RECT 65.205 133.255 65.615 133.695 ;
        RECT 65.785 133.315 66.800 133.515 ;
        RECT 63.075 132.885 64.325 133.055 ;
        RECT 63.075 132.765 63.405 132.885 ;
        RECT 61.735 132.375 63.635 132.545 ;
        RECT 61.375 132.035 63.295 132.205 ;
        RECT 61.375 132.015 61.695 132.035 ;
        RECT 60.925 131.355 61.255 131.865 ;
        RECT 61.525 131.405 61.695 132.015 ;
        RECT 63.465 131.865 63.635 132.375 ;
        RECT 63.805 132.305 63.985 132.715 ;
        RECT 64.155 132.125 64.325 132.885 ;
        RECT 61.865 131.145 62.195 131.835 ;
        RECT 62.425 131.695 63.635 131.865 ;
        RECT 63.805 131.815 64.325 132.125 ;
        RECT 64.495 132.715 64.915 133.055 ;
        RECT 65.205 132.715 65.615 133.045 ;
        RECT 64.495 131.945 64.685 132.715 ;
        RECT 65.785 132.585 65.955 133.315 ;
        RECT 67.100 133.145 67.270 133.475 ;
        RECT 67.440 133.315 67.770 133.695 ;
        RECT 66.125 132.765 66.475 133.135 ;
        RECT 65.785 132.545 66.205 132.585 ;
        RECT 64.855 132.375 66.205 132.545 ;
        RECT 64.855 132.215 65.105 132.375 ;
        RECT 65.615 131.945 65.865 132.205 ;
        RECT 64.495 131.695 65.865 131.945 ;
        RECT 62.425 131.405 62.665 131.695 ;
        RECT 63.465 131.615 63.635 131.695 ;
        RECT 62.865 131.145 63.285 131.525 ;
        RECT 63.465 131.365 64.095 131.615 ;
        RECT 64.565 131.145 64.895 131.525 ;
        RECT 65.065 131.405 65.235 131.695 ;
        RECT 66.035 131.530 66.205 132.375 ;
        RECT 66.655 132.205 66.875 133.075 ;
        RECT 67.100 132.955 67.795 133.145 ;
        RECT 66.375 131.825 66.875 132.205 ;
        RECT 67.045 132.155 67.455 132.775 ;
        RECT 67.625 131.985 67.795 132.955 ;
        RECT 67.100 131.815 67.795 131.985 ;
        RECT 65.415 131.145 65.795 131.525 ;
        RECT 66.035 131.360 66.865 131.530 ;
        RECT 67.100 131.315 67.270 131.815 ;
        RECT 67.440 131.145 67.770 131.645 ;
        RECT 67.985 131.315 68.210 133.435 ;
        RECT 68.380 133.315 68.710 133.695 ;
        RECT 68.880 133.145 69.050 133.435 ;
        RECT 68.385 132.975 69.050 133.145 ;
        RECT 69.310 133.020 69.570 133.525 ;
        RECT 69.750 133.315 70.080 133.695 ;
        RECT 70.260 133.145 70.430 133.525 ;
        RECT 70.700 133.195 71.030 133.695 ;
        RECT 68.385 131.985 68.615 132.975 ;
        RECT 68.785 132.155 69.135 132.805 ;
        RECT 69.310 132.220 69.480 133.020 ;
        RECT 69.765 132.975 70.430 133.145 ;
        RECT 71.230 133.125 71.400 133.475 ;
        RECT 71.600 133.295 71.930 133.695 ;
        RECT 72.100 133.125 72.270 133.475 ;
        RECT 72.440 133.295 72.820 133.695 ;
        RECT 69.765 132.720 69.935 132.975 ;
        RECT 69.650 132.390 69.935 132.720 ;
        RECT 70.170 132.425 70.500 132.795 ;
        RECT 70.695 132.455 71.045 133.025 ;
        RECT 71.230 132.955 72.840 133.125 ;
        RECT 73.010 133.020 73.280 133.365 ;
        RECT 72.670 132.785 72.840 132.955 ;
        RECT 69.765 132.245 69.935 132.390 ;
        RECT 68.385 131.815 69.050 131.985 ;
        RECT 68.380 131.145 68.710 131.645 ;
        RECT 68.880 131.315 69.050 131.815 ;
        RECT 69.310 131.315 69.580 132.220 ;
        RECT 69.765 132.075 70.430 132.245 ;
        RECT 69.750 131.145 70.080 131.905 ;
        RECT 70.260 131.315 70.430 132.075 ;
        RECT 70.695 131.995 71.015 132.285 ;
        RECT 71.215 132.165 71.925 132.785 ;
        RECT 72.095 132.455 72.500 132.785 ;
        RECT 72.670 132.455 72.940 132.785 ;
        RECT 72.670 132.285 72.840 132.455 ;
        RECT 73.110 132.285 73.280 133.020 ;
        RECT 73.450 132.970 73.740 133.695 ;
        RECT 74.370 132.895 74.710 133.525 ;
        RECT 74.880 132.895 75.130 133.695 ;
        RECT 75.320 133.045 75.650 133.525 ;
        RECT 75.820 133.235 76.045 133.695 ;
        RECT 76.215 133.045 76.545 133.525 ;
        RECT 74.370 132.845 74.600 132.895 ;
        RECT 75.320 132.875 76.545 133.045 ;
        RECT 77.175 132.915 77.675 133.525 ;
        RECT 72.115 132.115 72.840 132.285 ;
        RECT 72.115 131.995 72.285 132.115 ;
        RECT 70.695 131.825 72.285 131.995 ;
        RECT 70.695 131.365 72.350 131.655 ;
        RECT 72.520 131.145 72.800 131.945 ;
        RECT 73.010 131.315 73.280 132.285 ;
        RECT 73.450 131.145 73.740 132.310 ;
        RECT 74.370 132.285 74.545 132.845 ;
        RECT 74.715 132.535 75.410 132.705 ;
        RECT 75.240 132.285 75.410 132.535 ;
        RECT 75.585 132.505 76.005 132.705 ;
        RECT 76.175 132.505 76.505 132.705 ;
        RECT 76.675 132.505 77.005 132.705 ;
        RECT 77.175 132.285 77.345 132.915 ;
        RECT 78.110 132.875 78.320 133.695 ;
        RECT 78.490 132.895 78.820 133.525 ;
        RECT 77.530 132.455 77.880 132.705 ;
        RECT 78.490 132.295 78.740 132.895 ;
        RECT 78.990 132.875 79.220 133.695 ;
        RECT 79.805 132.985 80.060 133.515 ;
        RECT 80.240 133.235 80.525 133.695 ;
        RECT 78.910 132.455 79.240 132.705 ;
        RECT 74.370 131.315 74.710 132.285 ;
        RECT 74.880 131.145 75.050 132.285 ;
        RECT 75.240 132.115 77.675 132.285 ;
        RECT 75.320 131.145 75.570 131.945 ;
        RECT 76.215 131.315 76.545 132.115 ;
        RECT 76.845 131.145 77.175 131.945 ;
        RECT 77.345 131.315 77.675 132.115 ;
        RECT 78.110 131.145 78.320 132.285 ;
        RECT 78.490 131.315 78.820 132.295 ;
        RECT 78.990 131.145 79.220 132.285 ;
        RECT 79.805 132.125 79.985 132.985 ;
        RECT 80.705 132.785 80.955 133.435 ;
        RECT 80.155 132.455 80.955 132.785 ;
        RECT 79.805 131.995 80.060 132.125 ;
        RECT 79.720 131.825 80.060 131.995 ;
        RECT 79.805 131.455 80.060 131.825 ;
        RECT 80.240 131.145 80.525 131.945 ;
        RECT 80.705 131.865 80.955 132.455 ;
        RECT 81.155 133.100 81.475 133.430 ;
        RECT 81.655 133.215 82.315 133.695 ;
        RECT 82.515 133.305 83.365 133.475 ;
        RECT 81.155 132.205 81.345 133.100 ;
        RECT 81.665 132.775 82.325 133.045 ;
        RECT 81.995 132.715 82.325 132.775 ;
        RECT 81.515 132.545 81.845 132.605 ;
        RECT 82.515 132.545 82.685 133.305 ;
        RECT 83.925 133.235 84.245 133.695 ;
        RECT 84.445 133.055 84.695 133.485 ;
        RECT 84.985 133.255 85.395 133.695 ;
        RECT 85.565 133.315 86.580 133.515 ;
        RECT 82.855 132.885 84.105 133.055 ;
        RECT 82.855 132.765 83.185 132.885 ;
        RECT 81.515 132.375 83.415 132.545 ;
        RECT 81.155 132.035 83.075 132.205 ;
        RECT 81.155 132.015 81.475 132.035 ;
        RECT 80.705 131.355 81.035 131.865 ;
        RECT 81.305 131.405 81.475 132.015 ;
        RECT 83.245 131.865 83.415 132.375 ;
        RECT 83.585 132.305 83.765 132.715 ;
        RECT 83.935 132.125 84.105 132.885 ;
        RECT 81.645 131.145 81.975 131.835 ;
        RECT 82.205 131.695 83.415 131.865 ;
        RECT 83.585 131.815 84.105 132.125 ;
        RECT 84.275 132.715 84.695 133.055 ;
        RECT 84.985 132.715 85.395 133.045 ;
        RECT 84.275 131.945 84.465 132.715 ;
        RECT 85.565 132.585 85.735 133.315 ;
        RECT 86.880 133.145 87.050 133.475 ;
        RECT 87.220 133.315 87.550 133.695 ;
        RECT 85.905 132.765 86.255 133.135 ;
        RECT 85.565 132.545 85.985 132.585 ;
        RECT 84.635 132.375 85.985 132.545 ;
        RECT 84.635 132.215 84.885 132.375 ;
        RECT 85.395 131.945 85.645 132.205 ;
        RECT 84.275 131.695 85.645 131.945 ;
        RECT 82.205 131.405 82.445 131.695 ;
        RECT 83.245 131.615 83.415 131.695 ;
        RECT 82.645 131.145 83.065 131.525 ;
        RECT 83.245 131.365 83.875 131.615 ;
        RECT 84.345 131.145 84.675 131.525 ;
        RECT 84.845 131.405 85.015 131.695 ;
        RECT 85.815 131.530 85.985 132.375 ;
        RECT 86.435 132.205 86.655 133.075 ;
        RECT 86.880 132.955 87.575 133.145 ;
        RECT 86.155 131.825 86.655 132.205 ;
        RECT 86.825 132.155 87.235 132.775 ;
        RECT 87.405 131.985 87.575 132.955 ;
        RECT 86.880 131.815 87.575 131.985 ;
        RECT 85.195 131.145 85.575 131.525 ;
        RECT 85.815 131.360 86.645 131.530 ;
        RECT 86.880 131.315 87.050 131.815 ;
        RECT 87.220 131.145 87.550 131.645 ;
        RECT 87.765 131.315 87.990 133.435 ;
        RECT 88.160 133.315 88.490 133.695 ;
        RECT 88.660 133.145 88.830 133.435 ;
        RECT 89.925 133.355 90.180 133.515 ;
        RECT 89.840 133.185 90.180 133.355 ;
        RECT 90.360 133.235 90.645 133.695 ;
        RECT 88.165 132.975 88.830 133.145 ;
        RECT 89.925 132.985 90.180 133.185 ;
        RECT 88.165 131.985 88.395 132.975 ;
        RECT 88.565 132.155 88.915 132.805 ;
        RECT 89.925 132.125 90.105 132.985 ;
        RECT 90.825 132.785 91.075 133.435 ;
        RECT 90.275 132.455 91.075 132.785 ;
        RECT 88.165 131.815 88.830 131.985 ;
        RECT 88.160 131.145 88.490 131.645 ;
        RECT 88.660 131.315 88.830 131.815 ;
        RECT 89.925 131.455 90.180 132.125 ;
        RECT 90.360 131.145 90.645 131.945 ;
        RECT 90.825 131.865 91.075 132.455 ;
        RECT 91.275 133.100 91.595 133.430 ;
        RECT 91.775 133.215 92.435 133.695 ;
        RECT 92.635 133.305 93.485 133.475 ;
        RECT 91.275 132.205 91.465 133.100 ;
        RECT 91.785 132.775 92.445 133.045 ;
        RECT 92.115 132.715 92.445 132.775 ;
        RECT 91.635 132.545 91.965 132.605 ;
        RECT 92.635 132.545 92.805 133.305 ;
        RECT 94.045 133.235 94.365 133.695 ;
        RECT 94.565 133.055 94.815 133.485 ;
        RECT 95.105 133.255 95.515 133.695 ;
        RECT 95.685 133.315 96.700 133.515 ;
        RECT 92.975 132.885 94.225 133.055 ;
        RECT 92.975 132.765 93.305 132.885 ;
        RECT 91.635 132.375 93.535 132.545 ;
        RECT 91.275 132.035 93.195 132.205 ;
        RECT 91.275 132.015 91.595 132.035 ;
        RECT 90.825 131.355 91.155 131.865 ;
        RECT 91.425 131.405 91.595 132.015 ;
        RECT 93.365 131.865 93.535 132.375 ;
        RECT 93.705 132.305 93.885 132.715 ;
        RECT 94.055 132.125 94.225 132.885 ;
        RECT 91.765 131.145 92.095 131.835 ;
        RECT 92.325 131.695 93.535 131.865 ;
        RECT 93.705 131.815 94.225 132.125 ;
        RECT 94.395 132.715 94.815 133.055 ;
        RECT 95.105 132.715 95.515 133.045 ;
        RECT 94.395 131.945 94.585 132.715 ;
        RECT 95.685 132.585 95.855 133.315 ;
        RECT 97.000 133.145 97.170 133.475 ;
        RECT 97.340 133.315 97.670 133.695 ;
        RECT 96.025 132.765 96.375 133.135 ;
        RECT 95.685 132.545 96.105 132.585 ;
        RECT 94.755 132.375 96.105 132.545 ;
        RECT 94.755 132.215 95.005 132.375 ;
        RECT 95.515 131.945 95.765 132.205 ;
        RECT 94.395 131.695 95.765 131.945 ;
        RECT 92.325 131.405 92.565 131.695 ;
        RECT 93.365 131.615 93.535 131.695 ;
        RECT 92.765 131.145 93.185 131.525 ;
        RECT 93.365 131.365 93.995 131.615 ;
        RECT 94.465 131.145 94.795 131.525 ;
        RECT 94.965 131.405 95.135 131.695 ;
        RECT 95.935 131.530 96.105 132.375 ;
        RECT 96.555 132.205 96.775 133.075 ;
        RECT 97.000 132.955 97.695 133.145 ;
        RECT 96.275 131.825 96.775 132.205 ;
        RECT 96.945 132.155 97.355 132.775 ;
        RECT 97.525 131.985 97.695 132.955 ;
        RECT 97.000 131.815 97.695 131.985 ;
        RECT 95.315 131.145 95.695 131.525 ;
        RECT 95.935 131.360 96.765 131.530 ;
        RECT 97.000 131.315 97.170 131.815 ;
        RECT 97.340 131.145 97.670 131.645 ;
        RECT 97.885 131.315 98.110 133.435 ;
        RECT 98.280 133.315 98.610 133.695 ;
        RECT 98.780 133.145 98.950 133.435 ;
        RECT 98.285 132.975 98.950 133.145 ;
        RECT 98.285 131.985 98.515 132.975 ;
        RECT 99.210 132.970 99.500 133.695 ;
        RECT 99.730 132.875 99.940 133.695 ;
        RECT 100.110 132.895 100.440 133.525 ;
        RECT 98.685 132.155 99.035 132.805 ;
        RECT 98.285 131.815 98.950 131.985 ;
        RECT 98.280 131.145 98.610 131.645 ;
        RECT 98.780 131.315 98.950 131.815 ;
        RECT 99.210 131.145 99.500 132.310 ;
        RECT 100.110 132.295 100.360 132.895 ;
        RECT 100.610 132.875 100.840 133.695 ;
        RECT 101.785 132.885 102.030 133.490 ;
        RECT 102.250 133.160 102.760 133.695 ;
        RECT 101.510 132.715 102.740 132.885 ;
        RECT 100.530 132.455 100.860 132.705 ;
        RECT 99.730 131.145 99.940 132.285 ;
        RECT 100.110 131.315 100.440 132.295 ;
        RECT 100.610 131.145 100.840 132.285 ;
        RECT 101.510 131.905 101.850 132.715 ;
        RECT 102.020 132.150 102.770 132.340 ;
        RECT 101.510 131.495 102.025 131.905 ;
        RECT 102.260 131.145 102.430 131.905 ;
        RECT 102.600 131.485 102.770 132.150 ;
        RECT 102.940 132.165 103.130 133.525 ;
        RECT 103.300 132.675 103.575 133.525 ;
        RECT 103.765 133.160 104.295 133.525 ;
        RECT 104.720 133.295 105.050 133.695 ;
        RECT 104.120 133.125 104.295 133.160 ;
        RECT 103.300 132.505 103.580 132.675 ;
        RECT 103.300 132.365 103.575 132.505 ;
        RECT 103.780 132.165 103.950 132.965 ;
        RECT 102.940 131.995 103.950 132.165 ;
        RECT 104.120 132.955 105.050 133.125 ;
        RECT 105.220 132.955 105.475 133.525 ;
        RECT 106.660 133.145 106.830 133.525 ;
        RECT 107.010 133.315 107.340 133.695 ;
        RECT 106.660 132.975 107.325 133.145 ;
        RECT 107.520 133.020 107.780 133.525 ;
        RECT 104.120 131.825 104.290 132.955 ;
        RECT 104.880 132.785 105.050 132.955 ;
        RECT 103.165 131.655 104.290 131.825 ;
        RECT 104.460 132.455 104.655 132.785 ;
        RECT 104.880 132.455 105.135 132.785 ;
        RECT 104.460 131.485 104.630 132.455 ;
        RECT 105.305 132.285 105.475 132.955 ;
        RECT 106.590 132.425 106.920 132.795 ;
        RECT 107.155 132.720 107.325 132.975 ;
        RECT 102.600 131.315 104.630 131.485 ;
        RECT 104.800 131.145 104.970 132.285 ;
        RECT 105.140 131.315 105.475 132.285 ;
        RECT 107.155 132.390 107.440 132.720 ;
        RECT 107.155 132.245 107.325 132.390 ;
        RECT 106.660 132.075 107.325 132.245 ;
        RECT 107.610 132.220 107.780 133.020 ;
        RECT 108.410 132.925 111.000 133.695 ;
        RECT 111.170 132.945 112.380 133.695 ;
        RECT 106.660 131.315 106.830 132.075 ;
        RECT 107.010 131.145 107.340 131.905 ;
        RECT 107.510 131.315 107.780 132.220 ;
        RECT 108.410 132.235 109.620 132.755 ;
        RECT 109.790 132.405 111.000 132.925 ;
        RECT 111.170 132.235 111.690 132.775 ;
        RECT 111.860 132.405 112.380 132.945 ;
        RECT 108.410 131.145 111.000 132.235 ;
        RECT 111.170 131.145 112.380 132.235 ;
        RECT 18.165 130.975 112.465 131.145 ;
        RECT 18.250 129.885 19.460 130.975 ;
        RECT 19.745 130.345 20.030 130.805 ;
        RECT 20.200 130.515 20.470 130.975 ;
        RECT 19.745 130.125 20.700 130.345 ;
        RECT 18.250 129.175 18.770 129.715 ;
        RECT 18.940 129.345 19.460 129.885 ;
        RECT 19.630 129.395 20.320 129.955 ;
        RECT 20.490 129.225 20.700 130.125 ;
        RECT 18.250 128.425 19.460 129.175 ;
        RECT 19.745 129.055 20.700 129.225 ;
        RECT 20.870 129.955 21.270 130.805 ;
        RECT 21.460 130.345 21.740 130.805 ;
        RECT 22.260 130.515 22.585 130.975 ;
        RECT 21.460 130.125 22.585 130.345 ;
        RECT 20.870 129.395 21.965 129.955 ;
        RECT 22.135 129.665 22.585 130.125 ;
        RECT 22.755 129.835 23.140 130.805 ;
        RECT 19.745 128.595 20.030 129.055 ;
        RECT 20.200 128.425 20.470 128.885 ;
        RECT 20.870 128.595 21.270 129.395 ;
        RECT 22.135 129.335 22.690 129.665 ;
        RECT 22.135 129.225 22.585 129.335 ;
        RECT 21.460 129.055 22.585 129.225 ;
        RECT 22.860 129.165 23.140 129.835 ;
        RECT 23.310 129.885 24.520 130.975 ;
        RECT 23.310 129.345 23.830 129.885 ;
        RECT 24.695 129.835 25.030 130.805 ;
        RECT 25.200 129.835 25.370 130.975 ;
        RECT 25.540 130.635 27.570 130.805 ;
        RECT 24.000 129.175 24.520 129.715 ;
        RECT 21.460 128.595 21.740 129.055 ;
        RECT 22.260 128.425 22.585 128.885 ;
        RECT 22.755 128.595 23.140 129.165 ;
        RECT 23.310 128.425 24.520 129.175 ;
        RECT 24.695 129.165 24.865 129.835 ;
        RECT 25.540 129.665 25.710 130.635 ;
        RECT 25.035 129.335 25.290 129.665 ;
        RECT 25.515 129.335 25.710 129.665 ;
        RECT 25.880 130.295 27.005 130.465 ;
        RECT 25.120 129.165 25.290 129.335 ;
        RECT 25.880 129.165 26.050 130.295 ;
        RECT 24.695 128.595 24.950 129.165 ;
        RECT 25.120 128.995 26.050 129.165 ;
        RECT 26.220 129.955 27.230 130.125 ;
        RECT 26.220 129.155 26.390 129.955 ;
        RECT 25.875 128.960 26.050 128.995 ;
        RECT 25.120 128.425 25.450 128.825 ;
        RECT 25.875 128.595 26.405 128.960 ;
        RECT 26.595 128.935 26.870 129.755 ;
        RECT 26.590 128.765 26.870 128.935 ;
        RECT 26.595 128.595 26.870 128.765 ;
        RECT 27.040 128.595 27.230 129.955 ;
        RECT 27.400 129.970 27.570 130.635 ;
        RECT 27.740 130.215 27.910 130.975 ;
        RECT 28.145 130.215 28.660 130.625 ;
        RECT 27.400 129.780 28.150 129.970 ;
        RECT 28.320 129.405 28.660 130.215 ;
        RECT 27.430 129.235 28.660 129.405 ;
        RECT 28.830 129.885 30.040 130.975 ;
        RECT 28.830 129.345 29.350 129.885 ;
        RECT 30.270 129.835 30.480 130.975 ;
        RECT 30.650 129.825 30.980 130.805 ;
        RECT 31.150 129.835 31.380 130.975 ;
        RECT 32.050 129.885 34.640 130.975 ;
        RECT 27.410 128.425 27.920 128.960 ;
        RECT 28.140 128.630 28.385 129.235 ;
        RECT 29.520 129.175 30.040 129.715 ;
        RECT 28.830 128.425 30.040 129.175 ;
        RECT 30.270 128.425 30.480 129.245 ;
        RECT 30.650 129.225 30.900 129.825 ;
        RECT 31.070 129.415 31.400 129.665 ;
        RECT 32.050 129.365 33.260 129.885 ;
        RECT 34.810 129.810 35.100 130.975 ;
        RECT 35.730 129.900 36.000 130.805 ;
        RECT 36.170 130.215 36.500 130.975 ;
        RECT 36.680 130.045 36.850 130.805 ;
        RECT 37.310 130.305 37.590 130.975 ;
        RECT 30.650 128.595 30.980 129.225 ;
        RECT 31.150 128.425 31.380 129.245 ;
        RECT 33.430 129.195 34.640 129.715 ;
        RECT 32.050 128.425 34.640 129.195 ;
        RECT 34.810 128.425 35.100 129.150 ;
        RECT 35.730 129.100 35.900 129.900 ;
        RECT 36.185 129.875 36.850 130.045 ;
        RECT 37.760 130.085 38.060 130.635 ;
        RECT 38.260 130.255 38.590 130.975 ;
        RECT 38.780 130.255 39.240 130.805 ;
        RECT 39.415 130.465 41.070 130.755 ;
        RECT 36.185 129.730 36.355 129.875 ;
        RECT 36.070 129.400 36.355 129.730 ;
        RECT 36.185 129.145 36.355 129.400 ;
        RECT 36.590 129.325 36.920 129.695 ;
        RECT 37.125 129.665 37.390 130.025 ;
        RECT 37.760 129.915 38.700 130.085 ;
        RECT 38.530 129.665 38.700 129.915 ;
        RECT 37.125 129.415 37.800 129.665 ;
        RECT 38.020 129.415 38.360 129.665 ;
        RECT 38.530 129.335 38.820 129.665 ;
        RECT 38.530 129.245 38.700 129.335 ;
        RECT 35.730 128.595 35.990 129.100 ;
        RECT 36.185 128.975 36.850 129.145 ;
        RECT 36.170 128.425 36.500 128.805 ;
        RECT 36.680 128.595 36.850 128.975 ;
        RECT 37.310 129.055 38.700 129.245 ;
        RECT 37.310 128.695 37.640 129.055 ;
        RECT 38.990 128.885 39.240 130.255 ;
        RECT 39.415 130.125 41.005 130.295 ;
        RECT 41.240 130.175 41.520 130.975 ;
        RECT 39.415 129.835 39.735 130.125 ;
        RECT 40.835 130.005 41.005 130.125 ;
        RECT 39.415 129.095 39.765 129.665 ;
        RECT 39.935 129.335 40.645 129.955 ;
        RECT 40.835 129.835 41.560 130.005 ;
        RECT 41.730 129.835 42.000 130.805 ;
        RECT 42.175 130.465 43.830 130.755 ;
        RECT 42.175 130.125 43.765 130.295 ;
        RECT 44.000 130.175 44.280 130.975 ;
        RECT 42.175 129.835 42.495 130.125 ;
        RECT 43.595 130.005 43.765 130.125 ;
        RECT 41.390 129.665 41.560 129.835 ;
        RECT 40.815 129.335 41.220 129.665 ;
        RECT 41.390 129.335 41.660 129.665 ;
        RECT 41.390 129.165 41.560 129.335 ;
        RECT 39.950 128.995 41.560 129.165 ;
        RECT 41.830 129.100 42.000 129.835 ;
        RECT 38.260 128.425 38.510 128.885 ;
        RECT 38.680 128.595 39.240 128.885 ;
        RECT 39.420 128.425 39.750 128.925 ;
        RECT 39.950 128.645 40.120 128.995 ;
        RECT 40.320 128.425 40.650 128.825 ;
        RECT 40.820 128.645 40.990 128.995 ;
        RECT 41.160 128.425 41.540 128.825 ;
        RECT 41.730 128.755 42.000 129.100 ;
        RECT 42.175 129.095 42.525 129.665 ;
        RECT 42.695 129.335 43.405 129.955 ;
        RECT 43.595 129.835 44.320 130.005 ;
        RECT 44.490 129.835 44.760 130.805 ;
        RECT 44.150 129.665 44.320 129.835 ;
        RECT 43.575 129.335 43.980 129.665 ;
        RECT 44.150 129.335 44.420 129.665 ;
        RECT 44.150 129.165 44.320 129.335 ;
        RECT 42.710 128.995 44.320 129.165 ;
        RECT 44.590 129.100 44.760 129.835 ;
        RECT 42.180 128.425 42.510 128.925 ;
        RECT 42.710 128.645 42.880 128.995 ;
        RECT 43.080 128.425 43.410 128.825 ;
        RECT 43.580 128.645 43.750 128.995 ;
        RECT 43.920 128.425 44.300 128.825 ;
        RECT 44.490 128.755 44.760 129.100 ;
        RECT 44.930 129.835 45.200 130.805 ;
        RECT 45.410 130.175 45.690 130.975 ;
        RECT 45.860 130.465 47.515 130.755 ;
        RECT 45.925 130.125 47.515 130.295 ;
        RECT 45.925 130.005 46.095 130.125 ;
        RECT 45.370 129.835 46.095 130.005 ;
        RECT 44.930 129.100 45.100 129.835 ;
        RECT 45.370 129.665 45.540 129.835 ;
        RECT 46.285 129.785 47.000 129.955 ;
        RECT 47.195 129.835 47.515 130.125 ;
        RECT 48.150 129.835 48.490 130.805 ;
        RECT 48.660 129.835 48.830 130.975 ;
        RECT 49.100 130.175 49.350 130.975 ;
        RECT 49.995 130.005 50.325 130.805 ;
        RECT 50.625 130.175 50.955 130.975 ;
        RECT 51.125 130.005 51.455 130.805 ;
        RECT 49.020 129.835 51.455 130.005 ;
        RECT 51.830 129.835 52.170 130.805 ;
        RECT 52.340 129.835 52.510 130.975 ;
        RECT 52.780 130.175 53.030 130.975 ;
        RECT 53.675 130.005 54.005 130.805 ;
        RECT 54.305 130.175 54.635 130.975 ;
        RECT 54.805 130.005 55.135 130.805 ;
        RECT 52.700 129.835 55.135 130.005 ;
        RECT 56.430 130.215 56.945 130.625 ;
        RECT 57.180 130.215 57.350 130.975 ;
        RECT 57.520 130.635 59.550 130.805 ;
        RECT 45.270 129.335 45.540 129.665 ;
        RECT 45.710 129.335 46.115 129.665 ;
        RECT 46.285 129.335 46.995 129.785 ;
        RECT 45.370 129.165 45.540 129.335 ;
        RECT 44.930 128.755 45.200 129.100 ;
        RECT 45.370 128.995 46.980 129.165 ;
        RECT 47.165 129.095 47.515 129.665 ;
        RECT 48.150 129.275 48.325 129.835 ;
        RECT 49.020 129.585 49.190 129.835 ;
        RECT 48.495 129.415 49.190 129.585 ;
        RECT 49.365 129.415 49.785 129.615 ;
        RECT 49.955 129.415 50.285 129.615 ;
        RECT 50.455 129.415 50.785 129.615 ;
        RECT 48.150 129.225 48.380 129.275 ;
        RECT 45.390 128.425 45.770 128.825 ;
        RECT 45.940 128.645 46.110 128.995 ;
        RECT 46.280 128.425 46.610 128.825 ;
        RECT 46.810 128.645 46.980 128.995 ;
        RECT 47.180 128.425 47.510 128.925 ;
        RECT 48.150 128.595 48.490 129.225 ;
        RECT 48.660 128.425 48.910 129.225 ;
        RECT 49.100 129.075 50.325 129.245 ;
        RECT 49.100 128.595 49.430 129.075 ;
        RECT 49.600 128.425 49.825 128.885 ;
        RECT 49.995 128.595 50.325 129.075 ;
        RECT 50.955 129.205 51.125 129.835 ;
        RECT 51.310 129.415 51.660 129.665 ;
        RECT 51.830 129.275 52.005 129.835 ;
        RECT 52.700 129.585 52.870 129.835 ;
        RECT 52.175 129.415 52.870 129.585 ;
        RECT 53.045 129.415 53.465 129.615 ;
        RECT 53.635 129.415 53.965 129.615 ;
        RECT 54.135 129.415 54.465 129.615 ;
        RECT 51.830 129.225 52.060 129.275 ;
        RECT 50.955 128.595 51.455 129.205 ;
        RECT 51.830 128.595 52.170 129.225 ;
        RECT 52.340 128.425 52.590 129.225 ;
        RECT 52.780 129.075 54.005 129.245 ;
        RECT 52.780 128.595 53.110 129.075 ;
        RECT 53.280 128.425 53.505 128.885 ;
        RECT 53.675 128.595 54.005 129.075 ;
        RECT 54.635 129.205 54.805 129.835 ;
        RECT 54.990 129.415 55.340 129.665 ;
        RECT 56.430 129.405 56.770 130.215 ;
        RECT 57.520 129.970 57.690 130.635 ;
        RECT 58.085 130.295 59.210 130.465 ;
        RECT 56.940 129.780 57.690 129.970 ;
        RECT 57.860 129.955 58.870 130.125 ;
        RECT 56.430 129.235 57.660 129.405 ;
        RECT 54.635 128.595 55.135 129.205 ;
        RECT 56.705 128.630 56.950 129.235 ;
        RECT 57.170 128.425 57.680 128.960 ;
        RECT 57.860 128.595 58.050 129.955 ;
        RECT 58.220 129.615 58.495 129.755 ;
        RECT 58.220 129.445 58.500 129.615 ;
        RECT 58.220 128.595 58.495 129.445 ;
        RECT 58.700 129.155 58.870 129.955 ;
        RECT 59.040 129.165 59.210 130.295 ;
        RECT 59.380 129.665 59.550 130.635 ;
        RECT 59.720 129.835 59.890 130.975 ;
        RECT 60.060 129.835 60.395 130.805 ;
        RECT 59.380 129.335 59.575 129.665 ;
        RECT 59.800 129.335 60.055 129.665 ;
        RECT 59.800 129.165 59.970 129.335 ;
        RECT 60.225 129.165 60.395 129.835 ;
        RECT 60.570 129.810 60.860 130.975 ;
        RECT 61.405 129.995 61.660 130.665 ;
        RECT 61.840 130.175 62.125 130.975 ;
        RECT 62.305 130.255 62.635 130.765 ;
        RECT 59.040 128.995 59.970 129.165 ;
        RECT 59.040 128.960 59.215 128.995 ;
        RECT 58.685 128.595 59.215 128.960 ;
        RECT 59.640 128.425 59.970 128.825 ;
        RECT 60.140 128.595 60.395 129.165 ;
        RECT 60.570 128.425 60.860 129.150 ;
        RECT 61.405 129.135 61.585 129.995 ;
        RECT 62.305 129.665 62.555 130.255 ;
        RECT 62.905 130.105 63.075 130.715 ;
        RECT 63.245 130.285 63.575 130.975 ;
        RECT 63.805 130.425 64.045 130.715 ;
        RECT 64.245 130.595 64.665 130.975 ;
        RECT 64.845 130.505 65.475 130.755 ;
        RECT 65.945 130.595 66.275 130.975 ;
        RECT 64.845 130.425 65.015 130.505 ;
        RECT 66.445 130.425 66.615 130.715 ;
        RECT 66.795 130.595 67.175 130.975 ;
        RECT 67.415 130.590 68.245 130.760 ;
        RECT 63.805 130.255 65.015 130.425 ;
        RECT 61.755 129.335 62.555 129.665 ;
        RECT 61.405 128.935 61.660 129.135 ;
        RECT 61.320 128.765 61.660 128.935 ;
        RECT 61.405 128.605 61.660 128.765 ;
        RECT 61.840 128.425 62.125 128.885 ;
        RECT 62.305 128.685 62.555 129.335 ;
        RECT 62.755 130.085 63.075 130.105 ;
        RECT 62.755 129.915 64.675 130.085 ;
        RECT 62.755 129.020 62.945 129.915 ;
        RECT 64.845 129.745 65.015 130.255 ;
        RECT 65.185 129.995 65.705 130.305 ;
        RECT 63.115 129.575 65.015 129.745 ;
        RECT 63.115 129.515 63.445 129.575 ;
        RECT 63.595 129.345 63.925 129.405 ;
        RECT 63.265 129.075 63.925 129.345 ;
        RECT 62.755 128.690 63.075 129.020 ;
        RECT 63.255 128.425 63.915 128.905 ;
        RECT 64.115 128.815 64.285 129.575 ;
        RECT 65.185 129.405 65.365 129.815 ;
        RECT 64.455 129.235 64.785 129.355 ;
        RECT 65.535 129.235 65.705 129.995 ;
        RECT 64.455 129.065 65.705 129.235 ;
        RECT 65.875 130.175 67.245 130.425 ;
        RECT 65.875 129.405 66.065 130.175 ;
        RECT 66.995 129.915 67.245 130.175 ;
        RECT 66.235 129.745 66.485 129.905 ;
        RECT 67.415 129.745 67.585 130.590 ;
        RECT 68.480 130.305 68.650 130.805 ;
        RECT 68.820 130.475 69.150 130.975 ;
        RECT 67.755 129.915 68.255 130.295 ;
        RECT 68.480 130.135 69.175 130.305 ;
        RECT 66.235 129.575 67.585 129.745 ;
        RECT 67.165 129.535 67.585 129.575 ;
        RECT 65.875 129.065 66.295 129.405 ;
        RECT 66.585 129.075 66.995 129.405 ;
        RECT 64.115 128.645 64.965 128.815 ;
        RECT 65.525 128.425 65.845 128.885 ;
        RECT 66.045 128.635 66.295 129.065 ;
        RECT 66.585 128.425 66.995 128.865 ;
        RECT 67.165 128.805 67.335 129.535 ;
        RECT 67.505 128.985 67.855 129.355 ;
        RECT 68.035 129.045 68.255 129.915 ;
        RECT 68.425 129.345 68.835 129.965 ;
        RECT 69.005 129.165 69.175 130.135 ;
        RECT 68.480 128.975 69.175 129.165 ;
        RECT 67.165 128.605 68.180 128.805 ;
        RECT 68.480 128.645 68.650 128.975 ;
        RECT 68.820 128.425 69.150 128.805 ;
        RECT 69.365 128.685 69.590 130.805 ;
        RECT 69.760 130.475 70.090 130.975 ;
        RECT 70.260 130.305 70.430 130.805 ;
        RECT 69.765 130.135 70.430 130.305 ;
        RECT 70.690 130.255 71.150 130.805 ;
        RECT 71.340 130.255 71.670 130.975 ;
        RECT 69.765 129.145 69.995 130.135 ;
        RECT 70.165 129.315 70.515 129.965 ;
        RECT 69.765 128.975 70.430 129.145 ;
        RECT 69.760 128.425 70.090 128.805 ;
        RECT 70.260 128.685 70.430 128.975 ;
        RECT 70.690 128.885 70.940 130.255 ;
        RECT 71.870 130.085 72.170 130.635 ;
        RECT 72.340 130.305 72.620 130.975 ;
        RECT 71.230 129.915 72.170 130.085 ;
        RECT 71.230 129.665 71.400 129.915 ;
        RECT 72.540 129.665 72.805 130.025 ;
        RECT 71.110 129.335 71.400 129.665 ;
        RECT 71.570 129.415 71.910 129.665 ;
        RECT 72.130 129.415 72.805 129.665 ;
        RECT 72.990 129.835 73.330 130.805 ;
        RECT 73.500 129.835 73.670 130.975 ;
        RECT 73.940 130.175 74.190 130.975 ;
        RECT 74.835 130.005 75.165 130.805 ;
        RECT 75.465 130.175 75.795 130.975 ;
        RECT 75.965 130.005 76.295 130.805 ;
        RECT 73.860 129.835 76.295 130.005 ;
        RECT 77.045 129.995 77.300 130.665 ;
        RECT 77.480 130.175 77.765 130.975 ;
        RECT 77.945 130.255 78.275 130.765 ;
        RECT 71.230 129.245 71.400 129.335 ;
        RECT 71.230 129.055 72.620 129.245 ;
        RECT 70.690 128.595 71.250 128.885 ;
        RECT 71.420 128.425 71.670 128.885 ;
        RECT 72.290 128.695 72.620 129.055 ;
        RECT 72.990 129.225 73.165 129.835 ;
        RECT 73.860 129.585 74.030 129.835 ;
        RECT 73.335 129.415 74.030 129.585 ;
        RECT 74.205 129.415 74.625 129.615 ;
        RECT 74.795 129.415 75.125 129.615 ;
        RECT 75.295 129.415 75.625 129.615 ;
        RECT 72.990 128.595 73.330 129.225 ;
        RECT 73.500 128.425 73.750 129.225 ;
        RECT 73.940 129.075 75.165 129.245 ;
        RECT 73.940 128.595 74.270 129.075 ;
        RECT 74.440 128.425 74.665 128.885 ;
        RECT 74.835 128.595 75.165 129.075 ;
        RECT 75.795 129.205 75.965 129.835 ;
        RECT 76.150 129.415 76.500 129.665 ;
        RECT 75.795 128.595 76.295 129.205 ;
        RECT 77.045 129.135 77.225 129.995 ;
        RECT 77.945 129.665 78.195 130.255 ;
        RECT 78.545 130.105 78.715 130.715 ;
        RECT 78.885 130.285 79.215 130.975 ;
        RECT 79.445 130.425 79.685 130.715 ;
        RECT 79.885 130.595 80.305 130.975 ;
        RECT 80.485 130.505 81.115 130.755 ;
        RECT 81.585 130.595 81.915 130.975 ;
        RECT 80.485 130.425 80.655 130.505 ;
        RECT 82.085 130.425 82.255 130.715 ;
        RECT 82.435 130.595 82.815 130.975 ;
        RECT 83.055 130.590 83.885 130.760 ;
        RECT 79.445 130.255 80.655 130.425 ;
        RECT 77.395 129.335 78.195 129.665 ;
        RECT 77.045 128.935 77.300 129.135 ;
        RECT 76.960 128.765 77.300 128.935 ;
        RECT 77.045 128.605 77.300 128.765 ;
        RECT 77.480 128.425 77.765 128.885 ;
        RECT 77.945 128.685 78.195 129.335 ;
        RECT 78.395 130.085 78.715 130.105 ;
        RECT 78.395 129.915 80.315 130.085 ;
        RECT 78.395 129.020 78.585 129.915 ;
        RECT 80.485 129.745 80.655 130.255 ;
        RECT 80.825 129.995 81.345 130.305 ;
        RECT 78.755 129.575 80.655 129.745 ;
        RECT 78.755 129.515 79.085 129.575 ;
        RECT 79.235 129.345 79.565 129.405 ;
        RECT 78.905 129.075 79.565 129.345 ;
        RECT 78.395 128.690 78.715 129.020 ;
        RECT 78.895 128.425 79.555 128.905 ;
        RECT 79.755 128.815 79.925 129.575 ;
        RECT 80.825 129.405 81.005 129.815 ;
        RECT 80.095 129.235 80.425 129.355 ;
        RECT 81.175 129.235 81.345 129.995 ;
        RECT 80.095 129.065 81.345 129.235 ;
        RECT 81.515 130.175 82.885 130.425 ;
        RECT 81.515 129.405 81.705 130.175 ;
        RECT 82.635 129.915 82.885 130.175 ;
        RECT 81.875 129.745 82.125 129.905 ;
        RECT 83.055 129.745 83.225 130.590 ;
        RECT 84.120 130.305 84.290 130.805 ;
        RECT 84.460 130.475 84.790 130.975 ;
        RECT 83.395 129.915 83.895 130.295 ;
        RECT 84.120 130.135 84.815 130.305 ;
        RECT 81.875 129.575 83.225 129.745 ;
        RECT 82.805 129.535 83.225 129.575 ;
        RECT 81.515 129.065 81.935 129.405 ;
        RECT 82.225 129.075 82.635 129.405 ;
        RECT 79.755 128.645 80.605 128.815 ;
        RECT 81.165 128.425 81.485 128.885 ;
        RECT 81.685 128.635 81.935 129.065 ;
        RECT 82.225 128.425 82.635 128.865 ;
        RECT 82.805 128.805 82.975 129.535 ;
        RECT 83.145 128.985 83.495 129.355 ;
        RECT 83.675 129.045 83.895 129.915 ;
        RECT 84.065 129.345 84.475 129.965 ;
        RECT 84.645 129.165 84.815 130.135 ;
        RECT 84.120 128.975 84.815 129.165 ;
        RECT 82.805 128.605 83.820 128.805 ;
        RECT 84.120 128.645 84.290 128.975 ;
        RECT 84.460 128.425 84.790 128.805 ;
        RECT 85.005 128.685 85.230 130.805 ;
        RECT 85.400 130.475 85.730 130.975 ;
        RECT 85.900 130.305 86.070 130.805 ;
        RECT 85.405 130.135 86.070 130.305 ;
        RECT 85.405 129.145 85.635 130.135 ;
        RECT 85.805 129.315 86.155 129.965 ;
        RECT 86.330 129.810 86.620 130.975 ;
        RECT 86.850 129.835 87.060 130.975 ;
        RECT 87.230 129.825 87.560 130.805 ;
        RECT 87.730 129.835 87.960 130.975 ;
        RECT 88.545 130.295 88.800 130.665 ;
        RECT 88.460 130.125 88.800 130.295 ;
        RECT 88.980 130.175 89.265 130.975 ;
        RECT 89.445 130.255 89.775 130.765 ;
        RECT 88.545 129.995 88.800 130.125 ;
        RECT 85.405 128.975 86.070 129.145 ;
        RECT 85.400 128.425 85.730 128.805 ;
        RECT 85.900 128.685 86.070 128.975 ;
        RECT 86.330 128.425 86.620 129.150 ;
        RECT 86.850 128.425 87.060 129.245 ;
        RECT 87.230 129.225 87.480 129.825 ;
        RECT 87.650 129.415 87.980 129.665 ;
        RECT 87.230 128.595 87.560 129.225 ;
        RECT 87.730 128.425 87.960 129.245 ;
        RECT 88.545 129.135 88.725 129.995 ;
        RECT 89.445 129.665 89.695 130.255 ;
        RECT 90.045 130.105 90.215 130.715 ;
        RECT 90.385 130.285 90.715 130.975 ;
        RECT 90.945 130.425 91.185 130.715 ;
        RECT 91.385 130.595 91.805 130.975 ;
        RECT 91.985 130.505 92.615 130.755 ;
        RECT 93.085 130.595 93.415 130.975 ;
        RECT 91.985 130.425 92.155 130.505 ;
        RECT 93.585 130.425 93.755 130.715 ;
        RECT 93.935 130.595 94.315 130.975 ;
        RECT 94.555 130.590 95.385 130.760 ;
        RECT 90.945 130.255 92.155 130.425 ;
        RECT 88.895 129.335 89.695 129.665 ;
        RECT 88.545 128.605 88.800 129.135 ;
        RECT 88.980 128.425 89.265 128.885 ;
        RECT 89.445 128.685 89.695 129.335 ;
        RECT 89.895 130.085 90.215 130.105 ;
        RECT 89.895 129.915 91.815 130.085 ;
        RECT 89.895 129.020 90.085 129.915 ;
        RECT 91.985 129.745 92.155 130.255 ;
        RECT 92.325 129.995 92.845 130.305 ;
        RECT 90.255 129.575 92.155 129.745 ;
        RECT 90.255 129.515 90.585 129.575 ;
        RECT 90.735 129.345 91.065 129.405 ;
        RECT 90.405 129.075 91.065 129.345 ;
        RECT 89.895 128.690 90.215 129.020 ;
        RECT 90.395 128.425 91.055 128.905 ;
        RECT 91.255 128.815 91.425 129.575 ;
        RECT 92.325 129.405 92.505 129.815 ;
        RECT 91.595 129.235 91.925 129.355 ;
        RECT 92.675 129.235 92.845 129.995 ;
        RECT 91.595 129.065 92.845 129.235 ;
        RECT 93.015 130.175 94.385 130.425 ;
        RECT 93.015 129.405 93.205 130.175 ;
        RECT 94.135 129.915 94.385 130.175 ;
        RECT 93.375 129.745 93.625 129.905 ;
        RECT 94.555 129.745 94.725 130.590 ;
        RECT 95.620 130.305 95.790 130.805 ;
        RECT 95.960 130.475 96.290 130.975 ;
        RECT 94.895 129.915 95.395 130.295 ;
        RECT 95.620 130.135 96.315 130.305 ;
        RECT 93.375 129.575 94.725 129.745 ;
        RECT 94.305 129.535 94.725 129.575 ;
        RECT 93.015 129.065 93.435 129.405 ;
        RECT 93.725 129.075 94.135 129.405 ;
        RECT 91.255 128.645 92.105 128.815 ;
        RECT 92.665 128.425 92.985 128.885 ;
        RECT 93.185 128.635 93.435 129.065 ;
        RECT 93.725 128.425 94.135 128.865 ;
        RECT 94.305 128.805 94.475 129.535 ;
        RECT 94.645 128.985 94.995 129.355 ;
        RECT 95.175 129.045 95.395 129.915 ;
        RECT 95.565 129.345 95.975 129.965 ;
        RECT 96.145 129.165 96.315 130.135 ;
        RECT 95.620 128.975 96.315 129.165 ;
        RECT 94.305 128.605 95.320 128.805 ;
        RECT 95.620 128.645 95.790 128.975 ;
        RECT 95.960 128.425 96.290 128.805 ;
        RECT 96.505 128.685 96.730 130.805 ;
        RECT 96.900 130.475 97.230 130.975 ;
        RECT 97.400 130.305 97.570 130.805 ;
        RECT 96.905 130.135 97.570 130.305 ;
        RECT 96.905 129.145 97.135 130.135 ;
        RECT 97.305 129.315 97.655 129.965 ;
        RECT 97.830 129.900 98.100 130.805 ;
        RECT 98.270 130.215 98.600 130.975 ;
        RECT 98.780 130.045 98.950 130.805 ;
        RECT 96.905 128.975 97.570 129.145 ;
        RECT 96.900 128.425 97.230 128.805 ;
        RECT 97.400 128.685 97.570 128.975 ;
        RECT 97.830 129.100 98.000 129.900 ;
        RECT 98.285 129.875 98.950 130.045 ;
        RECT 99.670 129.900 99.940 130.805 ;
        RECT 100.110 130.215 100.440 130.975 ;
        RECT 100.620 130.045 100.790 130.805 ;
        RECT 98.285 129.730 98.455 129.875 ;
        RECT 98.170 129.400 98.455 129.730 ;
        RECT 98.285 129.145 98.455 129.400 ;
        RECT 98.690 129.325 99.020 129.695 ;
        RECT 97.830 128.595 98.090 129.100 ;
        RECT 98.285 128.975 98.950 129.145 ;
        RECT 98.270 128.425 98.600 128.805 ;
        RECT 98.780 128.595 98.950 128.975 ;
        RECT 99.670 129.100 99.840 129.900 ;
        RECT 100.125 129.875 100.790 130.045 ;
        RECT 101.970 129.885 105.480 130.975 ;
        RECT 105.655 130.540 111.000 130.975 ;
        RECT 100.125 129.730 100.295 129.875 ;
        RECT 100.010 129.400 100.295 129.730 ;
        RECT 100.125 129.145 100.295 129.400 ;
        RECT 100.530 129.325 100.860 129.695 ;
        RECT 101.970 129.365 103.660 129.885 ;
        RECT 103.830 129.195 105.480 129.715 ;
        RECT 107.245 129.290 107.595 130.540 ;
        RECT 111.170 129.885 112.380 130.975 ;
        RECT 99.670 128.595 99.930 129.100 ;
        RECT 100.125 128.975 100.790 129.145 ;
        RECT 100.110 128.425 100.440 128.805 ;
        RECT 100.620 128.595 100.790 128.975 ;
        RECT 101.970 128.425 105.480 129.195 ;
        RECT 109.075 128.970 109.415 129.800 ;
        RECT 111.170 129.345 111.690 129.885 ;
        RECT 111.860 129.175 112.380 129.715 ;
        RECT 105.655 128.425 111.000 128.970 ;
        RECT 111.170 128.425 112.380 129.175 ;
        RECT 18.165 128.255 112.465 128.425 ;
        RECT 18.250 127.505 19.460 128.255 ;
        RECT 18.250 126.965 18.770 127.505 ;
        RECT 20.610 127.435 20.820 128.255 ;
        RECT 20.990 127.455 21.320 128.085 ;
        RECT 18.940 126.795 19.460 127.335 ;
        RECT 20.990 126.855 21.240 127.455 ;
        RECT 21.490 127.435 21.720 128.255 ;
        RECT 21.930 127.530 22.220 128.255 ;
        RECT 22.765 127.545 23.020 128.075 ;
        RECT 23.200 127.795 23.485 128.255 ;
        RECT 21.410 127.015 21.740 127.265 ;
        RECT 18.250 125.705 19.460 126.795 ;
        RECT 20.610 125.705 20.820 126.845 ;
        RECT 20.990 125.875 21.320 126.855 ;
        RECT 21.490 125.705 21.720 126.845 ;
        RECT 21.930 125.705 22.220 126.870 ;
        RECT 22.765 126.685 22.945 127.545 ;
        RECT 23.665 127.345 23.915 127.995 ;
        RECT 23.115 127.015 23.915 127.345 ;
        RECT 22.765 126.215 23.020 126.685 ;
        RECT 22.680 126.045 23.020 126.215 ;
        RECT 22.765 126.015 23.020 126.045 ;
        RECT 23.200 125.705 23.485 126.505 ;
        RECT 23.665 126.425 23.915 127.015 ;
        RECT 24.115 127.660 24.435 127.990 ;
        RECT 24.615 127.775 25.275 128.255 ;
        RECT 25.475 127.865 26.325 128.035 ;
        RECT 24.115 126.765 24.305 127.660 ;
        RECT 24.625 127.335 25.285 127.605 ;
        RECT 24.955 127.275 25.285 127.335 ;
        RECT 24.475 127.105 24.805 127.165 ;
        RECT 25.475 127.105 25.645 127.865 ;
        RECT 26.885 127.795 27.205 128.255 ;
        RECT 27.405 127.615 27.655 128.045 ;
        RECT 27.945 127.815 28.355 128.255 ;
        RECT 28.525 127.875 29.540 128.075 ;
        RECT 25.815 127.445 27.065 127.615 ;
        RECT 25.815 127.325 26.145 127.445 ;
        RECT 24.475 126.935 26.375 127.105 ;
        RECT 24.115 126.595 26.035 126.765 ;
        RECT 24.115 126.575 24.435 126.595 ;
        RECT 23.665 125.915 23.995 126.425 ;
        RECT 24.265 125.965 24.435 126.575 ;
        RECT 26.205 126.425 26.375 126.935 ;
        RECT 26.545 126.865 26.725 127.275 ;
        RECT 26.895 126.685 27.065 127.445 ;
        RECT 24.605 125.705 24.935 126.395 ;
        RECT 25.165 126.255 26.375 126.425 ;
        RECT 26.545 126.375 27.065 126.685 ;
        RECT 27.235 127.275 27.655 127.615 ;
        RECT 27.945 127.275 28.355 127.605 ;
        RECT 27.235 126.505 27.425 127.275 ;
        RECT 28.525 127.145 28.695 127.875 ;
        RECT 29.840 127.705 30.010 128.035 ;
        RECT 30.180 127.875 30.510 128.255 ;
        RECT 28.865 127.325 29.215 127.695 ;
        RECT 28.525 127.105 28.945 127.145 ;
        RECT 27.595 126.935 28.945 127.105 ;
        RECT 27.595 126.775 27.845 126.935 ;
        RECT 28.355 126.505 28.605 126.765 ;
        RECT 27.235 126.255 28.605 126.505 ;
        RECT 25.165 125.965 25.405 126.255 ;
        RECT 26.205 126.175 26.375 126.255 ;
        RECT 25.605 125.705 26.025 126.085 ;
        RECT 26.205 125.925 26.835 126.175 ;
        RECT 27.305 125.705 27.635 126.085 ;
        RECT 27.805 125.965 27.975 126.255 ;
        RECT 28.775 126.090 28.945 126.935 ;
        RECT 29.395 126.765 29.615 127.635 ;
        RECT 29.840 127.515 30.535 127.705 ;
        RECT 29.115 126.385 29.615 126.765 ;
        RECT 29.785 126.715 30.195 127.335 ;
        RECT 30.365 126.545 30.535 127.515 ;
        RECT 29.840 126.375 30.535 126.545 ;
        RECT 28.155 125.705 28.535 126.085 ;
        RECT 28.775 125.920 29.605 126.090 ;
        RECT 29.840 125.875 30.010 126.375 ;
        RECT 30.180 125.705 30.510 126.205 ;
        RECT 30.725 125.875 30.950 127.995 ;
        RECT 31.120 127.875 31.450 128.255 ;
        RECT 31.620 127.705 31.790 127.995 ;
        RECT 31.125 127.535 31.790 127.705 ;
        RECT 31.125 126.545 31.355 127.535 ;
        RECT 32.325 127.445 32.570 128.050 ;
        RECT 32.790 127.720 33.300 128.255 ;
        RECT 31.525 126.715 31.875 127.365 ;
        RECT 32.050 127.275 33.280 127.445 ;
        RECT 31.125 126.375 31.790 126.545 ;
        RECT 31.120 125.705 31.450 126.205 ;
        RECT 31.620 125.875 31.790 126.375 ;
        RECT 32.050 126.465 32.390 127.275 ;
        RECT 32.560 126.710 33.310 126.900 ;
        RECT 32.050 126.055 32.565 126.465 ;
        RECT 32.800 125.705 32.970 126.465 ;
        RECT 33.140 126.045 33.310 126.710 ;
        RECT 33.480 126.725 33.670 128.085 ;
        RECT 33.840 127.915 34.115 128.085 ;
        RECT 33.840 127.745 34.120 127.915 ;
        RECT 33.840 126.925 34.115 127.745 ;
        RECT 34.305 127.720 34.835 128.085 ;
        RECT 35.260 127.855 35.590 128.255 ;
        RECT 34.660 127.685 34.835 127.720 ;
        RECT 34.320 126.725 34.490 127.525 ;
        RECT 33.480 126.555 34.490 126.725 ;
        RECT 34.660 127.515 35.590 127.685 ;
        RECT 35.760 127.515 36.015 128.085 ;
        RECT 36.740 127.705 36.910 128.085 ;
        RECT 37.090 127.875 37.420 128.255 ;
        RECT 36.740 127.535 37.405 127.705 ;
        RECT 37.600 127.580 37.860 128.085 ;
        RECT 34.660 126.385 34.830 127.515 ;
        RECT 35.420 127.345 35.590 127.515 ;
        RECT 33.705 126.215 34.830 126.385 ;
        RECT 35.000 127.015 35.195 127.345 ;
        RECT 35.420 127.015 35.675 127.345 ;
        RECT 35.000 126.045 35.170 127.015 ;
        RECT 35.845 126.845 36.015 127.515 ;
        RECT 36.670 126.985 37.000 127.355 ;
        RECT 37.235 127.280 37.405 127.535 ;
        RECT 33.140 125.875 35.170 126.045 ;
        RECT 35.340 125.705 35.510 126.845 ;
        RECT 35.680 125.875 36.015 126.845 ;
        RECT 37.235 126.950 37.520 127.280 ;
        RECT 37.235 126.805 37.405 126.950 ;
        RECT 36.740 126.635 37.405 126.805 ;
        RECT 37.690 126.780 37.860 127.580 ;
        RECT 36.740 125.875 36.910 126.635 ;
        RECT 37.090 125.705 37.420 126.465 ;
        RECT 37.590 125.875 37.860 126.780 ;
        RECT 38.035 127.515 38.290 128.085 ;
        RECT 38.460 127.855 38.790 128.255 ;
        RECT 39.215 127.720 39.745 128.085 ;
        RECT 39.215 127.685 39.390 127.720 ;
        RECT 38.460 127.515 39.390 127.685 ;
        RECT 39.935 127.575 40.210 128.085 ;
        RECT 38.035 126.845 38.205 127.515 ;
        RECT 38.460 127.345 38.630 127.515 ;
        RECT 38.375 127.015 38.630 127.345 ;
        RECT 38.855 127.015 39.050 127.345 ;
        RECT 38.035 125.875 38.370 126.845 ;
        RECT 38.540 125.705 38.710 126.845 ;
        RECT 38.880 126.045 39.050 127.015 ;
        RECT 39.220 126.385 39.390 127.515 ;
        RECT 39.560 126.725 39.730 127.525 ;
        RECT 39.930 127.405 40.210 127.575 ;
        RECT 39.935 126.925 40.210 127.405 ;
        RECT 40.380 126.725 40.570 128.085 ;
        RECT 40.750 127.720 41.260 128.255 ;
        RECT 41.480 127.445 41.725 128.050 ;
        RECT 42.830 127.625 43.160 127.985 ;
        RECT 43.780 127.795 44.030 128.255 ;
        RECT 44.200 127.795 44.760 128.085 ;
        RECT 40.770 127.275 42.000 127.445 ;
        RECT 42.830 127.435 44.220 127.625 ;
        RECT 39.560 126.555 40.570 126.725 ;
        RECT 40.740 126.710 41.490 126.900 ;
        RECT 39.220 126.215 40.345 126.385 ;
        RECT 40.740 126.045 40.910 126.710 ;
        RECT 41.660 126.465 42.000 127.275 ;
        RECT 44.050 127.345 44.220 127.435 ;
        RECT 42.645 127.015 43.320 127.265 ;
        RECT 43.540 127.015 43.880 127.265 ;
        RECT 44.050 127.015 44.340 127.345 ;
        RECT 42.645 126.655 42.910 127.015 ;
        RECT 44.050 126.765 44.220 127.015 ;
        RECT 38.880 125.875 40.910 126.045 ;
        RECT 41.080 125.705 41.250 126.465 ;
        RECT 41.485 126.055 42.000 126.465 ;
        RECT 43.280 126.595 44.220 126.765 ;
        RECT 42.830 125.705 43.110 126.375 ;
        RECT 43.280 126.045 43.580 126.595 ;
        RECT 44.510 126.425 44.760 127.795 ;
        RECT 43.780 125.705 44.110 126.425 ;
        RECT 44.300 125.875 44.760 126.425 ;
        RECT 44.930 127.580 45.200 127.925 ;
        RECT 45.390 127.855 45.770 128.255 ;
        RECT 45.940 127.685 46.110 128.035 ;
        RECT 46.280 127.855 46.610 128.255 ;
        RECT 46.810 127.685 46.980 128.035 ;
        RECT 47.180 127.755 47.510 128.255 ;
        RECT 44.930 126.845 45.100 127.580 ;
        RECT 45.370 127.515 46.980 127.685 ;
        RECT 45.370 127.345 45.540 127.515 ;
        RECT 45.270 127.015 45.540 127.345 ;
        RECT 45.710 127.015 46.115 127.345 ;
        RECT 45.370 126.845 45.540 127.015 ;
        RECT 44.930 125.875 45.200 126.845 ;
        RECT 45.370 126.675 46.095 126.845 ;
        RECT 46.285 126.725 46.995 127.345 ;
        RECT 47.165 127.015 47.515 127.585 ;
        RECT 47.690 127.530 47.980 128.255 ;
        RECT 49.130 127.775 49.410 128.255 ;
        RECT 49.580 127.605 49.840 127.995 ;
        RECT 50.015 127.775 50.270 128.255 ;
        RECT 50.440 127.605 50.735 127.995 ;
        RECT 50.915 127.775 51.190 128.255 ;
        RECT 51.360 127.755 51.660 128.085 ;
        RECT 49.085 127.435 50.735 127.605 ;
        RECT 49.085 126.925 49.490 127.435 ;
        RECT 49.660 127.095 50.800 127.265 ;
        RECT 45.925 126.555 46.095 126.675 ;
        RECT 47.195 126.555 47.515 126.845 ;
        RECT 45.410 125.705 45.690 126.505 ;
        RECT 45.925 126.385 47.515 126.555 ;
        RECT 45.860 125.925 47.515 126.215 ;
        RECT 47.690 125.705 47.980 126.870 ;
        RECT 49.085 126.755 49.840 126.925 ;
        RECT 49.125 125.705 49.410 126.575 ;
        RECT 49.580 126.505 49.840 126.755 ;
        RECT 50.630 126.845 50.800 127.095 ;
        RECT 50.970 127.015 51.320 127.585 ;
        RECT 51.490 126.845 51.660 127.755 ;
        RECT 50.630 126.675 51.660 126.845 ;
        RECT 49.580 126.335 50.700 126.505 ;
        RECT 49.580 125.875 49.840 126.335 ;
        RECT 50.015 125.705 50.270 126.165 ;
        RECT 50.440 125.875 50.700 126.335 ;
        RECT 50.870 125.705 51.180 126.505 ;
        RECT 51.350 125.875 51.660 126.675 ;
        RECT 51.830 127.455 52.170 128.085 ;
        RECT 52.340 127.455 52.590 128.255 ;
        RECT 52.780 127.605 53.110 128.085 ;
        RECT 53.280 127.795 53.505 128.255 ;
        RECT 53.675 127.605 54.005 128.085 ;
        RECT 51.830 126.895 52.005 127.455 ;
        RECT 52.780 127.435 54.005 127.605 ;
        RECT 54.635 127.475 55.135 128.085 ;
        RECT 55.885 127.915 56.140 128.075 ;
        RECT 55.800 127.745 56.140 127.915 ;
        RECT 56.320 127.795 56.605 128.255 ;
        RECT 55.885 127.545 56.140 127.745 ;
        RECT 52.175 127.095 52.870 127.265 ;
        RECT 51.830 126.845 52.060 126.895 ;
        RECT 52.700 126.845 52.870 127.095 ;
        RECT 53.045 127.065 53.465 127.265 ;
        RECT 53.635 127.065 53.965 127.265 ;
        RECT 54.135 127.065 54.465 127.265 ;
        RECT 54.635 126.845 54.805 127.475 ;
        RECT 54.990 127.015 55.340 127.265 ;
        RECT 51.830 125.875 52.170 126.845 ;
        RECT 52.340 125.705 52.510 126.845 ;
        RECT 52.700 126.675 55.135 126.845 ;
        RECT 52.780 125.705 53.030 126.505 ;
        RECT 53.675 125.875 54.005 126.675 ;
        RECT 54.305 125.705 54.635 126.505 ;
        RECT 54.805 125.875 55.135 126.675 ;
        RECT 55.885 126.685 56.065 127.545 ;
        RECT 56.785 127.345 57.035 127.995 ;
        RECT 56.235 127.015 57.035 127.345 ;
        RECT 55.885 126.015 56.140 126.685 ;
        RECT 56.320 125.705 56.605 126.505 ;
        RECT 56.785 126.425 57.035 127.015 ;
        RECT 57.235 127.660 57.555 127.990 ;
        RECT 57.735 127.775 58.395 128.255 ;
        RECT 58.595 127.865 59.445 128.035 ;
        RECT 57.235 126.765 57.425 127.660 ;
        RECT 57.745 127.335 58.405 127.605 ;
        RECT 58.075 127.275 58.405 127.335 ;
        RECT 57.595 127.105 57.925 127.165 ;
        RECT 58.595 127.105 58.765 127.865 ;
        RECT 60.005 127.795 60.325 128.255 ;
        RECT 60.525 127.615 60.775 128.045 ;
        RECT 61.065 127.815 61.475 128.255 ;
        RECT 61.645 127.875 62.660 128.075 ;
        RECT 58.935 127.445 60.185 127.615 ;
        RECT 58.935 127.325 59.265 127.445 ;
        RECT 57.595 126.935 59.495 127.105 ;
        RECT 57.235 126.595 59.155 126.765 ;
        RECT 57.235 126.575 57.555 126.595 ;
        RECT 56.785 125.915 57.115 126.425 ;
        RECT 57.385 125.965 57.555 126.575 ;
        RECT 59.325 126.425 59.495 126.935 ;
        RECT 59.665 126.865 59.845 127.275 ;
        RECT 60.015 126.685 60.185 127.445 ;
        RECT 57.725 125.705 58.055 126.395 ;
        RECT 58.285 126.255 59.495 126.425 ;
        RECT 59.665 126.375 60.185 126.685 ;
        RECT 60.355 127.275 60.775 127.615 ;
        RECT 61.065 127.275 61.475 127.605 ;
        RECT 60.355 126.505 60.545 127.275 ;
        RECT 61.645 127.145 61.815 127.875 ;
        RECT 62.960 127.705 63.130 128.035 ;
        RECT 63.300 127.875 63.630 128.255 ;
        RECT 61.985 127.325 62.335 127.695 ;
        RECT 61.645 127.105 62.065 127.145 ;
        RECT 60.715 126.935 62.065 127.105 ;
        RECT 60.715 126.775 60.965 126.935 ;
        RECT 61.475 126.505 61.725 126.765 ;
        RECT 60.355 126.255 61.725 126.505 ;
        RECT 58.285 125.965 58.525 126.255 ;
        RECT 59.325 126.175 59.495 126.255 ;
        RECT 58.725 125.705 59.145 126.085 ;
        RECT 59.325 125.925 59.955 126.175 ;
        RECT 60.425 125.705 60.755 126.085 ;
        RECT 60.925 125.965 61.095 126.255 ;
        RECT 61.895 126.090 62.065 126.935 ;
        RECT 62.515 126.765 62.735 127.635 ;
        RECT 62.960 127.515 63.655 127.705 ;
        RECT 62.235 126.385 62.735 126.765 ;
        RECT 62.905 126.715 63.315 127.335 ;
        RECT 63.485 126.545 63.655 127.515 ;
        RECT 62.960 126.375 63.655 126.545 ;
        RECT 61.275 125.705 61.655 126.085 ;
        RECT 61.895 125.920 62.725 126.090 ;
        RECT 62.960 125.875 63.130 126.375 ;
        RECT 63.300 125.705 63.630 126.205 ;
        RECT 63.845 125.875 64.070 127.995 ;
        RECT 64.240 127.875 64.570 128.255 ;
        RECT 64.740 127.705 64.910 127.995 ;
        RECT 64.245 127.535 64.910 127.705 ;
        RECT 65.170 127.755 65.430 128.085 ;
        RECT 65.640 127.775 65.915 128.255 ;
        RECT 64.245 126.545 64.475 127.535 ;
        RECT 64.645 126.715 64.995 127.365 ;
        RECT 65.170 126.845 65.340 127.755 ;
        RECT 66.125 127.685 66.330 128.085 ;
        RECT 66.500 127.855 66.835 128.255 ;
        RECT 65.510 127.015 65.870 127.595 ;
        RECT 66.125 127.515 66.810 127.685 ;
        RECT 66.050 126.845 66.300 127.345 ;
        RECT 65.170 126.675 66.300 126.845 ;
        RECT 64.245 126.375 64.910 126.545 ;
        RECT 64.240 125.705 64.570 126.205 ;
        RECT 64.740 125.875 64.910 126.375 ;
        RECT 65.170 125.905 65.440 126.675 ;
        RECT 66.470 126.485 66.810 127.515 ;
        RECT 65.610 125.705 65.940 126.485 ;
        RECT 66.145 126.310 66.810 126.485 ;
        RECT 67.010 127.580 67.280 127.925 ;
        RECT 67.470 127.855 67.850 128.255 ;
        RECT 68.020 127.685 68.190 128.035 ;
        RECT 68.360 127.855 68.690 128.255 ;
        RECT 68.890 127.685 69.060 128.035 ;
        RECT 69.260 127.755 69.590 128.255 ;
        RECT 67.010 126.845 67.180 127.580 ;
        RECT 67.450 127.515 69.060 127.685 ;
        RECT 67.450 127.345 67.620 127.515 ;
        RECT 67.350 127.015 67.620 127.345 ;
        RECT 67.790 127.015 68.195 127.345 ;
        RECT 67.450 126.845 67.620 127.015 ;
        RECT 68.365 126.895 69.075 127.345 ;
        RECT 69.245 127.015 69.595 127.585 ;
        RECT 69.770 127.455 70.110 128.085 ;
        RECT 70.280 127.455 70.530 128.255 ;
        RECT 70.720 127.605 71.050 128.085 ;
        RECT 71.220 127.795 71.445 128.255 ;
        RECT 71.615 127.605 71.945 128.085 ;
        RECT 66.145 125.905 66.330 126.310 ;
        RECT 66.500 125.705 66.835 126.130 ;
        RECT 67.010 125.875 67.280 126.845 ;
        RECT 67.450 126.675 68.175 126.845 ;
        RECT 68.365 126.725 69.080 126.895 ;
        RECT 69.770 126.845 69.945 127.455 ;
        RECT 70.720 127.435 71.945 127.605 ;
        RECT 72.575 127.475 73.075 128.085 ;
        RECT 73.450 127.530 73.740 128.255 ;
        RECT 74.830 127.795 75.390 128.085 ;
        RECT 75.560 127.795 75.810 128.255 ;
        RECT 70.115 127.095 70.810 127.265 ;
        RECT 70.640 126.845 70.810 127.095 ;
        RECT 70.985 127.065 71.405 127.265 ;
        RECT 71.575 127.065 71.905 127.265 ;
        RECT 72.075 127.065 72.405 127.265 ;
        RECT 72.575 126.845 72.745 127.475 ;
        RECT 72.930 127.015 73.280 127.265 ;
        RECT 68.005 126.555 68.175 126.675 ;
        RECT 69.275 126.555 69.595 126.845 ;
        RECT 67.490 125.705 67.770 126.505 ;
        RECT 68.005 126.385 69.595 126.555 ;
        RECT 67.940 125.925 69.595 126.215 ;
        RECT 69.770 125.875 70.110 126.845 ;
        RECT 70.280 125.705 70.450 126.845 ;
        RECT 70.640 126.675 73.075 126.845 ;
        RECT 70.720 125.705 70.970 126.505 ;
        RECT 71.615 125.875 71.945 126.675 ;
        RECT 72.245 125.705 72.575 126.505 ;
        RECT 72.745 125.875 73.075 126.675 ;
        RECT 73.450 125.705 73.740 126.870 ;
        RECT 74.830 126.425 75.080 127.795 ;
        RECT 76.430 127.625 76.760 127.985 ;
        RECT 75.370 127.435 76.760 127.625 ;
        RECT 77.405 127.445 77.650 128.050 ;
        RECT 77.870 127.720 78.380 128.255 ;
        RECT 75.370 127.345 75.540 127.435 ;
        RECT 75.250 127.015 75.540 127.345 ;
        RECT 77.130 127.275 78.360 127.445 ;
        RECT 75.710 127.015 76.050 127.265 ;
        RECT 76.270 127.015 76.945 127.265 ;
        RECT 75.370 126.765 75.540 127.015 ;
        RECT 75.370 126.595 76.310 126.765 ;
        RECT 76.680 126.655 76.945 127.015 ;
        RECT 74.830 125.875 75.290 126.425 ;
        RECT 75.480 125.705 75.810 126.425 ;
        RECT 76.010 126.045 76.310 126.595 ;
        RECT 77.130 126.465 77.470 127.275 ;
        RECT 77.640 126.710 78.390 126.900 ;
        RECT 76.480 125.705 76.760 126.375 ;
        RECT 77.130 126.055 77.645 126.465 ;
        RECT 77.880 125.705 78.050 126.465 ;
        RECT 78.220 126.045 78.390 126.710 ;
        RECT 78.560 126.725 78.750 128.085 ;
        RECT 78.920 127.575 79.195 128.085 ;
        RECT 79.385 127.720 79.915 128.085 ;
        RECT 80.340 127.855 80.670 128.255 ;
        RECT 79.740 127.685 79.915 127.720 ;
        RECT 78.920 127.405 79.200 127.575 ;
        RECT 78.920 126.925 79.195 127.405 ;
        RECT 79.400 126.725 79.570 127.525 ;
        RECT 78.560 126.555 79.570 126.725 ;
        RECT 79.740 127.515 80.670 127.685 ;
        RECT 80.840 127.515 81.095 128.085 ;
        RECT 81.730 127.745 82.035 128.255 ;
        RECT 79.740 126.385 79.910 127.515 ;
        RECT 80.500 127.345 80.670 127.515 ;
        RECT 78.785 126.215 79.910 126.385 ;
        RECT 80.080 127.015 80.275 127.345 ;
        RECT 80.500 127.015 80.755 127.345 ;
        RECT 80.080 126.045 80.250 127.015 ;
        RECT 80.925 126.845 81.095 127.515 ;
        RECT 81.730 127.015 82.045 127.575 ;
        RECT 82.215 127.265 82.465 128.075 ;
        RECT 82.635 127.730 82.895 128.255 ;
        RECT 83.075 127.265 83.325 128.075 ;
        RECT 83.495 127.695 83.755 128.255 ;
        RECT 83.925 127.605 84.185 128.060 ;
        RECT 84.355 127.775 84.615 128.255 ;
        RECT 84.785 127.605 85.045 128.060 ;
        RECT 85.215 127.775 85.475 128.255 ;
        RECT 85.645 127.605 85.905 128.060 ;
        RECT 86.075 127.775 86.320 128.255 ;
        RECT 86.490 127.605 86.765 128.060 ;
        RECT 86.935 127.775 87.180 128.255 ;
        RECT 87.350 127.605 87.610 128.060 ;
        RECT 87.790 127.775 88.040 128.255 ;
        RECT 88.210 127.605 88.470 128.060 ;
        RECT 88.650 127.775 88.900 128.255 ;
        RECT 89.070 127.605 89.330 128.060 ;
        RECT 89.510 127.775 89.770 128.255 ;
        RECT 89.940 127.605 90.200 128.060 ;
        RECT 90.370 127.775 90.670 128.255 ;
        RECT 83.925 127.435 90.670 127.605 ;
        RECT 82.215 127.015 89.335 127.265 ;
        RECT 78.220 125.875 80.250 126.045 ;
        RECT 80.420 125.705 80.590 126.845 ;
        RECT 80.760 125.875 81.095 126.845 ;
        RECT 81.740 125.705 82.035 126.515 ;
        RECT 82.215 125.875 82.460 127.015 ;
        RECT 82.635 125.705 82.895 126.515 ;
        RECT 83.075 125.880 83.325 127.015 ;
        RECT 89.505 126.845 90.670 127.435 ;
        RECT 83.925 126.620 90.670 126.845 ;
        RECT 90.930 127.580 91.190 128.085 ;
        RECT 91.370 127.875 91.700 128.255 ;
        RECT 91.880 127.705 92.050 128.085 ;
        RECT 90.930 126.780 91.100 127.580 ;
        RECT 91.385 127.535 92.050 127.705 ;
        RECT 91.385 127.280 91.555 127.535 ;
        RECT 92.770 127.485 94.440 128.255 ;
        RECT 91.270 126.950 91.555 127.280 ;
        RECT 91.790 126.985 92.120 127.355 ;
        RECT 91.385 126.805 91.555 126.950 ;
        RECT 83.925 126.605 89.330 126.620 ;
        RECT 83.495 125.710 83.755 126.505 ;
        RECT 83.925 125.880 84.185 126.605 ;
        RECT 84.355 125.710 84.615 126.435 ;
        RECT 84.785 125.880 85.045 126.605 ;
        RECT 85.215 125.710 85.475 126.435 ;
        RECT 85.645 125.880 85.905 126.605 ;
        RECT 86.075 125.710 86.335 126.435 ;
        RECT 86.505 125.880 86.765 126.605 ;
        RECT 86.935 125.710 87.180 126.435 ;
        RECT 87.350 125.880 87.610 126.605 ;
        RECT 87.795 125.710 88.040 126.435 ;
        RECT 88.210 125.880 88.470 126.605 ;
        RECT 88.655 125.710 88.900 126.435 ;
        RECT 89.070 125.880 89.330 126.605 ;
        RECT 89.515 125.710 89.770 126.435 ;
        RECT 89.940 125.880 90.230 126.620 ;
        RECT 83.495 125.705 89.770 125.710 ;
        RECT 90.400 125.705 90.670 126.450 ;
        RECT 90.930 125.875 91.200 126.780 ;
        RECT 91.385 126.635 92.050 126.805 ;
        RECT 91.370 125.705 91.700 126.465 ;
        RECT 91.880 125.875 92.050 126.635 ;
        RECT 92.770 126.795 93.520 127.315 ;
        RECT 93.690 126.965 94.440 127.485 ;
        RECT 94.810 127.625 95.140 127.985 ;
        RECT 95.760 127.795 96.010 128.255 ;
        RECT 96.180 127.795 96.740 128.085 ;
        RECT 94.810 127.435 96.200 127.625 ;
        RECT 96.030 127.345 96.200 127.435 ;
        RECT 94.625 127.015 95.300 127.265 ;
        RECT 95.520 127.015 95.860 127.265 ;
        RECT 96.030 127.015 96.320 127.345 ;
        RECT 92.770 125.705 94.440 126.795 ;
        RECT 94.625 126.655 94.890 127.015 ;
        RECT 96.030 126.765 96.200 127.015 ;
        RECT 95.260 126.595 96.200 126.765 ;
        RECT 94.810 125.705 95.090 126.375 ;
        RECT 95.260 126.045 95.560 126.595 ;
        RECT 96.490 126.425 96.740 127.795 ;
        RECT 97.110 127.625 97.440 127.985 ;
        RECT 98.060 127.795 98.310 128.255 ;
        RECT 98.480 127.795 99.040 128.085 ;
        RECT 97.110 127.435 98.500 127.625 ;
        RECT 98.330 127.345 98.500 127.435 ;
        RECT 96.925 127.015 97.600 127.265 ;
        RECT 97.820 127.015 98.160 127.265 ;
        RECT 98.330 127.015 98.620 127.345 ;
        RECT 96.925 126.655 97.190 127.015 ;
        RECT 98.330 126.765 98.500 127.015 ;
        RECT 95.760 125.705 96.090 126.425 ;
        RECT 96.280 125.875 96.740 126.425 ;
        RECT 97.560 126.595 98.500 126.765 ;
        RECT 97.110 125.705 97.390 126.375 ;
        RECT 97.560 126.045 97.860 126.595 ;
        RECT 98.790 126.425 99.040 127.795 ;
        RECT 99.210 127.530 99.500 128.255 ;
        RECT 99.670 127.505 100.880 128.255 ;
        RECT 98.060 125.705 98.390 126.425 ;
        RECT 98.580 125.875 99.040 126.425 ;
        RECT 99.210 125.705 99.500 126.870 ;
        RECT 99.670 126.795 100.190 127.335 ;
        RECT 100.360 126.965 100.880 127.505 ;
        RECT 101.050 127.485 104.560 128.255 ;
        RECT 101.050 126.795 102.740 127.315 ;
        RECT 102.910 126.965 104.560 127.485 ;
        RECT 104.770 127.435 105.000 128.255 ;
        RECT 105.170 127.455 105.500 128.085 ;
        RECT 104.750 127.015 105.080 127.265 ;
        RECT 105.250 126.855 105.500 127.455 ;
        RECT 105.670 127.435 105.880 128.255 ;
        RECT 107.120 127.705 107.290 128.085 ;
        RECT 107.470 127.875 107.800 128.255 ;
        RECT 107.120 127.535 107.785 127.705 ;
        RECT 107.980 127.580 108.240 128.085 ;
        RECT 107.050 126.985 107.380 127.355 ;
        RECT 107.615 127.280 107.785 127.535 ;
        RECT 99.670 125.705 100.880 126.795 ;
        RECT 101.050 125.705 104.560 126.795 ;
        RECT 104.770 125.705 105.000 126.845 ;
        RECT 105.170 125.875 105.500 126.855 ;
        RECT 107.615 126.950 107.900 127.280 ;
        RECT 105.670 125.705 105.880 126.845 ;
        RECT 107.615 126.805 107.785 126.950 ;
        RECT 107.120 126.635 107.785 126.805 ;
        RECT 108.070 126.780 108.240 127.580 ;
        RECT 108.410 127.485 111.000 128.255 ;
        RECT 111.170 127.505 112.380 128.255 ;
        RECT 107.120 125.875 107.290 126.635 ;
        RECT 107.470 125.705 107.800 126.465 ;
        RECT 107.970 125.875 108.240 126.780 ;
        RECT 108.410 126.795 109.620 127.315 ;
        RECT 109.790 126.965 111.000 127.485 ;
        RECT 111.170 126.795 111.690 127.335 ;
        RECT 111.860 126.965 112.380 127.505 ;
        RECT 108.410 125.705 111.000 126.795 ;
        RECT 111.170 125.705 112.380 126.795 ;
        RECT 18.165 125.535 112.465 125.705 ;
        RECT 18.250 124.445 19.460 125.535 ;
        RECT 18.250 123.735 18.770 124.275 ;
        RECT 18.940 123.905 19.460 124.445 ;
        RECT 19.720 124.605 19.890 125.365 ;
        RECT 20.070 124.775 20.400 125.535 ;
        RECT 19.720 124.435 20.385 124.605 ;
        RECT 20.570 124.460 20.840 125.365 ;
        RECT 20.215 124.290 20.385 124.435 ;
        RECT 19.650 123.885 19.980 124.255 ;
        RECT 20.215 123.960 20.500 124.290 ;
        RECT 18.250 122.985 19.460 123.735 ;
        RECT 20.215 123.705 20.385 123.960 ;
        RECT 19.720 123.535 20.385 123.705 ;
        RECT 20.670 123.660 20.840 124.460 ;
        RECT 19.720 123.155 19.890 123.535 ;
        RECT 20.070 122.985 20.400 123.365 ;
        RECT 20.580 123.155 20.840 123.660 ;
        RECT 21.015 124.395 21.350 125.365 ;
        RECT 21.520 124.395 21.690 125.535 ;
        RECT 21.860 125.195 23.890 125.365 ;
        RECT 21.015 123.725 21.185 124.395 ;
        RECT 21.860 124.225 22.030 125.195 ;
        RECT 21.355 123.895 21.610 124.225 ;
        RECT 21.835 123.895 22.030 124.225 ;
        RECT 22.200 124.855 23.325 125.025 ;
        RECT 21.440 123.725 21.610 123.895 ;
        RECT 22.200 123.725 22.370 124.855 ;
        RECT 21.015 123.155 21.270 123.725 ;
        RECT 21.440 123.555 22.370 123.725 ;
        RECT 22.540 124.515 23.550 124.685 ;
        RECT 22.540 123.715 22.710 124.515 ;
        RECT 22.915 124.175 23.190 124.315 ;
        RECT 22.910 124.005 23.190 124.175 ;
        RECT 22.195 123.520 22.370 123.555 ;
        RECT 21.440 122.985 21.770 123.385 ;
        RECT 22.195 123.155 22.725 123.520 ;
        RECT 22.915 123.155 23.190 124.005 ;
        RECT 23.360 123.155 23.550 124.515 ;
        RECT 23.720 124.530 23.890 125.195 ;
        RECT 24.060 124.775 24.230 125.535 ;
        RECT 25.525 125.195 25.780 125.225 ;
        RECT 24.465 124.775 24.980 125.185 ;
        RECT 25.440 125.025 25.780 125.195 ;
        RECT 23.720 124.340 24.470 124.530 ;
        RECT 24.640 123.965 24.980 124.775 ;
        RECT 23.750 123.795 24.980 123.965 ;
        RECT 25.525 124.555 25.780 125.025 ;
        RECT 25.960 124.735 26.245 125.535 ;
        RECT 26.425 124.815 26.755 125.325 ;
        RECT 23.730 122.985 24.240 123.520 ;
        RECT 24.460 123.190 24.705 123.795 ;
        RECT 25.525 123.695 25.705 124.555 ;
        RECT 26.425 124.225 26.675 124.815 ;
        RECT 27.025 124.665 27.195 125.275 ;
        RECT 27.365 124.845 27.695 125.535 ;
        RECT 27.925 124.985 28.165 125.275 ;
        RECT 28.365 125.155 28.785 125.535 ;
        RECT 28.965 125.065 29.595 125.315 ;
        RECT 30.065 125.155 30.395 125.535 ;
        RECT 28.965 124.985 29.135 125.065 ;
        RECT 30.565 124.985 30.735 125.275 ;
        RECT 30.915 125.155 31.295 125.535 ;
        RECT 31.535 125.150 32.365 125.320 ;
        RECT 27.925 124.815 29.135 124.985 ;
        RECT 25.875 123.895 26.675 124.225 ;
        RECT 25.525 123.165 25.780 123.695 ;
        RECT 25.960 122.985 26.245 123.445 ;
        RECT 26.425 123.245 26.675 123.895 ;
        RECT 26.875 124.645 27.195 124.665 ;
        RECT 26.875 124.475 28.795 124.645 ;
        RECT 26.875 123.580 27.065 124.475 ;
        RECT 28.965 124.305 29.135 124.815 ;
        RECT 29.305 124.555 29.825 124.865 ;
        RECT 27.235 124.135 29.135 124.305 ;
        RECT 27.235 124.075 27.565 124.135 ;
        RECT 27.715 123.905 28.045 123.965 ;
        RECT 27.385 123.635 28.045 123.905 ;
        RECT 26.875 123.250 27.195 123.580 ;
        RECT 27.375 122.985 28.035 123.465 ;
        RECT 28.235 123.375 28.405 124.135 ;
        RECT 29.305 123.965 29.485 124.375 ;
        RECT 28.575 123.795 28.905 123.915 ;
        RECT 29.655 123.795 29.825 124.555 ;
        RECT 28.575 123.625 29.825 123.795 ;
        RECT 29.995 124.735 31.365 124.985 ;
        RECT 29.995 123.965 30.185 124.735 ;
        RECT 31.115 124.475 31.365 124.735 ;
        RECT 30.355 124.305 30.605 124.465 ;
        RECT 31.535 124.305 31.705 125.150 ;
        RECT 32.600 124.865 32.770 125.365 ;
        RECT 32.940 125.035 33.270 125.535 ;
        RECT 31.875 124.475 32.375 124.855 ;
        RECT 32.600 124.695 33.295 124.865 ;
        RECT 30.355 124.135 31.705 124.305 ;
        RECT 31.285 124.095 31.705 124.135 ;
        RECT 29.995 123.625 30.415 123.965 ;
        RECT 30.705 123.635 31.115 123.965 ;
        RECT 28.235 123.205 29.085 123.375 ;
        RECT 29.645 122.985 29.965 123.445 ;
        RECT 30.165 123.195 30.415 123.625 ;
        RECT 30.705 122.985 31.115 123.425 ;
        RECT 31.285 123.365 31.455 124.095 ;
        RECT 31.625 123.545 31.975 123.915 ;
        RECT 32.155 123.605 32.375 124.475 ;
        RECT 32.545 123.905 32.955 124.525 ;
        RECT 33.125 123.725 33.295 124.695 ;
        RECT 32.600 123.535 33.295 123.725 ;
        RECT 31.285 123.165 32.300 123.365 ;
        RECT 32.600 123.205 32.770 123.535 ;
        RECT 32.940 122.985 33.270 123.365 ;
        RECT 33.485 123.245 33.710 125.365 ;
        RECT 33.880 125.035 34.210 125.535 ;
        RECT 34.380 124.865 34.550 125.365 ;
        RECT 33.885 124.695 34.550 124.865 ;
        RECT 33.885 123.705 34.115 124.695 ;
        RECT 34.285 123.875 34.635 124.525 ;
        RECT 34.810 124.370 35.100 125.535 ;
        RECT 35.360 124.790 35.630 125.535 ;
        RECT 36.260 125.530 42.535 125.535 ;
        RECT 35.800 124.620 36.090 125.360 ;
        RECT 36.260 124.805 36.515 125.530 ;
        RECT 36.700 124.635 36.960 125.360 ;
        RECT 37.130 124.805 37.375 125.530 ;
        RECT 37.560 124.635 37.820 125.360 ;
        RECT 37.990 124.805 38.235 125.530 ;
        RECT 38.420 124.635 38.680 125.360 ;
        RECT 38.850 124.805 39.095 125.530 ;
        RECT 39.265 124.635 39.525 125.360 ;
        RECT 39.695 124.805 39.955 125.530 ;
        RECT 40.125 124.635 40.385 125.360 ;
        RECT 40.555 124.805 40.815 125.530 ;
        RECT 40.985 124.635 41.245 125.360 ;
        RECT 41.415 124.805 41.675 125.530 ;
        RECT 41.845 124.635 42.105 125.360 ;
        RECT 42.275 124.735 42.535 125.530 ;
        RECT 36.700 124.620 42.105 124.635 ;
        RECT 35.360 124.395 42.105 124.620 ;
        RECT 35.360 123.805 36.525 124.395 ;
        RECT 42.705 124.225 42.955 125.360 ;
        RECT 43.135 124.725 43.395 125.535 ;
        RECT 43.570 124.225 43.815 125.365 ;
        RECT 43.995 124.725 44.290 125.535 ;
        RECT 44.470 124.815 44.930 125.365 ;
        RECT 45.120 124.815 45.450 125.535 ;
        RECT 36.695 123.975 43.815 124.225 ;
        RECT 33.885 123.535 34.550 123.705 ;
        RECT 33.880 122.985 34.210 123.365 ;
        RECT 34.380 123.245 34.550 123.535 ;
        RECT 34.810 122.985 35.100 123.710 ;
        RECT 35.360 123.635 42.105 123.805 ;
        RECT 35.360 122.985 35.660 123.465 ;
        RECT 35.830 123.180 36.090 123.635 ;
        RECT 36.260 122.985 36.520 123.465 ;
        RECT 36.700 123.180 36.960 123.635 ;
        RECT 37.130 122.985 37.380 123.465 ;
        RECT 37.560 123.180 37.820 123.635 ;
        RECT 37.990 122.985 38.240 123.465 ;
        RECT 38.420 123.180 38.680 123.635 ;
        RECT 38.850 122.985 39.095 123.465 ;
        RECT 39.265 123.180 39.540 123.635 ;
        RECT 39.710 122.985 39.955 123.465 ;
        RECT 40.125 123.180 40.385 123.635 ;
        RECT 40.555 122.985 40.815 123.465 ;
        RECT 40.985 123.180 41.245 123.635 ;
        RECT 41.415 122.985 41.675 123.465 ;
        RECT 41.845 123.180 42.105 123.635 ;
        RECT 42.275 122.985 42.535 123.545 ;
        RECT 42.705 123.165 42.955 123.975 ;
        RECT 43.135 122.985 43.395 123.510 ;
        RECT 43.565 123.165 43.815 123.975 ;
        RECT 43.985 123.665 44.300 124.225 ;
        RECT 43.995 122.985 44.300 123.495 ;
        RECT 44.470 123.445 44.720 124.815 ;
        RECT 45.650 124.645 45.950 125.195 ;
        RECT 46.120 124.865 46.400 125.535 ;
        RECT 45.010 124.475 45.950 124.645 ;
        RECT 46.770 124.815 47.230 125.365 ;
        RECT 47.420 124.815 47.750 125.535 ;
        RECT 45.010 124.225 45.180 124.475 ;
        RECT 46.320 124.225 46.585 124.585 ;
        RECT 44.890 123.895 45.180 124.225 ;
        RECT 45.350 123.975 45.690 124.225 ;
        RECT 45.910 123.975 46.585 124.225 ;
        RECT 45.010 123.805 45.180 123.895 ;
        RECT 45.010 123.615 46.400 123.805 ;
        RECT 44.470 123.155 45.030 123.445 ;
        RECT 45.200 122.985 45.450 123.445 ;
        RECT 46.070 123.255 46.400 123.615 ;
        RECT 46.770 123.445 47.020 124.815 ;
        RECT 47.950 124.645 48.250 125.195 ;
        RECT 48.420 124.865 48.700 125.535 ;
        RECT 47.310 124.475 48.250 124.645 ;
        RECT 47.310 124.225 47.480 124.475 ;
        RECT 48.620 124.225 48.885 124.585 ;
        RECT 47.190 123.895 47.480 124.225 ;
        RECT 47.650 123.975 47.990 124.225 ;
        RECT 48.210 123.975 48.885 124.225 ;
        RECT 49.075 124.395 49.410 125.365 ;
        RECT 49.580 124.395 49.750 125.535 ;
        RECT 49.920 125.195 51.950 125.365 ;
        RECT 47.310 123.805 47.480 123.895 ;
        RECT 47.310 123.615 48.700 123.805 ;
        RECT 46.770 123.155 47.330 123.445 ;
        RECT 47.500 122.985 47.750 123.445 ;
        RECT 48.370 123.255 48.700 123.615 ;
        RECT 49.075 123.725 49.245 124.395 ;
        RECT 49.920 124.225 50.090 125.195 ;
        RECT 49.415 123.895 49.670 124.225 ;
        RECT 49.895 123.895 50.090 124.225 ;
        RECT 50.260 124.855 51.385 125.025 ;
        RECT 49.500 123.725 49.670 123.895 ;
        RECT 50.260 123.725 50.430 124.855 ;
        RECT 49.075 123.155 49.330 123.725 ;
        RECT 49.500 123.555 50.430 123.725 ;
        RECT 50.600 124.515 51.610 124.685 ;
        RECT 50.600 123.715 50.770 124.515 ;
        RECT 50.255 123.520 50.430 123.555 ;
        RECT 49.500 122.985 49.830 123.385 ;
        RECT 50.255 123.155 50.785 123.520 ;
        RECT 50.975 123.495 51.250 124.315 ;
        RECT 50.970 123.325 51.250 123.495 ;
        RECT 50.975 123.155 51.250 123.325 ;
        RECT 51.420 123.155 51.610 124.515 ;
        RECT 51.780 124.530 51.950 125.195 ;
        RECT 52.120 124.775 52.290 125.535 ;
        RECT 52.525 124.775 53.040 125.185 ;
        RECT 53.310 125.075 53.480 125.535 ;
        RECT 51.780 124.340 52.530 124.530 ;
        RECT 52.700 123.965 53.040 124.775 ;
        RECT 53.650 124.585 53.980 125.365 ;
        RECT 54.150 124.735 54.320 125.535 ;
        RECT 51.810 123.795 53.040 123.965 ;
        RECT 53.210 124.565 53.980 124.585 ;
        RECT 54.490 124.565 54.820 125.365 ;
        RECT 54.990 124.735 55.160 125.535 ;
        RECT 55.330 124.565 55.660 125.365 ;
        RECT 53.210 124.395 55.660 124.565 ;
        RECT 55.920 124.395 56.215 125.535 ;
        RECT 56.435 124.395 56.770 125.365 ;
        RECT 56.940 124.395 57.110 125.535 ;
        RECT 57.280 125.195 59.310 125.365 ;
        RECT 53.210 123.805 53.560 124.395 ;
        RECT 53.730 123.975 56.240 124.225 ;
        RECT 51.790 122.985 52.300 123.520 ;
        RECT 52.520 123.190 52.765 123.795 ;
        RECT 53.210 123.625 55.580 123.805 ;
        RECT 53.310 122.985 53.560 123.450 ;
        RECT 53.730 123.155 53.900 123.625 ;
        RECT 54.150 122.985 54.320 123.445 ;
        RECT 54.570 123.155 54.740 123.625 ;
        RECT 54.990 122.985 55.160 123.445 ;
        RECT 55.410 123.155 55.580 123.625 ;
        RECT 56.435 123.725 56.605 124.395 ;
        RECT 57.280 124.225 57.450 125.195 ;
        RECT 56.775 123.895 57.030 124.225 ;
        RECT 57.255 123.895 57.450 124.225 ;
        RECT 57.620 124.855 58.745 125.025 ;
        RECT 56.860 123.725 57.030 123.895 ;
        RECT 57.620 123.725 57.790 124.855 ;
        RECT 55.950 122.985 56.215 123.445 ;
        RECT 56.435 123.155 56.690 123.725 ;
        RECT 56.860 123.555 57.790 123.725 ;
        RECT 57.960 124.515 58.970 124.685 ;
        RECT 57.960 123.715 58.130 124.515 ;
        RECT 58.335 124.175 58.610 124.315 ;
        RECT 58.330 124.005 58.610 124.175 ;
        RECT 57.615 123.520 57.790 123.555 ;
        RECT 56.860 122.985 57.190 123.385 ;
        RECT 57.615 123.155 58.145 123.520 ;
        RECT 58.335 123.155 58.610 124.005 ;
        RECT 58.780 123.155 58.970 124.515 ;
        RECT 59.140 124.530 59.310 125.195 ;
        RECT 59.480 124.775 59.650 125.535 ;
        RECT 59.885 124.775 60.400 125.185 ;
        RECT 59.140 124.340 59.890 124.530 ;
        RECT 60.060 123.965 60.400 124.775 ;
        RECT 60.570 124.370 60.860 125.535 ;
        RECT 61.490 124.815 61.950 125.365 ;
        RECT 62.140 124.815 62.470 125.535 ;
        RECT 59.170 123.795 60.400 123.965 ;
        RECT 59.150 122.985 59.660 123.520 ;
        RECT 59.880 123.190 60.125 123.795 ;
        RECT 60.570 122.985 60.860 123.710 ;
        RECT 61.490 123.445 61.740 124.815 ;
        RECT 62.670 124.645 62.970 125.195 ;
        RECT 63.140 124.865 63.420 125.535 ;
        RECT 63.990 124.865 64.270 125.535 ;
        RECT 62.030 124.475 62.970 124.645 ;
        RECT 64.440 124.645 64.740 125.195 ;
        RECT 64.940 124.815 65.270 125.535 ;
        RECT 65.460 124.815 65.920 125.365 ;
        RECT 62.030 124.225 62.200 124.475 ;
        RECT 63.340 124.225 63.605 124.585 ;
        RECT 61.910 123.895 62.200 124.225 ;
        RECT 62.370 123.975 62.710 124.225 ;
        RECT 62.930 123.975 63.605 124.225 ;
        RECT 63.805 124.225 64.070 124.585 ;
        RECT 64.440 124.475 65.380 124.645 ;
        RECT 65.210 124.225 65.380 124.475 ;
        RECT 63.805 123.975 64.480 124.225 ;
        RECT 64.700 123.975 65.040 124.225 ;
        RECT 62.030 123.805 62.200 123.895 ;
        RECT 65.210 123.895 65.500 124.225 ;
        RECT 65.210 123.805 65.380 123.895 ;
        RECT 62.030 123.615 63.420 123.805 ;
        RECT 61.490 123.155 62.050 123.445 ;
        RECT 62.220 122.985 62.470 123.445 ;
        RECT 63.090 123.255 63.420 123.615 ;
        RECT 63.990 123.615 65.380 123.805 ;
        RECT 63.990 123.255 64.320 123.615 ;
        RECT 65.670 123.445 65.920 124.815 ;
        RECT 64.940 122.985 65.190 123.445 ;
        RECT 65.360 123.155 65.920 123.445 ;
        RECT 66.090 124.395 66.360 125.365 ;
        RECT 66.570 124.735 66.850 125.535 ;
        RECT 67.020 125.025 68.675 125.315 ;
        RECT 67.085 124.685 68.675 124.855 ;
        RECT 67.085 124.565 67.255 124.685 ;
        RECT 66.530 124.395 67.255 124.565 ;
        RECT 66.090 123.660 66.260 124.395 ;
        RECT 66.530 124.225 66.700 124.395 ;
        RECT 67.445 124.345 68.160 124.515 ;
        RECT 68.355 124.395 68.675 124.685 ;
        RECT 68.850 124.565 69.160 125.365 ;
        RECT 69.330 124.735 69.640 125.535 ;
        RECT 69.810 124.905 70.070 125.365 ;
        RECT 70.240 125.075 70.495 125.535 ;
        RECT 70.670 124.905 70.930 125.365 ;
        RECT 69.810 124.735 70.930 124.905 ;
        RECT 68.850 124.395 69.880 124.565 ;
        RECT 66.430 123.895 66.700 124.225 ;
        RECT 66.870 123.895 67.275 124.225 ;
        RECT 67.445 123.895 68.155 124.345 ;
        RECT 66.530 123.725 66.700 123.895 ;
        RECT 66.090 123.315 66.360 123.660 ;
        RECT 66.530 123.555 68.140 123.725 ;
        RECT 68.325 123.655 68.675 124.225 ;
        RECT 66.550 122.985 66.930 123.385 ;
        RECT 67.100 123.205 67.270 123.555 ;
        RECT 67.440 122.985 67.770 123.385 ;
        RECT 67.970 123.205 68.140 123.555 ;
        RECT 68.850 123.485 69.020 124.395 ;
        RECT 69.190 123.655 69.540 124.225 ;
        RECT 69.710 124.145 69.880 124.395 ;
        RECT 70.670 124.485 70.930 124.735 ;
        RECT 71.100 124.665 71.385 125.535 ;
        RECT 71.700 124.790 71.970 125.535 ;
        RECT 72.600 125.530 78.875 125.535 ;
        RECT 72.140 124.620 72.430 125.360 ;
        RECT 72.600 124.805 72.855 125.530 ;
        RECT 73.040 124.635 73.300 125.360 ;
        RECT 73.470 124.805 73.715 125.530 ;
        RECT 73.900 124.635 74.160 125.360 ;
        RECT 74.330 124.805 74.575 125.530 ;
        RECT 74.760 124.635 75.020 125.360 ;
        RECT 75.190 124.805 75.435 125.530 ;
        RECT 75.605 124.635 75.865 125.360 ;
        RECT 76.035 124.805 76.295 125.530 ;
        RECT 76.465 124.635 76.725 125.360 ;
        RECT 76.895 124.805 77.155 125.530 ;
        RECT 77.325 124.635 77.585 125.360 ;
        RECT 77.755 124.805 78.015 125.530 ;
        RECT 78.185 124.635 78.445 125.360 ;
        RECT 78.615 124.735 78.875 125.530 ;
        RECT 73.040 124.620 78.445 124.635 ;
        RECT 70.670 124.315 71.425 124.485 ;
        RECT 69.710 123.975 70.850 124.145 ;
        RECT 71.020 123.805 71.425 124.315 ;
        RECT 69.775 123.635 71.425 123.805 ;
        RECT 71.700 124.395 78.445 124.620 ;
        RECT 71.700 123.805 72.865 124.395 ;
        RECT 79.045 124.225 79.295 125.360 ;
        RECT 79.475 124.725 79.735 125.535 ;
        RECT 79.910 124.225 80.155 125.365 ;
        RECT 80.335 124.725 80.630 125.535 ;
        RECT 80.810 124.460 81.080 125.365 ;
        RECT 81.250 124.775 81.580 125.535 ;
        RECT 81.760 124.605 81.930 125.365 ;
        RECT 73.035 123.975 80.155 124.225 ;
        RECT 71.700 123.635 78.445 123.805 ;
        RECT 68.340 122.985 68.670 123.485 ;
        RECT 68.850 123.155 69.150 123.485 ;
        RECT 69.320 122.985 69.595 123.465 ;
        RECT 69.775 123.245 70.070 123.635 ;
        RECT 70.240 122.985 70.495 123.465 ;
        RECT 70.670 123.245 70.930 123.635 ;
        RECT 71.100 122.985 71.380 123.465 ;
        RECT 71.700 122.985 72.000 123.465 ;
        RECT 72.170 123.180 72.430 123.635 ;
        RECT 72.600 122.985 72.860 123.465 ;
        RECT 73.040 123.180 73.300 123.635 ;
        RECT 73.470 122.985 73.720 123.465 ;
        RECT 73.900 123.180 74.160 123.635 ;
        RECT 74.330 122.985 74.580 123.465 ;
        RECT 74.760 123.180 75.020 123.635 ;
        RECT 75.190 122.985 75.435 123.465 ;
        RECT 75.605 123.180 75.880 123.635 ;
        RECT 76.050 122.985 76.295 123.465 ;
        RECT 76.465 123.180 76.725 123.635 ;
        RECT 76.895 122.985 77.155 123.465 ;
        RECT 77.325 123.180 77.585 123.635 ;
        RECT 77.755 122.985 78.015 123.465 ;
        RECT 78.185 123.180 78.445 123.635 ;
        RECT 78.615 122.985 78.875 123.545 ;
        RECT 79.045 123.165 79.295 123.975 ;
        RECT 79.475 122.985 79.735 123.510 ;
        RECT 79.905 123.165 80.155 123.975 ;
        RECT 80.325 123.665 80.640 124.225 ;
        RECT 80.810 123.660 80.980 124.460 ;
        RECT 81.265 124.435 81.930 124.605 ;
        RECT 82.190 124.775 82.705 125.185 ;
        RECT 82.940 124.775 83.110 125.535 ;
        RECT 83.280 125.195 85.310 125.365 ;
        RECT 81.265 124.290 81.435 124.435 ;
        RECT 81.150 123.960 81.435 124.290 ;
        RECT 81.265 123.705 81.435 123.960 ;
        RECT 81.670 123.885 82.000 124.255 ;
        RECT 82.190 123.965 82.530 124.775 ;
        RECT 83.280 124.530 83.450 125.195 ;
        RECT 83.845 124.855 84.970 125.025 ;
        RECT 82.700 124.340 83.450 124.530 ;
        RECT 83.620 124.515 84.630 124.685 ;
        RECT 82.190 123.795 83.420 123.965 ;
        RECT 80.335 122.985 80.640 123.495 ;
        RECT 80.810 123.155 81.070 123.660 ;
        RECT 81.265 123.535 81.930 123.705 ;
        RECT 81.250 122.985 81.580 123.365 ;
        RECT 81.760 123.155 81.930 123.535 ;
        RECT 82.465 123.190 82.710 123.795 ;
        RECT 82.930 122.985 83.440 123.520 ;
        RECT 83.620 123.155 83.810 124.515 ;
        RECT 83.980 123.495 84.255 124.315 ;
        RECT 84.460 123.715 84.630 124.515 ;
        RECT 84.800 123.725 84.970 124.855 ;
        RECT 85.140 124.225 85.310 125.195 ;
        RECT 85.480 124.395 85.650 125.535 ;
        RECT 85.820 124.395 86.155 125.365 ;
        RECT 85.140 123.895 85.335 124.225 ;
        RECT 85.560 123.895 85.815 124.225 ;
        RECT 85.560 123.725 85.730 123.895 ;
        RECT 85.985 123.725 86.155 124.395 ;
        RECT 86.330 124.370 86.620 125.535 ;
        RECT 87.450 124.865 87.730 125.535 ;
        RECT 87.900 124.645 88.200 125.195 ;
        RECT 88.400 124.815 88.730 125.535 ;
        RECT 88.920 124.815 89.380 125.365 ;
        RECT 87.265 124.225 87.530 124.585 ;
        RECT 87.900 124.475 88.840 124.645 ;
        RECT 88.670 124.225 88.840 124.475 ;
        RECT 87.265 123.975 87.940 124.225 ;
        RECT 88.160 123.975 88.500 124.225 ;
        RECT 88.670 123.895 88.960 124.225 ;
        RECT 88.670 123.805 88.840 123.895 ;
        RECT 84.800 123.555 85.730 123.725 ;
        RECT 84.800 123.520 84.975 123.555 ;
        RECT 83.980 123.325 84.260 123.495 ;
        RECT 83.980 123.155 84.255 123.325 ;
        RECT 84.445 123.155 84.975 123.520 ;
        RECT 85.400 122.985 85.730 123.385 ;
        RECT 85.900 123.155 86.155 123.725 ;
        RECT 86.330 122.985 86.620 123.710 ;
        RECT 87.450 123.615 88.840 123.805 ;
        RECT 87.450 123.255 87.780 123.615 ;
        RECT 89.130 123.445 89.380 124.815 ;
        RECT 88.400 122.985 88.650 123.445 ;
        RECT 88.820 123.155 89.380 123.445 ;
        RECT 89.550 124.815 90.010 125.365 ;
        RECT 90.200 124.815 90.530 125.535 ;
        RECT 89.550 123.445 89.800 124.815 ;
        RECT 90.730 124.645 91.030 125.195 ;
        RECT 91.200 124.865 91.480 125.535 ;
        RECT 92.510 124.865 92.790 125.535 ;
        RECT 90.090 124.475 91.030 124.645 ;
        RECT 92.960 124.645 93.260 125.195 ;
        RECT 93.460 124.815 93.790 125.535 ;
        RECT 93.980 124.815 94.440 125.365 ;
        RECT 90.090 124.225 90.260 124.475 ;
        RECT 91.400 124.225 91.665 124.585 ;
        RECT 89.970 123.895 90.260 124.225 ;
        RECT 90.430 123.975 90.770 124.225 ;
        RECT 90.990 123.975 91.665 124.225 ;
        RECT 92.325 124.225 92.590 124.585 ;
        RECT 92.960 124.475 93.900 124.645 ;
        RECT 93.730 124.225 93.900 124.475 ;
        RECT 92.325 123.975 93.000 124.225 ;
        RECT 93.220 123.975 93.560 124.225 ;
        RECT 90.090 123.805 90.260 123.895 ;
        RECT 93.730 123.895 94.020 124.225 ;
        RECT 93.730 123.805 93.900 123.895 ;
        RECT 90.090 123.615 91.480 123.805 ;
        RECT 89.550 123.155 90.110 123.445 ;
        RECT 90.280 122.985 90.530 123.445 ;
        RECT 91.150 123.255 91.480 123.615 ;
        RECT 92.510 123.615 93.900 123.805 ;
        RECT 92.510 123.255 92.840 123.615 ;
        RECT 94.190 123.445 94.440 124.815 ;
        RECT 93.460 122.985 93.710 123.445 ;
        RECT 93.880 123.155 94.440 123.445 ;
        RECT 94.610 124.815 95.070 125.365 ;
        RECT 95.260 124.815 95.590 125.535 ;
        RECT 94.610 123.445 94.860 124.815 ;
        RECT 95.790 124.645 96.090 125.195 ;
        RECT 96.260 124.865 96.540 125.535 ;
        RECT 95.150 124.475 96.090 124.645 ;
        RECT 97.370 124.775 97.885 125.185 ;
        RECT 98.120 124.775 98.290 125.535 ;
        RECT 98.460 125.195 100.490 125.365 ;
        RECT 95.150 124.225 95.320 124.475 ;
        RECT 96.460 124.225 96.725 124.585 ;
        RECT 95.030 123.895 95.320 124.225 ;
        RECT 95.490 123.975 95.830 124.225 ;
        RECT 96.050 123.975 96.725 124.225 ;
        RECT 95.150 123.805 95.320 123.895 ;
        RECT 97.370 123.965 97.710 124.775 ;
        RECT 98.460 124.530 98.630 125.195 ;
        RECT 99.025 124.855 100.150 125.025 ;
        RECT 97.880 124.340 98.630 124.530 ;
        RECT 98.800 124.515 99.810 124.685 ;
        RECT 95.150 123.615 96.540 123.805 ;
        RECT 97.370 123.795 98.600 123.965 ;
        RECT 94.610 123.155 95.170 123.445 ;
        RECT 95.340 122.985 95.590 123.445 ;
        RECT 96.210 123.255 96.540 123.615 ;
        RECT 97.645 123.190 97.890 123.795 ;
        RECT 98.110 122.985 98.620 123.520 ;
        RECT 98.800 123.155 98.990 124.515 ;
        RECT 99.160 123.495 99.435 124.315 ;
        RECT 99.640 123.715 99.810 124.515 ;
        RECT 99.980 123.725 100.150 124.855 ;
        RECT 100.320 124.225 100.490 125.195 ;
        RECT 100.660 124.395 100.830 125.535 ;
        RECT 101.000 124.395 101.335 125.365 ;
        RECT 100.320 123.895 100.515 124.225 ;
        RECT 100.740 123.895 100.995 124.225 ;
        RECT 100.740 123.725 100.910 123.895 ;
        RECT 101.165 123.725 101.335 124.395 ;
        RECT 99.980 123.555 100.910 123.725 ;
        RECT 99.980 123.520 100.155 123.555 ;
        RECT 99.160 123.325 99.440 123.495 ;
        RECT 99.160 123.155 99.435 123.325 ;
        RECT 99.625 123.155 100.155 123.520 ;
        RECT 100.580 122.985 100.910 123.385 ;
        RECT 101.080 123.155 101.335 123.725 ;
        RECT 101.885 124.555 102.140 125.225 ;
        RECT 102.320 124.735 102.605 125.535 ;
        RECT 102.785 124.815 103.115 125.325 ;
        RECT 101.885 123.695 102.065 124.555 ;
        RECT 102.785 124.225 103.035 124.815 ;
        RECT 103.385 124.665 103.555 125.275 ;
        RECT 103.725 124.845 104.055 125.535 ;
        RECT 104.285 124.985 104.525 125.275 ;
        RECT 104.725 125.155 105.145 125.535 ;
        RECT 105.325 125.065 105.955 125.315 ;
        RECT 106.425 125.155 106.755 125.535 ;
        RECT 105.325 124.985 105.495 125.065 ;
        RECT 106.925 124.985 107.095 125.275 ;
        RECT 107.275 125.155 107.655 125.535 ;
        RECT 107.895 125.150 108.725 125.320 ;
        RECT 104.285 124.815 105.495 124.985 ;
        RECT 102.235 123.895 103.035 124.225 ;
        RECT 101.885 123.495 102.140 123.695 ;
        RECT 101.800 123.325 102.140 123.495 ;
        RECT 101.885 123.165 102.140 123.325 ;
        RECT 102.320 122.985 102.605 123.445 ;
        RECT 102.785 123.245 103.035 123.895 ;
        RECT 103.235 124.645 103.555 124.665 ;
        RECT 103.235 124.475 105.155 124.645 ;
        RECT 103.235 123.580 103.425 124.475 ;
        RECT 105.325 124.305 105.495 124.815 ;
        RECT 105.665 124.555 106.185 124.865 ;
        RECT 103.595 124.135 105.495 124.305 ;
        RECT 103.595 124.075 103.925 124.135 ;
        RECT 104.075 123.905 104.405 123.965 ;
        RECT 103.745 123.635 104.405 123.905 ;
        RECT 103.235 123.250 103.555 123.580 ;
        RECT 103.735 122.985 104.395 123.465 ;
        RECT 104.595 123.375 104.765 124.135 ;
        RECT 105.665 123.965 105.845 124.375 ;
        RECT 104.935 123.795 105.265 123.915 ;
        RECT 106.015 123.795 106.185 124.555 ;
        RECT 104.935 123.625 106.185 123.795 ;
        RECT 106.355 124.735 107.725 124.985 ;
        RECT 106.355 123.965 106.545 124.735 ;
        RECT 107.475 124.475 107.725 124.735 ;
        RECT 106.715 124.305 106.965 124.465 ;
        RECT 107.895 124.305 108.065 125.150 ;
        RECT 108.960 124.865 109.130 125.365 ;
        RECT 109.300 125.035 109.630 125.535 ;
        RECT 108.235 124.475 108.735 124.855 ;
        RECT 108.960 124.695 109.655 124.865 ;
        RECT 106.715 124.135 108.065 124.305 ;
        RECT 107.645 124.095 108.065 124.135 ;
        RECT 106.355 123.625 106.775 123.965 ;
        RECT 107.065 123.635 107.475 123.965 ;
        RECT 104.595 123.205 105.445 123.375 ;
        RECT 106.005 122.985 106.325 123.445 ;
        RECT 106.525 123.195 106.775 123.625 ;
        RECT 107.065 122.985 107.475 123.425 ;
        RECT 107.645 123.365 107.815 124.095 ;
        RECT 107.985 123.545 108.335 123.915 ;
        RECT 108.515 123.605 108.735 124.475 ;
        RECT 108.905 123.905 109.315 124.525 ;
        RECT 109.485 123.725 109.655 124.695 ;
        RECT 108.960 123.535 109.655 123.725 ;
        RECT 107.645 123.165 108.660 123.365 ;
        RECT 108.960 123.205 109.130 123.535 ;
        RECT 109.300 122.985 109.630 123.365 ;
        RECT 109.845 123.245 110.070 125.365 ;
        RECT 110.240 125.035 110.570 125.535 ;
        RECT 110.740 124.865 110.910 125.365 ;
        RECT 110.245 124.695 110.910 124.865 ;
        RECT 110.245 123.705 110.475 124.695 ;
        RECT 110.645 123.875 110.995 124.525 ;
        RECT 111.170 124.445 112.380 125.535 ;
        RECT 111.170 123.905 111.690 124.445 ;
        RECT 111.860 123.735 112.380 124.275 ;
        RECT 110.245 123.535 110.910 123.705 ;
        RECT 110.240 122.985 110.570 123.365 ;
        RECT 110.740 123.245 110.910 123.535 ;
        RECT 111.170 122.985 112.380 123.735 ;
        RECT 18.165 122.815 112.465 122.985 ;
        RECT 18.250 122.065 19.460 122.815 ;
        RECT 20.640 122.265 20.810 122.645 ;
        RECT 20.990 122.435 21.320 122.815 ;
        RECT 20.640 122.095 21.305 122.265 ;
        RECT 21.500 122.140 21.760 122.645 ;
        RECT 18.250 121.525 18.770 122.065 ;
        RECT 18.940 121.355 19.460 121.895 ;
        RECT 20.570 121.545 20.900 121.915 ;
        RECT 21.135 121.840 21.305 122.095 ;
        RECT 21.135 121.510 21.420 121.840 ;
        RECT 21.135 121.365 21.305 121.510 ;
        RECT 18.250 120.265 19.460 121.355 ;
        RECT 20.640 121.195 21.305 121.365 ;
        RECT 21.590 121.340 21.760 122.140 ;
        RECT 21.930 122.090 22.220 122.815 ;
        RECT 22.765 122.105 23.020 122.635 ;
        RECT 23.200 122.355 23.485 122.815 ;
        RECT 20.640 120.435 20.810 121.195 ;
        RECT 20.990 120.265 21.320 121.025 ;
        RECT 21.490 120.435 21.760 121.340 ;
        RECT 21.930 120.265 22.220 121.430 ;
        RECT 22.765 121.245 22.945 122.105 ;
        RECT 23.665 121.905 23.915 122.555 ;
        RECT 23.115 121.575 23.915 121.905 ;
        RECT 22.765 120.775 23.020 121.245 ;
        RECT 22.680 120.605 23.020 120.775 ;
        RECT 22.765 120.575 23.020 120.605 ;
        RECT 23.200 120.265 23.485 121.065 ;
        RECT 23.665 120.985 23.915 121.575 ;
        RECT 24.115 122.220 24.435 122.550 ;
        RECT 24.615 122.335 25.275 122.815 ;
        RECT 25.475 122.425 26.325 122.595 ;
        RECT 24.115 121.325 24.305 122.220 ;
        RECT 24.625 121.895 25.285 122.165 ;
        RECT 24.955 121.835 25.285 121.895 ;
        RECT 24.475 121.665 24.805 121.725 ;
        RECT 25.475 121.665 25.645 122.425 ;
        RECT 26.885 122.355 27.205 122.815 ;
        RECT 27.405 122.175 27.655 122.605 ;
        RECT 27.945 122.375 28.355 122.815 ;
        RECT 28.525 122.435 29.540 122.635 ;
        RECT 25.815 122.005 27.065 122.175 ;
        RECT 25.815 121.885 26.145 122.005 ;
        RECT 24.475 121.495 26.375 121.665 ;
        RECT 24.115 121.155 26.035 121.325 ;
        RECT 24.115 121.135 24.435 121.155 ;
        RECT 23.665 120.475 23.995 120.985 ;
        RECT 24.265 120.525 24.435 121.135 ;
        RECT 26.205 120.985 26.375 121.495 ;
        RECT 26.545 121.425 26.725 121.835 ;
        RECT 26.895 121.245 27.065 122.005 ;
        RECT 24.605 120.265 24.935 120.955 ;
        RECT 25.165 120.815 26.375 120.985 ;
        RECT 26.545 120.935 27.065 121.245 ;
        RECT 27.235 121.835 27.655 122.175 ;
        RECT 27.945 121.835 28.355 122.165 ;
        RECT 27.235 121.065 27.425 121.835 ;
        RECT 28.525 121.705 28.695 122.435 ;
        RECT 29.840 122.265 30.010 122.595 ;
        RECT 30.180 122.435 30.510 122.815 ;
        RECT 28.865 121.885 29.215 122.255 ;
        RECT 28.525 121.665 28.945 121.705 ;
        RECT 27.595 121.495 28.945 121.665 ;
        RECT 27.595 121.335 27.845 121.495 ;
        RECT 28.355 121.065 28.605 121.325 ;
        RECT 27.235 120.815 28.605 121.065 ;
        RECT 25.165 120.525 25.405 120.815 ;
        RECT 26.205 120.735 26.375 120.815 ;
        RECT 25.605 120.265 26.025 120.645 ;
        RECT 26.205 120.485 26.835 120.735 ;
        RECT 27.305 120.265 27.635 120.645 ;
        RECT 27.805 120.525 27.975 120.815 ;
        RECT 28.775 120.650 28.945 121.495 ;
        RECT 29.395 121.325 29.615 122.195 ;
        RECT 29.840 122.075 30.535 122.265 ;
        RECT 29.115 120.945 29.615 121.325 ;
        RECT 29.785 121.275 30.195 121.895 ;
        RECT 30.365 121.105 30.535 122.075 ;
        RECT 29.840 120.935 30.535 121.105 ;
        RECT 28.155 120.265 28.535 120.645 ;
        RECT 28.775 120.480 29.605 120.650 ;
        RECT 29.840 120.435 30.010 120.935 ;
        RECT 30.180 120.265 30.510 120.765 ;
        RECT 30.725 120.435 30.950 122.555 ;
        RECT 31.120 122.435 31.450 122.815 ;
        RECT 31.620 122.265 31.790 122.555 ;
        RECT 32.425 122.475 32.680 122.635 ;
        RECT 32.340 122.305 32.680 122.475 ;
        RECT 32.860 122.355 33.145 122.815 ;
        RECT 31.125 122.095 31.790 122.265 ;
        RECT 32.425 122.105 32.680 122.305 ;
        RECT 31.125 121.105 31.355 122.095 ;
        RECT 31.525 121.275 31.875 121.925 ;
        RECT 32.425 121.245 32.605 122.105 ;
        RECT 33.325 121.905 33.575 122.555 ;
        RECT 32.775 121.575 33.575 121.905 ;
        RECT 31.125 120.935 31.790 121.105 ;
        RECT 31.120 120.265 31.450 120.765 ;
        RECT 31.620 120.435 31.790 120.935 ;
        RECT 32.425 120.575 32.680 121.245 ;
        RECT 32.860 120.265 33.145 121.065 ;
        RECT 33.325 120.985 33.575 121.575 ;
        RECT 33.775 122.220 34.095 122.550 ;
        RECT 34.275 122.335 34.935 122.815 ;
        RECT 35.135 122.425 35.985 122.595 ;
        RECT 33.775 121.325 33.965 122.220 ;
        RECT 34.285 121.895 34.945 122.165 ;
        RECT 34.615 121.835 34.945 121.895 ;
        RECT 34.135 121.665 34.465 121.725 ;
        RECT 35.135 121.665 35.305 122.425 ;
        RECT 36.545 122.355 36.865 122.815 ;
        RECT 37.065 122.175 37.315 122.605 ;
        RECT 37.605 122.375 38.015 122.815 ;
        RECT 38.185 122.435 39.200 122.635 ;
        RECT 35.475 122.005 36.725 122.175 ;
        RECT 35.475 121.885 35.805 122.005 ;
        RECT 34.135 121.495 36.035 121.665 ;
        RECT 33.775 121.155 35.695 121.325 ;
        RECT 33.775 121.135 34.095 121.155 ;
        RECT 33.325 120.475 33.655 120.985 ;
        RECT 33.925 120.525 34.095 121.135 ;
        RECT 35.865 120.985 36.035 121.495 ;
        RECT 36.205 121.425 36.385 121.835 ;
        RECT 36.555 121.245 36.725 122.005 ;
        RECT 34.265 120.265 34.595 120.955 ;
        RECT 34.825 120.815 36.035 120.985 ;
        RECT 36.205 120.935 36.725 121.245 ;
        RECT 36.895 121.835 37.315 122.175 ;
        RECT 37.605 121.835 38.015 122.165 ;
        RECT 36.895 121.065 37.085 121.835 ;
        RECT 38.185 121.705 38.355 122.435 ;
        RECT 39.500 122.265 39.670 122.595 ;
        RECT 39.840 122.435 40.170 122.815 ;
        RECT 38.525 121.885 38.875 122.255 ;
        RECT 38.185 121.665 38.605 121.705 ;
        RECT 37.255 121.495 38.605 121.665 ;
        RECT 37.255 121.335 37.505 121.495 ;
        RECT 38.015 121.065 38.265 121.325 ;
        RECT 36.895 120.815 38.265 121.065 ;
        RECT 34.825 120.525 35.065 120.815 ;
        RECT 35.865 120.735 36.035 120.815 ;
        RECT 35.265 120.265 35.685 120.645 ;
        RECT 35.865 120.485 36.495 120.735 ;
        RECT 36.965 120.265 37.295 120.645 ;
        RECT 37.465 120.525 37.635 120.815 ;
        RECT 38.435 120.650 38.605 121.495 ;
        RECT 39.055 121.325 39.275 122.195 ;
        RECT 39.500 122.075 40.195 122.265 ;
        RECT 38.775 120.945 39.275 121.325 ;
        RECT 39.445 121.275 39.855 121.895 ;
        RECT 40.025 121.105 40.195 122.075 ;
        RECT 39.500 120.935 40.195 121.105 ;
        RECT 37.815 120.265 38.195 120.645 ;
        RECT 38.435 120.480 39.265 120.650 ;
        RECT 39.500 120.435 39.670 120.935 ;
        RECT 39.840 120.265 40.170 120.765 ;
        RECT 40.385 120.435 40.610 122.555 ;
        RECT 40.780 122.435 41.110 122.815 ;
        RECT 41.280 122.265 41.450 122.555 ;
        RECT 41.710 122.310 41.995 122.815 ;
        RECT 40.785 122.095 41.450 122.265 ;
        RECT 42.165 122.140 42.490 122.645 ;
        RECT 40.785 121.105 41.015 122.095 ;
        RECT 41.185 121.275 41.535 121.925 ;
        RECT 41.710 121.610 42.490 122.140 ;
        RECT 40.785 120.935 41.450 121.105 ;
        RECT 40.780 120.265 41.110 120.765 ;
        RECT 41.280 120.435 41.450 120.935 ;
        RECT 41.710 120.265 41.990 121.235 ;
        RECT 42.160 120.435 42.490 121.610 ;
        RECT 42.680 121.575 42.920 122.525 ;
        RECT 43.550 122.355 44.110 122.645 ;
        RECT 44.280 122.355 44.530 122.815 ;
        RECT 42.660 120.265 42.920 121.235 ;
        RECT 43.550 120.985 43.800 122.355 ;
        RECT 45.150 122.185 45.480 122.545 ;
        RECT 44.090 121.995 45.480 122.185 ;
        RECT 46.400 122.265 46.570 122.645 ;
        RECT 46.750 122.435 47.080 122.815 ;
        RECT 46.400 122.095 47.065 122.265 ;
        RECT 47.260 122.140 47.520 122.645 ;
        RECT 44.090 121.905 44.260 121.995 ;
        RECT 43.970 121.575 44.260 121.905 ;
        RECT 44.430 121.575 44.770 121.825 ;
        RECT 44.990 121.575 45.665 121.825 ;
        RECT 44.090 121.325 44.260 121.575 ;
        RECT 44.090 121.155 45.030 121.325 ;
        RECT 45.400 121.215 45.665 121.575 ;
        RECT 46.330 121.545 46.660 121.915 ;
        RECT 46.895 121.840 47.065 122.095 ;
        RECT 46.895 121.510 47.180 121.840 ;
        RECT 46.895 121.365 47.065 121.510 ;
        RECT 43.550 120.435 44.010 120.985 ;
        RECT 44.200 120.265 44.530 120.985 ;
        RECT 44.730 120.605 45.030 121.155 ;
        RECT 46.400 121.195 47.065 121.365 ;
        RECT 47.350 121.340 47.520 122.140 ;
        RECT 47.690 122.090 47.980 122.815 ;
        RECT 48.150 122.305 48.455 122.815 ;
        RECT 48.150 121.575 48.465 122.135 ;
        RECT 48.635 121.825 48.885 122.635 ;
        RECT 49.055 122.290 49.315 122.815 ;
        RECT 49.495 121.825 49.745 122.635 ;
        RECT 49.915 122.255 50.175 122.815 ;
        RECT 50.345 122.165 50.605 122.620 ;
        RECT 50.775 122.335 51.035 122.815 ;
        RECT 51.205 122.165 51.465 122.620 ;
        RECT 51.635 122.335 51.895 122.815 ;
        RECT 52.065 122.165 52.325 122.620 ;
        RECT 52.495 122.335 52.740 122.815 ;
        RECT 52.910 122.165 53.185 122.620 ;
        RECT 53.355 122.335 53.600 122.815 ;
        RECT 53.770 122.165 54.030 122.620 ;
        RECT 54.210 122.335 54.460 122.815 ;
        RECT 54.630 122.165 54.890 122.620 ;
        RECT 55.070 122.335 55.320 122.815 ;
        RECT 55.490 122.165 55.750 122.620 ;
        RECT 55.930 122.335 56.190 122.815 ;
        RECT 56.360 122.165 56.620 122.620 ;
        RECT 56.790 122.335 57.090 122.815 ;
        RECT 58.185 122.475 58.440 122.635 ;
        RECT 58.100 122.305 58.440 122.475 ;
        RECT 58.620 122.355 58.905 122.815 ;
        RECT 50.345 121.995 57.090 122.165 ;
        RECT 48.635 121.575 55.755 121.825 ;
        RECT 45.200 120.265 45.480 120.935 ;
        RECT 46.400 120.435 46.570 121.195 ;
        RECT 46.750 120.265 47.080 121.025 ;
        RECT 47.250 120.435 47.520 121.340 ;
        RECT 47.690 120.265 47.980 121.430 ;
        RECT 48.160 120.265 48.455 121.075 ;
        RECT 48.635 120.435 48.880 121.575 ;
        RECT 49.055 120.265 49.315 121.075 ;
        RECT 49.495 120.440 49.745 121.575 ;
        RECT 55.925 121.455 57.090 121.995 ;
        RECT 58.185 122.105 58.440 122.305 ;
        RECT 55.925 121.405 57.120 121.455 ;
        RECT 50.345 121.285 57.120 121.405 ;
        RECT 50.345 121.180 57.090 121.285 ;
        RECT 58.185 121.245 58.365 122.105 ;
        RECT 59.085 121.905 59.335 122.555 ;
        RECT 58.535 121.575 59.335 121.905 ;
        RECT 50.345 121.165 55.750 121.180 ;
        RECT 49.915 120.270 50.175 121.065 ;
        RECT 50.345 120.440 50.605 121.165 ;
        RECT 50.775 120.270 51.035 120.995 ;
        RECT 51.205 120.440 51.465 121.165 ;
        RECT 51.635 120.270 51.895 120.995 ;
        RECT 52.065 120.440 52.325 121.165 ;
        RECT 52.495 120.270 52.755 120.995 ;
        RECT 52.925 120.440 53.185 121.165 ;
        RECT 53.355 120.270 53.600 120.995 ;
        RECT 53.770 120.440 54.030 121.165 ;
        RECT 54.215 120.270 54.460 120.995 ;
        RECT 54.630 120.440 54.890 121.165 ;
        RECT 55.075 120.270 55.320 120.995 ;
        RECT 55.490 120.440 55.750 121.165 ;
        RECT 55.935 120.270 56.190 120.995 ;
        RECT 56.360 120.440 56.650 121.180 ;
        RECT 49.915 120.265 56.190 120.270 ;
        RECT 56.820 120.265 57.090 121.010 ;
        RECT 58.185 120.575 58.440 121.245 ;
        RECT 58.620 120.265 58.905 121.065 ;
        RECT 59.085 120.985 59.335 121.575 ;
        RECT 59.535 122.220 59.855 122.550 ;
        RECT 60.035 122.335 60.695 122.815 ;
        RECT 60.895 122.425 61.745 122.595 ;
        RECT 59.535 121.325 59.725 122.220 ;
        RECT 60.045 121.895 60.705 122.165 ;
        RECT 60.375 121.835 60.705 121.895 ;
        RECT 59.895 121.665 60.225 121.725 ;
        RECT 60.895 121.665 61.065 122.425 ;
        RECT 62.305 122.355 62.625 122.815 ;
        RECT 62.825 122.175 63.075 122.605 ;
        RECT 63.365 122.375 63.775 122.815 ;
        RECT 63.945 122.435 64.960 122.635 ;
        RECT 61.235 122.005 62.485 122.175 ;
        RECT 61.235 121.885 61.565 122.005 ;
        RECT 59.895 121.495 61.795 121.665 ;
        RECT 59.535 121.155 61.455 121.325 ;
        RECT 59.535 121.135 59.855 121.155 ;
        RECT 59.085 120.475 59.415 120.985 ;
        RECT 59.685 120.525 59.855 121.135 ;
        RECT 61.625 120.985 61.795 121.495 ;
        RECT 61.965 121.425 62.145 121.835 ;
        RECT 62.315 121.245 62.485 122.005 ;
        RECT 60.025 120.265 60.355 120.955 ;
        RECT 60.585 120.815 61.795 120.985 ;
        RECT 61.965 120.935 62.485 121.245 ;
        RECT 62.655 121.835 63.075 122.175 ;
        RECT 63.365 121.835 63.775 122.165 ;
        RECT 62.655 121.065 62.845 121.835 ;
        RECT 63.945 121.705 64.115 122.435 ;
        RECT 65.260 122.265 65.430 122.595 ;
        RECT 65.600 122.435 65.930 122.815 ;
        RECT 64.285 121.885 64.635 122.255 ;
        RECT 63.945 121.665 64.365 121.705 ;
        RECT 63.015 121.495 64.365 121.665 ;
        RECT 63.015 121.335 63.265 121.495 ;
        RECT 63.775 121.065 64.025 121.325 ;
        RECT 62.655 120.815 64.025 121.065 ;
        RECT 60.585 120.525 60.825 120.815 ;
        RECT 61.625 120.735 61.795 120.815 ;
        RECT 61.025 120.265 61.445 120.645 ;
        RECT 61.625 120.485 62.255 120.735 ;
        RECT 62.725 120.265 63.055 120.645 ;
        RECT 63.225 120.525 63.395 120.815 ;
        RECT 64.195 120.650 64.365 121.495 ;
        RECT 64.815 121.325 65.035 122.195 ;
        RECT 65.260 122.075 65.955 122.265 ;
        RECT 64.535 120.945 65.035 121.325 ;
        RECT 65.205 121.275 65.615 121.895 ;
        RECT 65.785 121.105 65.955 122.075 ;
        RECT 65.260 120.935 65.955 121.105 ;
        RECT 63.575 120.265 63.955 120.645 ;
        RECT 64.195 120.480 65.025 120.650 ;
        RECT 65.260 120.435 65.430 120.935 ;
        RECT 65.600 120.265 65.930 120.765 ;
        RECT 66.145 120.435 66.370 122.555 ;
        RECT 66.540 122.435 66.870 122.815 ;
        RECT 67.040 122.265 67.210 122.555 ;
        RECT 66.545 122.095 67.210 122.265 ;
        RECT 67.470 122.315 67.730 122.645 ;
        RECT 67.940 122.335 68.215 122.815 ;
        RECT 66.545 121.105 66.775 122.095 ;
        RECT 66.945 121.275 67.295 121.925 ;
        RECT 67.470 121.405 67.640 122.315 ;
        RECT 68.425 122.245 68.630 122.645 ;
        RECT 68.800 122.415 69.135 122.815 ;
        RECT 67.810 121.575 68.170 122.155 ;
        RECT 68.425 122.075 69.110 122.245 ;
        RECT 68.350 121.405 68.600 121.905 ;
        RECT 67.470 121.235 68.600 121.405 ;
        RECT 66.545 120.935 67.210 121.105 ;
        RECT 66.540 120.265 66.870 120.765 ;
        RECT 67.040 120.435 67.210 120.935 ;
        RECT 67.470 120.465 67.740 121.235 ;
        RECT 68.770 121.045 69.110 122.075 ;
        RECT 69.585 122.005 69.830 122.610 ;
        RECT 70.050 122.280 70.560 122.815 ;
        RECT 67.910 120.265 68.240 121.045 ;
        RECT 68.445 120.870 69.110 121.045 ;
        RECT 69.310 121.835 70.540 122.005 ;
        RECT 69.310 121.025 69.650 121.835 ;
        RECT 69.820 121.270 70.570 121.460 ;
        RECT 68.445 120.465 68.630 120.870 ;
        RECT 68.800 120.265 69.135 120.690 ;
        RECT 69.310 120.615 69.825 121.025 ;
        RECT 70.060 120.265 70.230 121.025 ;
        RECT 70.400 120.605 70.570 121.270 ;
        RECT 70.740 121.285 70.930 122.645 ;
        RECT 71.100 122.475 71.375 122.645 ;
        RECT 71.100 122.305 71.380 122.475 ;
        RECT 71.100 121.485 71.375 122.305 ;
        RECT 71.565 122.280 72.095 122.645 ;
        RECT 72.520 122.415 72.850 122.815 ;
        RECT 71.920 122.245 72.095 122.280 ;
        RECT 71.580 121.285 71.750 122.085 ;
        RECT 70.740 121.115 71.750 121.285 ;
        RECT 71.920 122.075 72.850 122.245 ;
        RECT 73.020 122.075 73.275 122.645 ;
        RECT 73.450 122.090 73.740 122.815 ;
        RECT 74.430 122.345 74.730 122.815 ;
        RECT 74.900 122.175 75.155 122.620 ;
        RECT 75.325 122.345 75.585 122.815 ;
        RECT 75.755 122.175 76.015 122.620 ;
        RECT 76.185 122.345 76.480 122.815 ;
        RECT 77.220 122.265 77.390 122.555 ;
        RECT 77.560 122.435 77.890 122.815 ;
        RECT 71.920 120.945 72.090 122.075 ;
        RECT 72.680 121.905 72.850 122.075 ;
        RECT 70.965 120.775 72.090 120.945 ;
        RECT 72.260 121.575 72.455 121.905 ;
        RECT 72.680 121.575 72.935 121.905 ;
        RECT 72.260 120.605 72.430 121.575 ;
        RECT 73.105 121.405 73.275 122.075 ;
        RECT 73.910 122.005 76.940 122.175 ;
        RECT 77.220 122.095 77.885 122.265 ;
        RECT 73.910 121.440 74.210 122.005 ;
        RECT 74.385 121.610 76.600 121.835 ;
        RECT 76.770 121.440 76.940 122.005 ;
        RECT 70.400 120.435 72.430 120.605 ;
        RECT 72.600 120.265 72.770 121.405 ;
        RECT 72.940 120.435 73.275 121.405 ;
        RECT 73.450 120.265 73.740 121.430 ;
        RECT 73.910 121.270 76.940 121.440 ;
        RECT 77.135 121.275 77.485 121.925 ;
        RECT 73.910 120.265 74.295 121.100 ;
        RECT 74.465 120.465 74.725 121.270 ;
        RECT 74.895 120.265 75.155 121.100 ;
        RECT 75.325 120.465 75.580 121.270 ;
        RECT 75.755 120.265 76.015 121.100 ;
        RECT 76.185 120.465 76.440 121.270 ;
        RECT 77.655 121.105 77.885 122.095 ;
        RECT 76.615 120.265 76.960 121.100 ;
        RECT 77.220 120.935 77.885 121.105 ;
        RECT 77.220 120.435 77.390 120.935 ;
        RECT 77.560 120.265 77.890 120.765 ;
        RECT 78.060 120.435 78.285 122.555 ;
        RECT 78.500 122.435 78.830 122.815 ;
        RECT 79.000 122.265 79.170 122.595 ;
        RECT 79.470 122.435 80.485 122.635 ;
        RECT 78.475 122.075 79.170 122.265 ;
        RECT 78.475 121.105 78.645 122.075 ;
        RECT 78.815 121.275 79.225 121.895 ;
        RECT 79.395 121.325 79.615 122.195 ;
        RECT 79.795 121.885 80.145 122.255 ;
        RECT 80.315 121.705 80.485 122.435 ;
        RECT 80.655 122.375 81.065 122.815 ;
        RECT 81.355 122.175 81.605 122.605 ;
        RECT 81.805 122.355 82.125 122.815 ;
        RECT 82.685 122.425 83.535 122.595 ;
        RECT 80.655 121.835 81.065 122.165 ;
        RECT 81.355 121.835 81.775 122.175 ;
        RECT 80.065 121.665 80.485 121.705 ;
        RECT 80.065 121.495 81.415 121.665 ;
        RECT 78.475 120.935 79.170 121.105 ;
        RECT 79.395 120.945 79.895 121.325 ;
        RECT 78.500 120.265 78.830 120.765 ;
        RECT 79.000 120.435 79.170 120.935 ;
        RECT 80.065 120.650 80.235 121.495 ;
        RECT 81.165 121.335 81.415 121.495 ;
        RECT 80.405 121.065 80.655 121.325 ;
        RECT 81.585 121.065 81.775 121.835 ;
        RECT 80.405 120.815 81.775 121.065 ;
        RECT 81.945 122.005 83.195 122.175 ;
        RECT 81.945 121.245 82.115 122.005 ;
        RECT 82.865 121.885 83.195 122.005 ;
        RECT 82.285 121.425 82.465 121.835 ;
        RECT 83.365 121.665 83.535 122.425 ;
        RECT 83.735 122.335 84.395 122.815 ;
        RECT 84.575 122.220 84.895 122.550 ;
        RECT 83.725 121.895 84.385 122.165 ;
        RECT 83.725 121.835 84.055 121.895 ;
        RECT 84.205 121.665 84.535 121.725 ;
        RECT 82.635 121.495 84.535 121.665 ;
        RECT 81.945 120.935 82.465 121.245 ;
        RECT 82.635 120.985 82.805 121.495 ;
        RECT 84.705 121.325 84.895 122.220 ;
        RECT 82.975 121.155 84.895 121.325 ;
        RECT 84.575 121.135 84.895 121.155 ;
        RECT 85.095 121.905 85.345 122.555 ;
        RECT 85.525 122.355 85.810 122.815 ;
        RECT 85.990 122.105 86.245 122.635 ;
        RECT 85.095 121.575 85.895 121.905 ;
        RECT 82.635 120.815 83.845 120.985 ;
        RECT 79.405 120.480 80.235 120.650 ;
        RECT 80.475 120.265 80.855 120.645 ;
        RECT 81.035 120.525 81.205 120.815 ;
        RECT 82.635 120.735 82.805 120.815 ;
        RECT 81.375 120.265 81.705 120.645 ;
        RECT 82.175 120.485 82.805 120.735 ;
        RECT 82.985 120.265 83.405 120.645 ;
        RECT 83.605 120.525 83.845 120.815 ;
        RECT 84.075 120.265 84.405 120.955 ;
        RECT 84.575 120.525 84.745 121.135 ;
        RECT 85.095 120.985 85.345 121.575 ;
        RECT 86.065 121.455 86.245 122.105 ;
        RECT 86.790 122.065 88.000 122.815 ;
        RECT 86.065 121.285 86.330 121.455 ;
        RECT 86.790 121.355 87.310 121.895 ;
        RECT 87.480 121.525 88.000 122.065 ;
        RECT 88.445 122.005 88.690 122.610 ;
        RECT 88.910 122.280 89.420 122.815 ;
        RECT 88.170 121.835 89.400 122.005 ;
        RECT 86.065 121.245 86.245 121.285 ;
        RECT 85.015 120.475 85.345 120.985 ;
        RECT 85.525 120.265 85.810 121.065 ;
        RECT 85.990 120.575 86.245 121.245 ;
        RECT 86.790 120.265 88.000 121.355 ;
        RECT 88.170 121.025 88.510 121.835 ;
        RECT 88.680 121.270 89.430 121.460 ;
        RECT 88.170 120.615 88.685 121.025 ;
        RECT 88.920 120.265 89.090 121.025 ;
        RECT 89.260 120.605 89.430 121.270 ;
        RECT 89.600 121.285 89.790 122.645 ;
        RECT 89.960 121.795 90.235 122.645 ;
        RECT 90.425 122.280 90.955 122.645 ;
        RECT 91.380 122.415 91.710 122.815 ;
        RECT 90.780 122.245 90.955 122.280 ;
        RECT 89.960 121.625 90.240 121.795 ;
        RECT 89.960 121.485 90.235 121.625 ;
        RECT 90.440 121.285 90.610 122.085 ;
        RECT 89.600 121.115 90.610 121.285 ;
        RECT 90.780 122.075 91.710 122.245 ;
        RECT 91.880 122.075 92.135 122.645 ;
        RECT 90.780 120.945 90.950 122.075 ;
        RECT 91.540 121.905 91.710 122.075 ;
        RECT 89.825 120.775 90.950 120.945 ;
        RECT 91.120 121.575 91.315 121.905 ;
        RECT 91.540 121.575 91.795 121.905 ;
        RECT 91.120 120.605 91.290 121.575 ;
        RECT 91.965 121.405 92.135 122.075 ;
        RECT 92.370 121.995 92.580 122.815 ;
        RECT 92.750 122.015 93.080 122.645 ;
        RECT 92.750 121.415 93.000 122.015 ;
        RECT 93.250 121.995 93.480 122.815 ;
        RECT 93.780 122.265 93.950 122.645 ;
        RECT 94.130 122.435 94.460 122.815 ;
        RECT 93.780 122.095 94.445 122.265 ;
        RECT 94.640 122.140 94.900 122.645 ;
        RECT 93.170 121.575 93.500 121.825 ;
        RECT 93.710 121.545 94.040 121.915 ;
        RECT 94.275 121.840 94.445 122.095 ;
        RECT 94.275 121.510 94.560 121.840 ;
        RECT 89.260 120.435 91.290 120.605 ;
        RECT 91.460 120.265 91.630 121.405 ;
        RECT 91.800 120.435 92.135 121.405 ;
        RECT 92.370 120.265 92.580 121.405 ;
        RECT 92.750 120.435 93.080 121.415 ;
        RECT 93.250 120.265 93.480 121.405 ;
        RECT 94.275 121.365 94.445 121.510 ;
        RECT 93.780 121.195 94.445 121.365 ;
        RECT 94.730 121.340 94.900 122.140 ;
        RECT 95.345 122.005 95.590 122.610 ;
        RECT 95.810 122.280 96.320 122.815 ;
        RECT 93.780 120.435 93.950 121.195 ;
        RECT 94.130 120.265 94.460 121.025 ;
        RECT 94.630 120.435 94.900 121.340 ;
        RECT 95.070 121.835 96.300 122.005 ;
        RECT 95.070 121.025 95.410 121.835 ;
        RECT 95.580 121.270 96.330 121.460 ;
        RECT 95.070 120.615 95.585 121.025 ;
        RECT 95.820 120.265 95.990 121.025 ;
        RECT 96.160 120.605 96.330 121.270 ;
        RECT 96.500 121.285 96.690 122.645 ;
        RECT 96.860 122.475 97.135 122.645 ;
        RECT 96.860 122.305 97.140 122.475 ;
        RECT 96.860 121.485 97.135 122.305 ;
        RECT 97.325 122.280 97.855 122.645 ;
        RECT 98.280 122.415 98.610 122.815 ;
        RECT 97.680 122.245 97.855 122.280 ;
        RECT 97.340 121.285 97.510 122.085 ;
        RECT 96.500 121.115 97.510 121.285 ;
        RECT 97.680 122.075 98.610 122.245 ;
        RECT 98.780 122.075 99.035 122.645 ;
        RECT 99.210 122.090 99.500 122.815 ;
        RECT 97.680 120.945 97.850 122.075 ;
        RECT 98.440 121.905 98.610 122.075 ;
        RECT 96.725 120.775 97.850 120.945 ;
        RECT 98.020 121.575 98.215 121.905 ;
        RECT 98.440 121.575 98.695 121.905 ;
        RECT 98.020 120.605 98.190 121.575 ;
        RECT 98.865 121.405 99.035 122.075 ;
        RECT 99.730 121.995 99.940 122.815 ;
        RECT 100.110 122.015 100.440 122.645 ;
        RECT 96.160 120.435 98.190 120.605 ;
        RECT 98.360 120.265 98.530 121.405 ;
        RECT 98.700 120.435 99.035 121.405 ;
        RECT 99.210 120.265 99.500 121.430 ;
        RECT 100.110 121.415 100.360 122.015 ;
        RECT 100.610 121.995 100.840 122.815 ;
        RECT 101.425 122.475 101.680 122.635 ;
        RECT 101.340 122.305 101.680 122.475 ;
        RECT 101.860 122.355 102.145 122.815 ;
        RECT 101.425 122.105 101.680 122.305 ;
        RECT 100.530 121.575 100.860 121.825 ;
        RECT 99.730 120.265 99.940 121.405 ;
        RECT 100.110 120.435 100.440 121.415 ;
        RECT 100.610 120.265 100.840 121.405 ;
        RECT 101.425 121.245 101.605 122.105 ;
        RECT 102.325 121.905 102.575 122.555 ;
        RECT 101.775 121.575 102.575 121.905 ;
        RECT 101.425 120.575 101.680 121.245 ;
        RECT 101.860 120.265 102.145 121.065 ;
        RECT 102.325 120.985 102.575 121.575 ;
        RECT 102.775 122.220 103.095 122.550 ;
        RECT 103.275 122.335 103.935 122.815 ;
        RECT 104.135 122.425 104.985 122.595 ;
        RECT 102.775 121.325 102.965 122.220 ;
        RECT 103.285 121.895 103.945 122.165 ;
        RECT 103.615 121.835 103.945 121.895 ;
        RECT 103.135 121.665 103.465 121.725 ;
        RECT 104.135 121.665 104.305 122.425 ;
        RECT 105.545 122.355 105.865 122.815 ;
        RECT 106.065 122.175 106.315 122.605 ;
        RECT 106.605 122.375 107.015 122.815 ;
        RECT 107.185 122.435 108.200 122.635 ;
        RECT 104.475 122.005 105.725 122.175 ;
        RECT 104.475 121.885 104.805 122.005 ;
        RECT 103.135 121.495 105.035 121.665 ;
        RECT 102.775 121.155 104.695 121.325 ;
        RECT 102.775 121.135 103.095 121.155 ;
        RECT 102.325 120.475 102.655 120.985 ;
        RECT 102.925 120.525 103.095 121.135 ;
        RECT 104.865 120.985 105.035 121.495 ;
        RECT 105.205 121.425 105.385 121.835 ;
        RECT 105.555 121.245 105.725 122.005 ;
        RECT 103.265 120.265 103.595 120.955 ;
        RECT 103.825 120.815 105.035 120.985 ;
        RECT 105.205 120.935 105.725 121.245 ;
        RECT 105.895 121.835 106.315 122.175 ;
        RECT 106.605 121.835 107.015 122.165 ;
        RECT 105.895 121.065 106.085 121.835 ;
        RECT 107.185 121.705 107.355 122.435 ;
        RECT 108.500 122.265 108.670 122.595 ;
        RECT 108.840 122.435 109.170 122.815 ;
        RECT 107.525 121.885 107.875 122.255 ;
        RECT 107.185 121.665 107.605 121.705 ;
        RECT 106.255 121.495 107.605 121.665 ;
        RECT 106.255 121.335 106.505 121.495 ;
        RECT 107.015 121.065 107.265 121.325 ;
        RECT 105.895 120.815 107.265 121.065 ;
        RECT 103.825 120.525 104.065 120.815 ;
        RECT 104.865 120.735 105.035 120.815 ;
        RECT 104.265 120.265 104.685 120.645 ;
        RECT 104.865 120.485 105.495 120.735 ;
        RECT 105.965 120.265 106.295 120.645 ;
        RECT 106.465 120.525 106.635 120.815 ;
        RECT 107.435 120.650 107.605 121.495 ;
        RECT 108.055 121.325 108.275 122.195 ;
        RECT 108.500 122.075 109.195 122.265 ;
        RECT 107.775 120.945 108.275 121.325 ;
        RECT 108.445 121.275 108.855 121.895 ;
        RECT 109.025 121.105 109.195 122.075 ;
        RECT 108.500 120.935 109.195 121.105 ;
        RECT 106.815 120.265 107.195 120.645 ;
        RECT 107.435 120.480 108.265 120.650 ;
        RECT 108.500 120.435 108.670 120.935 ;
        RECT 108.840 120.265 109.170 120.765 ;
        RECT 109.385 120.435 109.610 122.555 ;
        RECT 109.780 122.435 110.110 122.815 ;
        RECT 110.280 122.265 110.450 122.555 ;
        RECT 109.785 122.095 110.450 122.265 ;
        RECT 109.785 121.105 110.015 122.095 ;
        RECT 111.170 122.065 112.380 122.815 ;
        RECT 110.185 121.275 110.535 121.925 ;
        RECT 111.170 121.355 111.690 121.895 ;
        RECT 111.860 121.525 112.380 122.065 ;
        RECT 109.785 120.935 110.450 121.105 ;
        RECT 109.780 120.265 110.110 120.765 ;
        RECT 110.280 120.435 110.450 120.935 ;
        RECT 111.170 120.265 112.380 121.355 ;
        RECT 18.165 120.095 112.465 120.265 ;
        RECT 18.250 119.005 19.460 120.095 ;
        RECT 18.250 118.295 18.770 118.835 ;
        RECT 18.940 118.465 19.460 119.005 ;
        RECT 19.630 119.005 21.300 120.095 ;
        RECT 19.630 118.485 20.380 119.005 ;
        RECT 21.510 118.955 21.740 120.095 ;
        RECT 21.910 118.945 22.240 119.925 ;
        RECT 22.410 118.955 22.620 120.095 ;
        RECT 22.855 118.955 23.190 119.925 ;
        RECT 23.360 118.955 23.530 120.095 ;
        RECT 23.700 119.755 25.730 119.925 ;
        RECT 20.550 118.315 21.300 118.835 ;
        RECT 21.490 118.535 21.820 118.785 ;
        RECT 18.250 117.545 19.460 118.295 ;
        RECT 19.630 117.545 21.300 118.315 ;
        RECT 21.510 117.545 21.740 118.365 ;
        RECT 21.990 118.345 22.240 118.945 ;
        RECT 21.910 117.715 22.240 118.345 ;
        RECT 22.410 117.545 22.620 118.365 ;
        RECT 22.855 118.285 23.025 118.955 ;
        RECT 23.700 118.785 23.870 119.755 ;
        RECT 23.195 118.455 23.450 118.785 ;
        RECT 23.675 118.455 23.870 118.785 ;
        RECT 24.040 119.415 25.165 119.585 ;
        RECT 23.280 118.285 23.450 118.455 ;
        RECT 24.040 118.285 24.210 119.415 ;
        RECT 22.855 117.715 23.110 118.285 ;
        RECT 23.280 118.115 24.210 118.285 ;
        RECT 24.380 119.075 25.390 119.245 ;
        RECT 24.380 118.275 24.550 119.075 ;
        RECT 24.755 118.735 25.030 118.875 ;
        RECT 24.750 118.565 25.030 118.735 ;
        RECT 24.035 118.080 24.210 118.115 ;
        RECT 23.280 117.545 23.610 117.945 ;
        RECT 24.035 117.715 24.565 118.080 ;
        RECT 24.755 117.715 25.030 118.565 ;
        RECT 25.200 117.715 25.390 119.075 ;
        RECT 25.560 119.090 25.730 119.755 ;
        RECT 25.900 119.335 26.070 120.095 ;
        RECT 26.305 119.335 26.820 119.745 ;
        RECT 25.560 118.900 26.310 119.090 ;
        RECT 26.480 118.525 26.820 119.335 ;
        RECT 25.590 118.355 26.820 118.525 ;
        RECT 26.990 119.335 27.505 119.745 ;
        RECT 27.740 119.335 27.910 120.095 ;
        RECT 28.080 119.755 30.110 119.925 ;
        RECT 26.990 118.525 27.330 119.335 ;
        RECT 28.080 119.090 28.250 119.755 ;
        RECT 28.645 119.415 29.770 119.585 ;
        RECT 27.500 118.900 28.250 119.090 ;
        RECT 28.420 119.075 29.430 119.245 ;
        RECT 26.990 118.355 28.220 118.525 ;
        RECT 25.570 117.545 26.080 118.080 ;
        RECT 26.300 117.750 26.545 118.355 ;
        RECT 27.265 117.750 27.510 118.355 ;
        RECT 27.730 117.545 28.240 118.080 ;
        RECT 28.420 117.715 28.610 119.075 ;
        RECT 28.780 118.735 29.055 118.875 ;
        RECT 28.780 118.565 29.060 118.735 ;
        RECT 28.780 117.715 29.055 118.565 ;
        RECT 29.260 118.275 29.430 119.075 ;
        RECT 29.600 118.285 29.770 119.415 ;
        RECT 29.940 118.785 30.110 119.755 ;
        RECT 30.280 118.955 30.450 120.095 ;
        RECT 30.620 118.955 30.955 119.925 ;
        RECT 31.170 118.955 31.400 120.095 ;
        RECT 29.940 118.455 30.135 118.785 ;
        RECT 30.360 118.455 30.615 118.785 ;
        RECT 30.360 118.285 30.530 118.455 ;
        RECT 30.785 118.285 30.955 118.955 ;
        RECT 31.570 118.945 31.900 119.925 ;
        RECT 32.070 118.955 32.280 120.095 ;
        RECT 32.710 119.425 32.990 120.095 ;
        RECT 33.160 119.205 33.460 119.755 ;
        RECT 33.660 119.375 33.990 120.095 ;
        RECT 34.180 119.375 34.640 119.925 ;
        RECT 31.150 118.535 31.480 118.785 ;
        RECT 29.600 118.115 30.530 118.285 ;
        RECT 29.600 118.080 29.775 118.115 ;
        RECT 29.245 117.715 29.775 118.080 ;
        RECT 30.200 117.545 30.530 117.945 ;
        RECT 30.700 117.715 30.955 118.285 ;
        RECT 31.170 117.545 31.400 118.365 ;
        RECT 31.650 118.345 31.900 118.945 ;
        RECT 32.525 118.785 32.790 119.145 ;
        RECT 33.160 119.035 34.100 119.205 ;
        RECT 33.930 118.785 34.100 119.035 ;
        RECT 32.525 118.535 33.200 118.785 ;
        RECT 33.420 118.535 33.760 118.785 ;
        RECT 33.930 118.455 34.220 118.785 ;
        RECT 33.930 118.365 34.100 118.455 ;
        RECT 31.570 117.715 31.900 118.345 ;
        RECT 32.070 117.545 32.280 118.365 ;
        RECT 32.710 118.175 34.100 118.365 ;
        RECT 32.710 117.815 33.040 118.175 ;
        RECT 34.390 118.005 34.640 119.375 ;
        RECT 34.810 118.930 35.100 120.095 ;
        RECT 35.930 119.425 36.210 120.095 ;
        RECT 36.380 119.205 36.680 119.755 ;
        RECT 36.880 119.375 37.210 120.095 ;
        RECT 37.400 119.375 37.860 119.925 ;
        RECT 39.150 119.425 39.430 120.095 ;
        RECT 35.745 118.785 36.010 119.145 ;
        RECT 36.380 119.035 37.320 119.205 ;
        RECT 37.150 118.785 37.320 119.035 ;
        RECT 35.745 118.535 36.420 118.785 ;
        RECT 36.640 118.535 36.980 118.785 ;
        RECT 37.150 118.455 37.440 118.785 ;
        RECT 37.150 118.365 37.320 118.455 ;
        RECT 33.660 117.545 33.910 118.005 ;
        RECT 34.080 117.715 34.640 118.005 ;
        RECT 34.810 117.545 35.100 118.270 ;
        RECT 35.930 118.175 37.320 118.365 ;
        RECT 35.930 117.815 36.260 118.175 ;
        RECT 37.610 118.005 37.860 119.375 ;
        RECT 39.600 119.205 39.900 119.755 ;
        RECT 40.100 119.375 40.430 120.095 ;
        RECT 40.620 119.375 41.080 119.925 ;
        RECT 38.965 118.785 39.230 119.145 ;
        RECT 39.600 119.035 40.540 119.205 ;
        RECT 40.370 118.785 40.540 119.035 ;
        RECT 38.965 118.535 39.640 118.785 ;
        RECT 39.860 118.535 40.200 118.785 ;
        RECT 40.370 118.455 40.660 118.785 ;
        RECT 40.370 118.365 40.540 118.455 ;
        RECT 36.880 117.545 37.130 118.005 ;
        RECT 37.300 117.715 37.860 118.005 ;
        RECT 39.150 118.175 40.540 118.365 ;
        RECT 39.150 117.815 39.480 118.175 ;
        RECT 40.830 118.005 41.080 119.375 ;
        RECT 40.100 117.545 40.350 118.005 ;
        RECT 40.520 117.715 41.080 118.005 ;
        RECT 41.250 119.375 41.710 119.925 ;
        RECT 41.900 119.375 42.230 120.095 ;
        RECT 41.250 118.005 41.500 119.375 ;
        RECT 42.430 119.205 42.730 119.755 ;
        RECT 42.900 119.425 43.180 120.095 ;
        RECT 41.790 119.035 42.730 119.205 ;
        RECT 43.550 119.335 44.065 119.745 ;
        RECT 44.300 119.335 44.470 120.095 ;
        RECT 44.640 119.755 46.670 119.925 ;
        RECT 41.790 118.785 41.960 119.035 ;
        RECT 43.100 118.785 43.365 119.145 ;
        RECT 41.670 118.455 41.960 118.785 ;
        RECT 42.130 118.535 42.470 118.785 ;
        RECT 42.690 118.535 43.365 118.785 ;
        RECT 41.790 118.365 41.960 118.455 ;
        RECT 43.550 118.525 43.890 119.335 ;
        RECT 44.640 119.090 44.810 119.755 ;
        RECT 45.205 119.415 46.330 119.585 ;
        RECT 44.060 118.900 44.810 119.090 ;
        RECT 44.980 119.075 45.990 119.245 ;
        RECT 41.790 118.175 43.180 118.365 ;
        RECT 43.550 118.355 44.780 118.525 ;
        RECT 41.250 117.715 41.810 118.005 ;
        RECT 41.980 117.545 42.230 118.005 ;
        RECT 42.850 117.815 43.180 118.175 ;
        RECT 43.825 117.750 44.070 118.355 ;
        RECT 44.290 117.545 44.800 118.080 ;
        RECT 44.980 117.715 45.170 119.075 ;
        RECT 45.340 118.055 45.615 118.875 ;
        RECT 45.820 118.275 45.990 119.075 ;
        RECT 46.160 118.285 46.330 119.415 ;
        RECT 46.500 118.785 46.670 119.755 ;
        RECT 46.840 118.955 47.010 120.095 ;
        RECT 47.180 118.955 47.515 119.925 ;
        RECT 46.500 118.455 46.695 118.785 ;
        RECT 46.920 118.455 47.175 118.785 ;
        RECT 46.920 118.285 47.090 118.455 ;
        RECT 47.345 118.285 47.515 118.955 ;
        RECT 48.150 119.335 48.665 119.745 ;
        RECT 48.900 119.335 49.070 120.095 ;
        RECT 49.240 119.755 51.270 119.925 ;
        RECT 48.150 118.525 48.490 119.335 ;
        RECT 49.240 119.090 49.410 119.755 ;
        RECT 49.805 119.415 50.930 119.585 ;
        RECT 48.660 118.900 49.410 119.090 ;
        RECT 49.580 119.075 50.590 119.245 ;
        RECT 48.150 118.355 49.380 118.525 ;
        RECT 46.160 118.115 47.090 118.285 ;
        RECT 46.160 118.080 46.335 118.115 ;
        RECT 45.340 117.885 45.620 118.055 ;
        RECT 45.340 117.715 45.615 117.885 ;
        RECT 45.805 117.715 46.335 118.080 ;
        RECT 46.760 117.545 47.090 117.945 ;
        RECT 47.260 117.715 47.515 118.285 ;
        RECT 48.425 117.750 48.670 118.355 ;
        RECT 48.890 117.545 49.400 118.080 ;
        RECT 49.580 117.715 49.770 119.075 ;
        RECT 49.940 118.395 50.215 118.875 ;
        RECT 49.940 118.225 50.220 118.395 ;
        RECT 50.420 118.275 50.590 119.075 ;
        RECT 50.760 118.285 50.930 119.415 ;
        RECT 51.100 118.785 51.270 119.755 ;
        RECT 51.440 118.955 51.610 120.095 ;
        RECT 51.780 118.955 52.115 119.925 ;
        RECT 52.380 119.165 52.550 119.925 ;
        RECT 52.730 119.335 53.060 120.095 ;
        RECT 52.380 118.995 53.045 119.165 ;
        RECT 53.230 119.020 53.500 119.925 ;
        RECT 51.100 118.455 51.295 118.785 ;
        RECT 51.520 118.455 51.775 118.785 ;
        RECT 51.520 118.285 51.690 118.455 ;
        RECT 51.945 118.285 52.115 118.955 ;
        RECT 52.875 118.850 53.045 118.995 ;
        RECT 52.310 118.445 52.640 118.815 ;
        RECT 52.875 118.520 53.160 118.850 ;
        RECT 49.940 117.715 50.215 118.225 ;
        RECT 50.760 118.115 51.690 118.285 ;
        RECT 50.760 118.080 50.935 118.115 ;
        RECT 50.405 117.715 50.935 118.080 ;
        RECT 51.360 117.545 51.690 117.945 ;
        RECT 51.860 117.715 52.115 118.285 ;
        RECT 52.875 118.265 53.045 118.520 ;
        RECT 52.380 118.095 53.045 118.265 ;
        RECT 53.330 118.220 53.500 119.020 ;
        RECT 53.760 119.165 53.930 119.925 ;
        RECT 54.110 119.335 54.440 120.095 ;
        RECT 53.760 118.995 54.425 119.165 ;
        RECT 54.610 119.020 54.880 119.925 ;
        RECT 54.255 118.850 54.425 118.995 ;
        RECT 53.690 118.445 54.020 118.815 ;
        RECT 54.255 118.520 54.540 118.850 ;
        RECT 54.255 118.265 54.425 118.520 ;
        RECT 52.380 117.715 52.550 118.095 ;
        RECT 52.730 117.545 53.060 117.925 ;
        RECT 53.240 117.715 53.500 118.220 ;
        RECT 53.760 118.095 54.425 118.265 ;
        RECT 54.710 118.220 54.880 119.020 ;
        RECT 55.090 118.955 55.320 120.095 ;
        RECT 55.490 118.945 55.820 119.925 ;
        RECT 55.990 118.955 56.200 120.095 ;
        RECT 56.430 119.335 56.945 119.745 ;
        RECT 57.180 119.335 57.350 120.095 ;
        RECT 57.520 119.755 59.550 119.925 ;
        RECT 55.070 118.535 55.400 118.785 ;
        RECT 53.760 117.715 53.930 118.095 ;
        RECT 54.110 117.545 54.440 117.925 ;
        RECT 54.620 117.715 54.880 118.220 ;
        RECT 55.090 117.545 55.320 118.365 ;
        RECT 55.570 118.345 55.820 118.945 ;
        RECT 56.430 118.525 56.770 119.335 ;
        RECT 57.520 119.090 57.690 119.755 ;
        RECT 58.085 119.415 59.210 119.585 ;
        RECT 56.940 118.900 57.690 119.090 ;
        RECT 57.860 119.075 58.870 119.245 ;
        RECT 55.490 117.715 55.820 118.345 ;
        RECT 55.990 117.545 56.200 118.365 ;
        RECT 56.430 118.355 57.660 118.525 ;
        RECT 56.705 117.750 56.950 118.355 ;
        RECT 57.170 117.545 57.680 118.080 ;
        RECT 57.860 117.715 58.050 119.075 ;
        RECT 58.220 118.735 58.495 118.875 ;
        RECT 58.220 118.565 58.500 118.735 ;
        RECT 58.220 117.715 58.495 118.565 ;
        RECT 58.700 118.275 58.870 119.075 ;
        RECT 59.040 118.285 59.210 119.415 ;
        RECT 59.380 118.785 59.550 119.755 ;
        RECT 59.720 118.955 59.890 120.095 ;
        RECT 60.060 118.955 60.395 119.925 ;
        RECT 59.380 118.455 59.575 118.785 ;
        RECT 59.800 118.455 60.055 118.785 ;
        RECT 59.800 118.285 59.970 118.455 ;
        RECT 60.225 118.285 60.395 118.955 ;
        RECT 60.570 118.930 60.860 120.095 ;
        RECT 61.035 118.955 61.370 119.925 ;
        RECT 61.540 118.955 61.710 120.095 ;
        RECT 61.880 119.755 63.910 119.925 ;
        RECT 59.040 118.115 59.970 118.285 ;
        RECT 59.040 118.080 59.215 118.115 ;
        RECT 58.685 117.715 59.215 118.080 ;
        RECT 59.640 117.545 59.970 117.945 ;
        RECT 60.140 117.715 60.395 118.285 ;
        RECT 61.035 118.285 61.205 118.955 ;
        RECT 61.880 118.785 62.050 119.755 ;
        RECT 61.375 118.455 61.630 118.785 ;
        RECT 61.855 118.455 62.050 118.785 ;
        RECT 62.220 119.415 63.345 119.585 ;
        RECT 61.460 118.285 61.630 118.455 ;
        RECT 62.220 118.285 62.390 119.415 ;
        RECT 60.570 117.545 60.860 118.270 ;
        RECT 61.035 117.715 61.290 118.285 ;
        RECT 61.460 118.115 62.390 118.285 ;
        RECT 62.560 119.075 63.570 119.245 ;
        RECT 62.560 118.275 62.730 119.075 ;
        RECT 62.935 118.395 63.210 118.875 ;
        RECT 62.930 118.225 63.210 118.395 ;
        RECT 62.215 118.080 62.390 118.115 ;
        RECT 61.460 117.545 61.790 117.945 ;
        RECT 62.215 117.715 62.745 118.080 ;
        RECT 62.935 117.715 63.210 118.225 ;
        RECT 63.380 117.715 63.570 119.075 ;
        RECT 63.740 119.090 63.910 119.755 ;
        RECT 64.080 119.335 64.250 120.095 ;
        RECT 64.485 119.335 65.000 119.745 ;
        RECT 63.740 118.900 64.490 119.090 ;
        RECT 64.660 118.525 65.000 119.335 ;
        RECT 65.210 118.955 65.440 120.095 ;
        RECT 65.610 118.945 65.940 119.925 ;
        RECT 66.110 118.955 66.320 120.095 ;
        RECT 66.610 118.955 66.820 120.095 ;
        RECT 65.190 118.535 65.520 118.785 ;
        RECT 63.770 118.355 65.000 118.525 ;
        RECT 63.750 117.545 64.260 118.080 ;
        RECT 64.480 117.750 64.725 118.355 ;
        RECT 65.210 117.545 65.440 118.365 ;
        RECT 65.690 118.345 65.940 118.945 ;
        RECT 66.990 118.945 67.320 119.925 ;
        RECT 67.490 118.955 67.720 120.095 ;
        RECT 69.225 119.755 69.480 119.785 ;
        RECT 69.140 119.585 69.480 119.755 ;
        RECT 69.225 119.115 69.480 119.585 ;
        RECT 69.660 119.295 69.945 120.095 ;
        RECT 70.125 119.375 70.455 119.885 ;
        RECT 65.610 117.715 65.940 118.345 ;
        RECT 66.110 117.545 66.320 118.365 ;
        RECT 66.610 117.545 66.820 118.365 ;
        RECT 66.990 118.345 67.240 118.945 ;
        RECT 67.410 118.535 67.740 118.785 ;
        RECT 66.990 117.715 67.320 118.345 ;
        RECT 67.490 117.545 67.720 118.365 ;
        RECT 69.225 118.255 69.405 119.115 ;
        RECT 70.125 118.785 70.375 119.375 ;
        RECT 70.725 119.225 70.895 119.835 ;
        RECT 71.065 119.405 71.395 120.095 ;
        RECT 71.625 119.545 71.865 119.835 ;
        RECT 72.065 119.715 72.485 120.095 ;
        RECT 72.665 119.625 73.295 119.875 ;
        RECT 73.765 119.715 74.095 120.095 ;
        RECT 72.665 119.545 72.835 119.625 ;
        RECT 74.265 119.545 74.435 119.835 ;
        RECT 74.615 119.715 74.995 120.095 ;
        RECT 75.235 119.710 76.065 119.880 ;
        RECT 71.625 119.375 72.835 119.545 ;
        RECT 69.575 118.455 70.375 118.785 ;
        RECT 69.225 117.725 69.480 118.255 ;
        RECT 69.660 117.545 69.945 118.005 ;
        RECT 70.125 117.805 70.375 118.455 ;
        RECT 70.575 119.205 70.895 119.225 ;
        RECT 70.575 119.035 72.495 119.205 ;
        RECT 70.575 118.140 70.765 119.035 ;
        RECT 72.665 118.865 72.835 119.375 ;
        RECT 73.005 119.115 73.525 119.425 ;
        RECT 70.935 118.695 72.835 118.865 ;
        RECT 70.935 118.635 71.265 118.695 ;
        RECT 71.415 118.465 71.745 118.525 ;
        RECT 71.085 118.195 71.745 118.465 ;
        RECT 70.575 117.810 70.895 118.140 ;
        RECT 71.075 117.545 71.735 118.025 ;
        RECT 71.935 117.935 72.105 118.695 ;
        RECT 73.005 118.525 73.185 118.935 ;
        RECT 72.275 118.355 72.605 118.475 ;
        RECT 73.355 118.355 73.525 119.115 ;
        RECT 72.275 118.185 73.525 118.355 ;
        RECT 73.695 119.295 75.065 119.545 ;
        RECT 73.695 118.525 73.885 119.295 ;
        RECT 74.815 119.035 75.065 119.295 ;
        RECT 74.055 118.865 74.305 119.025 ;
        RECT 75.235 118.865 75.405 119.710 ;
        RECT 76.300 119.425 76.470 119.925 ;
        RECT 76.640 119.595 76.970 120.095 ;
        RECT 75.575 119.035 76.075 119.415 ;
        RECT 76.300 119.255 76.995 119.425 ;
        RECT 74.055 118.695 75.405 118.865 ;
        RECT 74.985 118.655 75.405 118.695 ;
        RECT 73.695 118.185 74.115 118.525 ;
        RECT 74.405 118.195 74.815 118.525 ;
        RECT 71.935 117.765 72.785 117.935 ;
        RECT 73.345 117.545 73.665 118.005 ;
        RECT 73.865 117.755 74.115 118.185 ;
        RECT 74.405 117.545 74.815 117.985 ;
        RECT 74.985 117.925 75.155 118.655 ;
        RECT 75.325 118.105 75.675 118.475 ;
        RECT 75.855 118.165 76.075 119.035 ;
        RECT 76.245 118.465 76.655 119.085 ;
        RECT 76.825 118.285 76.995 119.255 ;
        RECT 76.300 118.095 76.995 118.285 ;
        RECT 74.985 117.725 76.000 117.925 ;
        RECT 76.300 117.765 76.470 118.095 ;
        RECT 76.640 117.545 76.970 117.925 ;
        RECT 77.185 117.805 77.410 119.925 ;
        RECT 77.580 119.595 77.910 120.095 ;
        RECT 78.080 119.425 78.250 119.925 ;
        RECT 77.585 119.255 78.250 119.425 ;
        RECT 78.510 119.375 78.970 119.925 ;
        RECT 79.160 119.375 79.490 120.095 ;
        RECT 77.585 118.265 77.815 119.255 ;
        RECT 77.985 118.435 78.335 119.085 ;
        RECT 77.585 118.095 78.250 118.265 ;
        RECT 77.580 117.545 77.910 117.925 ;
        RECT 78.080 117.805 78.250 118.095 ;
        RECT 78.510 118.005 78.760 119.375 ;
        RECT 79.690 119.205 79.990 119.755 ;
        RECT 80.160 119.425 80.440 120.095 ;
        RECT 79.050 119.035 79.990 119.205 ;
        RECT 79.050 118.785 79.220 119.035 ;
        RECT 80.360 118.785 80.625 119.145 ;
        RECT 78.930 118.455 79.220 118.785 ;
        RECT 79.390 118.535 79.730 118.785 ;
        RECT 79.950 118.535 80.625 118.785 ;
        RECT 80.810 119.020 81.080 119.925 ;
        RECT 81.250 119.335 81.580 120.095 ;
        RECT 81.760 119.165 81.930 119.925 ;
        RECT 79.050 118.365 79.220 118.455 ;
        RECT 79.050 118.175 80.440 118.365 ;
        RECT 78.510 117.715 79.070 118.005 ;
        RECT 79.240 117.545 79.490 118.005 ;
        RECT 80.110 117.815 80.440 118.175 ;
        RECT 80.810 118.220 80.980 119.020 ;
        RECT 81.265 118.995 81.930 119.165 ;
        RECT 82.190 119.335 82.705 119.745 ;
        RECT 82.940 119.335 83.110 120.095 ;
        RECT 83.280 119.755 85.310 119.925 ;
        RECT 81.265 118.850 81.435 118.995 ;
        RECT 81.150 118.520 81.435 118.850 ;
        RECT 81.265 118.265 81.435 118.520 ;
        RECT 81.670 118.445 82.000 118.815 ;
        RECT 82.190 118.525 82.530 119.335 ;
        RECT 83.280 119.090 83.450 119.755 ;
        RECT 83.845 119.415 84.970 119.585 ;
        RECT 82.700 118.900 83.450 119.090 ;
        RECT 83.620 119.075 84.630 119.245 ;
        RECT 82.190 118.355 83.420 118.525 ;
        RECT 80.810 117.715 81.070 118.220 ;
        RECT 81.265 118.095 81.930 118.265 ;
        RECT 81.250 117.545 81.580 117.925 ;
        RECT 81.760 117.715 81.930 118.095 ;
        RECT 82.465 117.750 82.710 118.355 ;
        RECT 82.930 117.545 83.440 118.080 ;
        RECT 83.620 117.715 83.810 119.075 ;
        RECT 83.980 118.055 84.255 118.875 ;
        RECT 84.460 118.275 84.630 119.075 ;
        RECT 84.800 118.285 84.970 119.415 ;
        RECT 85.140 118.785 85.310 119.755 ;
        RECT 85.480 118.955 85.650 120.095 ;
        RECT 85.820 118.955 86.155 119.925 ;
        RECT 85.140 118.455 85.335 118.785 ;
        RECT 85.560 118.455 85.815 118.785 ;
        RECT 85.560 118.285 85.730 118.455 ;
        RECT 85.985 118.285 86.155 118.955 ;
        RECT 86.330 118.930 86.620 120.095 ;
        RECT 88.085 119.755 88.340 119.785 ;
        RECT 88.000 119.585 88.340 119.755 ;
        RECT 88.085 119.115 88.340 119.585 ;
        RECT 88.520 119.295 88.805 120.095 ;
        RECT 88.985 119.375 89.315 119.885 ;
        RECT 84.800 118.115 85.730 118.285 ;
        RECT 84.800 118.080 84.975 118.115 ;
        RECT 83.980 117.885 84.260 118.055 ;
        RECT 83.980 117.715 84.255 117.885 ;
        RECT 84.445 117.715 84.975 118.080 ;
        RECT 85.400 117.545 85.730 117.945 ;
        RECT 85.900 117.715 86.155 118.285 ;
        RECT 86.330 117.545 86.620 118.270 ;
        RECT 88.085 118.255 88.265 119.115 ;
        RECT 88.985 118.785 89.235 119.375 ;
        RECT 89.585 119.225 89.755 119.835 ;
        RECT 89.925 119.405 90.255 120.095 ;
        RECT 90.485 119.545 90.725 119.835 ;
        RECT 90.925 119.715 91.345 120.095 ;
        RECT 91.525 119.625 92.155 119.875 ;
        RECT 92.625 119.715 92.955 120.095 ;
        RECT 91.525 119.545 91.695 119.625 ;
        RECT 93.125 119.545 93.295 119.835 ;
        RECT 93.475 119.715 93.855 120.095 ;
        RECT 94.095 119.710 94.925 119.880 ;
        RECT 90.485 119.375 91.695 119.545 ;
        RECT 88.435 118.455 89.235 118.785 ;
        RECT 88.085 117.725 88.340 118.255 ;
        RECT 88.520 117.545 88.805 118.005 ;
        RECT 88.985 117.805 89.235 118.455 ;
        RECT 89.435 119.205 89.755 119.225 ;
        RECT 89.435 119.035 91.355 119.205 ;
        RECT 89.435 118.140 89.625 119.035 ;
        RECT 91.525 118.865 91.695 119.375 ;
        RECT 91.865 119.115 92.385 119.425 ;
        RECT 89.795 118.695 91.695 118.865 ;
        RECT 89.795 118.635 90.125 118.695 ;
        RECT 90.275 118.465 90.605 118.525 ;
        RECT 89.945 118.195 90.605 118.465 ;
        RECT 89.435 117.810 89.755 118.140 ;
        RECT 89.935 117.545 90.595 118.025 ;
        RECT 90.795 117.935 90.965 118.695 ;
        RECT 91.865 118.525 92.045 118.935 ;
        RECT 91.135 118.355 91.465 118.475 ;
        RECT 92.215 118.355 92.385 119.115 ;
        RECT 91.135 118.185 92.385 118.355 ;
        RECT 92.555 119.295 93.925 119.545 ;
        RECT 92.555 118.525 92.745 119.295 ;
        RECT 93.675 119.035 93.925 119.295 ;
        RECT 92.915 118.865 93.165 119.025 ;
        RECT 94.095 118.865 94.265 119.710 ;
        RECT 95.160 119.425 95.330 119.925 ;
        RECT 95.500 119.595 95.830 120.095 ;
        RECT 94.435 119.035 94.935 119.415 ;
        RECT 95.160 119.255 95.855 119.425 ;
        RECT 92.915 118.695 94.265 118.865 ;
        RECT 93.845 118.655 94.265 118.695 ;
        RECT 92.555 118.185 92.975 118.525 ;
        RECT 93.265 118.195 93.675 118.525 ;
        RECT 90.795 117.765 91.645 117.935 ;
        RECT 92.205 117.545 92.525 118.005 ;
        RECT 92.725 117.755 92.975 118.185 ;
        RECT 93.265 117.545 93.675 117.985 ;
        RECT 93.845 117.925 94.015 118.655 ;
        RECT 94.185 118.105 94.535 118.475 ;
        RECT 94.715 118.165 94.935 119.035 ;
        RECT 95.105 118.465 95.515 119.085 ;
        RECT 95.685 118.285 95.855 119.255 ;
        RECT 95.160 118.095 95.855 118.285 ;
        RECT 93.845 117.725 94.860 117.925 ;
        RECT 95.160 117.765 95.330 118.095 ;
        RECT 95.500 117.545 95.830 117.925 ;
        RECT 96.045 117.805 96.270 119.925 ;
        RECT 96.440 119.595 96.770 120.095 ;
        RECT 96.940 119.425 97.110 119.925 ;
        RECT 96.445 119.255 97.110 119.425 ;
        RECT 97.370 119.335 97.885 119.745 ;
        RECT 98.120 119.335 98.290 120.095 ;
        RECT 98.460 119.755 100.490 119.925 ;
        RECT 96.445 118.265 96.675 119.255 ;
        RECT 96.845 118.435 97.195 119.085 ;
        RECT 97.370 118.525 97.710 119.335 ;
        RECT 98.460 119.090 98.630 119.755 ;
        RECT 99.025 119.415 100.150 119.585 ;
        RECT 97.880 118.900 98.630 119.090 ;
        RECT 98.800 119.075 99.810 119.245 ;
        RECT 97.370 118.355 98.600 118.525 ;
        RECT 96.445 118.095 97.110 118.265 ;
        RECT 96.440 117.545 96.770 117.925 ;
        RECT 96.940 117.805 97.110 118.095 ;
        RECT 97.645 117.750 97.890 118.355 ;
        RECT 98.110 117.545 98.620 118.080 ;
        RECT 98.800 117.715 98.990 119.075 ;
        RECT 99.160 118.055 99.435 118.875 ;
        RECT 99.640 118.275 99.810 119.075 ;
        RECT 99.980 118.285 100.150 119.415 ;
        RECT 100.320 118.785 100.490 119.755 ;
        RECT 100.660 118.955 100.830 120.095 ;
        RECT 101.000 118.955 101.335 119.925 ;
        RECT 100.320 118.455 100.515 118.785 ;
        RECT 100.740 118.455 100.995 118.785 ;
        RECT 100.740 118.285 100.910 118.455 ;
        RECT 101.165 118.285 101.335 118.955 ;
        RECT 101.510 119.335 102.025 119.745 ;
        RECT 102.260 119.335 102.430 120.095 ;
        RECT 102.600 119.755 104.630 119.925 ;
        RECT 101.510 118.525 101.850 119.335 ;
        RECT 102.600 119.090 102.770 119.755 ;
        RECT 103.165 119.415 104.290 119.585 ;
        RECT 102.020 118.900 102.770 119.090 ;
        RECT 102.940 119.075 103.950 119.245 ;
        RECT 101.510 118.355 102.740 118.525 ;
        RECT 99.980 118.115 100.910 118.285 ;
        RECT 99.980 118.080 100.155 118.115 ;
        RECT 99.160 117.885 99.440 118.055 ;
        RECT 99.160 117.715 99.435 117.885 ;
        RECT 99.625 117.715 100.155 118.080 ;
        RECT 100.580 117.545 100.910 117.945 ;
        RECT 101.080 117.715 101.335 118.285 ;
        RECT 101.785 117.750 102.030 118.355 ;
        RECT 102.250 117.545 102.760 118.080 ;
        RECT 102.940 117.715 103.130 119.075 ;
        RECT 103.300 118.735 103.575 118.875 ;
        RECT 103.300 118.565 103.580 118.735 ;
        RECT 103.300 117.715 103.575 118.565 ;
        RECT 103.780 118.275 103.950 119.075 ;
        RECT 104.120 118.285 104.290 119.415 ;
        RECT 104.460 118.785 104.630 119.755 ;
        RECT 104.800 118.955 104.970 120.095 ;
        RECT 105.140 118.955 105.475 119.925 ;
        RECT 105.690 118.955 105.920 120.095 ;
        RECT 104.460 118.455 104.655 118.785 ;
        RECT 104.880 118.455 105.135 118.785 ;
        RECT 104.880 118.285 105.050 118.455 ;
        RECT 105.305 118.285 105.475 118.955 ;
        RECT 106.090 118.945 106.420 119.925 ;
        RECT 106.590 118.955 106.800 120.095 ;
        RECT 107.120 119.165 107.290 119.925 ;
        RECT 107.470 119.335 107.800 120.095 ;
        RECT 107.120 118.995 107.785 119.165 ;
        RECT 107.970 119.020 108.240 119.925 ;
        RECT 105.670 118.535 106.000 118.785 ;
        RECT 104.120 118.115 105.050 118.285 ;
        RECT 104.120 118.080 104.295 118.115 ;
        RECT 103.765 117.715 104.295 118.080 ;
        RECT 104.720 117.545 105.050 117.945 ;
        RECT 105.220 117.715 105.475 118.285 ;
        RECT 105.690 117.545 105.920 118.365 ;
        RECT 106.170 118.345 106.420 118.945 ;
        RECT 107.615 118.850 107.785 118.995 ;
        RECT 107.050 118.445 107.380 118.815 ;
        RECT 107.615 118.520 107.900 118.850 ;
        RECT 106.090 117.715 106.420 118.345 ;
        RECT 106.590 117.545 106.800 118.365 ;
        RECT 107.615 118.265 107.785 118.520 ;
        RECT 107.120 118.095 107.785 118.265 ;
        RECT 108.070 118.220 108.240 119.020 ;
        RECT 108.410 119.005 111.000 120.095 ;
        RECT 111.170 119.005 112.380 120.095 ;
        RECT 108.410 118.485 109.620 119.005 ;
        RECT 109.790 118.315 111.000 118.835 ;
        RECT 111.170 118.465 111.690 119.005 ;
        RECT 107.120 117.715 107.290 118.095 ;
        RECT 107.470 117.545 107.800 117.925 ;
        RECT 107.980 117.715 108.240 118.220 ;
        RECT 108.410 117.545 111.000 118.315 ;
        RECT 111.860 118.295 112.380 118.835 ;
        RECT 111.170 117.545 112.380 118.295 ;
        RECT 18.165 117.375 112.465 117.545 ;
        RECT 18.250 116.625 19.460 117.375 ;
        RECT 18.250 116.085 18.770 116.625 ;
        RECT 20.610 116.555 20.820 117.375 ;
        RECT 20.990 116.575 21.320 117.205 ;
        RECT 18.940 115.915 19.460 116.455 ;
        RECT 20.990 115.975 21.240 116.575 ;
        RECT 21.490 116.555 21.720 117.375 ;
        RECT 21.930 116.650 22.220 117.375 ;
        RECT 22.480 116.825 22.650 117.115 ;
        RECT 22.820 116.995 23.150 117.375 ;
        RECT 22.480 116.655 23.145 116.825 ;
        RECT 21.410 116.135 21.740 116.385 ;
        RECT 18.250 114.825 19.460 115.915 ;
        RECT 20.610 114.825 20.820 115.965 ;
        RECT 20.990 114.995 21.320 115.975 ;
        RECT 21.490 114.825 21.720 115.965 ;
        RECT 21.930 114.825 22.220 115.990 ;
        RECT 22.395 115.835 22.745 116.485 ;
        RECT 22.915 115.665 23.145 116.655 ;
        RECT 22.480 115.495 23.145 115.665 ;
        RECT 22.480 114.995 22.650 115.495 ;
        RECT 22.820 114.825 23.150 115.325 ;
        RECT 23.320 114.995 23.545 117.115 ;
        RECT 23.760 116.995 24.090 117.375 ;
        RECT 24.260 116.825 24.430 117.155 ;
        RECT 24.730 116.995 25.745 117.195 ;
        RECT 23.735 116.635 24.430 116.825 ;
        RECT 23.735 115.665 23.905 116.635 ;
        RECT 24.075 115.835 24.485 116.455 ;
        RECT 24.655 115.885 24.875 116.755 ;
        RECT 25.055 116.445 25.405 116.815 ;
        RECT 25.575 116.265 25.745 116.995 ;
        RECT 25.915 116.935 26.325 117.375 ;
        RECT 26.615 116.735 26.865 117.165 ;
        RECT 27.065 116.915 27.385 117.375 ;
        RECT 27.945 116.985 28.795 117.155 ;
        RECT 25.915 116.395 26.325 116.725 ;
        RECT 26.615 116.395 27.035 116.735 ;
        RECT 25.325 116.225 25.745 116.265 ;
        RECT 25.325 116.055 26.675 116.225 ;
        RECT 23.735 115.495 24.430 115.665 ;
        RECT 24.655 115.505 25.155 115.885 ;
        RECT 23.760 114.825 24.090 115.325 ;
        RECT 24.260 114.995 24.430 115.495 ;
        RECT 25.325 115.210 25.495 116.055 ;
        RECT 26.425 115.895 26.675 116.055 ;
        RECT 25.665 115.625 25.915 115.885 ;
        RECT 26.845 115.625 27.035 116.395 ;
        RECT 25.665 115.375 27.035 115.625 ;
        RECT 27.205 116.565 28.455 116.735 ;
        RECT 27.205 115.805 27.375 116.565 ;
        RECT 28.125 116.445 28.455 116.565 ;
        RECT 27.545 115.985 27.725 116.395 ;
        RECT 28.625 116.225 28.795 116.985 ;
        RECT 28.995 116.895 29.655 117.375 ;
        RECT 29.835 116.780 30.155 117.110 ;
        RECT 28.985 116.455 29.645 116.725 ;
        RECT 28.985 116.395 29.315 116.455 ;
        RECT 29.465 116.225 29.795 116.285 ;
        RECT 27.895 116.055 29.795 116.225 ;
        RECT 27.205 115.495 27.725 115.805 ;
        RECT 27.895 115.545 28.065 116.055 ;
        RECT 29.965 115.885 30.155 116.780 ;
        RECT 28.235 115.715 30.155 115.885 ;
        RECT 29.835 115.695 30.155 115.715 ;
        RECT 30.355 116.465 30.605 117.115 ;
        RECT 30.785 116.915 31.070 117.375 ;
        RECT 31.250 116.665 31.505 117.195 ;
        RECT 30.355 116.135 31.155 116.465 ;
        RECT 27.895 115.375 29.105 115.545 ;
        RECT 24.665 115.040 25.495 115.210 ;
        RECT 25.735 114.825 26.115 115.205 ;
        RECT 26.295 115.085 26.465 115.375 ;
        RECT 27.895 115.295 28.065 115.375 ;
        RECT 26.635 114.825 26.965 115.205 ;
        RECT 27.435 115.045 28.065 115.295 ;
        RECT 28.245 114.825 28.665 115.205 ;
        RECT 28.865 115.085 29.105 115.375 ;
        RECT 29.335 114.825 29.665 115.515 ;
        RECT 29.835 115.085 30.005 115.695 ;
        RECT 30.355 115.545 30.605 116.135 ;
        RECT 31.325 115.805 31.505 116.665 ;
        RECT 32.550 116.555 32.780 117.375 ;
        RECT 32.950 116.575 33.280 117.205 ;
        RECT 32.530 116.135 32.860 116.385 ;
        RECT 33.030 115.975 33.280 116.575 ;
        RECT 33.450 116.555 33.660 117.375 ;
        RECT 33.895 116.635 34.150 117.205 ;
        RECT 34.320 116.975 34.650 117.375 ;
        RECT 35.075 116.840 35.605 117.205 ;
        RECT 35.075 116.805 35.250 116.840 ;
        RECT 34.320 116.635 35.250 116.805 ;
        RECT 30.275 115.035 30.605 115.545 ;
        RECT 30.785 114.825 31.070 115.625 ;
        RECT 31.250 115.335 31.505 115.805 ;
        RECT 31.250 115.165 31.590 115.335 ;
        RECT 31.250 115.135 31.505 115.165 ;
        RECT 32.550 114.825 32.780 115.965 ;
        RECT 32.950 114.995 33.280 115.975 ;
        RECT 33.895 115.965 34.065 116.635 ;
        RECT 34.320 116.465 34.490 116.635 ;
        RECT 34.235 116.135 34.490 116.465 ;
        RECT 34.715 116.135 34.910 116.465 ;
        RECT 33.450 114.825 33.660 115.965 ;
        RECT 33.895 114.995 34.230 115.965 ;
        RECT 34.400 114.825 34.570 115.965 ;
        RECT 34.740 115.165 34.910 116.135 ;
        RECT 35.080 115.505 35.250 116.635 ;
        RECT 35.420 115.845 35.590 116.645 ;
        RECT 35.795 116.355 36.070 117.205 ;
        RECT 35.790 116.185 36.070 116.355 ;
        RECT 35.795 116.045 36.070 116.185 ;
        RECT 36.240 115.845 36.430 117.205 ;
        RECT 36.610 116.840 37.120 117.375 ;
        RECT 37.340 116.565 37.585 117.170 ;
        RECT 38.405 117.035 38.660 117.195 ;
        RECT 38.320 116.865 38.660 117.035 ;
        RECT 38.840 116.915 39.125 117.375 ;
        RECT 38.405 116.665 38.660 116.865 ;
        RECT 36.630 116.395 37.860 116.565 ;
        RECT 35.420 115.675 36.430 115.845 ;
        RECT 36.600 115.830 37.350 116.020 ;
        RECT 35.080 115.335 36.205 115.505 ;
        RECT 36.600 115.165 36.770 115.830 ;
        RECT 37.520 115.585 37.860 116.395 ;
        RECT 34.740 114.995 36.770 115.165 ;
        RECT 36.940 114.825 37.110 115.585 ;
        RECT 37.345 115.175 37.860 115.585 ;
        RECT 38.405 115.805 38.585 116.665 ;
        RECT 39.305 116.465 39.555 117.115 ;
        RECT 38.755 116.135 39.555 116.465 ;
        RECT 38.405 115.135 38.660 115.805 ;
        RECT 38.840 114.825 39.125 115.625 ;
        RECT 39.305 115.545 39.555 116.135 ;
        RECT 39.755 116.780 40.075 117.110 ;
        RECT 40.255 116.895 40.915 117.375 ;
        RECT 41.115 116.985 41.965 117.155 ;
        RECT 39.755 115.885 39.945 116.780 ;
        RECT 40.265 116.455 40.925 116.725 ;
        RECT 40.595 116.395 40.925 116.455 ;
        RECT 40.115 116.225 40.445 116.285 ;
        RECT 41.115 116.225 41.285 116.985 ;
        RECT 42.525 116.915 42.845 117.375 ;
        RECT 43.045 116.735 43.295 117.165 ;
        RECT 43.585 116.935 43.995 117.375 ;
        RECT 44.165 116.995 45.180 117.195 ;
        RECT 41.455 116.565 42.705 116.735 ;
        RECT 41.455 116.445 41.785 116.565 ;
        RECT 40.115 116.055 42.015 116.225 ;
        RECT 39.755 115.715 41.675 115.885 ;
        RECT 39.755 115.695 40.075 115.715 ;
        RECT 39.305 115.035 39.635 115.545 ;
        RECT 39.905 115.085 40.075 115.695 ;
        RECT 41.845 115.545 42.015 116.055 ;
        RECT 42.185 115.985 42.365 116.395 ;
        RECT 42.535 115.805 42.705 116.565 ;
        RECT 40.245 114.825 40.575 115.515 ;
        RECT 40.805 115.375 42.015 115.545 ;
        RECT 42.185 115.495 42.705 115.805 ;
        RECT 42.875 116.395 43.295 116.735 ;
        RECT 43.585 116.395 43.995 116.725 ;
        RECT 42.875 115.625 43.065 116.395 ;
        RECT 44.165 116.265 44.335 116.995 ;
        RECT 45.480 116.825 45.650 117.155 ;
        RECT 45.820 116.995 46.150 117.375 ;
        RECT 44.505 116.445 44.855 116.815 ;
        RECT 44.165 116.225 44.585 116.265 ;
        RECT 43.235 116.055 44.585 116.225 ;
        RECT 43.235 115.895 43.485 116.055 ;
        RECT 43.995 115.625 44.245 115.885 ;
        RECT 42.875 115.375 44.245 115.625 ;
        RECT 40.805 115.085 41.045 115.375 ;
        RECT 41.845 115.295 42.015 115.375 ;
        RECT 41.245 114.825 41.665 115.205 ;
        RECT 41.845 115.045 42.475 115.295 ;
        RECT 42.945 114.825 43.275 115.205 ;
        RECT 43.445 115.085 43.615 115.375 ;
        RECT 44.415 115.210 44.585 116.055 ;
        RECT 45.035 115.885 45.255 116.755 ;
        RECT 45.480 116.635 46.175 116.825 ;
        RECT 44.755 115.505 45.255 115.885 ;
        RECT 45.425 115.835 45.835 116.455 ;
        RECT 46.005 115.665 46.175 116.635 ;
        RECT 45.480 115.495 46.175 115.665 ;
        RECT 43.795 114.825 44.175 115.205 ;
        RECT 44.415 115.040 45.245 115.210 ;
        RECT 45.480 114.995 45.650 115.495 ;
        RECT 45.820 114.825 46.150 115.325 ;
        RECT 46.365 114.995 46.590 117.115 ;
        RECT 46.760 116.995 47.090 117.375 ;
        RECT 47.260 116.825 47.430 117.115 ;
        RECT 46.765 116.655 47.430 116.825 ;
        RECT 46.765 115.665 46.995 116.655 ;
        RECT 47.690 116.650 47.980 117.375 ;
        RECT 48.525 117.035 48.780 117.195 ;
        RECT 48.440 116.865 48.780 117.035 ;
        RECT 48.960 116.915 49.245 117.375 ;
        RECT 48.525 116.665 48.780 116.865 ;
        RECT 47.165 115.835 47.515 116.485 ;
        RECT 46.765 115.495 47.430 115.665 ;
        RECT 46.760 114.825 47.090 115.325 ;
        RECT 47.260 114.995 47.430 115.495 ;
        RECT 47.690 114.825 47.980 115.990 ;
        RECT 48.525 115.805 48.705 116.665 ;
        RECT 49.425 116.465 49.675 117.115 ;
        RECT 48.875 116.135 49.675 116.465 ;
        RECT 48.525 115.135 48.780 115.805 ;
        RECT 48.960 114.825 49.245 115.625 ;
        RECT 49.425 115.545 49.675 116.135 ;
        RECT 49.875 116.780 50.195 117.110 ;
        RECT 50.375 116.895 51.035 117.375 ;
        RECT 51.235 116.985 52.085 117.155 ;
        RECT 49.875 115.885 50.065 116.780 ;
        RECT 50.385 116.455 51.045 116.725 ;
        RECT 50.715 116.395 51.045 116.455 ;
        RECT 50.235 116.225 50.565 116.285 ;
        RECT 51.235 116.225 51.405 116.985 ;
        RECT 52.645 116.915 52.965 117.375 ;
        RECT 53.165 116.735 53.415 117.165 ;
        RECT 53.705 116.935 54.115 117.375 ;
        RECT 54.285 116.995 55.300 117.195 ;
        RECT 51.575 116.565 52.825 116.735 ;
        RECT 51.575 116.445 51.905 116.565 ;
        RECT 50.235 116.055 52.135 116.225 ;
        RECT 49.875 115.715 51.795 115.885 ;
        RECT 49.875 115.695 50.195 115.715 ;
        RECT 49.425 115.035 49.755 115.545 ;
        RECT 50.025 115.085 50.195 115.695 ;
        RECT 51.965 115.545 52.135 116.055 ;
        RECT 52.305 115.985 52.485 116.395 ;
        RECT 52.655 115.805 52.825 116.565 ;
        RECT 50.365 114.825 50.695 115.515 ;
        RECT 50.925 115.375 52.135 115.545 ;
        RECT 52.305 115.495 52.825 115.805 ;
        RECT 52.995 116.395 53.415 116.735 ;
        RECT 53.705 116.395 54.115 116.725 ;
        RECT 52.995 115.625 53.185 116.395 ;
        RECT 54.285 116.265 54.455 116.995 ;
        RECT 55.600 116.825 55.770 117.155 ;
        RECT 55.940 116.995 56.270 117.375 ;
        RECT 54.625 116.445 54.975 116.815 ;
        RECT 54.285 116.225 54.705 116.265 ;
        RECT 53.355 116.055 54.705 116.225 ;
        RECT 53.355 115.895 53.605 116.055 ;
        RECT 54.115 115.625 54.365 115.885 ;
        RECT 52.995 115.375 54.365 115.625 ;
        RECT 50.925 115.085 51.165 115.375 ;
        RECT 51.965 115.295 52.135 115.375 ;
        RECT 51.365 114.825 51.785 115.205 ;
        RECT 51.965 115.045 52.595 115.295 ;
        RECT 53.065 114.825 53.395 115.205 ;
        RECT 53.565 115.085 53.735 115.375 ;
        RECT 54.535 115.210 54.705 116.055 ;
        RECT 55.155 115.885 55.375 116.755 ;
        RECT 55.600 116.635 56.295 116.825 ;
        RECT 54.875 115.505 55.375 115.885 ;
        RECT 55.545 115.835 55.955 116.455 ;
        RECT 56.125 115.665 56.295 116.635 ;
        RECT 55.600 115.495 56.295 115.665 ;
        RECT 53.915 114.825 54.295 115.205 ;
        RECT 54.535 115.040 55.365 115.210 ;
        RECT 55.600 114.995 55.770 115.495 ;
        RECT 55.940 114.825 56.270 115.325 ;
        RECT 56.485 114.995 56.710 117.115 ;
        RECT 56.880 116.995 57.210 117.375 ;
        RECT 57.380 116.825 57.550 117.115 ;
        RECT 56.885 116.655 57.550 116.825 ;
        RECT 57.900 116.825 58.070 117.115 ;
        RECT 58.240 116.995 58.570 117.375 ;
        RECT 57.900 116.655 58.565 116.825 ;
        RECT 56.885 115.665 57.115 116.655 ;
        RECT 57.285 115.835 57.635 116.485 ;
        RECT 57.815 115.835 58.165 116.485 ;
        RECT 58.335 115.665 58.565 116.655 ;
        RECT 56.885 115.495 57.550 115.665 ;
        RECT 56.880 114.825 57.210 115.325 ;
        RECT 57.380 114.995 57.550 115.495 ;
        RECT 57.900 115.495 58.565 115.665 ;
        RECT 57.900 114.995 58.070 115.495 ;
        RECT 58.240 114.825 58.570 115.325 ;
        RECT 58.740 114.995 58.965 117.115 ;
        RECT 59.180 116.995 59.510 117.375 ;
        RECT 59.680 116.825 59.850 117.155 ;
        RECT 60.150 116.995 61.165 117.195 ;
        RECT 59.155 116.635 59.850 116.825 ;
        RECT 59.155 115.665 59.325 116.635 ;
        RECT 59.495 115.835 59.905 116.455 ;
        RECT 60.075 115.885 60.295 116.755 ;
        RECT 60.475 116.445 60.825 116.815 ;
        RECT 60.995 116.265 61.165 116.995 ;
        RECT 61.335 116.935 61.745 117.375 ;
        RECT 62.035 116.735 62.285 117.165 ;
        RECT 62.485 116.915 62.805 117.375 ;
        RECT 63.365 116.985 64.215 117.155 ;
        RECT 61.335 116.395 61.745 116.725 ;
        RECT 62.035 116.395 62.455 116.735 ;
        RECT 60.745 116.225 61.165 116.265 ;
        RECT 60.745 116.055 62.095 116.225 ;
        RECT 59.155 115.495 59.850 115.665 ;
        RECT 60.075 115.505 60.575 115.885 ;
        RECT 59.180 114.825 59.510 115.325 ;
        RECT 59.680 114.995 59.850 115.495 ;
        RECT 60.745 115.210 60.915 116.055 ;
        RECT 61.845 115.895 62.095 116.055 ;
        RECT 61.085 115.625 61.335 115.885 ;
        RECT 62.265 115.625 62.455 116.395 ;
        RECT 61.085 115.375 62.455 115.625 ;
        RECT 62.625 116.565 63.875 116.735 ;
        RECT 62.625 115.805 62.795 116.565 ;
        RECT 63.545 116.445 63.875 116.565 ;
        RECT 62.965 115.985 63.145 116.395 ;
        RECT 64.045 116.225 64.215 116.985 ;
        RECT 64.415 116.895 65.075 117.375 ;
        RECT 65.255 116.780 65.575 117.110 ;
        RECT 64.405 116.455 65.065 116.725 ;
        RECT 64.405 116.395 64.735 116.455 ;
        RECT 64.885 116.225 65.215 116.285 ;
        RECT 63.315 116.055 65.215 116.225 ;
        RECT 62.625 115.495 63.145 115.805 ;
        RECT 63.315 115.545 63.485 116.055 ;
        RECT 65.385 115.885 65.575 116.780 ;
        RECT 63.655 115.715 65.575 115.885 ;
        RECT 65.255 115.695 65.575 115.715 ;
        RECT 65.775 116.465 66.025 117.115 ;
        RECT 66.205 116.915 66.490 117.375 ;
        RECT 66.670 117.035 66.925 117.195 ;
        RECT 66.670 116.865 67.010 117.035 ;
        RECT 66.670 116.665 66.925 116.865 ;
        RECT 65.775 116.135 66.575 116.465 ;
        RECT 63.315 115.375 64.525 115.545 ;
        RECT 60.085 115.040 60.915 115.210 ;
        RECT 61.155 114.825 61.535 115.205 ;
        RECT 61.715 115.085 61.885 115.375 ;
        RECT 63.315 115.295 63.485 115.375 ;
        RECT 62.055 114.825 62.385 115.205 ;
        RECT 62.855 115.045 63.485 115.295 ;
        RECT 63.665 114.825 64.085 115.205 ;
        RECT 64.285 115.085 64.525 115.375 ;
        RECT 64.755 114.825 65.085 115.515 ;
        RECT 65.255 115.085 65.425 115.695 ;
        RECT 65.775 115.545 66.025 116.135 ;
        RECT 66.745 115.805 66.925 116.665 ;
        RECT 65.695 115.035 66.025 115.545 ;
        RECT 66.205 114.825 66.490 115.625 ;
        RECT 66.670 115.135 66.925 115.805 ;
        RECT 67.470 116.700 67.730 117.205 ;
        RECT 67.910 116.995 68.240 117.375 ;
        RECT 68.420 116.825 68.590 117.205 ;
        RECT 67.470 115.900 67.640 116.700 ;
        RECT 67.925 116.655 68.590 116.825 ;
        RECT 69.400 116.825 69.570 117.205 ;
        RECT 69.750 116.995 70.080 117.375 ;
        RECT 69.400 116.655 70.065 116.825 ;
        RECT 70.260 116.700 70.520 117.205 ;
        RECT 67.925 116.400 68.095 116.655 ;
        RECT 67.810 116.070 68.095 116.400 ;
        RECT 68.330 116.105 68.660 116.475 ;
        RECT 69.330 116.105 69.660 116.475 ;
        RECT 69.895 116.400 70.065 116.655 ;
        RECT 67.925 115.925 68.095 116.070 ;
        RECT 69.895 116.070 70.180 116.400 ;
        RECT 69.895 115.925 70.065 116.070 ;
        RECT 67.470 114.995 67.740 115.900 ;
        RECT 67.925 115.755 68.590 115.925 ;
        RECT 67.910 114.825 68.240 115.585 ;
        RECT 68.420 114.995 68.590 115.755 ;
        RECT 69.400 115.755 70.065 115.925 ;
        RECT 70.350 115.900 70.520 116.700 ;
        RECT 70.730 116.555 70.960 117.375 ;
        RECT 71.130 116.575 71.460 117.205 ;
        RECT 70.710 116.135 71.040 116.385 ;
        RECT 71.210 115.975 71.460 116.575 ;
        RECT 71.630 116.555 71.840 117.375 ;
        RECT 72.110 116.555 72.340 117.375 ;
        RECT 72.510 116.575 72.840 117.205 ;
        RECT 72.090 116.135 72.420 116.385 ;
        RECT 72.590 115.975 72.840 116.575 ;
        RECT 73.010 116.555 73.220 117.375 ;
        RECT 73.450 116.650 73.740 117.375 ;
        RECT 73.915 116.635 74.170 117.205 ;
        RECT 74.340 116.975 74.670 117.375 ;
        RECT 75.095 116.840 75.625 117.205 ;
        RECT 75.095 116.805 75.270 116.840 ;
        RECT 74.340 116.635 75.270 116.805 ;
        RECT 69.400 114.995 69.570 115.755 ;
        RECT 69.750 114.825 70.080 115.585 ;
        RECT 70.250 114.995 70.520 115.900 ;
        RECT 70.730 114.825 70.960 115.965 ;
        RECT 71.130 114.995 71.460 115.975 ;
        RECT 71.630 114.825 71.840 115.965 ;
        RECT 72.110 114.825 72.340 115.965 ;
        RECT 72.510 114.995 72.840 115.975 ;
        RECT 73.010 114.825 73.220 115.965 ;
        RECT 73.450 114.825 73.740 115.990 ;
        RECT 73.915 115.965 74.085 116.635 ;
        RECT 74.340 116.465 74.510 116.635 ;
        RECT 74.255 116.135 74.510 116.465 ;
        RECT 74.735 116.135 74.930 116.465 ;
        RECT 73.915 114.995 74.250 115.965 ;
        RECT 74.420 114.825 74.590 115.965 ;
        RECT 74.760 115.165 74.930 116.135 ;
        RECT 75.100 115.505 75.270 116.635 ;
        RECT 75.440 115.845 75.610 116.645 ;
        RECT 75.815 116.355 76.090 117.205 ;
        RECT 75.810 116.185 76.090 116.355 ;
        RECT 75.815 116.045 76.090 116.185 ;
        RECT 76.260 115.845 76.450 117.205 ;
        RECT 76.630 116.840 77.140 117.375 ;
        RECT 77.360 116.565 77.605 117.170 ;
        RECT 78.885 116.695 79.140 117.195 ;
        RECT 79.320 116.915 79.605 117.375 ;
        RECT 78.800 116.665 79.140 116.695 ;
        RECT 76.650 116.395 77.880 116.565 ;
        RECT 78.800 116.525 79.065 116.665 ;
        RECT 75.440 115.675 76.450 115.845 ;
        RECT 76.620 115.830 77.370 116.020 ;
        RECT 75.100 115.335 76.225 115.505 ;
        RECT 76.620 115.165 76.790 115.830 ;
        RECT 77.540 115.585 77.880 116.395 ;
        RECT 74.760 114.995 76.790 115.165 ;
        RECT 76.960 114.825 77.130 115.585 ;
        RECT 77.365 115.175 77.880 115.585 ;
        RECT 78.885 115.805 79.065 116.525 ;
        RECT 79.785 116.465 80.035 117.115 ;
        RECT 79.235 116.135 80.035 116.465 ;
        RECT 78.885 115.135 79.140 115.805 ;
        RECT 79.320 114.825 79.605 115.625 ;
        RECT 79.785 115.545 80.035 116.135 ;
        RECT 80.235 116.780 80.555 117.110 ;
        RECT 80.735 116.895 81.395 117.375 ;
        RECT 81.595 116.985 82.445 117.155 ;
        RECT 80.235 115.885 80.425 116.780 ;
        RECT 80.745 116.455 81.405 116.725 ;
        RECT 81.075 116.395 81.405 116.455 ;
        RECT 80.595 116.225 80.925 116.285 ;
        RECT 81.595 116.225 81.765 116.985 ;
        RECT 83.005 116.915 83.325 117.375 ;
        RECT 83.525 116.735 83.775 117.165 ;
        RECT 84.065 116.935 84.475 117.375 ;
        RECT 84.645 116.995 85.660 117.195 ;
        RECT 81.935 116.565 83.185 116.735 ;
        RECT 81.935 116.445 82.265 116.565 ;
        RECT 80.595 116.055 82.495 116.225 ;
        RECT 80.235 115.715 82.155 115.885 ;
        RECT 80.235 115.695 80.555 115.715 ;
        RECT 79.785 115.035 80.115 115.545 ;
        RECT 80.385 115.085 80.555 115.695 ;
        RECT 82.325 115.545 82.495 116.055 ;
        RECT 82.665 115.985 82.845 116.395 ;
        RECT 83.015 115.805 83.185 116.565 ;
        RECT 80.725 114.825 81.055 115.515 ;
        RECT 81.285 115.375 82.495 115.545 ;
        RECT 82.665 115.495 83.185 115.805 ;
        RECT 83.355 116.395 83.775 116.735 ;
        RECT 84.065 116.395 84.475 116.725 ;
        RECT 83.355 115.625 83.545 116.395 ;
        RECT 84.645 116.265 84.815 116.995 ;
        RECT 85.960 116.825 86.130 117.155 ;
        RECT 86.300 116.995 86.630 117.375 ;
        RECT 84.985 116.445 85.335 116.815 ;
        RECT 84.645 116.225 85.065 116.265 ;
        RECT 83.715 116.055 85.065 116.225 ;
        RECT 83.715 115.895 83.965 116.055 ;
        RECT 84.475 115.625 84.725 115.885 ;
        RECT 83.355 115.375 84.725 115.625 ;
        RECT 81.285 115.085 81.525 115.375 ;
        RECT 82.325 115.295 82.495 115.375 ;
        RECT 81.725 114.825 82.145 115.205 ;
        RECT 82.325 115.045 82.955 115.295 ;
        RECT 83.425 114.825 83.755 115.205 ;
        RECT 83.925 115.085 84.095 115.375 ;
        RECT 84.895 115.210 85.065 116.055 ;
        RECT 85.515 115.885 85.735 116.755 ;
        RECT 85.960 116.635 86.655 116.825 ;
        RECT 85.235 115.505 85.735 115.885 ;
        RECT 85.905 115.835 86.315 116.455 ;
        RECT 86.485 115.665 86.655 116.635 ;
        RECT 85.960 115.495 86.655 115.665 ;
        RECT 84.275 114.825 84.655 115.205 ;
        RECT 84.895 115.040 85.725 115.210 ;
        RECT 85.960 114.995 86.130 115.495 ;
        RECT 86.300 114.825 86.630 115.325 ;
        RECT 86.845 114.995 87.070 117.115 ;
        RECT 87.240 116.995 87.570 117.375 ;
        RECT 87.740 116.825 87.910 117.115 ;
        RECT 87.245 116.655 87.910 116.825 ;
        RECT 88.170 116.700 88.430 117.205 ;
        RECT 88.610 116.995 88.940 117.375 ;
        RECT 89.120 116.825 89.290 117.205 ;
        RECT 87.245 115.665 87.475 116.655 ;
        RECT 87.645 115.835 87.995 116.485 ;
        RECT 88.170 115.900 88.340 116.700 ;
        RECT 88.625 116.655 89.290 116.825 ;
        RECT 89.925 116.665 90.180 117.195 ;
        RECT 90.360 116.915 90.645 117.375 ;
        RECT 88.625 116.400 88.795 116.655 ;
        RECT 88.510 116.070 88.795 116.400 ;
        RECT 89.030 116.105 89.360 116.475 ;
        RECT 88.625 115.925 88.795 116.070 ;
        RECT 87.245 115.495 87.910 115.665 ;
        RECT 87.240 114.825 87.570 115.325 ;
        RECT 87.740 114.995 87.910 115.495 ;
        RECT 88.170 114.995 88.440 115.900 ;
        RECT 88.625 115.755 89.290 115.925 ;
        RECT 88.610 114.825 88.940 115.585 ;
        RECT 89.120 114.995 89.290 115.755 ;
        RECT 89.925 115.805 90.105 116.665 ;
        RECT 90.825 116.465 91.075 117.115 ;
        RECT 90.275 116.135 91.075 116.465 ;
        RECT 89.925 115.335 90.180 115.805 ;
        RECT 89.840 115.165 90.180 115.335 ;
        RECT 89.925 115.135 90.180 115.165 ;
        RECT 90.360 114.825 90.645 115.625 ;
        RECT 90.825 115.545 91.075 116.135 ;
        RECT 91.275 116.780 91.595 117.110 ;
        RECT 91.775 116.895 92.435 117.375 ;
        RECT 92.635 116.985 93.485 117.155 ;
        RECT 91.275 115.885 91.465 116.780 ;
        RECT 91.785 116.455 92.445 116.725 ;
        RECT 92.115 116.395 92.445 116.455 ;
        RECT 91.635 116.225 91.965 116.285 ;
        RECT 92.635 116.225 92.805 116.985 ;
        RECT 94.045 116.915 94.365 117.375 ;
        RECT 94.565 116.735 94.815 117.165 ;
        RECT 95.105 116.935 95.515 117.375 ;
        RECT 95.685 116.995 96.700 117.195 ;
        RECT 92.975 116.565 94.225 116.735 ;
        RECT 92.975 116.445 93.305 116.565 ;
        RECT 91.635 116.055 93.535 116.225 ;
        RECT 91.275 115.715 93.195 115.885 ;
        RECT 91.275 115.695 91.595 115.715 ;
        RECT 90.825 115.035 91.155 115.545 ;
        RECT 91.425 115.085 91.595 115.695 ;
        RECT 93.365 115.545 93.535 116.055 ;
        RECT 93.705 115.985 93.885 116.395 ;
        RECT 94.055 115.805 94.225 116.565 ;
        RECT 91.765 114.825 92.095 115.515 ;
        RECT 92.325 115.375 93.535 115.545 ;
        RECT 93.705 115.495 94.225 115.805 ;
        RECT 94.395 116.395 94.815 116.735 ;
        RECT 95.105 116.395 95.515 116.725 ;
        RECT 94.395 115.625 94.585 116.395 ;
        RECT 95.685 116.265 95.855 116.995 ;
        RECT 97.000 116.825 97.170 117.155 ;
        RECT 97.340 116.995 97.670 117.375 ;
        RECT 96.025 116.445 96.375 116.815 ;
        RECT 95.685 116.225 96.105 116.265 ;
        RECT 94.755 116.055 96.105 116.225 ;
        RECT 94.755 115.895 95.005 116.055 ;
        RECT 95.515 115.625 95.765 115.885 ;
        RECT 94.395 115.375 95.765 115.625 ;
        RECT 92.325 115.085 92.565 115.375 ;
        RECT 93.365 115.295 93.535 115.375 ;
        RECT 92.765 114.825 93.185 115.205 ;
        RECT 93.365 115.045 93.995 115.295 ;
        RECT 94.465 114.825 94.795 115.205 ;
        RECT 94.965 115.085 95.135 115.375 ;
        RECT 95.935 115.210 96.105 116.055 ;
        RECT 96.555 115.885 96.775 116.755 ;
        RECT 97.000 116.635 97.695 116.825 ;
        RECT 96.275 115.505 96.775 115.885 ;
        RECT 96.945 115.835 97.355 116.455 ;
        RECT 97.525 115.665 97.695 116.635 ;
        RECT 97.000 115.495 97.695 115.665 ;
        RECT 95.315 114.825 95.695 115.205 ;
        RECT 95.935 115.040 96.765 115.210 ;
        RECT 97.000 114.995 97.170 115.495 ;
        RECT 97.340 114.825 97.670 115.325 ;
        RECT 97.885 114.995 98.110 117.115 ;
        RECT 98.280 116.995 98.610 117.375 ;
        RECT 98.780 116.825 98.950 117.115 ;
        RECT 98.285 116.655 98.950 116.825 ;
        RECT 98.285 115.665 98.515 116.655 ;
        RECT 99.210 116.650 99.500 117.375 ;
        RECT 100.130 116.700 100.390 117.205 ;
        RECT 100.570 116.995 100.900 117.375 ;
        RECT 101.080 116.825 101.250 117.205 ;
        RECT 101.885 117.035 102.140 117.195 ;
        RECT 101.800 116.865 102.140 117.035 ;
        RECT 102.320 116.915 102.605 117.375 ;
        RECT 98.685 115.835 99.035 116.485 ;
        RECT 98.285 115.495 98.950 115.665 ;
        RECT 98.280 114.825 98.610 115.325 ;
        RECT 98.780 114.995 98.950 115.495 ;
        RECT 99.210 114.825 99.500 115.990 ;
        RECT 100.130 115.900 100.300 116.700 ;
        RECT 100.585 116.655 101.250 116.825 ;
        RECT 101.885 116.665 102.140 116.865 ;
        RECT 100.585 116.400 100.755 116.655 ;
        RECT 100.470 116.070 100.755 116.400 ;
        RECT 100.990 116.105 101.320 116.475 ;
        RECT 100.585 115.925 100.755 116.070 ;
        RECT 100.130 114.995 100.400 115.900 ;
        RECT 100.585 115.755 101.250 115.925 ;
        RECT 100.570 114.825 100.900 115.585 ;
        RECT 101.080 114.995 101.250 115.755 ;
        RECT 101.885 115.805 102.065 116.665 ;
        RECT 102.785 116.465 103.035 117.115 ;
        RECT 102.235 116.135 103.035 116.465 ;
        RECT 101.885 115.135 102.140 115.805 ;
        RECT 102.320 114.825 102.605 115.625 ;
        RECT 102.785 115.545 103.035 116.135 ;
        RECT 103.235 116.780 103.555 117.110 ;
        RECT 103.735 116.895 104.395 117.375 ;
        RECT 104.595 116.985 105.445 117.155 ;
        RECT 103.235 115.885 103.425 116.780 ;
        RECT 103.745 116.455 104.405 116.725 ;
        RECT 104.075 116.395 104.405 116.455 ;
        RECT 103.595 116.225 103.925 116.285 ;
        RECT 104.595 116.225 104.765 116.985 ;
        RECT 106.005 116.915 106.325 117.375 ;
        RECT 106.525 116.735 106.775 117.165 ;
        RECT 107.065 116.935 107.475 117.375 ;
        RECT 107.645 116.995 108.660 117.195 ;
        RECT 104.935 116.565 106.185 116.735 ;
        RECT 104.935 116.445 105.265 116.565 ;
        RECT 103.595 116.055 105.495 116.225 ;
        RECT 103.235 115.715 105.155 115.885 ;
        RECT 103.235 115.695 103.555 115.715 ;
        RECT 102.785 115.035 103.115 115.545 ;
        RECT 103.385 115.085 103.555 115.695 ;
        RECT 105.325 115.545 105.495 116.055 ;
        RECT 105.665 115.985 105.845 116.395 ;
        RECT 106.015 115.805 106.185 116.565 ;
        RECT 103.725 114.825 104.055 115.515 ;
        RECT 104.285 115.375 105.495 115.545 ;
        RECT 105.665 115.495 106.185 115.805 ;
        RECT 106.355 116.395 106.775 116.735 ;
        RECT 107.065 116.395 107.475 116.725 ;
        RECT 106.355 115.625 106.545 116.395 ;
        RECT 107.645 116.265 107.815 116.995 ;
        RECT 108.960 116.825 109.130 117.155 ;
        RECT 109.300 116.995 109.630 117.375 ;
        RECT 107.985 116.445 108.335 116.815 ;
        RECT 107.645 116.225 108.065 116.265 ;
        RECT 106.715 116.055 108.065 116.225 ;
        RECT 106.715 115.895 106.965 116.055 ;
        RECT 107.475 115.625 107.725 115.885 ;
        RECT 106.355 115.375 107.725 115.625 ;
        RECT 104.285 115.085 104.525 115.375 ;
        RECT 105.325 115.295 105.495 115.375 ;
        RECT 104.725 114.825 105.145 115.205 ;
        RECT 105.325 115.045 105.955 115.295 ;
        RECT 106.425 114.825 106.755 115.205 ;
        RECT 106.925 115.085 107.095 115.375 ;
        RECT 107.895 115.210 108.065 116.055 ;
        RECT 108.515 115.885 108.735 116.755 ;
        RECT 108.960 116.635 109.655 116.825 ;
        RECT 108.235 115.505 108.735 115.885 ;
        RECT 108.905 115.835 109.315 116.455 ;
        RECT 109.485 115.665 109.655 116.635 ;
        RECT 108.960 115.495 109.655 115.665 ;
        RECT 107.275 114.825 107.655 115.205 ;
        RECT 107.895 115.040 108.725 115.210 ;
        RECT 108.960 114.995 109.130 115.495 ;
        RECT 109.300 114.825 109.630 115.325 ;
        RECT 109.845 114.995 110.070 117.115 ;
        RECT 110.240 116.995 110.570 117.375 ;
        RECT 110.740 116.825 110.910 117.115 ;
        RECT 110.245 116.655 110.910 116.825 ;
        RECT 110.245 115.665 110.475 116.655 ;
        RECT 111.170 116.625 112.380 117.375 ;
        RECT 110.645 115.835 110.995 116.485 ;
        RECT 111.170 115.915 111.690 116.455 ;
        RECT 111.860 116.085 112.380 116.625 ;
        RECT 110.245 115.495 110.910 115.665 ;
        RECT 110.240 114.825 110.570 115.325 ;
        RECT 110.740 114.995 110.910 115.495 ;
        RECT 111.170 114.825 112.380 115.915 ;
        RECT 18.165 114.655 112.465 114.825 ;
        RECT 18.250 113.565 19.460 114.655 ;
        RECT 18.250 112.855 18.770 113.395 ;
        RECT 18.940 113.025 19.460 113.565 ;
        RECT 19.720 113.725 19.890 114.485 ;
        RECT 20.070 113.895 20.400 114.655 ;
        RECT 19.720 113.555 20.385 113.725 ;
        RECT 20.570 113.580 20.840 114.485 ;
        RECT 20.215 113.410 20.385 113.555 ;
        RECT 19.650 113.005 19.980 113.375 ;
        RECT 20.215 113.080 20.500 113.410 ;
        RECT 18.250 112.105 19.460 112.855 ;
        RECT 20.215 112.825 20.385 113.080 ;
        RECT 19.720 112.655 20.385 112.825 ;
        RECT 20.670 112.780 20.840 113.580 ;
        RECT 21.070 113.515 21.280 114.655 ;
        RECT 21.450 113.505 21.780 114.485 ;
        RECT 21.950 113.515 22.180 114.655 ;
        RECT 22.765 113.675 23.020 114.345 ;
        RECT 23.200 113.855 23.485 114.655 ;
        RECT 23.665 113.935 23.995 114.445 ;
        RECT 19.720 112.275 19.890 112.655 ;
        RECT 20.070 112.105 20.400 112.485 ;
        RECT 20.580 112.275 20.840 112.780 ;
        RECT 21.070 112.105 21.280 112.925 ;
        RECT 21.450 112.905 21.700 113.505 ;
        RECT 21.870 113.095 22.200 113.345 ;
        RECT 22.765 113.295 22.945 113.675 ;
        RECT 23.665 113.345 23.915 113.935 ;
        RECT 24.265 113.785 24.435 114.395 ;
        RECT 24.605 113.965 24.935 114.655 ;
        RECT 25.165 114.105 25.405 114.395 ;
        RECT 25.605 114.275 26.025 114.655 ;
        RECT 26.205 114.185 26.835 114.435 ;
        RECT 27.305 114.275 27.635 114.655 ;
        RECT 26.205 114.105 26.375 114.185 ;
        RECT 27.805 114.105 27.975 114.395 ;
        RECT 28.155 114.275 28.535 114.655 ;
        RECT 28.775 114.270 29.605 114.440 ;
        RECT 25.165 113.935 26.375 114.105 ;
        RECT 22.680 113.125 22.945 113.295 ;
        RECT 21.450 112.275 21.780 112.905 ;
        RECT 21.950 112.105 22.180 112.925 ;
        RECT 22.765 112.815 22.945 113.125 ;
        RECT 23.115 113.015 23.915 113.345 ;
        RECT 22.765 112.285 23.020 112.815 ;
        RECT 23.200 112.105 23.485 112.565 ;
        RECT 23.665 112.365 23.915 113.015 ;
        RECT 24.115 113.765 24.435 113.785 ;
        RECT 24.115 113.595 26.035 113.765 ;
        RECT 24.115 112.700 24.305 113.595 ;
        RECT 26.205 113.425 26.375 113.935 ;
        RECT 26.545 113.675 27.065 113.985 ;
        RECT 24.475 113.255 26.375 113.425 ;
        RECT 24.475 113.195 24.805 113.255 ;
        RECT 24.955 113.025 25.285 113.085 ;
        RECT 24.625 112.755 25.285 113.025 ;
        RECT 24.115 112.370 24.435 112.700 ;
        RECT 24.615 112.105 25.275 112.585 ;
        RECT 25.475 112.495 25.645 113.255 ;
        RECT 26.545 113.085 26.725 113.495 ;
        RECT 25.815 112.915 26.145 113.035 ;
        RECT 26.895 112.915 27.065 113.675 ;
        RECT 25.815 112.745 27.065 112.915 ;
        RECT 27.235 113.855 28.605 114.105 ;
        RECT 27.235 113.085 27.425 113.855 ;
        RECT 28.355 113.595 28.605 113.855 ;
        RECT 27.595 113.425 27.845 113.585 ;
        RECT 28.775 113.425 28.945 114.270 ;
        RECT 29.840 113.985 30.010 114.485 ;
        RECT 30.180 114.155 30.510 114.655 ;
        RECT 29.115 113.595 29.615 113.975 ;
        RECT 29.840 113.815 30.535 113.985 ;
        RECT 27.595 113.255 28.945 113.425 ;
        RECT 28.525 113.215 28.945 113.255 ;
        RECT 27.235 112.745 27.655 113.085 ;
        RECT 27.945 112.755 28.355 113.085 ;
        RECT 25.475 112.325 26.325 112.495 ;
        RECT 26.885 112.105 27.205 112.565 ;
        RECT 27.405 112.315 27.655 112.745 ;
        RECT 27.945 112.105 28.355 112.545 ;
        RECT 28.525 112.485 28.695 113.215 ;
        RECT 28.865 112.665 29.215 113.035 ;
        RECT 29.395 112.725 29.615 113.595 ;
        RECT 29.785 113.025 30.195 113.645 ;
        RECT 30.365 112.845 30.535 113.815 ;
        RECT 29.840 112.655 30.535 112.845 ;
        RECT 28.525 112.285 29.540 112.485 ;
        RECT 29.840 112.325 30.010 112.655 ;
        RECT 30.180 112.105 30.510 112.485 ;
        RECT 30.725 112.365 30.950 114.485 ;
        RECT 31.120 114.155 31.450 114.655 ;
        RECT 31.620 113.985 31.790 114.485 ;
        RECT 31.125 113.815 31.790 113.985 ;
        RECT 31.125 112.825 31.355 113.815 ;
        RECT 31.525 112.995 31.875 113.645 ;
        RECT 32.050 113.580 32.320 114.485 ;
        RECT 32.490 113.895 32.820 114.655 ;
        RECT 33.000 113.725 33.170 114.485 ;
        RECT 31.125 112.655 31.790 112.825 ;
        RECT 31.120 112.105 31.450 112.485 ;
        RECT 31.620 112.365 31.790 112.655 ;
        RECT 32.050 112.780 32.220 113.580 ;
        RECT 32.505 113.555 33.170 113.725 ;
        RECT 33.520 113.725 33.690 114.485 ;
        RECT 33.870 113.895 34.200 114.655 ;
        RECT 33.520 113.555 34.185 113.725 ;
        RECT 34.370 113.580 34.640 114.485 ;
        RECT 32.505 113.410 32.675 113.555 ;
        RECT 32.390 113.080 32.675 113.410 ;
        RECT 34.015 113.410 34.185 113.555 ;
        RECT 32.505 112.825 32.675 113.080 ;
        RECT 32.910 113.005 33.240 113.375 ;
        RECT 33.450 113.005 33.780 113.375 ;
        RECT 34.015 113.080 34.300 113.410 ;
        RECT 34.015 112.825 34.185 113.080 ;
        RECT 32.050 112.275 32.310 112.780 ;
        RECT 32.505 112.655 33.170 112.825 ;
        RECT 32.490 112.105 32.820 112.485 ;
        RECT 33.000 112.275 33.170 112.655 ;
        RECT 33.520 112.655 34.185 112.825 ;
        RECT 34.470 112.780 34.640 113.580 ;
        RECT 34.810 113.490 35.100 114.655 ;
        RECT 35.360 113.985 35.530 114.485 ;
        RECT 35.700 114.155 36.030 114.655 ;
        RECT 35.360 113.815 36.025 113.985 ;
        RECT 35.275 112.995 35.625 113.645 ;
        RECT 33.520 112.275 33.690 112.655 ;
        RECT 33.870 112.105 34.200 112.485 ;
        RECT 34.380 112.275 34.640 112.780 ;
        RECT 34.810 112.105 35.100 112.830 ;
        RECT 35.795 112.825 36.025 113.815 ;
        RECT 35.360 112.655 36.025 112.825 ;
        RECT 35.360 112.365 35.530 112.655 ;
        RECT 35.700 112.105 36.030 112.485 ;
        RECT 36.200 112.365 36.425 114.485 ;
        RECT 36.640 114.155 36.970 114.655 ;
        RECT 37.140 113.985 37.310 114.485 ;
        RECT 37.545 114.270 38.375 114.440 ;
        RECT 38.615 114.275 38.995 114.655 ;
        RECT 36.615 113.815 37.310 113.985 ;
        RECT 36.615 112.845 36.785 113.815 ;
        RECT 36.955 113.025 37.365 113.645 ;
        RECT 37.535 113.595 38.035 113.975 ;
        RECT 36.615 112.655 37.310 112.845 ;
        RECT 37.535 112.725 37.755 113.595 ;
        RECT 38.205 113.425 38.375 114.270 ;
        RECT 39.175 114.105 39.345 114.395 ;
        RECT 39.515 114.275 39.845 114.655 ;
        RECT 40.315 114.185 40.945 114.435 ;
        RECT 41.125 114.275 41.545 114.655 ;
        RECT 40.775 114.105 40.945 114.185 ;
        RECT 41.745 114.105 41.985 114.395 ;
        RECT 38.545 113.855 39.915 114.105 ;
        RECT 38.545 113.595 38.795 113.855 ;
        RECT 39.305 113.425 39.555 113.585 ;
        RECT 38.205 113.255 39.555 113.425 ;
        RECT 38.205 113.215 38.625 113.255 ;
        RECT 37.935 112.665 38.285 113.035 ;
        RECT 36.640 112.105 36.970 112.485 ;
        RECT 37.140 112.325 37.310 112.655 ;
        RECT 38.455 112.485 38.625 113.215 ;
        RECT 39.725 113.085 39.915 113.855 ;
        RECT 38.795 112.755 39.205 113.085 ;
        RECT 39.495 112.745 39.915 113.085 ;
        RECT 40.085 113.675 40.605 113.985 ;
        RECT 40.775 113.935 41.985 114.105 ;
        RECT 42.215 113.965 42.545 114.655 ;
        RECT 40.085 112.915 40.255 113.675 ;
        RECT 40.425 113.085 40.605 113.495 ;
        RECT 40.775 113.425 40.945 113.935 ;
        RECT 42.715 113.785 42.885 114.395 ;
        RECT 43.155 113.935 43.485 114.445 ;
        RECT 42.715 113.765 43.035 113.785 ;
        RECT 41.115 113.595 43.035 113.765 ;
        RECT 40.775 113.255 42.675 113.425 ;
        RECT 41.005 112.915 41.335 113.035 ;
        RECT 40.085 112.745 41.335 112.915 ;
        RECT 37.610 112.285 38.625 112.485 ;
        RECT 38.795 112.105 39.205 112.545 ;
        RECT 39.495 112.315 39.745 112.745 ;
        RECT 39.945 112.105 40.265 112.565 ;
        RECT 41.505 112.495 41.675 113.255 ;
        RECT 42.345 113.195 42.675 113.255 ;
        RECT 41.865 113.025 42.195 113.085 ;
        RECT 41.865 112.755 42.525 113.025 ;
        RECT 42.845 112.700 43.035 113.595 ;
        RECT 40.825 112.325 41.675 112.495 ;
        RECT 41.875 112.105 42.535 112.585 ;
        RECT 42.715 112.370 43.035 112.700 ;
        RECT 43.235 113.345 43.485 113.935 ;
        RECT 43.665 113.855 43.950 114.655 ;
        RECT 44.130 113.675 44.385 114.345 ;
        RECT 43.235 113.015 44.035 113.345 ;
        RECT 44.205 113.295 44.385 113.675 ;
        RECT 45.850 113.580 46.120 114.485 ;
        RECT 46.290 113.895 46.620 114.655 ;
        RECT 46.800 113.725 46.970 114.485 ;
        RECT 44.205 113.125 44.470 113.295 ;
        RECT 43.235 112.365 43.485 113.015 ;
        RECT 44.205 112.815 44.385 113.125 ;
        RECT 43.665 112.105 43.950 112.565 ;
        RECT 44.130 112.285 44.385 112.815 ;
        RECT 45.850 112.780 46.020 113.580 ;
        RECT 46.305 113.555 46.970 113.725 ;
        RECT 46.305 113.410 46.475 113.555 ;
        RECT 47.270 113.515 47.500 114.655 ;
        RECT 47.670 113.505 48.000 114.485 ;
        RECT 48.170 113.515 48.380 114.655 ;
        RECT 48.985 114.315 49.240 114.345 ;
        RECT 48.900 114.145 49.240 114.315 ;
        RECT 48.985 113.675 49.240 114.145 ;
        RECT 49.420 113.855 49.705 114.655 ;
        RECT 49.885 113.935 50.215 114.445 ;
        RECT 46.190 113.080 46.475 113.410 ;
        RECT 46.305 112.825 46.475 113.080 ;
        RECT 46.710 113.005 47.040 113.375 ;
        RECT 47.250 113.095 47.580 113.345 ;
        RECT 45.850 112.275 46.110 112.780 ;
        RECT 46.305 112.655 46.970 112.825 ;
        RECT 46.290 112.105 46.620 112.485 ;
        RECT 46.800 112.275 46.970 112.655 ;
        RECT 47.270 112.105 47.500 112.925 ;
        RECT 47.750 112.905 48.000 113.505 ;
        RECT 47.670 112.275 48.000 112.905 ;
        RECT 48.170 112.105 48.380 112.925 ;
        RECT 48.985 112.815 49.165 113.675 ;
        RECT 49.885 113.345 50.135 113.935 ;
        RECT 50.485 113.785 50.655 114.395 ;
        RECT 50.825 113.965 51.155 114.655 ;
        RECT 51.385 114.105 51.625 114.395 ;
        RECT 51.825 114.275 52.245 114.655 ;
        RECT 52.425 114.185 53.055 114.435 ;
        RECT 53.525 114.275 53.855 114.655 ;
        RECT 52.425 114.105 52.595 114.185 ;
        RECT 54.025 114.105 54.195 114.395 ;
        RECT 54.375 114.275 54.755 114.655 ;
        RECT 54.995 114.270 55.825 114.440 ;
        RECT 51.385 113.935 52.595 114.105 ;
        RECT 49.335 113.015 50.135 113.345 ;
        RECT 48.985 112.285 49.240 112.815 ;
        RECT 49.420 112.105 49.705 112.565 ;
        RECT 49.885 112.365 50.135 113.015 ;
        RECT 50.335 113.765 50.655 113.785 ;
        RECT 50.335 113.595 52.255 113.765 ;
        RECT 50.335 112.700 50.525 113.595 ;
        RECT 52.425 113.425 52.595 113.935 ;
        RECT 52.765 113.675 53.285 113.985 ;
        RECT 50.695 113.255 52.595 113.425 ;
        RECT 50.695 113.195 51.025 113.255 ;
        RECT 51.175 113.025 51.505 113.085 ;
        RECT 50.845 112.755 51.505 113.025 ;
        RECT 50.335 112.370 50.655 112.700 ;
        RECT 50.835 112.105 51.495 112.585 ;
        RECT 51.695 112.495 51.865 113.255 ;
        RECT 52.765 113.085 52.945 113.495 ;
        RECT 52.035 112.915 52.365 113.035 ;
        RECT 53.115 112.915 53.285 113.675 ;
        RECT 52.035 112.745 53.285 112.915 ;
        RECT 53.455 113.855 54.825 114.105 ;
        RECT 53.455 113.085 53.645 113.855 ;
        RECT 54.575 113.595 54.825 113.855 ;
        RECT 53.815 113.425 54.065 113.585 ;
        RECT 54.995 113.425 55.165 114.270 ;
        RECT 56.060 113.985 56.230 114.485 ;
        RECT 56.400 114.155 56.730 114.655 ;
        RECT 55.335 113.595 55.835 113.975 ;
        RECT 56.060 113.815 56.755 113.985 ;
        RECT 53.815 113.255 55.165 113.425 ;
        RECT 54.745 113.215 55.165 113.255 ;
        RECT 53.455 112.745 53.875 113.085 ;
        RECT 54.165 112.755 54.575 113.085 ;
        RECT 51.695 112.325 52.545 112.495 ;
        RECT 53.105 112.105 53.425 112.565 ;
        RECT 53.625 112.315 53.875 112.745 ;
        RECT 54.165 112.105 54.575 112.545 ;
        RECT 54.745 112.485 54.915 113.215 ;
        RECT 55.085 112.665 55.435 113.035 ;
        RECT 55.615 112.725 55.835 113.595 ;
        RECT 56.005 113.025 56.415 113.645 ;
        RECT 56.585 112.845 56.755 113.815 ;
        RECT 56.060 112.655 56.755 112.845 ;
        RECT 54.745 112.285 55.760 112.485 ;
        RECT 56.060 112.325 56.230 112.655 ;
        RECT 56.400 112.105 56.730 112.485 ;
        RECT 56.945 112.365 57.170 114.485 ;
        RECT 57.340 114.155 57.670 114.655 ;
        RECT 57.840 113.985 58.010 114.485 ;
        RECT 57.345 113.815 58.010 113.985 ;
        RECT 57.345 112.825 57.575 113.815 ;
        RECT 57.745 112.995 58.095 113.645 ;
        RECT 58.730 113.565 60.400 114.655 ;
        RECT 58.730 113.045 59.480 113.565 ;
        RECT 60.570 113.490 60.860 114.655 ;
        RECT 61.530 113.515 61.760 114.655 ;
        RECT 61.930 113.505 62.260 114.485 ;
        RECT 62.430 113.515 62.640 114.655 ;
        RECT 63.335 114.220 68.680 114.655 ;
        RECT 59.650 112.875 60.400 113.395 ;
        RECT 61.510 113.095 61.840 113.345 ;
        RECT 57.345 112.655 58.010 112.825 ;
        RECT 57.340 112.105 57.670 112.485 ;
        RECT 57.840 112.365 58.010 112.655 ;
        RECT 58.730 112.105 60.400 112.875 ;
        RECT 60.570 112.105 60.860 112.830 ;
        RECT 61.530 112.105 61.760 112.925 ;
        RECT 62.010 112.905 62.260 113.505 ;
        RECT 64.925 112.970 65.275 114.220 ;
        RECT 68.910 113.515 69.120 114.655 ;
        RECT 69.290 113.505 69.620 114.485 ;
        RECT 69.790 113.515 70.020 114.655 ;
        RECT 70.320 113.985 70.490 114.485 ;
        RECT 70.660 114.155 70.990 114.655 ;
        RECT 70.320 113.815 70.985 113.985 ;
        RECT 61.930 112.275 62.260 112.905 ;
        RECT 62.430 112.105 62.640 112.925 ;
        RECT 66.755 112.650 67.095 113.480 ;
        RECT 63.335 112.105 68.680 112.650 ;
        RECT 68.910 112.105 69.120 112.925 ;
        RECT 69.290 112.905 69.540 113.505 ;
        RECT 69.710 113.095 70.040 113.345 ;
        RECT 70.235 112.995 70.585 113.645 ;
        RECT 69.290 112.275 69.620 112.905 ;
        RECT 69.790 112.105 70.020 112.925 ;
        RECT 70.755 112.825 70.985 113.815 ;
        RECT 70.320 112.655 70.985 112.825 ;
        RECT 70.320 112.365 70.490 112.655 ;
        RECT 70.660 112.105 70.990 112.485 ;
        RECT 71.160 112.365 71.385 114.485 ;
        RECT 71.600 114.155 71.930 114.655 ;
        RECT 72.100 113.985 72.270 114.485 ;
        RECT 72.505 114.270 73.335 114.440 ;
        RECT 73.575 114.275 73.955 114.655 ;
        RECT 71.575 113.815 72.270 113.985 ;
        RECT 71.575 112.845 71.745 113.815 ;
        RECT 71.915 113.025 72.325 113.645 ;
        RECT 72.495 113.595 72.995 113.975 ;
        RECT 71.575 112.655 72.270 112.845 ;
        RECT 72.495 112.725 72.715 113.595 ;
        RECT 73.165 113.425 73.335 114.270 ;
        RECT 74.135 114.105 74.305 114.395 ;
        RECT 74.475 114.275 74.805 114.655 ;
        RECT 75.275 114.185 75.905 114.435 ;
        RECT 76.085 114.275 76.505 114.655 ;
        RECT 75.735 114.105 75.905 114.185 ;
        RECT 76.705 114.105 76.945 114.395 ;
        RECT 73.505 113.855 74.875 114.105 ;
        RECT 73.505 113.595 73.755 113.855 ;
        RECT 74.265 113.425 74.515 113.585 ;
        RECT 73.165 113.255 74.515 113.425 ;
        RECT 73.165 113.215 73.585 113.255 ;
        RECT 72.895 112.665 73.245 113.035 ;
        RECT 71.600 112.105 71.930 112.485 ;
        RECT 72.100 112.325 72.270 112.655 ;
        RECT 73.415 112.485 73.585 113.215 ;
        RECT 74.685 113.085 74.875 113.855 ;
        RECT 73.755 112.755 74.165 113.085 ;
        RECT 74.455 112.745 74.875 113.085 ;
        RECT 75.045 113.675 75.565 113.985 ;
        RECT 75.735 113.935 76.945 114.105 ;
        RECT 77.175 113.965 77.505 114.655 ;
        RECT 75.045 112.915 75.215 113.675 ;
        RECT 75.385 113.085 75.565 113.495 ;
        RECT 75.735 113.425 75.905 113.935 ;
        RECT 77.675 113.785 77.845 114.395 ;
        RECT 78.115 113.935 78.445 114.445 ;
        RECT 77.675 113.765 77.995 113.785 ;
        RECT 76.075 113.595 77.995 113.765 ;
        RECT 75.735 113.255 77.635 113.425 ;
        RECT 75.965 112.915 76.295 113.035 ;
        RECT 75.045 112.745 76.295 112.915 ;
        RECT 72.570 112.285 73.585 112.485 ;
        RECT 73.755 112.105 74.165 112.545 ;
        RECT 74.455 112.315 74.705 112.745 ;
        RECT 74.905 112.105 75.225 112.565 ;
        RECT 76.465 112.495 76.635 113.255 ;
        RECT 77.305 113.195 77.635 113.255 ;
        RECT 76.825 113.025 77.155 113.085 ;
        RECT 76.825 112.755 77.485 113.025 ;
        RECT 77.805 112.700 77.995 113.595 ;
        RECT 75.785 112.325 76.635 112.495 ;
        RECT 76.835 112.105 77.495 112.585 ;
        RECT 77.675 112.370 77.995 112.700 ;
        RECT 78.195 113.345 78.445 113.935 ;
        RECT 78.625 113.855 78.910 114.655 ;
        RECT 79.090 114.315 79.345 114.345 ;
        RECT 79.090 114.145 79.430 114.315 ;
        RECT 79.090 113.675 79.345 114.145 ;
        RECT 78.195 113.015 78.995 113.345 ;
        RECT 78.195 112.365 78.445 113.015 ;
        RECT 79.165 112.815 79.345 113.675 ;
        RECT 78.625 112.105 78.910 112.565 ;
        RECT 79.090 112.285 79.345 112.815 ;
        RECT 79.890 113.580 80.160 114.485 ;
        RECT 80.330 113.895 80.660 114.655 ;
        RECT 80.840 113.725 81.010 114.485 ;
        RECT 79.890 112.780 80.060 113.580 ;
        RECT 80.345 113.555 81.010 113.725 ;
        RECT 80.345 113.410 80.515 113.555 ;
        RECT 81.330 113.515 81.540 114.655 ;
        RECT 80.230 113.080 80.515 113.410 ;
        RECT 81.710 113.505 82.040 114.485 ;
        RECT 82.210 113.515 82.440 114.655 ;
        RECT 82.710 113.515 82.920 114.655 ;
        RECT 83.090 113.505 83.420 114.485 ;
        RECT 83.590 113.515 83.820 114.655 ;
        RECT 84.990 113.515 85.220 114.655 ;
        RECT 85.390 113.505 85.720 114.485 ;
        RECT 85.890 113.515 86.100 114.655 ;
        RECT 80.345 112.825 80.515 113.080 ;
        RECT 80.750 113.005 81.080 113.375 ;
        RECT 79.890 112.275 80.150 112.780 ;
        RECT 80.345 112.655 81.010 112.825 ;
        RECT 80.330 112.105 80.660 112.485 ;
        RECT 80.840 112.275 81.010 112.655 ;
        RECT 81.330 112.105 81.540 112.925 ;
        RECT 81.710 112.905 81.960 113.505 ;
        RECT 82.130 113.095 82.460 113.345 ;
        RECT 81.710 112.275 82.040 112.905 ;
        RECT 82.210 112.105 82.440 112.925 ;
        RECT 82.710 112.105 82.920 112.925 ;
        RECT 83.090 112.905 83.340 113.505 ;
        RECT 83.510 113.095 83.840 113.345 ;
        RECT 84.970 113.095 85.300 113.345 ;
        RECT 83.090 112.275 83.420 112.905 ;
        RECT 83.590 112.105 83.820 112.925 ;
        RECT 84.990 112.105 85.220 112.925 ;
        RECT 85.470 112.905 85.720 113.505 ;
        RECT 86.330 113.490 86.620 114.655 ;
        RECT 87.165 114.315 87.420 114.345 ;
        RECT 87.080 114.145 87.420 114.315 ;
        RECT 87.165 113.675 87.420 114.145 ;
        RECT 87.600 113.855 87.885 114.655 ;
        RECT 88.065 113.935 88.395 114.445 ;
        RECT 85.390 112.275 85.720 112.905 ;
        RECT 85.890 112.105 86.100 112.925 ;
        RECT 86.330 112.105 86.620 112.830 ;
        RECT 87.165 112.815 87.345 113.675 ;
        RECT 88.065 113.345 88.315 113.935 ;
        RECT 88.665 113.785 88.835 114.395 ;
        RECT 89.005 113.965 89.335 114.655 ;
        RECT 89.565 114.105 89.805 114.395 ;
        RECT 90.005 114.275 90.425 114.655 ;
        RECT 90.605 114.185 91.235 114.435 ;
        RECT 91.705 114.275 92.035 114.655 ;
        RECT 90.605 114.105 90.775 114.185 ;
        RECT 92.205 114.105 92.375 114.395 ;
        RECT 92.555 114.275 92.935 114.655 ;
        RECT 93.175 114.270 94.005 114.440 ;
        RECT 89.565 113.935 90.775 114.105 ;
        RECT 87.515 113.015 88.315 113.345 ;
        RECT 87.165 112.285 87.420 112.815 ;
        RECT 87.600 112.105 87.885 112.565 ;
        RECT 88.065 112.365 88.315 113.015 ;
        RECT 88.515 113.765 88.835 113.785 ;
        RECT 88.515 113.595 90.435 113.765 ;
        RECT 88.515 112.700 88.705 113.595 ;
        RECT 90.605 113.425 90.775 113.935 ;
        RECT 90.945 113.675 91.465 113.985 ;
        RECT 88.875 113.255 90.775 113.425 ;
        RECT 88.875 113.195 89.205 113.255 ;
        RECT 89.355 113.025 89.685 113.085 ;
        RECT 89.025 112.755 89.685 113.025 ;
        RECT 88.515 112.370 88.835 112.700 ;
        RECT 89.015 112.105 89.675 112.585 ;
        RECT 89.875 112.495 90.045 113.255 ;
        RECT 90.945 113.085 91.125 113.495 ;
        RECT 90.215 112.915 90.545 113.035 ;
        RECT 91.295 112.915 91.465 113.675 ;
        RECT 90.215 112.745 91.465 112.915 ;
        RECT 91.635 113.855 93.005 114.105 ;
        RECT 91.635 113.085 91.825 113.855 ;
        RECT 92.755 113.595 93.005 113.855 ;
        RECT 91.995 113.425 92.245 113.585 ;
        RECT 93.175 113.425 93.345 114.270 ;
        RECT 94.240 113.985 94.410 114.485 ;
        RECT 94.580 114.155 94.910 114.655 ;
        RECT 93.515 113.595 94.015 113.975 ;
        RECT 94.240 113.815 94.935 113.985 ;
        RECT 91.995 113.255 93.345 113.425 ;
        RECT 92.925 113.215 93.345 113.255 ;
        RECT 91.635 112.745 92.055 113.085 ;
        RECT 92.345 112.755 92.755 113.085 ;
        RECT 89.875 112.325 90.725 112.495 ;
        RECT 91.285 112.105 91.605 112.565 ;
        RECT 91.805 112.315 92.055 112.745 ;
        RECT 92.345 112.105 92.755 112.545 ;
        RECT 92.925 112.485 93.095 113.215 ;
        RECT 93.265 112.665 93.615 113.035 ;
        RECT 93.795 112.725 94.015 113.595 ;
        RECT 94.185 113.025 94.595 113.645 ;
        RECT 94.765 112.845 94.935 113.815 ;
        RECT 94.240 112.655 94.935 112.845 ;
        RECT 92.925 112.285 93.940 112.485 ;
        RECT 94.240 112.325 94.410 112.655 ;
        RECT 94.580 112.105 94.910 112.485 ;
        RECT 95.125 112.365 95.350 114.485 ;
        RECT 95.520 114.155 95.850 114.655 ;
        RECT 96.020 113.985 96.190 114.485 ;
        RECT 95.525 113.815 96.190 113.985 ;
        RECT 95.525 112.825 95.755 113.815 ;
        RECT 95.925 112.995 96.275 113.645 ;
        RECT 96.450 113.580 96.720 114.485 ;
        RECT 96.890 113.895 97.220 114.655 ;
        RECT 97.400 113.725 97.570 114.485 ;
        RECT 98.755 114.220 104.100 114.655 ;
        RECT 95.525 112.655 96.190 112.825 ;
        RECT 95.520 112.105 95.850 112.485 ;
        RECT 96.020 112.365 96.190 112.655 ;
        RECT 96.450 112.780 96.620 113.580 ;
        RECT 96.905 113.555 97.570 113.725 ;
        RECT 96.905 113.410 97.075 113.555 ;
        RECT 96.790 113.080 97.075 113.410 ;
        RECT 96.905 112.825 97.075 113.080 ;
        RECT 97.310 113.005 97.640 113.375 ;
        RECT 100.345 112.970 100.695 114.220 ;
        RECT 104.310 113.515 104.540 114.655 ;
        RECT 104.710 113.505 105.040 114.485 ;
        RECT 105.210 113.515 105.420 114.655 ;
        RECT 106.200 113.725 106.370 114.485 ;
        RECT 106.550 113.895 106.880 114.655 ;
        RECT 106.200 113.555 106.865 113.725 ;
        RECT 107.050 113.580 107.320 114.485 ;
        RECT 96.450 112.275 96.710 112.780 ;
        RECT 96.905 112.655 97.570 112.825 ;
        RECT 96.890 112.105 97.220 112.485 ;
        RECT 97.400 112.275 97.570 112.655 ;
        RECT 102.175 112.650 102.515 113.480 ;
        RECT 104.290 113.095 104.620 113.345 ;
        RECT 98.755 112.105 104.100 112.650 ;
        RECT 104.310 112.105 104.540 112.925 ;
        RECT 104.790 112.905 105.040 113.505 ;
        RECT 106.695 113.410 106.865 113.555 ;
        RECT 106.130 113.005 106.460 113.375 ;
        RECT 106.695 113.080 106.980 113.410 ;
        RECT 104.710 112.275 105.040 112.905 ;
        RECT 105.210 112.105 105.420 112.925 ;
        RECT 106.695 112.825 106.865 113.080 ;
        RECT 106.200 112.655 106.865 112.825 ;
        RECT 107.150 112.780 107.320 113.580 ;
        RECT 107.490 113.565 111.000 114.655 ;
        RECT 111.170 113.565 112.380 114.655 ;
        RECT 107.490 113.045 109.180 113.565 ;
        RECT 109.350 112.875 111.000 113.395 ;
        RECT 111.170 113.025 111.690 113.565 ;
        RECT 106.200 112.275 106.370 112.655 ;
        RECT 106.550 112.105 106.880 112.485 ;
        RECT 107.060 112.275 107.320 112.780 ;
        RECT 107.490 112.105 111.000 112.875 ;
        RECT 111.860 112.855 112.380 113.395 ;
        RECT 111.170 112.105 112.380 112.855 ;
        RECT 18.165 111.935 112.465 112.105 ;
        RECT 18.250 111.185 19.460 111.935 ;
        RECT 20.640 111.385 20.810 111.765 ;
        RECT 20.990 111.555 21.320 111.935 ;
        RECT 20.640 111.215 21.305 111.385 ;
        RECT 21.500 111.260 21.760 111.765 ;
        RECT 18.250 110.645 18.770 111.185 ;
        RECT 18.940 110.475 19.460 111.015 ;
        RECT 20.570 110.665 20.900 111.035 ;
        RECT 21.135 110.960 21.305 111.215 ;
        RECT 21.135 110.630 21.420 110.960 ;
        RECT 21.135 110.485 21.305 110.630 ;
        RECT 18.250 109.385 19.460 110.475 ;
        RECT 20.640 110.315 21.305 110.485 ;
        RECT 21.590 110.460 21.760 111.260 ;
        RECT 21.930 111.210 22.220 111.935 ;
        RECT 23.315 111.195 23.570 111.765 ;
        RECT 23.740 111.535 24.070 111.935 ;
        RECT 24.495 111.400 25.025 111.765 ;
        RECT 24.495 111.365 24.670 111.400 ;
        RECT 23.740 111.195 24.670 111.365 ;
        RECT 25.215 111.255 25.490 111.765 ;
        RECT 20.640 109.555 20.810 110.315 ;
        RECT 20.990 109.385 21.320 110.145 ;
        RECT 21.490 109.555 21.760 110.460 ;
        RECT 21.930 109.385 22.220 110.550 ;
        RECT 23.315 110.525 23.485 111.195 ;
        RECT 23.740 111.025 23.910 111.195 ;
        RECT 23.655 110.695 23.910 111.025 ;
        RECT 24.135 110.695 24.330 111.025 ;
        RECT 23.315 109.555 23.650 110.525 ;
        RECT 23.820 109.385 23.990 110.525 ;
        RECT 24.160 109.725 24.330 110.695 ;
        RECT 24.500 110.065 24.670 111.195 ;
        RECT 24.840 110.405 25.010 111.205 ;
        RECT 25.210 111.085 25.490 111.255 ;
        RECT 25.215 110.605 25.490 111.085 ;
        RECT 25.660 110.405 25.850 111.765 ;
        RECT 26.030 111.400 26.540 111.935 ;
        RECT 26.760 111.125 27.005 111.730 ;
        RECT 26.050 110.955 27.280 111.125 ;
        RECT 27.490 111.115 27.720 111.935 ;
        RECT 27.890 111.135 28.220 111.765 ;
        RECT 24.840 110.235 25.850 110.405 ;
        RECT 26.020 110.390 26.770 110.580 ;
        RECT 24.500 109.895 25.625 110.065 ;
        RECT 26.020 109.725 26.190 110.390 ;
        RECT 26.940 110.145 27.280 110.955 ;
        RECT 27.470 110.695 27.800 110.945 ;
        RECT 27.970 110.535 28.220 111.135 ;
        RECT 28.390 111.115 28.600 111.935 ;
        RECT 29.140 111.465 29.310 111.935 ;
        RECT 29.480 111.285 29.810 111.765 ;
        RECT 29.980 111.465 30.150 111.935 ;
        RECT 30.320 111.285 30.650 111.765 ;
        RECT 28.885 111.115 30.650 111.285 ;
        RECT 30.820 111.125 30.990 111.935 ;
        RECT 31.190 111.555 32.260 111.725 ;
        RECT 31.190 111.200 31.510 111.555 ;
        RECT 24.160 109.555 26.190 109.725 ;
        RECT 26.360 109.385 26.530 110.145 ;
        RECT 26.765 109.735 27.280 110.145 ;
        RECT 27.490 109.385 27.720 110.525 ;
        RECT 27.890 109.555 28.220 110.535 ;
        RECT 28.885 110.565 29.295 111.115 ;
        RECT 31.185 110.945 31.510 111.200 ;
        RECT 29.480 110.735 31.510 110.945 ;
        RECT 31.165 110.725 31.510 110.735 ;
        RECT 31.680 110.985 31.920 111.385 ;
        RECT 32.090 111.325 32.260 111.555 ;
        RECT 32.430 111.495 32.620 111.935 ;
        RECT 32.790 111.485 33.740 111.765 ;
        RECT 33.960 111.575 34.310 111.745 ;
        RECT 32.090 111.155 32.620 111.325 ;
        RECT 28.390 109.385 28.600 110.525 ;
        RECT 28.885 110.395 30.610 110.565 ;
        RECT 29.140 109.385 29.310 110.225 ;
        RECT 29.520 109.555 29.770 110.395 ;
        RECT 29.980 109.385 30.150 110.225 ;
        RECT 30.320 109.555 30.610 110.395 ;
        RECT 30.820 109.385 30.990 110.445 ;
        RECT 31.165 110.105 31.335 110.725 ;
        RECT 31.680 110.615 32.220 110.985 ;
        RECT 32.400 110.875 32.620 111.155 ;
        RECT 32.790 110.705 32.960 111.485 ;
        RECT 32.555 110.535 32.960 110.705 ;
        RECT 33.130 110.695 33.480 111.315 ;
        RECT 32.555 110.445 32.725 110.535 ;
        RECT 33.650 110.525 33.860 111.315 ;
        RECT 31.505 110.275 32.725 110.445 ;
        RECT 33.185 110.365 33.860 110.525 ;
        RECT 31.165 109.935 31.965 110.105 ;
        RECT 31.285 109.385 31.615 109.765 ;
        RECT 31.795 109.645 31.965 109.935 ;
        RECT 32.555 109.895 32.725 110.275 ;
        RECT 32.895 110.355 33.860 110.365 ;
        RECT 34.050 111.185 34.310 111.575 ;
        RECT 34.520 111.475 34.850 111.935 ;
        RECT 35.725 111.545 36.580 111.715 ;
        RECT 36.785 111.545 37.280 111.715 ;
        RECT 37.450 111.575 37.780 111.935 ;
        RECT 34.050 110.495 34.220 111.185 ;
        RECT 34.390 110.835 34.560 111.015 ;
        RECT 34.730 111.005 35.520 111.255 ;
        RECT 35.725 110.835 35.895 111.545 ;
        RECT 36.065 111.035 36.420 111.255 ;
        RECT 34.390 110.665 36.080 110.835 ;
        RECT 32.895 110.065 33.355 110.355 ;
        RECT 34.050 110.325 35.550 110.495 ;
        RECT 34.050 110.185 34.220 110.325 ;
        RECT 33.660 110.015 34.220 110.185 ;
        RECT 32.135 109.385 32.385 109.845 ;
        RECT 32.555 109.555 33.425 109.895 ;
        RECT 33.660 109.555 33.830 110.015 ;
        RECT 34.665 109.985 35.740 110.155 ;
        RECT 34.000 109.385 34.370 109.845 ;
        RECT 34.665 109.645 34.835 109.985 ;
        RECT 35.005 109.385 35.335 109.815 ;
        RECT 35.570 109.645 35.740 109.985 ;
        RECT 35.910 109.885 36.080 110.665 ;
        RECT 36.250 110.445 36.420 111.035 ;
        RECT 36.590 110.635 36.940 111.255 ;
        RECT 36.250 110.055 36.715 110.445 ;
        RECT 37.110 110.185 37.280 111.545 ;
        RECT 37.450 110.355 37.910 111.405 ;
        RECT 36.885 110.015 37.280 110.185 ;
        RECT 36.885 109.885 37.055 110.015 ;
        RECT 35.910 109.555 36.590 109.885 ;
        RECT 36.805 109.555 37.055 109.885 ;
        RECT 37.225 109.385 37.475 109.845 ;
        RECT 37.645 109.570 37.970 110.355 ;
        RECT 38.140 109.555 38.310 111.675 ;
        RECT 38.480 111.555 38.810 111.935 ;
        RECT 38.980 111.385 39.235 111.675 ;
        RECT 38.485 111.215 39.235 111.385 ;
        RECT 38.485 110.225 38.715 111.215 ;
        RECT 39.410 111.165 42.000 111.935 ;
        RECT 42.175 111.390 47.520 111.935 ;
        RECT 38.885 110.395 39.235 111.045 ;
        RECT 39.410 110.475 40.620 110.995 ;
        RECT 40.790 110.645 42.000 111.165 ;
        RECT 38.485 110.055 39.235 110.225 ;
        RECT 38.480 109.385 38.810 109.885 ;
        RECT 38.980 109.555 39.235 110.055 ;
        RECT 39.410 109.385 42.000 110.475 ;
        RECT 43.765 109.820 44.115 111.070 ;
        RECT 45.595 110.560 45.935 111.390 ;
        RECT 47.690 111.210 47.980 111.935 ;
        RECT 49.160 111.385 49.330 111.765 ;
        RECT 49.510 111.555 49.840 111.935 ;
        RECT 49.160 111.215 49.825 111.385 ;
        RECT 50.020 111.260 50.280 111.765 ;
        RECT 49.090 110.665 49.420 111.035 ;
        RECT 49.655 110.960 49.825 111.215 ;
        RECT 49.655 110.630 49.940 110.960 ;
        RECT 42.175 109.385 47.520 109.820 ;
        RECT 47.690 109.385 47.980 110.550 ;
        RECT 49.655 110.485 49.825 110.630 ;
        RECT 49.160 110.315 49.825 110.485 ;
        RECT 50.110 110.460 50.280 111.260 ;
        RECT 50.490 111.115 50.720 111.935 ;
        RECT 50.890 111.135 51.220 111.765 ;
        RECT 50.470 110.695 50.800 110.945 ;
        RECT 50.970 110.535 51.220 111.135 ;
        RECT 51.390 111.115 51.600 111.935 ;
        RECT 51.920 111.385 52.090 111.765 ;
        RECT 52.270 111.555 52.600 111.935 ;
        RECT 51.920 111.215 52.585 111.385 ;
        RECT 52.780 111.260 53.040 111.765 ;
        RECT 51.850 110.665 52.180 111.035 ;
        RECT 52.415 110.960 52.585 111.215 ;
        RECT 49.160 109.555 49.330 110.315 ;
        RECT 49.510 109.385 49.840 110.145 ;
        RECT 50.010 109.555 50.280 110.460 ;
        RECT 50.490 109.385 50.720 110.525 ;
        RECT 50.890 109.555 51.220 110.535 ;
        RECT 52.415 110.630 52.700 110.960 ;
        RECT 51.390 109.385 51.600 110.525 ;
        RECT 52.415 110.485 52.585 110.630 ;
        RECT 51.920 110.315 52.585 110.485 ;
        RECT 52.870 110.460 53.040 111.260 ;
        RECT 53.360 111.135 53.690 111.935 ;
        RECT 53.860 111.285 54.030 111.765 ;
        RECT 54.200 111.455 54.530 111.935 ;
        RECT 54.700 111.285 54.870 111.765 ;
        RECT 55.120 111.455 55.360 111.935 ;
        RECT 55.540 111.285 55.710 111.765 ;
        RECT 56.280 111.465 56.450 111.935 ;
        RECT 56.620 111.285 56.950 111.765 ;
        RECT 57.120 111.465 57.290 111.935 ;
        RECT 57.460 111.285 57.790 111.765 ;
        RECT 53.860 111.115 54.870 111.285 ;
        RECT 55.075 111.115 55.710 111.285 ;
        RECT 56.025 111.115 57.790 111.285 ;
        RECT 57.960 111.125 58.130 111.935 ;
        RECT 58.330 111.555 59.400 111.725 ;
        RECT 58.330 111.200 58.650 111.555 ;
        RECT 53.860 111.085 54.360 111.115 ;
        RECT 53.860 110.575 54.355 111.085 ;
        RECT 55.075 110.945 55.245 111.115 ;
        RECT 54.745 110.775 55.245 110.945 ;
        RECT 51.920 109.555 52.090 110.315 ;
        RECT 52.270 109.385 52.600 110.145 ;
        RECT 52.770 109.555 53.040 110.460 ;
        RECT 53.360 109.385 53.690 110.535 ;
        RECT 53.860 110.405 54.870 110.575 ;
        RECT 53.860 109.555 54.030 110.405 ;
        RECT 54.200 109.385 54.530 110.185 ;
        RECT 54.700 109.555 54.870 110.405 ;
        RECT 55.075 110.535 55.245 110.775 ;
        RECT 55.415 110.705 55.795 110.945 ;
        RECT 56.025 110.565 56.435 111.115 ;
        RECT 58.325 110.945 58.650 111.200 ;
        RECT 56.620 110.735 58.650 110.945 ;
        RECT 58.305 110.725 58.650 110.735 ;
        RECT 58.820 110.985 59.060 111.385 ;
        RECT 59.230 111.325 59.400 111.555 ;
        RECT 59.570 111.495 59.760 111.935 ;
        RECT 59.930 111.485 60.880 111.765 ;
        RECT 61.100 111.575 61.450 111.745 ;
        RECT 59.230 111.155 59.760 111.325 ;
        RECT 55.075 110.365 55.790 110.535 ;
        RECT 56.025 110.395 57.750 110.565 ;
        RECT 55.050 109.385 55.290 110.185 ;
        RECT 55.460 109.555 55.790 110.365 ;
        RECT 56.280 109.385 56.450 110.225 ;
        RECT 56.660 109.555 56.910 110.395 ;
        RECT 57.120 109.385 57.290 110.225 ;
        RECT 57.460 109.555 57.750 110.395 ;
        RECT 57.960 109.385 58.130 110.445 ;
        RECT 58.305 110.105 58.475 110.725 ;
        RECT 58.820 110.615 59.360 110.985 ;
        RECT 59.540 110.875 59.760 111.155 ;
        RECT 59.930 110.705 60.100 111.485 ;
        RECT 59.695 110.535 60.100 110.705 ;
        RECT 60.270 110.695 60.620 111.315 ;
        RECT 59.695 110.445 59.865 110.535 ;
        RECT 60.790 110.525 61.000 111.315 ;
        RECT 58.645 110.275 59.865 110.445 ;
        RECT 60.325 110.365 61.000 110.525 ;
        RECT 58.305 109.935 59.105 110.105 ;
        RECT 58.425 109.385 58.755 109.765 ;
        RECT 58.935 109.645 59.105 109.935 ;
        RECT 59.695 109.895 59.865 110.275 ;
        RECT 60.035 110.355 61.000 110.365 ;
        RECT 61.190 111.185 61.450 111.575 ;
        RECT 61.660 111.475 61.990 111.935 ;
        RECT 62.865 111.545 63.720 111.715 ;
        RECT 63.925 111.545 64.420 111.715 ;
        RECT 64.590 111.575 64.920 111.935 ;
        RECT 61.190 110.495 61.360 111.185 ;
        RECT 61.530 110.835 61.700 111.015 ;
        RECT 61.870 111.005 62.660 111.255 ;
        RECT 62.865 110.835 63.035 111.545 ;
        RECT 63.205 111.035 63.560 111.255 ;
        RECT 61.530 110.665 63.220 110.835 ;
        RECT 60.035 110.065 60.495 110.355 ;
        RECT 61.190 110.325 62.690 110.495 ;
        RECT 61.190 110.185 61.360 110.325 ;
        RECT 60.800 110.015 61.360 110.185 ;
        RECT 59.275 109.385 59.525 109.845 ;
        RECT 59.695 109.555 60.565 109.895 ;
        RECT 60.800 109.555 60.970 110.015 ;
        RECT 61.805 109.985 62.880 110.155 ;
        RECT 61.140 109.385 61.510 109.845 ;
        RECT 61.805 109.645 61.975 109.985 ;
        RECT 62.145 109.385 62.475 109.815 ;
        RECT 62.710 109.645 62.880 109.985 ;
        RECT 63.050 109.885 63.220 110.665 ;
        RECT 63.390 110.445 63.560 111.035 ;
        RECT 63.730 110.635 64.080 111.255 ;
        RECT 63.390 110.055 63.855 110.445 ;
        RECT 64.250 110.185 64.420 111.545 ;
        RECT 64.590 110.355 65.050 111.405 ;
        RECT 64.025 110.015 64.420 110.185 ;
        RECT 64.025 109.885 64.195 110.015 ;
        RECT 63.050 109.555 63.730 109.885 ;
        RECT 63.945 109.555 64.195 109.885 ;
        RECT 64.365 109.385 64.615 109.845 ;
        RECT 64.785 109.570 65.110 110.355 ;
        RECT 65.280 109.555 65.450 111.675 ;
        RECT 65.620 111.555 65.950 111.935 ;
        RECT 66.120 111.385 66.375 111.675 ;
        RECT 65.625 111.215 66.375 111.385 ;
        RECT 65.625 110.225 65.855 111.215 ;
        RECT 67.010 111.165 70.520 111.935 ;
        RECT 66.025 110.395 66.375 111.045 ;
        RECT 67.010 110.475 68.700 110.995 ;
        RECT 68.870 110.645 70.520 111.165 ;
        RECT 70.840 111.135 71.170 111.935 ;
        RECT 71.340 111.285 71.510 111.765 ;
        RECT 71.680 111.455 72.010 111.935 ;
        RECT 72.180 111.285 72.350 111.765 ;
        RECT 72.600 111.455 72.840 111.935 ;
        RECT 73.020 111.285 73.190 111.765 ;
        RECT 71.340 111.115 72.350 111.285 ;
        RECT 72.555 111.115 73.190 111.285 ;
        RECT 73.450 111.210 73.740 111.935 ;
        RECT 74.000 111.385 74.170 111.765 ;
        RECT 74.350 111.555 74.680 111.935 ;
        RECT 74.000 111.215 74.665 111.385 ;
        RECT 74.860 111.260 75.120 111.765 ;
        RECT 71.340 110.575 71.835 111.115 ;
        RECT 72.555 110.945 72.725 111.115 ;
        RECT 72.225 110.775 72.725 110.945 ;
        RECT 65.625 110.055 66.375 110.225 ;
        RECT 65.620 109.385 65.950 109.885 ;
        RECT 66.120 109.555 66.375 110.055 ;
        RECT 67.010 109.385 70.520 110.475 ;
        RECT 70.840 109.385 71.170 110.535 ;
        RECT 71.340 110.405 72.350 110.575 ;
        RECT 71.340 109.555 71.510 110.405 ;
        RECT 71.680 109.385 72.010 110.185 ;
        RECT 72.180 109.555 72.350 110.405 ;
        RECT 72.555 110.535 72.725 110.775 ;
        RECT 72.895 110.705 73.275 110.945 ;
        RECT 73.930 110.665 74.260 111.035 ;
        RECT 74.495 110.960 74.665 111.215 ;
        RECT 74.495 110.630 74.780 110.960 ;
        RECT 72.555 110.365 73.270 110.535 ;
        RECT 72.530 109.385 72.770 110.185 ;
        RECT 72.940 109.555 73.270 110.365 ;
        RECT 73.450 109.385 73.740 110.550 ;
        RECT 74.495 110.485 74.665 110.630 ;
        RECT 74.000 110.315 74.665 110.485 ;
        RECT 74.950 110.460 75.120 111.260 ;
        RECT 75.790 111.115 76.020 111.935 ;
        RECT 76.190 111.135 76.520 111.765 ;
        RECT 75.770 110.695 76.100 110.945 ;
        RECT 76.270 110.535 76.520 111.135 ;
        RECT 76.690 111.115 76.900 111.935 ;
        RECT 77.220 111.385 77.390 111.765 ;
        RECT 77.570 111.555 77.900 111.935 ;
        RECT 77.220 111.215 77.885 111.385 ;
        RECT 78.080 111.260 78.340 111.765 ;
        RECT 77.150 110.665 77.480 111.035 ;
        RECT 77.715 110.960 77.885 111.215 ;
        RECT 74.000 109.555 74.170 110.315 ;
        RECT 74.350 109.385 74.680 110.145 ;
        RECT 74.850 109.555 75.120 110.460 ;
        RECT 75.790 109.385 76.020 110.525 ;
        RECT 76.190 109.555 76.520 110.535 ;
        RECT 77.715 110.630 78.000 110.960 ;
        RECT 76.690 109.385 76.900 110.525 ;
        RECT 77.715 110.485 77.885 110.630 ;
        RECT 77.220 110.315 77.885 110.485 ;
        RECT 78.170 110.460 78.340 111.260 ;
        RECT 79.430 111.165 82.940 111.935 ;
        RECT 83.200 111.385 83.370 111.765 ;
        RECT 83.550 111.555 83.880 111.935 ;
        RECT 83.200 111.215 83.865 111.385 ;
        RECT 84.060 111.260 84.320 111.765 ;
        RECT 77.220 109.555 77.390 110.315 ;
        RECT 77.570 109.385 77.900 110.145 ;
        RECT 78.070 109.555 78.340 110.460 ;
        RECT 79.430 110.475 81.120 110.995 ;
        RECT 81.290 110.645 82.940 111.165 ;
        RECT 83.130 110.665 83.460 111.035 ;
        RECT 83.695 110.960 83.865 111.215 ;
        RECT 83.695 110.630 83.980 110.960 ;
        RECT 83.695 110.485 83.865 110.630 ;
        RECT 79.430 109.385 82.940 110.475 ;
        RECT 83.200 110.315 83.865 110.485 ;
        RECT 84.150 110.460 84.320 111.260 ;
        RECT 84.490 111.185 85.700 111.935 ;
        RECT 83.200 109.555 83.370 110.315 ;
        RECT 83.550 109.385 83.880 110.145 ;
        RECT 84.050 109.555 84.320 110.460 ;
        RECT 84.490 110.475 85.010 111.015 ;
        RECT 85.180 110.645 85.700 111.185 ;
        RECT 85.870 111.165 89.380 111.935 ;
        RECT 89.640 111.385 89.810 111.765 ;
        RECT 89.990 111.555 90.320 111.935 ;
        RECT 89.640 111.215 90.305 111.385 ;
        RECT 90.500 111.260 90.760 111.765 ;
        RECT 85.870 110.475 87.560 110.995 ;
        RECT 87.730 110.645 89.380 111.165 ;
        RECT 89.570 110.665 89.900 111.035 ;
        RECT 90.135 110.960 90.305 111.215 ;
        RECT 90.135 110.630 90.420 110.960 ;
        RECT 90.135 110.485 90.305 110.630 ;
        RECT 84.490 109.385 85.700 110.475 ;
        RECT 85.870 109.385 89.380 110.475 ;
        RECT 89.640 110.315 90.305 110.485 ;
        RECT 90.590 110.460 90.760 111.260 ;
        RECT 91.205 111.125 91.450 111.730 ;
        RECT 91.670 111.400 92.180 111.935 ;
        RECT 89.640 109.555 89.810 110.315 ;
        RECT 89.990 109.385 90.320 110.145 ;
        RECT 90.490 109.555 90.760 110.460 ;
        RECT 90.930 110.955 92.160 111.125 ;
        RECT 90.930 110.145 91.270 110.955 ;
        RECT 91.440 110.390 92.190 110.580 ;
        RECT 90.930 109.735 91.445 110.145 ;
        RECT 91.680 109.385 91.850 110.145 ;
        RECT 92.020 109.725 92.190 110.390 ;
        RECT 92.360 110.405 92.550 111.765 ;
        RECT 92.720 111.255 92.995 111.765 ;
        RECT 93.185 111.400 93.715 111.765 ;
        RECT 94.140 111.535 94.470 111.935 ;
        RECT 93.540 111.365 93.715 111.400 ;
        RECT 92.720 111.085 93.000 111.255 ;
        RECT 92.720 110.605 92.995 111.085 ;
        RECT 93.200 110.405 93.370 111.205 ;
        RECT 92.360 110.235 93.370 110.405 ;
        RECT 93.540 111.195 94.470 111.365 ;
        RECT 94.640 111.195 94.895 111.765 ;
        RECT 93.540 110.065 93.710 111.195 ;
        RECT 94.300 111.025 94.470 111.195 ;
        RECT 92.585 109.895 93.710 110.065 ;
        RECT 93.880 110.695 94.075 111.025 ;
        RECT 94.300 110.695 94.555 111.025 ;
        RECT 93.880 109.725 94.050 110.695 ;
        RECT 94.725 110.525 94.895 111.195 ;
        RECT 95.530 111.165 97.200 111.935 ;
        RECT 92.020 109.555 94.050 109.725 ;
        RECT 94.220 109.385 94.390 110.525 ;
        RECT 94.560 109.555 94.895 110.525 ;
        RECT 95.530 110.475 96.280 110.995 ;
        RECT 96.450 110.645 97.200 111.165 ;
        RECT 97.370 111.260 97.630 111.765 ;
        RECT 97.810 111.555 98.140 111.935 ;
        RECT 98.320 111.385 98.490 111.765 ;
        RECT 95.530 109.385 97.200 110.475 ;
        RECT 97.370 110.460 97.540 111.260 ;
        RECT 97.825 111.215 98.490 111.385 ;
        RECT 97.825 110.960 97.995 111.215 ;
        RECT 99.210 111.210 99.500 111.935 ;
        RECT 99.670 111.185 100.880 111.935 ;
        RECT 101.140 111.385 101.310 111.765 ;
        RECT 101.490 111.555 101.820 111.935 ;
        RECT 101.140 111.215 101.805 111.385 ;
        RECT 102.000 111.260 102.260 111.765 ;
        RECT 97.710 110.630 97.995 110.960 ;
        RECT 98.230 110.665 98.560 111.035 ;
        RECT 97.825 110.485 97.995 110.630 ;
        RECT 97.370 109.555 97.640 110.460 ;
        RECT 97.825 110.315 98.490 110.485 ;
        RECT 97.810 109.385 98.140 110.145 ;
        RECT 98.320 109.555 98.490 110.315 ;
        RECT 99.210 109.385 99.500 110.550 ;
        RECT 99.670 110.475 100.190 111.015 ;
        RECT 100.360 110.645 100.880 111.185 ;
        RECT 101.070 110.665 101.400 111.035 ;
        RECT 101.635 110.960 101.805 111.215 ;
        RECT 101.635 110.630 101.920 110.960 ;
        RECT 101.635 110.485 101.805 110.630 ;
        RECT 99.670 109.385 100.880 110.475 ;
        RECT 101.140 110.315 101.805 110.485 ;
        RECT 102.090 110.460 102.260 111.260 ;
        RECT 102.470 111.115 102.700 111.935 ;
        RECT 102.870 111.135 103.200 111.765 ;
        RECT 102.450 110.695 102.780 110.945 ;
        RECT 102.950 110.535 103.200 111.135 ;
        RECT 103.370 111.115 103.580 111.935 ;
        RECT 103.850 111.115 104.080 111.935 ;
        RECT 104.250 111.135 104.580 111.765 ;
        RECT 103.830 110.695 104.160 110.945 ;
        RECT 104.330 110.535 104.580 111.135 ;
        RECT 104.750 111.115 104.960 111.935 ;
        RECT 105.190 111.260 105.450 111.765 ;
        RECT 105.630 111.555 105.960 111.935 ;
        RECT 106.140 111.385 106.310 111.765 ;
        RECT 101.140 109.555 101.310 110.315 ;
        RECT 101.490 109.385 101.820 110.145 ;
        RECT 101.990 109.555 102.260 110.460 ;
        RECT 102.470 109.385 102.700 110.525 ;
        RECT 102.870 109.555 103.200 110.535 ;
        RECT 103.370 109.385 103.580 110.525 ;
        RECT 103.850 109.385 104.080 110.525 ;
        RECT 104.250 109.555 104.580 110.535 ;
        RECT 104.750 109.385 104.960 110.525 ;
        RECT 105.190 110.460 105.360 111.260 ;
        RECT 105.645 111.215 106.310 111.385 ;
        RECT 106.660 111.385 106.830 111.765 ;
        RECT 107.010 111.555 107.340 111.935 ;
        RECT 106.660 111.215 107.325 111.385 ;
        RECT 107.520 111.260 107.780 111.765 ;
        RECT 105.645 110.960 105.815 111.215 ;
        RECT 105.530 110.630 105.815 110.960 ;
        RECT 106.050 110.665 106.380 111.035 ;
        RECT 106.590 110.665 106.920 111.035 ;
        RECT 107.155 110.960 107.325 111.215 ;
        RECT 105.645 110.485 105.815 110.630 ;
        RECT 107.155 110.630 107.440 110.960 ;
        RECT 107.155 110.485 107.325 110.630 ;
        RECT 105.190 109.555 105.460 110.460 ;
        RECT 105.645 110.315 106.310 110.485 ;
        RECT 105.630 109.385 105.960 110.145 ;
        RECT 106.140 109.555 106.310 110.315 ;
        RECT 106.660 110.315 107.325 110.485 ;
        RECT 107.610 110.460 107.780 111.260 ;
        RECT 107.950 111.165 109.620 111.935 ;
        RECT 106.660 109.555 106.830 110.315 ;
        RECT 107.010 109.385 107.340 110.145 ;
        RECT 107.510 109.555 107.780 110.460 ;
        RECT 107.950 110.475 108.700 110.995 ;
        RECT 108.870 110.645 109.620 111.165 ;
        RECT 109.790 111.260 110.050 111.765 ;
        RECT 110.230 111.555 110.560 111.935 ;
        RECT 110.740 111.385 110.910 111.765 ;
        RECT 107.950 109.385 109.620 110.475 ;
        RECT 109.790 110.460 109.970 111.260 ;
        RECT 110.245 111.215 110.910 111.385 ;
        RECT 110.245 110.960 110.415 111.215 ;
        RECT 111.170 111.185 112.380 111.935 ;
        RECT 110.140 110.630 110.415 110.960 ;
        RECT 110.640 110.665 110.980 111.035 ;
        RECT 110.245 110.485 110.415 110.630 ;
        RECT 109.790 109.555 110.060 110.460 ;
        RECT 110.245 110.315 110.920 110.485 ;
        RECT 110.230 109.385 110.560 110.145 ;
        RECT 110.740 109.555 110.920 110.315 ;
        RECT 111.170 110.475 111.690 111.015 ;
        RECT 111.860 110.645 112.380 111.185 ;
        RECT 111.170 109.385 112.380 110.475 ;
        RECT 18.165 109.215 112.465 109.385 ;
        RECT 18.250 108.125 19.460 109.215 ;
        RECT 18.250 107.415 18.770 107.955 ;
        RECT 18.940 107.585 19.460 108.125 ;
        RECT 19.630 108.125 23.140 109.215 ;
        RECT 23.620 108.375 23.790 109.215 ;
        RECT 24.000 108.205 24.250 109.045 ;
        RECT 24.460 108.375 24.630 109.215 ;
        RECT 24.800 108.205 25.090 109.045 ;
        RECT 19.630 107.605 21.320 108.125 ;
        RECT 23.365 108.035 25.090 108.205 ;
        RECT 25.300 108.155 25.470 109.215 ;
        RECT 25.765 108.835 26.095 109.215 ;
        RECT 26.275 108.665 26.445 108.955 ;
        RECT 26.615 108.755 26.865 109.215 ;
        RECT 25.645 108.495 26.445 108.665 ;
        RECT 27.035 108.705 27.905 109.045 ;
        RECT 21.490 107.435 23.140 107.955 ;
        RECT 18.250 106.665 19.460 107.415 ;
        RECT 19.630 106.665 23.140 107.435 ;
        RECT 23.365 107.485 23.775 108.035 ;
        RECT 25.645 107.875 25.815 108.495 ;
        RECT 27.035 108.325 27.205 108.705 ;
        RECT 28.140 108.585 28.310 109.045 ;
        RECT 28.480 108.755 28.850 109.215 ;
        RECT 29.145 108.615 29.315 108.955 ;
        RECT 29.485 108.785 29.815 109.215 ;
        RECT 30.050 108.615 30.220 108.955 ;
        RECT 25.985 108.155 27.205 108.325 ;
        RECT 27.375 108.245 27.835 108.535 ;
        RECT 28.140 108.415 28.700 108.585 ;
        RECT 29.145 108.445 30.220 108.615 ;
        RECT 30.390 108.715 31.070 109.045 ;
        RECT 31.285 108.715 31.535 109.045 ;
        RECT 31.705 108.755 31.955 109.215 ;
        RECT 28.530 108.275 28.700 108.415 ;
        RECT 27.375 108.235 28.340 108.245 ;
        RECT 27.035 108.065 27.205 108.155 ;
        RECT 27.665 108.075 28.340 108.235 ;
        RECT 25.645 107.865 25.990 107.875 ;
        RECT 23.960 107.655 25.990 107.865 ;
        RECT 23.365 107.315 25.130 107.485 ;
        RECT 23.620 106.665 23.790 107.135 ;
        RECT 23.960 106.835 24.290 107.315 ;
        RECT 24.460 106.665 24.630 107.135 ;
        RECT 24.800 106.835 25.130 107.315 ;
        RECT 25.300 106.665 25.470 107.475 ;
        RECT 25.665 107.400 25.990 107.655 ;
        RECT 25.670 107.045 25.990 107.400 ;
        RECT 26.160 107.615 26.700 107.985 ;
        RECT 27.035 107.895 27.440 108.065 ;
        RECT 26.160 107.215 26.400 107.615 ;
        RECT 26.880 107.445 27.100 107.725 ;
        RECT 26.570 107.275 27.100 107.445 ;
        RECT 26.570 107.045 26.740 107.275 ;
        RECT 27.270 107.115 27.440 107.895 ;
        RECT 27.610 107.285 27.960 107.905 ;
        RECT 28.130 107.285 28.340 108.075 ;
        RECT 28.530 108.105 30.030 108.275 ;
        RECT 28.530 107.415 28.700 108.105 ;
        RECT 30.390 107.935 30.560 108.715 ;
        RECT 31.365 108.585 31.535 108.715 ;
        RECT 28.870 107.765 30.560 107.935 ;
        RECT 30.730 108.155 31.195 108.545 ;
        RECT 31.365 108.415 31.760 108.585 ;
        RECT 28.870 107.585 29.040 107.765 ;
        RECT 25.670 106.875 26.740 107.045 ;
        RECT 26.910 106.665 27.100 107.105 ;
        RECT 27.270 106.835 28.220 107.115 ;
        RECT 28.530 107.025 28.790 107.415 ;
        RECT 29.210 107.345 30.000 107.595 ;
        RECT 28.440 106.855 28.790 107.025 ;
        RECT 29.000 106.665 29.330 107.125 ;
        RECT 30.205 107.055 30.375 107.765 ;
        RECT 30.730 107.565 30.900 108.155 ;
        RECT 30.545 107.345 30.900 107.565 ;
        RECT 31.070 107.345 31.420 107.965 ;
        RECT 31.590 107.055 31.760 108.415 ;
        RECT 32.125 108.245 32.450 109.030 ;
        RECT 31.930 107.195 32.390 108.245 ;
        RECT 30.205 106.885 31.060 107.055 ;
        RECT 31.265 106.885 31.760 107.055 ;
        RECT 31.930 106.665 32.260 107.025 ;
        RECT 32.620 106.925 32.790 109.045 ;
        RECT 32.960 108.715 33.290 109.215 ;
        RECT 33.460 108.545 33.715 109.045 ;
        RECT 32.965 108.375 33.715 108.545 ;
        RECT 32.965 107.385 33.195 108.375 ;
        RECT 33.365 107.555 33.715 108.205 ;
        RECT 34.810 108.050 35.100 109.215 ;
        RECT 35.730 108.140 36.000 109.045 ;
        RECT 36.170 108.455 36.500 109.215 ;
        RECT 36.680 108.285 36.850 109.045 ;
        RECT 32.965 107.215 33.715 107.385 ;
        RECT 32.960 106.665 33.290 107.045 ;
        RECT 33.460 106.925 33.715 107.215 ;
        RECT 34.810 106.665 35.100 107.390 ;
        RECT 35.730 107.340 35.900 108.140 ;
        RECT 36.185 108.115 36.850 108.285 ;
        RECT 36.185 107.970 36.355 108.115 ;
        RECT 37.630 108.075 37.840 109.215 ;
        RECT 36.070 107.640 36.355 107.970 ;
        RECT 38.010 108.065 38.340 109.045 ;
        RECT 38.510 108.075 38.740 109.215 ;
        RECT 39.450 108.075 39.680 109.215 ;
        RECT 39.850 108.065 40.180 109.045 ;
        RECT 40.350 108.075 40.560 109.215 ;
        RECT 40.790 108.140 41.060 109.045 ;
        RECT 41.230 108.455 41.560 109.215 ;
        RECT 41.740 108.285 41.910 109.045 ;
        RECT 36.185 107.385 36.355 107.640 ;
        RECT 36.590 107.565 36.920 107.935 ;
        RECT 35.730 106.835 35.990 107.340 ;
        RECT 36.185 107.215 36.850 107.385 ;
        RECT 36.170 106.665 36.500 107.045 ;
        RECT 36.680 106.835 36.850 107.215 ;
        RECT 37.630 106.665 37.840 107.485 ;
        RECT 38.010 107.465 38.260 108.065 ;
        RECT 38.430 107.655 38.760 107.905 ;
        RECT 39.430 107.655 39.760 107.905 ;
        RECT 38.010 106.835 38.340 107.465 ;
        RECT 38.510 106.665 38.740 107.485 ;
        RECT 39.450 106.665 39.680 107.485 ;
        RECT 39.930 107.465 40.180 108.065 ;
        RECT 39.850 106.835 40.180 107.465 ;
        RECT 40.350 106.665 40.560 107.485 ;
        RECT 40.790 107.340 40.960 108.140 ;
        RECT 41.245 108.115 41.910 108.285 ;
        RECT 42.630 108.140 42.900 109.045 ;
        RECT 43.070 108.455 43.400 109.215 ;
        RECT 43.580 108.285 43.750 109.045 ;
        RECT 41.245 107.970 41.415 108.115 ;
        RECT 41.130 107.640 41.415 107.970 ;
        RECT 41.245 107.385 41.415 107.640 ;
        RECT 41.650 107.565 41.980 107.935 ;
        RECT 40.790 106.835 41.050 107.340 ;
        RECT 41.245 107.215 41.910 107.385 ;
        RECT 41.230 106.665 41.560 107.045 ;
        RECT 41.740 106.835 41.910 107.215 ;
        RECT 42.630 107.340 42.800 108.140 ;
        RECT 43.085 108.115 43.750 108.285 ;
        RECT 44.010 108.140 44.280 109.045 ;
        RECT 44.450 108.455 44.780 109.215 ;
        RECT 44.960 108.285 45.130 109.045 ;
        RECT 43.085 107.970 43.255 108.115 ;
        RECT 42.970 107.640 43.255 107.970 ;
        RECT 43.085 107.385 43.255 107.640 ;
        RECT 43.490 107.565 43.820 107.935 ;
        RECT 42.630 106.835 42.890 107.340 ;
        RECT 43.085 107.215 43.750 107.385 ;
        RECT 43.070 106.665 43.400 107.045 ;
        RECT 43.580 106.835 43.750 107.215 ;
        RECT 44.010 107.340 44.180 108.140 ;
        RECT 44.465 108.115 45.130 108.285 ;
        RECT 45.480 108.285 45.650 109.045 ;
        RECT 45.830 108.455 46.160 109.215 ;
        RECT 45.480 108.115 46.145 108.285 ;
        RECT 46.330 108.140 46.600 109.045 ;
        RECT 47.080 108.375 47.250 109.215 ;
        RECT 47.460 108.205 47.710 109.045 ;
        RECT 47.920 108.375 48.090 109.215 ;
        RECT 48.260 108.205 48.550 109.045 ;
        RECT 44.465 107.970 44.635 108.115 ;
        RECT 44.350 107.640 44.635 107.970 ;
        RECT 45.975 107.970 46.145 108.115 ;
        RECT 44.465 107.385 44.635 107.640 ;
        RECT 44.870 107.565 45.200 107.935 ;
        RECT 45.410 107.565 45.740 107.935 ;
        RECT 45.975 107.640 46.260 107.970 ;
        RECT 45.975 107.385 46.145 107.640 ;
        RECT 44.010 106.835 44.270 107.340 ;
        RECT 44.465 107.215 45.130 107.385 ;
        RECT 44.450 106.665 44.780 107.045 ;
        RECT 44.960 106.835 45.130 107.215 ;
        RECT 45.480 107.215 46.145 107.385 ;
        RECT 46.430 107.340 46.600 108.140 ;
        RECT 45.480 106.835 45.650 107.215 ;
        RECT 45.830 106.665 46.160 107.045 ;
        RECT 46.340 106.835 46.600 107.340 ;
        RECT 46.825 108.035 48.550 108.205 ;
        RECT 48.760 108.155 48.930 109.215 ;
        RECT 49.225 108.835 49.555 109.215 ;
        RECT 49.735 108.665 49.905 108.955 ;
        RECT 50.075 108.755 50.325 109.215 ;
        RECT 49.105 108.495 49.905 108.665 ;
        RECT 50.495 108.705 51.365 109.045 ;
        RECT 46.825 107.485 47.235 108.035 ;
        RECT 49.105 107.875 49.275 108.495 ;
        RECT 50.495 108.325 50.665 108.705 ;
        RECT 51.600 108.585 51.770 109.045 ;
        RECT 51.940 108.755 52.310 109.215 ;
        RECT 52.605 108.615 52.775 108.955 ;
        RECT 52.945 108.785 53.275 109.215 ;
        RECT 53.510 108.615 53.680 108.955 ;
        RECT 49.445 108.155 50.665 108.325 ;
        RECT 50.835 108.245 51.295 108.535 ;
        RECT 51.600 108.415 52.160 108.585 ;
        RECT 52.605 108.445 53.680 108.615 ;
        RECT 53.850 108.715 54.530 109.045 ;
        RECT 54.745 108.715 54.995 109.045 ;
        RECT 55.165 108.755 55.415 109.215 ;
        RECT 51.990 108.275 52.160 108.415 ;
        RECT 50.835 108.235 51.800 108.245 ;
        RECT 50.495 108.065 50.665 108.155 ;
        RECT 51.125 108.075 51.800 108.235 ;
        RECT 49.105 107.865 49.450 107.875 ;
        RECT 47.420 107.655 49.450 107.865 ;
        RECT 46.825 107.315 48.590 107.485 ;
        RECT 47.080 106.665 47.250 107.135 ;
        RECT 47.420 106.835 47.750 107.315 ;
        RECT 47.920 106.665 48.090 107.135 ;
        RECT 48.260 106.835 48.590 107.315 ;
        RECT 48.760 106.665 48.930 107.475 ;
        RECT 49.125 107.400 49.450 107.655 ;
        RECT 49.130 107.045 49.450 107.400 ;
        RECT 49.620 107.615 50.160 107.985 ;
        RECT 50.495 107.895 50.900 108.065 ;
        RECT 49.620 107.215 49.860 107.615 ;
        RECT 50.340 107.445 50.560 107.725 ;
        RECT 50.030 107.275 50.560 107.445 ;
        RECT 50.030 107.045 50.200 107.275 ;
        RECT 50.730 107.115 50.900 107.895 ;
        RECT 51.070 107.285 51.420 107.905 ;
        RECT 51.590 107.285 51.800 108.075 ;
        RECT 51.990 108.105 53.490 108.275 ;
        RECT 51.990 107.415 52.160 108.105 ;
        RECT 53.850 107.935 54.020 108.715 ;
        RECT 54.825 108.585 54.995 108.715 ;
        RECT 52.330 107.765 54.020 107.935 ;
        RECT 54.190 108.155 54.655 108.545 ;
        RECT 54.825 108.415 55.220 108.585 ;
        RECT 52.330 107.585 52.500 107.765 ;
        RECT 49.130 106.875 50.200 107.045 ;
        RECT 50.370 106.665 50.560 107.105 ;
        RECT 50.730 106.835 51.680 107.115 ;
        RECT 51.990 107.025 52.250 107.415 ;
        RECT 52.670 107.345 53.460 107.595 ;
        RECT 51.900 106.855 52.250 107.025 ;
        RECT 52.460 106.665 52.790 107.125 ;
        RECT 53.665 107.055 53.835 107.765 ;
        RECT 54.190 107.565 54.360 108.155 ;
        RECT 54.005 107.345 54.360 107.565 ;
        RECT 54.530 107.345 54.880 107.965 ;
        RECT 55.050 107.055 55.220 108.415 ;
        RECT 55.585 108.245 55.910 109.030 ;
        RECT 55.390 107.195 55.850 108.245 ;
        RECT 53.665 106.885 54.520 107.055 ;
        RECT 54.725 106.885 55.220 107.055 ;
        RECT 55.390 106.665 55.720 107.025 ;
        RECT 56.080 106.925 56.250 109.045 ;
        RECT 56.420 108.715 56.750 109.215 ;
        RECT 56.920 108.545 57.175 109.045 ;
        RECT 56.425 108.375 57.175 108.545 ;
        RECT 56.425 107.385 56.655 108.375 ;
        RECT 57.820 108.235 58.150 109.045 ;
        RECT 58.320 108.415 58.560 109.215 ;
        RECT 56.825 107.555 57.175 108.205 ;
        RECT 57.820 108.065 58.535 108.235 ;
        RECT 57.815 107.655 58.195 107.895 ;
        RECT 58.365 107.825 58.535 108.065 ;
        RECT 58.740 108.195 58.910 109.045 ;
        RECT 59.080 108.415 59.410 109.215 ;
        RECT 59.580 108.195 59.750 109.045 ;
        RECT 58.740 108.025 59.750 108.195 ;
        RECT 59.920 108.065 60.250 109.215 ;
        RECT 60.570 108.050 60.860 109.215 ;
        RECT 61.070 108.075 61.300 109.215 ;
        RECT 61.470 108.065 61.800 109.045 ;
        RECT 61.970 108.075 62.180 109.215 ;
        RECT 62.500 108.285 62.670 109.045 ;
        RECT 62.850 108.455 63.180 109.215 ;
        RECT 62.500 108.115 63.165 108.285 ;
        RECT 63.350 108.140 63.620 109.045 ;
        RECT 59.255 107.855 59.750 108.025 ;
        RECT 58.365 107.655 58.865 107.825 ;
        RECT 59.250 107.685 59.750 107.855 ;
        RECT 58.365 107.485 58.535 107.655 ;
        RECT 59.255 107.485 59.750 107.685 ;
        RECT 61.050 107.655 61.380 107.905 ;
        RECT 56.425 107.215 57.175 107.385 ;
        RECT 56.420 106.665 56.750 107.045 ;
        RECT 56.920 106.925 57.175 107.215 ;
        RECT 57.900 107.315 58.535 107.485 ;
        RECT 58.740 107.315 59.750 107.485 ;
        RECT 57.900 106.835 58.070 107.315 ;
        RECT 58.250 106.665 58.490 107.145 ;
        RECT 58.740 106.835 58.910 107.315 ;
        RECT 59.080 106.665 59.410 107.145 ;
        RECT 59.580 106.835 59.750 107.315 ;
        RECT 59.920 106.665 60.250 107.465 ;
        RECT 60.570 106.665 60.860 107.390 ;
        RECT 61.070 106.665 61.300 107.485 ;
        RECT 61.550 107.465 61.800 108.065 ;
        RECT 62.995 107.970 63.165 108.115 ;
        RECT 62.430 107.565 62.760 107.935 ;
        RECT 62.995 107.640 63.280 107.970 ;
        RECT 61.470 106.835 61.800 107.465 ;
        RECT 61.970 106.665 62.180 107.485 ;
        RECT 62.995 107.385 63.165 107.640 ;
        RECT 62.500 107.215 63.165 107.385 ;
        RECT 63.450 107.340 63.620 108.140 ;
        RECT 63.880 108.285 64.050 109.045 ;
        RECT 64.230 108.455 64.560 109.215 ;
        RECT 63.880 108.115 64.545 108.285 ;
        RECT 64.730 108.140 65.000 109.045 ;
        RECT 65.480 108.375 65.650 109.215 ;
        RECT 65.860 108.205 66.110 109.045 ;
        RECT 66.320 108.375 66.490 109.215 ;
        RECT 66.660 108.205 66.950 109.045 ;
        RECT 64.375 107.970 64.545 108.115 ;
        RECT 63.810 107.565 64.140 107.935 ;
        RECT 64.375 107.640 64.660 107.970 ;
        RECT 64.375 107.385 64.545 107.640 ;
        RECT 62.500 106.835 62.670 107.215 ;
        RECT 62.850 106.665 63.180 107.045 ;
        RECT 63.360 106.835 63.620 107.340 ;
        RECT 63.880 107.215 64.545 107.385 ;
        RECT 64.830 107.340 65.000 108.140 ;
        RECT 63.880 106.835 64.050 107.215 ;
        RECT 64.230 106.665 64.560 107.045 ;
        RECT 64.740 106.835 65.000 107.340 ;
        RECT 65.225 108.035 66.950 108.205 ;
        RECT 67.160 108.155 67.330 109.215 ;
        RECT 67.625 108.835 67.955 109.215 ;
        RECT 68.135 108.665 68.305 108.955 ;
        RECT 68.475 108.755 68.725 109.215 ;
        RECT 67.505 108.495 68.305 108.665 ;
        RECT 68.895 108.705 69.765 109.045 ;
        RECT 65.225 107.485 65.635 108.035 ;
        RECT 67.505 107.875 67.675 108.495 ;
        RECT 68.895 108.325 69.065 108.705 ;
        RECT 70.000 108.585 70.170 109.045 ;
        RECT 70.340 108.755 70.710 109.215 ;
        RECT 71.005 108.615 71.175 108.955 ;
        RECT 71.345 108.785 71.675 109.215 ;
        RECT 71.910 108.615 72.080 108.955 ;
        RECT 67.845 108.155 69.065 108.325 ;
        RECT 69.235 108.245 69.695 108.535 ;
        RECT 70.000 108.415 70.560 108.585 ;
        RECT 71.005 108.445 72.080 108.615 ;
        RECT 72.250 108.715 72.930 109.045 ;
        RECT 73.145 108.715 73.395 109.045 ;
        RECT 73.565 108.755 73.815 109.215 ;
        RECT 70.390 108.275 70.560 108.415 ;
        RECT 69.235 108.235 70.200 108.245 ;
        RECT 68.895 108.065 69.065 108.155 ;
        RECT 69.525 108.075 70.200 108.235 ;
        RECT 67.505 107.865 67.850 107.875 ;
        RECT 65.820 107.655 67.850 107.865 ;
        RECT 65.225 107.315 66.990 107.485 ;
        RECT 65.480 106.665 65.650 107.135 ;
        RECT 65.820 106.835 66.150 107.315 ;
        RECT 66.320 106.665 66.490 107.135 ;
        RECT 66.660 106.835 66.990 107.315 ;
        RECT 67.160 106.665 67.330 107.475 ;
        RECT 67.525 107.400 67.850 107.655 ;
        RECT 67.530 107.045 67.850 107.400 ;
        RECT 68.020 107.615 68.560 107.985 ;
        RECT 68.895 107.895 69.300 108.065 ;
        RECT 68.020 107.215 68.260 107.615 ;
        RECT 68.740 107.445 68.960 107.725 ;
        RECT 68.430 107.275 68.960 107.445 ;
        RECT 68.430 107.045 68.600 107.275 ;
        RECT 69.130 107.115 69.300 107.895 ;
        RECT 69.470 107.285 69.820 107.905 ;
        RECT 69.990 107.285 70.200 108.075 ;
        RECT 70.390 108.105 71.890 108.275 ;
        RECT 70.390 107.415 70.560 108.105 ;
        RECT 72.250 107.935 72.420 108.715 ;
        RECT 73.225 108.585 73.395 108.715 ;
        RECT 70.730 107.765 72.420 107.935 ;
        RECT 72.590 108.155 73.055 108.545 ;
        RECT 73.225 108.415 73.620 108.585 ;
        RECT 70.730 107.585 70.900 107.765 ;
        RECT 67.530 106.875 68.600 107.045 ;
        RECT 68.770 106.665 68.960 107.105 ;
        RECT 69.130 106.835 70.080 107.115 ;
        RECT 70.390 107.025 70.650 107.415 ;
        RECT 71.070 107.345 71.860 107.595 ;
        RECT 70.300 106.855 70.650 107.025 ;
        RECT 70.860 106.665 71.190 107.125 ;
        RECT 72.065 107.055 72.235 107.765 ;
        RECT 72.590 107.565 72.760 108.155 ;
        RECT 72.405 107.345 72.760 107.565 ;
        RECT 72.930 107.345 73.280 107.965 ;
        RECT 73.450 107.055 73.620 108.415 ;
        RECT 73.985 108.245 74.310 109.030 ;
        RECT 73.790 107.195 74.250 108.245 ;
        RECT 72.065 106.885 72.920 107.055 ;
        RECT 73.125 106.885 73.620 107.055 ;
        RECT 73.790 106.665 74.120 107.025 ;
        RECT 74.480 106.925 74.650 109.045 ;
        RECT 74.820 108.715 75.150 109.215 ;
        RECT 75.320 108.545 75.575 109.045 ;
        RECT 74.825 108.375 75.575 108.545 ;
        RECT 76.060 108.375 76.230 109.215 ;
        RECT 74.825 107.385 75.055 108.375 ;
        RECT 76.440 108.205 76.690 109.045 ;
        RECT 76.900 108.375 77.070 109.215 ;
        RECT 77.240 108.205 77.530 109.045 ;
        RECT 75.225 107.555 75.575 108.205 ;
        RECT 75.805 108.035 77.530 108.205 ;
        RECT 77.740 108.155 77.910 109.215 ;
        RECT 78.205 108.835 78.535 109.215 ;
        RECT 78.715 108.665 78.885 108.955 ;
        RECT 79.055 108.755 79.305 109.215 ;
        RECT 78.085 108.495 78.885 108.665 ;
        RECT 79.475 108.705 80.345 109.045 ;
        RECT 75.805 107.485 76.215 108.035 ;
        RECT 78.085 107.875 78.255 108.495 ;
        RECT 79.475 108.325 79.645 108.705 ;
        RECT 80.580 108.585 80.750 109.045 ;
        RECT 80.920 108.755 81.290 109.215 ;
        RECT 81.585 108.615 81.755 108.955 ;
        RECT 81.925 108.785 82.255 109.215 ;
        RECT 82.490 108.615 82.660 108.955 ;
        RECT 78.425 108.155 79.645 108.325 ;
        RECT 79.815 108.245 80.275 108.535 ;
        RECT 80.580 108.415 81.140 108.585 ;
        RECT 81.585 108.445 82.660 108.615 ;
        RECT 82.830 108.715 83.510 109.045 ;
        RECT 83.725 108.715 83.975 109.045 ;
        RECT 84.145 108.755 84.395 109.215 ;
        RECT 80.970 108.275 81.140 108.415 ;
        RECT 79.815 108.235 80.780 108.245 ;
        RECT 79.475 108.065 79.645 108.155 ;
        RECT 80.105 108.075 80.780 108.235 ;
        RECT 78.085 107.865 78.430 107.875 ;
        RECT 76.400 107.655 78.430 107.865 ;
        RECT 74.825 107.215 75.575 107.385 ;
        RECT 75.805 107.315 77.570 107.485 ;
        RECT 74.820 106.665 75.150 107.045 ;
        RECT 75.320 106.925 75.575 107.215 ;
        RECT 76.060 106.665 76.230 107.135 ;
        RECT 76.400 106.835 76.730 107.315 ;
        RECT 76.900 106.665 77.070 107.135 ;
        RECT 77.240 106.835 77.570 107.315 ;
        RECT 77.740 106.665 77.910 107.475 ;
        RECT 78.105 107.400 78.430 107.655 ;
        RECT 78.110 107.045 78.430 107.400 ;
        RECT 78.600 107.615 79.140 107.985 ;
        RECT 79.475 107.895 79.880 108.065 ;
        RECT 78.600 107.215 78.840 107.615 ;
        RECT 79.320 107.445 79.540 107.725 ;
        RECT 79.010 107.275 79.540 107.445 ;
        RECT 79.010 107.045 79.180 107.275 ;
        RECT 79.710 107.115 79.880 107.895 ;
        RECT 80.050 107.285 80.400 107.905 ;
        RECT 80.570 107.285 80.780 108.075 ;
        RECT 80.970 108.105 82.470 108.275 ;
        RECT 80.970 107.415 81.140 108.105 ;
        RECT 82.830 107.935 83.000 108.715 ;
        RECT 83.805 108.585 83.975 108.715 ;
        RECT 81.310 107.765 83.000 107.935 ;
        RECT 83.170 108.155 83.635 108.545 ;
        RECT 83.805 108.415 84.200 108.585 ;
        RECT 81.310 107.585 81.480 107.765 ;
        RECT 78.110 106.875 79.180 107.045 ;
        RECT 79.350 106.665 79.540 107.105 ;
        RECT 79.710 106.835 80.660 107.115 ;
        RECT 80.970 107.025 81.230 107.415 ;
        RECT 81.650 107.345 82.440 107.595 ;
        RECT 80.880 106.855 81.230 107.025 ;
        RECT 81.440 106.665 81.770 107.125 ;
        RECT 82.645 107.055 82.815 107.765 ;
        RECT 83.170 107.565 83.340 108.155 ;
        RECT 82.985 107.345 83.340 107.565 ;
        RECT 83.510 107.345 83.860 107.965 ;
        RECT 84.030 107.055 84.200 108.415 ;
        RECT 84.565 108.245 84.890 109.030 ;
        RECT 84.370 107.195 84.830 108.245 ;
        RECT 82.645 106.885 83.500 107.055 ;
        RECT 83.705 106.885 84.200 107.055 ;
        RECT 84.370 106.665 84.700 107.025 ;
        RECT 85.060 106.925 85.230 109.045 ;
        RECT 85.400 108.715 85.730 109.215 ;
        RECT 85.900 108.545 86.155 109.045 ;
        RECT 85.405 108.375 86.155 108.545 ;
        RECT 85.405 107.385 85.635 108.375 ;
        RECT 85.805 107.555 86.155 108.205 ;
        RECT 86.330 108.050 86.620 109.215 ;
        RECT 88.020 108.375 88.190 109.215 ;
        RECT 88.400 108.205 88.650 109.045 ;
        RECT 88.860 108.375 89.030 109.215 ;
        RECT 89.200 108.205 89.490 109.045 ;
        RECT 87.765 108.035 89.490 108.205 ;
        RECT 89.700 108.155 89.870 109.215 ;
        RECT 90.165 108.835 90.495 109.215 ;
        RECT 90.675 108.665 90.845 108.955 ;
        RECT 91.015 108.755 91.265 109.215 ;
        RECT 90.045 108.495 90.845 108.665 ;
        RECT 91.435 108.705 92.305 109.045 ;
        RECT 87.765 107.485 88.175 108.035 ;
        RECT 90.045 107.875 90.215 108.495 ;
        RECT 91.435 108.325 91.605 108.705 ;
        RECT 92.540 108.585 92.710 109.045 ;
        RECT 92.880 108.755 93.250 109.215 ;
        RECT 93.545 108.615 93.715 108.955 ;
        RECT 93.885 108.785 94.215 109.215 ;
        RECT 94.450 108.615 94.620 108.955 ;
        RECT 90.385 108.155 91.605 108.325 ;
        RECT 91.775 108.245 92.235 108.535 ;
        RECT 92.540 108.415 93.100 108.585 ;
        RECT 93.545 108.445 94.620 108.615 ;
        RECT 94.790 108.715 95.470 109.045 ;
        RECT 95.685 108.715 95.935 109.045 ;
        RECT 96.105 108.755 96.355 109.215 ;
        RECT 92.930 108.275 93.100 108.415 ;
        RECT 91.775 108.235 92.740 108.245 ;
        RECT 91.435 108.065 91.605 108.155 ;
        RECT 92.065 108.075 92.740 108.235 ;
        RECT 90.045 107.865 90.390 107.875 ;
        RECT 88.360 107.655 90.390 107.865 ;
        RECT 85.405 107.215 86.155 107.385 ;
        RECT 85.400 106.665 85.730 107.045 ;
        RECT 85.900 106.925 86.155 107.215 ;
        RECT 86.330 106.665 86.620 107.390 ;
        RECT 87.765 107.315 89.530 107.485 ;
        RECT 88.020 106.665 88.190 107.135 ;
        RECT 88.360 106.835 88.690 107.315 ;
        RECT 88.860 106.665 89.030 107.135 ;
        RECT 89.200 106.835 89.530 107.315 ;
        RECT 89.700 106.665 89.870 107.475 ;
        RECT 90.065 107.400 90.390 107.655 ;
        RECT 90.070 107.045 90.390 107.400 ;
        RECT 90.560 107.615 91.100 107.985 ;
        RECT 91.435 107.895 91.840 108.065 ;
        RECT 90.560 107.215 90.800 107.615 ;
        RECT 91.280 107.445 91.500 107.725 ;
        RECT 90.970 107.275 91.500 107.445 ;
        RECT 90.970 107.045 91.140 107.275 ;
        RECT 91.670 107.115 91.840 107.895 ;
        RECT 92.010 107.285 92.360 107.905 ;
        RECT 92.530 107.285 92.740 108.075 ;
        RECT 92.930 108.105 94.430 108.275 ;
        RECT 92.930 107.415 93.100 108.105 ;
        RECT 94.790 107.935 94.960 108.715 ;
        RECT 95.765 108.585 95.935 108.715 ;
        RECT 93.270 107.765 94.960 107.935 ;
        RECT 95.130 108.155 95.595 108.545 ;
        RECT 95.765 108.415 96.160 108.585 ;
        RECT 93.270 107.585 93.440 107.765 ;
        RECT 90.070 106.875 91.140 107.045 ;
        RECT 91.310 106.665 91.500 107.105 ;
        RECT 91.670 106.835 92.620 107.115 ;
        RECT 92.930 107.025 93.190 107.415 ;
        RECT 93.610 107.345 94.400 107.595 ;
        RECT 92.840 106.855 93.190 107.025 ;
        RECT 93.400 106.665 93.730 107.125 ;
        RECT 94.605 107.055 94.775 107.765 ;
        RECT 95.130 107.565 95.300 108.155 ;
        RECT 94.945 107.345 95.300 107.565 ;
        RECT 95.470 107.345 95.820 107.965 ;
        RECT 95.990 107.055 96.160 108.415 ;
        RECT 96.525 108.245 96.850 109.030 ;
        RECT 96.330 107.195 96.790 108.245 ;
        RECT 94.605 106.885 95.460 107.055 ;
        RECT 95.665 106.885 96.160 107.055 ;
        RECT 96.330 106.665 96.660 107.025 ;
        RECT 97.020 106.925 97.190 109.045 ;
        RECT 97.360 108.715 97.690 109.215 ;
        RECT 97.860 108.545 98.115 109.045 ;
        RECT 97.365 108.375 98.115 108.545 ;
        RECT 97.365 107.385 97.595 108.375 ;
        RECT 97.765 107.555 98.115 108.205 ;
        RECT 98.290 108.140 98.560 109.045 ;
        RECT 98.730 108.455 99.060 109.215 ;
        RECT 99.240 108.285 99.410 109.045 ;
        RECT 100.900 108.375 101.070 109.215 ;
        RECT 97.365 107.215 98.115 107.385 ;
        RECT 97.360 106.665 97.690 107.045 ;
        RECT 97.860 106.925 98.115 107.215 ;
        RECT 98.290 107.340 98.460 108.140 ;
        RECT 98.745 108.115 99.410 108.285 ;
        RECT 101.280 108.205 101.530 109.045 ;
        RECT 101.740 108.375 101.910 109.215 ;
        RECT 102.080 108.205 102.370 109.045 ;
        RECT 98.745 107.970 98.915 108.115 ;
        RECT 98.630 107.640 98.915 107.970 ;
        RECT 100.645 108.035 102.370 108.205 ;
        RECT 102.580 108.155 102.750 109.215 ;
        RECT 103.045 108.835 103.375 109.215 ;
        RECT 103.555 108.665 103.725 108.955 ;
        RECT 103.895 108.755 104.145 109.215 ;
        RECT 102.925 108.495 103.725 108.665 ;
        RECT 104.315 108.705 105.185 109.045 ;
        RECT 98.745 107.385 98.915 107.640 ;
        RECT 99.150 107.565 99.480 107.935 ;
        RECT 100.645 107.485 101.055 108.035 ;
        RECT 102.925 107.875 103.095 108.495 ;
        RECT 104.315 108.325 104.485 108.705 ;
        RECT 105.420 108.585 105.590 109.045 ;
        RECT 105.760 108.755 106.130 109.215 ;
        RECT 106.425 108.615 106.595 108.955 ;
        RECT 106.765 108.785 107.095 109.215 ;
        RECT 107.330 108.615 107.500 108.955 ;
        RECT 103.265 108.155 104.485 108.325 ;
        RECT 104.655 108.245 105.115 108.535 ;
        RECT 105.420 108.415 105.980 108.585 ;
        RECT 106.425 108.445 107.500 108.615 ;
        RECT 107.670 108.715 108.350 109.045 ;
        RECT 108.565 108.715 108.815 109.045 ;
        RECT 108.985 108.755 109.235 109.215 ;
        RECT 105.810 108.275 105.980 108.415 ;
        RECT 104.655 108.235 105.620 108.245 ;
        RECT 104.315 108.065 104.485 108.155 ;
        RECT 104.945 108.075 105.620 108.235 ;
        RECT 102.925 107.865 103.270 107.875 ;
        RECT 101.240 107.655 103.270 107.865 ;
        RECT 98.290 106.835 98.550 107.340 ;
        RECT 98.745 107.215 99.410 107.385 ;
        RECT 100.645 107.315 102.410 107.485 ;
        RECT 98.730 106.665 99.060 107.045 ;
        RECT 99.240 106.835 99.410 107.215 ;
        RECT 100.900 106.665 101.070 107.135 ;
        RECT 101.240 106.835 101.570 107.315 ;
        RECT 101.740 106.665 101.910 107.135 ;
        RECT 102.080 106.835 102.410 107.315 ;
        RECT 102.580 106.665 102.750 107.475 ;
        RECT 102.945 107.400 103.270 107.655 ;
        RECT 102.950 107.045 103.270 107.400 ;
        RECT 103.440 107.615 103.980 107.985 ;
        RECT 104.315 107.895 104.720 108.065 ;
        RECT 103.440 107.215 103.680 107.615 ;
        RECT 104.160 107.445 104.380 107.725 ;
        RECT 103.850 107.275 104.380 107.445 ;
        RECT 103.850 107.045 104.020 107.275 ;
        RECT 104.550 107.115 104.720 107.895 ;
        RECT 104.890 107.285 105.240 107.905 ;
        RECT 105.410 107.285 105.620 108.075 ;
        RECT 105.810 108.105 107.310 108.275 ;
        RECT 105.810 107.415 105.980 108.105 ;
        RECT 107.670 107.935 107.840 108.715 ;
        RECT 108.645 108.585 108.815 108.715 ;
        RECT 106.150 107.765 107.840 107.935 ;
        RECT 108.010 108.155 108.475 108.545 ;
        RECT 108.645 108.415 109.040 108.585 ;
        RECT 106.150 107.585 106.320 107.765 ;
        RECT 102.950 106.875 104.020 107.045 ;
        RECT 104.190 106.665 104.380 107.105 ;
        RECT 104.550 106.835 105.500 107.115 ;
        RECT 105.810 107.025 106.070 107.415 ;
        RECT 106.490 107.345 107.280 107.595 ;
        RECT 105.720 106.855 106.070 107.025 ;
        RECT 106.280 106.665 106.610 107.125 ;
        RECT 107.485 107.055 107.655 107.765 ;
        RECT 108.010 107.565 108.180 108.155 ;
        RECT 107.825 107.345 108.180 107.565 ;
        RECT 108.350 107.345 108.700 107.965 ;
        RECT 108.870 107.055 109.040 108.415 ;
        RECT 109.405 108.245 109.730 109.030 ;
        RECT 109.210 107.195 109.670 108.245 ;
        RECT 107.485 106.885 108.340 107.055 ;
        RECT 108.545 106.885 109.040 107.055 ;
        RECT 109.210 106.665 109.540 107.025 ;
        RECT 109.900 106.925 110.070 109.045 ;
        RECT 110.240 108.715 110.570 109.215 ;
        RECT 110.740 108.545 110.995 109.045 ;
        RECT 110.245 108.375 110.995 108.545 ;
        RECT 110.245 107.385 110.475 108.375 ;
        RECT 110.645 107.555 110.995 108.205 ;
        RECT 111.170 108.125 112.380 109.215 ;
        RECT 111.170 107.585 111.690 108.125 ;
        RECT 111.860 107.415 112.380 107.955 ;
        RECT 110.245 107.215 110.995 107.385 ;
        RECT 110.240 106.665 110.570 107.045 ;
        RECT 110.740 106.925 110.995 107.215 ;
        RECT 111.170 106.665 112.380 107.415 ;
        RECT 18.165 106.495 112.465 106.665 ;
        RECT 18.250 105.745 19.460 106.495 ;
        RECT 18.250 105.205 18.770 105.745 ;
        RECT 20.090 105.725 21.760 106.495 ;
        RECT 21.930 105.770 22.220 106.495 ;
        RECT 18.940 105.035 19.460 105.575 ;
        RECT 18.250 103.945 19.460 105.035 ;
        RECT 20.090 105.035 20.840 105.555 ;
        RECT 21.010 105.205 21.760 105.725 ;
        RECT 22.450 105.675 22.660 106.495 ;
        RECT 22.830 105.695 23.160 106.325 ;
        RECT 20.090 103.945 21.760 105.035 ;
        RECT 21.930 103.945 22.220 105.110 ;
        RECT 22.830 105.095 23.080 105.695 ;
        RECT 23.330 105.675 23.560 106.495 ;
        RECT 23.810 105.675 24.040 106.495 ;
        RECT 24.210 105.695 24.540 106.325 ;
        RECT 23.250 105.255 23.580 105.505 ;
        RECT 23.790 105.255 24.120 105.505 ;
        RECT 24.290 105.095 24.540 105.695 ;
        RECT 24.710 105.675 24.920 106.495 ;
        RECT 25.190 105.675 25.420 106.495 ;
        RECT 25.590 105.695 25.920 106.325 ;
        RECT 25.170 105.255 25.500 105.505 ;
        RECT 25.670 105.095 25.920 105.695 ;
        RECT 26.090 105.675 26.300 106.495 ;
        RECT 26.535 105.945 26.790 106.235 ;
        RECT 26.960 106.115 27.290 106.495 ;
        RECT 26.535 105.775 27.285 105.945 ;
        RECT 22.450 103.945 22.660 105.085 ;
        RECT 22.830 104.115 23.160 105.095 ;
        RECT 23.330 103.945 23.560 105.085 ;
        RECT 23.810 103.945 24.040 105.085 ;
        RECT 24.210 104.115 24.540 105.095 ;
        RECT 24.710 103.945 24.920 105.085 ;
        RECT 25.190 103.945 25.420 105.085 ;
        RECT 25.590 104.115 25.920 105.095 ;
        RECT 26.090 103.945 26.300 105.085 ;
        RECT 26.535 104.955 26.885 105.605 ;
        RECT 27.055 104.785 27.285 105.775 ;
        RECT 26.535 104.615 27.285 104.785 ;
        RECT 26.535 104.115 26.790 104.615 ;
        RECT 26.960 103.945 27.290 104.445 ;
        RECT 27.460 104.115 27.630 106.235 ;
        RECT 27.990 106.135 28.320 106.495 ;
        RECT 28.490 106.105 28.985 106.275 ;
        RECT 29.190 106.105 30.045 106.275 ;
        RECT 27.860 104.915 28.320 105.965 ;
        RECT 27.800 104.130 28.125 104.915 ;
        RECT 28.490 104.745 28.660 106.105 ;
        RECT 28.830 105.195 29.180 105.815 ;
        RECT 29.350 105.595 29.705 105.815 ;
        RECT 29.350 105.005 29.520 105.595 ;
        RECT 29.875 105.395 30.045 106.105 ;
        RECT 30.920 106.035 31.250 106.495 ;
        RECT 31.460 106.135 31.810 106.305 ;
        RECT 30.250 105.565 31.040 105.815 ;
        RECT 31.460 105.745 31.720 106.135 ;
        RECT 32.030 106.045 32.980 106.325 ;
        RECT 33.150 106.055 33.340 106.495 ;
        RECT 33.510 106.115 34.580 106.285 ;
        RECT 31.210 105.395 31.380 105.575 ;
        RECT 28.490 104.575 28.885 104.745 ;
        RECT 29.055 104.615 29.520 105.005 ;
        RECT 29.690 105.225 31.380 105.395 ;
        RECT 28.715 104.445 28.885 104.575 ;
        RECT 29.690 104.445 29.860 105.225 ;
        RECT 31.550 105.055 31.720 105.745 ;
        RECT 30.220 104.885 31.720 105.055 ;
        RECT 31.910 105.085 32.120 105.875 ;
        RECT 32.290 105.255 32.640 105.875 ;
        RECT 32.810 105.265 32.980 106.045 ;
        RECT 33.510 105.885 33.680 106.115 ;
        RECT 33.150 105.715 33.680 105.885 ;
        RECT 33.150 105.435 33.370 105.715 ;
        RECT 33.850 105.545 34.090 105.945 ;
        RECT 32.810 105.095 33.215 105.265 ;
        RECT 33.550 105.175 34.090 105.545 ;
        RECT 34.260 105.760 34.580 106.115 ;
        RECT 34.260 105.505 34.585 105.760 ;
        RECT 34.780 105.685 34.950 106.495 ;
        RECT 35.120 105.845 35.450 106.325 ;
        RECT 35.620 106.025 35.790 106.495 ;
        RECT 35.960 105.845 36.290 106.325 ;
        RECT 36.460 106.025 36.630 106.495 ;
        RECT 37.115 105.945 37.370 106.235 ;
        RECT 37.540 106.115 37.870 106.495 ;
        RECT 35.120 105.675 36.885 105.845 ;
        RECT 37.115 105.775 37.865 105.945 ;
        RECT 34.260 105.295 36.290 105.505 ;
        RECT 34.260 105.285 34.605 105.295 ;
        RECT 31.910 104.925 32.585 105.085 ;
        RECT 33.045 105.005 33.215 105.095 ;
        RECT 31.910 104.915 32.875 104.925 ;
        RECT 31.550 104.745 31.720 104.885 ;
        RECT 28.295 103.945 28.545 104.405 ;
        RECT 28.715 104.115 28.965 104.445 ;
        RECT 29.180 104.115 29.860 104.445 ;
        RECT 30.030 104.545 31.105 104.715 ;
        RECT 31.550 104.575 32.110 104.745 ;
        RECT 32.415 104.625 32.875 104.915 ;
        RECT 33.045 104.835 34.265 105.005 ;
        RECT 30.030 104.205 30.200 104.545 ;
        RECT 30.435 103.945 30.765 104.375 ;
        RECT 30.935 104.205 31.105 104.545 ;
        RECT 31.400 103.945 31.770 104.405 ;
        RECT 31.940 104.115 32.110 104.575 ;
        RECT 33.045 104.455 33.215 104.835 ;
        RECT 34.435 104.665 34.605 105.285 ;
        RECT 36.475 105.125 36.885 105.675 ;
        RECT 32.345 104.115 33.215 104.455 ;
        RECT 33.805 104.495 34.605 104.665 ;
        RECT 33.385 103.945 33.635 104.405 ;
        RECT 33.805 104.205 33.975 104.495 ;
        RECT 34.155 103.945 34.485 104.325 ;
        RECT 34.780 103.945 34.950 105.005 ;
        RECT 35.160 104.955 36.885 105.125 ;
        RECT 37.115 104.955 37.465 105.605 ;
        RECT 35.160 104.115 35.450 104.955 ;
        RECT 35.620 103.945 35.790 104.785 ;
        RECT 36.000 104.115 36.250 104.955 ;
        RECT 37.635 104.785 37.865 105.775 ;
        RECT 36.460 103.945 36.630 104.785 ;
        RECT 37.115 104.615 37.865 104.785 ;
        RECT 37.115 104.115 37.370 104.615 ;
        RECT 37.540 103.945 37.870 104.445 ;
        RECT 38.040 104.115 38.210 106.235 ;
        RECT 38.570 106.135 38.900 106.495 ;
        RECT 39.070 106.105 39.565 106.275 ;
        RECT 39.770 106.105 40.625 106.275 ;
        RECT 38.440 104.915 38.900 105.965 ;
        RECT 38.380 104.130 38.705 104.915 ;
        RECT 39.070 104.745 39.240 106.105 ;
        RECT 39.410 105.195 39.760 105.815 ;
        RECT 39.930 105.595 40.285 105.815 ;
        RECT 39.930 105.005 40.100 105.595 ;
        RECT 40.455 105.395 40.625 106.105 ;
        RECT 41.500 106.035 41.830 106.495 ;
        RECT 42.040 106.135 42.390 106.305 ;
        RECT 40.830 105.565 41.620 105.815 ;
        RECT 42.040 105.745 42.300 106.135 ;
        RECT 42.610 106.045 43.560 106.325 ;
        RECT 43.730 106.055 43.920 106.495 ;
        RECT 44.090 106.115 45.160 106.285 ;
        RECT 41.790 105.395 41.960 105.575 ;
        RECT 39.070 104.575 39.465 104.745 ;
        RECT 39.635 104.615 40.100 105.005 ;
        RECT 40.270 105.225 41.960 105.395 ;
        RECT 39.295 104.445 39.465 104.575 ;
        RECT 40.270 104.445 40.440 105.225 ;
        RECT 42.130 105.055 42.300 105.745 ;
        RECT 40.800 104.885 42.300 105.055 ;
        RECT 42.490 105.085 42.700 105.875 ;
        RECT 42.870 105.255 43.220 105.875 ;
        RECT 43.390 105.265 43.560 106.045 ;
        RECT 44.090 105.885 44.260 106.115 ;
        RECT 43.730 105.715 44.260 105.885 ;
        RECT 43.730 105.435 43.950 105.715 ;
        RECT 44.430 105.545 44.670 105.945 ;
        RECT 43.390 105.095 43.795 105.265 ;
        RECT 44.130 105.175 44.670 105.545 ;
        RECT 44.840 105.760 45.160 106.115 ;
        RECT 44.840 105.505 45.165 105.760 ;
        RECT 45.360 105.685 45.530 106.495 ;
        RECT 45.700 105.845 46.030 106.325 ;
        RECT 46.200 106.025 46.370 106.495 ;
        RECT 46.540 105.845 46.870 106.325 ;
        RECT 47.040 106.025 47.210 106.495 ;
        RECT 45.700 105.675 47.465 105.845 ;
        RECT 47.690 105.770 47.980 106.495 ;
        RECT 48.210 105.675 48.420 106.495 ;
        RECT 48.590 105.695 48.920 106.325 ;
        RECT 44.840 105.295 46.870 105.505 ;
        RECT 44.840 105.285 45.185 105.295 ;
        RECT 42.490 104.925 43.165 105.085 ;
        RECT 43.625 105.005 43.795 105.095 ;
        RECT 42.490 104.915 43.455 104.925 ;
        RECT 42.130 104.745 42.300 104.885 ;
        RECT 38.875 103.945 39.125 104.405 ;
        RECT 39.295 104.115 39.545 104.445 ;
        RECT 39.760 104.115 40.440 104.445 ;
        RECT 40.610 104.545 41.685 104.715 ;
        RECT 42.130 104.575 42.690 104.745 ;
        RECT 42.995 104.625 43.455 104.915 ;
        RECT 43.625 104.835 44.845 105.005 ;
        RECT 40.610 104.205 40.780 104.545 ;
        RECT 41.015 103.945 41.345 104.375 ;
        RECT 41.515 104.205 41.685 104.545 ;
        RECT 41.980 103.945 42.350 104.405 ;
        RECT 42.520 104.115 42.690 104.575 ;
        RECT 43.625 104.455 43.795 104.835 ;
        RECT 45.015 104.665 45.185 105.285 ;
        RECT 47.055 105.125 47.465 105.675 ;
        RECT 42.925 104.115 43.795 104.455 ;
        RECT 44.385 104.495 45.185 104.665 ;
        RECT 43.965 103.945 44.215 104.405 ;
        RECT 44.385 104.205 44.555 104.495 ;
        RECT 44.735 103.945 45.065 104.325 ;
        RECT 45.360 103.945 45.530 105.005 ;
        RECT 45.740 104.955 47.465 105.125 ;
        RECT 45.740 104.115 46.030 104.955 ;
        RECT 46.200 103.945 46.370 104.785 ;
        RECT 46.580 104.115 46.830 104.955 ;
        RECT 47.040 103.945 47.210 104.785 ;
        RECT 47.690 103.945 47.980 105.110 ;
        RECT 48.590 105.095 48.840 105.695 ;
        RECT 49.090 105.675 49.320 106.495 ;
        RECT 49.570 105.675 49.800 106.495 ;
        RECT 49.970 105.695 50.300 106.325 ;
        RECT 49.010 105.255 49.340 105.505 ;
        RECT 49.550 105.255 49.880 105.505 ;
        RECT 50.050 105.095 50.300 105.695 ;
        RECT 50.470 105.675 50.680 106.495 ;
        RECT 51.220 106.025 51.390 106.495 ;
        RECT 51.560 105.845 51.890 106.325 ;
        RECT 52.060 106.025 52.230 106.495 ;
        RECT 52.400 105.845 52.730 106.325 ;
        RECT 50.965 105.675 52.730 105.845 ;
        RECT 52.900 105.685 53.070 106.495 ;
        RECT 53.270 106.115 54.340 106.285 ;
        RECT 53.270 105.760 53.590 106.115 ;
        RECT 48.210 103.945 48.420 105.085 ;
        RECT 48.590 104.115 48.920 105.095 ;
        RECT 49.090 103.945 49.320 105.085 ;
        RECT 49.570 103.945 49.800 105.085 ;
        RECT 49.970 104.115 50.300 105.095 ;
        RECT 50.965 105.125 51.375 105.675 ;
        RECT 53.265 105.505 53.590 105.760 ;
        RECT 51.560 105.295 53.590 105.505 ;
        RECT 53.245 105.285 53.590 105.295 ;
        RECT 53.760 105.545 54.000 105.945 ;
        RECT 54.170 105.885 54.340 106.115 ;
        RECT 54.510 106.055 54.700 106.495 ;
        RECT 54.870 106.045 55.820 106.325 ;
        RECT 56.040 106.135 56.390 106.305 ;
        RECT 54.170 105.715 54.700 105.885 ;
        RECT 50.470 103.945 50.680 105.085 ;
        RECT 50.965 104.955 52.690 105.125 ;
        RECT 51.220 103.945 51.390 104.785 ;
        RECT 51.600 104.115 51.850 104.955 ;
        RECT 52.060 103.945 52.230 104.785 ;
        RECT 52.400 104.115 52.690 104.955 ;
        RECT 52.900 103.945 53.070 105.005 ;
        RECT 53.245 104.665 53.415 105.285 ;
        RECT 53.760 105.175 54.300 105.545 ;
        RECT 54.480 105.435 54.700 105.715 ;
        RECT 54.870 105.265 55.040 106.045 ;
        RECT 54.635 105.095 55.040 105.265 ;
        RECT 55.210 105.255 55.560 105.875 ;
        RECT 54.635 105.005 54.805 105.095 ;
        RECT 55.730 105.085 55.940 105.875 ;
        RECT 53.585 104.835 54.805 105.005 ;
        RECT 55.265 104.925 55.940 105.085 ;
        RECT 53.245 104.495 54.045 104.665 ;
        RECT 53.365 103.945 53.695 104.325 ;
        RECT 53.875 104.205 54.045 104.495 ;
        RECT 54.635 104.455 54.805 104.835 ;
        RECT 54.975 104.915 55.940 104.925 ;
        RECT 56.130 105.745 56.390 106.135 ;
        RECT 56.600 106.035 56.930 106.495 ;
        RECT 57.805 106.105 58.660 106.275 ;
        RECT 58.865 106.105 59.360 106.275 ;
        RECT 59.530 106.135 59.860 106.495 ;
        RECT 56.130 105.055 56.300 105.745 ;
        RECT 56.470 105.395 56.640 105.575 ;
        RECT 56.810 105.565 57.600 105.815 ;
        RECT 57.805 105.395 57.975 106.105 ;
        RECT 58.145 105.595 58.500 105.815 ;
        RECT 56.470 105.225 58.160 105.395 ;
        RECT 54.975 104.625 55.435 104.915 ;
        RECT 56.130 104.885 57.630 105.055 ;
        RECT 56.130 104.745 56.300 104.885 ;
        RECT 55.740 104.575 56.300 104.745 ;
        RECT 54.215 103.945 54.465 104.405 ;
        RECT 54.635 104.115 55.505 104.455 ;
        RECT 55.740 104.115 55.910 104.575 ;
        RECT 56.745 104.545 57.820 104.715 ;
        RECT 56.080 103.945 56.450 104.405 ;
        RECT 56.745 104.205 56.915 104.545 ;
        RECT 57.085 103.945 57.415 104.375 ;
        RECT 57.650 104.205 57.820 104.545 ;
        RECT 57.990 104.445 58.160 105.225 ;
        RECT 58.330 105.005 58.500 105.595 ;
        RECT 58.670 105.195 59.020 105.815 ;
        RECT 58.330 104.615 58.795 105.005 ;
        RECT 59.190 104.745 59.360 106.105 ;
        RECT 59.530 104.915 59.990 105.965 ;
        RECT 58.965 104.575 59.360 104.745 ;
        RECT 58.965 104.445 59.135 104.575 ;
        RECT 57.990 104.115 58.670 104.445 ;
        RECT 58.885 104.115 59.135 104.445 ;
        RECT 59.305 103.945 59.555 104.405 ;
        RECT 59.725 104.130 60.050 104.915 ;
        RECT 60.220 104.115 60.390 106.235 ;
        RECT 60.560 106.115 60.890 106.495 ;
        RECT 61.060 105.945 61.315 106.235 ;
        RECT 61.800 106.025 61.970 106.495 ;
        RECT 60.565 105.775 61.315 105.945 ;
        RECT 62.140 105.845 62.470 106.325 ;
        RECT 62.640 106.025 62.810 106.495 ;
        RECT 62.980 105.845 63.310 106.325 ;
        RECT 60.565 104.785 60.795 105.775 ;
        RECT 61.545 105.675 63.310 105.845 ;
        RECT 63.480 105.685 63.650 106.495 ;
        RECT 63.850 106.115 64.920 106.285 ;
        RECT 63.850 105.760 64.170 106.115 ;
        RECT 60.965 104.955 61.315 105.605 ;
        RECT 61.545 105.125 61.955 105.675 ;
        RECT 63.845 105.505 64.170 105.760 ;
        RECT 62.140 105.295 64.170 105.505 ;
        RECT 63.825 105.285 64.170 105.295 ;
        RECT 64.340 105.545 64.580 105.945 ;
        RECT 64.750 105.885 64.920 106.115 ;
        RECT 65.090 106.055 65.280 106.495 ;
        RECT 65.450 106.045 66.400 106.325 ;
        RECT 66.620 106.135 66.970 106.305 ;
        RECT 64.750 105.715 65.280 105.885 ;
        RECT 61.545 104.955 63.270 105.125 ;
        RECT 60.565 104.615 61.315 104.785 ;
        RECT 60.560 103.945 60.890 104.445 ;
        RECT 61.060 104.115 61.315 104.615 ;
        RECT 61.800 103.945 61.970 104.785 ;
        RECT 62.180 104.115 62.430 104.955 ;
        RECT 62.640 103.945 62.810 104.785 ;
        RECT 62.980 104.115 63.270 104.955 ;
        RECT 63.480 103.945 63.650 105.005 ;
        RECT 63.825 104.665 63.995 105.285 ;
        RECT 64.340 105.175 64.880 105.545 ;
        RECT 65.060 105.435 65.280 105.715 ;
        RECT 65.450 105.265 65.620 106.045 ;
        RECT 65.215 105.095 65.620 105.265 ;
        RECT 65.790 105.255 66.140 105.875 ;
        RECT 65.215 105.005 65.385 105.095 ;
        RECT 66.310 105.085 66.520 105.875 ;
        RECT 64.165 104.835 65.385 105.005 ;
        RECT 65.845 104.925 66.520 105.085 ;
        RECT 63.825 104.495 64.625 104.665 ;
        RECT 63.945 103.945 64.275 104.325 ;
        RECT 64.455 104.205 64.625 104.495 ;
        RECT 65.215 104.455 65.385 104.835 ;
        RECT 65.555 104.915 66.520 104.925 ;
        RECT 66.710 105.745 66.970 106.135 ;
        RECT 67.180 106.035 67.510 106.495 ;
        RECT 68.385 106.105 69.240 106.275 ;
        RECT 69.445 106.105 69.940 106.275 ;
        RECT 70.110 106.135 70.440 106.495 ;
        RECT 66.710 105.055 66.880 105.745 ;
        RECT 67.050 105.395 67.220 105.575 ;
        RECT 67.390 105.565 68.180 105.815 ;
        RECT 68.385 105.395 68.555 106.105 ;
        RECT 68.725 105.595 69.080 105.815 ;
        RECT 67.050 105.225 68.740 105.395 ;
        RECT 65.555 104.625 66.015 104.915 ;
        RECT 66.710 104.885 68.210 105.055 ;
        RECT 66.710 104.745 66.880 104.885 ;
        RECT 66.320 104.575 66.880 104.745 ;
        RECT 64.795 103.945 65.045 104.405 ;
        RECT 65.215 104.115 66.085 104.455 ;
        RECT 66.320 104.115 66.490 104.575 ;
        RECT 67.325 104.545 68.400 104.715 ;
        RECT 66.660 103.945 67.030 104.405 ;
        RECT 67.325 104.205 67.495 104.545 ;
        RECT 67.665 103.945 67.995 104.375 ;
        RECT 68.230 104.205 68.400 104.545 ;
        RECT 68.570 104.445 68.740 105.225 ;
        RECT 68.910 105.005 69.080 105.595 ;
        RECT 69.250 105.195 69.600 105.815 ;
        RECT 68.910 104.615 69.375 105.005 ;
        RECT 69.770 104.745 69.940 106.105 ;
        RECT 70.110 104.915 70.570 105.965 ;
        RECT 69.545 104.575 69.940 104.745 ;
        RECT 69.545 104.445 69.715 104.575 ;
        RECT 68.570 104.115 69.250 104.445 ;
        RECT 69.465 104.115 69.715 104.445 ;
        RECT 69.885 103.945 70.135 104.405 ;
        RECT 70.305 104.130 70.630 104.915 ;
        RECT 70.800 104.115 70.970 106.235 ;
        RECT 71.140 106.115 71.470 106.495 ;
        RECT 71.640 105.945 71.895 106.235 ;
        RECT 71.145 105.775 71.895 105.945 ;
        RECT 72.160 105.945 72.330 106.325 ;
        RECT 72.510 106.115 72.840 106.495 ;
        RECT 72.160 105.775 72.825 105.945 ;
        RECT 73.020 105.820 73.280 106.325 ;
        RECT 71.145 104.785 71.375 105.775 ;
        RECT 71.545 104.955 71.895 105.605 ;
        RECT 72.090 105.225 72.420 105.595 ;
        RECT 72.655 105.520 72.825 105.775 ;
        RECT 72.655 105.190 72.940 105.520 ;
        RECT 72.655 105.045 72.825 105.190 ;
        RECT 72.160 104.875 72.825 105.045 ;
        RECT 73.110 105.020 73.280 105.820 ;
        RECT 73.450 105.770 73.740 106.495 ;
        RECT 74.220 106.025 74.390 106.495 ;
        RECT 74.560 105.845 74.890 106.325 ;
        RECT 75.060 106.025 75.230 106.495 ;
        RECT 75.400 105.845 75.730 106.325 ;
        RECT 73.965 105.675 75.730 105.845 ;
        RECT 75.900 105.685 76.070 106.495 ;
        RECT 76.270 106.115 77.340 106.285 ;
        RECT 76.270 105.760 76.590 106.115 ;
        RECT 73.965 105.125 74.375 105.675 ;
        RECT 76.265 105.505 76.590 105.760 ;
        RECT 74.560 105.295 76.590 105.505 ;
        RECT 76.245 105.285 76.590 105.295 ;
        RECT 76.760 105.545 77.000 105.945 ;
        RECT 77.170 105.885 77.340 106.115 ;
        RECT 77.510 106.055 77.700 106.495 ;
        RECT 77.870 106.045 78.820 106.325 ;
        RECT 79.040 106.135 79.390 106.305 ;
        RECT 77.170 105.715 77.700 105.885 ;
        RECT 71.145 104.615 71.895 104.785 ;
        RECT 71.140 103.945 71.470 104.445 ;
        RECT 71.640 104.115 71.895 104.615 ;
        RECT 72.160 104.115 72.330 104.875 ;
        RECT 72.510 103.945 72.840 104.705 ;
        RECT 73.010 104.115 73.280 105.020 ;
        RECT 73.450 103.945 73.740 105.110 ;
        RECT 73.965 104.955 75.690 105.125 ;
        RECT 74.220 103.945 74.390 104.785 ;
        RECT 74.600 104.115 74.850 104.955 ;
        RECT 75.060 103.945 75.230 104.785 ;
        RECT 75.400 104.115 75.690 104.955 ;
        RECT 75.900 103.945 76.070 105.005 ;
        RECT 76.245 104.665 76.415 105.285 ;
        RECT 76.760 105.175 77.300 105.545 ;
        RECT 77.480 105.435 77.700 105.715 ;
        RECT 77.870 105.265 78.040 106.045 ;
        RECT 77.635 105.095 78.040 105.265 ;
        RECT 78.210 105.255 78.560 105.875 ;
        RECT 77.635 105.005 77.805 105.095 ;
        RECT 78.730 105.085 78.940 105.875 ;
        RECT 76.585 104.835 77.805 105.005 ;
        RECT 78.265 104.925 78.940 105.085 ;
        RECT 76.245 104.495 77.045 104.665 ;
        RECT 76.365 103.945 76.695 104.325 ;
        RECT 76.875 104.205 77.045 104.495 ;
        RECT 77.635 104.455 77.805 104.835 ;
        RECT 77.975 104.915 78.940 104.925 ;
        RECT 79.130 105.745 79.390 106.135 ;
        RECT 79.600 106.035 79.930 106.495 ;
        RECT 80.805 106.105 81.660 106.275 ;
        RECT 81.865 106.105 82.360 106.275 ;
        RECT 82.530 106.135 82.860 106.495 ;
        RECT 79.130 105.055 79.300 105.745 ;
        RECT 79.470 105.395 79.640 105.575 ;
        RECT 79.810 105.565 80.600 105.815 ;
        RECT 80.805 105.395 80.975 106.105 ;
        RECT 81.145 105.595 81.500 105.815 ;
        RECT 79.470 105.225 81.160 105.395 ;
        RECT 77.975 104.625 78.435 104.915 ;
        RECT 79.130 104.885 80.630 105.055 ;
        RECT 79.130 104.745 79.300 104.885 ;
        RECT 78.740 104.575 79.300 104.745 ;
        RECT 77.215 103.945 77.465 104.405 ;
        RECT 77.635 104.115 78.505 104.455 ;
        RECT 78.740 104.115 78.910 104.575 ;
        RECT 79.745 104.545 80.820 104.715 ;
        RECT 79.080 103.945 79.450 104.405 ;
        RECT 79.745 104.205 79.915 104.545 ;
        RECT 80.085 103.945 80.415 104.375 ;
        RECT 80.650 104.205 80.820 104.545 ;
        RECT 80.990 104.445 81.160 105.225 ;
        RECT 81.330 105.005 81.500 105.595 ;
        RECT 81.670 105.195 82.020 105.815 ;
        RECT 81.330 104.615 81.795 105.005 ;
        RECT 82.190 104.745 82.360 106.105 ;
        RECT 82.530 104.915 82.990 105.965 ;
        RECT 81.965 104.575 82.360 104.745 ;
        RECT 81.965 104.445 82.135 104.575 ;
        RECT 80.990 104.115 81.670 104.445 ;
        RECT 81.885 104.115 82.135 104.445 ;
        RECT 82.305 103.945 82.555 104.405 ;
        RECT 82.725 104.130 83.050 104.915 ;
        RECT 83.220 104.115 83.390 106.235 ;
        RECT 83.560 106.115 83.890 106.495 ;
        RECT 84.060 105.945 84.315 106.235 ;
        RECT 84.800 106.025 84.970 106.495 ;
        RECT 83.565 105.775 84.315 105.945 ;
        RECT 85.140 105.845 85.470 106.325 ;
        RECT 85.640 106.025 85.810 106.495 ;
        RECT 85.980 105.845 86.310 106.325 ;
        RECT 83.565 104.785 83.795 105.775 ;
        RECT 84.545 105.675 86.310 105.845 ;
        RECT 86.480 105.685 86.650 106.495 ;
        RECT 86.850 106.115 87.920 106.285 ;
        RECT 86.850 105.760 87.170 106.115 ;
        RECT 83.965 104.955 84.315 105.605 ;
        RECT 84.545 105.125 84.955 105.675 ;
        RECT 86.845 105.505 87.170 105.760 ;
        RECT 85.140 105.295 87.170 105.505 ;
        RECT 86.825 105.285 87.170 105.295 ;
        RECT 87.340 105.545 87.580 105.945 ;
        RECT 87.750 105.885 87.920 106.115 ;
        RECT 88.090 106.055 88.280 106.495 ;
        RECT 88.450 106.045 89.400 106.325 ;
        RECT 89.620 106.135 89.970 106.305 ;
        RECT 87.750 105.715 88.280 105.885 ;
        RECT 84.545 104.955 86.270 105.125 ;
        RECT 83.565 104.615 84.315 104.785 ;
        RECT 83.560 103.945 83.890 104.445 ;
        RECT 84.060 104.115 84.315 104.615 ;
        RECT 84.800 103.945 84.970 104.785 ;
        RECT 85.180 104.115 85.430 104.955 ;
        RECT 85.640 103.945 85.810 104.785 ;
        RECT 85.980 104.115 86.270 104.955 ;
        RECT 86.480 103.945 86.650 105.005 ;
        RECT 86.825 104.665 86.995 105.285 ;
        RECT 87.340 105.175 87.880 105.545 ;
        RECT 88.060 105.435 88.280 105.715 ;
        RECT 88.450 105.265 88.620 106.045 ;
        RECT 88.215 105.095 88.620 105.265 ;
        RECT 88.790 105.255 89.140 105.875 ;
        RECT 88.215 105.005 88.385 105.095 ;
        RECT 89.310 105.085 89.520 105.875 ;
        RECT 87.165 104.835 88.385 105.005 ;
        RECT 88.845 104.925 89.520 105.085 ;
        RECT 86.825 104.495 87.625 104.665 ;
        RECT 86.945 103.945 87.275 104.325 ;
        RECT 87.455 104.205 87.625 104.495 ;
        RECT 88.215 104.455 88.385 104.835 ;
        RECT 88.555 104.915 89.520 104.925 ;
        RECT 89.710 105.745 89.970 106.135 ;
        RECT 90.180 106.035 90.510 106.495 ;
        RECT 91.385 106.105 92.240 106.275 ;
        RECT 92.445 106.105 92.940 106.275 ;
        RECT 93.110 106.135 93.440 106.495 ;
        RECT 89.710 105.055 89.880 105.745 ;
        RECT 90.050 105.395 90.220 105.575 ;
        RECT 90.390 105.565 91.180 105.815 ;
        RECT 91.385 105.395 91.555 106.105 ;
        RECT 91.725 105.595 92.080 105.815 ;
        RECT 90.050 105.225 91.740 105.395 ;
        RECT 88.555 104.625 89.015 104.915 ;
        RECT 89.710 104.885 91.210 105.055 ;
        RECT 89.710 104.745 89.880 104.885 ;
        RECT 89.320 104.575 89.880 104.745 ;
        RECT 87.795 103.945 88.045 104.405 ;
        RECT 88.215 104.115 89.085 104.455 ;
        RECT 89.320 104.115 89.490 104.575 ;
        RECT 90.325 104.545 91.400 104.715 ;
        RECT 89.660 103.945 90.030 104.405 ;
        RECT 90.325 104.205 90.495 104.545 ;
        RECT 90.665 103.945 90.995 104.375 ;
        RECT 91.230 104.205 91.400 104.545 ;
        RECT 91.570 104.445 91.740 105.225 ;
        RECT 91.910 105.005 92.080 105.595 ;
        RECT 92.250 105.195 92.600 105.815 ;
        RECT 91.910 104.615 92.375 105.005 ;
        RECT 92.770 104.745 92.940 106.105 ;
        RECT 93.110 104.915 93.570 105.965 ;
        RECT 92.545 104.575 92.940 104.745 ;
        RECT 92.545 104.445 92.715 104.575 ;
        RECT 91.570 104.115 92.250 104.445 ;
        RECT 92.465 104.115 92.715 104.445 ;
        RECT 92.885 103.945 93.135 104.405 ;
        RECT 93.305 104.130 93.630 104.915 ;
        RECT 93.800 104.115 93.970 106.235 ;
        RECT 94.140 106.115 94.470 106.495 ;
        RECT 94.640 105.945 94.895 106.235 ;
        RECT 94.145 105.775 94.895 105.945 ;
        RECT 94.145 104.785 94.375 105.775 ;
        RECT 95.130 105.675 95.340 106.495 ;
        RECT 95.510 105.695 95.840 106.325 ;
        RECT 94.545 104.955 94.895 105.605 ;
        RECT 95.510 105.095 95.760 105.695 ;
        RECT 96.010 105.675 96.240 106.495 ;
        RECT 96.510 105.675 96.720 106.495 ;
        RECT 96.890 105.695 97.220 106.325 ;
        RECT 95.930 105.255 96.260 105.505 ;
        RECT 96.890 105.095 97.140 105.695 ;
        RECT 97.390 105.675 97.620 106.495 ;
        RECT 97.870 105.675 98.100 106.495 ;
        RECT 98.270 105.695 98.600 106.325 ;
        RECT 97.310 105.255 97.640 105.505 ;
        RECT 97.850 105.255 98.180 105.505 ;
        RECT 98.350 105.095 98.600 105.695 ;
        RECT 98.770 105.675 98.980 106.495 ;
        RECT 99.210 105.770 99.500 106.495 ;
        RECT 99.980 106.025 100.150 106.495 ;
        RECT 100.320 105.845 100.650 106.325 ;
        RECT 100.820 106.025 100.990 106.495 ;
        RECT 101.160 105.845 101.490 106.325 ;
        RECT 99.725 105.675 101.490 105.845 ;
        RECT 101.660 105.685 101.830 106.495 ;
        RECT 102.030 106.115 103.100 106.285 ;
        RECT 102.030 105.760 102.350 106.115 ;
        RECT 99.725 105.125 100.135 105.675 ;
        RECT 102.025 105.505 102.350 105.760 ;
        RECT 100.320 105.295 102.350 105.505 ;
        RECT 102.005 105.285 102.350 105.295 ;
        RECT 102.520 105.545 102.760 105.945 ;
        RECT 102.930 105.885 103.100 106.115 ;
        RECT 103.270 106.055 103.460 106.495 ;
        RECT 103.630 106.045 104.580 106.325 ;
        RECT 104.800 106.135 105.150 106.305 ;
        RECT 102.930 105.715 103.460 105.885 ;
        RECT 94.145 104.615 94.895 104.785 ;
        RECT 94.140 103.945 94.470 104.445 ;
        RECT 94.640 104.115 94.895 104.615 ;
        RECT 95.130 103.945 95.340 105.085 ;
        RECT 95.510 104.115 95.840 105.095 ;
        RECT 96.010 103.945 96.240 105.085 ;
        RECT 96.510 103.945 96.720 105.085 ;
        RECT 96.890 104.115 97.220 105.095 ;
        RECT 97.390 103.945 97.620 105.085 ;
        RECT 97.870 103.945 98.100 105.085 ;
        RECT 98.270 104.115 98.600 105.095 ;
        RECT 98.770 103.945 98.980 105.085 ;
        RECT 99.210 103.945 99.500 105.110 ;
        RECT 99.725 104.955 101.450 105.125 ;
        RECT 99.980 103.945 100.150 104.785 ;
        RECT 100.360 104.115 100.610 104.955 ;
        RECT 100.820 103.945 100.990 104.785 ;
        RECT 101.160 104.115 101.450 104.955 ;
        RECT 101.660 103.945 101.830 105.005 ;
        RECT 102.005 104.665 102.175 105.285 ;
        RECT 102.520 105.175 103.060 105.545 ;
        RECT 103.240 105.435 103.460 105.715 ;
        RECT 103.630 105.265 103.800 106.045 ;
        RECT 103.395 105.095 103.800 105.265 ;
        RECT 103.970 105.255 104.320 105.875 ;
        RECT 103.395 105.005 103.565 105.095 ;
        RECT 104.490 105.085 104.700 105.875 ;
        RECT 102.345 104.835 103.565 105.005 ;
        RECT 104.025 104.925 104.700 105.085 ;
        RECT 102.005 104.495 102.805 104.665 ;
        RECT 102.125 103.945 102.455 104.325 ;
        RECT 102.635 104.205 102.805 104.495 ;
        RECT 103.395 104.455 103.565 104.835 ;
        RECT 103.735 104.915 104.700 104.925 ;
        RECT 104.890 105.745 105.150 106.135 ;
        RECT 105.360 106.035 105.690 106.495 ;
        RECT 106.565 106.105 107.420 106.275 ;
        RECT 107.625 106.105 108.120 106.275 ;
        RECT 108.290 106.135 108.620 106.495 ;
        RECT 104.890 105.055 105.060 105.745 ;
        RECT 105.230 105.395 105.400 105.575 ;
        RECT 105.570 105.565 106.360 105.815 ;
        RECT 106.565 105.395 106.735 106.105 ;
        RECT 106.905 105.595 107.260 105.815 ;
        RECT 105.230 105.225 106.920 105.395 ;
        RECT 103.735 104.625 104.195 104.915 ;
        RECT 104.890 104.885 106.390 105.055 ;
        RECT 104.890 104.745 105.060 104.885 ;
        RECT 104.500 104.575 105.060 104.745 ;
        RECT 102.975 103.945 103.225 104.405 ;
        RECT 103.395 104.115 104.265 104.455 ;
        RECT 104.500 104.115 104.670 104.575 ;
        RECT 105.505 104.545 106.580 104.715 ;
        RECT 104.840 103.945 105.210 104.405 ;
        RECT 105.505 104.205 105.675 104.545 ;
        RECT 105.845 103.945 106.175 104.375 ;
        RECT 106.410 104.205 106.580 104.545 ;
        RECT 106.750 104.445 106.920 105.225 ;
        RECT 107.090 105.005 107.260 105.595 ;
        RECT 107.430 105.195 107.780 105.815 ;
        RECT 107.090 104.615 107.555 105.005 ;
        RECT 107.950 104.745 108.120 106.105 ;
        RECT 108.290 104.915 108.750 105.965 ;
        RECT 107.725 104.575 108.120 104.745 ;
        RECT 107.725 104.445 107.895 104.575 ;
        RECT 106.750 104.115 107.430 104.445 ;
        RECT 107.645 104.115 107.895 104.445 ;
        RECT 108.065 103.945 108.315 104.405 ;
        RECT 108.485 104.130 108.810 104.915 ;
        RECT 108.980 104.115 109.150 106.235 ;
        RECT 109.320 106.115 109.650 106.495 ;
        RECT 109.820 105.945 110.075 106.235 ;
        RECT 109.325 105.775 110.075 105.945 ;
        RECT 109.325 104.785 109.555 105.775 ;
        RECT 111.170 105.745 112.380 106.495 ;
        RECT 109.725 104.955 110.075 105.605 ;
        RECT 111.170 105.035 111.690 105.575 ;
        RECT 111.860 105.205 112.380 105.745 ;
        RECT 109.325 104.615 110.075 104.785 ;
        RECT 109.320 103.945 109.650 104.445 ;
        RECT 109.820 104.115 110.075 104.615 ;
        RECT 111.170 103.945 112.380 105.035 ;
        RECT 18.165 103.775 112.465 103.945 ;
        RECT 18.250 102.685 19.460 103.775 ;
        RECT 18.250 101.975 18.770 102.515 ;
        RECT 18.940 102.145 19.460 102.685 ;
        RECT 20.090 102.685 21.760 103.775 ;
        RECT 20.090 102.165 20.840 102.685 ;
        RECT 21.930 102.610 22.220 103.775 ;
        RECT 22.700 102.935 22.870 103.775 ;
        RECT 23.080 102.765 23.330 103.605 ;
        RECT 23.540 102.935 23.710 103.775 ;
        RECT 23.880 102.765 24.170 103.605 ;
        RECT 22.445 102.595 24.170 102.765 ;
        RECT 24.380 102.715 24.550 103.775 ;
        RECT 24.845 103.395 25.175 103.775 ;
        RECT 25.355 103.225 25.525 103.515 ;
        RECT 25.695 103.315 25.945 103.775 ;
        RECT 24.725 103.055 25.525 103.225 ;
        RECT 26.115 103.265 26.985 103.605 ;
        RECT 21.010 101.995 21.760 102.515 ;
        RECT 18.250 101.225 19.460 101.975 ;
        RECT 20.090 101.225 21.760 101.995 ;
        RECT 22.445 102.045 22.855 102.595 ;
        RECT 24.725 102.435 24.895 103.055 ;
        RECT 26.115 102.885 26.285 103.265 ;
        RECT 27.220 103.145 27.390 103.605 ;
        RECT 27.560 103.315 27.930 103.775 ;
        RECT 28.225 103.175 28.395 103.515 ;
        RECT 28.565 103.345 28.895 103.775 ;
        RECT 29.130 103.175 29.300 103.515 ;
        RECT 25.065 102.715 26.285 102.885 ;
        RECT 26.455 102.805 26.915 103.095 ;
        RECT 27.220 102.975 27.780 103.145 ;
        RECT 28.225 103.005 29.300 103.175 ;
        RECT 29.470 103.275 30.150 103.605 ;
        RECT 30.365 103.275 30.615 103.605 ;
        RECT 30.785 103.315 31.035 103.775 ;
        RECT 27.610 102.835 27.780 102.975 ;
        RECT 26.455 102.795 27.420 102.805 ;
        RECT 26.115 102.625 26.285 102.715 ;
        RECT 26.745 102.635 27.420 102.795 ;
        RECT 24.725 102.425 25.070 102.435 ;
        RECT 23.040 102.215 25.070 102.425 ;
        RECT 21.930 101.225 22.220 101.950 ;
        RECT 22.445 101.875 24.210 102.045 ;
        RECT 22.700 101.225 22.870 101.695 ;
        RECT 23.040 101.395 23.370 101.875 ;
        RECT 23.540 101.225 23.710 101.695 ;
        RECT 23.880 101.395 24.210 101.875 ;
        RECT 24.380 101.225 24.550 102.035 ;
        RECT 24.745 101.960 25.070 102.215 ;
        RECT 24.750 101.605 25.070 101.960 ;
        RECT 25.240 102.175 25.780 102.545 ;
        RECT 26.115 102.455 26.520 102.625 ;
        RECT 25.240 101.775 25.480 102.175 ;
        RECT 25.960 102.005 26.180 102.285 ;
        RECT 25.650 101.835 26.180 102.005 ;
        RECT 25.650 101.605 25.820 101.835 ;
        RECT 26.350 101.675 26.520 102.455 ;
        RECT 26.690 101.845 27.040 102.465 ;
        RECT 27.210 101.845 27.420 102.635 ;
        RECT 27.610 102.665 29.110 102.835 ;
        RECT 27.610 101.975 27.780 102.665 ;
        RECT 29.470 102.495 29.640 103.275 ;
        RECT 30.445 103.145 30.615 103.275 ;
        RECT 27.950 102.325 29.640 102.495 ;
        RECT 29.810 102.715 30.275 103.105 ;
        RECT 30.445 102.975 30.840 103.145 ;
        RECT 27.950 102.145 28.120 102.325 ;
        RECT 24.750 101.435 25.820 101.605 ;
        RECT 25.990 101.225 26.180 101.665 ;
        RECT 26.350 101.395 27.300 101.675 ;
        RECT 27.610 101.585 27.870 101.975 ;
        RECT 28.290 101.905 29.080 102.155 ;
        RECT 27.520 101.415 27.870 101.585 ;
        RECT 28.080 101.225 28.410 101.685 ;
        RECT 29.285 101.615 29.455 102.325 ;
        RECT 29.810 102.125 29.980 102.715 ;
        RECT 29.625 101.905 29.980 102.125 ;
        RECT 30.150 101.905 30.500 102.525 ;
        RECT 30.670 101.615 30.840 102.975 ;
        RECT 31.205 102.805 31.530 103.590 ;
        RECT 31.010 101.755 31.470 102.805 ;
        RECT 29.285 101.445 30.140 101.615 ;
        RECT 30.345 101.445 30.840 101.615 ;
        RECT 31.010 101.225 31.340 101.585 ;
        RECT 31.700 101.485 31.870 103.605 ;
        RECT 32.040 103.275 32.370 103.775 ;
        RECT 32.540 103.105 32.795 103.605 ;
        RECT 32.045 102.935 32.795 103.105 ;
        RECT 32.045 101.945 32.275 102.935 ;
        RECT 32.445 102.115 32.795 102.765 ;
        RECT 32.970 102.685 34.640 103.775 ;
        RECT 32.970 102.165 33.720 102.685 ;
        RECT 34.810 102.610 35.100 103.775 ;
        RECT 35.270 102.685 36.940 103.775 ;
        RECT 37.420 102.935 37.590 103.775 ;
        RECT 37.800 102.765 38.050 103.605 ;
        RECT 38.260 102.935 38.430 103.775 ;
        RECT 38.600 102.765 38.890 103.605 ;
        RECT 33.890 101.995 34.640 102.515 ;
        RECT 35.270 102.165 36.020 102.685 ;
        RECT 37.165 102.595 38.890 102.765 ;
        RECT 39.100 102.715 39.270 103.775 ;
        RECT 39.565 103.395 39.895 103.775 ;
        RECT 40.075 103.225 40.245 103.515 ;
        RECT 40.415 103.315 40.665 103.775 ;
        RECT 39.445 103.055 40.245 103.225 ;
        RECT 40.835 103.265 41.705 103.605 ;
        RECT 36.190 101.995 36.940 102.515 ;
        RECT 32.045 101.775 32.795 101.945 ;
        RECT 32.040 101.225 32.370 101.605 ;
        RECT 32.540 101.485 32.795 101.775 ;
        RECT 32.970 101.225 34.640 101.995 ;
        RECT 34.810 101.225 35.100 101.950 ;
        RECT 35.270 101.225 36.940 101.995 ;
        RECT 37.165 102.045 37.575 102.595 ;
        RECT 39.445 102.435 39.615 103.055 ;
        RECT 40.835 102.885 41.005 103.265 ;
        RECT 41.940 103.145 42.110 103.605 ;
        RECT 42.280 103.315 42.650 103.775 ;
        RECT 42.945 103.175 43.115 103.515 ;
        RECT 43.285 103.345 43.615 103.775 ;
        RECT 43.850 103.175 44.020 103.515 ;
        RECT 39.785 102.715 41.005 102.885 ;
        RECT 41.175 102.805 41.635 103.095 ;
        RECT 41.940 102.975 42.500 103.145 ;
        RECT 42.945 103.005 44.020 103.175 ;
        RECT 44.190 103.275 44.870 103.605 ;
        RECT 45.085 103.275 45.335 103.605 ;
        RECT 45.505 103.315 45.755 103.775 ;
        RECT 42.330 102.835 42.500 102.975 ;
        RECT 41.175 102.795 42.140 102.805 ;
        RECT 40.835 102.625 41.005 102.715 ;
        RECT 41.465 102.635 42.140 102.795 ;
        RECT 39.445 102.425 39.790 102.435 ;
        RECT 37.760 102.215 39.790 102.425 ;
        RECT 37.165 101.875 38.930 102.045 ;
        RECT 37.420 101.225 37.590 101.695 ;
        RECT 37.760 101.395 38.090 101.875 ;
        RECT 38.260 101.225 38.430 101.695 ;
        RECT 38.600 101.395 38.930 101.875 ;
        RECT 39.100 101.225 39.270 102.035 ;
        RECT 39.465 101.960 39.790 102.215 ;
        RECT 39.470 101.605 39.790 101.960 ;
        RECT 39.960 102.175 40.500 102.545 ;
        RECT 40.835 102.455 41.240 102.625 ;
        RECT 39.960 101.775 40.200 102.175 ;
        RECT 40.680 102.005 40.900 102.285 ;
        RECT 40.370 101.835 40.900 102.005 ;
        RECT 40.370 101.605 40.540 101.835 ;
        RECT 41.070 101.675 41.240 102.455 ;
        RECT 41.410 101.845 41.760 102.465 ;
        RECT 41.930 101.845 42.140 102.635 ;
        RECT 42.330 102.665 43.830 102.835 ;
        RECT 42.330 101.975 42.500 102.665 ;
        RECT 44.190 102.495 44.360 103.275 ;
        RECT 45.165 103.145 45.335 103.275 ;
        RECT 42.670 102.325 44.360 102.495 ;
        RECT 44.530 102.715 44.995 103.105 ;
        RECT 45.165 102.975 45.560 103.145 ;
        RECT 42.670 102.145 42.840 102.325 ;
        RECT 39.470 101.435 40.540 101.605 ;
        RECT 40.710 101.225 40.900 101.665 ;
        RECT 41.070 101.395 42.020 101.675 ;
        RECT 42.330 101.585 42.590 101.975 ;
        RECT 43.010 101.905 43.800 102.155 ;
        RECT 42.240 101.415 42.590 101.585 ;
        RECT 42.800 101.225 43.130 101.685 ;
        RECT 44.005 101.615 44.175 102.325 ;
        RECT 44.530 102.125 44.700 102.715 ;
        RECT 44.345 101.905 44.700 102.125 ;
        RECT 44.870 101.905 45.220 102.525 ;
        RECT 45.390 101.615 45.560 102.975 ;
        RECT 45.925 102.805 46.250 103.590 ;
        RECT 45.730 101.755 46.190 102.805 ;
        RECT 44.005 101.445 44.860 101.615 ;
        RECT 45.065 101.445 45.560 101.615 ;
        RECT 45.730 101.225 46.060 101.585 ;
        RECT 46.420 101.485 46.590 103.605 ;
        RECT 46.760 103.275 47.090 103.775 ;
        RECT 47.260 103.105 47.515 103.605 ;
        RECT 46.765 102.935 47.515 103.105 ;
        RECT 46.765 101.945 46.995 102.935 ;
        RECT 47.165 102.115 47.515 102.765 ;
        RECT 47.690 102.610 47.980 103.775 ;
        RECT 48.150 102.685 49.820 103.775 ;
        RECT 49.995 103.340 55.340 103.775 ;
        RECT 48.150 102.165 48.900 102.685 ;
        RECT 49.070 101.995 49.820 102.515 ;
        RECT 51.585 102.090 51.935 103.340 ;
        RECT 55.570 102.635 55.780 103.775 ;
        RECT 55.950 102.625 56.280 103.605 ;
        RECT 56.450 102.635 56.680 103.775 ;
        RECT 56.980 102.845 57.150 103.605 ;
        RECT 57.330 103.015 57.660 103.775 ;
        RECT 56.980 102.675 57.645 102.845 ;
        RECT 57.830 102.700 58.100 103.605 ;
        RECT 46.765 101.775 47.515 101.945 ;
        RECT 46.760 101.225 47.090 101.605 ;
        RECT 47.260 101.485 47.515 101.775 ;
        RECT 47.690 101.225 47.980 101.950 ;
        RECT 48.150 101.225 49.820 101.995 ;
        RECT 53.415 101.770 53.755 102.600 ;
        RECT 49.995 101.225 55.340 101.770 ;
        RECT 55.570 101.225 55.780 102.045 ;
        RECT 55.950 102.025 56.200 102.625 ;
        RECT 57.475 102.530 57.645 102.675 ;
        RECT 56.370 102.215 56.700 102.465 ;
        RECT 56.910 102.125 57.240 102.495 ;
        RECT 57.475 102.200 57.760 102.530 ;
        RECT 55.950 101.395 56.280 102.025 ;
        RECT 56.450 101.225 56.680 102.045 ;
        RECT 57.475 101.945 57.645 102.200 ;
        RECT 56.980 101.775 57.645 101.945 ;
        RECT 57.930 101.900 58.100 102.700 ;
        RECT 59.230 102.635 59.460 103.775 ;
        RECT 59.630 102.625 59.960 103.605 ;
        RECT 60.130 102.635 60.340 103.775 ;
        RECT 59.210 102.215 59.540 102.465 ;
        RECT 56.980 101.395 57.150 101.775 ;
        RECT 57.330 101.225 57.660 101.605 ;
        RECT 57.840 101.395 58.100 101.900 ;
        RECT 59.230 101.225 59.460 102.045 ;
        RECT 59.710 102.025 59.960 102.625 ;
        RECT 60.570 102.610 60.860 103.775 ;
        RECT 61.490 102.685 65.000 103.775 ;
        RECT 65.175 103.340 70.520 103.775 ;
        RECT 61.490 102.165 63.180 102.685 ;
        RECT 59.630 101.395 59.960 102.025 ;
        RECT 60.130 101.225 60.340 102.045 ;
        RECT 63.350 101.995 65.000 102.515 ;
        RECT 66.765 102.090 67.115 103.340 ;
        RECT 70.750 102.635 70.960 103.775 ;
        RECT 71.130 102.625 71.460 103.605 ;
        RECT 71.630 102.635 71.860 103.775 ;
        RECT 72.110 102.635 72.340 103.775 ;
        RECT 72.510 102.625 72.840 103.605 ;
        RECT 73.010 102.635 73.220 103.775 ;
        RECT 60.570 101.225 60.860 101.950 ;
        RECT 61.490 101.225 65.000 101.995 ;
        RECT 68.595 101.770 68.935 102.600 ;
        RECT 65.175 101.225 70.520 101.770 ;
        RECT 70.750 101.225 70.960 102.045 ;
        RECT 71.130 102.025 71.380 102.625 ;
        RECT 71.550 102.215 71.880 102.465 ;
        RECT 72.090 102.215 72.420 102.465 ;
        RECT 71.130 101.395 71.460 102.025 ;
        RECT 71.630 101.225 71.860 102.045 ;
        RECT 72.110 101.225 72.340 102.045 ;
        RECT 72.590 102.025 72.840 102.625 ;
        RECT 73.450 102.610 73.740 103.775 ;
        RECT 74.220 102.935 74.390 103.775 ;
        RECT 74.600 102.765 74.850 103.605 ;
        RECT 75.060 102.935 75.230 103.775 ;
        RECT 75.400 102.765 75.690 103.605 ;
        RECT 73.965 102.595 75.690 102.765 ;
        RECT 75.900 102.715 76.070 103.775 ;
        RECT 76.365 103.395 76.695 103.775 ;
        RECT 76.875 103.225 77.045 103.515 ;
        RECT 77.215 103.315 77.465 103.775 ;
        RECT 76.245 103.055 77.045 103.225 ;
        RECT 77.635 103.265 78.505 103.605 ;
        RECT 73.965 102.045 74.375 102.595 ;
        RECT 76.245 102.435 76.415 103.055 ;
        RECT 77.635 102.885 77.805 103.265 ;
        RECT 78.740 103.145 78.910 103.605 ;
        RECT 79.080 103.315 79.450 103.775 ;
        RECT 79.745 103.175 79.915 103.515 ;
        RECT 80.085 103.345 80.415 103.775 ;
        RECT 80.650 103.175 80.820 103.515 ;
        RECT 76.585 102.715 77.805 102.885 ;
        RECT 77.975 102.805 78.435 103.095 ;
        RECT 78.740 102.975 79.300 103.145 ;
        RECT 79.745 103.005 80.820 103.175 ;
        RECT 80.990 103.275 81.670 103.605 ;
        RECT 81.885 103.275 82.135 103.605 ;
        RECT 82.305 103.315 82.555 103.775 ;
        RECT 79.130 102.835 79.300 102.975 ;
        RECT 77.975 102.795 78.940 102.805 ;
        RECT 77.635 102.625 77.805 102.715 ;
        RECT 78.265 102.635 78.940 102.795 ;
        RECT 76.245 102.425 76.590 102.435 ;
        RECT 74.560 102.215 76.590 102.425 ;
        RECT 72.510 101.395 72.840 102.025 ;
        RECT 73.010 101.225 73.220 102.045 ;
        RECT 73.450 101.225 73.740 101.950 ;
        RECT 73.965 101.875 75.730 102.045 ;
        RECT 74.220 101.225 74.390 101.695 ;
        RECT 74.560 101.395 74.890 101.875 ;
        RECT 75.060 101.225 75.230 101.695 ;
        RECT 75.400 101.395 75.730 101.875 ;
        RECT 75.900 101.225 76.070 102.035 ;
        RECT 76.265 101.960 76.590 102.215 ;
        RECT 76.270 101.605 76.590 101.960 ;
        RECT 76.760 102.175 77.300 102.545 ;
        RECT 77.635 102.455 78.040 102.625 ;
        RECT 76.760 101.775 77.000 102.175 ;
        RECT 77.480 102.005 77.700 102.285 ;
        RECT 77.170 101.835 77.700 102.005 ;
        RECT 77.170 101.605 77.340 101.835 ;
        RECT 77.870 101.675 78.040 102.455 ;
        RECT 78.210 101.845 78.560 102.465 ;
        RECT 78.730 101.845 78.940 102.635 ;
        RECT 79.130 102.665 80.630 102.835 ;
        RECT 79.130 101.975 79.300 102.665 ;
        RECT 80.990 102.495 81.160 103.275 ;
        RECT 81.965 103.145 82.135 103.275 ;
        RECT 79.470 102.325 81.160 102.495 ;
        RECT 81.330 102.715 81.795 103.105 ;
        RECT 81.965 102.975 82.360 103.145 ;
        RECT 79.470 102.145 79.640 102.325 ;
        RECT 76.270 101.435 77.340 101.605 ;
        RECT 77.510 101.225 77.700 101.665 ;
        RECT 77.870 101.395 78.820 101.675 ;
        RECT 79.130 101.585 79.390 101.975 ;
        RECT 79.810 101.905 80.600 102.155 ;
        RECT 79.040 101.415 79.390 101.585 ;
        RECT 79.600 101.225 79.930 101.685 ;
        RECT 80.805 101.615 80.975 102.325 ;
        RECT 81.330 102.125 81.500 102.715 ;
        RECT 81.145 101.905 81.500 102.125 ;
        RECT 81.670 101.905 82.020 102.525 ;
        RECT 82.190 101.615 82.360 102.975 ;
        RECT 82.725 102.805 83.050 103.590 ;
        RECT 82.530 101.755 82.990 102.805 ;
        RECT 80.805 101.445 81.660 101.615 ;
        RECT 81.865 101.445 82.360 101.615 ;
        RECT 82.530 101.225 82.860 101.585 ;
        RECT 83.220 101.485 83.390 103.605 ;
        RECT 83.560 103.275 83.890 103.775 ;
        RECT 84.060 103.105 84.315 103.605 ;
        RECT 83.565 102.935 84.315 103.105 ;
        RECT 83.565 101.945 83.795 102.935 ;
        RECT 83.965 102.115 84.315 102.765 ;
        RECT 84.550 102.635 84.760 103.775 ;
        RECT 84.930 102.625 85.260 103.605 ;
        RECT 85.430 102.635 85.660 103.775 ;
        RECT 83.565 101.775 84.315 101.945 ;
        RECT 83.560 101.225 83.890 101.605 ;
        RECT 84.060 101.485 84.315 101.775 ;
        RECT 84.550 101.225 84.760 102.045 ;
        RECT 84.930 102.025 85.180 102.625 ;
        RECT 86.330 102.610 86.620 103.775 ;
        RECT 86.830 102.635 87.060 103.775 ;
        RECT 87.230 102.625 87.560 103.605 ;
        RECT 87.730 102.635 87.940 103.775 ;
        RECT 88.940 102.935 89.110 103.775 ;
        RECT 89.320 102.765 89.570 103.605 ;
        RECT 89.780 102.935 89.950 103.775 ;
        RECT 90.120 102.765 90.410 103.605 ;
        RECT 85.350 102.215 85.680 102.465 ;
        RECT 86.810 102.215 87.140 102.465 ;
        RECT 84.930 101.395 85.260 102.025 ;
        RECT 85.430 101.225 85.660 102.045 ;
        RECT 86.330 101.225 86.620 101.950 ;
        RECT 86.830 101.225 87.060 102.045 ;
        RECT 87.310 102.025 87.560 102.625 ;
        RECT 88.685 102.595 90.410 102.765 ;
        RECT 90.620 102.715 90.790 103.775 ;
        RECT 91.085 103.395 91.415 103.775 ;
        RECT 91.595 103.225 91.765 103.515 ;
        RECT 91.935 103.315 92.185 103.775 ;
        RECT 90.965 103.055 91.765 103.225 ;
        RECT 92.355 103.265 93.225 103.605 ;
        RECT 88.685 102.045 89.095 102.595 ;
        RECT 90.965 102.435 91.135 103.055 ;
        RECT 92.355 102.885 92.525 103.265 ;
        RECT 93.460 103.145 93.630 103.605 ;
        RECT 93.800 103.315 94.170 103.775 ;
        RECT 94.465 103.175 94.635 103.515 ;
        RECT 94.805 103.345 95.135 103.775 ;
        RECT 95.370 103.175 95.540 103.515 ;
        RECT 91.305 102.715 92.525 102.885 ;
        RECT 92.695 102.805 93.155 103.095 ;
        RECT 93.460 102.975 94.020 103.145 ;
        RECT 94.465 103.005 95.540 103.175 ;
        RECT 95.710 103.275 96.390 103.605 ;
        RECT 96.605 103.275 96.855 103.605 ;
        RECT 97.025 103.315 97.275 103.775 ;
        RECT 93.850 102.835 94.020 102.975 ;
        RECT 92.695 102.795 93.660 102.805 ;
        RECT 92.355 102.625 92.525 102.715 ;
        RECT 92.985 102.635 93.660 102.795 ;
        RECT 90.965 102.425 91.310 102.435 ;
        RECT 89.280 102.215 91.310 102.425 ;
        RECT 87.230 101.395 87.560 102.025 ;
        RECT 87.730 101.225 87.940 102.045 ;
        RECT 88.685 101.875 90.450 102.045 ;
        RECT 88.940 101.225 89.110 101.695 ;
        RECT 89.280 101.395 89.610 101.875 ;
        RECT 89.780 101.225 89.950 101.695 ;
        RECT 90.120 101.395 90.450 101.875 ;
        RECT 90.620 101.225 90.790 102.035 ;
        RECT 90.985 101.960 91.310 102.215 ;
        RECT 90.990 101.605 91.310 101.960 ;
        RECT 91.480 102.175 92.020 102.545 ;
        RECT 92.355 102.455 92.760 102.625 ;
        RECT 91.480 101.775 91.720 102.175 ;
        RECT 92.200 102.005 92.420 102.285 ;
        RECT 91.890 101.835 92.420 102.005 ;
        RECT 91.890 101.605 92.060 101.835 ;
        RECT 92.590 101.675 92.760 102.455 ;
        RECT 92.930 101.845 93.280 102.465 ;
        RECT 93.450 101.845 93.660 102.635 ;
        RECT 93.850 102.665 95.350 102.835 ;
        RECT 93.850 101.975 94.020 102.665 ;
        RECT 95.710 102.495 95.880 103.275 ;
        RECT 96.685 103.145 96.855 103.275 ;
        RECT 94.190 102.325 95.880 102.495 ;
        RECT 96.050 102.715 96.515 103.105 ;
        RECT 96.685 102.975 97.080 103.145 ;
        RECT 94.190 102.145 94.360 102.325 ;
        RECT 90.990 101.435 92.060 101.605 ;
        RECT 92.230 101.225 92.420 101.665 ;
        RECT 92.590 101.395 93.540 101.675 ;
        RECT 93.850 101.585 94.110 101.975 ;
        RECT 94.530 101.905 95.320 102.155 ;
        RECT 93.760 101.415 94.110 101.585 ;
        RECT 94.320 101.225 94.650 101.685 ;
        RECT 95.525 101.615 95.695 102.325 ;
        RECT 96.050 102.125 96.220 102.715 ;
        RECT 95.865 101.905 96.220 102.125 ;
        RECT 96.390 101.905 96.740 102.525 ;
        RECT 96.910 101.615 97.080 102.975 ;
        RECT 97.445 102.805 97.770 103.590 ;
        RECT 97.250 101.755 97.710 102.805 ;
        RECT 95.525 101.445 96.380 101.615 ;
        RECT 96.585 101.445 97.080 101.615 ;
        RECT 97.250 101.225 97.580 101.585 ;
        RECT 97.940 101.485 98.110 103.605 ;
        RECT 98.280 103.275 98.610 103.775 ;
        RECT 98.780 103.105 99.035 103.605 ;
        RECT 98.285 102.935 99.035 103.105 ;
        RECT 98.285 101.945 98.515 102.935 ;
        RECT 98.685 102.115 99.035 102.765 ;
        RECT 99.210 102.610 99.500 103.775 ;
        RECT 100.595 103.105 100.850 103.605 ;
        RECT 101.020 103.275 101.350 103.775 ;
        RECT 100.595 102.935 101.345 103.105 ;
        RECT 100.595 102.115 100.945 102.765 ;
        RECT 98.285 101.775 99.035 101.945 ;
        RECT 98.280 101.225 98.610 101.605 ;
        RECT 98.780 101.485 99.035 101.775 ;
        RECT 99.210 101.225 99.500 101.950 ;
        RECT 101.115 101.945 101.345 102.935 ;
        RECT 100.595 101.775 101.345 101.945 ;
        RECT 100.595 101.485 100.850 101.775 ;
        RECT 101.020 101.225 101.350 101.605 ;
        RECT 101.520 101.485 101.690 103.605 ;
        RECT 101.860 102.805 102.185 103.590 ;
        RECT 102.355 103.315 102.605 103.775 ;
        RECT 102.775 103.275 103.025 103.605 ;
        RECT 103.240 103.275 103.920 103.605 ;
        RECT 102.775 103.145 102.945 103.275 ;
        RECT 102.550 102.975 102.945 103.145 ;
        RECT 101.920 101.755 102.380 102.805 ;
        RECT 102.550 101.615 102.720 102.975 ;
        RECT 103.115 102.715 103.580 103.105 ;
        RECT 102.890 101.905 103.240 102.525 ;
        RECT 103.410 102.125 103.580 102.715 ;
        RECT 103.750 102.495 103.920 103.275 ;
        RECT 104.090 103.175 104.260 103.515 ;
        RECT 104.495 103.345 104.825 103.775 ;
        RECT 104.995 103.175 105.165 103.515 ;
        RECT 105.460 103.315 105.830 103.775 ;
        RECT 104.090 103.005 105.165 103.175 ;
        RECT 106.000 103.145 106.170 103.605 ;
        RECT 106.405 103.265 107.275 103.605 ;
        RECT 107.445 103.315 107.695 103.775 ;
        RECT 105.610 102.975 106.170 103.145 ;
        RECT 105.610 102.835 105.780 102.975 ;
        RECT 104.280 102.665 105.780 102.835 ;
        RECT 106.475 102.805 106.935 103.095 ;
        RECT 103.750 102.325 105.440 102.495 ;
        RECT 103.410 101.905 103.765 102.125 ;
        RECT 103.935 101.615 104.105 102.325 ;
        RECT 104.310 101.905 105.100 102.155 ;
        RECT 105.270 102.145 105.440 102.325 ;
        RECT 105.610 101.975 105.780 102.665 ;
        RECT 102.050 101.225 102.380 101.585 ;
        RECT 102.550 101.445 103.045 101.615 ;
        RECT 103.250 101.445 104.105 101.615 ;
        RECT 104.980 101.225 105.310 101.685 ;
        RECT 105.520 101.585 105.780 101.975 ;
        RECT 105.970 102.795 106.935 102.805 ;
        RECT 107.105 102.885 107.275 103.265 ;
        RECT 107.865 103.225 108.035 103.515 ;
        RECT 108.215 103.395 108.545 103.775 ;
        RECT 107.865 103.055 108.665 103.225 ;
        RECT 105.970 102.635 106.645 102.795 ;
        RECT 107.105 102.715 108.325 102.885 ;
        RECT 105.970 101.845 106.180 102.635 ;
        RECT 107.105 102.625 107.275 102.715 ;
        RECT 106.350 101.845 106.700 102.465 ;
        RECT 106.870 102.455 107.275 102.625 ;
        RECT 106.870 101.675 107.040 102.455 ;
        RECT 107.210 102.005 107.430 102.285 ;
        RECT 107.610 102.175 108.150 102.545 ;
        RECT 108.495 102.435 108.665 103.055 ;
        RECT 108.840 102.715 109.010 103.775 ;
        RECT 109.220 102.765 109.510 103.605 ;
        RECT 109.680 102.935 109.850 103.775 ;
        RECT 110.060 102.765 110.310 103.605 ;
        RECT 110.520 102.935 110.690 103.775 ;
        RECT 109.220 102.595 110.945 102.765 ;
        RECT 107.210 101.835 107.740 102.005 ;
        RECT 105.520 101.415 105.870 101.585 ;
        RECT 106.090 101.395 107.040 101.675 ;
        RECT 107.210 101.225 107.400 101.665 ;
        RECT 107.570 101.605 107.740 101.835 ;
        RECT 107.910 101.775 108.150 102.175 ;
        RECT 108.320 102.425 108.665 102.435 ;
        RECT 108.320 102.215 110.350 102.425 ;
        RECT 108.320 101.960 108.645 102.215 ;
        RECT 110.535 102.045 110.945 102.595 ;
        RECT 111.170 102.685 112.380 103.775 ;
        RECT 111.170 102.145 111.690 102.685 ;
        RECT 108.320 101.605 108.640 101.960 ;
        RECT 107.570 101.435 108.640 101.605 ;
        RECT 108.840 101.225 109.010 102.035 ;
        RECT 109.180 101.875 110.945 102.045 ;
        RECT 111.860 101.975 112.380 102.515 ;
        RECT 109.180 101.395 109.510 101.875 ;
        RECT 109.680 101.225 109.850 101.695 ;
        RECT 110.020 101.395 110.350 101.875 ;
        RECT 110.520 101.225 110.690 101.695 ;
        RECT 111.170 101.225 112.380 101.975 ;
        RECT 18.165 101.055 112.465 101.225 ;
        RECT 19.165 66.070 30.165 66.940 ;
        RECT 19.165 54.930 20.835 66.070 ;
        RECT 21.465 65.555 26.465 65.725 ;
        RECT 21.235 55.300 21.405 65.340 ;
        RECT 26.525 55.300 26.695 65.340 ;
        RECT 27.095 54.930 27.265 66.070 ;
        RECT 27.895 65.555 28.895 65.725 ;
        RECT 27.665 55.300 27.835 65.340 ;
        RECT 28.955 55.300 29.125 65.340 ;
        RECT 29.525 54.930 30.165 66.070 ;
        RECT 19.165 52.860 30.165 54.930 ;
        RECT 19.165 49.370 21.005 52.860 ;
        RECT 22.765 52.780 30.165 52.860 ;
        RECT 21.635 52.350 22.135 52.520 ;
        RECT 21.405 50.095 21.575 52.135 ;
        RECT 22.195 50.095 22.365 52.135 ;
        RECT 21.635 49.710 22.135 49.880 ;
        RECT 22.765 49.370 25.085 52.780 ;
        RECT 25.715 52.270 26.215 52.440 ;
        RECT 19.165 48.650 25.085 49.370 ;
        RECT 19.135 48.040 23.045 48.260 ;
        RECT 19.135 45.640 20.855 48.040 ;
        RECT 21.485 47.530 21.985 47.700 ;
        RECT 21.255 46.320 21.425 47.360 ;
        RECT 22.045 46.320 22.215 47.360 ;
        RECT 21.485 45.980 21.985 46.150 ;
        RECT 22.615 45.640 23.045 48.040 ;
        RECT 24.025 46.290 25.085 48.650 ;
        RECT 25.485 47.015 25.655 52.055 ;
        RECT 26.275 47.015 26.445 52.055 ;
        RECT 25.715 46.630 26.215 46.800 ;
        RECT 26.845 46.290 27.015 52.780 ;
        RECT 27.645 52.270 28.145 52.440 ;
        RECT 27.415 47.015 27.585 52.055 ;
        RECT 28.205 47.015 28.375 52.055 ;
        RECT 27.645 46.630 28.145 46.800 ;
        RECT 28.775 46.290 30.165 52.780 ;
        RECT 30.365 66.080 41.365 66.950 ;
        RECT 30.365 54.940 32.035 66.080 ;
        RECT 32.665 65.565 37.665 65.735 ;
        RECT 32.435 55.310 32.605 65.350 ;
        RECT 37.725 55.310 37.895 65.350 ;
        RECT 38.295 54.940 38.465 66.080 ;
        RECT 39.095 65.565 40.095 65.735 ;
        RECT 38.865 55.310 39.035 65.350 ;
        RECT 40.155 55.310 40.325 65.350 ;
        RECT 40.725 54.940 41.365 66.080 ;
        RECT 30.365 52.870 41.365 54.940 ;
        RECT 30.365 49.380 32.205 52.870 ;
        RECT 33.965 52.790 41.365 52.870 ;
        RECT 32.835 52.360 33.335 52.530 ;
        RECT 32.605 50.105 32.775 52.145 ;
        RECT 33.395 50.105 33.565 52.145 ;
        RECT 32.835 49.720 33.335 49.890 ;
        RECT 33.965 49.380 36.285 52.790 ;
        RECT 36.915 52.280 37.415 52.450 ;
        RECT 30.365 48.660 36.285 49.380 ;
        RECT 24.025 45.800 30.165 46.290 ;
        RECT 30.335 48.050 34.245 48.270 ;
        RECT 19.135 45.370 23.045 45.640 ;
        RECT 30.335 45.650 32.055 48.050 ;
        RECT 32.685 47.540 33.185 47.710 ;
        RECT 32.455 46.330 32.625 47.370 ;
        RECT 33.245 46.330 33.415 47.370 ;
        RECT 32.685 45.990 33.185 46.160 ;
        RECT 33.815 45.650 34.245 48.050 ;
        RECT 35.225 46.300 36.285 48.660 ;
        RECT 36.685 47.025 36.855 52.065 ;
        RECT 37.475 47.025 37.645 52.065 ;
        RECT 36.915 46.640 37.415 46.810 ;
        RECT 38.045 46.300 38.215 52.790 ;
        RECT 38.845 52.280 39.345 52.450 ;
        RECT 38.615 47.025 38.785 52.065 ;
        RECT 39.405 47.025 39.575 52.065 ;
        RECT 38.845 46.640 39.345 46.810 ;
        RECT 39.975 46.300 41.365 52.790 ;
        RECT 41.585 66.050 52.585 66.920 ;
        RECT 41.585 54.910 43.255 66.050 ;
        RECT 43.885 65.535 48.885 65.705 ;
        RECT 43.655 55.280 43.825 65.320 ;
        RECT 48.945 55.280 49.115 65.320 ;
        RECT 49.515 54.910 49.685 66.050 ;
        RECT 50.315 65.535 51.315 65.705 ;
        RECT 50.085 55.280 50.255 65.320 ;
        RECT 51.375 55.280 51.545 65.320 ;
        RECT 51.945 54.910 52.585 66.050 ;
        RECT 41.585 52.840 52.585 54.910 ;
        RECT 41.585 49.350 43.425 52.840 ;
        RECT 45.185 52.760 52.585 52.840 ;
        RECT 44.055 52.330 44.555 52.500 ;
        RECT 43.825 50.075 43.995 52.115 ;
        RECT 44.615 50.075 44.785 52.115 ;
        RECT 44.055 49.690 44.555 49.860 ;
        RECT 45.185 49.350 47.505 52.760 ;
        RECT 48.135 52.250 48.635 52.420 ;
        RECT 41.585 48.630 47.505 49.350 ;
        RECT 35.225 45.810 41.365 46.300 ;
        RECT 41.555 48.020 45.465 48.240 ;
        RECT 30.335 45.380 34.245 45.650 ;
        RECT 41.555 45.620 43.275 48.020 ;
        RECT 43.905 47.510 44.405 47.680 ;
        RECT 43.675 46.300 43.845 47.340 ;
        RECT 44.465 46.300 44.635 47.340 ;
        RECT 43.905 45.960 44.405 46.130 ;
        RECT 45.035 45.620 45.465 48.020 ;
        RECT 46.445 46.270 47.505 48.630 ;
        RECT 47.905 46.995 48.075 52.035 ;
        RECT 48.695 46.995 48.865 52.035 ;
        RECT 48.135 46.610 48.635 46.780 ;
        RECT 49.265 46.270 49.435 52.760 ;
        RECT 50.065 52.250 50.565 52.420 ;
        RECT 49.835 46.995 50.005 52.035 ;
        RECT 50.625 46.995 50.795 52.035 ;
        RECT 50.065 46.610 50.565 46.780 ;
        RECT 51.195 46.270 52.585 52.760 ;
        RECT 52.835 66.030 63.835 66.900 ;
        RECT 52.835 54.890 54.505 66.030 ;
        RECT 55.135 65.515 60.135 65.685 ;
        RECT 54.905 55.260 55.075 65.300 ;
        RECT 60.195 55.260 60.365 65.300 ;
        RECT 60.765 54.890 60.935 66.030 ;
        RECT 61.565 65.515 62.565 65.685 ;
        RECT 61.335 55.260 61.505 65.300 ;
        RECT 62.625 55.260 62.795 65.300 ;
        RECT 63.195 54.890 63.835 66.030 ;
        RECT 52.835 52.820 63.835 54.890 ;
        RECT 52.835 49.330 54.675 52.820 ;
        RECT 56.435 52.740 63.835 52.820 ;
        RECT 55.305 52.310 55.805 52.480 ;
        RECT 55.075 50.055 55.245 52.095 ;
        RECT 55.865 50.055 56.035 52.095 ;
        RECT 55.305 49.670 55.805 49.840 ;
        RECT 56.435 49.330 58.755 52.740 ;
        RECT 59.385 52.230 59.885 52.400 ;
        RECT 52.835 48.610 58.755 49.330 ;
        RECT 46.445 45.780 52.585 46.270 ;
        RECT 52.805 48.000 56.715 48.220 ;
        RECT 41.555 45.350 45.465 45.620 ;
        RECT 52.805 45.600 54.525 48.000 ;
        RECT 55.155 47.490 55.655 47.660 ;
        RECT 54.925 46.280 55.095 47.320 ;
        RECT 55.715 46.280 55.885 47.320 ;
        RECT 55.155 45.940 55.655 46.110 ;
        RECT 56.285 45.600 56.715 48.000 ;
        RECT 57.695 46.250 58.755 48.610 ;
        RECT 59.155 46.975 59.325 52.015 ;
        RECT 59.945 46.975 60.115 52.015 ;
        RECT 59.385 46.590 59.885 46.760 ;
        RECT 60.515 46.250 60.685 52.740 ;
        RECT 61.315 52.230 61.815 52.400 ;
        RECT 61.085 46.975 61.255 52.015 ;
        RECT 61.875 46.975 62.045 52.015 ;
        RECT 61.315 46.590 61.815 46.760 ;
        RECT 62.445 46.250 63.835 52.740 ;
        RECT 64.055 66.020 75.055 66.890 ;
        RECT 64.055 54.880 65.725 66.020 ;
        RECT 66.355 65.505 71.355 65.675 ;
        RECT 66.125 55.250 66.295 65.290 ;
        RECT 71.415 55.250 71.585 65.290 ;
        RECT 71.985 54.880 72.155 66.020 ;
        RECT 72.785 65.505 73.785 65.675 ;
        RECT 72.555 55.250 72.725 65.290 ;
        RECT 73.845 55.250 74.015 65.290 ;
        RECT 74.415 54.880 75.055 66.020 ;
        RECT 64.055 52.810 75.055 54.880 ;
        RECT 64.055 49.320 65.895 52.810 ;
        RECT 67.655 52.730 75.055 52.810 ;
        RECT 66.525 52.300 67.025 52.470 ;
        RECT 66.295 50.045 66.465 52.085 ;
        RECT 67.085 50.045 67.255 52.085 ;
        RECT 66.525 49.660 67.025 49.830 ;
        RECT 67.655 49.320 69.975 52.730 ;
        RECT 70.605 52.220 71.105 52.390 ;
        RECT 64.055 48.600 69.975 49.320 ;
        RECT 57.695 45.760 63.835 46.250 ;
        RECT 64.025 47.990 67.935 48.210 ;
        RECT 52.805 45.330 56.715 45.600 ;
        RECT 64.025 45.590 65.745 47.990 ;
        RECT 66.375 47.480 66.875 47.650 ;
        RECT 66.145 46.270 66.315 47.310 ;
        RECT 66.935 46.270 67.105 47.310 ;
        RECT 66.375 45.930 66.875 46.100 ;
        RECT 67.505 45.590 67.935 47.990 ;
        RECT 68.915 46.240 69.975 48.600 ;
        RECT 70.375 46.965 70.545 52.005 ;
        RECT 71.165 46.965 71.335 52.005 ;
        RECT 70.605 46.580 71.105 46.750 ;
        RECT 71.735 46.240 71.905 52.730 ;
        RECT 72.535 52.220 73.035 52.390 ;
        RECT 72.305 46.965 72.475 52.005 ;
        RECT 73.095 46.965 73.265 52.005 ;
        RECT 72.535 46.580 73.035 46.750 ;
        RECT 73.665 46.240 75.055 52.730 ;
        RECT 75.295 66.010 86.295 66.880 ;
        RECT 75.295 54.870 76.965 66.010 ;
        RECT 77.595 65.495 82.595 65.665 ;
        RECT 77.365 55.240 77.535 65.280 ;
        RECT 82.655 55.240 82.825 65.280 ;
        RECT 83.225 54.870 83.395 66.010 ;
        RECT 84.025 65.495 85.025 65.665 ;
        RECT 83.795 55.240 83.965 65.280 ;
        RECT 85.085 55.240 85.255 65.280 ;
        RECT 85.655 54.870 86.295 66.010 ;
        RECT 75.295 52.800 86.295 54.870 ;
        RECT 75.295 49.310 77.135 52.800 ;
        RECT 78.895 52.720 86.295 52.800 ;
        RECT 77.765 52.290 78.265 52.460 ;
        RECT 77.535 50.035 77.705 52.075 ;
        RECT 78.325 50.035 78.495 52.075 ;
        RECT 77.765 49.650 78.265 49.820 ;
        RECT 78.895 49.310 81.215 52.720 ;
        RECT 81.845 52.210 82.345 52.380 ;
        RECT 75.295 48.590 81.215 49.310 ;
        RECT 68.915 45.750 75.055 46.240 ;
        RECT 75.265 47.980 79.175 48.200 ;
        RECT 64.025 45.320 67.935 45.590 ;
        RECT 75.265 45.580 76.985 47.980 ;
        RECT 77.615 47.470 78.115 47.640 ;
        RECT 77.385 46.260 77.555 47.300 ;
        RECT 78.175 46.260 78.345 47.300 ;
        RECT 77.615 45.920 78.115 46.090 ;
        RECT 78.745 45.580 79.175 47.980 ;
        RECT 80.155 46.230 81.215 48.590 ;
        RECT 81.615 46.955 81.785 51.995 ;
        RECT 82.405 46.955 82.575 51.995 ;
        RECT 81.845 46.570 82.345 46.740 ;
        RECT 82.975 46.230 83.145 52.720 ;
        RECT 83.775 52.210 84.275 52.380 ;
        RECT 83.545 46.955 83.715 51.995 ;
        RECT 84.335 46.955 84.505 51.995 ;
        RECT 83.775 46.570 84.275 46.740 ;
        RECT 84.905 46.230 86.295 52.720 ;
        RECT 86.545 66.020 97.545 66.890 ;
        RECT 131.125 66.880 140.025 66.890 ;
        RECT 86.545 54.880 88.215 66.020 ;
        RECT 88.845 65.505 93.845 65.675 ;
        RECT 88.615 55.250 88.785 65.290 ;
        RECT 93.905 55.250 94.075 65.290 ;
        RECT 94.475 54.880 94.645 66.020 ;
        RECT 95.275 65.505 96.275 65.675 ;
        RECT 95.045 55.250 95.215 65.290 ;
        RECT 96.335 55.250 96.505 65.290 ;
        RECT 96.905 54.880 97.545 66.020 ;
        RECT 86.545 52.810 97.545 54.880 ;
        RECT 86.545 49.320 88.385 52.810 ;
        RECT 90.145 52.730 97.545 52.810 ;
        RECT 89.015 52.300 89.515 52.470 ;
        RECT 88.785 50.045 88.955 52.085 ;
        RECT 89.575 50.045 89.745 52.085 ;
        RECT 89.015 49.660 89.515 49.830 ;
        RECT 90.145 49.320 92.465 52.730 ;
        RECT 93.095 52.220 93.595 52.390 ;
        RECT 86.545 48.600 92.465 49.320 ;
        RECT 80.155 45.740 86.295 46.230 ;
        RECT 86.515 47.990 90.425 48.210 ;
        RECT 75.265 45.310 79.175 45.580 ;
        RECT 86.515 45.590 88.235 47.990 ;
        RECT 88.865 47.480 89.365 47.650 ;
        RECT 88.635 46.270 88.805 47.310 ;
        RECT 89.425 46.270 89.595 47.310 ;
        RECT 88.865 45.930 89.365 46.100 ;
        RECT 89.995 45.590 90.425 47.990 ;
        RECT 91.405 46.240 92.465 48.600 ;
        RECT 92.865 46.965 93.035 52.005 ;
        RECT 93.655 46.965 93.825 52.005 ;
        RECT 93.095 46.580 93.595 46.750 ;
        RECT 94.225 46.240 94.395 52.730 ;
        RECT 95.025 52.220 95.525 52.390 ;
        RECT 94.795 46.965 94.965 52.005 ;
        RECT 95.585 46.965 95.755 52.005 ;
        RECT 95.025 46.580 95.525 46.750 ;
        RECT 96.155 46.240 97.545 52.730 ;
        RECT 97.825 66.010 108.825 66.880 ;
        RECT 97.825 54.870 99.495 66.010 ;
        RECT 100.125 65.495 105.125 65.665 ;
        RECT 99.895 55.240 100.065 65.280 ;
        RECT 105.185 55.240 105.355 65.280 ;
        RECT 105.755 54.870 105.925 66.010 ;
        RECT 106.555 65.495 107.555 65.665 ;
        RECT 106.325 55.240 106.495 65.280 ;
        RECT 107.615 55.240 107.785 65.280 ;
        RECT 108.185 54.870 108.825 66.010 ;
        RECT 97.825 52.800 108.825 54.870 ;
        RECT 97.825 49.310 99.665 52.800 ;
        RECT 101.425 52.720 108.825 52.800 ;
        RECT 100.295 52.290 100.795 52.460 ;
        RECT 100.065 50.035 100.235 52.075 ;
        RECT 100.855 50.035 101.025 52.075 ;
        RECT 100.295 49.650 100.795 49.820 ;
        RECT 101.425 49.310 103.745 52.720 ;
        RECT 104.375 52.210 104.875 52.380 ;
        RECT 97.825 48.590 103.745 49.310 ;
        RECT 91.405 45.750 97.545 46.240 ;
        RECT 97.795 47.980 101.705 48.200 ;
        RECT 86.515 45.320 90.425 45.590 ;
        RECT 97.795 45.580 99.515 47.980 ;
        RECT 100.145 47.470 100.645 47.640 ;
        RECT 99.915 46.260 100.085 47.300 ;
        RECT 100.705 46.260 100.875 47.300 ;
        RECT 100.145 45.920 100.645 46.090 ;
        RECT 101.275 45.580 101.705 47.980 ;
        RECT 102.685 46.230 103.745 48.590 ;
        RECT 104.145 46.955 104.315 51.995 ;
        RECT 104.935 46.955 105.105 51.995 ;
        RECT 104.375 46.570 104.875 46.740 ;
        RECT 105.505 46.230 105.675 52.720 ;
        RECT 106.305 52.210 106.805 52.380 ;
        RECT 106.075 46.955 106.245 51.995 ;
        RECT 106.865 46.955 107.035 51.995 ;
        RECT 106.305 46.570 106.805 46.740 ;
        RECT 107.435 46.230 108.825 52.720 ;
        RECT 109.095 66.010 120.095 66.880 ;
        RECT 109.095 54.870 110.765 66.010 ;
        RECT 111.395 65.495 116.395 65.665 ;
        RECT 111.165 55.240 111.335 65.280 ;
        RECT 116.455 55.240 116.625 65.280 ;
        RECT 117.025 54.870 117.195 66.010 ;
        RECT 117.825 65.495 118.825 65.665 ;
        RECT 117.595 55.240 117.765 65.280 ;
        RECT 118.885 55.240 119.055 65.280 ;
        RECT 119.455 54.870 120.095 66.010 ;
        RECT 109.095 52.800 120.095 54.870 ;
        RECT 109.095 49.310 110.935 52.800 ;
        RECT 112.695 52.720 120.095 52.800 ;
        RECT 111.565 52.290 112.065 52.460 ;
        RECT 111.335 50.035 111.505 52.075 ;
        RECT 112.125 50.035 112.295 52.075 ;
        RECT 111.565 49.650 112.065 49.820 ;
        RECT 112.695 49.310 115.015 52.720 ;
        RECT 115.645 52.210 116.145 52.380 ;
        RECT 109.095 48.590 115.015 49.310 ;
        RECT 102.685 45.740 108.825 46.230 ;
        RECT 109.065 47.980 112.975 48.200 ;
        RECT 97.795 45.310 101.705 45.580 ;
        RECT 109.065 45.580 110.785 47.980 ;
        RECT 111.415 47.470 111.915 47.640 ;
        RECT 111.185 46.260 111.355 47.300 ;
        RECT 111.975 46.260 112.145 47.300 ;
        RECT 111.415 45.920 111.915 46.090 ;
        RECT 112.545 45.580 112.975 47.980 ;
        RECT 113.955 46.230 115.015 48.590 ;
        RECT 115.415 46.955 115.585 51.995 ;
        RECT 116.205 46.955 116.375 51.995 ;
        RECT 115.645 46.570 116.145 46.740 ;
        RECT 116.775 46.230 116.945 52.720 ;
        RECT 117.575 52.210 118.075 52.380 ;
        RECT 117.345 46.955 117.515 51.995 ;
        RECT 118.135 46.955 118.305 51.995 ;
        RECT 117.575 46.570 118.075 46.740 ;
        RECT 118.705 46.230 120.095 52.720 ;
        RECT 120.345 66.010 140.025 66.880 ;
        RECT 120.345 54.870 122.015 66.010 ;
        RECT 122.645 65.495 127.645 65.665 ;
        RECT 122.415 55.240 122.585 65.280 ;
        RECT 127.705 55.240 127.875 65.280 ;
        RECT 128.275 54.870 128.445 66.010 ;
        RECT 130.705 65.980 140.025 66.010 ;
        RECT 129.075 65.495 130.075 65.665 ;
        RECT 128.845 55.240 129.015 65.280 ;
        RECT 130.135 55.240 130.305 65.280 ;
        RECT 130.705 54.870 132.765 65.980 ;
        RECT 133.395 65.465 138.395 65.635 ;
        RECT 133.165 55.210 133.335 65.250 ;
        RECT 138.455 55.210 138.625 65.250 ;
        RECT 120.345 54.840 132.765 54.870 ;
        RECT 139.025 54.840 140.025 65.980 ;
        RECT 120.345 54.720 140.025 54.840 ;
        RECT 120.345 53.550 140.035 54.720 ;
        RECT 120.345 52.800 131.345 53.550 ;
        RECT 120.345 49.310 122.185 52.800 ;
        RECT 123.945 52.720 131.345 52.800 ;
        RECT 122.815 52.290 123.315 52.460 ;
        RECT 122.585 50.035 122.755 52.075 ;
        RECT 123.375 50.035 123.545 52.075 ;
        RECT 122.815 49.650 123.315 49.820 ;
        RECT 123.945 49.310 126.265 52.720 ;
        RECT 126.895 52.210 127.395 52.380 ;
        RECT 120.345 48.590 126.265 49.310 ;
        RECT 113.955 45.740 120.095 46.230 ;
        RECT 120.315 47.980 124.225 48.200 ;
        RECT 109.065 45.310 112.975 45.580 ;
        RECT 120.315 45.580 122.035 47.980 ;
        RECT 122.665 47.470 123.165 47.640 ;
        RECT 122.435 46.260 122.605 47.300 ;
        RECT 123.225 46.260 123.395 47.300 ;
        RECT 122.665 45.920 123.165 46.090 ;
        RECT 123.795 45.580 124.225 47.980 ;
        RECT 125.205 46.230 126.265 48.590 ;
        RECT 126.665 46.955 126.835 51.995 ;
        RECT 127.455 46.955 127.625 51.995 ;
        RECT 126.895 46.570 127.395 46.740 ;
        RECT 128.025 46.230 128.195 52.720 ;
        RECT 128.825 52.210 129.325 52.380 ;
        RECT 128.595 46.955 128.765 51.995 ;
        RECT 129.385 46.955 129.555 51.995 ;
        RECT 128.825 46.570 129.325 46.740 ;
        RECT 129.955 46.230 131.345 52.720 ;
        RECT 125.205 45.740 131.345 46.230 ;
        RECT 120.315 45.310 124.225 45.580 ;
        RECT 25.695 39.770 29.605 40.040 ;
        RECT 18.575 39.120 24.715 39.610 ;
        RECT 18.575 32.630 19.965 39.120 ;
        RECT 20.595 38.610 21.095 38.780 ;
        RECT 20.365 33.355 20.535 38.395 ;
        RECT 21.155 33.355 21.325 38.395 ;
        RECT 20.595 32.970 21.095 33.140 ;
        RECT 21.725 32.630 21.895 39.120 ;
        RECT 22.525 38.610 23.025 38.780 ;
        RECT 22.295 33.355 22.465 38.395 ;
        RECT 23.085 33.355 23.255 38.395 ;
        RECT 23.655 36.760 24.715 39.120 ;
        RECT 25.695 37.370 26.125 39.770 ;
        RECT 26.755 39.260 27.255 39.430 ;
        RECT 26.525 38.050 26.695 39.090 ;
        RECT 27.315 38.050 27.485 39.090 ;
        RECT 26.755 37.710 27.255 37.880 ;
        RECT 27.885 37.370 29.605 39.770 ;
        RECT 36.975 39.770 40.885 40.040 ;
        RECT 25.695 37.150 29.605 37.370 ;
        RECT 29.855 39.120 35.995 39.610 ;
        RECT 23.655 36.040 29.575 36.760 ;
        RECT 22.525 32.970 23.025 33.140 ;
        RECT 23.655 32.630 25.975 36.040 ;
        RECT 26.605 35.530 27.105 35.700 ;
        RECT 26.375 33.275 26.545 35.315 ;
        RECT 27.165 33.275 27.335 35.315 ;
        RECT 26.605 32.890 27.105 33.060 ;
        RECT 18.575 32.550 25.975 32.630 ;
        RECT 27.735 32.550 29.575 36.040 ;
        RECT 18.575 30.480 29.575 32.550 ;
        RECT 18.575 19.340 19.215 30.480 ;
        RECT 19.615 20.070 19.785 30.110 ;
        RECT 20.905 20.070 21.075 30.110 ;
        RECT 19.845 19.685 20.845 19.855 ;
        RECT 21.475 19.340 21.645 30.480 ;
        RECT 22.045 20.070 22.215 30.110 ;
        RECT 27.335 20.070 27.505 30.110 ;
        RECT 22.275 19.685 27.275 19.855 ;
        RECT 27.905 19.340 29.575 30.480 ;
        RECT 18.575 18.470 29.575 19.340 ;
        RECT 29.855 32.630 31.245 39.120 ;
        RECT 31.875 38.610 32.375 38.780 ;
        RECT 31.645 33.355 31.815 38.395 ;
        RECT 32.435 33.355 32.605 38.395 ;
        RECT 31.875 32.970 32.375 33.140 ;
        RECT 33.005 32.630 33.175 39.120 ;
        RECT 33.805 38.610 34.305 38.780 ;
        RECT 33.575 33.355 33.745 38.395 ;
        RECT 34.365 33.355 34.535 38.395 ;
        RECT 34.935 36.760 35.995 39.120 ;
        RECT 36.975 37.370 37.405 39.770 ;
        RECT 38.035 39.260 38.535 39.430 ;
        RECT 37.805 38.050 37.975 39.090 ;
        RECT 38.595 38.050 38.765 39.090 ;
        RECT 38.035 37.710 38.535 37.880 ;
        RECT 39.165 37.370 40.885 39.770 ;
        RECT 48.265 39.750 52.175 40.020 ;
        RECT 36.975 37.150 40.885 37.370 ;
        RECT 41.145 39.100 47.285 39.590 ;
        RECT 34.935 36.040 40.855 36.760 ;
        RECT 33.805 32.970 34.305 33.140 ;
        RECT 34.935 32.630 37.255 36.040 ;
        RECT 37.885 35.530 38.385 35.700 ;
        RECT 37.655 33.275 37.825 35.315 ;
        RECT 38.445 33.275 38.615 35.315 ;
        RECT 37.885 32.890 38.385 33.060 ;
        RECT 29.855 32.550 37.255 32.630 ;
        RECT 39.015 32.550 40.855 36.040 ;
        RECT 29.855 30.480 40.855 32.550 ;
        RECT 29.855 19.340 30.495 30.480 ;
        RECT 30.895 20.070 31.065 30.110 ;
        RECT 32.185 20.070 32.355 30.110 ;
        RECT 31.125 19.685 32.125 19.855 ;
        RECT 32.755 19.340 32.925 30.480 ;
        RECT 33.325 20.070 33.495 30.110 ;
        RECT 38.615 20.070 38.785 30.110 ;
        RECT 33.555 19.685 38.555 19.855 ;
        RECT 39.185 19.340 40.855 30.480 ;
        RECT 29.855 18.470 40.855 19.340 ;
        RECT 41.145 32.610 42.535 39.100 ;
        RECT 43.165 38.590 43.665 38.760 ;
        RECT 42.935 33.335 43.105 38.375 ;
        RECT 43.725 33.335 43.895 38.375 ;
        RECT 43.165 32.950 43.665 33.120 ;
        RECT 44.295 32.610 44.465 39.100 ;
        RECT 45.095 38.590 45.595 38.760 ;
        RECT 44.865 33.335 45.035 38.375 ;
        RECT 45.655 33.335 45.825 38.375 ;
        RECT 46.225 36.740 47.285 39.100 ;
        RECT 48.265 37.350 48.695 39.750 ;
        RECT 49.325 39.240 49.825 39.410 ;
        RECT 49.095 38.030 49.265 39.070 ;
        RECT 49.885 38.030 50.055 39.070 ;
        RECT 49.325 37.690 49.825 37.860 ;
        RECT 50.455 37.350 52.175 39.750 ;
        RECT 59.485 39.750 63.395 40.020 ;
        RECT 48.265 37.130 52.175 37.350 ;
        RECT 52.365 39.100 58.505 39.590 ;
        RECT 46.225 36.020 52.145 36.740 ;
        RECT 45.095 32.950 45.595 33.120 ;
        RECT 46.225 32.610 48.545 36.020 ;
        RECT 49.175 35.510 49.675 35.680 ;
        RECT 48.945 33.255 49.115 35.295 ;
        RECT 49.735 33.255 49.905 35.295 ;
        RECT 49.175 32.870 49.675 33.040 ;
        RECT 41.145 32.530 48.545 32.610 ;
        RECT 50.305 32.530 52.145 36.020 ;
        RECT 41.145 30.460 52.145 32.530 ;
        RECT 41.145 19.320 41.785 30.460 ;
        RECT 42.185 20.050 42.355 30.090 ;
        RECT 43.475 20.050 43.645 30.090 ;
        RECT 42.415 19.665 43.415 19.835 ;
        RECT 44.045 19.320 44.215 30.460 ;
        RECT 44.615 20.050 44.785 30.090 ;
        RECT 49.905 20.050 50.075 30.090 ;
        RECT 44.845 19.665 49.845 19.835 ;
        RECT 50.475 19.320 52.145 30.460 ;
        RECT 41.145 18.450 52.145 19.320 ;
        RECT 52.365 32.610 53.755 39.100 ;
        RECT 54.385 38.590 54.885 38.760 ;
        RECT 54.155 33.335 54.325 38.375 ;
        RECT 54.945 33.335 55.115 38.375 ;
        RECT 54.385 32.950 54.885 33.120 ;
        RECT 55.515 32.610 55.685 39.100 ;
        RECT 56.315 38.590 56.815 38.760 ;
        RECT 56.085 33.335 56.255 38.375 ;
        RECT 56.875 33.335 57.045 38.375 ;
        RECT 57.445 36.740 58.505 39.100 ;
        RECT 59.485 37.350 59.915 39.750 ;
        RECT 60.545 39.240 61.045 39.410 ;
        RECT 60.315 38.030 60.485 39.070 ;
        RECT 61.105 38.030 61.275 39.070 ;
        RECT 60.545 37.690 61.045 37.860 ;
        RECT 61.675 37.350 63.395 39.750 ;
        RECT 70.685 39.750 74.595 40.020 ;
        RECT 59.485 37.130 63.395 37.350 ;
        RECT 63.565 39.100 69.705 39.590 ;
        RECT 57.445 36.020 63.365 36.740 ;
        RECT 56.315 32.950 56.815 33.120 ;
        RECT 57.445 32.610 59.765 36.020 ;
        RECT 60.395 35.510 60.895 35.680 ;
        RECT 60.165 33.255 60.335 35.295 ;
        RECT 60.955 33.255 61.125 35.295 ;
        RECT 60.395 32.870 60.895 33.040 ;
        RECT 52.365 32.530 59.765 32.610 ;
        RECT 61.525 32.530 63.365 36.020 ;
        RECT 52.365 30.460 63.365 32.530 ;
        RECT 52.365 19.320 53.005 30.460 ;
        RECT 53.405 20.050 53.575 30.090 ;
        RECT 54.695 20.050 54.865 30.090 ;
        RECT 53.635 19.665 54.635 19.835 ;
        RECT 55.265 19.320 55.435 30.460 ;
        RECT 55.835 20.050 56.005 30.090 ;
        RECT 61.125 20.050 61.295 30.090 ;
        RECT 56.065 19.665 61.065 19.835 ;
        RECT 61.695 19.320 63.365 30.460 ;
        RECT 52.365 18.450 63.365 19.320 ;
        RECT 63.565 32.610 64.955 39.100 ;
        RECT 65.585 38.590 66.085 38.760 ;
        RECT 65.355 33.335 65.525 38.375 ;
        RECT 66.145 33.335 66.315 38.375 ;
        RECT 65.585 32.950 66.085 33.120 ;
        RECT 66.715 32.610 66.885 39.100 ;
        RECT 67.515 38.590 68.015 38.760 ;
        RECT 67.285 33.335 67.455 38.375 ;
        RECT 68.075 33.335 68.245 38.375 ;
        RECT 68.645 36.740 69.705 39.100 ;
        RECT 70.685 37.350 71.115 39.750 ;
        RECT 71.745 39.240 72.245 39.410 ;
        RECT 71.515 38.030 71.685 39.070 ;
        RECT 72.305 38.030 72.475 39.070 ;
        RECT 71.745 37.690 72.245 37.860 ;
        RECT 72.875 37.350 74.595 39.750 ;
        RECT 81.975 39.740 85.885 40.010 ;
        RECT 70.685 37.130 74.595 37.350 ;
        RECT 74.855 39.090 80.995 39.580 ;
        RECT 68.645 36.020 74.565 36.740 ;
        RECT 67.515 32.950 68.015 33.120 ;
        RECT 68.645 32.610 70.965 36.020 ;
        RECT 71.595 35.510 72.095 35.680 ;
        RECT 71.365 33.255 71.535 35.295 ;
        RECT 72.155 33.255 72.325 35.295 ;
        RECT 71.595 32.870 72.095 33.040 ;
        RECT 63.565 32.530 70.965 32.610 ;
        RECT 72.725 32.530 74.565 36.020 ;
        RECT 63.565 30.460 74.565 32.530 ;
        RECT 63.565 19.320 64.205 30.460 ;
        RECT 64.605 20.050 64.775 30.090 ;
        RECT 65.895 20.050 66.065 30.090 ;
        RECT 64.835 19.665 65.835 19.835 ;
        RECT 66.465 19.320 66.635 30.460 ;
        RECT 67.035 20.050 67.205 30.090 ;
        RECT 72.325 20.050 72.495 30.090 ;
        RECT 67.265 19.665 72.265 19.835 ;
        RECT 72.895 19.320 74.565 30.460 ;
        RECT 63.565 18.450 74.565 19.320 ;
        RECT 74.855 32.600 76.245 39.090 ;
        RECT 76.875 38.580 77.375 38.750 ;
        RECT 76.645 33.325 76.815 38.365 ;
        RECT 77.435 33.325 77.605 38.365 ;
        RECT 76.875 32.940 77.375 33.110 ;
        RECT 78.005 32.600 78.175 39.090 ;
        RECT 78.805 38.580 79.305 38.750 ;
        RECT 78.575 33.325 78.745 38.365 ;
        RECT 79.365 33.325 79.535 38.365 ;
        RECT 79.935 36.730 80.995 39.090 ;
        RECT 81.975 37.340 82.405 39.740 ;
        RECT 83.035 39.230 83.535 39.400 ;
        RECT 82.805 38.020 82.975 39.060 ;
        RECT 83.595 38.020 83.765 39.060 ;
        RECT 83.035 37.680 83.535 37.850 ;
        RECT 84.165 37.340 85.885 39.740 ;
        RECT 93.215 39.760 97.125 40.030 ;
        RECT 81.975 37.120 85.885 37.340 ;
        RECT 86.095 39.110 92.235 39.600 ;
        RECT 79.935 36.010 85.855 36.730 ;
        RECT 78.805 32.940 79.305 33.110 ;
        RECT 79.935 32.600 82.255 36.010 ;
        RECT 82.885 35.500 83.385 35.670 ;
        RECT 82.655 33.245 82.825 35.285 ;
        RECT 83.445 33.245 83.615 35.285 ;
        RECT 82.885 32.860 83.385 33.030 ;
        RECT 74.855 32.520 82.255 32.600 ;
        RECT 84.015 32.520 85.855 36.010 ;
        RECT 74.855 30.450 85.855 32.520 ;
        RECT 74.855 19.310 75.495 30.450 ;
        RECT 75.895 20.040 76.065 30.080 ;
        RECT 77.185 20.040 77.355 30.080 ;
        RECT 76.125 19.655 77.125 19.825 ;
        RECT 77.755 19.310 77.925 30.450 ;
        RECT 78.325 20.040 78.495 30.080 ;
        RECT 83.615 20.040 83.785 30.080 ;
        RECT 78.555 19.655 83.555 19.825 ;
        RECT 84.185 19.310 85.855 30.450 ;
        RECT 74.855 18.440 85.855 19.310 ;
        RECT 86.095 32.620 87.485 39.110 ;
        RECT 88.115 38.600 88.615 38.770 ;
        RECT 87.885 33.345 88.055 38.385 ;
        RECT 88.675 33.345 88.845 38.385 ;
        RECT 88.115 32.960 88.615 33.130 ;
        RECT 89.245 32.620 89.415 39.110 ;
        RECT 90.045 38.600 90.545 38.770 ;
        RECT 89.815 33.345 89.985 38.385 ;
        RECT 90.605 33.345 90.775 38.385 ;
        RECT 91.175 36.750 92.235 39.110 ;
        RECT 93.215 37.360 93.645 39.760 ;
        RECT 94.275 39.250 94.775 39.420 ;
        RECT 94.045 38.040 94.215 39.080 ;
        RECT 94.835 38.040 95.005 39.080 ;
        RECT 94.275 37.700 94.775 37.870 ;
        RECT 95.405 37.360 97.125 39.760 ;
        RECT 104.425 39.780 108.335 40.050 ;
        RECT 93.215 37.140 97.125 37.360 ;
        RECT 97.305 39.130 103.445 39.620 ;
        RECT 91.175 36.030 97.095 36.750 ;
        RECT 90.045 32.960 90.545 33.130 ;
        RECT 91.175 32.620 93.495 36.030 ;
        RECT 94.125 35.520 94.625 35.690 ;
        RECT 93.895 33.265 94.065 35.305 ;
        RECT 94.685 33.265 94.855 35.305 ;
        RECT 94.125 32.880 94.625 33.050 ;
        RECT 86.095 32.540 93.495 32.620 ;
        RECT 95.255 32.540 97.095 36.030 ;
        RECT 86.095 30.470 97.095 32.540 ;
        RECT 86.095 19.330 86.735 30.470 ;
        RECT 87.135 20.060 87.305 30.100 ;
        RECT 88.425 20.060 88.595 30.100 ;
        RECT 87.365 19.675 88.365 19.845 ;
        RECT 88.995 19.330 89.165 30.470 ;
        RECT 89.565 20.060 89.735 30.100 ;
        RECT 94.855 20.060 95.025 30.100 ;
        RECT 89.795 19.675 94.795 19.845 ;
        RECT 95.425 19.330 97.095 30.470 ;
        RECT 86.095 18.460 97.095 19.330 ;
        RECT 97.305 32.640 98.695 39.130 ;
        RECT 99.325 38.620 99.825 38.790 ;
        RECT 99.095 33.365 99.265 38.405 ;
        RECT 99.885 33.365 100.055 38.405 ;
        RECT 99.325 32.980 99.825 33.150 ;
        RECT 100.455 32.640 100.625 39.130 ;
        RECT 101.255 38.620 101.755 38.790 ;
        RECT 101.025 33.365 101.195 38.405 ;
        RECT 101.815 33.365 101.985 38.405 ;
        RECT 102.385 36.770 103.445 39.130 ;
        RECT 104.425 37.380 104.855 39.780 ;
        RECT 105.485 39.270 105.985 39.440 ;
        RECT 105.255 38.060 105.425 39.100 ;
        RECT 106.045 38.060 106.215 39.100 ;
        RECT 105.485 37.720 105.985 37.890 ;
        RECT 106.615 37.380 108.335 39.780 ;
        RECT 115.625 39.820 119.535 40.090 ;
        RECT 104.425 37.160 108.335 37.380 ;
        RECT 108.505 39.170 114.645 39.660 ;
        RECT 102.385 36.050 108.305 36.770 ;
        RECT 101.255 32.980 101.755 33.150 ;
        RECT 102.385 32.640 104.705 36.050 ;
        RECT 105.335 35.540 105.835 35.710 ;
        RECT 105.105 33.285 105.275 35.325 ;
        RECT 105.895 33.285 106.065 35.325 ;
        RECT 105.335 32.900 105.835 33.070 ;
        RECT 97.305 32.560 104.705 32.640 ;
        RECT 106.465 32.560 108.305 36.050 ;
        RECT 97.305 30.490 108.305 32.560 ;
        RECT 97.305 19.350 97.945 30.490 ;
        RECT 98.345 20.080 98.515 30.120 ;
        RECT 99.635 20.080 99.805 30.120 ;
        RECT 98.575 19.695 99.575 19.865 ;
        RECT 100.205 19.350 100.375 30.490 ;
        RECT 100.775 20.080 100.945 30.120 ;
        RECT 106.065 20.080 106.235 30.120 ;
        RECT 101.005 19.695 106.005 19.865 ;
        RECT 106.635 19.350 108.305 30.490 ;
        RECT 97.305 18.480 108.305 19.350 ;
        RECT 108.505 32.680 109.895 39.170 ;
        RECT 110.525 38.660 111.025 38.830 ;
        RECT 110.295 33.405 110.465 38.445 ;
        RECT 111.085 33.405 111.255 38.445 ;
        RECT 110.525 33.020 111.025 33.190 ;
        RECT 111.655 32.680 111.825 39.170 ;
        RECT 112.455 38.660 112.955 38.830 ;
        RECT 112.225 33.405 112.395 38.445 ;
        RECT 113.015 33.405 113.185 38.445 ;
        RECT 113.585 36.810 114.645 39.170 ;
        RECT 115.625 37.420 116.055 39.820 ;
        RECT 116.685 39.310 117.185 39.480 ;
        RECT 116.455 38.100 116.625 39.140 ;
        RECT 117.245 38.100 117.415 39.140 ;
        RECT 116.685 37.760 117.185 37.930 ;
        RECT 117.815 37.420 119.535 39.820 ;
        RECT 126.835 39.840 130.745 40.110 ;
        RECT 115.625 37.200 119.535 37.420 ;
        RECT 119.715 39.190 125.855 39.680 ;
        RECT 113.585 36.090 119.505 36.810 ;
        RECT 112.455 33.020 112.955 33.190 ;
        RECT 113.585 32.680 115.905 36.090 ;
        RECT 116.535 35.580 117.035 35.750 ;
        RECT 116.305 33.325 116.475 35.365 ;
        RECT 117.095 33.325 117.265 35.365 ;
        RECT 116.535 32.940 117.035 33.110 ;
        RECT 108.505 32.600 115.905 32.680 ;
        RECT 117.665 32.600 119.505 36.090 ;
        RECT 108.505 30.530 119.505 32.600 ;
        RECT 108.505 19.390 109.145 30.530 ;
        RECT 109.545 20.120 109.715 30.160 ;
        RECT 110.835 20.120 111.005 30.160 ;
        RECT 109.775 19.735 110.775 19.905 ;
        RECT 111.405 19.390 111.575 30.530 ;
        RECT 111.975 20.120 112.145 30.160 ;
        RECT 117.265 20.120 117.435 30.160 ;
        RECT 112.205 19.735 117.205 19.905 ;
        RECT 117.835 19.390 119.505 30.530 ;
        RECT 108.505 18.520 119.505 19.390 ;
        RECT 119.715 32.700 121.105 39.190 ;
        RECT 121.735 38.680 122.235 38.850 ;
        RECT 121.505 33.425 121.675 38.465 ;
        RECT 122.295 33.425 122.465 38.465 ;
        RECT 121.735 33.040 122.235 33.210 ;
        RECT 122.865 32.700 123.035 39.190 ;
        RECT 123.665 38.680 124.165 38.850 ;
        RECT 123.435 33.425 123.605 38.465 ;
        RECT 124.225 33.425 124.395 38.465 ;
        RECT 124.795 36.830 125.855 39.190 ;
        RECT 126.835 37.440 127.265 39.840 ;
        RECT 127.895 39.330 128.395 39.500 ;
        RECT 127.665 38.120 127.835 39.160 ;
        RECT 128.455 38.120 128.625 39.160 ;
        RECT 127.895 37.780 128.395 37.950 ;
        RECT 129.025 37.440 130.745 39.840 ;
        RECT 126.835 37.220 130.745 37.440 ;
        RECT 124.795 36.110 130.715 36.830 ;
        RECT 123.665 33.040 124.165 33.210 ;
        RECT 124.795 32.700 127.115 36.110 ;
        RECT 127.745 35.600 128.245 35.770 ;
        RECT 127.515 33.345 127.685 35.385 ;
        RECT 128.305 33.345 128.475 35.385 ;
        RECT 127.745 32.960 128.245 33.130 ;
        RECT 119.715 32.620 127.115 32.700 ;
        RECT 128.875 32.620 130.715 36.110 ;
        RECT 119.715 31.140 130.715 32.620 ;
        RECT 119.715 30.550 139.465 31.140 ;
        RECT 119.715 19.410 120.355 30.550 ;
        RECT 120.755 20.140 120.925 30.180 ;
        RECT 122.045 20.140 122.215 30.180 ;
        RECT 120.985 19.755 121.985 19.925 ;
        RECT 122.615 19.410 122.785 30.550 ;
        RECT 129.045 30.520 139.465 30.550 ;
        RECT 123.185 20.140 123.355 30.180 ;
        RECT 128.475 20.140 128.645 30.180 ;
        RECT 123.415 19.755 128.415 19.925 ;
        RECT 129.045 19.410 132.075 30.520 ;
        RECT 132.475 20.110 132.645 30.150 ;
        RECT 137.765 20.110 137.935 30.150 ;
        RECT 132.705 19.725 137.705 19.895 ;
        RECT 119.715 19.380 132.075 19.410 ;
        RECT 138.335 19.380 139.465 30.520 ;
        RECT 119.715 18.540 139.465 19.380 ;
        RECT 131.925 18.520 139.465 18.540 ;
      LAYER met1 ;
        RECT 135.340 223.880 136.790 225.180 ;
        RECT 17.370 193.380 112.465 193.860 ;
        RECT 18.165 190.660 112.465 191.140 ;
        RECT 59.635 189.440 59.955 189.500 ;
        RECT 69.310 189.440 69.600 189.485 ;
        RECT 59.635 189.300 69.600 189.440 ;
        RECT 59.635 189.240 59.955 189.300 ;
        RECT 69.310 189.255 69.600 189.300 ;
        RECT 68.835 188.560 69.155 188.820 ;
        RECT 17.370 187.940 112.465 188.420 ;
        RECT 68.390 187.740 68.680 187.785 ;
        RECT 66.625 187.600 68.680 187.740 ;
        RECT 66.625 187.445 66.765 187.600 ;
        RECT 68.390 187.555 68.680 187.600 ;
        RECT 58.270 187.400 58.560 187.445 ;
        RECT 60.670 187.400 60.960 187.445 ;
        RECT 63.910 187.400 64.560 187.445 ;
        RECT 58.270 187.260 64.560 187.400 ;
        RECT 58.270 187.215 58.560 187.260 ;
        RECT 60.670 187.215 61.260 187.260 ;
        RECT 63.910 187.215 64.560 187.260 ;
        RECT 66.550 187.215 66.840 187.445 ;
        RECT 57.350 187.060 57.640 187.105 ;
        RECT 57.810 187.060 58.100 187.105 ;
        RECT 59.635 187.060 59.955 187.120 ;
        RECT 57.350 186.920 59.955 187.060 ;
        RECT 57.350 186.875 57.640 186.920 ;
        RECT 57.810 186.875 58.100 186.920 ;
        RECT 59.635 186.860 59.955 186.920 ;
        RECT 60.970 186.900 61.260 187.215 ;
        RECT 62.050 187.060 62.340 187.105 ;
        RECT 65.630 187.060 65.920 187.105 ;
        RECT 67.465 187.060 67.755 187.105 ;
        RECT 62.050 186.920 67.755 187.060 ;
        RECT 62.050 186.875 62.340 186.920 ;
        RECT 65.630 186.875 65.920 186.920 ;
        RECT 67.465 186.875 67.755 186.920 ;
        RECT 70.215 186.860 70.535 187.120 ;
        RECT 92.295 187.060 92.615 187.120 ;
        RECT 95.070 187.060 95.360 187.105 ;
        RECT 92.295 186.920 95.360 187.060 ;
        RECT 92.295 186.860 92.615 186.920 ;
        RECT 95.070 186.875 95.360 186.920 ;
        RECT 67.930 186.535 68.220 186.765 ;
        RECT 69.295 186.720 69.615 186.780 ;
        RECT 69.770 186.720 70.060 186.765 ;
        RECT 69.295 186.580 70.060 186.720 ;
        RECT 62.050 186.380 62.340 186.425 ;
        RECT 65.170 186.380 65.460 186.425 ;
        RECT 67.060 186.380 67.350 186.425 ;
        RECT 62.050 186.240 67.350 186.380 ;
        RECT 68.005 186.380 68.145 186.535 ;
        RECT 69.295 186.520 69.615 186.580 ;
        RECT 69.770 186.535 70.060 186.580 ;
        RECT 73.895 186.380 74.215 186.440 ;
        RECT 68.005 186.240 74.215 186.380 ;
        RECT 62.050 186.195 62.340 186.240 ;
        RECT 65.170 186.195 65.460 186.240 ;
        RECT 67.060 186.195 67.350 186.240 ;
        RECT 73.895 186.180 74.215 186.240 ;
        RECT 56.415 186.040 56.735 186.100 ;
        RECT 56.890 186.040 57.180 186.085 ;
        RECT 56.415 185.900 57.180 186.040 ;
        RECT 56.415 185.840 56.735 185.900 ;
        RECT 56.890 185.855 57.180 185.900 ;
        RECT 59.175 185.840 59.495 186.100 ;
        RECT 80.795 186.040 81.115 186.100 ;
        RECT 93.675 186.040 93.995 186.100 ;
        RECT 80.795 185.900 93.995 186.040 ;
        RECT 80.795 185.840 81.115 185.900 ;
        RECT 93.675 185.840 93.995 185.900 ;
        RECT 95.530 186.040 95.820 186.085 ;
        RECT 95.975 186.040 96.295 186.100 ;
        RECT 95.530 185.900 96.295 186.040 ;
        RECT 95.530 185.855 95.820 185.900 ;
        RECT 95.975 185.840 96.295 185.900 ;
        RECT 18.165 185.220 112.465 185.700 ;
        RECT 61.475 185.020 61.795 185.080 ;
        RECT 61.950 185.020 62.240 185.065 ;
        RECT 70.215 185.020 70.535 185.080 ;
        RECT 61.475 184.880 70.535 185.020 ;
        RECT 61.475 184.820 61.795 184.880 ;
        RECT 61.950 184.835 62.240 184.880 ;
        RECT 70.215 184.820 70.535 184.880 ;
        RECT 78.585 184.880 87.005 185.020 ;
        RECT 52.240 184.680 52.530 184.725 ;
        RECT 54.130 184.680 54.420 184.725 ;
        RECT 57.250 184.680 57.540 184.725 ;
        RECT 52.240 184.540 57.540 184.680 ;
        RECT 52.240 184.495 52.530 184.540 ;
        RECT 54.130 184.495 54.420 184.540 ;
        RECT 57.250 184.495 57.540 184.540 ;
        RECT 63.790 184.495 64.080 184.725 ;
        RECT 68.030 184.680 68.320 184.725 ;
        RECT 71.150 184.680 71.440 184.725 ;
        RECT 73.040 184.680 73.330 184.725 ;
        RECT 68.030 184.540 73.330 184.680 ;
        RECT 68.030 184.495 68.320 184.540 ;
        RECT 71.150 184.495 71.440 184.540 ;
        RECT 73.040 184.495 73.330 184.540 ;
        RECT 52.750 184.340 53.040 184.385 ;
        RECT 63.865 184.340 64.005 184.495 ;
        RECT 52.750 184.200 64.005 184.340 ;
        RECT 52.750 184.155 53.040 184.200 ;
        RECT 73.895 184.140 74.215 184.400 ;
        RECT 51.370 183.815 51.660 184.045 ;
        RECT 51.835 184.000 52.125 184.045 ;
        RECT 53.670 184.000 53.960 184.045 ;
        RECT 57.250 184.000 57.540 184.045 ;
        RECT 51.835 183.860 57.540 184.000 ;
        RECT 51.835 183.815 52.125 183.860 ;
        RECT 53.670 183.815 53.960 183.860 ;
        RECT 57.250 183.815 57.540 183.860 ;
        RECT 51.445 183.660 51.585 183.815 ;
        RECT 52.275 183.660 52.595 183.720 ;
        RECT 51.445 183.520 52.595 183.660 ;
        RECT 52.275 183.460 52.595 183.520 ;
        RECT 55.030 183.660 55.680 183.705 ;
        RECT 56.415 183.660 56.735 183.720 ;
        RECT 58.330 183.705 58.620 184.020 ;
        RECT 59.175 184.000 59.495 184.060 ;
        RECT 61.030 184.000 61.320 184.045 ;
        RECT 59.175 183.860 61.320 184.000 ;
        RECT 59.175 183.800 59.495 183.860 ;
        RECT 61.030 183.815 61.320 183.860 ;
        RECT 64.710 184.000 65.000 184.045 ;
        RECT 66.075 184.000 66.395 184.060 ;
        RECT 64.710 183.860 66.395 184.000 ;
        RECT 64.710 183.815 65.000 183.860 ;
        RECT 66.075 183.800 66.395 183.860 ;
        RECT 66.950 183.705 67.240 184.020 ;
        RECT 68.030 184.000 68.320 184.045 ;
        RECT 71.610 184.000 71.900 184.045 ;
        RECT 73.445 184.000 73.735 184.045 ;
        RECT 68.030 183.860 73.735 184.000 ;
        RECT 68.030 183.815 68.320 183.860 ;
        RECT 71.610 183.815 71.900 183.860 ;
        RECT 73.445 183.815 73.735 183.860 ;
        RECT 58.330 183.660 58.920 183.705 ;
        RECT 55.030 183.520 58.920 183.660 ;
        RECT 55.030 183.475 55.680 183.520 ;
        RECT 56.415 183.460 56.735 183.520 ;
        RECT 58.630 183.475 58.920 183.520 ;
        RECT 66.650 183.660 67.240 183.705 ;
        RECT 68.835 183.660 69.155 183.720 ;
        RECT 69.890 183.660 70.540 183.705 ;
        RECT 66.650 183.520 70.540 183.660 ;
        RECT 66.650 183.475 66.940 183.520 ;
        RECT 68.835 183.460 69.155 183.520 ;
        RECT 69.890 183.475 70.540 183.520 ;
        RECT 72.530 183.475 72.820 183.705 ;
        RECT 73.985 183.660 74.125 184.140 ;
        RECT 74.355 183.800 74.675 184.060 ;
        RECT 78.585 184.045 78.725 184.880 ;
        RECT 83.570 184.495 83.860 184.725 ;
        RECT 80.795 184.140 81.115 184.400 ;
        RECT 78.510 183.815 78.800 184.045 ;
        RECT 81.270 184.000 81.560 184.045 ;
        RECT 81.715 184.000 82.035 184.060 ;
        RECT 81.270 183.860 82.035 184.000 ;
        RECT 83.645 184.000 83.785 184.495 ;
        RECT 86.865 184.340 87.005 184.880 ;
        RECT 89.040 184.680 89.330 184.725 ;
        RECT 90.930 184.680 91.220 184.725 ;
        RECT 94.050 184.680 94.340 184.725 ;
        RECT 89.040 184.540 94.340 184.680 ;
        RECT 89.040 184.495 89.330 184.540 ;
        RECT 90.930 184.495 91.220 184.540 ;
        RECT 94.050 184.495 94.340 184.540 ;
        RECT 100.230 184.680 100.520 184.725 ;
        RECT 103.350 184.680 103.640 184.725 ;
        RECT 105.240 184.680 105.530 184.725 ;
        RECT 100.230 184.540 105.530 184.680 ;
        RECT 100.230 184.495 100.520 184.540 ;
        RECT 103.350 184.495 103.640 184.540 ;
        RECT 105.240 184.495 105.530 184.540 ;
        RECT 92.295 184.340 92.615 184.400 ;
        RECT 86.865 184.200 92.615 184.340 ;
        RECT 86.865 184.045 87.005 184.200 ;
        RECT 92.295 184.140 92.615 184.200 ;
        RECT 84.030 184.000 84.320 184.045 ;
        RECT 83.645 183.860 84.320 184.000 ;
        RECT 81.270 183.815 81.560 183.860 ;
        RECT 81.715 183.800 82.035 183.860 ;
        RECT 84.030 183.815 84.320 183.860 ;
        RECT 86.790 183.815 87.080 184.045 ;
        RECT 88.170 183.815 88.460 184.045 ;
        RECT 88.635 184.000 88.925 184.045 ;
        RECT 90.470 184.000 90.760 184.045 ;
        RECT 94.050 184.000 94.340 184.045 ;
        RECT 88.635 183.860 94.340 184.000 ;
        RECT 88.635 183.815 88.925 183.860 ;
        RECT 90.470 183.815 90.760 183.860 ;
        RECT 94.050 183.815 94.340 183.860 ;
        RECT 83.095 183.660 83.415 183.720 ;
        RECT 88.245 183.660 88.385 183.815 ;
        RECT 73.985 183.520 88.385 183.660 ;
        RECT 89.550 183.660 89.840 183.705 ;
        RECT 89.995 183.660 90.315 183.720 ;
        RECT 95.130 183.705 95.420 184.020 ;
        RECT 91.830 183.660 92.480 183.705 ;
        RECT 95.130 183.660 95.720 183.705 ;
        RECT 89.550 183.520 90.315 183.660 ;
        RECT 60.095 183.120 60.415 183.380 ;
        RECT 63.775 183.320 64.095 183.380 ;
        RECT 65.170 183.320 65.460 183.365 ;
        RECT 63.775 183.180 65.460 183.320 ;
        RECT 72.605 183.320 72.745 183.475 ;
        RECT 83.095 183.460 83.415 183.520 ;
        RECT 89.550 183.475 89.840 183.520 ;
        RECT 89.995 183.460 90.315 183.520 ;
        RECT 91.005 183.520 95.720 183.660 ;
        RECT 74.830 183.320 75.120 183.365 ;
        RECT 72.605 183.180 75.120 183.320 ;
        RECT 63.775 183.120 64.095 183.180 ;
        RECT 65.170 183.135 65.460 183.180 ;
        RECT 74.830 183.135 75.120 183.180 ;
        RECT 78.955 183.120 79.275 183.380 ;
        RECT 79.415 183.320 79.735 183.380 ;
        RECT 81.730 183.320 82.020 183.365 ;
        RECT 79.415 183.180 82.020 183.320 ;
        RECT 79.415 183.120 79.735 183.180 ;
        RECT 81.730 183.135 82.020 183.180 ;
        RECT 84.950 183.320 85.240 183.365 ;
        RECT 85.395 183.320 85.715 183.380 ;
        RECT 84.950 183.180 85.715 183.320 ;
        RECT 84.950 183.135 85.240 183.180 ;
        RECT 85.395 183.120 85.715 183.180 ;
        RECT 87.250 183.320 87.540 183.365 ;
        RECT 91.005 183.320 91.145 183.520 ;
        RECT 91.830 183.475 92.480 183.520 ;
        RECT 95.430 183.475 95.720 183.520 ;
        RECT 95.975 183.660 96.295 183.720 ;
        RECT 99.150 183.705 99.440 184.020 ;
        RECT 100.230 184.000 100.520 184.045 ;
        RECT 103.810 184.000 104.100 184.045 ;
        RECT 105.645 184.000 105.935 184.045 ;
        RECT 100.230 183.860 105.935 184.000 ;
        RECT 100.230 183.815 100.520 183.860 ;
        RECT 103.810 183.815 104.100 183.860 ;
        RECT 105.645 183.815 105.935 183.860 ;
        RECT 106.095 183.800 106.415 184.060 ;
        RECT 98.850 183.660 99.440 183.705 ;
        RECT 102.090 183.660 102.740 183.705 ;
        RECT 95.975 183.520 102.740 183.660 ;
        RECT 95.975 183.460 96.295 183.520 ;
        RECT 98.850 183.475 99.140 183.520 ;
        RECT 102.090 183.475 102.740 183.520 ;
        RECT 104.730 183.475 105.020 183.705 ;
        RECT 87.250 183.180 91.145 183.320 ;
        RECT 87.250 183.135 87.540 183.180 ;
        RECT 96.895 183.120 97.215 183.380 ;
        RECT 97.370 183.320 97.660 183.365 ;
        RECT 97.815 183.320 98.135 183.380 ;
        RECT 97.370 183.180 98.135 183.320 ;
        RECT 97.370 183.135 97.660 183.180 ;
        RECT 97.815 183.120 98.135 183.180 ;
        RECT 100.575 183.320 100.895 183.380 ;
        RECT 104.805 183.320 104.945 183.475 ;
        RECT 100.575 183.180 104.945 183.320 ;
        RECT 100.575 183.120 100.895 183.180 ;
        RECT 17.370 182.500 112.465 182.980 ;
        RECT 59.190 182.300 59.480 182.345 ;
        RECT 63.775 182.300 64.095 182.360 ;
        RECT 64.250 182.300 64.540 182.345 ;
        RECT 59.190 182.160 64.540 182.300 ;
        RECT 59.190 182.115 59.480 182.160 ;
        RECT 63.775 182.100 64.095 182.160 ;
        RECT 64.250 182.115 64.540 182.160 ;
        RECT 68.375 182.300 68.695 182.360 ;
        RECT 70.560 182.300 70.850 182.345 ;
        RECT 68.375 182.160 70.850 182.300 ;
        RECT 61.490 181.960 61.780 182.005 ;
        RECT 57.425 181.820 61.780 181.960 ;
        RECT 55.035 181.620 55.355 181.680 ;
        RECT 57.425 181.665 57.565 181.820 ;
        RECT 61.490 181.775 61.780 181.820 ;
        RECT 57.350 181.620 57.640 181.665 ;
        RECT 55.035 181.480 57.640 181.620 ;
        RECT 55.035 181.420 55.355 181.480 ;
        RECT 57.350 181.435 57.640 181.480 ;
        RECT 58.730 181.620 59.020 181.665 ;
        RECT 59.175 181.620 59.495 181.680 ;
        RECT 58.730 181.480 59.495 181.620 ;
        RECT 58.730 181.435 59.020 181.480 ;
        RECT 59.175 181.420 59.495 181.480 ;
        RECT 59.775 181.620 60.065 181.665 ;
        RECT 64.325 181.620 64.465 182.115 ;
        RECT 68.375 182.100 68.695 182.160 ;
        RECT 70.560 182.115 70.850 182.160 ;
        RECT 89.550 182.300 89.840 182.345 ;
        RECT 89.995 182.300 90.315 182.360 ;
        RECT 89.550 182.160 90.315 182.300 ;
        RECT 89.550 182.115 89.840 182.160 ;
        RECT 89.995 182.100 90.315 182.160 ;
        RECT 100.575 182.100 100.895 182.360 ;
        RECT 65.615 181.960 65.935 182.020 ;
        RECT 67.470 181.960 67.760 182.005 ;
        RECT 69.295 181.960 69.615 182.020 ;
        RECT 71.610 181.960 71.900 182.005 ;
        RECT 65.615 181.820 69.065 181.960 ;
        RECT 65.615 181.760 65.935 181.820 ;
        RECT 67.085 181.665 67.225 181.820 ;
        RECT 67.470 181.775 67.760 181.820 ;
        RECT 66.090 181.620 66.380 181.665 ;
        RECT 59.775 181.480 60.785 181.620 ;
        RECT 64.325 181.480 66.380 181.620 ;
        RECT 59.775 181.435 60.065 181.480 ;
        RECT 60.645 181.340 60.785 181.480 ;
        RECT 66.090 181.435 66.380 181.480 ;
        RECT 67.010 181.435 67.300 181.665 ;
        RECT 68.390 181.435 68.680 181.665 ;
        RECT 68.925 181.620 69.065 181.820 ;
        RECT 69.295 181.820 71.900 181.960 ;
        RECT 69.295 181.760 69.615 181.820 ;
        RECT 71.610 181.775 71.900 181.820 ;
        RECT 78.955 181.960 79.275 182.020 ;
        RECT 79.530 181.960 79.820 182.005 ;
        RECT 82.770 181.960 83.420 182.005 ;
        RECT 78.955 181.820 83.420 181.960 ;
        RECT 78.955 181.760 79.275 181.820 ;
        RECT 79.530 181.775 80.120 181.820 ;
        RECT 82.770 181.775 83.420 181.820 ;
        RECT 72.055 181.620 72.375 181.680 ;
        RECT 73.895 181.620 74.215 181.680 ;
        RECT 68.925 181.480 74.215 181.620 ;
        RECT 60.555 181.280 60.875 181.340 ;
        RECT 63.790 181.280 64.080 181.325 ;
        RECT 60.555 181.140 64.080 181.280 ;
        RECT 60.555 181.080 60.875 181.140 ;
        RECT 63.790 181.095 64.080 181.140 ;
        RECT 67.915 181.280 68.235 181.340 ;
        RECT 68.465 181.280 68.605 181.435 ;
        RECT 72.055 181.420 72.375 181.480 ;
        RECT 73.895 181.420 74.215 181.480 ;
        RECT 74.355 181.620 74.675 181.680 ;
        RECT 76.670 181.620 76.960 181.665 ;
        RECT 74.355 181.480 76.960 181.620 ;
        RECT 74.355 181.420 74.675 181.480 ;
        RECT 76.670 181.435 76.960 181.480 ;
        RECT 79.830 181.460 80.120 181.775 ;
        RECT 85.395 181.760 85.715 182.020 ;
        RECT 90.915 181.960 91.235 182.020 ;
        RECT 93.230 181.960 93.520 182.005 ;
        RECT 96.895 181.960 97.215 182.020 ;
        RECT 90.915 181.820 97.215 181.960 ;
        RECT 90.915 181.760 91.235 181.820 ;
        RECT 93.230 181.775 93.520 181.820 ;
        RECT 96.895 181.760 97.215 181.820 ;
        RECT 80.910 181.620 81.200 181.665 ;
        RECT 84.490 181.620 84.780 181.665 ;
        RECT 86.325 181.620 86.615 181.665 ;
        RECT 80.910 181.480 86.615 181.620 ;
        RECT 80.910 181.435 81.200 181.480 ;
        RECT 84.490 181.435 84.780 181.480 ;
        RECT 86.325 181.435 86.615 181.480 ;
        RECT 90.470 181.620 90.760 181.665 ;
        RECT 92.770 181.620 93.060 181.665 ;
        RECT 95.055 181.620 95.375 181.680 ;
        RECT 99.670 181.620 99.960 181.665 ;
        RECT 90.470 181.480 91.145 181.620 ;
        RECT 90.470 181.435 90.760 181.480 ;
        RECT 70.215 181.280 70.535 181.340 ;
        RECT 67.915 181.140 70.535 181.280 ;
        RECT 67.915 181.080 68.235 181.140 ;
        RECT 70.215 181.080 70.535 181.140 ;
        RECT 78.050 181.280 78.340 181.325 ;
        RECT 81.715 181.280 82.035 181.340 ;
        RECT 78.050 181.140 82.035 181.280 ;
        RECT 78.050 181.095 78.340 181.140 ;
        RECT 81.715 181.080 82.035 181.140 ;
        RECT 83.555 181.280 83.875 181.340 ;
        RECT 86.790 181.280 87.080 181.325 ;
        RECT 83.555 181.140 87.080 181.280 ;
        RECT 83.555 181.080 83.875 181.140 ;
        RECT 86.790 181.095 87.080 181.140 ;
        RECT 61.475 180.740 61.795 181.000 ;
        RECT 66.535 180.940 66.855 181.000 ;
        RECT 91.005 180.985 91.145 181.480 ;
        RECT 92.770 181.480 95.375 181.620 ;
        RECT 92.770 181.435 93.060 181.480 ;
        RECT 69.770 180.940 70.060 180.985 ;
        RECT 66.535 180.800 70.060 180.940 ;
        RECT 66.535 180.740 66.855 180.800 ;
        RECT 69.770 180.755 70.060 180.800 ;
        RECT 80.910 180.940 81.200 180.985 ;
        RECT 84.030 180.940 84.320 180.985 ;
        RECT 85.920 180.940 86.210 180.985 ;
        RECT 80.910 180.800 86.210 180.940 ;
        RECT 80.910 180.755 81.200 180.800 ;
        RECT 84.030 180.755 84.320 180.800 ;
        RECT 85.920 180.755 86.210 180.800 ;
        RECT 90.930 180.755 91.220 180.985 ;
        RECT 60.555 180.400 60.875 180.660 ;
        RECT 65.155 180.400 65.475 180.660 ;
        RECT 69.310 180.600 69.600 180.645 ;
        RECT 70.690 180.600 70.980 180.645 ;
        RECT 69.310 180.460 70.980 180.600 ;
        RECT 69.310 180.415 69.600 180.460 ;
        RECT 70.690 180.415 70.980 180.460 ;
        RECT 77.130 180.600 77.420 180.645 ;
        RECT 78.035 180.600 78.355 180.660 ;
        RECT 77.130 180.460 78.355 180.600 ;
        RECT 77.130 180.415 77.420 180.460 ;
        RECT 78.035 180.400 78.355 180.460 ;
        RECT 81.715 180.600 82.035 180.660 ;
        RECT 92.845 180.600 92.985 181.435 ;
        RECT 95.055 181.420 95.375 181.480 ;
        RECT 98.825 181.480 99.960 181.620 ;
        RECT 93.675 181.280 93.995 181.340 ;
        RECT 95.530 181.280 95.820 181.325 ;
        RECT 93.675 181.140 95.820 181.280 ;
        RECT 93.675 181.080 93.995 181.140 ;
        RECT 95.530 181.095 95.820 181.140 ;
        RECT 96.435 181.280 96.755 181.340 ;
        RECT 97.815 181.280 98.135 181.340 ;
        RECT 96.435 181.140 98.135 181.280 ;
        RECT 96.435 181.080 96.755 181.140 ;
        RECT 97.815 181.080 98.135 181.140 ;
        RECT 98.825 180.985 98.965 181.480 ;
        RECT 99.670 181.435 99.960 181.480 ;
        RECT 98.750 180.755 99.040 180.985 ;
        RECT 81.715 180.460 92.985 180.600 ;
        RECT 81.715 180.400 82.035 180.460 ;
        RECT 18.165 179.780 112.465 180.260 ;
        RECT 62.855 179.380 63.175 179.640 ;
        RECT 66.075 179.580 66.395 179.640 ;
        RECT 66.995 179.580 67.315 179.640 ;
        RECT 63.405 179.440 67.315 179.580 ;
        RECT 48.105 179.240 48.395 179.285 ;
        RECT 50.885 179.240 51.175 179.285 ;
        RECT 52.745 179.240 53.035 179.285 ;
        RECT 48.105 179.100 53.035 179.240 ;
        RECT 48.105 179.055 48.395 179.100 ;
        RECT 50.885 179.055 51.175 179.100 ;
        RECT 52.745 179.055 53.035 179.100 ;
        RECT 60.110 179.240 60.400 179.285 ;
        RECT 63.405 179.240 63.545 179.440 ;
        RECT 66.075 179.380 66.395 179.440 ;
        RECT 66.995 179.380 67.315 179.440 ;
        RECT 69.295 179.380 69.615 179.640 ;
        RECT 60.110 179.100 63.545 179.240 ;
        RECT 60.110 179.055 60.400 179.100 ;
        RECT 63.775 179.040 64.095 179.300 ;
        RECT 78.925 179.240 79.215 179.285 ;
        RECT 81.705 179.240 81.995 179.285 ;
        RECT 83.565 179.240 83.855 179.285 ;
        RECT 78.925 179.100 83.855 179.240 ;
        RECT 78.925 179.055 79.215 179.100 ;
        RECT 81.705 179.055 81.995 179.100 ;
        RECT 83.565 179.055 83.855 179.100 ;
        RECT 84.490 179.055 84.780 179.285 ;
        RECT 96.550 179.240 96.840 179.285 ;
        RECT 99.670 179.240 99.960 179.285 ;
        RECT 101.560 179.240 101.850 179.285 ;
        RECT 102.890 179.240 103.180 179.285 ;
        RECT 96.550 179.100 101.850 179.240 ;
        RECT 96.550 179.055 96.840 179.100 ;
        RECT 99.670 179.055 99.960 179.100 ;
        RECT 101.560 179.055 101.850 179.100 ;
        RECT 102.045 179.100 103.180 179.240 ;
        RECT 49.055 178.900 49.375 178.960 ;
        RECT 43.625 178.760 49.375 178.900 ;
        RECT 43.625 178.605 43.765 178.760 ;
        RECT 49.055 178.700 49.375 178.760 ;
        RECT 52.275 178.900 52.595 178.960 ;
        RECT 53.210 178.900 53.500 178.945 ;
        RECT 52.275 178.760 53.500 178.900 ;
        RECT 52.275 178.700 52.595 178.760 ;
        RECT 53.210 178.715 53.500 178.760 ;
        RECT 61.475 178.900 61.795 178.960 ;
        RECT 65.170 178.900 65.460 178.945 ;
        RECT 61.475 178.760 65.460 178.900 ;
        RECT 61.475 178.700 61.795 178.760 ;
        RECT 65.170 178.715 65.460 178.760 ;
        RECT 65.615 178.700 65.935 178.960 ;
        RECT 66.075 178.700 66.395 178.960 ;
        RECT 66.550 178.900 66.840 178.945 ;
        RECT 66.995 178.900 67.315 178.960 ;
        RECT 72.055 178.900 72.375 178.960 ;
        RECT 79.415 178.900 79.735 178.960 ;
        RECT 66.550 178.760 67.315 178.900 ;
        RECT 66.550 178.715 66.840 178.760 ;
        RECT 66.995 178.700 67.315 178.760 ;
        RECT 69.385 178.760 72.375 178.900 ;
        RECT 43.550 178.375 43.840 178.605 ;
        RECT 48.105 178.560 48.395 178.605 ;
        RECT 48.105 178.420 50.640 178.560 ;
        RECT 48.105 178.375 48.395 178.420 ;
        RECT 46.245 178.220 46.535 178.265 ;
        RECT 48.595 178.220 48.915 178.280 ;
        RECT 50.425 178.265 50.640 178.420 ;
        RECT 51.355 178.360 51.675 178.620 ;
        RECT 59.190 178.560 59.480 178.605 ;
        RECT 60.095 178.560 60.415 178.620 ;
        RECT 59.190 178.420 60.415 178.560 ;
        RECT 59.190 178.375 59.480 178.420 ;
        RECT 60.095 178.360 60.415 178.420 ;
        RECT 63.775 178.560 64.095 178.620 ;
        RECT 68.390 178.560 68.680 178.605 ;
        RECT 63.775 178.420 68.680 178.560 ;
        RECT 63.775 178.360 64.095 178.420 ;
        RECT 68.390 178.375 68.680 178.420 ;
        RECT 68.885 178.560 69.175 178.605 ;
        RECT 69.385 178.560 69.525 178.760 ;
        RECT 72.055 178.700 72.375 178.760 ;
        RECT 76.745 178.760 79.735 178.900 ;
        RECT 68.885 178.420 69.525 178.560 ;
        RECT 69.770 178.560 70.060 178.605 ;
        RECT 70.215 178.560 70.535 178.620 ;
        RECT 69.770 178.420 70.535 178.560 ;
        RECT 68.885 178.375 69.175 178.420 ;
        RECT 69.770 178.375 70.060 178.420 ;
        RECT 70.215 178.360 70.535 178.420 ;
        RECT 49.505 178.220 49.795 178.265 ;
        RECT 46.245 178.080 49.795 178.220 ;
        RECT 46.245 178.035 46.535 178.080 ;
        RECT 48.595 178.020 48.915 178.080 ;
        RECT 49.505 178.035 49.795 178.080 ;
        RECT 50.425 178.220 50.715 178.265 ;
        RECT 52.285 178.220 52.575 178.265 ;
        RECT 50.425 178.080 52.575 178.220 ;
        RECT 50.425 178.035 50.715 178.080 ;
        RECT 52.285 178.035 52.575 178.080 ;
        RECT 61.950 178.220 62.240 178.265 ;
        RECT 73.895 178.220 74.215 178.280 ;
        RECT 75.060 178.220 75.350 178.265 ;
        RECT 76.745 178.220 76.885 178.760 ;
        RECT 79.415 178.700 79.735 178.760 ;
        RECT 83.095 178.900 83.415 178.960 ;
        RECT 84.030 178.900 84.320 178.945 ;
        RECT 83.095 178.760 84.320 178.900 ;
        RECT 83.095 178.700 83.415 178.760 ;
        RECT 84.030 178.715 84.320 178.760 ;
        RECT 78.925 178.560 79.215 178.605 ;
        RECT 82.190 178.560 82.480 178.605 ;
        RECT 84.565 178.560 84.705 179.055 ;
        RECT 91.375 178.900 91.695 178.960 ;
        RECT 93.675 178.900 93.995 178.960 ;
        RECT 91.375 178.760 93.995 178.900 ;
        RECT 91.375 178.700 91.695 178.760 ;
        RECT 93.675 178.700 93.995 178.760 ;
        RECT 101.050 178.900 101.340 178.945 ;
        RECT 102.045 178.900 102.185 179.100 ;
        RECT 102.890 179.055 103.180 179.100 ;
        RECT 106.095 178.900 106.415 178.960 ;
        RECT 101.050 178.760 102.185 178.900 ;
        RECT 102.505 178.760 106.415 178.900 ;
        RECT 101.050 178.715 101.340 178.760 ;
        RECT 78.925 178.420 81.460 178.560 ;
        RECT 78.925 178.375 79.215 178.420 ;
        RECT 61.950 178.080 68.605 178.220 ;
        RECT 61.950 178.035 62.240 178.080 ;
        RECT 68.465 177.940 68.605 178.080 ;
        RECT 73.895 178.080 76.885 178.220 ;
        RECT 77.065 178.220 77.355 178.265 ;
        RECT 78.035 178.220 78.355 178.280 ;
        RECT 81.245 178.265 81.460 178.420 ;
        RECT 82.190 178.420 84.705 178.560 ;
        RECT 82.190 178.375 82.480 178.420 ;
        RECT 85.410 178.375 85.700 178.605 ;
        RECT 80.325 178.220 80.615 178.265 ;
        RECT 77.065 178.080 80.615 178.220 ;
        RECT 73.895 178.020 74.215 178.080 ;
        RECT 75.060 178.035 75.350 178.080 ;
        RECT 77.065 178.035 77.355 178.080 ;
        RECT 78.035 178.020 78.355 178.080 ;
        RECT 80.325 178.035 80.615 178.080 ;
        RECT 81.245 178.220 81.535 178.265 ;
        RECT 83.105 178.220 83.395 178.265 ;
        RECT 81.245 178.080 83.395 178.220 ;
        RECT 81.245 178.035 81.535 178.080 ;
        RECT 83.105 178.035 83.395 178.080 ;
        RECT 43.090 177.880 43.380 177.925 ;
        RECT 43.535 177.880 43.855 177.940 ;
        RECT 43.090 177.740 43.855 177.880 ;
        RECT 43.090 177.695 43.380 177.740 ;
        RECT 43.535 177.680 43.855 177.740 ;
        RECT 43.995 177.925 44.315 177.940 ;
        RECT 43.995 177.695 44.530 177.925 ;
        RECT 63.000 177.880 63.290 177.925 ;
        RECT 64.250 177.880 64.540 177.925 ;
        RECT 63.000 177.740 64.540 177.880 ;
        RECT 63.000 177.695 63.290 177.740 ;
        RECT 64.250 177.695 64.540 177.740 ;
        RECT 66.535 177.880 66.855 177.940 ;
        RECT 67.470 177.880 67.760 177.925 ;
        RECT 66.535 177.740 67.760 177.880 ;
        RECT 43.995 177.680 44.315 177.695 ;
        RECT 66.535 177.680 66.855 177.740 ;
        RECT 67.470 177.695 67.760 177.740 ;
        RECT 68.375 177.680 68.695 177.940 ;
        RECT 72.975 177.880 73.295 177.940 ;
        RECT 85.485 177.880 85.625 178.375 ;
        RECT 92.295 178.360 92.615 178.620 ;
        RECT 102.505 178.605 102.645 178.760 ;
        RECT 106.095 178.700 106.415 178.760 ;
        RECT 95.470 178.265 95.760 178.580 ;
        RECT 96.550 178.560 96.840 178.605 ;
        RECT 100.130 178.560 100.420 178.605 ;
        RECT 101.965 178.560 102.255 178.605 ;
        RECT 96.550 178.420 102.255 178.560 ;
        RECT 96.550 178.375 96.840 178.420 ;
        RECT 100.130 178.375 100.420 178.420 ;
        RECT 101.965 178.375 102.255 178.420 ;
        RECT 102.430 178.375 102.720 178.605 ;
        RECT 103.810 178.375 104.100 178.605 ;
        RECT 92.770 178.220 93.060 178.265 ;
        RECT 95.170 178.220 95.760 178.265 ;
        RECT 98.410 178.220 99.060 178.265 ;
        RECT 92.770 178.080 99.060 178.220 ;
        RECT 92.770 178.035 93.060 178.080 ;
        RECT 95.170 178.035 95.460 178.080 ;
        RECT 98.410 178.035 99.060 178.080 ;
        RECT 99.655 178.220 99.975 178.280 ;
        RECT 102.505 178.220 102.645 178.375 ;
        RECT 99.655 178.080 102.645 178.220 ;
        RECT 99.655 178.020 99.975 178.080 ;
        RECT 72.975 177.740 85.625 177.880 ;
        RECT 72.975 177.680 73.295 177.740 ;
        RECT 93.675 177.680 93.995 177.940 ;
        RECT 99.195 177.880 99.515 177.940 ;
        RECT 103.885 177.880 104.025 178.375 ;
        RECT 99.195 177.740 104.025 177.880 ;
        RECT 99.195 177.680 99.515 177.740 ;
        RECT 17.370 177.060 112.465 177.540 ;
        RECT 48.595 176.660 48.915 176.920 ;
        RECT 51.355 176.660 51.675 176.920 ;
        RECT 53.210 176.675 53.500 176.905 ;
        RECT 65.615 176.860 65.935 176.920 ;
        RECT 66.995 176.860 67.315 176.920 ;
        RECT 55.125 176.720 67.315 176.860 ;
        RECT 43.535 176.565 43.855 176.580 ;
        RECT 40.265 176.520 40.555 176.565 ;
        RECT 43.525 176.520 43.855 176.565 ;
        RECT 40.265 176.380 43.855 176.520 ;
        RECT 40.265 176.335 40.555 176.380 ;
        RECT 43.525 176.335 43.855 176.380 ;
        RECT 43.535 176.320 43.855 176.335 ;
        RECT 44.445 176.520 44.735 176.565 ;
        RECT 46.305 176.520 46.595 176.565 ;
        RECT 53.285 176.520 53.425 176.675 ;
        RECT 55.125 176.580 55.265 176.720 ;
        RECT 65.615 176.660 65.935 176.720 ;
        RECT 66.995 176.660 67.315 176.720 ;
        RECT 68.375 176.660 68.695 176.920 ;
        RECT 72.975 176.660 73.295 176.920 ;
        RECT 74.355 176.860 74.675 176.920 ;
        RECT 89.995 176.860 90.315 176.920 ;
        RECT 74.355 176.720 101.725 176.860 ;
        RECT 74.355 176.660 74.675 176.720 ;
        RECT 44.445 176.380 46.595 176.520 ;
        RECT 44.445 176.335 44.735 176.380 ;
        RECT 46.305 176.335 46.595 176.380 ;
        RECT 48.685 176.380 53.425 176.520 ;
        RECT 42.125 176.180 42.415 176.225 ;
        RECT 44.445 176.180 44.660 176.335 ;
        RECT 42.125 176.040 44.660 176.180 ;
        RECT 45.390 176.180 45.680 176.225 ;
        RECT 48.685 176.180 48.825 176.380 ;
        RECT 55.035 176.320 55.355 176.580 ;
        RECT 57.910 176.520 58.200 176.565 ;
        RECT 58.715 176.520 59.035 176.580 ;
        RECT 61.150 176.520 61.800 176.565 ;
        RECT 57.910 176.380 61.800 176.520 ;
        RECT 57.910 176.335 58.500 176.380 ;
        RECT 45.390 176.040 48.825 176.180 ;
        RECT 42.125 175.995 42.415 176.040 ;
        RECT 45.390 175.995 45.680 176.040 ;
        RECT 49.055 175.980 49.375 176.240 ;
        RECT 50.435 175.980 50.755 176.240 ;
        RECT 51.355 176.180 51.675 176.240 ;
        RECT 52.750 176.180 53.040 176.225 ;
        RECT 51.355 176.040 53.040 176.180 ;
        RECT 51.355 175.980 51.675 176.040 ;
        RECT 52.750 175.995 53.040 176.040 ;
        RECT 53.195 176.180 53.515 176.240 ;
        RECT 54.130 176.180 54.420 176.225 ;
        RECT 53.195 176.040 54.420 176.180 ;
        RECT 53.195 175.980 53.515 176.040 ;
        RECT 54.130 175.995 54.420 176.040 ;
        RECT 58.210 176.020 58.500 176.335 ;
        RECT 58.715 176.320 59.035 176.380 ;
        RECT 61.150 176.335 61.800 176.380 ;
        RECT 63.790 176.520 64.080 176.565 ;
        RECT 66.535 176.520 66.855 176.580 ;
        RECT 63.790 176.380 66.855 176.520 ;
        RECT 67.085 176.520 67.225 176.660 ;
        RECT 70.215 176.520 70.535 176.580 ;
        RECT 67.085 176.380 70.535 176.520 ;
        RECT 63.790 176.335 64.080 176.380 ;
        RECT 66.535 176.320 66.855 176.380 ;
        RECT 70.215 176.320 70.535 176.380 ;
        RECT 70.690 176.520 70.980 176.565 ;
        RECT 73.895 176.520 74.215 176.580 ;
        RECT 70.690 176.380 74.215 176.520 ;
        RECT 70.690 176.335 70.980 176.380 ;
        RECT 73.895 176.320 74.215 176.380 ;
        RECT 75.275 176.520 75.595 176.580 ;
        RECT 76.145 176.520 76.435 176.565 ;
        RECT 79.405 176.520 79.695 176.565 ;
        RECT 75.275 176.380 79.695 176.520 ;
        RECT 75.275 176.320 75.595 176.380 ;
        RECT 76.145 176.335 76.435 176.380 ;
        RECT 79.405 176.335 79.695 176.380 ;
        RECT 80.325 176.520 80.615 176.565 ;
        RECT 82.185 176.520 82.475 176.565 ;
        RECT 80.325 176.380 82.475 176.520 ;
        RECT 80.325 176.335 80.615 176.380 ;
        RECT 82.185 176.335 82.475 176.380 ;
        RECT 59.290 176.180 59.580 176.225 ;
        RECT 62.870 176.180 63.160 176.225 ;
        RECT 64.705 176.180 64.995 176.225 ;
        RECT 59.290 176.040 64.995 176.180 ;
        RECT 59.290 175.995 59.580 176.040 ;
        RECT 62.870 175.995 63.160 176.040 ;
        RECT 64.705 175.995 64.995 176.040 ;
        RECT 65.615 175.980 65.935 176.240 ;
        RECT 71.150 176.180 71.440 176.225 ;
        RECT 78.005 176.180 78.295 176.225 ;
        RECT 80.325 176.180 80.540 176.335 ;
        RECT 71.150 176.040 74.355 176.180 ;
        RECT 71.150 175.995 71.440 176.040 ;
        RECT 38.260 175.840 38.550 175.885 ;
        RECT 38.935 175.840 39.255 175.900 ;
        RECT 38.260 175.700 39.255 175.840 ;
        RECT 38.260 175.655 38.550 175.700 ;
        RECT 38.935 175.640 39.255 175.700 ;
        RECT 47.230 175.840 47.520 175.885 ;
        RECT 52.275 175.840 52.595 175.900 ;
        RECT 57.335 175.840 57.655 175.900 ;
        RECT 65.170 175.840 65.460 175.885 ;
        RECT 47.230 175.700 65.460 175.840 ;
        RECT 47.230 175.655 47.520 175.700 ;
        RECT 52.275 175.640 52.595 175.700 ;
        RECT 57.335 175.640 57.655 175.700 ;
        RECT 65.170 175.655 65.460 175.700 ;
        RECT 66.995 175.640 67.315 175.900 ;
        RECT 70.230 175.655 70.520 175.885 ;
        RECT 42.125 175.500 42.415 175.545 ;
        RECT 44.905 175.500 45.195 175.545 ;
        RECT 46.765 175.500 47.055 175.545 ;
        RECT 52.735 175.500 53.055 175.560 ;
        RECT 42.125 175.360 47.055 175.500 ;
        RECT 42.125 175.315 42.415 175.360 ;
        RECT 44.905 175.315 45.195 175.360 ;
        RECT 46.765 175.315 47.055 175.360 ;
        RECT 47.305 175.360 53.055 175.500 ;
        RECT 47.305 175.220 47.445 175.360 ;
        RECT 52.735 175.300 53.055 175.360 ;
        RECT 59.290 175.500 59.580 175.545 ;
        RECT 62.410 175.500 62.700 175.545 ;
        RECT 64.300 175.500 64.590 175.545 ;
        RECT 59.290 175.360 64.590 175.500 ;
        RECT 70.305 175.500 70.445 175.655 ;
        RECT 72.975 175.500 73.295 175.560 ;
        RECT 70.305 175.360 73.295 175.500 ;
        RECT 59.290 175.315 59.580 175.360 ;
        RECT 62.410 175.315 62.700 175.360 ;
        RECT 64.300 175.315 64.590 175.360 ;
        RECT 72.975 175.300 73.295 175.360 ;
        RECT 47.215 174.960 47.535 175.220 ;
        RECT 49.055 175.160 49.375 175.220 ;
        RECT 51.355 175.160 51.675 175.220 ;
        RECT 49.055 175.020 51.675 175.160 ;
        RECT 49.055 174.960 49.375 175.020 ;
        RECT 51.355 174.960 51.675 175.020 ;
        RECT 51.815 175.160 52.135 175.220 ;
        RECT 52.290 175.160 52.580 175.205 ;
        RECT 51.815 175.020 52.580 175.160 ;
        RECT 51.815 174.960 52.135 175.020 ;
        RECT 52.290 174.975 52.580 175.020 ;
        RECT 61.475 175.160 61.795 175.220 ;
        RECT 66.090 175.160 66.380 175.205 ;
        RECT 71.135 175.160 71.455 175.220 ;
        RECT 74.215 175.205 74.355 176.040 ;
        RECT 78.005 176.040 80.540 176.180 ;
        RECT 85.025 176.180 85.165 176.720 ;
        RECT 89.995 176.660 90.315 176.720 ;
        RECT 85.395 176.520 85.715 176.580 ;
        RECT 90.570 176.520 90.860 176.565 ;
        RECT 93.810 176.520 94.460 176.565 ;
        RECT 85.395 176.380 94.460 176.520 ;
        RECT 85.395 176.320 85.715 176.380 ;
        RECT 90.570 176.335 91.160 176.380 ;
        RECT 93.810 176.335 94.460 176.380 ;
        RECT 85.870 176.180 86.160 176.225 ;
        RECT 85.025 176.040 86.160 176.180 ;
        RECT 78.005 175.995 78.295 176.040 ;
        RECT 85.870 175.995 86.160 176.040 ;
        RECT 87.695 175.980 88.015 176.240 ;
        RECT 90.870 176.020 91.160 176.335 ;
        RECT 91.950 176.180 92.240 176.225 ;
        RECT 95.530 176.180 95.820 176.225 ;
        RECT 97.365 176.180 97.655 176.225 ;
        RECT 91.950 176.040 97.655 176.180 ;
        RECT 101.585 176.180 101.725 176.720 ;
        RECT 101.970 176.180 102.260 176.225 ;
        RECT 104.255 176.180 104.575 176.240 ;
        RECT 101.585 176.040 104.575 176.180 ;
        RECT 91.950 175.995 92.240 176.040 ;
        RECT 95.530 175.995 95.820 176.040 ;
        RECT 97.365 175.995 97.655 176.040 ;
        RECT 101.970 175.995 102.260 176.040 ;
        RECT 104.255 175.980 104.575 176.040 ;
        RECT 81.270 175.840 81.560 175.885 ;
        RECT 81.715 175.840 82.035 175.900 ;
        RECT 81.270 175.700 82.035 175.840 ;
        RECT 81.270 175.655 81.560 175.700 ;
        RECT 81.715 175.640 82.035 175.700 ;
        RECT 83.095 175.640 83.415 175.900 ;
        RECT 86.330 175.840 86.620 175.885 ;
        RECT 88.615 175.840 88.935 175.900 ;
        RECT 86.330 175.700 88.935 175.840 ;
        RECT 86.330 175.655 86.620 175.700 ;
        RECT 88.615 175.640 88.935 175.700 ;
        RECT 95.975 175.840 96.295 175.900 ;
        RECT 97.830 175.840 98.120 175.885 ;
        RECT 99.655 175.840 99.975 175.900 ;
        RECT 95.975 175.700 99.975 175.840 ;
        RECT 95.975 175.640 96.295 175.700 ;
        RECT 97.830 175.655 98.120 175.700 ;
        RECT 99.655 175.640 99.975 175.700 ;
        RECT 102.430 175.840 102.720 175.885 ;
        RECT 102.875 175.840 103.195 175.900 ;
        RECT 102.430 175.700 103.195 175.840 ;
        RECT 102.430 175.655 102.720 175.700 ;
        RECT 102.875 175.640 103.195 175.700 ;
        RECT 103.810 175.840 104.100 175.885 ;
        RECT 104.715 175.840 105.035 175.900 ;
        RECT 103.810 175.700 105.035 175.840 ;
        RECT 103.810 175.655 104.100 175.700 ;
        RECT 104.715 175.640 105.035 175.700 ;
        RECT 78.005 175.500 78.295 175.545 ;
        RECT 80.785 175.500 81.075 175.545 ;
        RECT 82.645 175.500 82.935 175.545 ;
        RECT 78.005 175.360 82.935 175.500 ;
        RECT 78.005 175.315 78.295 175.360 ;
        RECT 80.785 175.315 81.075 175.360 ;
        RECT 82.645 175.315 82.935 175.360 ;
        RECT 89.090 175.500 89.380 175.545 ;
        RECT 90.455 175.500 90.775 175.560 ;
        RECT 89.090 175.360 90.775 175.500 ;
        RECT 89.090 175.315 89.380 175.360 ;
        RECT 90.455 175.300 90.775 175.360 ;
        RECT 91.950 175.500 92.240 175.545 ;
        RECT 95.070 175.500 95.360 175.545 ;
        RECT 96.960 175.500 97.250 175.545 ;
        RECT 91.950 175.360 97.250 175.500 ;
        RECT 91.950 175.315 92.240 175.360 ;
        RECT 95.070 175.315 95.360 175.360 ;
        RECT 96.960 175.315 97.250 175.360 ;
        RECT 61.475 175.020 71.455 175.160 ;
        RECT 61.475 174.960 61.795 175.020 ;
        RECT 66.090 174.975 66.380 175.020 ;
        RECT 71.135 174.960 71.455 175.020 ;
        RECT 74.140 175.160 74.430 175.205 ;
        RECT 74.815 175.160 75.135 175.220 ;
        RECT 74.140 175.020 75.135 175.160 ;
        RECT 74.140 174.975 74.430 175.020 ;
        RECT 74.815 174.960 75.135 175.020 ;
        RECT 88.630 175.160 88.920 175.205 ;
        RECT 94.135 175.160 94.455 175.220 ;
        RECT 88.630 175.020 94.455 175.160 ;
        RECT 88.630 174.975 88.920 175.020 ;
        RECT 94.135 174.960 94.455 175.020 ;
        RECT 96.545 175.160 96.835 175.205 ;
        RECT 97.355 175.160 97.675 175.220 ;
        RECT 96.545 175.020 97.675 175.160 ;
        RECT 96.545 174.975 96.835 175.020 ;
        RECT 97.355 174.960 97.675 175.020 ;
        RECT 18.165 174.340 112.465 174.820 ;
        RECT 135.635 174.550 136.775 223.880 ;
        RECT 138.130 223.810 139.580 225.110 ;
        RECT 143.180 223.840 144.630 225.140 ;
        RECT 43.550 174.140 43.840 174.185 ;
        RECT 47.215 174.140 47.535 174.200 ;
        RECT 43.550 174.000 47.535 174.140 ;
        RECT 43.550 173.955 43.840 174.000 ;
        RECT 47.215 173.940 47.535 174.000 ;
        RECT 58.715 174.140 59.035 174.200 ;
        RECT 59.650 174.140 59.940 174.185 ;
        RECT 58.715 174.000 59.940 174.140 ;
        RECT 58.715 173.940 59.035 174.000 ;
        RECT 59.650 173.955 59.940 174.000 ;
        RECT 63.775 174.140 64.095 174.200 ;
        RECT 64.710 174.140 65.000 174.185 ;
        RECT 63.775 174.000 65.000 174.140 ;
        RECT 63.775 173.940 64.095 174.000 ;
        RECT 64.710 173.955 65.000 174.000 ;
        RECT 66.995 173.940 67.315 174.200 ;
        RECT 67.915 174.140 68.235 174.200 ;
        RECT 74.370 174.140 74.660 174.185 ;
        RECT 75.275 174.140 75.595 174.200 ;
        RECT 67.915 174.000 72.745 174.140 ;
        RECT 67.915 173.940 68.235 174.000 ;
        RECT 47.690 173.800 47.980 173.845 ;
        RECT 50.435 173.800 50.755 173.860 ;
        RECT 47.690 173.660 50.755 173.800 ;
        RECT 47.690 173.615 47.980 173.660 ;
        RECT 50.435 173.600 50.755 173.660 ;
        RECT 52.245 173.800 52.535 173.845 ;
        RECT 55.025 173.800 55.315 173.845 ;
        RECT 56.885 173.800 57.175 173.845 ;
        RECT 52.245 173.660 57.175 173.800 ;
        RECT 52.245 173.615 52.535 173.660 ;
        RECT 55.025 173.615 55.315 173.660 ;
        RECT 56.885 173.615 57.175 173.660 ;
        RECT 62.855 173.800 63.175 173.860 ;
        RECT 71.150 173.800 71.440 173.845 ;
        RECT 62.855 173.660 71.440 173.800 ;
        RECT 62.855 173.600 63.175 173.660 ;
        RECT 40.790 173.460 41.080 173.505 ;
        RECT 44.930 173.460 45.220 173.505 ;
        RECT 49.515 173.460 49.835 173.520 ;
        RECT 40.790 173.320 49.835 173.460 ;
        RECT 40.790 173.275 41.080 173.320 ;
        RECT 44.930 173.275 45.220 173.320 ;
        RECT 49.515 173.260 49.835 173.320 ;
        RECT 57.335 173.260 57.655 173.520 ;
        RECT 65.630 173.460 65.920 173.505 ;
        RECT 67.915 173.460 68.235 173.520 ;
        RECT 68.925 173.505 69.065 173.660 ;
        RECT 71.150 173.615 71.440 173.660 ;
        RECT 72.605 173.505 72.745 174.000 ;
        RECT 74.370 174.000 75.595 174.140 ;
        RECT 74.370 173.955 74.660 174.000 ;
        RECT 75.275 173.940 75.595 174.000 ;
        RECT 81.715 173.940 82.035 174.200 ;
        RECT 85.395 173.940 85.715 174.200 ;
        RECT 91.375 174.140 91.695 174.200 ;
        RECT 99.195 174.140 99.515 174.200 ;
        RECT 99.670 174.140 99.960 174.185 ;
        RECT 91.375 174.000 96.665 174.140 ;
        RECT 91.375 173.940 91.695 174.000 ;
        RECT 89.650 173.800 89.940 173.845 ;
        RECT 92.770 173.800 93.060 173.845 ;
        RECT 94.660 173.800 94.950 173.845 ;
        RECT 89.650 173.660 94.950 173.800 ;
        RECT 89.650 173.615 89.940 173.660 ;
        RECT 92.770 173.615 93.060 173.660 ;
        RECT 94.660 173.615 94.950 173.660 ;
        RECT 65.630 173.320 68.235 173.460 ;
        RECT 65.630 173.275 65.920 173.320 ;
        RECT 67.915 173.260 68.235 173.320 ;
        RECT 68.850 173.275 69.140 173.505 ;
        RECT 72.530 173.275 72.820 173.505 ;
        RECT 72.975 173.460 73.295 173.520 ;
        RECT 76.210 173.460 76.500 173.505 ;
        RECT 78.495 173.460 78.815 173.520 ;
        RECT 92.295 173.460 92.615 173.520 ;
        RECT 72.975 173.320 78.815 173.460 ;
        RECT 72.975 173.260 73.295 173.320 ;
        RECT 76.210 173.275 76.500 173.320 ;
        RECT 78.495 173.260 78.815 173.320 ;
        RECT 85.025 173.320 92.615 173.460 ;
        RECT 85.025 173.180 85.165 173.320 ;
        RECT 92.295 173.260 92.615 173.320 ;
        RECT 94.135 173.260 94.455 173.520 ;
        RECT 96.525 173.505 96.665 174.000 ;
        RECT 99.195 174.000 99.960 174.140 ;
        RECT 99.195 173.940 99.515 174.000 ;
        RECT 99.670 173.955 99.960 174.000 ;
        RECT 103.910 173.800 104.200 173.845 ;
        RECT 107.030 173.800 107.320 173.845 ;
        RECT 108.920 173.800 109.210 173.845 ;
        RECT 103.910 173.660 109.210 173.800 ;
        RECT 103.910 173.615 104.200 173.660 ;
        RECT 107.030 173.615 107.320 173.660 ;
        RECT 108.920 173.615 109.210 173.660 ;
        RECT 96.450 173.275 96.740 173.505 ;
        RECT 135.580 173.430 136.830 174.550 ;
        RECT 135.635 173.420 136.775 173.430 ;
        RECT 25.135 173.120 25.455 173.180 ;
        RECT 38.490 173.120 38.780 173.165 ;
        RECT 25.135 172.980 38.780 173.120 ;
        RECT 25.135 172.920 25.455 172.980 ;
        RECT 38.490 172.935 38.780 172.980 ;
        RECT 38.935 173.120 39.255 173.180 ;
        RECT 52.245 173.120 52.535 173.165 ;
        RECT 38.935 172.980 41.465 173.120 ;
        RECT 38.935 172.920 39.255 172.980 ;
        RECT 38.935 172.240 39.255 172.500 ;
        RECT 41.325 172.485 41.465 172.980 ;
        RECT 52.245 172.980 54.780 173.120 ;
        RECT 52.245 172.935 52.535 172.980 ;
        RECT 41.710 172.780 42.000 172.825 ;
        RECT 43.535 172.780 43.855 172.840 ;
        RECT 45.390 172.780 45.680 172.825 ;
        RECT 41.710 172.640 45.680 172.780 ;
        RECT 41.710 172.595 42.000 172.640 ;
        RECT 43.535 172.580 43.855 172.640 ;
        RECT 45.390 172.595 45.680 172.640 ;
        RECT 50.385 172.780 50.675 172.825 ;
        RECT 51.815 172.780 52.135 172.840 ;
        RECT 54.565 172.825 54.780 172.980 ;
        RECT 55.495 172.920 55.815 173.180 ;
        RECT 59.635 173.120 59.955 173.180 ;
        RECT 60.110 173.120 60.400 173.165 ;
        RECT 62.870 173.120 63.160 173.165 ;
        RECT 63.315 173.120 63.635 173.180 ;
        RECT 59.635 172.980 63.635 173.120 ;
        RECT 59.635 172.920 59.955 172.980 ;
        RECT 60.110 172.935 60.400 172.980 ;
        RECT 62.870 172.935 63.160 172.980 ;
        RECT 63.315 172.920 63.635 172.980 ;
        RECT 64.250 173.120 64.540 173.165 ;
        RECT 68.375 173.120 68.695 173.180 ;
        RECT 64.250 172.980 68.695 173.120 ;
        RECT 64.250 172.935 64.540 172.980 ;
        RECT 68.375 172.920 68.695 172.980 ;
        RECT 69.310 172.935 69.600 173.165 ;
        RECT 70.215 173.120 70.535 173.180 ;
        RECT 70.690 173.120 70.980 173.165 ;
        RECT 70.215 172.980 70.980 173.120 ;
        RECT 53.645 172.780 53.935 172.825 ;
        RECT 50.385 172.640 53.935 172.780 ;
        RECT 50.385 172.595 50.675 172.640 ;
        RECT 51.815 172.580 52.135 172.640 ;
        RECT 53.645 172.595 53.935 172.640 ;
        RECT 54.565 172.780 54.855 172.825 ;
        RECT 56.425 172.780 56.715 172.825 ;
        RECT 54.565 172.640 56.715 172.780 ;
        RECT 54.565 172.595 54.855 172.640 ;
        RECT 56.425 172.595 56.715 172.640 ;
        RECT 58.715 172.780 59.035 172.840 ;
        RECT 69.385 172.780 69.525 172.935 ;
        RECT 70.215 172.920 70.535 172.980 ;
        RECT 70.690 172.935 70.980 172.980 ;
        RECT 71.135 172.920 71.455 173.180 ;
        RECT 73.910 173.120 74.200 173.165 ;
        RECT 74.355 173.120 74.675 173.180 ;
        RECT 73.910 172.980 74.675 173.120 ;
        RECT 73.910 172.935 74.200 172.980 ;
        RECT 74.355 172.920 74.675 172.980 ;
        RECT 79.875 173.120 80.195 173.180 ;
        RECT 81.270 173.120 81.560 173.165 ;
        RECT 79.875 172.980 81.560 173.120 ;
        RECT 79.875 172.920 80.195 172.980 ;
        RECT 81.270 172.935 81.560 172.980 ;
        RECT 82.650 172.935 82.940 173.165 ;
        RECT 82.725 172.780 82.865 172.935 ;
        RECT 84.935 172.920 85.255 173.180 ;
        RECT 88.615 173.140 88.935 173.180 ;
        RECT 88.570 172.920 88.935 173.140 ;
        RECT 89.650 173.120 89.940 173.165 ;
        RECT 93.230 173.120 93.520 173.165 ;
        RECT 95.065 173.120 95.355 173.165 ;
        RECT 89.650 172.980 95.355 173.120 ;
        RECT 89.650 172.935 89.940 172.980 ;
        RECT 93.230 172.935 93.520 172.980 ;
        RECT 95.065 172.935 95.355 172.980 ;
        RECT 95.515 172.920 95.835 173.180 ;
        RECT 102.875 173.140 103.195 173.180 ;
        RECT 102.830 172.920 103.195 173.140 ;
        RECT 103.910 173.120 104.200 173.165 ;
        RECT 107.490 173.120 107.780 173.165 ;
        RECT 109.325 173.120 109.615 173.165 ;
        RECT 103.910 172.980 109.615 173.120 ;
        RECT 103.910 172.935 104.200 172.980 ;
        RECT 107.490 172.935 107.780 172.980 ;
        RECT 109.325 172.935 109.615 172.980 ;
        RECT 109.775 172.920 110.095 173.180 ;
        RECT 88.570 172.825 88.860 172.920 ;
        RECT 58.715 172.640 69.525 172.780 ;
        RECT 79.045 172.640 82.865 172.780 ;
        RECT 88.270 172.780 88.860 172.825 ;
        RECT 91.510 172.780 92.160 172.825 ;
        RECT 96.435 172.780 96.755 172.840 ;
        RECT 102.830 172.825 103.120 172.920 ;
        RECT 97.830 172.780 98.120 172.825 ;
        RECT 88.270 172.640 92.160 172.780 ;
        RECT 58.715 172.580 59.035 172.640 ;
        RECT 41.250 172.440 41.540 172.485 ;
        RECT 44.915 172.440 45.235 172.500 ;
        RECT 41.250 172.300 45.235 172.440 ;
        RECT 41.250 172.255 41.540 172.300 ;
        RECT 44.915 172.240 45.235 172.300 ;
        RECT 45.850 172.440 46.140 172.485 ;
        RECT 46.295 172.440 46.615 172.500 ;
        RECT 48.380 172.440 48.670 172.485 ;
        RECT 45.850 172.300 48.670 172.440 ;
        RECT 45.850 172.255 46.140 172.300 ;
        RECT 46.295 172.240 46.615 172.300 ;
        RECT 48.380 172.255 48.670 172.300 ;
        RECT 62.410 172.440 62.700 172.485 ;
        RECT 62.855 172.440 63.175 172.500 ;
        RECT 62.410 172.300 63.175 172.440 ;
        RECT 62.410 172.255 62.700 172.300 ;
        RECT 62.855 172.240 63.175 172.300 ;
        RECT 66.535 172.440 66.855 172.500 ;
        RECT 67.470 172.440 67.760 172.485 ;
        RECT 66.535 172.300 67.760 172.440 ;
        RECT 66.535 172.240 66.855 172.300 ;
        RECT 67.470 172.255 67.760 172.300 ;
        RECT 68.375 172.440 68.695 172.500 ;
        RECT 71.610 172.440 71.900 172.485 ;
        RECT 72.055 172.440 72.375 172.500 ;
        RECT 68.375 172.300 72.375 172.440 ;
        RECT 68.375 172.240 68.695 172.300 ;
        RECT 71.610 172.255 71.900 172.300 ;
        RECT 72.055 172.240 72.375 172.300 ;
        RECT 74.815 172.440 75.135 172.500 ;
        RECT 76.670 172.440 76.960 172.485 ;
        RECT 74.815 172.300 76.960 172.440 ;
        RECT 74.815 172.240 75.135 172.300 ;
        RECT 76.670 172.255 76.960 172.300 ;
        RECT 77.130 172.440 77.420 172.485 ;
        RECT 78.035 172.440 78.355 172.500 ;
        RECT 79.045 172.485 79.185 172.640 ;
        RECT 88.270 172.595 88.560 172.640 ;
        RECT 91.510 172.595 92.160 172.640 ;
        RECT 92.385 172.640 98.120 172.780 ;
        RECT 92.385 172.500 92.525 172.640 ;
        RECT 96.435 172.580 96.755 172.640 ;
        RECT 97.830 172.595 98.120 172.640 ;
        RECT 102.530 172.780 103.120 172.825 ;
        RECT 105.770 172.780 106.420 172.825 ;
        RECT 102.530 172.640 106.420 172.780 ;
        RECT 102.530 172.595 102.820 172.640 ;
        RECT 105.770 172.595 106.420 172.640 ;
        RECT 108.395 172.580 108.715 172.840 ;
        RECT 77.130 172.300 78.355 172.440 ;
        RECT 77.130 172.255 77.420 172.300 ;
        RECT 78.035 172.240 78.355 172.300 ;
        RECT 78.970 172.255 79.260 172.485 ;
        RECT 80.335 172.240 80.655 172.500 ;
        RECT 86.775 172.240 87.095 172.500 ;
        RECT 92.295 172.240 92.615 172.500 ;
        RECT 94.135 172.440 94.455 172.500 ;
        RECT 97.370 172.440 97.660 172.485 ;
        RECT 94.135 172.300 97.660 172.440 ;
        RECT 94.135 172.240 94.455 172.300 ;
        RECT 97.370 172.255 97.660 172.300 ;
        RECT 98.275 172.440 98.595 172.500 ;
        RECT 101.050 172.440 101.340 172.485 ;
        RECT 98.275 172.300 101.340 172.440 ;
        RECT 98.275 172.240 98.595 172.300 ;
        RECT 101.050 172.255 101.340 172.300 ;
        RECT 133.700 172.190 134.930 172.680 ;
        RECT 17.370 171.620 112.465 172.100 ;
        RECT 133.700 171.930 136.690 172.190 ;
        RECT 138.330 171.930 139.470 223.810 ;
        RECT 29.290 171.420 29.580 171.465 ;
        RECT 39.395 171.420 39.715 171.480 ;
        RECT 42.170 171.420 42.460 171.465 ;
        RECT 29.290 171.280 33.185 171.420 ;
        RECT 29.290 171.235 29.580 171.280 ;
        RECT 33.045 171.080 33.185 171.280 ;
        RECT 39.395 171.280 42.460 171.420 ;
        RECT 39.395 171.220 39.715 171.280 ;
        RECT 42.170 171.235 42.460 171.280 ;
        RECT 55.050 171.420 55.340 171.465 ;
        RECT 55.495 171.420 55.815 171.480 ;
        RECT 55.050 171.280 55.815 171.420 ;
        RECT 55.050 171.235 55.340 171.280 ;
        RECT 55.495 171.220 55.815 171.280 ;
        RECT 58.715 171.220 59.035 171.480 ;
        RECT 63.315 171.420 63.635 171.480 ;
        RECT 84.935 171.420 85.255 171.480 ;
        RECT 63.315 171.280 85.255 171.420 ;
        RECT 63.315 171.220 63.635 171.280 ;
        RECT 34.810 171.080 35.100 171.125 ;
        RECT 33.045 170.940 35.100 171.080 ;
        RECT 34.810 170.895 35.100 170.940 ;
        RECT 37.090 171.080 37.740 171.125 ;
        RECT 40.690 171.080 40.980 171.125 ;
        RECT 37.090 170.940 40.980 171.080 ;
        RECT 37.090 170.895 37.740 170.940 ;
        RECT 40.390 170.895 40.980 170.940 ;
        RECT 46.295 171.080 46.615 171.140 ;
        RECT 51.370 171.080 51.660 171.125 ;
        RECT 46.295 170.940 51.660 171.080 ;
        RECT 25.135 170.740 25.455 170.800 ;
        RECT 25.610 170.740 25.900 170.785 ;
        RECT 26.990 170.740 27.280 170.785 ;
        RECT 25.135 170.600 27.280 170.740 ;
        RECT 25.135 170.540 25.455 170.600 ;
        RECT 25.610 170.555 25.900 170.600 ;
        RECT 26.990 170.555 27.280 170.600 ;
        RECT 28.370 170.740 28.660 170.785 ;
        RECT 28.815 170.740 29.135 170.800 ;
        RECT 28.370 170.600 29.135 170.740 ;
        RECT 28.370 170.555 28.660 170.600 ;
        RECT 28.815 170.540 29.135 170.600 ;
        RECT 31.115 170.540 31.435 170.800 ;
        RECT 31.590 170.555 31.880 170.785 ;
        RECT 27.895 170.400 28.215 170.460 ;
        RECT 29.750 170.400 30.040 170.445 ;
        RECT 27.895 170.260 30.040 170.400 ;
        RECT 27.895 170.200 28.215 170.260 ;
        RECT 29.750 170.215 30.040 170.260 ;
        RECT 26.070 170.060 26.360 170.105 ;
        RECT 28.355 170.060 28.675 170.120 ;
        RECT 26.070 169.920 28.675 170.060 ;
        RECT 31.665 170.060 31.805 170.555 ;
        RECT 32.035 170.540 32.355 170.800 ;
        RECT 32.955 170.540 33.275 170.800 ;
        RECT 33.895 170.740 34.185 170.785 ;
        RECT 35.730 170.740 36.020 170.785 ;
        RECT 39.310 170.740 39.600 170.785 ;
        RECT 33.895 170.600 39.600 170.740 ;
        RECT 33.895 170.555 34.185 170.600 ;
        RECT 35.730 170.555 36.020 170.600 ;
        RECT 39.310 170.555 39.600 170.600 ;
        RECT 40.390 170.580 40.680 170.895 ;
        RECT 46.295 170.880 46.615 170.940 ;
        RECT 51.370 170.895 51.660 170.940 ;
        RECT 60.670 171.080 60.960 171.125 ;
        RECT 62.855 171.080 63.175 171.140 ;
        RECT 63.910 171.080 64.560 171.125 ;
        RECT 60.670 170.940 64.560 171.080 ;
        RECT 60.670 170.895 61.260 170.940 ;
        RECT 44.455 170.740 44.775 170.800 ;
        RECT 46.770 170.740 47.060 170.785 ;
        RECT 44.455 170.600 47.060 170.740 ;
        RECT 33.415 170.200 33.735 170.460 ;
        RECT 39.855 170.400 40.175 170.460 ;
        RECT 33.965 170.260 40.175 170.400 ;
        RECT 33.965 170.060 34.105 170.260 ;
        RECT 39.855 170.200 40.175 170.260 ;
        RECT 31.665 169.920 34.105 170.060 ;
        RECT 34.300 170.060 34.590 170.105 ;
        RECT 36.190 170.060 36.480 170.105 ;
        RECT 39.310 170.060 39.600 170.105 ;
        RECT 34.300 169.920 39.600 170.060 ;
        RECT 26.070 169.875 26.360 169.920 ;
        RECT 28.355 169.860 28.675 169.920 ;
        RECT 34.300 169.875 34.590 169.920 ;
        RECT 36.190 169.875 36.480 169.920 ;
        RECT 39.310 169.875 39.600 169.920 ;
        RECT 27.450 169.720 27.740 169.765 ;
        RECT 40.405 169.720 40.545 170.580 ;
        RECT 44.455 170.540 44.775 170.600 ;
        RECT 46.770 170.555 47.060 170.600 ;
        RECT 48.135 170.740 48.455 170.800 ;
        RECT 48.610 170.740 48.900 170.785 ;
        RECT 49.055 170.740 49.375 170.800 ;
        RECT 48.135 170.600 49.375 170.740 ;
        RECT 48.135 170.540 48.455 170.600 ;
        RECT 48.610 170.555 48.900 170.600 ;
        RECT 49.055 170.540 49.375 170.600 ;
        RECT 50.435 170.740 50.755 170.800 ;
        RECT 51.830 170.740 52.120 170.785 ;
        RECT 54.130 170.740 54.420 170.785 ;
        RECT 50.435 170.600 52.120 170.740 ;
        RECT 50.435 170.540 50.755 170.600 ;
        RECT 51.830 170.555 52.120 170.600 ;
        RECT 53.745 170.600 54.420 170.740 ;
        RECT 49.515 170.400 49.835 170.460 ;
        RECT 50.910 170.400 51.200 170.445 ;
        RECT 49.515 170.260 51.200 170.400 ;
        RECT 49.515 170.200 49.835 170.260 ;
        RECT 50.910 170.215 51.200 170.260 ;
        RECT 53.745 170.105 53.885 170.600 ;
        RECT 54.130 170.555 54.420 170.600 ;
        RECT 60.970 170.580 61.260 170.895 ;
        RECT 62.855 170.880 63.175 170.940 ;
        RECT 63.910 170.895 64.560 170.940 ;
        RECT 66.535 170.880 66.855 171.140 ;
        RECT 69.845 171.125 69.985 171.280 ;
        RECT 84.935 171.220 85.255 171.280 ;
        RECT 87.695 171.220 88.015 171.480 ;
        RECT 92.295 171.420 92.615 171.480 ;
        RECT 94.150 171.420 94.440 171.465 ;
        RECT 92.295 171.280 94.440 171.420 ;
        RECT 92.295 171.220 92.615 171.280 ;
        RECT 94.150 171.235 94.440 171.280 ;
        RECT 96.450 171.235 96.740 171.465 ;
        RECT 96.910 171.420 97.200 171.465 ;
        RECT 97.355 171.420 97.675 171.480 ;
        RECT 96.910 171.280 97.675 171.420 ;
        RECT 96.910 171.235 97.200 171.280 ;
        RECT 69.770 170.895 70.060 171.125 ;
        RECT 75.735 171.080 76.055 171.140 ;
        RECT 77.690 171.080 77.980 171.125 ;
        RECT 80.930 171.080 81.580 171.125 ;
        RECT 75.735 170.940 81.580 171.080 ;
        RECT 75.735 170.880 76.055 170.940 ;
        RECT 77.690 170.895 78.280 170.940 ;
        RECT 80.930 170.895 81.580 170.940 ;
        RECT 62.050 170.740 62.340 170.785 ;
        RECT 65.630 170.740 65.920 170.785 ;
        RECT 67.465 170.740 67.755 170.785 ;
        RECT 62.050 170.600 67.755 170.740 ;
        RECT 62.050 170.555 62.340 170.600 ;
        RECT 65.630 170.555 65.920 170.600 ;
        RECT 67.465 170.555 67.755 170.600 ;
        RECT 68.390 170.740 68.680 170.785 ;
        RECT 68.835 170.740 69.155 170.800 ;
        RECT 68.390 170.600 69.155 170.740 ;
        RECT 68.390 170.555 68.680 170.600 ;
        RECT 68.835 170.540 69.155 170.600 ;
        RECT 73.435 170.740 73.755 170.800 ;
        RECT 74.355 170.740 74.675 170.800 ;
        RECT 74.830 170.740 75.120 170.785 ;
        RECT 73.435 170.600 75.120 170.740 ;
        RECT 73.435 170.540 73.755 170.600 ;
        RECT 74.355 170.540 74.675 170.600 ;
        RECT 74.830 170.555 75.120 170.600 ;
        RECT 77.990 170.580 78.280 170.895 ;
        RECT 83.555 170.880 83.875 171.140 ;
        RECT 89.550 171.080 89.840 171.125 ;
        RECT 90.455 171.080 90.775 171.140 ;
        RECT 92.385 171.080 92.525 171.220 ;
        RECT 89.550 170.940 92.525 171.080 ;
        RECT 89.550 170.895 89.840 170.940 ;
        RECT 90.455 170.880 90.775 170.940 ;
        RECT 79.070 170.740 79.360 170.785 ;
        RECT 82.650 170.740 82.940 170.785 ;
        RECT 84.485 170.740 84.775 170.785 ;
        RECT 79.070 170.600 84.775 170.740 ;
        RECT 79.070 170.555 79.360 170.600 ;
        RECT 82.650 170.555 82.940 170.600 ;
        RECT 84.485 170.555 84.775 170.600 ;
        RECT 94.135 170.740 94.455 170.800 ;
        RECT 94.610 170.740 94.900 170.785 ;
        RECT 94.135 170.600 94.900 170.740 ;
        RECT 96.525 170.740 96.665 171.235 ;
        RECT 97.355 171.220 97.675 171.280 ;
        RECT 108.395 171.420 108.715 171.480 ;
        RECT 109.790 171.420 110.080 171.465 ;
        RECT 108.395 171.280 110.080 171.420 ;
        RECT 108.395 171.220 108.715 171.280 ;
        RECT 109.790 171.235 110.080 171.280 ;
        RECT 102.070 171.080 102.360 171.125 ;
        RECT 104.715 171.080 105.035 171.140 ;
        RECT 105.310 171.080 105.960 171.125 ;
        RECT 102.070 170.940 105.960 171.080 ;
        RECT 102.070 170.895 102.660 170.940 ;
        RECT 97.830 170.740 98.120 170.785 ;
        RECT 96.525 170.600 98.120 170.740 ;
        RECT 94.135 170.540 94.455 170.600 ;
        RECT 94.610 170.555 94.900 170.600 ;
        RECT 97.830 170.555 98.120 170.600 ;
        RECT 102.370 170.580 102.660 170.895 ;
        RECT 104.715 170.880 105.035 170.940 ;
        RECT 105.310 170.895 105.960 170.940 ;
        RECT 107.935 170.880 108.255 171.140 ;
        RECT 103.450 170.740 103.740 170.785 ;
        RECT 107.030 170.740 107.320 170.785 ;
        RECT 108.865 170.740 109.155 170.785 ;
        RECT 103.450 170.600 109.155 170.740 ;
        RECT 103.450 170.555 103.740 170.600 ;
        RECT 107.030 170.555 107.320 170.600 ;
        RECT 108.865 170.555 109.155 170.600 ;
        RECT 110.695 170.540 111.015 170.800 ;
        RECT 133.700 170.790 139.470 171.930 ;
        RECT 133.700 170.600 136.690 170.790 ;
        RECT 55.970 170.400 56.260 170.445 ;
        RECT 67.930 170.400 68.220 170.445 ;
        RECT 70.215 170.400 70.535 170.460 ;
        RECT 55.970 170.260 59.405 170.400 ;
        RECT 55.970 170.215 56.260 170.260 ;
        RECT 53.670 169.875 53.960 170.105 ;
        RECT 27.450 169.580 40.545 169.720 ;
        RECT 43.995 169.720 44.315 169.780 ;
        RECT 45.850 169.720 46.140 169.765 ;
        RECT 43.995 169.580 46.140 169.720 ;
        RECT 27.450 169.535 27.740 169.580 ;
        RECT 43.995 169.520 44.315 169.580 ;
        RECT 45.850 169.535 46.140 169.580 ;
        RECT 49.055 169.520 49.375 169.780 ;
        RECT 59.265 169.765 59.405 170.260 ;
        RECT 67.930 170.260 70.535 170.400 ;
        RECT 67.930 170.215 68.220 170.260 ;
        RECT 70.215 170.200 70.535 170.260 ;
        RECT 80.795 170.400 81.115 170.460 ;
        RECT 83.095 170.400 83.415 170.460 ;
        RECT 84.950 170.400 85.240 170.445 ;
        RECT 80.795 170.260 85.240 170.400 ;
        RECT 80.795 170.200 81.115 170.260 ;
        RECT 83.095 170.200 83.415 170.260 ;
        RECT 84.950 170.215 85.240 170.260 ;
        RECT 86.775 170.400 87.095 170.460 ;
        RECT 90.010 170.400 90.300 170.445 ;
        RECT 86.775 170.260 90.300 170.400 ;
        RECT 86.775 170.200 87.095 170.260 ;
        RECT 90.010 170.215 90.300 170.260 ;
        RECT 90.470 170.400 90.760 170.445 ;
        RECT 91.375 170.400 91.695 170.460 ;
        RECT 93.230 170.400 93.520 170.445 ;
        RECT 90.470 170.260 93.520 170.400 ;
        RECT 90.470 170.215 90.760 170.260 ;
        RECT 62.050 170.060 62.340 170.105 ;
        RECT 65.170 170.060 65.460 170.105 ;
        RECT 67.060 170.060 67.350 170.105 ;
        RECT 62.050 169.920 67.350 170.060 ;
        RECT 62.050 169.875 62.340 169.920 ;
        RECT 65.170 169.875 65.460 169.920 ;
        RECT 67.060 169.875 67.350 169.920 ;
        RECT 74.355 170.060 74.675 170.120 ;
        RECT 76.210 170.060 76.500 170.105 ;
        RECT 74.355 169.920 76.500 170.060 ;
        RECT 74.355 169.860 74.675 169.920 ;
        RECT 76.210 169.875 76.500 169.920 ;
        RECT 79.070 170.060 79.360 170.105 ;
        RECT 82.190 170.060 82.480 170.105 ;
        RECT 84.080 170.060 84.370 170.105 ;
        RECT 79.070 169.920 84.370 170.060 ;
        RECT 79.070 169.875 79.360 169.920 ;
        RECT 82.190 169.875 82.480 169.920 ;
        RECT 84.080 169.875 84.370 169.920 ;
        RECT 59.190 169.720 59.480 169.765 ;
        RECT 63.775 169.720 64.095 169.780 ;
        RECT 59.190 169.580 64.095 169.720 ;
        RECT 59.190 169.535 59.480 169.580 ;
        RECT 63.775 169.520 64.095 169.580 ;
        RECT 75.275 169.520 75.595 169.780 ;
        RECT 78.495 169.720 78.815 169.780 ;
        RECT 90.545 169.720 90.685 170.215 ;
        RECT 91.375 170.200 91.695 170.260 ;
        RECT 93.230 170.215 93.520 170.260 ;
        RECT 95.515 170.400 95.835 170.460 ;
        RECT 109.330 170.400 109.620 170.445 ;
        RECT 109.775 170.400 110.095 170.460 ;
        RECT 95.515 170.260 110.095 170.400 ;
        RECT 95.515 170.200 95.835 170.260 ;
        RECT 109.330 170.215 109.620 170.260 ;
        RECT 109.775 170.200 110.095 170.260 ;
        RECT 133.700 170.120 134.930 170.600 ;
        RECT 103.450 170.060 103.740 170.105 ;
        RECT 106.570 170.060 106.860 170.105 ;
        RECT 108.460 170.060 108.750 170.105 ;
        RECT 103.450 169.920 108.750 170.060 ;
        RECT 103.450 169.875 103.740 169.920 ;
        RECT 106.570 169.875 106.860 169.920 ;
        RECT 108.460 169.875 108.750 169.920 ;
        RECT 78.495 169.580 90.685 169.720 ;
        RECT 99.195 169.720 99.515 169.780 ;
        RECT 100.590 169.720 100.880 169.765 ;
        RECT 99.195 169.580 100.880 169.720 ;
        RECT 78.495 169.520 78.815 169.580 ;
        RECT 99.195 169.520 99.515 169.580 ;
        RECT 100.590 169.535 100.880 169.580 ;
        RECT 18.165 168.900 112.465 169.380 ;
        RECT 38.475 168.700 38.795 168.760 ;
        RECT 45.850 168.700 46.140 168.745 ;
        RECT 38.475 168.560 46.140 168.700 ;
        RECT 38.475 168.500 38.795 168.560 ;
        RECT 45.850 168.515 46.140 168.560 ;
        RECT 78.495 168.700 78.815 168.760 ;
        RECT 83.555 168.700 83.875 168.760 ;
        RECT 86.790 168.700 87.080 168.745 ;
        RECT 95.515 168.700 95.835 168.760 ;
        RECT 78.495 168.560 82.405 168.700 ;
        RECT 78.495 168.500 78.815 168.560 ;
        RECT 26.480 168.360 26.770 168.405 ;
        RECT 28.370 168.360 28.660 168.405 ;
        RECT 31.490 168.360 31.780 168.405 ;
        RECT 26.480 168.220 31.780 168.360 ;
        RECT 26.480 168.175 26.770 168.220 ;
        RECT 28.370 168.175 28.660 168.220 ;
        RECT 31.490 168.175 31.780 168.220 ;
        RECT 39.510 168.360 39.800 168.405 ;
        RECT 42.630 168.360 42.920 168.405 ;
        RECT 44.520 168.360 44.810 168.405 ;
        RECT 57.335 168.360 57.655 168.420 ;
        RECT 39.510 168.220 44.810 168.360 ;
        RECT 39.510 168.175 39.800 168.220 ;
        RECT 42.630 168.175 42.920 168.220 ;
        RECT 44.520 168.175 44.810 168.220 ;
        RECT 45.465 168.220 57.655 168.360 ;
        RECT 32.955 168.020 33.275 168.080 ;
        RECT 40.315 168.020 40.635 168.080 ;
        RECT 32.955 167.880 40.635 168.020 ;
        RECT 32.955 167.820 33.275 167.880 ;
        RECT 40.315 167.820 40.635 167.880 ;
        RECT 43.995 167.820 44.315 168.080 ;
        RECT 45.465 168.065 45.605 168.220 ;
        RECT 57.335 168.160 57.655 168.220 ;
        RECT 75.850 168.360 76.140 168.405 ;
        RECT 78.970 168.360 79.260 168.405 ;
        RECT 80.860 168.360 81.150 168.405 ;
        RECT 75.850 168.220 81.150 168.360 ;
        RECT 75.850 168.175 76.140 168.220 ;
        RECT 78.970 168.175 79.260 168.220 ;
        RECT 80.860 168.175 81.150 168.220 ;
        RECT 45.390 167.835 45.680 168.065 ;
        RECT 46.755 168.020 47.075 168.080 ;
        RECT 49.515 168.020 49.835 168.080 ;
        RECT 50.910 168.020 51.200 168.065 ;
        RECT 46.755 167.880 49.285 168.020 ;
        RECT 46.755 167.820 47.075 167.880 ;
        RECT 25.595 167.480 25.915 167.740 ;
        RECT 26.075 167.680 26.365 167.725 ;
        RECT 27.910 167.680 28.200 167.725 ;
        RECT 31.490 167.680 31.780 167.725 ;
        RECT 26.075 167.540 31.780 167.680 ;
        RECT 26.075 167.495 26.365 167.540 ;
        RECT 27.910 167.495 28.200 167.540 ;
        RECT 31.490 167.495 31.780 167.540 ;
        RECT 26.975 167.140 27.295 167.400 ;
        RECT 28.355 167.340 28.675 167.400 ;
        RECT 32.570 167.385 32.860 167.700 ;
        RECT 36.175 167.480 36.495 167.740 ;
        RECT 38.430 167.385 38.720 167.700 ;
        RECT 39.510 167.680 39.800 167.725 ;
        RECT 43.090 167.680 43.380 167.725 ;
        RECT 44.925 167.680 45.215 167.725 ;
        RECT 39.510 167.540 45.215 167.680 ;
        RECT 39.510 167.495 39.800 167.540 ;
        RECT 43.090 167.495 43.380 167.540 ;
        RECT 44.925 167.495 45.215 167.540 ;
        RECT 47.215 167.480 47.535 167.740 ;
        RECT 47.675 167.480 47.995 167.740 ;
        RECT 49.145 167.725 49.285 167.880 ;
        RECT 49.515 167.880 51.200 168.020 ;
        RECT 49.515 167.820 49.835 167.880 ;
        RECT 50.910 167.835 51.200 167.880 ;
        RECT 71.610 168.020 71.900 168.065 ;
        RECT 73.435 168.020 73.755 168.080 ;
        RECT 71.610 167.880 73.755 168.020 ;
        RECT 71.610 167.835 71.900 167.880 ;
        RECT 73.435 167.820 73.755 167.880 ;
        RECT 80.335 167.820 80.655 168.080 ;
        RECT 82.265 168.020 82.405 168.560 ;
        RECT 83.555 168.560 87.080 168.700 ;
        RECT 83.555 168.500 83.875 168.560 ;
        RECT 86.790 168.515 87.080 168.560 ;
        RECT 91.925 168.560 95.835 168.700 ;
        RECT 85.870 168.175 86.160 168.405 ;
        RECT 82.650 168.020 82.940 168.065 ;
        RECT 82.265 167.880 82.940 168.020 ;
        RECT 82.650 167.835 82.940 167.880 ;
        RECT 48.150 167.495 48.440 167.725 ;
        RECT 49.070 167.495 49.360 167.725 ;
        RECT 55.050 167.680 55.340 167.725 ;
        RECT 54.205 167.540 55.340 167.680 ;
        RECT 29.270 167.340 29.920 167.385 ;
        RECT 32.570 167.340 33.160 167.385 ;
        RECT 28.355 167.200 33.160 167.340 ;
        RECT 28.355 167.140 28.675 167.200 ;
        RECT 29.270 167.155 29.920 167.200 ;
        RECT 32.870 167.155 33.160 167.200 ;
        RECT 38.130 167.340 38.720 167.385 ;
        RECT 38.935 167.340 39.255 167.400 ;
        RECT 41.370 167.340 42.020 167.385 ;
        RECT 48.225 167.340 48.365 167.495 ;
        RECT 38.130 167.200 42.020 167.340 ;
        RECT 38.130 167.155 38.420 167.200 ;
        RECT 38.935 167.140 39.255 167.200 ;
        RECT 41.370 167.155 42.020 167.200 ;
        RECT 47.765 167.200 48.365 167.340 ;
        RECT 48.595 167.340 48.915 167.400 ;
        RECT 52.290 167.340 52.580 167.385 ;
        RECT 48.595 167.200 52.580 167.340 ;
        RECT 34.335 166.800 34.655 167.060 ;
        RECT 35.255 166.800 35.575 167.060 ;
        RECT 36.635 166.800 36.955 167.060 ;
        RECT 39.395 167.000 39.715 167.060 ;
        RECT 47.765 167.000 47.905 167.200 ;
        RECT 48.595 167.140 48.915 167.200 ;
        RECT 52.290 167.155 52.580 167.200 ;
        RECT 39.395 166.860 47.905 167.000 ;
        RECT 50.435 167.000 50.755 167.060 ;
        RECT 54.205 167.045 54.345 167.540 ;
        RECT 55.050 167.495 55.340 167.540 ;
        RECT 61.015 167.680 61.335 167.740 ;
        RECT 68.835 167.680 69.155 167.740 ;
        RECT 70.230 167.680 70.520 167.725 ;
        RECT 61.015 167.540 70.520 167.680 ;
        RECT 61.015 167.480 61.335 167.540 ;
        RECT 68.835 167.480 69.155 167.540 ;
        RECT 70.230 167.495 70.520 167.540 ;
        RECT 74.770 167.385 75.060 167.700 ;
        RECT 75.850 167.680 76.140 167.725 ;
        RECT 79.430 167.680 79.720 167.725 ;
        RECT 81.265 167.680 81.555 167.725 ;
        RECT 75.850 167.540 81.555 167.680 ;
        RECT 75.850 167.495 76.140 167.540 ;
        RECT 79.430 167.495 79.720 167.540 ;
        RECT 81.265 167.495 81.555 167.540 ;
        RECT 81.730 167.495 82.020 167.725 ;
        RECT 85.945 167.680 86.085 168.175 ;
        RECT 89.995 168.020 90.315 168.080 ;
        RECT 89.995 167.880 90.685 168.020 ;
        RECT 89.995 167.820 90.315 167.880 ;
        RECT 90.545 167.725 90.685 167.880 ;
        RECT 91.925 167.725 92.065 168.560 ;
        RECT 95.515 168.500 95.835 168.560 ;
        RECT 106.570 168.700 106.860 168.745 ;
        RECT 107.935 168.700 108.255 168.760 ;
        RECT 106.570 168.560 108.255 168.700 ;
        RECT 106.570 168.515 106.860 168.560 ;
        RECT 107.935 168.500 108.255 168.560 ;
        RECT 92.720 168.360 93.010 168.405 ;
        RECT 94.610 168.360 94.900 168.405 ;
        RECT 97.730 168.360 98.020 168.405 ;
        RECT 92.720 168.220 98.020 168.360 ;
        RECT 92.720 168.175 93.010 168.220 ;
        RECT 94.610 168.175 94.900 168.220 ;
        RECT 97.730 168.175 98.020 168.220 ;
        RECT 104.730 168.360 105.020 168.405 ;
        RECT 110.695 168.360 111.015 168.420 ;
        RECT 104.730 168.220 111.015 168.360 ;
        RECT 104.730 168.175 105.020 168.220 ;
        RECT 110.695 168.160 111.015 168.220 ;
        RECT 100.115 168.020 100.435 168.080 ;
        RECT 100.590 168.020 100.880 168.065 ;
        RECT 100.115 167.880 100.880 168.020 ;
        RECT 100.115 167.820 100.435 167.880 ;
        RECT 100.590 167.835 100.880 167.880 ;
        RECT 101.035 168.020 101.355 168.080 ;
        RECT 101.510 168.020 101.800 168.065 ;
        RECT 101.035 167.880 101.800 168.020 ;
        RECT 101.035 167.820 101.355 167.880 ;
        RECT 101.510 167.835 101.800 167.880 ;
        RECT 87.710 167.680 88.000 167.725 ;
        RECT 85.945 167.540 88.000 167.680 ;
        RECT 87.710 167.495 88.000 167.540 ;
        RECT 89.090 167.680 89.380 167.725 ;
        RECT 90.470 167.680 90.760 167.725 ;
        RECT 89.090 167.540 90.760 167.680 ;
        RECT 89.090 167.495 89.380 167.540 ;
        RECT 90.470 167.495 90.760 167.540 ;
        RECT 91.850 167.495 92.140 167.725 ;
        RECT 92.315 167.680 92.605 167.725 ;
        RECT 94.150 167.680 94.440 167.725 ;
        RECT 97.730 167.680 98.020 167.725 ;
        RECT 92.315 167.540 98.020 167.680 ;
        RECT 92.315 167.495 92.605 167.540 ;
        RECT 94.150 167.495 94.440 167.540 ;
        RECT 97.730 167.495 98.020 167.540 ;
        RECT 74.470 167.340 75.060 167.385 ;
        RECT 75.275 167.340 75.595 167.400 ;
        RECT 77.710 167.340 78.360 167.385 ;
        RECT 74.470 167.200 78.360 167.340 ;
        RECT 74.470 167.155 74.760 167.200 ;
        RECT 75.275 167.140 75.595 167.200 ;
        RECT 77.710 167.155 78.360 167.200 ;
        RECT 80.795 167.340 81.115 167.400 ;
        RECT 81.805 167.340 81.945 167.495 ;
        RECT 80.795 167.200 81.945 167.340 ;
        RECT 89.995 167.340 90.315 167.400 ;
        RECT 91.925 167.340 92.065 167.495 ;
        RECT 89.995 167.200 92.065 167.340 ;
        RECT 80.795 167.140 81.115 167.200 ;
        RECT 89.995 167.140 90.315 167.200 ;
        RECT 93.215 167.140 93.535 167.400 ;
        RECT 98.810 167.385 99.100 167.700 ;
        RECT 103.795 167.680 104.115 167.740 ;
        RECT 105.650 167.680 105.940 167.725 ;
        RECT 103.795 167.540 105.940 167.680 ;
        RECT 103.795 167.480 104.115 167.540 ;
        RECT 105.650 167.495 105.940 167.540 ;
        RECT 95.510 167.340 96.160 167.385 ;
        RECT 98.810 167.340 99.400 167.385 ;
        RECT 94.685 167.200 99.400 167.340 ;
        RECT 51.830 167.000 52.120 167.045 ;
        RECT 50.435 166.860 52.120 167.000 ;
        RECT 39.395 166.800 39.715 166.860 ;
        RECT 50.435 166.800 50.755 166.860 ;
        RECT 51.830 166.815 52.120 166.860 ;
        RECT 54.130 166.815 54.420 167.045 ;
        RECT 55.970 167.000 56.260 167.045 ;
        RECT 56.875 167.000 57.195 167.060 ;
        RECT 55.970 166.860 57.195 167.000 ;
        RECT 55.970 166.815 56.260 166.860 ;
        RECT 56.875 166.800 57.195 166.860 ;
        RECT 71.135 167.000 71.455 167.060 ;
        RECT 72.990 167.000 73.280 167.045 ;
        RECT 71.135 166.860 73.280 167.000 ;
        RECT 71.135 166.800 71.455 166.860 ;
        RECT 72.990 166.815 73.280 166.860 ;
        RECT 80.335 167.000 80.655 167.060 ;
        RECT 83.570 167.000 83.860 167.045 ;
        RECT 80.335 166.860 83.860 167.000 ;
        RECT 80.335 166.800 80.655 166.860 ;
        RECT 83.570 166.815 83.860 166.860 ;
        RECT 84.030 167.000 84.320 167.045 ;
        RECT 86.775 167.000 87.095 167.060 ;
        RECT 84.030 166.860 87.095 167.000 ;
        RECT 84.030 166.815 84.320 166.860 ;
        RECT 86.775 166.800 87.095 166.860 ;
        RECT 87.695 167.000 88.015 167.060 ;
        RECT 88.630 167.000 88.920 167.045 ;
        RECT 87.695 166.860 88.920 167.000 ;
        RECT 87.695 166.800 88.015 166.860 ;
        RECT 88.630 166.815 88.920 166.860 ;
        RECT 90.930 167.000 91.220 167.045 ;
        RECT 94.685 167.000 94.825 167.200 ;
        RECT 95.510 167.155 96.160 167.200 ;
        RECT 99.110 167.155 99.400 167.200 ;
        RECT 100.575 167.340 100.895 167.400 ;
        RECT 102.890 167.340 103.180 167.385 ;
        RECT 100.575 167.200 103.180 167.340 ;
        RECT 100.575 167.140 100.895 167.200 ;
        RECT 102.890 167.155 103.180 167.200 ;
        RECT 90.930 166.860 94.825 167.000 ;
        RECT 98.275 167.000 98.595 167.060 ;
        RECT 102.430 167.000 102.720 167.045 ;
        RECT 98.275 166.860 102.720 167.000 ;
        RECT 90.930 166.815 91.220 166.860 ;
        RECT 98.275 166.800 98.595 166.860 ;
        RECT 102.430 166.815 102.720 166.860 ;
        RECT 17.370 166.180 112.465 166.660 ;
        RECT 23.310 165.980 23.600 166.025 ;
        RECT 26.975 165.980 27.295 166.040 ;
        RECT 36.635 165.980 36.955 166.040 ;
        RECT 42.170 165.980 42.460 166.025 ;
        RECT 23.310 165.840 27.295 165.980 ;
        RECT 23.310 165.795 23.600 165.840 ;
        RECT 26.975 165.780 27.295 165.840 ;
        RECT 35.805 165.840 42.460 165.980 ;
        RECT 21.455 165.640 21.775 165.700 ;
        RECT 27.435 165.685 27.755 165.700 ;
        RECT 25.150 165.640 25.440 165.685 ;
        RECT 21.455 165.500 25.440 165.640 ;
        RECT 21.455 165.440 21.775 165.500 ;
        RECT 25.150 165.455 25.440 165.500 ;
        RECT 27.430 165.640 28.080 165.685 ;
        RECT 31.030 165.640 31.320 165.685 ;
        RECT 27.430 165.500 31.320 165.640 ;
        RECT 27.430 165.455 28.080 165.500 ;
        RECT 30.730 165.455 31.320 165.500 ;
        RECT 27.435 165.440 27.755 165.455 ;
        RECT 22.390 165.115 22.680 165.345 ;
        RECT 24.235 165.300 24.525 165.345 ;
        RECT 26.070 165.300 26.360 165.345 ;
        RECT 29.650 165.300 29.940 165.345 ;
        RECT 24.235 165.160 29.940 165.300 ;
        RECT 24.235 165.115 24.525 165.160 ;
        RECT 26.070 165.115 26.360 165.160 ;
        RECT 29.650 165.115 29.940 165.160 ;
        RECT 30.730 165.140 31.020 165.455 ;
        RECT 32.495 165.300 32.815 165.360 ;
        RECT 33.430 165.300 33.720 165.345 ;
        RECT 35.805 165.300 35.945 165.840 ;
        RECT 36.635 165.780 36.955 165.840 ;
        RECT 42.170 165.795 42.460 165.840 ;
        RECT 44.455 165.780 44.775 166.040 ;
        RECT 67.455 165.980 67.775 166.040 ;
        RECT 68.375 165.980 68.695 166.040 ;
        RECT 71.595 165.980 71.915 166.040 ;
        RECT 67.455 165.840 71.915 165.980 ;
        RECT 67.455 165.780 67.775 165.840 ;
        RECT 68.375 165.780 68.695 165.840 ;
        RECT 71.595 165.780 71.915 165.840 ;
        RECT 75.290 165.980 75.580 166.025 ;
        RECT 75.735 165.980 76.055 166.040 ;
        RECT 75.290 165.840 76.055 165.980 ;
        RECT 75.290 165.795 75.580 165.840 ;
        RECT 75.735 165.780 76.055 165.840 ;
        RECT 79.875 165.780 80.195 166.040 ;
        RECT 83.555 165.980 83.875 166.040 ;
        RECT 85.410 165.980 85.700 166.025 ;
        RECT 86.315 165.980 86.635 166.040 ;
        RECT 96.450 165.980 96.740 166.025 ;
        RECT 83.555 165.840 96.740 165.980 ;
        RECT 83.555 165.780 83.875 165.840 ;
        RECT 85.410 165.795 85.700 165.840 ;
        RECT 86.315 165.780 86.635 165.840 ;
        RECT 96.450 165.795 96.740 165.840 ;
        RECT 103.795 165.780 104.115 166.040 ;
        RECT 36.190 165.640 36.480 165.685 ;
        RECT 38.490 165.640 38.780 165.685 ;
        RECT 36.190 165.500 38.780 165.640 ;
        RECT 36.190 165.455 36.480 165.500 ;
        RECT 38.490 165.455 38.780 165.500 ;
        RECT 39.855 165.640 40.175 165.700 ;
        RECT 47.675 165.640 47.995 165.700 ;
        RECT 39.855 165.500 47.995 165.640 ;
        RECT 39.855 165.440 40.175 165.500 ;
        RECT 47.675 165.440 47.995 165.500 ;
        RECT 49.055 165.640 49.375 165.700 ;
        RECT 52.225 165.640 52.515 165.685 ;
        RECT 55.485 165.640 55.775 165.685 ;
        RECT 49.055 165.500 55.775 165.640 ;
        RECT 49.055 165.440 49.375 165.500 ;
        RECT 52.225 165.455 52.515 165.500 ;
        RECT 55.485 165.455 55.775 165.500 ;
        RECT 56.405 165.640 56.695 165.685 ;
        RECT 58.265 165.640 58.555 165.685 ;
        RECT 70.675 165.640 70.995 165.700 ;
        RECT 74.355 165.640 74.675 165.700 ;
        RECT 78.050 165.640 78.340 165.685 ;
        RECT 80.335 165.640 80.655 165.700 ;
        RECT 56.405 165.500 58.555 165.640 ;
        RECT 56.405 165.455 56.695 165.500 ;
        RECT 58.265 165.455 58.555 165.500 ;
        RECT 68.005 165.500 70.445 165.640 ;
        RECT 32.495 165.160 35.945 165.300 ;
        RECT 42.630 165.300 42.920 165.345 ;
        RECT 44.915 165.300 45.235 165.360 ;
        RECT 42.630 165.160 45.235 165.300 ;
        RECT 22.465 164.280 22.605 165.115 ;
        RECT 32.495 165.100 32.815 165.160 ;
        RECT 33.430 165.115 33.720 165.160 ;
        RECT 42.630 165.115 42.920 165.160 ;
        RECT 44.915 165.100 45.235 165.160 ;
        RECT 46.310 165.300 46.600 165.345 ;
        RECT 48.135 165.300 48.455 165.360 ;
        RECT 50.895 165.300 51.215 165.360 ;
        RECT 46.310 165.160 51.215 165.300 ;
        RECT 46.310 165.115 46.600 165.160 ;
        RECT 48.135 165.100 48.455 165.160 ;
        RECT 50.895 165.100 51.215 165.160 ;
        RECT 54.085 165.300 54.375 165.345 ;
        RECT 56.405 165.300 56.620 165.455 ;
        RECT 68.005 165.360 68.145 165.500 ;
        RECT 54.085 165.160 56.620 165.300 ;
        RECT 56.875 165.300 57.195 165.360 ;
        RECT 57.350 165.300 57.640 165.345 ;
        RECT 56.875 165.160 57.640 165.300 ;
        RECT 54.085 165.115 54.375 165.160 ;
        RECT 56.875 165.100 57.195 165.160 ;
        RECT 57.350 165.115 57.640 165.160 ;
        RECT 57.795 165.300 58.115 165.360 ;
        RECT 59.190 165.300 59.480 165.345 ;
        RECT 57.795 165.160 59.480 165.300 ;
        RECT 57.795 165.100 58.115 165.160 ;
        RECT 59.190 165.115 59.480 165.160 ;
        RECT 60.095 165.300 60.415 165.360 ;
        RECT 60.570 165.300 60.860 165.345 ;
        RECT 61.015 165.300 61.335 165.360 ;
        RECT 60.095 165.160 61.335 165.300 ;
        RECT 60.095 165.100 60.415 165.160 ;
        RECT 60.570 165.115 60.860 165.160 ;
        RECT 61.015 165.100 61.335 165.160 ;
        RECT 63.775 165.300 64.095 165.360 ;
        RECT 64.710 165.300 65.000 165.345 ;
        RECT 67.010 165.300 67.300 165.345 ;
        RECT 63.775 165.160 67.300 165.300 ;
        RECT 63.775 165.100 64.095 165.160 ;
        RECT 64.710 165.115 65.000 165.160 ;
        RECT 67.010 165.115 67.300 165.160 ;
        RECT 67.915 165.100 68.235 165.360 ;
        RECT 68.375 165.100 68.695 165.360 ;
        RECT 69.755 165.100 70.075 165.360 ;
        RECT 70.305 165.345 70.445 165.500 ;
        RECT 70.675 165.500 80.655 165.640 ;
        RECT 70.675 165.440 70.995 165.500 ;
        RECT 74.355 165.440 74.675 165.500 ;
        RECT 78.050 165.455 78.340 165.500 ;
        RECT 80.335 165.440 80.655 165.500 ;
        RECT 86.890 165.640 87.180 165.685 ;
        RECT 87.695 165.640 88.015 165.700 ;
        RECT 90.130 165.640 90.780 165.685 ;
        RECT 86.890 165.500 90.780 165.640 ;
        RECT 86.890 165.455 87.480 165.500 ;
        RECT 70.230 165.115 70.520 165.345 ;
        RECT 71.150 165.300 71.440 165.345 ;
        RECT 71.595 165.300 71.915 165.360 ;
        RECT 71.150 165.160 71.915 165.300 ;
        RECT 71.150 165.115 71.440 165.160 ;
        RECT 71.595 165.100 71.915 165.160 ;
        RECT 73.435 165.300 73.755 165.360 ;
        RECT 74.830 165.300 75.120 165.345 ;
        RECT 78.495 165.300 78.815 165.360 ;
        RECT 73.435 165.160 75.120 165.300 ;
        RECT 73.435 165.100 73.755 165.160 ;
        RECT 74.830 165.115 75.120 165.160 ;
        RECT 77.205 165.160 78.815 165.300 ;
        RECT 23.770 164.960 24.060 165.005 ;
        RECT 25.595 164.960 25.915 165.020 ;
        RECT 31.575 164.960 31.895 165.020 ;
        RECT 23.770 164.820 31.895 164.960 ;
        RECT 23.770 164.775 24.060 164.820 ;
        RECT 25.595 164.760 25.915 164.820 ;
        RECT 31.575 164.760 31.895 164.820 ;
        RECT 37.095 164.960 37.415 165.020 ;
        RECT 38.950 164.960 39.240 165.005 ;
        RECT 39.395 164.960 39.715 165.020 ;
        RECT 37.095 164.820 39.715 164.960 ;
        RECT 37.095 164.760 37.415 164.820 ;
        RECT 38.950 164.775 39.240 164.820 ;
        RECT 39.395 164.760 39.715 164.820 ;
        RECT 39.870 164.960 40.160 165.005 ;
        RECT 41.250 164.960 41.540 165.005 ;
        RECT 49.055 164.960 49.375 165.020 ;
        RECT 50.435 165.005 50.755 165.020 ;
        RECT 39.870 164.820 49.375 164.960 ;
        RECT 39.870 164.775 40.160 164.820 ;
        RECT 41.250 164.775 41.540 164.820 ;
        RECT 24.640 164.620 24.930 164.665 ;
        RECT 26.530 164.620 26.820 164.665 ;
        RECT 29.650 164.620 29.940 164.665 ;
        RECT 24.640 164.480 29.940 164.620 ;
        RECT 24.640 164.435 24.930 164.480 ;
        RECT 26.530 164.435 26.820 164.480 ;
        RECT 29.650 164.435 29.940 164.480 ;
        RECT 32.510 164.620 32.800 164.665 ;
        RECT 37.555 164.620 37.875 164.680 ;
        RECT 32.510 164.480 37.875 164.620 ;
        RECT 32.510 164.435 32.800 164.480 ;
        RECT 37.555 164.420 37.875 164.480 ;
        RECT 38.015 164.620 38.335 164.680 ;
        RECT 39.945 164.620 40.085 164.775 ;
        RECT 49.055 164.760 49.375 164.820 ;
        RECT 50.220 164.775 50.755 165.005 ;
        RECT 50.435 164.760 50.755 164.775 ;
        RECT 62.395 164.960 62.715 165.020 ;
        RECT 67.470 164.960 67.760 165.005 ;
        RECT 69.845 164.960 69.985 165.100 ;
        RECT 62.395 164.820 69.985 164.960 ;
        RECT 70.690 164.960 70.980 165.005 ;
        RECT 72.055 164.960 72.375 165.020 ;
        RECT 70.690 164.820 72.375 164.960 ;
        RECT 62.395 164.760 62.715 164.820 ;
        RECT 67.470 164.775 67.760 164.820 ;
        RECT 70.690 164.775 70.980 164.820 ;
        RECT 38.015 164.480 40.085 164.620 ;
        RECT 54.085 164.620 54.375 164.665 ;
        RECT 56.865 164.620 57.155 164.665 ;
        RECT 58.725 164.620 59.015 164.665 ;
        RECT 54.085 164.480 59.015 164.620 ;
        RECT 38.015 164.420 38.335 164.480 ;
        RECT 54.085 164.435 54.375 164.480 ;
        RECT 56.865 164.435 57.155 164.480 ;
        RECT 58.725 164.435 59.015 164.480 ;
        RECT 65.170 164.620 65.460 164.665 ;
        RECT 66.535 164.620 66.855 164.680 ;
        RECT 65.170 164.480 66.855 164.620 ;
        RECT 65.170 164.435 65.460 164.480 ;
        RECT 66.535 164.420 66.855 164.480 ;
        RECT 68.375 164.620 68.695 164.680 ;
        RECT 70.765 164.620 70.905 164.775 ;
        RECT 72.055 164.760 72.375 164.820 ;
        RECT 75.735 164.960 76.055 165.020 ;
        RECT 76.670 164.960 76.960 165.005 ;
        RECT 77.205 164.960 77.345 165.160 ;
        RECT 78.495 165.100 78.815 165.160 ;
        RECT 80.795 165.100 81.115 165.360 ;
        RECT 84.490 165.115 84.780 165.345 ;
        RECT 87.190 165.140 87.480 165.455 ;
        RECT 87.695 165.440 88.015 165.500 ;
        RECT 90.130 165.455 90.780 165.500 ;
        RECT 92.755 165.440 93.075 165.700 ;
        RECT 100.115 165.640 100.435 165.700 ;
        RECT 101.970 165.640 102.260 165.685 ;
        RECT 96.985 165.500 102.260 165.640 ;
        RECT 88.270 165.300 88.560 165.345 ;
        RECT 91.850 165.300 92.140 165.345 ;
        RECT 93.685 165.300 93.975 165.345 ;
        RECT 88.270 165.160 93.975 165.300 ;
        RECT 88.270 165.115 88.560 165.160 ;
        RECT 91.850 165.115 92.140 165.160 ;
        RECT 93.685 165.115 93.975 165.160 ;
        RECT 75.735 164.820 77.345 164.960 ;
        RECT 77.590 164.960 77.880 165.005 ;
        RECT 78.035 164.960 78.355 165.020 ;
        RECT 77.590 164.820 78.355 164.960 ;
        RECT 84.565 164.960 84.705 165.115 ;
        RECT 87.695 164.960 88.015 165.020 ;
        RECT 84.565 164.820 88.015 164.960 ;
        RECT 75.735 164.760 76.055 164.820 ;
        RECT 76.670 164.775 76.960 164.820 ;
        RECT 77.590 164.775 77.880 164.820 ;
        RECT 68.375 164.480 70.905 164.620 ;
        RECT 71.135 164.620 71.455 164.680 ;
        RECT 77.665 164.620 77.805 164.775 ;
        RECT 78.035 164.760 78.355 164.820 ;
        RECT 87.695 164.760 88.015 164.820 ;
        RECT 89.995 164.960 90.315 165.020 ;
        RECT 94.150 164.960 94.440 165.005 ;
        RECT 89.995 164.820 94.440 164.960 ;
        RECT 89.995 164.760 90.315 164.820 ;
        RECT 94.150 164.775 94.440 164.820 ;
        RECT 96.435 164.960 96.755 165.020 ;
        RECT 96.985 165.005 97.125 165.500 ;
        RECT 100.115 165.440 100.435 165.500 ;
        RECT 101.970 165.455 102.260 165.500 ;
        RECT 135.580 165.470 136.830 166.590 ;
        RECT 99.195 165.300 99.515 165.360 ;
        RECT 100.575 165.300 100.895 165.360 ;
        RECT 101.510 165.300 101.800 165.345 ;
        RECT 99.195 165.160 101.800 165.300 ;
        RECT 99.195 165.100 99.515 165.160 ;
        RECT 100.575 165.100 100.895 165.160 ;
        RECT 101.510 165.115 101.800 165.160 ;
        RECT 104.255 165.100 104.575 165.360 ;
        RECT 106.555 165.100 106.875 165.360 ;
        RECT 96.910 164.960 97.200 165.005 ;
        RECT 96.435 164.820 97.200 164.960 ;
        RECT 96.435 164.760 96.755 164.820 ;
        RECT 96.910 164.775 97.200 164.820 ;
        RECT 97.815 164.960 98.135 165.020 ;
        RECT 101.035 164.960 101.355 165.020 ;
        RECT 97.815 164.820 101.355 164.960 ;
        RECT 97.815 164.760 98.135 164.820 ;
        RECT 101.035 164.760 101.355 164.820 ;
        RECT 71.135 164.480 77.805 164.620 ;
        RECT 88.270 164.620 88.560 164.665 ;
        RECT 91.390 164.620 91.680 164.665 ;
        RECT 93.280 164.620 93.570 164.665 ;
        RECT 88.270 164.480 93.570 164.620 ;
        RECT 68.375 164.420 68.695 164.480 ;
        RECT 71.135 164.420 71.455 164.480 ;
        RECT 88.270 164.435 88.560 164.480 ;
        RECT 91.390 164.435 91.680 164.480 ;
        RECT 93.280 164.435 93.570 164.480 ;
        RECT 26.055 164.280 26.375 164.340 ;
        RECT 22.465 164.140 26.375 164.280 ;
        RECT 26.055 164.080 26.375 164.140 ;
        RECT 28.815 164.280 29.135 164.340 ;
        RECT 36.650 164.280 36.940 164.325 ;
        RECT 28.815 164.140 36.940 164.280 ;
        RECT 28.815 164.080 29.135 164.140 ;
        RECT 36.650 164.095 36.940 164.140 ;
        RECT 46.755 164.080 47.075 164.340 ;
        RECT 59.175 164.280 59.495 164.340 ;
        RECT 60.110 164.280 60.400 164.325 ;
        RECT 59.175 164.140 60.400 164.280 ;
        RECT 59.175 164.080 59.495 164.140 ;
        RECT 60.110 164.095 60.400 164.140 ;
        RECT 63.775 164.280 64.095 164.340 ;
        RECT 66.090 164.280 66.380 164.325 ;
        RECT 63.775 164.140 66.380 164.280 ;
        RECT 63.775 164.080 64.095 164.140 ;
        RECT 66.090 164.095 66.380 164.140 ;
        RECT 72.070 164.280 72.360 164.325 ;
        RECT 72.975 164.280 73.295 164.340 ;
        RECT 72.070 164.140 73.295 164.280 ;
        RECT 72.070 164.095 72.360 164.140 ;
        RECT 72.975 164.080 73.295 164.140 ;
        RECT 79.875 164.280 80.195 164.340 ;
        RECT 84.030 164.280 84.320 164.325 ;
        RECT 79.875 164.140 84.320 164.280 ;
        RECT 79.875 164.080 80.195 164.140 ;
        RECT 84.030 164.095 84.320 164.140 ;
        RECT 94.595 164.080 94.915 164.340 ;
        RECT 102.875 164.280 103.195 164.340 ;
        RECT 104.730 164.280 105.020 164.325 ;
        RECT 102.875 164.140 105.020 164.280 ;
        RECT 102.875 164.080 103.195 164.140 ;
        RECT 104.730 164.095 105.020 164.140 ;
        RECT 107.490 164.280 107.780 164.325 ;
        RECT 108.395 164.280 108.715 164.340 ;
        RECT 107.490 164.140 108.715 164.280 ;
        RECT 107.490 164.095 107.780 164.140 ;
        RECT 108.395 164.080 108.715 164.140 ;
        RECT 18.165 163.460 112.465 163.940 ;
        RECT 26.055 163.260 26.375 163.320 ;
        RECT 35.270 163.260 35.560 163.305 ;
        RECT 26.055 163.120 35.560 163.260 ;
        RECT 26.055 163.060 26.375 163.120 ;
        RECT 35.270 163.075 35.560 163.120 ;
        RECT 52.275 163.260 52.595 163.320 ;
        RECT 71.150 163.260 71.440 163.305 ;
        RECT 75.735 163.260 76.055 163.320 ;
        RECT 52.275 163.120 58.945 163.260 ;
        RECT 52.275 163.060 52.595 163.120 ;
        RECT 21.930 162.920 22.220 162.965 ;
        RECT 27.435 162.920 27.755 162.980 ;
        RECT 21.930 162.780 27.755 162.920 ;
        RECT 21.930 162.735 22.220 162.780 ;
        RECT 27.435 162.720 27.755 162.780 ;
        RECT 28.470 162.920 28.760 162.965 ;
        RECT 31.590 162.920 31.880 162.965 ;
        RECT 33.480 162.920 33.770 162.965 ;
        RECT 28.470 162.780 33.770 162.920 ;
        RECT 28.470 162.735 28.760 162.780 ;
        RECT 31.590 162.735 31.880 162.780 ;
        RECT 33.480 162.735 33.770 162.780 ;
        RECT 35.715 162.920 36.035 162.980 ;
        RECT 39.855 162.920 40.175 162.980 ;
        RECT 35.715 162.780 40.175 162.920 ;
        RECT 35.715 162.720 36.035 162.780 ;
        RECT 39.855 162.720 40.175 162.780 ;
        RECT 51.785 162.920 52.075 162.965 ;
        RECT 54.565 162.920 54.855 162.965 ;
        RECT 56.425 162.920 56.715 162.965 ;
        RECT 51.785 162.780 56.715 162.920 ;
        RECT 51.785 162.735 52.075 162.780 ;
        RECT 54.565 162.735 54.855 162.780 ;
        RECT 56.425 162.735 56.715 162.780 ;
        RECT 57.810 162.735 58.100 162.965 ;
        RECT 32.970 162.580 33.260 162.625 ;
        RECT 35.255 162.580 35.575 162.640 ;
        RECT 32.970 162.440 35.575 162.580 ;
        RECT 32.970 162.395 33.260 162.440 ;
        RECT 35.255 162.380 35.575 162.440 ;
        RECT 36.635 162.580 36.955 162.640 ;
        RECT 38.015 162.580 38.335 162.640 ;
        RECT 36.635 162.440 38.335 162.580 ;
        RECT 39.945 162.580 40.085 162.720 ;
        RECT 39.945 162.440 41.925 162.580 ;
        RECT 36.635 162.380 36.955 162.440 ;
        RECT 38.015 162.380 38.335 162.440 ;
        RECT 21.470 162.055 21.760 162.285 ;
        RECT 21.545 161.900 21.685 162.055 ;
        RECT 23.295 162.040 23.615 162.300 ;
        RECT 23.755 162.240 24.075 162.300 ;
        RECT 25.135 162.240 25.455 162.300 ;
        RECT 23.755 162.100 25.455 162.240 ;
        RECT 23.755 162.040 24.075 162.100 ;
        RECT 25.135 162.040 25.455 162.100 ;
        RECT 23.845 161.900 23.985 162.040 ;
        RECT 27.390 161.945 27.680 162.260 ;
        RECT 28.470 162.240 28.760 162.285 ;
        RECT 32.050 162.240 32.340 162.285 ;
        RECT 33.885 162.240 34.175 162.285 ;
        RECT 28.470 162.100 34.175 162.240 ;
        RECT 28.470 162.055 28.760 162.100 ;
        RECT 32.050 162.055 32.340 162.100 ;
        RECT 33.885 162.055 34.175 162.100 ;
        RECT 34.350 162.055 34.640 162.285 ;
        RECT 21.545 161.760 23.985 161.900 ;
        RECT 27.090 161.900 27.680 161.945 ;
        RECT 27.895 161.900 28.215 161.960 ;
        RECT 30.330 161.900 30.980 161.945 ;
        RECT 27.090 161.760 30.980 161.900 ;
        RECT 27.090 161.715 27.380 161.760 ;
        RECT 27.895 161.700 28.215 161.760 ;
        RECT 30.330 161.715 30.980 161.760 ;
        RECT 31.575 161.900 31.895 161.960 ;
        RECT 34.425 161.900 34.565 162.055 ;
        RECT 37.095 162.040 37.415 162.300 ;
        RECT 40.315 162.040 40.635 162.300 ;
        RECT 41.785 162.285 41.925 162.440 ;
        RECT 43.535 162.380 43.855 162.640 ;
        RECT 44.010 162.580 44.300 162.625 ;
        RECT 44.455 162.580 44.775 162.640 ;
        RECT 44.010 162.440 44.775 162.580 ;
        RECT 44.010 162.395 44.300 162.440 ;
        RECT 44.455 162.380 44.775 162.440 ;
        RECT 44.915 162.580 45.235 162.640 ;
        RECT 56.890 162.580 57.180 162.625 ;
        RECT 57.335 162.580 57.655 162.640 ;
        RECT 44.915 162.440 46.525 162.580 ;
        RECT 44.915 162.380 45.235 162.440 ;
        RECT 41.250 162.240 41.540 162.285 ;
        RECT 40.865 162.100 41.540 162.240 ;
        RECT 40.865 161.900 41.005 162.100 ;
        RECT 41.250 162.055 41.540 162.100 ;
        RECT 41.710 162.055 42.000 162.285 ;
        RECT 42.170 162.240 42.460 162.285 ;
        RECT 42.615 162.240 42.935 162.300 ;
        RECT 42.170 162.100 42.935 162.240 ;
        RECT 42.170 162.055 42.460 162.100 ;
        RECT 31.575 161.760 34.565 161.900 ;
        RECT 37.645 161.760 41.005 161.900 ;
        RECT 31.575 161.700 31.895 161.760 ;
        RECT 25.595 161.360 25.915 161.620 ;
        RECT 32.495 161.560 32.815 161.620 ;
        RECT 34.335 161.560 34.655 161.620 ;
        RECT 37.645 161.605 37.785 161.760 ;
        RECT 37.570 161.560 37.860 161.605 ;
        RECT 32.495 161.420 37.860 161.560 ;
        RECT 32.495 161.360 32.815 161.420 ;
        RECT 34.335 161.360 34.655 161.420 ;
        RECT 37.570 161.375 37.860 161.420 ;
        RECT 38.475 161.560 38.795 161.620 ;
        RECT 42.245 161.560 42.385 162.055 ;
        RECT 42.615 162.040 42.935 162.100 ;
        RECT 45.375 162.040 45.695 162.300 ;
        RECT 45.835 162.040 46.155 162.300 ;
        RECT 46.385 162.285 46.525 162.440 ;
        RECT 56.890 162.440 57.655 162.580 ;
        RECT 56.890 162.395 57.180 162.440 ;
        RECT 57.335 162.380 57.655 162.440 ;
        RECT 46.310 162.055 46.600 162.285 ;
        RECT 47.215 162.040 47.535 162.300 ;
        RECT 51.785 162.240 52.075 162.285 ;
        RECT 55.050 162.240 55.340 162.285 ;
        RECT 57.885 162.240 58.025 162.735 ;
        RECT 58.805 162.285 58.945 163.120 ;
        RECT 71.150 163.120 76.055 163.260 ;
        RECT 71.150 163.075 71.440 163.120 ;
        RECT 75.735 163.060 76.055 163.120 ;
        RECT 80.335 163.260 80.655 163.320 ;
        RECT 87.250 163.260 87.540 163.305 ;
        RECT 80.335 163.120 87.540 163.260 ;
        RECT 80.335 163.060 80.655 163.120 ;
        RECT 87.250 163.075 87.540 163.120 ;
        RECT 91.850 163.260 92.140 163.305 ;
        RECT 92.755 163.260 93.075 163.320 ;
        RECT 91.850 163.120 93.075 163.260 ;
        RECT 91.850 163.075 92.140 163.120 ;
        RECT 92.755 163.060 93.075 163.120 ;
        RECT 93.215 163.260 93.535 163.320 ;
        RECT 95.530 163.260 95.820 163.305 ;
        RECT 106.555 163.260 106.875 163.320 ;
        RECT 93.215 163.120 95.820 163.260 ;
        RECT 93.215 163.060 93.535 163.120 ;
        RECT 95.530 163.075 95.820 163.120 ;
        RECT 101.355 163.120 106.875 163.260 ;
        RECT 65.170 162.920 65.460 162.965 ;
        RECT 68.375 162.920 68.695 162.980 ;
        RECT 63.405 162.780 68.695 162.920 ;
        RECT 62.395 162.380 62.715 162.640 ;
        RECT 63.405 162.625 63.545 162.780 ;
        RECT 65.170 162.735 65.460 162.780 ;
        RECT 68.375 162.720 68.695 162.780 ;
        RECT 70.215 162.920 70.535 162.980 ;
        RECT 78.510 162.920 78.800 162.965 ;
        RECT 80.795 162.920 81.115 162.980 ;
        RECT 70.215 162.780 81.115 162.920 ;
        RECT 70.215 162.720 70.535 162.780 ;
        RECT 78.510 162.735 78.800 162.780 ;
        RECT 80.795 162.720 81.115 162.780 ;
        RECT 85.870 162.735 86.160 162.965 ;
        RECT 100.590 162.920 100.880 162.965 ;
        RECT 101.355 162.920 101.495 163.120 ;
        RECT 106.555 163.060 106.875 163.120 ;
        RECT 100.590 162.780 101.495 162.920 ;
        RECT 103.910 162.920 104.200 162.965 ;
        RECT 107.030 162.920 107.320 162.965 ;
        RECT 108.920 162.920 109.210 162.965 ;
        RECT 103.910 162.780 109.210 162.920 ;
        RECT 100.590 162.735 100.880 162.780 ;
        RECT 103.910 162.735 104.200 162.780 ;
        RECT 107.030 162.735 107.320 162.780 ;
        RECT 108.920 162.735 109.210 162.780 ;
        RECT 63.330 162.395 63.620 162.625 ;
        RECT 63.790 162.580 64.080 162.625 ;
        RECT 67.915 162.580 68.235 162.640 ;
        RECT 63.790 162.440 68.235 162.580 ;
        RECT 63.790 162.395 64.080 162.440 ;
        RECT 67.915 162.380 68.235 162.440 ;
        RECT 83.110 162.395 83.400 162.625 ;
        RECT 51.785 162.100 54.320 162.240 ;
        RECT 51.785 162.055 52.075 162.100 ;
        RECT 46.755 161.900 47.075 161.960 ;
        RECT 54.105 161.945 54.320 162.100 ;
        RECT 55.050 162.100 58.025 162.240 ;
        RECT 55.050 162.055 55.340 162.100 ;
        RECT 58.730 162.055 59.020 162.285 ;
        RECT 59.190 162.055 59.480 162.285 ;
        RECT 49.925 161.900 50.215 161.945 ;
        RECT 53.185 161.900 53.475 161.945 ;
        RECT 46.755 161.760 53.475 161.900 ;
        RECT 46.755 161.700 47.075 161.760 ;
        RECT 49.925 161.715 50.215 161.760 ;
        RECT 53.185 161.715 53.475 161.760 ;
        RECT 54.105 161.900 54.395 161.945 ;
        RECT 55.965 161.900 56.255 161.945 ;
        RECT 54.105 161.760 56.255 161.900 ;
        RECT 54.105 161.715 54.395 161.760 ;
        RECT 55.965 161.715 56.255 161.760 ;
        RECT 58.255 161.900 58.575 161.960 ;
        RECT 59.265 161.900 59.405 162.055 ;
        RECT 61.490 161.900 61.780 161.945 ;
        RECT 58.255 161.760 61.780 161.900 ;
        RECT 62.485 161.900 62.625 162.380 ;
        RECT 62.870 162.240 63.160 162.285 ;
        RECT 67.455 162.240 67.775 162.300 ;
        RECT 62.870 162.100 67.775 162.240 ;
        RECT 62.870 162.055 63.160 162.100 ;
        RECT 67.455 162.040 67.775 162.100 ;
        RECT 68.850 162.240 69.140 162.285 ;
        RECT 69.295 162.240 69.615 162.300 ;
        RECT 68.850 162.100 69.615 162.240 ;
        RECT 68.850 162.055 69.140 162.100 ;
        RECT 69.295 162.040 69.615 162.100 ;
        RECT 72.055 162.040 72.375 162.300 ;
        RECT 83.185 162.240 83.325 162.395 ;
        RECT 83.555 162.380 83.875 162.640 ;
        RECT 85.945 162.580 86.085 162.735 ;
        RECT 85.945 162.440 91.145 162.580 ;
        RECT 84.935 162.240 85.255 162.300 ;
        RECT 83.185 162.100 85.255 162.240 ;
        RECT 84.935 162.040 85.255 162.100 ;
        RECT 87.695 162.240 88.015 162.300 ;
        RECT 87.695 162.100 89.765 162.240 ;
        RECT 87.695 162.040 88.015 162.100 ;
        RECT 65.170 161.900 65.460 161.945 ;
        RECT 66.995 161.900 67.315 161.960 ;
        RECT 62.485 161.760 67.315 161.900 ;
        RECT 58.255 161.700 58.575 161.760 ;
        RECT 61.490 161.715 61.780 161.760 ;
        RECT 65.170 161.715 65.460 161.760 ;
        RECT 66.995 161.700 67.315 161.760 ;
        RECT 69.755 161.700 70.075 161.960 ;
        RECT 71.595 161.900 71.915 161.960 ;
        RECT 89.625 161.900 89.765 162.100 ;
        RECT 89.995 162.040 90.315 162.300 ;
        RECT 91.005 162.285 91.145 162.440 ;
        RECT 97.815 162.380 98.135 162.640 ;
        RECT 108.395 162.380 108.715 162.640 ;
        RECT 109.775 162.380 110.095 162.640 ;
        RECT 90.930 162.055 91.220 162.285 ;
        RECT 91.375 162.040 91.695 162.300 ;
        RECT 94.595 162.240 94.915 162.300 ;
        RECT 96.450 162.240 96.740 162.285 ;
        RECT 94.595 162.100 96.740 162.240 ;
        RECT 94.595 162.040 94.915 162.100 ;
        RECT 96.450 162.055 96.740 162.100 ;
        RECT 98.275 162.240 98.595 162.300 ;
        RECT 102.875 162.260 103.195 162.300 ;
        RECT 98.275 162.100 98.965 162.240 ;
        RECT 98.275 162.040 98.595 162.100 ;
        RECT 91.465 161.900 91.605 162.040 ;
        RECT 98.825 161.945 98.965 162.100 ;
        RECT 102.830 162.040 103.195 162.260 ;
        RECT 103.910 162.240 104.200 162.285 ;
        RECT 107.490 162.240 107.780 162.285 ;
        RECT 109.325 162.240 109.615 162.285 ;
        RECT 103.910 162.100 109.615 162.240 ;
        RECT 103.910 162.055 104.200 162.100 ;
        RECT 107.490 162.055 107.780 162.100 ;
        RECT 109.325 162.055 109.615 162.100 ;
        RECT 102.830 161.945 103.120 162.040 ;
        RECT 71.595 161.760 87.925 161.900 ;
        RECT 89.625 161.760 91.605 161.900 ;
        RECT 71.595 161.700 71.915 161.760 ;
        RECT 87.785 161.620 87.925 161.760 ;
        RECT 98.750 161.715 99.040 161.945 ;
        RECT 102.530 161.900 103.120 161.945 ;
        RECT 105.770 161.900 106.420 161.945 ;
        RECT 102.530 161.760 106.420 161.900 ;
        RECT 102.530 161.715 102.820 161.760 ;
        RECT 105.770 161.715 106.420 161.760 ;
        RECT 38.475 161.420 42.385 161.560 ;
        RECT 47.920 161.560 48.210 161.605 ;
        RECT 48.595 161.560 48.915 161.620 ;
        RECT 47.920 161.420 48.915 161.560 ;
        RECT 38.475 161.360 38.795 161.420 ;
        RECT 47.920 161.375 48.210 161.420 ;
        RECT 48.595 161.360 48.915 161.420 ;
        RECT 50.895 161.560 51.215 161.620 ;
        RECT 52.735 161.560 53.055 161.620 ;
        RECT 50.895 161.420 53.055 161.560 ;
        RECT 50.895 161.360 51.215 161.420 ;
        RECT 52.735 161.360 53.055 161.420 ;
        RECT 60.110 161.560 60.400 161.605 ;
        RECT 61.015 161.560 61.335 161.620 ;
        RECT 63.315 161.560 63.635 161.620 ;
        RECT 60.110 161.420 63.635 161.560 ;
        RECT 60.110 161.375 60.400 161.420 ;
        RECT 61.015 161.360 61.335 161.420 ;
        RECT 63.315 161.360 63.635 161.420 ;
        RECT 84.015 161.360 84.335 161.620 ;
        RECT 87.695 161.360 88.015 161.620 ;
        RECT 97.815 161.560 98.135 161.620 ;
        RECT 98.290 161.560 98.580 161.605 ;
        RECT 101.050 161.560 101.340 161.605 ;
        RECT 97.815 161.420 101.340 161.560 ;
        RECT 97.815 161.360 98.135 161.420 ;
        RECT 98.290 161.375 98.580 161.420 ;
        RECT 101.050 161.375 101.340 161.420 ;
        RECT 17.370 160.740 112.465 161.220 ;
        RECT 21.455 160.340 21.775 160.600 ;
        RECT 25.610 160.540 25.900 160.585 ;
        RECT 22.925 160.400 25.900 160.540 ;
        RECT 20.550 159.860 20.840 159.905 ;
        RECT 22.925 159.860 23.065 160.400 ;
        RECT 25.610 160.355 25.900 160.400 ;
        RECT 27.910 160.540 28.200 160.585 ;
        RECT 37.555 160.540 37.875 160.600 ;
        RECT 49.990 160.540 50.280 160.585 ;
        RECT 27.910 160.400 40.545 160.540 ;
        RECT 27.910 160.355 28.200 160.400 ;
        RECT 37.555 160.340 37.875 160.400 ;
        RECT 23.755 160.000 24.075 160.260 ;
        RECT 31.115 160.200 31.435 160.260 ;
        RECT 33.530 160.200 33.820 160.245 ;
        RECT 36.770 160.200 37.420 160.245 ;
        RECT 31.115 160.060 37.420 160.200 ;
        RECT 31.115 160.000 31.435 160.060 ;
        RECT 33.530 160.015 34.120 160.060 ;
        RECT 36.770 160.015 37.420 160.060 ;
        RECT 39.410 160.200 39.700 160.245 ;
        RECT 39.855 160.200 40.175 160.260 ;
        RECT 39.410 160.060 40.175 160.200 ;
        RECT 40.405 160.200 40.545 160.400 ;
        RECT 43.165 160.400 50.280 160.540 ;
        RECT 43.165 160.200 43.305 160.400 ;
        RECT 49.990 160.355 50.280 160.400 ;
        RECT 51.830 160.540 52.120 160.585 ;
        RECT 52.275 160.540 52.595 160.600 ;
        RECT 51.830 160.400 52.595 160.540 ;
        RECT 51.830 160.355 52.120 160.400 ;
        RECT 52.275 160.340 52.595 160.400 ;
        RECT 54.575 160.540 54.895 160.600 ;
        RECT 58.730 160.540 59.020 160.585 ;
        RECT 71.595 160.540 71.915 160.600 ;
        RECT 54.575 160.400 71.915 160.540 ;
        RECT 54.575 160.340 54.895 160.400 ;
        RECT 58.730 160.355 59.020 160.400 ;
        RECT 71.595 160.340 71.915 160.400 ;
        RECT 72.515 160.540 72.835 160.600 ;
        RECT 75.060 160.540 75.350 160.585 ;
        RECT 84.015 160.540 84.335 160.600 ;
        RECT 72.515 160.400 84.335 160.540 ;
        RECT 72.515 160.340 72.835 160.400 ;
        RECT 75.060 160.355 75.350 160.400 ;
        RECT 84.015 160.340 84.335 160.400 ;
        RECT 84.490 160.355 84.780 160.585 ;
        RECT 87.695 160.540 88.015 160.600 ;
        RECT 92.755 160.540 93.075 160.600 ;
        RECT 87.695 160.400 101.265 160.540 ;
        RECT 80.335 160.245 80.655 160.260 ;
        RECT 40.405 160.060 43.305 160.200 ;
        RECT 56.890 160.200 57.180 160.245 ;
        RECT 65.630 160.200 65.920 160.245 ;
        RECT 71.150 160.200 71.440 160.245 ;
        RECT 56.890 160.060 71.440 160.200 ;
        RECT 39.410 160.015 39.700 160.060 ;
        RECT 20.550 159.720 23.065 159.860 ;
        RECT 20.550 159.675 20.840 159.720 ;
        RECT 25.150 159.675 25.440 159.905 ;
        RECT 25.595 159.860 25.915 159.920 ;
        RECT 27.450 159.860 27.740 159.905 ;
        RECT 32.035 159.860 32.355 159.920 ;
        RECT 25.595 159.720 32.355 159.860 ;
        RECT 25.225 159.180 25.365 159.675 ;
        RECT 25.595 159.660 25.915 159.720 ;
        RECT 27.450 159.675 27.740 159.720 ;
        RECT 32.035 159.660 32.355 159.720 ;
        RECT 33.830 159.700 34.120 160.015 ;
        RECT 39.855 160.000 40.175 160.060 ;
        RECT 56.890 160.015 57.180 160.060 ;
        RECT 65.630 160.015 65.920 160.060 ;
        RECT 71.150 160.015 71.440 160.060 ;
        RECT 77.065 160.200 77.355 160.245 ;
        RECT 80.325 160.200 80.655 160.245 ;
        RECT 77.065 160.060 80.655 160.200 ;
        RECT 77.065 160.015 77.355 160.060 ;
        RECT 80.325 160.015 80.655 160.060 ;
        RECT 80.335 160.000 80.655 160.015 ;
        RECT 81.245 160.200 81.535 160.245 ;
        RECT 83.105 160.200 83.395 160.245 ;
        RECT 81.245 160.060 83.395 160.200 ;
        RECT 81.245 160.015 81.535 160.060 ;
        RECT 83.105 160.015 83.395 160.060 ;
        RECT 34.910 159.860 35.200 159.905 ;
        RECT 38.490 159.860 38.780 159.905 ;
        RECT 40.325 159.860 40.615 159.905 ;
        RECT 34.910 159.720 40.615 159.860 ;
        RECT 34.910 159.675 35.200 159.720 ;
        RECT 38.490 159.675 38.780 159.720 ;
        RECT 40.325 159.675 40.615 159.720 ;
        RECT 43.075 159.660 43.395 159.920 ;
        RECT 45.375 159.660 45.695 159.920 ;
        RECT 45.835 159.660 46.155 159.920 ;
        RECT 46.295 159.660 46.615 159.920 ;
        RECT 47.215 159.660 47.535 159.920 ;
        RECT 48.595 159.860 48.915 159.920 ;
        RECT 49.530 159.860 49.820 159.905 ;
        RECT 48.595 159.720 49.820 159.860 ;
        RECT 48.595 159.660 48.915 159.720 ;
        RECT 49.530 159.675 49.820 159.720 ;
        RECT 52.275 159.660 52.595 159.920 ;
        RECT 52.735 159.860 53.055 159.920 ;
        RECT 53.670 159.860 53.960 159.905 ;
        RECT 55.035 159.860 55.355 159.920 ;
        RECT 52.735 159.720 55.355 159.860 ;
        RECT 52.735 159.660 53.055 159.720 ;
        RECT 53.670 159.675 53.960 159.720 ;
        RECT 55.035 159.660 55.355 159.720 ;
        RECT 59.650 159.860 59.940 159.905 ;
        RECT 60.555 159.860 60.875 159.920 ;
        RECT 61.475 159.860 61.795 159.920 ;
        RECT 59.650 159.720 61.795 159.860 ;
        RECT 59.650 159.675 59.940 159.720 ;
        RECT 60.555 159.660 60.875 159.720 ;
        RECT 61.475 159.660 61.795 159.720 ;
        RECT 61.935 159.660 62.255 159.920 ;
        RECT 63.315 159.660 63.635 159.920 ;
        RECT 64.695 159.660 65.015 159.920 ;
        RECT 65.170 159.860 65.460 159.905 ;
        RECT 66.535 159.860 66.855 159.920 ;
        RECT 65.170 159.720 66.855 159.860 ;
        RECT 65.170 159.675 65.460 159.720 ;
        RECT 66.535 159.660 66.855 159.720 ;
        RECT 66.995 159.660 67.315 159.920 ;
        RECT 67.455 159.660 67.775 159.920 ;
        RECT 67.915 159.660 68.235 159.920 ;
        RECT 68.375 159.660 68.695 159.920 ;
        RECT 78.925 159.860 79.215 159.905 ;
        RECT 81.245 159.860 81.460 160.015 ;
        RECT 78.925 159.720 81.460 159.860 ;
        RECT 82.190 159.860 82.480 159.905 ;
        RECT 84.565 159.860 84.705 160.355 ;
        RECT 87.695 160.340 88.015 160.400 ;
        RECT 92.755 160.340 93.075 160.400 ;
        RECT 84.935 160.200 85.255 160.260 ;
        RECT 91.390 160.200 91.680 160.245 ;
        RECT 93.215 160.200 93.535 160.260 ;
        RECT 84.935 160.060 90.685 160.200 ;
        RECT 84.935 160.000 85.255 160.060 ;
        RECT 82.190 159.720 84.705 159.860 ;
        RECT 78.925 159.675 79.215 159.720 ;
        RECT 82.190 159.675 82.480 159.720 ;
        RECT 85.395 159.660 85.715 159.920 ;
        RECT 85.855 159.660 86.175 159.920 ;
        RECT 86.315 159.860 86.635 159.920 ;
        RECT 86.790 159.860 87.080 159.905 ;
        RECT 86.315 159.720 87.080 159.860 ;
        RECT 86.315 159.660 86.635 159.720 ;
        RECT 86.790 159.675 87.080 159.720 ;
        RECT 87.235 159.660 87.555 159.920 ;
        RECT 87.710 159.675 88.000 159.905 ;
        RECT 90.545 159.860 90.685 160.060 ;
        RECT 91.390 160.060 93.535 160.200 ;
        RECT 91.390 160.015 91.680 160.060 ;
        RECT 93.215 160.000 93.535 160.060 ;
        RECT 97.445 159.905 97.585 160.400 ;
        RECT 98.275 160.200 98.595 160.260 ;
        RECT 98.275 160.060 100.805 160.200 ;
        RECT 98.275 160.000 98.595 160.060 ;
        RECT 93.690 159.860 93.980 159.905 ;
        RECT 90.545 159.720 91.605 159.860 ;
        RECT 28.830 159.520 29.120 159.565 ;
        RECT 32.955 159.520 33.275 159.580 ;
        RECT 36.635 159.520 36.955 159.580 ;
        RECT 28.830 159.380 36.955 159.520 ;
        RECT 28.830 159.335 29.120 159.380 ;
        RECT 32.955 159.320 33.275 159.380 ;
        RECT 36.635 159.320 36.955 159.380 ;
        RECT 40.775 159.320 41.095 159.580 ;
        RECT 41.695 159.520 42.015 159.580 ;
        RECT 45.925 159.520 46.065 159.660 ;
        RECT 41.695 159.380 46.065 159.520 ;
        RECT 41.695 159.320 42.015 159.380 ;
        RECT 33.875 159.180 34.195 159.240 ;
        RECT 25.225 159.040 34.195 159.180 ;
        RECT 33.875 158.980 34.195 159.040 ;
        RECT 34.910 159.180 35.200 159.225 ;
        RECT 38.030 159.180 38.320 159.225 ;
        RECT 39.920 159.180 40.210 159.225 ;
        RECT 34.910 159.040 40.210 159.180 ;
        RECT 45.925 159.180 46.065 159.380 ;
        RECT 49.055 159.520 49.375 159.580 ;
        RECT 55.510 159.520 55.800 159.565 ;
        RECT 80.795 159.520 81.115 159.580 ;
        RECT 84.030 159.520 84.320 159.565 ;
        RECT 84.475 159.520 84.795 159.580 ;
        RECT 87.785 159.520 87.925 159.675 ;
        RECT 90.545 159.565 90.685 159.720 ;
        RECT 49.055 159.380 55.800 159.520 ;
        RECT 49.055 159.320 49.375 159.380 ;
        RECT 55.510 159.335 55.800 159.380 ;
        RECT 60.645 159.380 65.385 159.520 ;
        RECT 54.575 159.180 54.895 159.240 ;
        RECT 60.645 159.225 60.785 159.380 ;
        RECT 65.245 159.240 65.385 159.380 ;
        RECT 80.795 159.380 84.795 159.520 ;
        RECT 80.795 159.320 81.115 159.380 ;
        RECT 84.030 159.335 84.320 159.380 ;
        RECT 84.475 159.320 84.795 159.380 ;
        RECT 85.945 159.380 87.925 159.520 ;
        RECT 60.570 159.180 60.860 159.225 ;
        RECT 45.925 159.040 54.895 159.180 ;
        RECT 34.910 158.995 35.200 159.040 ;
        RECT 38.030 158.995 38.320 159.040 ;
        RECT 39.920 158.995 40.210 159.040 ;
        RECT 54.575 158.980 54.895 159.040 ;
        RECT 55.125 159.040 60.860 159.180 ;
        RECT 28.815 158.840 29.135 158.900 ;
        RECT 32.050 158.840 32.340 158.885 ;
        RECT 28.815 158.700 32.340 158.840 ;
        RECT 28.815 158.640 29.135 158.700 ;
        RECT 32.050 158.655 32.340 158.700 ;
        RECT 36.635 158.840 36.955 158.900 ;
        RECT 41.710 158.840 42.000 158.885 ;
        RECT 36.635 158.700 42.000 158.840 ;
        RECT 36.635 158.640 36.955 158.700 ;
        RECT 41.710 158.655 42.000 158.700 ;
        RECT 44.010 158.840 44.300 158.885 ;
        RECT 44.915 158.840 45.235 158.900 ;
        RECT 44.010 158.700 45.235 158.840 ;
        RECT 44.010 158.655 44.300 158.700 ;
        RECT 44.915 158.640 45.235 158.700 ;
        RECT 47.675 158.840 47.995 158.900 ;
        RECT 55.125 158.840 55.265 159.040 ;
        RECT 60.570 158.995 60.860 159.040 ;
        RECT 62.855 158.980 63.175 159.240 ;
        RECT 63.315 159.180 63.635 159.240 ;
        RECT 63.790 159.180 64.080 159.225 ;
        RECT 63.315 159.040 64.080 159.180 ;
        RECT 63.315 158.980 63.635 159.040 ;
        RECT 63.790 158.995 64.080 159.040 ;
        RECT 65.155 158.980 65.475 159.240 ;
        RECT 65.615 159.180 65.935 159.240 ;
        RECT 66.090 159.180 66.380 159.225 ;
        RECT 65.615 159.040 66.380 159.180 ;
        RECT 65.615 158.980 65.935 159.040 ;
        RECT 66.090 158.995 66.380 159.040 ;
        RECT 72.530 159.180 72.820 159.225 ;
        RECT 75.275 159.180 75.595 159.240 ;
        RECT 72.530 159.040 75.595 159.180 ;
        RECT 72.530 158.995 72.820 159.040 ;
        RECT 75.275 158.980 75.595 159.040 ;
        RECT 78.925 159.180 79.215 159.225 ;
        RECT 81.705 159.180 81.995 159.225 ;
        RECT 83.565 159.180 83.855 159.225 ;
        RECT 78.925 159.040 83.855 159.180 ;
        RECT 78.925 158.995 79.215 159.040 ;
        RECT 81.705 158.995 81.995 159.040 ;
        RECT 83.565 158.995 83.855 159.040 ;
        RECT 47.675 158.700 55.265 158.840 ;
        RECT 56.875 158.840 57.195 158.900 ;
        RECT 85.945 158.840 86.085 159.380 ;
        RECT 90.470 159.335 90.760 159.565 ;
        RECT 90.930 159.335 91.220 159.565 ;
        RECT 89.535 159.180 89.855 159.240 ;
        RECT 91.005 159.180 91.145 159.335 ;
        RECT 89.535 159.040 91.145 159.180 ;
        RECT 89.535 158.980 89.855 159.040 ;
        RECT 87.235 158.840 87.555 158.900 ;
        RECT 56.875 158.700 87.555 158.840 ;
        RECT 47.675 158.640 47.995 158.700 ;
        RECT 56.875 158.640 57.195 158.700 ;
        RECT 87.235 158.640 87.555 158.700 ;
        RECT 87.695 158.840 88.015 158.900 ;
        RECT 89.090 158.840 89.380 158.885 ;
        RECT 87.695 158.700 89.380 158.840 ;
        RECT 91.465 158.840 91.605 159.720 ;
        RECT 93.305 159.720 93.980 159.860 ;
        RECT 93.305 159.225 93.445 159.720 ;
        RECT 93.690 159.675 93.980 159.720 ;
        RECT 96.910 159.675 97.200 159.905 ;
        RECT 97.370 159.675 97.660 159.905 ;
        RECT 93.230 158.995 93.520 159.225 ;
        RECT 96.985 159.180 97.125 159.675 ;
        RECT 97.815 159.660 98.135 159.920 ;
        RECT 98.735 159.860 99.055 159.920 ;
        RECT 100.665 159.905 100.805 160.060 ;
        RECT 101.125 159.905 101.265 160.400 ;
        RECT 99.670 159.860 99.960 159.905 ;
        RECT 98.735 159.720 99.960 159.860 ;
        RECT 98.735 159.660 99.055 159.720 ;
        RECT 99.670 159.675 99.960 159.720 ;
        RECT 100.590 159.675 100.880 159.905 ;
        RECT 101.050 159.675 101.340 159.905 ;
        RECT 101.510 159.860 101.800 159.905 ;
        RECT 101.955 159.860 102.275 159.920 ;
        RECT 101.510 159.720 102.275 159.860 ;
        RECT 101.510 159.675 101.800 159.720 ;
        RECT 101.585 159.180 101.725 159.675 ;
        RECT 101.955 159.660 102.275 159.720 ;
        RECT 104.255 159.660 104.575 159.920 ;
        RECT 107.950 159.860 108.240 159.905 ;
        RECT 111.155 159.860 111.475 159.920 ;
        RECT 107.950 159.720 111.475 159.860 ;
        RECT 107.950 159.675 108.240 159.720 ;
        RECT 111.155 159.660 111.475 159.720 ;
        RECT 93.765 159.040 96.205 159.180 ;
        RECT 96.985 159.040 101.725 159.180 ;
        RECT 105.635 159.180 105.955 159.240 ;
        RECT 107.030 159.180 107.320 159.225 ;
        RECT 105.635 159.040 107.320 159.180 ;
        RECT 93.765 158.840 93.905 159.040 ;
        RECT 91.465 158.700 93.905 158.840 ;
        RECT 87.695 158.640 88.015 158.700 ;
        RECT 89.090 158.655 89.380 158.700 ;
        RECT 94.595 158.640 94.915 158.900 ;
        RECT 95.055 158.840 95.375 158.900 ;
        RECT 95.530 158.840 95.820 158.885 ;
        RECT 95.055 158.700 95.820 158.840 ;
        RECT 96.065 158.840 96.205 159.040 ;
        RECT 105.635 158.980 105.955 159.040 ;
        RECT 107.030 158.995 107.320 159.040 ;
        RECT 97.355 158.840 97.675 158.900 ;
        RECT 96.065 158.700 97.675 158.840 ;
        RECT 95.055 158.640 95.375 158.700 ;
        RECT 95.530 158.655 95.820 158.700 ;
        RECT 97.355 158.640 97.675 158.700 ;
        RECT 102.875 158.640 103.195 158.900 ;
        RECT 104.715 158.640 105.035 158.900 ;
        RECT 18.165 158.020 112.465 158.500 ;
        RECT 27.895 157.820 28.215 157.880 ;
        RECT 29.750 157.820 30.040 157.865 ;
        RECT 27.895 157.680 30.040 157.820 ;
        RECT 27.895 157.620 28.215 157.680 ;
        RECT 29.750 157.635 30.040 157.680 ;
        RECT 34.350 157.820 34.640 157.865 ;
        RECT 36.175 157.820 36.495 157.880 ;
        RECT 52.275 157.820 52.595 157.880 ;
        RECT 34.350 157.680 36.495 157.820 ;
        RECT 34.350 157.635 34.640 157.680 ;
        RECT 36.175 157.620 36.495 157.680 ;
        RECT 42.705 157.680 52.595 157.820 ;
        RECT 22.490 157.480 22.780 157.525 ;
        RECT 25.610 157.480 25.900 157.525 ;
        RECT 27.500 157.480 27.790 157.525 ;
        RECT 22.490 157.340 27.790 157.480 ;
        RECT 22.490 157.295 22.780 157.340 ;
        RECT 25.610 157.295 25.900 157.340 ;
        RECT 27.500 157.295 27.790 157.340 ;
        RECT 33.875 157.480 34.195 157.540 ;
        RECT 40.315 157.480 40.635 157.540 ;
        RECT 42.705 157.480 42.845 157.680 ;
        RECT 52.275 157.620 52.595 157.680 ;
        RECT 66.995 157.820 67.315 157.880 ;
        RECT 85.395 157.820 85.715 157.880 ;
        RECT 66.995 157.680 70.905 157.820 ;
        RECT 66.995 157.620 67.315 157.680 ;
        RECT 33.875 157.340 42.845 157.480 ;
        RECT 43.075 157.480 43.395 157.540 ;
        RECT 67.930 157.480 68.220 157.525 ;
        RECT 69.755 157.480 70.075 157.540 ;
        RECT 70.765 157.525 70.905 157.680 ;
        RECT 79.045 157.680 85.715 157.820 ;
        RECT 43.075 157.340 70.075 157.480 ;
        RECT 33.875 157.280 34.195 157.340 ;
        RECT 40.315 157.280 40.635 157.340 ;
        RECT 43.075 157.280 43.395 157.340 ;
        RECT 67.930 157.295 68.220 157.340 ;
        RECT 69.755 157.280 70.075 157.340 ;
        RECT 70.690 157.295 70.980 157.525 ;
        RECT 74.830 157.480 75.120 157.525 ;
        RECT 79.045 157.480 79.185 157.680 ;
        RECT 85.395 157.620 85.715 157.680 ;
        RECT 95.975 157.820 96.295 157.880 ;
        RECT 98.735 157.820 99.055 157.880 ;
        RECT 95.975 157.680 99.055 157.820 ;
        RECT 95.975 157.620 96.295 157.680 ;
        RECT 98.735 157.620 99.055 157.680 ;
        RECT 74.830 157.340 79.185 157.480 ;
        RECT 79.385 157.480 79.675 157.525 ;
        RECT 82.165 157.480 82.455 157.525 ;
        RECT 84.025 157.480 84.315 157.525 ;
        RECT 79.385 157.340 84.315 157.480 ;
        RECT 74.830 157.295 75.120 157.340 ;
        RECT 79.385 157.295 79.675 157.340 ;
        RECT 82.165 157.295 82.455 157.340 ;
        RECT 84.025 157.295 84.315 157.340 ;
        RECT 84.950 157.295 85.240 157.525 ;
        RECT 90.885 157.480 91.175 157.525 ;
        RECT 93.665 157.480 93.955 157.525 ;
        RECT 95.525 157.480 95.815 157.525 ;
        RECT 90.885 157.340 95.815 157.480 ;
        RECT 90.885 157.295 91.175 157.340 ;
        RECT 93.665 157.295 93.955 157.340 ;
        RECT 95.525 157.295 95.815 157.340 ;
        RECT 105.145 157.480 105.435 157.525 ;
        RECT 107.925 157.480 108.215 157.525 ;
        RECT 109.785 157.480 110.075 157.525 ;
        RECT 105.145 157.340 110.075 157.480 ;
        RECT 105.145 157.295 105.435 157.340 ;
        RECT 107.925 157.295 108.215 157.340 ;
        RECT 109.785 157.295 110.075 157.340 ;
        RECT 20.535 157.140 20.855 157.200 ;
        RECT 23.755 157.140 24.075 157.200 ;
        RECT 31.590 157.140 31.880 157.185 ;
        RECT 32.955 157.140 33.275 157.200 ;
        RECT 48.595 157.140 48.915 157.200 ;
        RECT 20.535 157.000 30.425 157.140 ;
        RECT 20.535 156.940 20.855 157.000 ;
        RECT 23.755 156.940 24.075 157.000 ;
        RECT 30.285 156.845 30.425 157.000 ;
        RECT 31.590 157.000 33.275 157.140 ;
        RECT 31.590 156.955 31.880 157.000 ;
        RECT 32.955 156.940 33.275 157.000 ;
        RECT 36.725 157.000 39.625 157.140 ;
        RECT 21.410 156.505 21.700 156.820 ;
        RECT 22.490 156.800 22.780 156.845 ;
        RECT 26.070 156.800 26.360 156.845 ;
        RECT 27.905 156.800 28.195 156.845 ;
        RECT 22.490 156.660 28.195 156.800 ;
        RECT 22.490 156.615 22.780 156.660 ;
        RECT 26.070 156.615 26.360 156.660 ;
        RECT 27.905 156.615 28.195 156.660 ;
        RECT 28.370 156.615 28.660 156.845 ;
        RECT 30.210 156.615 30.500 156.845 ;
        RECT 21.110 156.460 21.700 156.505 ;
        RECT 23.295 156.460 23.615 156.520 ;
        RECT 24.350 156.460 25.000 156.505 ;
        RECT 21.110 156.320 25.000 156.460 ;
        RECT 21.110 156.275 21.400 156.320 ;
        RECT 23.295 156.260 23.615 156.320 ;
        RECT 24.350 156.275 25.000 156.320 ;
        RECT 26.975 156.260 27.295 156.520 ;
        RECT 28.445 156.460 28.585 156.615 ;
        RECT 32.495 156.600 32.815 156.860 ;
        RECT 36.725 156.845 36.865 157.000 ;
        RECT 39.485 156.860 39.625 157.000 ;
        RECT 41.325 157.000 48.915 157.140 ;
        RECT 36.650 156.615 36.940 156.845 ;
        RECT 37.555 156.600 37.875 156.860 ;
        RECT 38.030 156.615 38.320 156.845 ;
        RECT 31.575 156.460 31.895 156.520 ;
        RECT 28.445 156.320 31.895 156.460 ;
        RECT 31.575 156.260 31.895 156.320 ;
        RECT 35.715 156.460 36.035 156.520 ;
        RECT 38.105 156.460 38.245 156.615 ;
        RECT 38.475 156.600 38.795 156.860 ;
        RECT 39.395 156.800 39.715 156.860 ;
        RECT 41.325 156.845 41.465 157.000 ;
        RECT 48.595 156.940 48.915 157.000 ;
        RECT 61.475 157.140 61.795 157.200 ;
        RECT 63.315 157.140 63.635 157.200 ;
        RECT 61.475 157.000 63.635 157.140 ;
        RECT 61.475 156.940 61.795 157.000 ;
        RECT 63.315 156.940 63.635 157.000 ;
        RECT 64.695 157.140 65.015 157.200 ;
        RECT 68.375 157.140 68.695 157.200 ;
        RECT 64.695 157.000 68.695 157.140 ;
        RECT 64.695 156.940 65.015 157.000 ;
        RECT 68.375 156.940 68.695 157.000 ;
        RECT 72.070 156.955 72.360 157.185 ;
        RECT 40.330 156.800 40.620 156.845 ;
        RECT 39.395 156.660 40.620 156.800 ;
        RECT 39.395 156.600 39.715 156.660 ;
        RECT 40.330 156.615 40.620 156.660 ;
        RECT 41.250 156.615 41.540 156.845 ;
        RECT 41.695 156.600 42.015 156.860 ;
        RECT 42.170 156.800 42.460 156.845 ;
        RECT 45.375 156.800 45.695 156.860 ;
        RECT 49.515 156.800 49.835 156.860 ;
        RECT 42.170 156.660 49.835 156.800 ;
        RECT 42.170 156.615 42.460 156.660 ;
        RECT 45.375 156.600 45.695 156.660 ;
        RECT 49.515 156.600 49.835 156.660 ;
        RECT 52.735 156.600 53.055 156.860 ;
        RECT 55.970 156.800 56.260 156.845 ;
        RECT 57.335 156.800 57.655 156.860 ;
        RECT 55.970 156.660 57.655 156.800 ;
        RECT 55.970 156.615 56.260 156.660 ;
        RECT 35.715 156.320 38.245 156.460 ;
        RECT 35.715 156.260 36.035 156.320 ;
        RECT 19.630 156.120 19.920 156.165 ;
        RECT 26.515 156.120 26.835 156.180 ;
        RECT 19.630 155.980 26.835 156.120 ;
        RECT 19.630 155.935 19.920 155.980 ;
        RECT 26.515 155.920 26.835 155.980 ;
        RECT 32.035 155.920 32.355 156.180 ;
        RECT 38.105 156.120 38.245 156.320 ;
        RECT 39.870 156.460 40.160 156.505 ;
        RECT 44.915 156.460 45.235 156.520 ;
        RECT 56.045 156.460 56.185 156.615 ;
        RECT 57.335 156.600 57.655 156.660 ;
        RECT 57.810 156.800 58.100 156.845 ;
        RECT 58.255 156.800 58.575 156.860 ;
        RECT 57.810 156.660 58.575 156.800 ;
        RECT 57.810 156.615 58.100 156.660 ;
        RECT 58.255 156.600 58.575 156.660 ;
        RECT 59.190 156.800 59.480 156.845 ;
        RECT 59.635 156.800 59.955 156.860 ;
        RECT 59.190 156.660 59.955 156.800 ;
        RECT 59.190 156.615 59.480 156.660 ;
        RECT 59.635 156.600 59.955 156.660 ;
        RECT 61.015 156.800 61.335 156.860 ;
        RECT 61.950 156.800 62.240 156.845 ;
        RECT 61.015 156.660 62.240 156.800 ;
        RECT 61.015 156.600 61.335 156.660 ;
        RECT 61.950 156.615 62.240 156.660 ;
        RECT 62.395 156.800 62.715 156.860 ;
        RECT 66.075 156.800 66.395 156.860 ;
        RECT 62.395 156.660 66.395 156.800 ;
        RECT 62.395 156.600 62.715 156.660 ;
        RECT 66.075 156.600 66.395 156.660 ;
        RECT 66.995 156.600 67.315 156.860 ;
        RECT 67.930 156.615 68.220 156.845 ;
        RECT 68.465 156.800 68.605 156.940 ;
        RECT 69.310 156.800 69.600 156.845 ;
        RECT 68.465 156.660 69.600 156.800 ;
        RECT 72.145 156.800 72.285 156.955 ;
        RECT 72.515 156.940 72.835 157.200 ;
        RECT 84.475 156.940 84.795 157.200 ;
        RECT 75.275 156.800 75.595 156.860 ;
        RECT 72.145 156.660 75.595 156.800 ;
        RECT 69.310 156.615 69.600 156.660 ;
        RECT 68.005 156.460 68.145 156.615 ;
        RECT 75.275 156.600 75.595 156.660 ;
        RECT 79.385 156.800 79.675 156.845 ;
        RECT 82.650 156.800 82.940 156.845 ;
        RECT 85.025 156.800 85.165 157.295 ;
        RECT 87.020 157.140 87.310 157.185 ;
        RECT 89.535 157.140 89.855 157.200 ;
        RECT 79.385 156.660 81.920 156.800 ;
        RECT 79.385 156.615 79.675 156.660 ;
        RECT 39.870 156.320 45.235 156.460 ;
        RECT 39.870 156.275 40.160 156.320 ;
        RECT 44.915 156.260 45.235 156.320 ;
        RECT 46.385 156.320 56.185 156.460 ;
        RECT 60.185 156.320 68.145 156.460 ;
        RECT 77.525 156.460 77.815 156.505 ;
        RECT 79.875 156.460 80.195 156.520 ;
        RECT 81.705 156.505 81.920 156.660 ;
        RECT 82.650 156.660 85.165 156.800 ;
        RECT 85.485 157.000 89.855 157.140 ;
        RECT 82.650 156.615 82.940 156.660 ;
        RECT 80.785 156.460 81.075 156.505 ;
        RECT 77.525 156.320 81.075 156.460 ;
        RECT 43.075 156.120 43.395 156.180 ;
        RECT 38.105 155.980 43.395 156.120 ;
        RECT 43.075 155.920 43.395 155.980 ;
        RECT 43.535 155.920 43.855 156.180 ;
        RECT 46.385 156.165 46.525 156.320 ;
        RECT 46.310 155.935 46.600 156.165 ;
        RECT 49.515 156.120 49.835 156.180 ;
        RECT 56.875 156.120 57.195 156.180 ;
        RECT 60.185 156.165 60.325 156.320 ;
        RECT 77.525 156.275 77.815 156.320 ;
        RECT 79.875 156.260 80.195 156.320 ;
        RECT 80.785 156.275 81.075 156.320 ;
        RECT 81.705 156.460 81.995 156.505 ;
        RECT 83.565 156.460 83.855 156.505 ;
        RECT 81.705 156.320 83.855 156.460 ;
        RECT 81.705 156.275 81.995 156.320 ;
        RECT 83.565 156.275 83.855 156.320 ;
        RECT 84.015 156.460 84.335 156.520 ;
        RECT 85.485 156.460 85.625 157.000 ;
        RECT 87.020 156.955 87.310 157.000 ;
        RECT 89.535 156.940 89.855 157.000 ;
        RECT 89.995 157.140 90.315 157.200 ;
        RECT 94.150 157.140 94.440 157.185 ;
        RECT 94.595 157.140 94.915 157.200 ;
        RECT 89.995 157.000 93.905 157.140 ;
        RECT 89.995 156.940 90.315 157.000 ;
        RECT 85.870 156.615 86.160 156.845 ;
        RECT 90.885 156.800 91.175 156.845 ;
        RECT 93.765 156.800 93.905 157.000 ;
        RECT 94.150 157.000 94.915 157.140 ;
        RECT 94.150 156.955 94.440 157.000 ;
        RECT 94.595 156.940 94.915 157.000 ;
        RECT 97.355 156.940 97.675 157.200 ;
        RECT 95.990 156.800 96.280 156.845 ;
        RECT 101.280 156.800 101.570 156.845 ;
        RECT 90.885 156.660 93.420 156.800 ;
        RECT 93.765 156.660 96.280 156.800 ;
        RECT 90.885 156.615 91.175 156.660 ;
        RECT 84.015 156.320 85.625 156.460 ;
        RECT 84.015 156.260 84.335 156.320 ;
        RECT 49.515 155.980 57.195 156.120 ;
        RECT 49.515 155.920 49.835 155.980 ;
        RECT 56.875 155.920 57.195 155.980 ;
        RECT 60.110 155.935 60.400 156.165 ;
        RECT 61.475 156.120 61.795 156.180 ;
        RECT 62.870 156.120 63.160 156.165 ;
        RECT 61.475 155.980 63.160 156.120 ;
        RECT 61.475 155.920 61.795 155.980 ;
        RECT 62.870 155.935 63.160 155.980 ;
        RECT 63.315 156.120 63.635 156.180 ;
        RECT 65.170 156.120 65.460 156.165 ;
        RECT 63.315 155.980 65.460 156.120 ;
        RECT 63.315 155.920 63.635 155.980 ;
        RECT 65.170 155.935 65.460 155.980 ;
        RECT 72.990 156.120 73.280 156.165 ;
        RECT 73.435 156.120 73.755 156.180 ;
        RECT 75.520 156.120 75.810 156.165 ;
        RECT 78.035 156.120 78.355 156.180 ;
        RECT 72.990 155.980 78.355 156.120 ;
        RECT 72.990 155.935 73.280 155.980 ;
        RECT 73.435 155.920 73.755 155.980 ;
        RECT 75.520 155.935 75.810 155.980 ;
        RECT 78.035 155.920 78.355 155.980 ;
        RECT 80.335 156.120 80.655 156.180 ;
        RECT 85.945 156.120 86.085 156.615 ;
        RECT 89.025 156.460 89.315 156.505 ;
        RECT 90.455 156.460 90.775 156.520 ;
        RECT 93.205 156.505 93.420 156.660 ;
        RECT 95.990 156.615 96.280 156.660 ;
        RECT 99.285 156.660 101.570 156.800 ;
        RECT 92.285 156.460 92.575 156.505 ;
        RECT 89.025 156.320 92.575 156.460 ;
        RECT 89.025 156.275 89.315 156.320 ;
        RECT 90.455 156.260 90.775 156.320 ;
        RECT 92.285 156.275 92.575 156.320 ;
        RECT 93.205 156.460 93.495 156.505 ;
        RECT 95.065 156.460 95.355 156.505 ;
        RECT 93.205 156.320 95.355 156.460 ;
        RECT 93.205 156.275 93.495 156.320 ;
        RECT 95.065 156.275 95.355 156.320 ;
        RECT 97.815 156.460 98.135 156.520 ;
        RECT 98.750 156.460 99.040 156.505 ;
        RECT 97.815 156.320 99.040 156.460 ;
        RECT 97.815 156.260 98.135 156.320 ;
        RECT 98.750 156.275 99.040 156.320 ;
        RECT 80.335 155.980 86.085 156.120 ;
        RECT 93.675 156.120 93.995 156.180 ;
        RECT 98.290 156.120 98.580 156.165 ;
        RECT 99.285 156.120 99.425 156.660 ;
        RECT 101.280 156.615 101.570 156.660 ;
        RECT 105.145 156.800 105.435 156.845 ;
        RECT 105.145 156.660 107.680 156.800 ;
        RECT 105.145 156.615 105.435 156.660 ;
        RECT 103.285 156.460 103.575 156.505 ;
        RECT 104.715 156.460 105.035 156.520 ;
        RECT 107.465 156.505 107.680 156.660 ;
        RECT 108.395 156.600 108.715 156.860 ;
        RECT 109.775 156.800 110.095 156.860 ;
        RECT 110.250 156.800 110.540 156.845 ;
        RECT 109.775 156.660 110.540 156.800 ;
        RECT 109.775 156.600 110.095 156.660 ;
        RECT 110.250 156.615 110.540 156.660 ;
        RECT 106.545 156.460 106.835 156.505 ;
        RECT 103.285 156.320 106.835 156.460 ;
        RECT 103.285 156.275 103.575 156.320 ;
        RECT 104.715 156.260 105.035 156.320 ;
        RECT 106.545 156.275 106.835 156.320 ;
        RECT 107.465 156.460 107.755 156.505 ;
        RECT 109.325 156.460 109.615 156.505 ;
        RECT 107.465 156.320 109.615 156.460 ;
        RECT 107.465 156.275 107.755 156.320 ;
        RECT 109.325 156.275 109.615 156.320 ;
        RECT 93.675 155.980 99.425 156.120 ;
        RECT 100.590 156.120 100.880 156.165 ;
        RECT 101.035 156.120 101.355 156.180 ;
        RECT 100.590 155.980 101.355 156.120 ;
        RECT 80.335 155.920 80.655 155.980 ;
        RECT 93.675 155.920 93.995 155.980 ;
        RECT 98.290 155.935 98.580 155.980 ;
        RECT 100.590 155.935 100.880 155.980 ;
        RECT 101.035 155.920 101.355 155.980 ;
        RECT 17.370 155.300 112.465 155.780 ;
        RECT 39.855 155.100 40.175 155.160 ;
        RECT 40.775 155.100 41.095 155.160 ;
        RECT 39.855 154.960 41.095 155.100 ;
        RECT 39.855 154.900 40.175 154.960 ;
        RECT 40.775 154.900 41.095 154.960 ;
        RECT 45.835 155.100 46.155 155.160 ;
        RECT 45.835 154.960 47.905 155.100 ;
        RECT 66.995 155.010 67.315 155.160 ;
        RECT 45.835 154.900 46.155 154.960 ;
        RECT 26.070 154.760 26.360 154.805 ;
        RECT 27.435 154.760 27.755 154.820 ;
        RECT 26.070 154.620 27.755 154.760 ;
        RECT 26.070 154.575 26.360 154.620 ;
        RECT 27.435 154.560 27.755 154.620 ;
        RECT 38.935 154.560 39.255 154.820 ;
        RECT 39.395 154.760 39.715 154.820 ;
        RECT 47.765 154.760 47.905 154.960 ;
        RECT 66.855 154.900 67.315 155.010 ;
        RECT 67.915 154.900 68.235 155.160 ;
        RECT 73.895 155.100 74.215 155.160 ;
        RECT 70.765 154.960 74.215 155.100 ;
        RECT 66.855 154.870 67.225 154.900 ;
        RECT 58.715 154.805 59.035 154.820 ;
        RECT 55.445 154.760 55.735 154.805 ;
        RECT 58.705 154.760 59.035 154.805 ;
        RECT 39.395 154.620 45.145 154.760 ;
        RECT 47.765 154.620 50.205 154.760 ;
        RECT 39.395 154.560 39.715 154.620 ;
        RECT 22.850 154.420 23.140 154.465 ;
        RECT 26.515 154.420 26.835 154.480 ;
        RECT 28.355 154.420 28.675 154.480 ;
        RECT 22.850 154.280 24.445 154.420 ;
        RECT 22.850 154.235 23.140 154.280 ;
        RECT 24.305 153.785 24.445 154.280 ;
        RECT 26.515 154.280 28.675 154.420 ;
        RECT 26.515 154.220 26.835 154.280 ;
        RECT 28.355 154.220 28.675 154.280 ;
        RECT 38.475 154.420 38.795 154.480 ;
        RECT 42.615 154.420 42.935 154.480 ;
        RECT 43.090 154.420 43.380 154.465 ;
        RECT 38.475 154.280 43.380 154.420 ;
        RECT 38.475 154.220 38.795 154.280 ;
        RECT 42.615 154.220 42.935 154.280 ;
        RECT 43.090 154.235 43.380 154.280 ;
        RECT 43.535 154.220 43.855 154.480 ;
        RECT 45.005 154.465 45.145 154.620 ;
        RECT 44.010 154.235 44.300 154.465 ;
        RECT 44.930 154.235 45.220 154.465 ;
        RECT 27.450 153.895 27.740 154.125 ;
        RECT 32.035 154.080 32.355 154.140 ;
        RECT 44.085 154.080 44.225 154.235 ;
        RECT 32.035 153.940 44.225 154.080 ;
        RECT 24.230 153.555 24.520 153.785 ;
        RECT 27.525 153.740 27.665 153.895 ;
        RECT 32.035 153.880 32.355 153.940 ;
        RECT 45.005 153.740 45.145 154.235 ;
        RECT 49.515 154.220 49.835 154.480 ;
        RECT 50.065 154.465 50.205 154.620 ;
        RECT 55.445 154.620 59.035 154.760 ;
        RECT 55.445 154.575 55.735 154.620 ;
        RECT 58.705 154.575 59.035 154.620 ;
        RECT 58.715 154.560 59.035 154.575 ;
        RECT 59.625 154.760 59.915 154.805 ;
        RECT 61.485 154.760 61.775 154.805 ;
        RECT 59.625 154.620 61.775 154.760 ;
        RECT 59.625 154.575 59.915 154.620 ;
        RECT 61.485 154.575 61.775 154.620 ;
        RECT 62.395 154.760 62.715 154.820 ;
        RECT 62.395 154.620 64.925 154.760 ;
        RECT 49.990 154.235 50.280 154.465 ;
        RECT 50.435 154.220 50.755 154.480 ;
        RECT 51.370 154.235 51.660 154.465 ;
        RECT 57.305 154.420 57.595 154.465 ;
        RECT 59.625 154.420 59.840 154.575 ;
        RECT 62.395 154.560 62.715 154.620 ;
        RECT 57.305 154.280 59.840 154.420 ;
        RECT 57.305 154.235 57.595 154.280 ;
        RECT 47.215 154.080 47.535 154.140 ;
        RECT 51.445 154.080 51.585 154.235 ;
        RECT 60.555 154.220 60.875 154.480 ;
        RECT 61.935 154.420 62.255 154.480 ;
        RECT 62.870 154.420 63.160 154.465 ;
        RECT 61.935 154.280 63.160 154.420 ;
        RECT 64.785 154.450 64.925 154.620 ;
        RECT 66.855 154.480 66.995 154.870 ;
        RECT 68.005 154.760 68.145 154.900 ;
        RECT 70.765 154.760 70.905 154.960 ;
        RECT 73.895 154.900 74.215 154.960 ;
        RECT 78.035 154.900 78.355 155.160 ;
        RECT 80.335 154.900 80.655 155.160 ;
        RECT 87.235 155.100 87.555 155.160 ;
        RECT 101.955 155.100 102.275 155.160 ;
        RECT 87.235 154.960 87.925 155.100 ;
        RECT 87.235 154.900 87.555 154.960 ;
        RECT 75.275 154.760 75.595 154.820 ;
        RECT 81.255 154.760 81.575 154.820 ;
        RECT 84.935 154.760 85.255 154.820 ;
        RECT 68.005 154.620 70.905 154.760 ;
        RECT 71.225 154.620 74.585 154.760 ;
        RECT 65.600 154.450 65.890 154.465 ;
        RECT 64.785 154.310 65.890 154.450 ;
        RECT 61.935 154.220 62.255 154.280 ;
        RECT 62.870 154.235 63.160 154.280 ;
        RECT 65.600 154.235 65.890 154.310 ;
        RECT 66.090 154.235 66.380 154.465 ;
        RECT 66.855 154.300 67.275 154.480 ;
        RECT 66.985 154.250 67.275 154.300 ;
        RECT 67.470 154.235 67.760 154.465 ;
        RECT 67.930 154.435 68.220 154.465 ;
        RECT 68.465 154.435 68.605 154.620 ;
        RECT 67.930 154.295 68.605 154.435 ;
        RECT 67.930 154.235 68.220 154.295 ;
        RECT 51.815 154.080 52.135 154.140 ;
        RECT 47.215 153.940 52.135 154.080 ;
        RECT 47.215 153.880 47.535 153.940 ;
        RECT 51.815 153.880 52.135 153.940 ;
        RECT 57.795 154.080 58.115 154.140 ;
        RECT 62.410 154.080 62.700 154.125 ;
        RECT 57.795 153.940 62.700 154.080 ;
        RECT 57.795 153.880 58.115 153.940 ;
        RECT 62.410 153.895 62.700 153.940 ;
        RECT 63.315 154.080 63.635 154.140 ;
        RECT 66.165 154.080 66.305 154.235 ;
        RECT 63.315 153.940 66.305 154.080 ;
        RECT 66.535 154.080 66.855 154.140 ;
        RECT 67.545 154.080 67.685 154.235 ;
        RECT 69.755 154.220 70.075 154.480 ;
        RECT 71.225 154.465 71.365 154.620 ;
        RECT 70.690 154.420 70.980 154.465 ;
        RECT 70.635 154.235 70.980 154.420 ;
        RECT 71.150 154.235 71.440 154.465 ;
        RECT 71.610 154.420 71.900 154.465 ;
        RECT 73.895 154.420 74.215 154.480 ;
        RECT 71.610 154.280 74.215 154.420 ;
        RECT 74.445 154.420 74.585 154.620 ;
        RECT 75.275 154.620 85.255 154.760 ;
        RECT 75.275 154.560 75.595 154.620 ;
        RECT 74.445 154.280 75.505 154.420 ;
        RECT 71.610 154.235 71.900 154.280 ;
        RECT 66.535 153.940 67.685 154.080 ;
        RECT 63.315 153.880 63.635 153.940 ;
        RECT 66.535 153.880 66.855 153.940 ;
        RECT 57.305 153.740 57.595 153.785 ;
        RECT 60.085 153.740 60.375 153.785 ;
        RECT 61.945 153.740 62.235 153.785 ;
        RECT 27.525 153.600 32.265 153.740 ;
        RECT 45.005 153.600 57.105 153.740 ;
        RECT 32.125 153.460 32.265 153.600 ;
        RECT 23.770 153.400 24.060 153.445 ;
        RECT 26.975 153.400 27.295 153.460 ;
        RECT 23.770 153.260 27.295 153.400 ;
        RECT 23.770 153.215 24.060 153.260 ;
        RECT 26.975 153.200 27.295 153.260 ;
        RECT 31.575 153.200 31.895 153.460 ;
        RECT 32.035 153.200 32.355 153.460 ;
        RECT 39.395 153.400 39.715 153.460 ;
        RECT 41.710 153.400 42.000 153.445 ;
        RECT 39.395 153.260 42.000 153.400 ;
        RECT 39.395 153.200 39.715 153.260 ;
        RECT 41.710 153.215 42.000 153.260 ;
        RECT 47.215 153.400 47.535 153.460 ;
        RECT 48.150 153.400 48.440 153.445 ;
        RECT 47.215 153.260 48.440 153.400 ;
        RECT 47.215 153.200 47.535 153.260 ;
        RECT 48.150 153.215 48.440 153.260 ;
        RECT 53.440 153.400 53.730 153.445 ;
        RECT 54.575 153.400 54.895 153.460 ;
        RECT 53.440 153.260 54.895 153.400 ;
        RECT 56.965 153.400 57.105 153.600 ;
        RECT 57.305 153.600 62.235 153.740 ;
        RECT 57.305 153.555 57.595 153.600 ;
        RECT 60.085 153.555 60.375 153.600 ;
        RECT 61.945 153.555 62.235 153.600 ;
        RECT 63.790 153.740 64.080 153.785 ;
        RECT 66.995 153.740 67.315 153.800 ;
        RECT 63.790 153.600 67.315 153.740 ;
        RECT 69.845 153.740 69.985 154.220 ;
        RECT 70.635 154.080 70.775 154.235 ;
        RECT 73.895 154.220 74.215 154.280 ;
        RECT 75.365 154.140 75.505 154.280 ;
        RECT 75.735 154.220 76.055 154.480 ;
        RECT 73.435 154.080 73.755 154.140 ;
        RECT 70.635 153.940 73.755 154.080 ;
        RECT 73.435 153.880 73.755 153.940 ;
        RECT 75.275 153.880 75.595 154.140 ;
        RECT 77.665 154.125 77.805 154.620 ;
        RECT 81.255 154.560 81.575 154.620 ;
        RECT 84.935 154.560 85.255 154.620 ;
        RECT 78.510 154.420 78.800 154.465 ;
        RECT 78.955 154.420 79.275 154.480 ;
        RECT 78.510 154.280 79.275 154.420 ;
        RECT 78.510 154.235 78.800 154.280 ;
        RECT 78.955 154.220 79.275 154.280 ;
        RECT 81.715 154.220 82.035 154.480 ;
        RECT 87.785 154.420 87.925 154.960 ;
        RECT 97.445 154.960 102.275 155.100 ;
        RECT 88.615 154.760 88.935 154.820 ;
        RECT 91.375 154.760 91.695 154.820 ;
        RECT 97.445 154.760 97.585 154.960 ;
        RECT 88.615 154.620 91.695 154.760 ;
        RECT 88.615 154.560 88.935 154.620 ;
        RECT 91.375 154.560 91.695 154.620 ;
        RECT 92.385 154.620 97.585 154.760 ;
        RECT 92.385 154.465 92.525 154.620 ;
        RECT 92.310 154.420 92.600 154.465 ;
        RECT 87.785 154.280 92.600 154.420 ;
        RECT 92.310 154.235 92.600 154.280 ;
        RECT 92.755 154.220 93.075 154.480 ;
        RECT 93.215 154.220 93.535 154.480 ;
        RECT 94.150 154.420 94.440 154.465 ;
        RECT 95.530 154.420 95.820 154.465 ;
        RECT 95.975 154.420 96.295 154.480 ;
        RECT 94.150 154.280 96.295 154.420 ;
        RECT 94.150 154.235 94.440 154.280 ;
        RECT 95.530 154.235 95.820 154.280 ;
        RECT 77.590 153.895 77.880 154.125 ;
        RECT 85.855 154.080 86.175 154.140 ;
        RECT 94.225 154.080 94.365 154.235 ;
        RECT 95.975 154.220 96.295 154.280 ;
        RECT 96.435 154.220 96.755 154.480 ;
        RECT 97.445 154.465 97.585 154.620 ;
        RECT 98.275 154.760 98.595 154.820 ;
        RECT 98.750 154.760 99.040 154.805 ;
        RECT 98.275 154.620 99.040 154.760 ;
        RECT 98.275 154.560 98.595 154.620 ;
        RECT 98.750 154.575 99.040 154.620 ;
        RECT 99.195 154.760 99.515 154.820 ;
        RECT 99.195 154.620 100.805 154.760 ;
        RECT 99.195 154.560 99.515 154.620 ;
        RECT 100.665 154.465 100.805 154.620 ;
        RECT 101.585 154.465 101.725 154.960 ;
        RECT 101.955 154.900 102.275 154.960 ;
        RECT 104.255 154.760 104.575 154.820 ;
        RECT 102.045 154.620 104.575 154.760 ;
        RECT 102.045 154.480 102.185 154.620 ;
        RECT 104.255 154.560 104.575 154.620 ;
        RECT 96.910 154.235 97.200 154.465 ;
        RECT 97.370 154.235 97.660 154.465 ;
        RECT 99.670 154.420 99.960 154.465 ;
        RECT 98.825 154.280 99.960 154.420 ;
        RECT 85.855 153.940 94.365 154.080 ;
        RECT 85.855 153.880 86.175 153.940 ;
        RECT 72.515 153.740 72.835 153.800 ;
        RECT 69.845 153.600 72.835 153.740 ;
        RECT 63.790 153.555 64.080 153.600 ;
        RECT 66.995 153.540 67.315 153.600 ;
        RECT 72.515 153.540 72.835 153.600 ;
        RECT 88.615 153.740 88.935 153.800 ;
        RECT 94.135 153.740 94.455 153.800 ;
        RECT 88.615 153.600 94.455 153.740 ;
        RECT 96.985 153.740 97.125 154.235 ;
        RECT 98.825 154.140 98.965 154.280 ;
        RECT 99.670 154.235 99.960 154.280 ;
        RECT 100.590 154.235 100.880 154.465 ;
        RECT 101.050 154.235 101.340 154.465 ;
        RECT 101.510 154.235 101.800 154.465 ;
        RECT 98.735 153.880 99.055 154.140 ;
        RECT 101.125 153.740 101.265 154.235 ;
        RECT 101.955 154.220 102.275 154.480 ;
        RECT 102.415 154.420 102.735 154.480 ;
        RECT 105.635 154.420 105.955 154.480 ;
        RECT 102.415 154.280 105.955 154.420 ;
        RECT 102.415 154.220 102.735 154.280 ;
        RECT 105.635 154.220 105.955 154.280 ;
        RECT 106.110 154.235 106.400 154.465 ;
        RECT 96.985 153.600 101.265 153.740 ;
        RECT 101.495 153.740 101.815 153.800 ;
        RECT 106.185 153.740 106.325 154.235 ;
        RECT 101.495 153.600 106.325 153.740 ;
        RECT 107.030 153.740 107.320 153.785 ;
        RECT 108.395 153.740 108.715 153.800 ;
        RECT 107.030 153.600 108.715 153.740 ;
        RECT 88.615 153.540 88.935 153.600 ;
        RECT 94.135 153.540 94.455 153.600 ;
        RECT 63.315 153.400 63.635 153.460 ;
        RECT 56.965 153.260 63.635 153.400 ;
        RECT 53.440 153.215 53.730 153.260 ;
        RECT 54.575 153.200 54.895 153.260 ;
        RECT 63.315 153.200 63.635 153.260 ;
        RECT 64.695 153.400 65.015 153.460 ;
        RECT 68.835 153.400 69.155 153.460 ;
        RECT 64.695 153.260 69.155 153.400 ;
        RECT 64.695 153.200 65.015 153.260 ;
        RECT 68.835 153.200 69.155 153.260 ;
        RECT 69.310 153.400 69.600 153.445 ;
        RECT 69.755 153.400 70.075 153.460 ;
        RECT 69.310 153.260 70.075 153.400 ;
        RECT 69.310 153.215 69.600 153.260 ;
        RECT 69.755 153.200 70.075 153.260 ;
        RECT 72.055 153.400 72.375 153.460 ;
        RECT 72.990 153.400 73.280 153.445 ;
        RECT 72.055 153.260 73.280 153.400 ;
        RECT 72.055 153.200 72.375 153.260 ;
        RECT 72.990 153.215 73.280 153.260 ;
        RECT 73.435 153.400 73.755 153.460 ;
        RECT 74.370 153.400 74.660 153.445 ;
        RECT 73.435 153.260 74.660 153.400 ;
        RECT 73.435 153.200 73.755 153.260 ;
        RECT 74.370 153.215 74.660 153.260 ;
        RECT 85.855 153.400 86.175 153.460 ;
        RECT 88.170 153.400 88.460 153.445 ;
        RECT 89.995 153.400 90.315 153.460 ;
        RECT 85.855 153.260 90.315 153.400 ;
        RECT 85.855 153.200 86.175 153.260 ;
        RECT 88.170 153.215 88.460 153.260 ;
        RECT 89.995 153.200 90.315 153.260 ;
        RECT 90.930 153.400 91.220 153.445 ;
        RECT 91.375 153.400 91.695 153.460 ;
        RECT 90.930 153.260 91.695 153.400 ;
        RECT 90.930 153.215 91.220 153.260 ;
        RECT 91.375 153.200 91.695 153.260 ;
        RECT 92.755 153.400 93.075 153.460 ;
        RECT 97.445 153.400 97.585 153.600 ;
        RECT 101.495 153.540 101.815 153.600 ;
        RECT 107.030 153.555 107.320 153.600 ;
        RECT 108.395 153.540 108.715 153.600 ;
        RECT 92.755 153.260 97.585 153.400 ;
        RECT 97.815 153.400 98.135 153.460 ;
        RECT 102.890 153.400 103.180 153.445 ;
        RECT 97.815 153.260 103.180 153.400 ;
        RECT 92.755 153.200 93.075 153.260 ;
        RECT 97.815 153.200 98.135 153.260 ;
        RECT 102.890 153.215 103.180 153.260 ;
        RECT 18.165 152.580 112.465 153.060 ;
        RECT 28.355 152.380 28.675 152.440 ;
        RECT 51.815 152.380 52.135 152.440 ;
        RECT 60.555 152.380 60.875 152.440 ;
        RECT 61.030 152.380 61.320 152.425 ;
        RECT 28.355 152.240 40.085 152.380 ;
        RECT 28.355 152.180 28.675 152.240 ;
        RECT 21.880 152.040 22.170 152.085 ;
        RECT 23.770 152.040 24.060 152.085 ;
        RECT 26.890 152.040 27.180 152.085 ;
        RECT 21.880 151.900 27.180 152.040 ;
        RECT 21.880 151.855 22.170 151.900 ;
        RECT 23.770 151.855 24.060 151.900 ;
        RECT 26.890 151.855 27.180 151.900 ;
        RECT 27.435 152.040 27.755 152.100 ;
        RECT 29.750 152.040 30.040 152.085 ;
        RECT 38.475 152.040 38.795 152.100 ;
        RECT 27.435 151.900 38.795 152.040 ;
        RECT 27.435 151.840 27.755 151.900 ;
        RECT 29.750 151.855 30.040 151.900 ;
        RECT 38.475 151.840 38.795 151.900 ;
        RECT 20.090 151.700 20.380 151.745 ;
        RECT 28.355 151.700 28.675 151.760 ;
        RECT 31.590 151.700 31.880 151.745 ;
        RECT 32.035 151.700 32.355 151.760 ;
        RECT 36.635 151.700 36.955 151.760 ;
        RECT 20.090 151.560 28.125 151.700 ;
        RECT 20.090 151.515 20.380 151.560 ;
        RECT 20.535 151.160 20.855 151.420 ;
        RECT 21.010 151.175 21.300 151.405 ;
        RECT 21.475 151.360 21.765 151.405 ;
        RECT 23.310 151.360 23.600 151.405 ;
        RECT 26.890 151.360 27.180 151.405 ;
        RECT 27.985 151.380 28.125 151.560 ;
        RECT 28.355 151.560 36.955 151.700 ;
        RECT 28.355 151.500 28.675 151.560 ;
        RECT 31.590 151.515 31.880 151.560 ;
        RECT 32.035 151.500 32.355 151.560 ;
        RECT 36.635 151.500 36.955 151.560 ;
        RECT 21.475 151.220 27.180 151.360 ;
        RECT 21.475 151.175 21.765 151.220 ;
        RECT 23.310 151.175 23.600 151.220 ;
        RECT 26.890 151.175 27.180 151.220 ;
        RECT 21.085 150.680 21.225 151.175 ;
        RECT 22.375 150.820 22.695 151.080 ;
        RECT 27.970 151.065 28.260 151.380 ;
        RECT 28.815 151.360 29.135 151.420 ;
        RECT 32.510 151.360 32.800 151.405 ;
        RECT 37.095 151.360 37.415 151.420 ;
        RECT 28.815 151.220 37.415 151.360 ;
        RECT 28.815 151.160 29.135 151.220 ;
        RECT 32.510 151.175 32.800 151.220 ;
        RECT 37.095 151.160 37.415 151.220 ;
        RECT 37.570 151.360 37.860 151.405 ;
        RECT 39.025 151.360 39.165 152.240 ;
        RECT 39.410 151.855 39.700 152.085 ;
        RECT 39.945 152.040 40.085 152.240 ;
        RECT 51.815 152.240 60.325 152.380 ;
        RECT 51.815 152.180 52.135 152.240 ;
        RECT 55.005 152.040 55.295 152.085 ;
        RECT 57.785 152.040 58.075 152.085 ;
        RECT 59.645 152.040 59.935 152.085 ;
        RECT 39.945 151.900 46.525 152.040 ;
        RECT 37.570 151.220 39.165 151.360 ;
        RECT 39.485 151.360 39.625 151.855 ;
        RECT 40.790 151.360 41.080 151.405 ;
        RECT 39.485 151.220 41.080 151.360 ;
        RECT 37.570 151.175 37.860 151.220 ;
        RECT 40.790 151.175 41.080 151.220 ;
        RECT 42.615 151.360 42.935 151.420 ;
        RECT 43.090 151.360 43.380 151.405 ;
        RECT 42.615 151.220 43.380 151.360 ;
        RECT 42.615 151.160 42.935 151.220 ;
        RECT 43.090 151.175 43.380 151.220 ;
        RECT 43.535 151.160 43.855 151.420 ;
        RECT 43.995 151.160 44.315 151.420 ;
        RECT 46.385 151.405 46.525 151.900 ;
        RECT 55.005 151.900 59.935 152.040 ;
        RECT 60.185 152.040 60.325 152.240 ;
        RECT 60.555 152.240 61.320 152.380 ;
        RECT 60.555 152.180 60.875 152.240 ;
        RECT 61.030 152.195 61.320 152.240 ;
        RECT 61.475 152.380 61.795 152.440 ;
        RECT 65.170 152.380 65.460 152.425 ;
        RECT 61.475 152.240 65.460 152.380 ;
        RECT 61.475 152.180 61.795 152.240 ;
        RECT 65.170 152.195 65.460 152.240 ;
        RECT 72.515 152.380 72.835 152.440 ;
        RECT 88.170 152.380 88.460 152.425 ;
        RECT 90.455 152.380 90.775 152.440 ;
        RECT 72.515 152.240 75.965 152.380 ;
        RECT 72.515 152.180 72.835 152.240 ;
        RECT 64.695 152.040 65.015 152.100 ;
        RECT 60.185 151.900 65.015 152.040 ;
        RECT 55.005 151.855 55.295 151.900 ;
        RECT 57.785 151.855 58.075 151.900 ;
        RECT 59.645 151.855 59.935 151.900 ;
        RECT 64.695 151.840 65.015 151.900 ;
        RECT 66.075 152.040 66.395 152.100 ;
        RECT 75.275 152.040 75.595 152.100 ;
        RECT 66.075 151.900 75.595 152.040 ;
        RECT 66.075 151.840 66.395 151.900 ;
        RECT 58.270 151.700 58.560 151.745 ;
        RECT 60.555 151.700 60.875 151.760 ;
        RECT 58.270 151.560 60.875 151.700 ;
        RECT 58.270 151.515 58.560 151.560 ;
        RECT 60.555 151.500 60.875 151.560 ;
        RECT 62.855 151.700 63.175 151.760 ;
        RECT 62.855 151.560 66.305 151.700 ;
        RECT 62.855 151.500 63.175 151.560 ;
        RECT 44.930 151.360 45.220 151.405 ;
        RECT 45.390 151.360 45.680 151.405 ;
        RECT 44.930 151.220 45.680 151.360 ;
        RECT 44.930 151.175 45.220 151.220 ;
        RECT 45.390 151.175 45.680 151.220 ;
        RECT 46.310 151.175 46.600 151.405 ;
        RECT 24.670 151.020 25.320 151.065 ;
        RECT 27.970 151.020 28.560 151.065 ;
        RECT 24.670 150.880 28.560 151.020 ;
        RECT 24.670 150.835 25.320 150.880 ;
        RECT 28.270 150.835 28.560 150.880 ;
        RECT 32.050 151.020 32.340 151.065 ;
        RECT 45.465 151.020 45.605 151.175 ;
        RECT 46.755 151.160 47.075 151.420 ;
        RECT 47.230 151.360 47.520 151.405 ;
        RECT 47.675 151.360 47.995 151.420 ;
        RECT 47.230 151.220 47.995 151.360 ;
        RECT 47.230 151.175 47.520 151.220 ;
        RECT 47.675 151.160 47.995 151.220 ;
        RECT 55.005 151.360 55.295 151.405 ;
        RECT 57.795 151.360 58.115 151.420 ;
        RECT 60.110 151.360 60.400 151.405 ;
        RECT 55.005 151.220 57.540 151.360 ;
        RECT 55.005 151.175 55.295 151.220 ;
        RECT 48.135 151.020 48.455 151.080 ;
        RECT 57.325 151.065 57.540 151.220 ;
        RECT 57.795 151.220 60.400 151.360 ;
        RECT 57.795 151.160 58.115 151.220 ;
        RECT 60.110 151.175 60.400 151.220 ;
        RECT 61.935 151.160 62.255 151.420 ;
        RECT 63.315 151.160 63.635 151.420 ;
        RECT 66.165 151.405 66.305 151.560 ;
        RECT 64.250 151.175 64.540 151.405 ;
        RECT 66.090 151.175 66.380 151.405 ;
        RECT 68.835 151.360 69.155 151.420 ;
        RECT 70.765 151.405 70.905 151.900 ;
        RECT 71.225 151.560 73.665 151.700 ;
        RECT 71.225 151.405 71.365 151.560 ;
        RECT 70.230 151.360 70.520 151.405 ;
        RECT 68.835 151.220 70.520 151.360 ;
        RECT 32.050 150.880 39.165 151.020 ;
        RECT 45.465 150.880 48.455 151.020 ;
        RECT 32.050 150.835 32.340 150.880 ;
        RECT 39.025 150.740 39.165 150.880 ;
        RECT 48.135 150.820 48.455 150.880 ;
        RECT 53.145 151.020 53.435 151.065 ;
        RECT 56.405 151.020 56.695 151.065 ;
        RECT 57.325 151.020 57.615 151.065 ;
        RECT 59.185 151.020 59.475 151.065 ;
        RECT 53.145 150.880 57.105 151.020 ;
        RECT 53.145 150.835 53.435 150.880 ;
        RECT 56.405 150.835 56.695 150.880 ;
        RECT 31.575 150.680 31.895 150.740 ;
        RECT 21.085 150.540 31.895 150.680 ;
        RECT 31.575 150.480 31.895 150.540 ;
        RECT 34.335 150.480 34.655 150.740 ;
        RECT 37.095 150.480 37.415 150.740 ;
        RECT 38.935 150.480 39.255 150.740 ;
        RECT 39.870 150.680 40.160 150.725 ;
        RECT 40.775 150.680 41.095 150.740 ;
        RECT 39.870 150.540 41.095 150.680 ;
        RECT 39.870 150.495 40.160 150.540 ;
        RECT 40.775 150.480 41.095 150.540 ;
        RECT 41.710 150.680 42.000 150.725 ;
        RECT 42.615 150.680 42.935 150.740 ;
        RECT 41.710 150.540 42.935 150.680 ;
        RECT 41.710 150.495 42.000 150.540 ;
        RECT 42.615 150.480 42.935 150.540 ;
        RECT 48.610 150.680 48.900 150.725 ;
        RECT 49.055 150.680 49.375 150.740 ;
        RECT 48.610 150.540 49.375 150.680 ;
        RECT 48.610 150.495 48.900 150.540 ;
        RECT 49.055 150.480 49.375 150.540 ;
        RECT 50.895 150.725 51.215 150.740 ;
        RECT 50.895 150.495 51.430 150.725 ;
        RECT 56.965 150.680 57.105 150.880 ;
        RECT 57.325 150.880 59.475 151.020 ;
        RECT 57.325 150.835 57.615 150.880 ;
        RECT 59.185 150.835 59.475 150.880 ;
        RECT 59.635 151.020 59.955 151.080 ;
        RECT 64.325 151.020 64.465 151.175 ;
        RECT 68.835 151.160 69.155 151.220 ;
        RECT 70.230 151.175 70.520 151.220 ;
        RECT 70.690 151.175 70.980 151.405 ;
        RECT 71.150 151.175 71.440 151.405 ;
        RECT 72.070 151.360 72.360 151.405 ;
        RECT 72.515 151.360 72.835 151.420 ;
        RECT 72.070 151.220 72.835 151.360 ;
        RECT 72.070 151.175 72.360 151.220 ;
        RECT 72.515 151.160 72.835 151.220 ;
        RECT 71.595 151.020 71.915 151.080 ;
        RECT 59.635 150.880 71.915 151.020 ;
        RECT 59.635 150.820 59.955 150.880 ;
        RECT 71.595 150.820 71.915 150.880 ;
        RECT 62.870 150.680 63.160 150.725 ;
        RECT 56.965 150.540 63.160 150.680 ;
        RECT 62.870 150.495 63.160 150.540 ;
        RECT 67.010 150.680 67.300 150.725 ;
        RECT 67.455 150.680 67.775 150.740 ;
        RECT 67.010 150.540 67.775 150.680 ;
        RECT 67.010 150.495 67.300 150.540 ;
        RECT 50.895 150.480 51.215 150.495 ;
        RECT 67.455 150.480 67.775 150.540 ;
        RECT 68.835 150.480 69.155 150.740 ;
        RECT 72.515 150.480 72.835 150.740 ;
        RECT 73.525 150.680 73.665 151.560 ;
        RECT 73.895 151.160 74.215 151.420 ;
        RECT 74.445 151.405 74.585 151.900 ;
        RECT 75.275 151.840 75.595 151.900 ;
        RECT 75.825 151.405 75.965 152.240 ;
        RECT 88.170 152.240 90.775 152.380 ;
        RECT 88.170 152.195 88.460 152.240 ;
        RECT 90.455 152.180 90.775 152.240 ;
        RECT 93.215 152.380 93.535 152.440 ;
        RECT 95.515 152.380 95.835 152.440 ;
        RECT 93.215 152.240 95.835 152.380 ;
        RECT 93.215 152.180 93.535 152.240 ;
        RECT 95.515 152.180 95.835 152.240 ;
        RECT 80.305 152.040 80.595 152.085 ;
        RECT 83.085 152.040 83.375 152.085 ;
        RECT 84.945 152.040 85.235 152.085 ;
        RECT 90.915 152.040 91.235 152.100 ;
        RECT 80.305 151.900 85.235 152.040 ;
        RECT 80.305 151.855 80.595 151.900 ;
        RECT 83.085 151.855 83.375 151.900 ;
        RECT 84.945 151.855 85.235 151.900 ;
        RECT 90.085 151.900 91.235 152.040 ;
        RECT 74.370 151.175 74.660 151.405 ;
        RECT 74.830 151.175 75.120 151.405 ;
        RECT 75.750 151.175 76.040 151.405 ;
        RECT 80.305 151.360 80.595 151.405 ;
        RECT 83.570 151.360 83.860 151.405 ;
        RECT 84.935 151.360 85.255 151.420 ;
        RECT 80.305 151.220 82.840 151.360 ;
        RECT 80.305 151.175 80.595 151.220 ;
        RECT 73.895 150.680 74.215 150.740 ;
        RECT 73.525 150.540 74.215 150.680 ;
        RECT 74.905 150.680 75.045 151.175 ;
        RECT 78.445 151.020 78.735 151.065 ;
        RECT 79.875 151.020 80.195 151.080 ;
        RECT 82.625 151.065 82.840 151.220 ;
        RECT 83.570 151.220 85.255 151.360 ;
        RECT 83.570 151.175 83.860 151.220 ;
        RECT 84.935 151.160 85.255 151.220 ;
        RECT 85.410 151.360 85.700 151.405 ;
        RECT 85.855 151.360 86.175 151.420 ;
        RECT 85.410 151.220 86.175 151.360 ;
        RECT 85.410 151.175 85.700 151.220 ;
        RECT 85.855 151.160 86.175 151.220 ;
        RECT 87.710 151.360 88.000 151.405 ;
        RECT 88.615 151.360 88.935 151.420 ;
        RECT 87.710 151.220 88.935 151.360 ;
        RECT 87.710 151.175 88.000 151.220 ;
        RECT 81.705 151.020 81.995 151.065 ;
        RECT 78.445 150.880 81.995 151.020 ;
        RECT 78.445 150.835 78.735 150.880 ;
        RECT 79.875 150.820 80.195 150.880 ;
        RECT 81.705 150.835 81.995 150.880 ;
        RECT 82.625 151.020 82.915 151.065 ;
        RECT 84.485 151.020 84.775 151.065 ;
        RECT 82.625 150.880 84.775 151.020 ;
        RECT 82.625 150.835 82.915 150.880 ;
        RECT 84.485 150.835 84.775 150.880 ;
        RECT 76.440 150.680 76.730 150.725 ;
        RECT 78.955 150.680 79.275 150.740 ;
        RECT 82.175 150.680 82.495 150.740 ;
        RECT 74.905 150.540 82.495 150.680 ;
        RECT 73.895 150.480 74.215 150.540 ;
        RECT 76.440 150.495 76.730 150.540 ;
        RECT 78.955 150.480 79.275 150.540 ;
        RECT 82.175 150.480 82.495 150.540 ;
        RECT 83.095 150.680 83.415 150.740 ;
        RECT 87.785 150.680 87.925 151.175 ;
        RECT 88.615 151.160 88.935 151.220 ;
        RECT 89.090 151.360 89.380 151.405 ;
        RECT 89.535 151.360 89.855 151.420 ;
        RECT 90.085 151.405 90.225 151.900 ;
        RECT 90.915 151.840 91.235 151.900 ;
        RECT 104.370 152.040 104.660 152.085 ;
        RECT 107.490 152.040 107.780 152.085 ;
        RECT 109.380 152.040 109.670 152.085 ;
        RECT 104.370 151.900 109.670 152.040 ;
        RECT 104.370 151.855 104.660 151.900 ;
        RECT 107.490 151.855 107.780 151.900 ;
        RECT 109.380 151.855 109.670 151.900 ;
        RECT 96.435 151.700 96.755 151.760 ;
        RECT 90.545 151.560 94.365 151.700 ;
        RECT 90.545 151.420 90.685 151.560 ;
        RECT 89.090 151.220 89.855 151.360 ;
        RECT 89.090 151.175 89.380 151.220 ;
        RECT 89.535 151.160 89.855 151.220 ;
        RECT 90.010 151.175 90.300 151.405 ;
        RECT 90.455 151.160 90.775 151.420 ;
        RECT 90.915 151.160 91.235 151.420 ;
        RECT 92.755 151.160 93.075 151.420 ;
        RECT 93.675 151.160 93.995 151.420 ;
        RECT 94.225 151.405 94.365 151.560 ;
        RECT 96.435 151.560 99.425 151.700 ;
        RECT 96.435 151.500 96.755 151.560 ;
        RECT 94.595 151.405 94.915 151.420 ;
        RECT 94.150 151.175 94.440 151.405 ;
        RECT 94.595 151.175 95.000 151.405 ;
        RECT 95.515 151.360 95.835 151.420 ;
        RECT 97.370 151.360 97.660 151.405 ;
        RECT 95.515 151.220 97.660 151.360 ;
        RECT 94.595 151.160 94.915 151.175 ;
        RECT 95.515 151.160 95.835 151.220 ;
        RECT 97.370 151.175 97.660 151.220 ;
        RECT 98.290 151.175 98.580 151.405 ;
        RECT 98.365 151.020 98.505 151.175 ;
        RECT 98.735 151.160 99.055 151.420 ;
        RECT 99.285 151.405 99.425 151.560 ;
        RECT 110.235 151.500 110.555 151.760 ;
        RECT 99.210 151.175 99.500 151.405 ;
        RECT 103.290 151.065 103.580 151.380 ;
        RECT 104.370 151.360 104.660 151.405 ;
        RECT 107.950 151.360 108.240 151.405 ;
        RECT 109.785 151.360 110.075 151.405 ;
        RECT 104.370 151.220 110.075 151.360 ;
        RECT 104.370 151.175 104.660 151.220 ;
        RECT 107.950 151.175 108.240 151.220 ;
        RECT 109.785 151.175 110.075 151.220 ;
        RECT 102.990 151.020 103.580 151.065 ;
        RECT 106.095 151.065 106.415 151.080 ;
        RECT 106.095 151.020 106.880 151.065 ;
        RECT 98.365 150.880 101.725 151.020 ;
        RECT 83.095 150.540 87.925 150.680 ;
        RECT 92.310 150.680 92.600 150.725 ;
        RECT 93.675 150.680 93.995 150.740 ;
        RECT 92.310 150.540 93.995 150.680 ;
        RECT 83.095 150.480 83.415 150.540 ;
        RECT 92.310 150.495 92.600 150.540 ;
        RECT 93.675 150.480 93.995 150.540 ;
        RECT 95.975 150.480 96.295 150.740 ;
        RECT 99.195 150.680 99.515 150.740 ;
        RECT 101.585 150.725 101.725 150.880 ;
        RECT 102.990 150.880 106.880 151.020 ;
        RECT 102.990 150.835 103.280 150.880 ;
        RECT 106.095 150.835 106.880 150.880 ;
        RECT 106.095 150.820 106.415 150.835 ;
        RECT 108.855 150.820 109.175 151.080 ;
        RECT 100.590 150.680 100.880 150.725 ;
        RECT 99.195 150.540 100.880 150.680 ;
        RECT 99.195 150.480 99.515 150.540 ;
        RECT 100.590 150.495 100.880 150.540 ;
        RECT 101.510 150.680 101.800 150.725 ;
        RECT 104.255 150.680 104.575 150.740 ;
        RECT 101.510 150.540 104.575 150.680 ;
        RECT 101.510 150.495 101.800 150.540 ;
        RECT 104.255 150.480 104.575 150.540 ;
        RECT 17.370 149.860 112.465 150.340 ;
        RECT 22.375 149.660 22.695 149.720 ;
        RECT 23.770 149.660 24.060 149.705 ;
        RECT 22.375 149.520 24.060 149.660 ;
        RECT 22.375 149.460 22.695 149.520 ;
        RECT 23.770 149.475 24.060 149.520 ;
        RECT 25.150 149.475 25.440 149.705 ;
        RECT 20.535 148.980 20.855 149.040 ;
        RECT 22.390 148.980 22.680 149.025 ;
        RECT 20.535 148.840 22.680 148.980 ;
        RECT 20.535 148.780 20.855 148.840 ;
        RECT 22.390 148.795 22.680 148.840 ;
        RECT 24.690 148.980 24.980 149.025 ;
        RECT 25.225 148.980 25.365 149.475 ;
        RECT 27.435 149.460 27.755 149.720 ;
        RECT 29.750 149.660 30.040 149.705 ;
        RECT 31.115 149.660 31.435 149.720 ;
        RECT 29.750 149.520 31.435 149.660 ;
        RECT 29.750 149.475 30.040 149.520 ;
        RECT 31.115 149.460 31.435 149.520 ;
        RECT 53.670 149.660 53.960 149.705 ;
        RECT 54.575 149.660 54.895 149.720 ;
        RECT 53.670 149.520 54.895 149.660 ;
        RECT 53.670 149.475 53.960 149.520 ;
        RECT 54.575 149.460 54.895 149.520 ;
        RECT 60.110 149.475 60.400 149.705 ;
        RECT 31.595 149.320 31.885 149.365 ;
        RECT 33.455 149.320 33.745 149.365 ;
        RECT 31.595 149.180 33.745 149.320 ;
        RECT 31.595 149.135 31.885 149.180 ;
        RECT 33.455 149.135 33.745 149.180 ;
        RECT 34.375 149.320 34.665 149.365 ;
        RECT 35.255 149.320 35.575 149.380 ;
        RECT 37.635 149.320 37.925 149.365 ;
        RECT 34.375 149.180 37.925 149.320 ;
        RECT 34.375 149.135 34.665 149.180 ;
        RECT 24.690 148.840 25.365 148.980 ;
        RECT 24.690 148.795 24.980 148.840 ;
        RECT 22.465 148.640 22.605 148.795 ;
        RECT 26.975 148.780 27.295 149.040 ;
        RECT 29.290 148.980 29.580 149.025 ;
        RECT 32.035 148.980 32.355 149.040 ;
        RECT 27.525 148.840 32.355 148.980 ;
        RECT 27.525 148.640 27.665 148.840 ;
        RECT 29.290 148.795 29.580 148.840 ;
        RECT 32.035 148.780 32.355 148.840 ;
        RECT 32.510 148.980 32.800 149.025 ;
        RECT 32.955 148.980 33.275 149.040 ;
        RECT 32.510 148.840 33.275 148.980 ;
        RECT 33.530 148.980 33.745 149.135 ;
        RECT 35.255 149.120 35.575 149.180 ;
        RECT 37.635 149.135 37.925 149.180 ;
        RECT 38.475 149.320 38.795 149.380 ;
        RECT 54.130 149.320 54.420 149.365 ;
        RECT 57.810 149.320 58.100 149.365 ;
        RECT 38.475 149.180 46.525 149.320 ;
        RECT 38.475 149.120 38.795 149.180 ;
        RECT 35.775 148.980 36.065 149.025 ;
        RECT 33.530 148.840 36.065 148.980 ;
        RECT 32.510 148.795 32.800 148.840 ;
        RECT 32.955 148.780 33.275 148.840 ;
        RECT 35.775 148.795 36.065 148.840 ;
        RECT 40.315 148.980 40.635 149.040 ;
        RECT 40.790 148.980 41.080 149.025 ;
        RECT 40.315 148.840 41.080 148.980 ;
        RECT 40.315 148.780 40.635 148.840 ;
        RECT 40.790 148.795 41.080 148.840 ;
        RECT 45.375 148.780 45.695 149.040 ;
        RECT 45.835 148.780 46.155 149.040 ;
        RECT 46.385 149.025 46.525 149.180 ;
        RECT 50.985 149.180 58.100 149.320 ;
        RECT 50.985 149.040 51.125 149.180 ;
        RECT 54.130 149.135 54.420 149.180 ;
        RECT 57.810 149.135 58.100 149.180 ;
        RECT 46.310 148.795 46.600 149.025 ;
        RECT 47.230 148.980 47.520 149.025 ;
        RECT 48.135 148.980 48.455 149.040 ;
        RECT 47.230 148.840 48.455 148.980 ;
        RECT 47.230 148.795 47.520 148.840 ;
        RECT 48.135 148.780 48.455 148.840 ;
        RECT 49.975 148.780 50.295 149.040 ;
        RECT 50.435 148.780 50.755 149.040 ;
        RECT 50.895 148.780 51.215 149.040 ;
        RECT 51.830 148.980 52.120 149.025 ;
        RECT 52.275 148.980 52.595 149.040 ;
        RECT 51.830 148.840 52.595 148.980 ;
        RECT 51.830 148.795 52.120 148.840 ;
        RECT 52.275 148.780 52.595 148.840 ;
        RECT 58.270 148.980 58.560 149.025 ;
        RECT 58.715 148.980 59.035 149.040 ;
        RECT 58.270 148.840 59.035 148.980 ;
        RECT 60.185 148.980 60.325 149.475 ;
        RECT 60.555 149.460 60.875 149.720 ;
        RECT 61.475 149.660 61.795 149.720 ;
        RECT 64.250 149.660 64.540 149.705 ;
        RECT 61.475 149.520 64.540 149.660 ;
        RECT 61.475 149.460 61.795 149.520 ;
        RECT 64.250 149.475 64.540 149.520 ;
        RECT 71.595 149.660 71.915 149.720 ;
        RECT 72.070 149.660 72.360 149.705 ;
        RECT 71.595 149.520 72.360 149.660 ;
        RECT 71.595 149.460 71.915 149.520 ;
        RECT 72.070 149.475 72.360 149.520 ;
        RECT 79.875 149.460 80.195 149.720 ;
        RECT 82.175 149.460 82.495 149.720 ;
        RECT 84.490 149.475 84.780 149.705 ;
        RECT 62.395 149.320 62.715 149.380 ;
        RECT 73.895 149.320 74.215 149.380 ;
        RECT 82.650 149.320 82.940 149.365 ;
        RECT 84.015 149.320 84.335 149.380 ;
        RECT 62.395 149.180 69.525 149.320 ;
        RECT 62.395 149.120 62.715 149.180 ;
        RECT 61.490 148.980 61.780 149.025 ;
        RECT 60.185 148.840 61.780 148.980 ;
        RECT 58.270 148.795 58.560 148.840 ;
        RECT 58.715 148.780 59.035 148.840 ;
        RECT 61.490 148.795 61.780 148.840 ;
        RECT 61.950 148.795 62.240 149.025 ;
        RECT 62.855 148.980 63.175 149.040 ;
        RECT 63.330 148.980 63.620 149.025 ;
        RECT 62.855 148.840 63.620 148.980 ;
        RECT 22.465 148.500 27.665 148.640 ;
        RECT 28.355 148.440 28.675 148.700 ;
        RECT 30.670 148.640 30.960 148.685 ;
        RECT 31.575 148.640 31.895 148.700 ;
        RECT 40.405 148.640 40.545 148.780 ;
        RECT 47.675 148.640 47.995 148.700 ;
        RECT 53.210 148.640 53.500 148.685 ;
        RECT 57.335 148.640 57.655 148.700 ;
        RECT 30.670 148.500 40.545 148.640 ;
        RECT 45.925 148.500 49.285 148.640 ;
        RECT 30.670 148.455 30.960 148.500 ;
        RECT 31.575 148.440 31.895 148.500 ;
        RECT 22.835 148.100 23.155 148.360 ;
        RECT 26.055 148.300 26.375 148.360 ;
        RECT 28.445 148.300 28.585 148.440 ;
        RECT 26.055 148.160 28.585 148.300 ;
        RECT 31.135 148.300 31.425 148.345 ;
        RECT 32.995 148.300 33.285 148.345 ;
        RECT 35.775 148.300 36.065 148.345 ;
        RECT 31.135 148.160 36.065 148.300 ;
        RECT 26.055 148.100 26.375 148.160 ;
        RECT 31.135 148.115 31.425 148.160 ;
        RECT 32.995 148.115 33.285 148.160 ;
        RECT 35.775 148.115 36.065 148.160 ;
        RECT 38.935 148.300 39.255 148.360 ;
        RECT 39.640 148.300 39.930 148.345 ;
        RECT 38.935 148.160 39.930 148.300 ;
        RECT 38.935 148.100 39.255 148.160 ;
        RECT 39.640 148.115 39.930 148.160 ;
        RECT 43.535 148.300 43.855 148.360 ;
        RECT 44.010 148.300 44.300 148.345 ;
        RECT 43.535 148.160 44.300 148.300 ;
        RECT 43.535 148.100 43.855 148.160 ;
        RECT 44.010 148.115 44.300 148.160 ;
        RECT 45.375 148.300 45.695 148.360 ;
        RECT 45.925 148.300 46.065 148.500 ;
        RECT 47.675 148.440 47.995 148.500 ;
        RECT 45.375 148.160 46.065 148.300 ;
        RECT 45.375 148.100 45.695 148.160 ;
        RECT 48.595 148.100 48.915 148.360 ;
        RECT 49.145 148.300 49.285 148.500 ;
        RECT 53.210 148.500 57.655 148.640 ;
        RECT 53.210 148.455 53.500 148.500 ;
        RECT 57.335 148.440 57.655 148.500 ;
        RECT 60.095 148.640 60.415 148.700 ;
        RECT 62.025 148.640 62.165 148.795 ;
        RECT 62.855 148.780 63.175 148.840 ;
        RECT 63.330 148.795 63.620 148.840 ;
        RECT 64.235 148.980 64.555 149.040 ;
        RECT 65.170 148.980 65.460 149.025 ;
        RECT 64.235 148.840 65.460 148.980 ;
        RECT 64.235 148.780 64.555 148.840 ;
        RECT 65.170 148.795 65.460 148.840 ;
        RECT 66.075 148.780 66.395 149.040 ;
        RECT 66.535 148.780 66.855 149.040 ;
        RECT 66.995 148.780 67.315 149.040 ;
        RECT 60.095 148.500 62.165 148.640 ;
        RECT 69.385 148.640 69.525 149.180 ;
        RECT 69.845 149.180 73.205 149.320 ;
        RECT 69.845 149.025 69.985 149.180 ;
        RECT 73.065 149.040 73.205 149.180 ;
        RECT 73.895 149.180 84.335 149.320 ;
        RECT 73.895 149.120 74.215 149.180 ;
        RECT 82.650 149.135 82.940 149.180 ;
        RECT 84.015 149.120 84.335 149.180 ;
        RECT 69.770 148.795 70.060 149.025 ;
        RECT 70.230 148.795 70.520 149.025 ;
        RECT 70.675 148.980 70.995 149.040 ;
        RECT 71.595 148.980 71.915 149.040 ;
        RECT 70.675 148.840 71.915 148.980 ;
        RECT 70.305 148.640 70.445 148.795 ;
        RECT 70.675 148.780 70.995 148.840 ;
        RECT 71.595 148.780 71.915 148.840 ;
        RECT 72.975 148.780 73.295 149.040 ;
        RECT 78.970 148.980 79.260 149.025 ;
        RECT 79.430 148.980 79.720 149.025 ;
        RECT 83.095 148.980 83.415 149.040 ;
        RECT 78.970 148.840 83.415 148.980 ;
        RECT 84.565 148.980 84.705 149.475 ;
        RECT 84.935 149.460 85.255 149.720 ;
        RECT 90.915 149.660 91.235 149.720 ;
        RECT 89.625 149.520 91.235 149.660 ;
        RECT 85.870 148.980 86.160 149.025 ;
        RECT 89.625 148.980 89.765 149.520 ;
        RECT 90.915 149.460 91.235 149.520 ;
        RECT 92.295 149.660 92.615 149.720 ;
        RECT 94.135 149.660 94.455 149.720 ;
        RECT 92.295 149.520 93.905 149.660 ;
        RECT 92.295 149.460 92.615 149.520 ;
        RECT 89.995 149.320 90.315 149.380 ;
        RECT 89.995 149.180 92.525 149.320 ;
        RECT 89.995 149.120 90.315 149.180 ;
        RECT 92.385 149.025 92.525 149.180 ;
        RECT 90.470 148.980 90.760 149.025 ;
        RECT 84.565 148.840 86.160 148.980 ;
        RECT 78.970 148.795 79.260 148.840 ;
        RECT 79.430 148.795 79.720 148.840 ;
        RECT 83.095 148.780 83.415 148.840 ;
        RECT 85.870 148.795 86.160 148.840 ;
        RECT 88.705 148.840 90.760 148.980 ;
        RECT 72.515 148.640 72.835 148.700 ;
        RECT 69.385 148.500 72.835 148.640 ;
        RECT 60.095 148.440 60.415 148.500 ;
        RECT 72.515 148.440 72.835 148.500 ;
        RECT 78.125 148.500 81.485 148.640 ;
        RECT 55.970 148.300 56.260 148.345 ;
        RECT 61.935 148.300 62.255 148.360 ;
        RECT 49.145 148.160 55.725 148.300 ;
        RECT 55.585 147.960 55.725 148.160 ;
        RECT 55.970 148.160 62.255 148.300 ;
        RECT 55.970 148.115 56.260 148.160 ;
        RECT 61.935 148.100 62.255 148.160 ;
        RECT 62.395 148.100 62.715 148.360 ;
        RECT 67.455 148.300 67.775 148.360 ;
        RECT 70.675 148.300 70.995 148.360 ;
        RECT 71.150 148.300 71.440 148.345 ;
        RECT 78.125 148.300 78.265 148.500 ;
        RECT 63.405 148.160 70.445 148.300 ;
        RECT 63.405 147.960 63.545 148.160 ;
        RECT 67.455 148.100 67.775 148.160 ;
        RECT 55.585 147.820 63.545 147.960 ;
        RECT 67.930 147.960 68.220 148.005 ;
        RECT 68.375 147.960 68.695 148.020 ;
        RECT 67.930 147.820 68.695 147.960 ;
        RECT 67.930 147.775 68.220 147.820 ;
        RECT 68.375 147.760 68.695 147.820 ;
        RECT 68.835 147.760 69.155 148.020 ;
        RECT 70.305 147.960 70.445 148.160 ;
        RECT 70.675 148.160 71.440 148.300 ;
        RECT 70.675 148.100 70.995 148.160 ;
        RECT 71.150 148.115 71.440 148.160 ;
        RECT 71.685 148.160 78.265 148.300 ;
        RECT 78.510 148.300 78.800 148.345 ;
        RECT 78.955 148.300 79.275 148.360 ;
        RECT 78.510 148.160 79.275 148.300 ;
        RECT 81.345 148.300 81.485 148.500 ;
        RECT 81.715 148.440 82.035 148.700 ;
        RECT 88.705 148.360 88.845 148.840 ;
        RECT 90.470 148.795 90.760 148.840 ;
        RECT 90.930 148.795 91.220 149.025 ;
        RECT 91.390 148.795 91.680 149.025 ;
        RECT 92.310 148.980 92.600 149.025 ;
        RECT 92.755 148.980 93.075 149.040 ;
        RECT 93.765 149.025 93.905 149.520 ;
        RECT 94.135 149.520 100.345 149.660 ;
        RECT 94.135 149.460 94.455 149.520 ;
        RECT 92.310 148.840 93.075 148.980 ;
        RECT 92.310 148.795 92.600 148.840 ;
        RECT 88.615 148.300 88.935 148.360 ;
        RECT 81.345 148.160 88.935 148.300 ;
        RECT 71.685 147.960 71.825 148.160 ;
        RECT 78.510 148.115 78.800 148.160 ;
        RECT 78.955 148.100 79.275 148.160 ;
        RECT 88.615 148.100 88.935 148.160 ;
        RECT 90.455 148.300 90.775 148.360 ;
        RECT 91.005 148.300 91.145 148.795 ;
        RECT 91.465 148.640 91.605 148.795 ;
        RECT 92.755 148.780 93.075 148.840 ;
        RECT 93.690 148.795 93.980 149.025 ;
        RECT 94.135 148.780 94.455 149.040 ;
        RECT 94.595 148.780 94.915 149.040 ;
        RECT 96.450 148.980 96.740 149.025 ;
        RECT 97.355 148.980 97.675 149.040 ;
        RECT 96.450 148.840 97.675 148.980 ;
        RECT 96.450 148.795 96.740 148.840 ;
        RECT 97.355 148.780 97.675 148.840 ;
        RECT 97.815 148.780 98.135 149.040 ;
        RECT 100.205 149.025 100.345 149.520 ;
        RECT 100.590 149.320 100.880 149.365 ;
        RECT 103.745 149.320 104.035 149.365 ;
        RECT 107.005 149.320 107.295 149.365 ;
        RECT 100.590 149.180 107.295 149.320 ;
        RECT 100.590 149.135 100.880 149.180 ;
        RECT 103.745 149.135 104.035 149.180 ;
        RECT 107.005 149.135 107.295 149.180 ;
        RECT 107.925 149.320 108.215 149.365 ;
        RECT 109.785 149.320 110.075 149.365 ;
        RECT 107.925 149.180 110.075 149.320 ;
        RECT 107.925 149.135 108.215 149.180 ;
        RECT 109.785 149.135 110.075 149.180 ;
        RECT 100.130 148.980 100.420 149.025 ;
        RECT 101.955 148.980 102.275 149.040 ;
        RECT 104.715 148.980 105.035 149.040 ;
        RECT 100.130 148.840 105.035 148.980 ;
        RECT 100.130 148.795 100.420 148.840 ;
        RECT 101.955 148.780 102.275 148.840 ;
        RECT 104.715 148.780 105.035 148.840 ;
        RECT 105.605 148.980 105.895 149.025 ;
        RECT 107.925 148.980 108.140 149.135 ;
        RECT 105.605 148.840 108.140 148.980 ;
        RECT 110.235 148.980 110.555 149.040 ;
        RECT 110.710 148.980 111.000 149.025 ;
        RECT 110.235 148.840 111.000 148.980 ;
        RECT 105.605 148.795 105.895 148.840 ;
        RECT 110.235 148.780 110.555 148.840 ;
        RECT 110.710 148.795 111.000 148.840 ;
        RECT 93.215 148.640 93.535 148.700 ;
        RECT 91.465 148.500 93.535 148.640 ;
        RECT 93.215 148.440 93.535 148.500 ;
        RECT 96.895 148.440 97.215 148.700 ;
        RECT 108.870 148.640 109.160 148.685 ;
        RECT 109.315 148.640 109.635 148.700 ;
        RECT 108.870 148.500 109.635 148.640 ;
        RECT 108.870 148.455 109.160 148.500 ;
        RECT 109.315 148.440 109.635 148.500 ;
        RECT 94.135 148.300 94.455 148.360 ;
        RECT 90.455 148.160 94.455 148.300 ;
        RECT 90.455 148.100 90.775 148.160 ;
        RECT 94.135 148.100 94.455 148.160 ;
        RECT 94.595 148.300 94.915 148.360 ;
        RECT 95.990 148.300 96.280 148.345 ;
        RECT 94.595 148.160 96.280 148.300 ;
        RECT 94.595 148.100 94.915 148.160 ;
        RECT 95.990 148.115 96.280 148.160 ;
        RECT 98.750 148.300 99.040 148.345 ;
        RECT 99.655 148.300 99.975 148.360 ;
        RECT 98.750 148.160 99.975 148.300 ;
        RECT 98.750 148.115 99.040 148.160 ;
        RECT 99.655 148.100 99.975 148.160 ;
        RECT 105.605 148.300 105.895 148.345 ;
        RECT 108.385 148.300 108.675 148.345 ;
        RECT 110.245 148.300 110.535 148.345 ;
        RECT 105.605 148.160 110.535 148.300 ;
        RECT 105.605 148.115 105.895 148.160 ;
        RECT 108.385 148.115 108.675 148.160 ;
        RECT 110.245 148.115 110.535 148.160 ;
        RECT 70.305 147.820 71.825 147.960 ;
        RECT 89.090 147.960 89.380 148.005 ;
        RECT 89.995 147.960 90.315 148.020 ;
        RECT 89.090 147.820 90.315 147.960 ;
        RECT 89.090 147.775 89.380 147.820 ;
        RECT 89.995 147.760 90.315 147.820 ;
        RECT 97.815 147.760 98.135 148.020 ;
        RECT 101.740 147.960 102.030 148.005 ;
        RECT 103.795 147.960 104.115 148.020 ;
        RECT 101.740 147.820 104.115 147.960 ;
        RECT 101.740 147.775 102.030 147.820 ;
        RECT 103.795 147.760 104.115 147.820 ;
        RECT 18.165 147.140 112.465 147.620 ;
        RECT 32.955 146.940 33.275 147.000 ;
        RECT 33.430 146.940 33.720 146.985 ;
        RECT 70.675 146.940 70.995 147.000 ;
        RECT 89.535 146.940 89.855 147.000 ;
        RECT 32.955 146.800 33.720 146.940 ;
        RECT 32.955 146.740 33.275 146.800 ;
        RECT 33.430 146.755 33.720 146.800 ;
        RECT 49.605 146.800 89.855 146.940 ;
        RECT 23.870 146.600 24.160 146.645 ;
        RECT 26.990 146.600 27.280 146.645 ;
        RECT 28.880 146.600 29.170 146.645 ;
        RECT 23.870 146.460 29.170 146.600 ;
        RECT 23.870 146.415 24.160 146.460 ;
        RECT 26.990 146.415 27.280 146.460 ;
        RECT 28.880 146.415 29.170 146.460 ;
        RECT 32.510 146.600 32.800 146.645 ;
        RECT 35.255 146.600 35.575 146.660 ;
        RECT 32.510 146.460 35.575 146.600 ;
        RECT 32.510 146.415 32.800 146.460 ;
        RECT 35.255 146.400 35.575 146.460 ;
        RECT 37.095 146.600 37.415 146.660 ;
        RECT 37.095 146.460 43.765 146.600 ;
        RECT 37.095 146.400 37.415 146.460 ;
        RECT 29.750 146.260 30.040 146.305 ;
        RECT 31.575 146.260 31.895 146.320 ;
        RECT 29.750 146.120 31.895 146.260 ;
        RECT 29.750 146.075 30.040 146.120 ;
        RECT 31.575 146.060 31.895 146.120 ;
        RECT 36.635 146.260 36.955 146.320 ;
        RECT 38.030 146.260 38.320 146.305 ;
        RECT 36.635 146.120 38.320 146.260 ;
        RECT 36.635 146.060 36.955 146.120 ;
        RECT 38.030 146.075 38.320 146.120 ;
        RECT 22.835 145.940 23.155 145.980 ;
        RECT 22.790 145.720 23.155 145.940 ;
        RECT 23.870 145.920 24.160 145.965 ;
        RECT 27.450 145.920 27.740 145.965 ;
        RECT 29.285 145.920 29.575 145.965 ;
        RECT 23.870 145.780 29.575 145.920 ;
        RECT 23.870 145.735 24.160 145.780 ;
        RECT 27.450 145.735 27.740 145.780 ;
        RECT 29.285 145.735 29.575 145.780 ;
        RECT 31.115 145.720 31.435 145.980 ;
        RECT 32.035 145.720 32.355 145.980 ;
        RECT 34.335 145.720 34.655 145.980 ;
        RECT 37.110 145.920 37.400 145.965 ;
        RECT 37.555 145.920 37.875 145.980 ;
        RECT 37.110 145.780 37.875 145.920 ;
        RECT 37.110 145.735 37.400 145.780 ;
        RECT 37.555 145.720 37.875 145.780 ;
        RECT 39.395 145.920 39.715 145.980 ;
        RECT 42.630 145.920 42.920 145.965 ;
        RECT 39.395 145.780 42.920 145.920 ;
        RECT 39.395 145.720 39.715 145.780 ;
        RECT 42.630 145.735 42.920 145.780 ;
        RECT 43.075 145.720 43.395 145.980 ;
        RECT 43.625 145.965 43.765 146.460 ;
        RECT 43.995 146.260 44.315 146.320 ;
        RECT 47.675 146.260 47.995 146.320 ;
        RECT 49.070 146.260 49.360 146.305 ;
        RECT 43.995 146.120 47.445 146.260 ;
        RECT 43.995 146.060 44.315 146.120 ;
        RECT 43.550 145.735 43.840 145.965 ;
        RECT 44.470 145.735 44.760 145.965 ;
        RECT 45.375 145.920 45.695 145.980 ;
        RECT 46.310 145.920 46.600 145.965 ;
        RECT 45.375 145.780 46.600 145.920 ;
        RECT 22.790 145.625 23.080 145.720 ;
        RECT 22.490 145.580 23.080 145.625 ;
        RECT 25.730 145.580 26.380 145.625 ;
        RECT 22.490 145.440 26.380 145.580 ;
        RECT 22.490 145.395 22.780 145.440 ;
        RECT 25.730 145.395 26.380 145.440 ;
        RECT 28.370 145.395 28.660 145.625 ;
        RECT 41.250 145.580 41.540 145.625 ;
        RECT 43.995 145.580 44.315 145.640 ;
        RECT 41.250 145.440 44.315 145.580 ;
        RECT 44.545 145.580 44.685 145.735 ;
        RECT 45.375 145.720 45.695 145.780 ;
        RECT 46.310 145.735 46.600 145.780 ;
        RECT 46.755 145.720 47.075 145.980 ;
        RECT 47.305 145.965 47.445 146.120 ;
        RECT 47.675 146.120 49.360 146.260 ;
        RECT 47.675 146.060 47.995 146.120 ;
        RECT 49.070 146.075 49.360 146.120 ;
        RECT 47.230 145.735 47.520 145.965 ;
        RECT 48.135 145.920 48.455 145.980 ;
        RECT 49.605 145.920 49.745 146.800 ;
        RECT 70.675 146.740 70.995 146.800 ;
        RECT 54.575 146.600 54.895 146.660 ;
        RECT 51.445 146.460 54.895 146.600 ;
        RECT 48.135 145.780 49.745 145.920 ;
        RECT 49.975 145.920 50.295 145.980 ;
        RECT 50.450 145.920 50.740 145.965 ;
        RECT 49.975 145.780 50.740 145.920 ;
        RECT 48.135 145.720 48.455 145.780 ;
        RECT 49.975 145.720 50.295 145.780 ;
        RECT 50.450 145.735 50.740 145.780 ;
        RECT 50.895 145.720 51.215 145.980 ;
        RECT 51.445 145.965 51.585 146.460 ;
        RECT 54.575 146.400 54.895 146.460 ;
        RECT 55.970 146.600 56.260 146.645 ;
        RECT 64.235 146.600 64.555 146.660 ;
        RECT 55.970 146.460 64.555 146.600 ;
        RECT 55.970 146.415 56.260 146.460 ;
        RECT 64.235 146.400 64.555 146.460 ;
        RECT 65.125 146.600 65.415 146.645 ;
        RECT 67.905 146.600 68.195 146.645 ;
        RECT 69.765 146.600 70.055 146.645 ;
        RECT 65.125 146.460 70.055 146.600 ;
        RECT 65.125 146.415 65.415 146.460 ;
        RECT 67.905 146.415 68.195 146.460 ;
        RECT 69.765 146.415 70.055 146.460 ;
        RECT 79.990 146.600 80.280 146.645 ;
        RECT 83.110 146.600 83.400 146.645 ;
        RECT 85.000 146.600 85.290 146.645 ;
        RECT 79.990 146.460 85.290 146.600 ;
        RECT 79.990 146.415 80.280 146.460 ;
        RECT 83.110 146.415 83.400 146.460 ;
        RECT 85.000 146.415 85.290 146.460 ;
        RECT 56.875 146.060 57.195 146.320 ;
        RECT 68.375 146.060 68.695 146.320 ;
        RECT 70.215 146.060 70.535 146.320 ;
        RECT 85.855 146.060 86.175 146.320 ;
        RECT 51.370 145.735 51.660 145.965 ;
        RECT 51.815 145.920 52.135 145.980 ;
        RECT 52.290 145.920 52.580 145.965 ;
        RECT 51.815 145.780 52.580 145.920 ;
        RECT 51.815 145.720 52.135 145.780 ;
        RECT 52.290 145.735 52.580 145.780 ;
        RECT 52.735 145.920 53.055 145.980 ;
        RECT 58.270 145.920 58.560 145.965 ;
        RECT 61.260 145.920 61.550 145.965 ;
        RECT 52.735 145.780 61.550 145.920 ;
        RECT 52.735 145.720 53.055 145.780 ;
        RECT 58.270 145.735 58.560 145.780 ;
        RECT 61.260 145.735 61.550 145.780 ;
        RECT 65.125 145.920 65.415 145.965 ;
        RECT 78.955 145.940 79.275 145.980 ;
        RECT 65.125 145.780 67.660 145.920 ;
        RECT 65.125 145.735 65.415 145.780 ;
        RECT 49.515 145.580 49.835 145.640 ;
        RECT 60.555 145.580 60.875 145.640 ;
        RECT 62.395 145.580 62.715 145.640 ;
        RECT 67.445 145.625 67.660 145.780 ;
        RECT 78.910 145.720 79.275 145.940 ;
        RECT 79.990 145.920 80.280 145.965 ;
        RECT 83.570 145.920 83.860 145.965 ;
        RECT 85.405 145.920 85.695 145.965 ;
        RECT 79.990 145.780 85.695 145.920 ;
        RECT 86.405 145.920 86.545 146.800 ;
        RECT 89.535 146.740 89.855 146.800 ;
        RECT 95.990 146.940 96.280 146.985 ;
        RECT 96.895 146.940 97.215 147.000 ;
        RECT 95.990 146.800 97.215 146.940 ;
        RECT 95.990 146.755 96.280 146.800 ;
        RECT 96.895 146.740 97.215 146.800 ;
        RECT 97.355 146.940 97.675 147.000 ;
        RECT 97.830 146.940 98.120 146.985 ;
        RECT 97.355 146.800 98.120 146.940 ;
        RECT 97.355 146.740 97.675 146.800 ;
        RECT 97.830 146.755 98.120 146.800 ;
        RECT 106.095 146.740 106.415 147.000 ;
        RECT 107.950 146.940 108.240 146.985 ;
        RECT 108.855 146.940 109.175 147.000 ;
        RECT 107.950 146.800 109.175 146.940 ;
        RECT 107.950 146.755 108.240 146.800 ;
        RECT 108.855 146.740 109.175 146.800 ;
        RECT 109.315 146.740 109.635 147.000 ;
        RECT 93.215 146.600 93.535 146.660 ;
        RECT 103.335 146.600 103.655 146.660 ;
        RECT 93.215 146.460 101.725 146.600 ;
        RECT 93.215 146.400 93.535 146.460 ;
        RECT 86.775 146.260 87.095 146.320 ;
        RECT 90.455 146.260 90.775 146.320 ;
        RECT 86.775 146.120 88.385 146.260 ;
        RECT 86.775 146.060 87.095 146.120 ;
        RECT 88.245 145.965 88.385 146.120 ;
        RECT 88.705 146.120 90.775 146.260 ;
        RECT 88.705 145.965 88.845 146.120 ;
        RECT 90.455 146.060 90.775 146.120 ;
        RECT 91.835 146.260 92.155 146.320 ;
        RECT 91.835 146.120 93.905 146.260 ;
        RECT 91.835 146.060 92.155 146.120 ;
        RECT 87.250 145.920 87.540 145.965 ;
        RECT 86.405 145.780 87.540 145.920 ;
        RECT 79.990 145.735 80.280 145.780 ;
        RECT 83.570 145.735 83.860 145.780 ;
        RECT 85.405 145.735 85.695 145.780 ;
        RECT 87.250 145.735 87.540 145.780 ;
        RECT 88.170 145.735 88.460 145.965 ;
        RECT 88.630 145.735 88.920 145.965 ;
        RECT 78.910 145.625 79.200 145.720 ;
        RECT 63.265 145.580 63.555 145.625 ;
        RECT 66.525 145.580 66.815 145.625 ;
        RECT 44.545 145.440 48.825 145.580 ;
        RECT 41.250 145.395 41.540 145.440 ;
        RECT 21.010 145.240 21.300 145.285 ;
        RECT 26.975 145.240 27.295 145.300 ;
        RECT 21.010 145.100 27.295 145.240 ;
        RECT 28.445 145.240 28.585 145.395 ;
        RECT 43.995 145.380 44.315 145.440 ;
        RECT 30.210 145.240 30.500 145.285 ;
        RECT 28.445 145.100 30.500 145.240 ;
        RECT 21.010 145.055 21.300 145.100 ;
        RECT 26.975 145.040 27.295 145.100 ;
        RECT 30.210 145.055 30.500 145.100 ;
        RECT 35.270 145.240 35.560 145.285 ;
        RECT 36.175 145.240 36.495 145.300 ;
        RECT 35.270 145.100 36.495 145.240 ;
        RECT 35.270 145.055 35.560 145.100 ;
        RECT 36.175 145.040 36.495 145.100 ;
        RECT 37.555 145.040 37.875 145.300 ;
        RECT 43.075 145.240 43.395 145.300 ;
        RECT 44.930 145.240 45.220 145.285 ;
        RECT 43.075 145.100 45.220 145.240 ;
        RECT 48.685 145.240 48.825 145.440 ;
        RECT 49.515 145.440 62.165 145.580 ;
        RECT 49.515 145.380 49.835 145.440 ;
        RECT 60.555 145.380 60.875 145.440 ;
        RECT 53.195 145.240 53.515 145.300 ;
        RECT 55.495 145.240 55.815 145.300 ;
        RECT 48.685 145.100 55.815 145.240 ;
        RECT 43.075 145.040 43.395 145.100 ;
        RECT 44.930 145.055 45.220 145.100 ;
        RECT 53.195 145.040 53.515 145.100 ;
        RECT 55.495 145.040 55.815 145.100 ;
        RECT 57.795 145.040 58.115 145.300 ;
        RECT 60.110 145.240 60.400 145.285 ;
        RECT 61.015 145.240 61.335 145.300 ;
        RECT 60.110 145.100 61.335 145.240 ;
        RECT 62.025 145.240 62.165 145.440 ;
        RECT 62.395 145.440 66.815 145.580 ;
        RECT 62.395 145.380 62.715 145.440 ;
        RECT 63.265 145.395 63.555 145.440 ;
        RECT 66.525 145.395 66.815 145.440 ;
        RECT 67.445 145.580 67.735 145.625 ;
        RECT 69.305 145.580 69.595 145.625 ;
        RECT 78.610 145.580 79.200 145.625 ;
        RECT 81.850 145.580 82.500 145.625 ;
        RECT 67.445 145.440 69.595 145.580 ;
        RECT 67.445 145.395 67.735 145.440 ;
        RECT 69.305 145.395 69.595 145.440 ;
        RECT 76.745 145.440 78.265 145.580 ;
        RECT 76.745 145.240 76.885 145.440 ;
        RECT 62.025 145.100 76.885 145.240 ;
        RECT 60.110 145.055 60.400 145.100 ;
        RECT 61.015 145.040 61.335 145.100 ;
        RECT 77.115 145.040 77.435 145.300 ;
        RECT 78.125 145.240 78.265 145.440 ;
        RECT 78.610 145.440 82.500 145.580 ;
        RECT 78.610 145.395 78.900 145.440 ;
        RECT 81.850 145.395 82.500 145.440 ;
        RECT 84.475 145.380 84.795 145.640 ;
        RECT 88.705 145.240 88.845 145.735 ;
        RECT 89.075 145.720 89.395 145.980 ;
        RECT 89.535 145.920 89.855 145.980 ;
        RECT 93.765 145.965 93.905 146.120 ;
        RECT 92.770 145.920 93.060 145.965 ;
        RECT 89.535 145.780 93.060 145.920 ;
        RECT 89.535 145.720 89.855 145.780 ;
        RECT 92.770 145.735 93.060 145.780 ;
        RECT 93.690 145.735 93.980 145.965 ;
        RECT 94.135 145.720 94.455 145.980 ;
        RECT 94.610 145.735 94.900 145.965 ;
        RECT 97.355 145.920 97.675 145.980 ;
        RECT 99.210 145.920 99.500 145.965 ;
        RECT 97.355 145.780 99.500 145.920 ;
        RECT 89.165 145.580 89.305 145.720 ;
        RECT 94.685 145.580 94.825 145.735 ;
        RECT 97.355 145.720 97.675 145.780 ;
        RECT 99.210 145.735 99.500 145.780 ;
        RECT 99.670 145.735 99.960 145.965 ;
        RECT 100.130 145.735 100.420 145.965 ;
        RECT 100.575 145.920 100.895 145.980 ;
        RECT 101.050 145.920 101.340 145.965 ;
        RECT 100.575 145.780 101.340 145.920 ;
        RECT 101.585 145.920 101.725 146.460 ;
        RECT 102.505 146.460 103.655 146.600 ;
        RECT 102.505 146.305 102.645 146.460 ;
        RECT 103.335 146.400 103.655 146.460 ;
        RECT 105.190 146.415 105.480 146.645 ;
        RECT 102.430 146.075 102.720 146.305 ;
        RECT 105.265 146.260 105.405 146.415 ;
        RECT 105.265 146.120 107.245 146.260 ;
        RECT 103.350 145.920 103.640 145.965 ;
        RECT 101.585 145.780 103.640 145.920 ;
        RECT 98.735 145.580 99.055 145.640 ;
        RECT 99.745 145.580 99.885 145.735 ;
        RECT 89.165 145.440 94.825 145.580 ;
        RECT 96.985 145.440 99.885 145.580 ;
        RECT 100.205 145.580 100.345 145.735 ;
        RECT 100.575 145.720 100.895 145.780 ;
        RECT 101.050 145.735 101.340 145.780 ;
        RECT 103.350 145.735 103.640 145.780 ;
        RECT 104.715 145.920 105.035 145.980 ;
        RECT 106.555 145.920 106.875 145.980 ;
        RECT 107.105 145.965 107.245 146.120 ;
        RECT 104.715 145.780 106.875 145.920 ;
        RECT 104.715 145.720 105.035 145.780 ;
        RECT 106.555 145.720 106.875 145.780 ;
        RECT 107.030 145.735 107.320 145.965 ;
        RECT 108.395 145.720 108.715 145.980 ;
        RECT 103.795 145.580 104.115 145.640 ;
        RECT 100.205 145.440 104.115 145.580 ;
        RECT 96.985 145.300 97.125 145.440 ;
        RECT 98.735 145.380 99.055 145.440 ;
        RECT 103.795 145.380 104.115 145.440 ;
        RECT 78.125 145.100 88.845 145.240 ;
        RECT 90.455 145.040 90.775 145.300 ;
        RECT 96.895 145.040 97.215 145.300 ;
        RECT 102.890 145.240 103.180 145.285 ;
        RECT 104.255 145.240 104.575 145.300 ;
        RECT 102.890 145.100 104.575 145.240 ;
        RECT 102.890 145.055 103.180 145.100 ;
        RECT 104.255 145.040 104.575 145.100 ;
        RECT 17.370 144.420 112.465 144.900 ;
        RECT 28.830 144.220 29.120 144.265 ;
        RECT 31.115 144.220 31.435 144.280 ;
        RECT 28.830 144.080 31.435 144.220 ;
        RECT 28.830 144.035 29.120 144.080 ;
        RECT 31.115 144.020 31.435 144.080 ;
        RECT 31.590 144.220 31.880 144.265 ;
        RECT 37.555 144.220 37.875 144.280 ;
        RECT 31.590 144.080 37.875 144.220 ;
        RECT 31.590 144.035 31.880 144.080 ;
        RECT 37.555 144.020 37.875 144.080 ;
        RECT 38.475 144.220 38.795 144.280 ;
        RECT 41.250 144.220 41.540 144.265 ;
        RECT 44.455 144.220 44.775 144.280 ;
        RECT 38.475 144.080 41.540 144.220 ;
        RECT 38.475 144.020 38.795 144.080 ;
        RECT 41.250 144.035 41.540 144.080 ;
        RECT 42.245 144.080 44.775 144.220 ;
        RECT 26.515 143.880 26.835 143.940 ;
        RECT 26.990 143.880 27.280 143.925 ;
        RECT 26.515 143.740 27.280 143.880 ;
        RECT 26.515 143.680 26.835 143.740 ;
        RECT 26.990 143.695 27.280 143.740 ;
        RECT 30.670 143.880 30.960 143.925 ;
        RECT 33.070 143.880 33.360 143.925 ;
        RECT 36.310 143.880 36.960 143.925 ;
        RECT 30.670 143.740 36.960 143.880 ;
        RECT 30.670 143.695 30.960 143.740 ;
        RECT 33.070 143.695 33.660 143.740 ;
        RECT 36.310 143.695 36.960 143.740 ;
        RECT 39.395 143.880 39.715 143.940 ;
        RECT 41.695 143.880 42.015 143.940 ;
        RECT 39.395 143.740 42.015 143.880 ;
        RECT 23.755 143.540 24.075 143.600 ;
        RECT 30.210 143.540 30.500 143.585 ;
        RECT 31.115 143.540 31.435 143.600 ;
        RECT 23.755 143.400 29.965 143.540 ;
        RECT 23.755 143.340 24.075 143.400 ;
        RECT 26.055 143.000 26.375 143.260 ;
        RECT 26.530 143.200 26.820 143.245 ;
        RECT 26.975 143.200 27.295 143.260 ;
        RECT 26.530 143.060 27.295 143.200 ;
        RECT 29.825 143.200 29.965 143.400 ;
        RECT 30.210 143.400 31.435 143.540 ;
        RECT 30.210 143.355 30.500 143.400 ;
        RECT 31.115 143.340 31.435 143.400 ;
        RECT 33.370 143.380 33.660 143.695 ;
        RECT 39.395 143.680 39.715 143.740 ;
        RECT 41.695 143.680 42.015 143.740 ;
        RECT 34.450 143.540 34.740 143.585 ;
        RECT 38.030 143.540 38.320 143.585 ;
        RECT 39.865 143.540 40.155 143.585 ;
        RECT 34.450 143.400 40.155 143.540 ;
        RECT 34.450 143.355 34.740 143.400 ;
        RECT 38.030 143.355 38.320 143.400 ;
        RECT 39.865 143.355 40.155 143.400 ;
        RECT 40.315 143.340 40.635 143.600 ;
        RECT 42.245 143.585 42.385 144.080 ;
        RECT 44.455 144.020 44.775 144.080 ;
        RECT 46.755 144.220 47.075 144.280 ;
        RECT 49.515 144.220 49.835 144.280 ;
        RECT 46.755 144.080 49.835 144.220 ;
        RECT 46.755 144.020 47.075 144.080 ;
        RECT 49.515 144.020 49.835 144.080 ;
        RECT 50.435 144.220 50.755 144.280 ;
        RECT 56.875 144.220 57.195 144.280 ;
        RECT 67.470 144.220 67.760 144.265 ;
        RECT 50.435 144.080 54.345 144.220 ;
        RECT 50.435 144.020 50.755 144.080 ;
        RECT 43.550 143.880 43.840 143.925 ;
        RECT 48.610 143.880 48.900 143.925 ;
        RECT 52.735 143.880 53.055 143.940 ;
        RECT 43.550 143.740 48.900 143.880 ;
        RECT 43.550 143.695 43.840 143.740 ;
        RECT 48.610 143.695 48.900 143.740 ;
        RECT 50.985 143.740 53.055 143.880 ;
        RECT 42.170 143.355 42.460 143.585 ;
        RECT 42.630 143.540 42.920 143.585 ;
        RECT 43.075 143.540 43.395 143.600 ;
        RECT 42.630 143.400 43.395 143.540 ;
        RECT 42.630 143.355 42.920 143.400 ;
        RECT 43.075 143.340 43.395 143.400 ;
        RECT 44.010 143.540 44.300 143.585 ;
        RECT 44.455 143.540 44.775 143.600 ;
        RECT 44.010 143.400 44.775 143.540 ;
        RECT 44.010 143.355 44.300 143.400 ;
        RECT 44.455 143.340 44.775 143.400 ;
        RECT 44.930 143.355 45.220 143.585 ;
        RECT 45.390 143.355 45.680 143.585 ;
        RECT 38.475 143.200 38.795 143.260 ;
        RECT 29.825 143.060 38.795 143.200 ;
        RECT 26.530 143.015 26.820 143.060 ;
        RECT 26.605 142.520 26.745 143.015 ;
        RECT 26.975 143.000 27.295 143.060 ;
        RECT 38.475 143.000 38.795 143.060 ;
        RECT 38.935 143.000 39.255 143.260 ;
        RECT 41.235 143.200 41.555 143.260 ;
        RECT 43.535 143.200 43.855 143.260 ;
        RECT 41.235 143.060 43.855 143.200 ;
        RECT 41.235 143.000 41.555 143.060 ;
        RECT 43.535 143.000 43.855 143.060 ;
        RECT 34.450 142.860 34.740 142.905 ;
        RECT 37.570 142.860 37.860 142.905 ;
        RECT 39.460 142.860 39.750 142.905 ;
        RECT 45.005 142.860 45.145 143.355 ;
        RECT 45.465 143.200 45.605 143.355 ;
        RECT 45.835 143.340 46.155 143.600 ;
        RECT 46.755 143.340 47.075 143.600 ;
        RECT 49.975 143.340 50.295 143.600 ;
        RECT 50.435 143.340 50.755 143.600 ;
        RECT 50.985 143.585 51.125 143.740 ;
        RECT 52.735 143.680 53.055 143.740 ;
        RECT 50.910 143.355 51.200 143.585 ;
        RECT 51.830 143.540 52.120 143.585 ;
        RECT 53.195 143.540 53.515 143.600 ;
        RECT 54.205 143.585 54.345 144.080 ;
        RECT 56.875 144.080 67.760 144.220 ;
        RECT 56.875 144.020 57.195 144.080 ;
        RECT 67.470 144.035 67.760 144.080 ;
        RECT 77.115 144.220 77.435 144.280 ;
        RECT 80.810 144.220 81.100 144.265 ;
        RECT 83.110 144.220 83.400 144.265 ;
        RECT 77.115 144.080 82.405 144.220 ;
        RECT 77.115 144.020 77.435 144.080 ;
        RECT 80.810 144.035 81.100 144.080 ;
        RECT 58.715 143.880 59.035 143.940 ;
        RECT 54.665 143.740 59.035 143.880 ;
        RECT 54.665 143.585 54.805 143.740 ;
        RECT 58.715 143.680 59.035 143.740 ;
        RECT 64.235 143.880 64.555 143.940 ;
        RECT 68.375 143.880 68.695 143.940 ;
        RECT 64.235 143.740 68.695 143.880 ;
        RECT 64.235 143.680 64.555 143.740 ;
        RECT 68.375 143.680 68.695 143.740 ;
        RECT 68.850 143.880 69.140 143.925 ;
        RECT 72.070 143.880 72.360 143.925 ;
        RECT 74.370 143.880 74.660 143.925 ;
        RECT 68.850 143.740 74.660 143.880 ;
        RECT 68.850 143.695 69.140 143.740 ;
        RECT 72.070 143.695 72.360 143.740 ;
        RECT 74.370 143.695 74.660 143.740 ;
        RECT 51.830 143.400 53.515 143.540 ;
        RECT 51.830 143.355 52.120 143.400 ;
        RECT 53.195 143.340 53.515 143.400 ;
        RECT 53.670 143.355 53.960 143.585 ;
        RECT 54.130 143.355 54.420 143.585 ;
        RECT 54.590 143.355 54.880 143.585 ;
        RECT 46.845 143.200 46.985 143.340 ;
        RECT 45.465 143.060 46.985 143.200 ;
        RECT 50.065 143.200 50.205 143.340 ;
        RECT 53.745 143.200 53.885 143.355 ;
        RECT 50.065 143.060 53.885 143.200 ;
        RECT 34.450 142.720 39.750 142.860 ;
        RECT 34.450 142.675 34.740 142.720 ;
        RECT 37.570 142.675 37.860 142.720 ;
        RECT 39.460 142.675 39.750 142.720 ;
        RECT 39.945 142.720 45.145 142.860 ;
        RECT 39.945 142.520 40.085 142.720 ;
        RECT 26.605 142.380 40.085 142.520 ;
        RECT 43.075 142.320 43.395 142.580 ;
        RECT 44.455 142.520 44.775 142.580 ;
        RECT 45.835 142.520 46.155 142.580 ;
        RECT 44.455 142.380 46.155 142.520 ;
        RECT 44.455 142.320 44.775 142.380 ;
        RECT 45.835 142.320 46.155 142.380 ;
        RECT 46.295 142.520 46.615 142.580 ;
        RECT 47.230 142.520 47.520 142.565 ;
        RECT 46.295 142.380 47.520 142.520 ;
        RECT 46.295 142.320 46.615 142.380 ;
        RECT 47.230 142.335 47.520 142.380 ;
        RECT 51.815 142.520 52.135 142.580 ;
        RECT 52.290 142.520 52.580 142.565 ;
        RECT 51.815 142.380 52.580 142.520 ;
        RECT 53.745 142.520 53.885 143.060 ;
        RECT 54.205 142.860 54.345 143.355 ;
        RECT 55.495 143.340 55.815 143.600 ;
        RECT 56.415 143.340 56.735 143.600 ;
        RECT 65.155 143.340 65.475 143.600 ;
        RECT 66.995 143.540 67.315 143.600 ;
        RECT 69.770 143.540 70.060 143.585 ;
        RECT 66.995 143.400 70.060 143.540 ;
        RECT 66.995 143.340 67.315 143.400 ;
        RECT 69.770 143.355 70.060 143.400 ;
        RECT 71.610 143.540 71.900 143.585 ;
        RECT 72.515 143.540 72.835 143.600 ;
        RECT 71.610 143.400 72.835 143.540 ;
        RECT 71.610 143.355 71.900 143.400 ;
        RECT 68.375 143.200 68.695 143.260 ;
        RECT 62.945 143.060 68.695 143.200 ;
        RECT 62.945 142.860 63.085 143.060 ;
        RECT 68.375 143.000 68.695 143.060 ;
        RECT 69.295 143.200 69.615 143.260 ;
        RECT 70.230 143.200 70.520 143.245 ;
        RECT 69.295 143.060 70.520 143.200 ;
        RECT 69.295 143.000 69.615 143.060 ;
        RECT 70.230 143.015 70.520 143.060 ;
        RECT 71.150 143.015 71.440 143.245 ;
        RECT 54.205 142.720 63.085 142.860 ;
        RECT 63.315 142.860 63.635 142.920 ;
        RECT 66.075 142.860 66.395 142.920 ;
        RECT 71.225 142.860 71.365 143.015 ;
        RECT 63.315 142.720 71.365 142.860 ;
        RECT 63.315 142.660 63.635 142.720 ;
        RECT 66.075 142.660 66.395 142.720 ;
        RECT 64.235 142.520 64.555 142.580 ;
        RECT 53.745 142.380 64.555 142.520 ;
        RECT 51.815 142.320 52.135 142.380 ;
        RECT 52.290 142.335 52.580 142.380 ;
        RECT 64.235 142.320 64.555 142.380 ;
        RECT 64.695 142.520 65.015 142.580 ;
        RECT 71.685 142.520 71.825 143.355 ;
        RECT 72.515 143.340 72.835 143.400 ;
        RECT 80.795 143.540 81.115 143.600 ;
        RECT 81.270 143.540 81.560 143.585 ;
        RECT 80.795 143.400 81.560 143.540 ;
        RECT 82.265 143.540 82.405 144.080 ;
        RECT 83.110 144.080 83.785 144.220 ;
        RECT 83.110 144.035 83.400 144.080 ;
        RECT 83.645 143.585 83.785 144.080 ;
        RECT 84.475 144.020 84.795 144.280 ;
        RECT 96.895 144.220 97.215 144.280 ;
        RECT 92.845 144.080 97.215 144.220 ;
        RECT 88.170 143.880 88.460 143.925 ;
        RECT 90.930 143.880 91.220 143.925 ;
        RECT 88.170 143.740 91.220 143.880 ;
        RECT 88.170 143.695 88.460 143.740 ;
        RECT 90.930 143.695 91.220 143.740 ;
        RECT 92.845 143.600 92.985 144.080 ;
        RECT 96.895 144.020 97.215 144.080 ;
        RECT 98.275 144.220 98.595 144.280 ;
        RECT 98.275 144.080 101.265 144.220 ;
        RECT 98.275 144.020 98.595 144.080 ;
        RECT 93.675 143.880 93.995 143.940 ;
        RECT 99.195 143.880 99.515 143.940 ;
        RECT 99.670 143.880 99.960 143.925 ;
        RECT 93.675 143.740 98.045 143.880 ;
        RECT 93.675 143.680 93.995 143.740 ;
        RECT 82.265 143.400 83.325 143.540 ;
        RECT 80.795 143.340 81.115 143.400 ;
        RECT 81.270 143.355 81.560 143.400 ;
        RECT 75.750 143.200 76.040 143.245 ;
        RECT 79.890 143.200 80.180 143.245 ;
        RECT 75.750 143.060 80.180 143.200 ;
        RECT 83.185 143.200 83.325 143.400 ;
        RECT 83.570 143.355 83.860 143.585 ;
        RECT 87.695 143.540 88.015 143.600 ;
        RECT 89.550 143.540 89.840 143.585 ;
        RECT 87.695 143.400 89.840 143.540 ;
        RECT 87.695 143.340 88.015 143.400 ;
        RECT 89.550 143.355 89.840 143.400 ;
        RECT 92.295 143.340 92.615 143.600 ;
        RECT 92.755 143.340 93.075 143.600 ;
        RECT 93.215 143.340 93.535 143.600 ;
        RECT 94.135 143.540 94.455 143.600 ;
        RECT 95.515 143.540 95.835 143.600 ;
        RECT 94.135 143.400 95.835 143.540 ;
        RECT 94.135 143.340 94.455 143.400 ;
        RECT 95.515 143.340 95.835 143.400 ;
        RECT 96.450 143.355 96.740 143.585 ;
        RECT 89.090 143.200 89.380 143.245 ;
        RECT 89.995 143.200 90.315 143.260 ;
        RECT 83.185 143.060 88.845 143.200 ;
        RECT 75.750 143.015 76.040 143.060 ;
        RECT 79.890 143.015 80.180 143.060 ;
        RECT 79.965 142.860 80.105 143.015 ;
        RECT 81.255 142.860 81.575 142.920 ;
        RECT 79.965 142.720 81.575 142.860 ;
        RECT 88.705 142.860 88.845 143.060 ;
        RECT 89.090 143.060 90.315 143.200 ;
        RECT 89.090 143.015 89.380 143.060 ;
        RECT 89.995 143.000 90.315 143.060 ;
        RECT 93.305 142.860 93.445 143.340 ;
        RECT 96.525 143.200 96.665 143.355 ;
        RECT 96.895 143.340 97.215 143.600 ;
        RECT 97.355 143.340 97.675 143.600 ;
        RECT 97.905 143.540 98.045 143.740 ;
        RECT 99.195 143.740 99.960 143.880 ;
        RECT 99.195 143.680 99.515 143.740 ;
        RECT 99.670 143.695 99.960 143.740 ;
        RECT 101.125 143.585 101.265 144.080 ;
        RECT 104.255 144.020 104.575 144.280 ;
        RECT 106.110 144.220 106.400 144.265 ;
        RECT 108.395 144.220 108.715 144.280 ;
        RECT 106.110 144.080 108.715 144.220 ;
        RECT 106.110 144.035 106.400 144.080 ;
        RECT 108.395 144.020 108.715 144.080 ;
        RECT 100.590 143.540 100.880 143.585 ;
        RECT 97.905 143.400 100.880 143.540 ;
        RECT 100.590 143.355 100.880 143.400 ;
        RECT 101.050 143.355 101.340 143.585 ;
        RECT 102.415 143.200 102.735 143.260 ;
        RECT 96.525 143.060 102.735 143.200 ;
        RECT 102.415 143.000 102.735 143.060 ;
        RECT 103.335 143.000 103.655 143.260 ;
        RECT 103.810 143.200 104.100 143.245 ;
        RECT 104.255 143.200 104.575 143.260 ;
        RECT 103.810 143.060 104.575 143.200 ;
        RECT 103.810 143.015 104.100 143.060 ;
        RECT 104.255 143.000 104.575 143.060 ;
        RECT 88.705 142.720 93.445 142.860 ;
        RECT 96.435 142.860 96.755 142.920 ;
        RECT 96.435 142.720 99.885 142.860 ;
        RECT 81.255 142.660 81.575 142.720 ;
        RECT 96.435 142.660 96.755 142.720 ;
        RECT 64.695 142.380 71.825 142.520 ;
        RECT 89.550 142.520 89.840 142.565 ;
        RECT 89.995 142.520 90.315 142.580 ;
        RECT 89.550 142.380 90.315 142.520 ;
        RECT 64.695 142.320 65.015 142.380 ;
        RECT 89.550 142.335 89.840 142.380 ;
        RECT 89.995 142.320 90.315 142.380 ;
        RECT 90.470 142.520 90.760 142.565 ;
        RECT 91.835 142.520 92.155 142.580 ;
        RECT 90.470 142.380 92.155 142.520 ;
        RECT 90.470 142.335 90.760 142.380 ;
        RECT 91.835 142.320 92.155 142.380 ;
        RECT 98.735 142.320 99.055 142.580 ;
        RECT 99.745 142.565 99.885 142.720 ;
        RECT 99.670 142.335 99.960 142.565 ;
        RECT 101.970 142.520 102.260 142.565 ;
        RECT 106.095 142.520 106.415 142.580 ;
        RECT 101.970 142.380 106.415 142.520 ;
        RECT 101.970 142.335 102.260 142.380 ;
        RECT 106.095 142.320 106.415 142.380 ;
        RECT 18.165 141.700 112.465 142.180 ;
        RECT 37.110 141.500 37.400 141.545 ;
        RECT 38.935 141.500 39.255 141.560 ;
        RECT 37.110 141.360 39.255 141.500 ;
        RECT 37.110 141.315 37.400 141.360 ;
        RECT 38.935 141.300 39.255 141.360 ;
        RECT 39.395 141.500 39.715 141.560 ;
        RECT 40.330 141.500 40.620 141.545 ;
        RECT 48.135 141.500 48.455 141.560 ;
        RECT 48.610 141.500 48.900 141.545 ;
        RECT 55.035 141.500 55.355 141.560 ;
        RECT 39.395 141.360 40.620 141.500 ;
        RECT 39.395 141.300 39.715 141.360 ;
        RECT 40.330 141.315 40.620 141.360 ;
        RECT 40.865 141.360 46.065 141.500 ;
        RECT 22.490 141.160 22.780 141.205 ;
        RECT 25.610 141.160 25.900 141.205 ;
        RECT 27.500 141.160 27.790 141.205 ;
        RECT 37.555 141.160 37.875 141.220 ;
        RECT 40.865 141.160 41.005 141.360 ;
        RECT 22.490 141.020 27.790 141.160 ;
        RECT 22.490 140.975 22.780 141.020 ;
        RECT 25.610 140.975 25.900 141.020 ;
        RECT 27.500 140.975 27.790 141.020 ;
        RECT 29.365 141.020 41.005 141.160 ;
        RECT 19.630 140.820 19.920 140.865 ;
        RECT 26.515 140.820 26.835 140.880 ;
        RECT 29.365 140.865 29.505 141.020 ;
        RECT 37.555 140.960 37.875 141.020 ;
        RECT 41.695 140.960 42.015 141.220 ;
        RECT 42.630 141.160 42.920 141.205 ;
        RECT 44.455 141.160 44.775 141.220 ;
        RECT 45.375 141.160 45.695 141.220 ;
        RECT 42.630 141.020 44.775 141.160 ;
        RECT 42.630 140.975 42.920 141.020 ;
        RECT 44.455 140.960 44.775 141.020 ;
        RECT 45.070 141.020 45.695 141.160 ;
        RECT 19.630 140.680 26.835 140.820 ;
        RECT 19.630 140.635 19.920 140.680 ;
        RECT 26.515 140.620 26.835 140.680 ;
        RECT 29.290 140.635 29.580 140.865 ;
        RECT 31.115 140.820 31.435 140.880 ;
        RECT 35.715 140.820 36.035 140.880 ;
        RECT 38.490 140.820 38.780 140.865 ;
        RECT 40.315 140.820 40.635 140.880 ;
        RECT 31.115 140.680 38.780 140.820 ;
        RECT 31.115 140.620 31.435 140.680 ;
        RECT 35.715 140.620 36.035 140.680 ;
        RECT 38.490 140.635 38.780 140.680 ;
        RECT 39.945 140.680 40.635 140.820 ;
        RECT 21.410 140.185 21.700 140.500 ;
        RECT 22.490 140.480 22.780 140.525 ;
        RECT 26.070 140.480 26.360 140.525 ;
        RECT 27.905 140.480 28.195 140.525 ;
        RECT 22.490 140.340 28.195 140.480 ;
        RECT 22.490 140.295 22.780 140.340 ;
        RECT 26.070 140.295 26.360 140.340 ;
        RECT 27.905 140.295 28.195 140.340 ;
        RECT 28.370 140.480 28.660 140.525 ;
        RECT 31.575 140.480 31.895 140.540 ;
        RECT 28.370 140.340 31.895 140.480 ;
        RECT 28.370 140.295 28.660 140.340 ;
        RECT 31.575 140.280 31.895 140.340 ;
        RECT 33.875 140.480 34.195 140.540 ;
        RECT 34.350 140.480 34.640 140.525 ;
        RECT 33.875 140.340 34.640 140.480 ;
        RECT 33.875 140.280 34.195 140.340 ;
        RECT 34.350 140.295 34.640 140.340 ;
        RECT 36.175 140.280 36.495 140.540 ;
        RECT 39.945 140.525 40.085 140.680 ;
        RECT 40.315 140.620 40.635 140.680 ;
        RECT 41.235 140.620 41.555 140.880 ;
        RECT 41.785 140.820 41.925 140.960 ;
        RECT 41.785 140.680 44.685 140.820 ;
        RECT 39.870 140.295 40.160 140.525 ;
        RECT 41.710 140.480 42.000 140.525 ;
        RECT 42.155 140.480 42.475 140.540 ;
        RECT 44.545 140.525 44.685 140.680 ;
        RECT 45.070 140.525 45.210 141.020 ;
        RECT 45.375 140.960 45.695 141.020 ;
        RECT 45.925 140.820 46.065 141.360 ;
        RECT 48.135 141.360 48.900 141.500 ;
        RECT 48.135 141.300 48.455 141.360 ;
        RECT 48.610 141.315 48.900 141.360 ;
        RECT 49.145 141.360 55.355 141.500 ;
        RECT 49.145 141.160 49.285 141.360 ;
        RECT 55.035 141.300 55.355 141.360 ;
        RECT 55.495 141.500 55.815 141.560 ;
        RECT 62.855 141.500 63.175 141.560 ;
        RECT 63.790 141.500 64.080 141.545 ;
        RECT 55.495 141.360 64.080 141.500 ;
        RECT 55.495 141.300 55.815 141.360 ;
        RECT 62.855 141.300 63.175 141.360 ;
        RECT 63.790 141.315 64.080 141.360 ;
        RECT 64.235 141.500 64.555 141.560 ;
        RECT 66.090 141.500 66.380 141.545 ;
        RECT 64.235 141.360 66.380 141.500 ;
        RECT 64.235 141.300 64.555 141.360 ;
        RECT 66.090 141.315 66.380 141.360 ;
        RECT 68.835 141.500 69.155 141.560 ;
        RECT 70.675 141.500 70.995 141.560 ;
        RECT 72.975 141.500 73.295 141.560 ;
        RECT 90.470 141.500 90.760 141.545 ;
        RECT 90.915 141.500 91.235 141.560 ;
        RECT 68.835 141.360 72.745 141.500 ;
        RECT 68.835 141.300 69.155 141.360 ;
        RECT 70.675 141.300 70.995 141.360 ;
        RECT 45.465 140.680 46.065 140.820 ;
        RECT 48.225 141.020 49.285 141.160 ;
        RECT 54.230 141.160 54.520 141.205 ;
        RECT 57.350 141.160 57.640 141.205 ;
        RECT 59.240 141.160 59.530 141.205 ;
        RECT 54.230 141.020 59.530 141.160 ;
        RECT 45.465 140.525 45.605 140.680 ;
        RECT 41.710 140.340 42.475 140.480 ;
        RECT 41.710 140.295 42.000 140.340 ;
        RECT 42.155 140.280 42.475 140.340 ;
        RECT 44.470 140.295 44.760 140.525 ;
        RECT 44.930 140.295 45.220 140.525 ;
        RECT 45.390 140.295 45.680 140.525 ;
        RECT 45.835 140.480 46.155 140.540 ;
        RECT 46.310 140.480 46.600 140.525 ;
        RECT 45.835 140.340 46.600 140.480 ;
        RECT 21.110 140.140 21.700 140.185 ;
        RECT 23.295 140.140 23.615 140.200 ;
        RECT 24.350 140.140 25.000 140.185 ;
        RECT 21.110 140.000 25.000 140.140 ;
        RECT 21.110 139.955 21.400 140.000 ;
        RECT 23.295 139.940 23.615 140.000 ;
        RECT 24.350 139.955 25.000 140.000 ;
        RECT 26.975 139.940 27.295 140.200 ;
        RECT 36.635 140.140 36.955 140.200 ;
        RECT 27.985 140.000 36.955 140.140 ;
        RECT 27.985 139.860 28.125 140.000 ;
        RECT 36.635 139.940 36.955 140.000 ;
        RECT 40.330 140.140 40.620 140.185 ;
        RECT 40.775 140.140 41.095 140.200 ;
        RECT 40.330 140.000 41.095 140.140 ;
        RECT 44.545 140.140 44.685 140.295 ;
        RECT 45.835 140.280 46.155 140.340 ;
        RECT 46.310 140.295 46.600 140.340 ;
        RECT 47.230 140.480 47.520 140.525 ;
        RECT 48.225 140.480 48.365 141.020 ;
        RECT 54.230 140.975 54.520 141.020 ;
        RECT 57.350 140.975 57.640 141.020 ;
        RECT 59.240 140.975 59.530 141.020 ;
        RECT 61.950 141.160 62.240 141.205 ;
        RECT 61.950 141.020 72.285 141.160 ;
        RECT 61.950 140.975 62.240 141.020 ;
        RECT 49.055 140.620 49.375 140.880 ;
        RECT 49.515 140.820 49.835 140.880 ;
        RECT 62.025 140.820 62.165 140.975 ;
        RECT 49.515 140.680 62.165 140.820 ;
        RECT 67.915 140.820 68.235 140.880 ;
        RECT 68.850 140.820 69.140 140.865 ;
        RECT 67.915 140.680 69.140 140.820 ;
        RECT 49.515 140.620 49.835 140.680 ;
        RECT 67.915 140.620 68.235 140.680 ;
        RECT 68.850 140.635 69.140 140.680 ;
        RECT 47.230 140.340 48.365 140.480 ;
        RECT 47.230 140.295 47.520 140.340 ;
        RECT 48.595 140.280 48.915 140.540 ;
        RECT 49.975 140.280 50.295 140.540 ;
        RECT 46.755 140.140 47.075 140.200 ;
        RECT 53.150 140.185 53.440 140.500 ;
        RECT 54.230 140.480 54.520 140.525 ;
        RECT 57.810 140.480 58.100 140.525 ;
        RECT 59.645 140.480 59.935 140.525 ;
        RECT 54.230 140.340 59.935 140.480 ;
        RECT 54.230 140.295 54.520 140.340 ;
        RECT 57.810 140.295 58.100 140.340 ;
        RECT 59.645 140.295 59.935 140.340 ;
        RECT 60.095 140.280 60.415 140.540 ;
        RECT 62.395 140.480 62.715 140.540 ;
        RECT 62.870 140.480 63.160 140.525 ;
        RECT 64.695 140.480 65.015 140.540 ;
        RECT 62.395 140.340 65.015 140.480 ;
        RECT 62.395 140.280 62.715 140.340 ;
        RECT 62.870 140.295 63.160 140.340 ;
        RECT 64.695 140.280 65.015 140.340 ;
        RECT 65.170 140.480 65.460 140.525 ;
        RECT 66.995 140.480 67.315 140.540 ;
        RECT 65.170 140.340 67.315 140.480 ;
        RECT 65.170 140.295 65.460 140.340 ;
        RECT 66.995 140.280 67.315 140.340 ;
        RECT 70.230 140.295 70.520 140.525 ;
        RECT 44.545 140.000 47.075 140.140 ;
        RECT 40.330 139.955 40.620 140.000 ;
        RECT 40.775 139.940 41.095 140.000 ;
        RECT 46.755 139.940 47.075 140.000 ;
        RECT 47.690 140.140 47.980 140.185 ;
        RECT 52.850 140.140 53.440 140.185 ;
        RECT 56.090 140.140 56.740 140.185 ;
        RECT 47.690 140.000 56.740 140.140 ;
        RECT 47.690 139.955 47.980 140.000 ;
        RECT 52.850 139.955 53.140 140.000 ;
        RECT 56.090 139.955 56.740 140.000 ;
        RECT 58.730 140.140 59.020 140.185 ;
        RECT 59.175 140.140 59.495 140.200 ;
        RECT 58.730 140.000 59.495 140.140 ;
        RECT 58.730 139.955 59.020 140.000 ;
        RECT 59.175 139.940 59.495 140.000 ;
        RECT 61.475 140.140 61.795 140.200 ;
        RECT 70.305 140.140 70.445 140.295 ;
        RECT 70.675 140.280 70.995 140.540 ;
        RECT 71.150 140.480 71.440 140.525 ;
        RECT 71.595 140.480 71.915 140.540 ;
        RECT 72.145 140.525 72.285 141.020 ;
        RECT 72.605 140.820 72.745 141.360 ;
        RECT 72.975 141.360 90.225 141.500 ;
        RECT 72.975 141.300 73.295 141.360 ;
        RECT 75.735 141.160 76.055 141.220 ;
        RECT 74.445 141.020 76.055 141.160 ;
        RECT 74.445 140.820 74.585 141.020 ;
        RECT 75.735 140.960 76.055 141.020 ;
        RECT 80.765 141.160 81.055 141.205 ;
        RECT 83.545 141.160 83.835 141.205 ;
        RECT 85.405 141.160 85.695 141.205 ;
        RECT 80.765 141.020 85.695 141.160 ;
        RECT 90.085 141.160 90.225 141.360 ;
        RECT 90.470 141.360 91.235 141.500 ;
        RECT 90.470 141.315 90.760 141.360 ;
        RECT 90.915 141.300 91.235 141.360 ;
        RECT 92.295 141.500 92.615 141.560 ;
        RECT 93.675 141.500 93.995 141.560 ;
        RECT 99.670 141.500 99.960 141.545 ;
        RECT 92.295 141.360 93.445 141.500 ;
        RECT 92.295 141.300 92.615 141.360 ;
        RECT 92.755 141.160 93.075 141.220 ;
        RECT 90.085 141.020 93.075 141.160 ;
        RECT 80.765 140.975 81.055 141.020 ;
        RECT 83.545 140.975 83.835 141.020 ;
        RECT 85.405 140.975 85.695 141.020 ;
        RECT 92.755 140.960 93.075 141.020 ;
        RECT 72.605 140.680 74.585 140.820 ;
        RECT 71.150 140.340 71.915 140.480 ;
        RECT 71.150 140.295 71.440 140.340 ;
        RECT 71.595 140.280 71.915 140.340 ;
        RECT 72.070 140.480 72.360 140.525 ;
        RECT 72.975 140.480 73.295 140.540 ;
        RECT 74.445 140.525 74.585 140.680 ;
        RECT 90.010 140.820 90.300 140.865 ;
        RECT 90.455 140.820 90.775 140.880 ;
        RECT 90.010 140.680 90.775 140.820 ;
        RECT 90.010 140.635 90.300 140.680 ;
        RECT 90.455 140.620 90.775 140.680 ;
        RECT 72.070 140.340 73.295 140.480 ;
        RECT 72.070 140.295 72.360 140.340 ;
        RECT 72.975 140.280 73.295 140.340 ;
        RECT 73.910 140.295 74.200 140.525 ;
        RECT 74.370 140.295 74.660 140.525 ;
        RECT 74.830 140.490 75.120 140.525 ;
        RECT 74.830 140.350 75.505 140.490 ;
        RECT 74.830 140.295 75.120 140.350 ;
        RECT 73.985 140.140 74.125 140.295 ;
        RECT 61.475 140.000 74.125 140.140 ;
        RECT 61.475 139.940 61.795 140.000 ;
        RECT 27.895 139.600 28.215 139.860 ;
        RECT 32.035 139.600 32.355 139.860 ;
        RECT 32.495 139.800 32.815 139.860 ;
        RECT 33.430 139.800 33.720 139.845 ;
        RECT 32.495 139.660 33.720 139.800 ;
        RECT 32.495 139.600 32.815 139.660 ;
        RECT 33.430 139.615 33.720 139.660 ;
        RECT 43.090 139.800 43.380 139.845 ;
        RECT 43.535 139.800 43.855 139.860 ;
        RECT 43.090 139.660 43.855 139.800 ;
        RECT 43.090 139.615 43.380 139.660 ;
        RECT 43.535 139.600 43.855 139.660 ;
        RECT 49.975 139.800 50.295 139.860 ;
        RECT 50.910 139.800 51.200 139.845 ;
        RECT 49.975 139.660 51.200 139.800 ;
        RECT 49.975 139.600 50.295 139.660 ;
        RECT 50.910 139.615 51.200 139.660 ;
        RECT 51.370 139.800 51.660 139.845 ;
        RECT 53.655 139.800 53.975 139.860 ;
        RECT 57.795 139.800 58.115 139.860 ;
        RECT 51.370 139.660 58.115 139.800 ;
        RECT 51.370 139.615 51.660 139.660 ;
        RECT 53.655 139.600 53.975 139.660 ;
        RECT 57.795 139.600 58.115 139.660 ;
        RECT 67.930 139.800 68.220 139.845 ;
        RECT 68.375 139.800 68.695 139.860 ;
        RECT 67.930 139.660 68.695 139.800 ;
        RECT 70.305 139.800 70.445 140.000 ;
        RECT 70.675 139.800 70.995 139.860 ;
        RECT 70.305 139.660 70.995 139.800 ;
        RECT 67.930 139.615 68.220 139.660 ;
        RECT 68.375 139.600 68.695 139.660 ;
        RECT 70.675 139.600 70.995 139.660 ;
        RECT 72.530 139.800 72.820 139.845 ;
        RECT 73.895 139.800 74.215 139.860 ;
        RECT 72.530 139.660 74.215 139.800 ;
        RECT 72.530 139.615 72.820 139.660 ;
        RECT 73.895 139.600 74.215 139.660 ;
        RECT 74.355 139.800 74.675 139.860 ;
        RECT 75.365 139.800 75.505 140.350 ;
        RECT 75.750 140.480 76.040 140.525 ;
        RECT 76.655 140.480 76.975 140.540 ;
        RECT 75.750 140.340 76.975 140.480 ;
        RECT 75.750 140.295 76.040 140.340 ;
        RECT 76.655 140.280 76.975 140.340 ;
        RECT 80.765 140.480 81.055 140.525 ;
        RECT 84.030 140.480 84.320 140.525 ;
        RECT 85.395 140.480 85.715 140.540 ;
        RECT 80.765 140.340 83.300 140.480 ;
        RECT 80.765 140.295 81.055 140.340 ;
        RECT 83.085 140.185 83.300 140.340 ;
        RECT 84.030 140.340 85.715 140.480 ;
        RECT 84.030 140.295 84.320 140.340 ;
        RECT 85.395 140.280 85.715 140.340 ;
        RECT 85.870 140.480 86.160 140.525 ;
        RECT 87.235 140.480 87.555 140.540 ;
        RECT 85.870 140.340 87.555 140.480 ;
        RECT 85.870 140.295 86.160 140.340 ;
        RECT 87.235 140.280 87.555 140.340 ;
        RECT 89.090 140.480 89.380 140.525 ;
        RECT 91.375 140.480 91.695 140.540 ;
        RECT 89.090 140.340 91.695 140.480 ;
        RECT 89.090 140.295 89.380 140.340 ;
        RECT 91.375 140.280 91.695 140.340 ;
        RECT 92.295 140.280 92.615 140.540 ;
        RECT 92.845 140.525 92.985 140.960 ;
        RECT 93.305 140.820 93.445 141.360 ;
        RECT 93.675 141.360 99.960 141.500 ;
        RECT 93.675 141.300 93.995 141.360 ;
        RECT 99.670 141.315 99.960 141.360 ;
        RECT 135.635 141.220 136.775 165.470 ;
        RECT 95.515 141.160 95.835 141.220 ;
        RECT 101.970 141.160 102.260 141.205 ;
        RECT 95.515 141.020 102.260 141.160 ;
        RECT 95.515 140.960 95.835 141.020 ;
        RECT 101.970 140.975 102.260 141.020 ;
        RECT 106.110 140.975 106.400 141.205 ;
        RECT 95.975 140.820 96.295 140.880 ;
        RECT 100.130 140.820 100.420 140.865 ;
        RECT 93.305 140.680 94.825 140.820 ;
        RECT 92.770 140.295 93.060 140.525 ;
        RECT 78.905 140.140 79.195 140.185 ;
        RECT 82.165 140.140 82.455 140.185 ;
        RECT 83.085 140.140 83.375 140.185 ;
        RECT 84.945 140.140 85.235 140.185 ;
        RECT 78.905 140.000 82.865 140.140 ;
        RECT 78.905 139.955 79.195 140.000 ;
        RECT 82.165 139.955 82.455 140.000 ;
        RECT 74.355 139.660 75.505 139.800 ;
        RECT 76.900 139.800 77.190 139.845 ;
        RECT 80.795 139.800 81.115 139.860 ;
        RECT 76.900 139.660 81.115 139.800 ;
        RECT 82.725 139.800 82.865 140.000 ;
        RECT 83.085 140.000 85.235 140.140 ;
        RECT 83.085 139.955 83.375 140.000 ;
        RECT 84.945 139.955 85.235 140.000 ;
        RECT 90.470 140.140 90.760 140.185 ;
        RECT 90.930 140.140 91.220 140.185 ;
        RECT 90.470 140.000 91.220 140.140 ;
        RECT 92.845 140.140 92.985 140.295 ;
        RECT 93.215 140.280 93.535 140.540 ;
        RECT 94.135 140.280 94.455 140.540 ;
        RECT 94.685 140.480 94.825 140.680 ;
        RECT 95.975 140.680 100.420 140.820 ;
        RECT 95.975 140.620 96.295 140.680 ;
        RECT 100.130 140.635 100.420 140.680 ;
        RECT 103.335 140.620 103.655 140.880 ;
        RECT 106.185 140.820 106.325 140.975 ;
        RECT 106.185 140.680 108.165 140.820 ;
        RECT 97.355 140.480 97.675 140.540 ;
        RECT 94.685 140.340 97.675 140.480 ;
        RECT 97.355 140.280 97.675 140.340 ;
        RECT 97.830 140.295 98.120 140.525 ;
        RECT 98.290 140.295 98.580 140.525 ;
        RECT 92.845 140.000 96.665 140.140 ;
        RECT 90.470 139.955 90.760 140.000 ;
        RECT 90.930 139.955 91.220 140.000 ;
        RECT 84.475 139.800 84.795 139.860 ;
        RECT 82.725 139.660 84.795 139.800 ;
        RECT 74.355 139.600 74.675 139.660 ;
        RECT 76.900 139.615 77.190 139.660 ;
        RECT 80.795 139.600 81.115 139.660 ;
        RECT 84.475 139.600 84.795 139.660 ;
        RECT 87.695 139.800 88.015 139.860 ;
        RECT 88.170 139.800 88.460 139.845 ;
        RECT 87.695 139.660 88.460 139.800 ;
        RECT 87.695 139.600 88.015 139.660 ;
        RECT 88.170 139.615 88.460 139.660 ;
        RECT 95.975 139.600 96.295 139.860 ;
        RECT 96.525 139.800 96.665 140.000 ;
        RECT 97.905 139.800 98.045 140.295 ;
        RECT 96.525 139.660 98.045 139.800 ;
        RECT 98.365 139.800 98.505 140.295 ;
        RECT 99.195 140.280 99.515 140.540 ;
        RECT 101.050 140.480 101.340 140.525 ;
        RECT 102.875 140.480 103.195 140.540 ;
        RECT 101.050 140.340 103.195 140.480 ;
        RECT 101.050 140.295 101.340 140.340 ;
        RECT 102.875 140.280 103.195 140.340 ;
        RECT 104.255 140.280 104.575 140.540 ;
        RECT 104.715 140.480 105.035 140.540 ;
        RECT 106.555 140.480 106.875 140.540 ;
        RECT 108.025 140.525 108.165 140.680 ;
        RECT 104.715 140.340 106.875 140.480 ;
        RECT 104.715 140.280 105.035 140.340 ;
        RECT 106.555 140.280 106.875 140.340 ;
        RECT 107.950 140.295 108.240 140.525 ;
        RECT 135.580 140.230 136.830 141.220 ;
        RECT 98.735 140.140 99.055 140.200 ;
        RECT 99.670 140.140 99.960 140.185 ;
        RECT 98.735 140.000 99.960 140.140 ;
        RECT 98.735 139.940 99.055 140.000 ;
        RECT 99.670 139.955 99.960 140.000 ;
        RECT 102.415 140.140 102.735 140.200 ;
        RECT 103.810 140.140 104.100 140.185 ;
        RECT 135.635 140.155 136.775 140.230 ;
        RECT 102.415 140.000 104.100 140.140 ;
        RECT 102.415 139.940 102.735 140.000 ;
        RECT 103.810 139.955 104.100 140.000 ;
        RECT 102.875 139.800 103.195 139.860 ;
        RECT 98.365 139.660 103.195 139.800 ;
        RECT 102.875 139.600 103.195 139.660 ;
        RECT 106.555 139.800 106.875 139.860 ;
        RECT 107.030 139.800 107.320 139.845 ;
        RECT 106.555 139.660 107.320 139.800 ;
        RECT 106.555 139.600 106.875 139.660 ;
        RECT 107.030 139.615 107.320 139.660 ;
        RECT 108.855 139.600 109.175 139.860 ;
        RECT 17.370 138.980 112.465 139.460 ;
        RECT 132.510 139.190 135.210 140.010 ;
        RECT 143.370 139.390 144.510 223.840 ;
        RECT 137.240 139.380 144.510 139.390 ;
        RECT 136.210 139.190 144.510 139.380 ;
        RECT 22.850 138.780 23.140 138.825 ;
        RECT 23.295 138.780 23.615 138.840 ;
        RECT 22.850 138.640 23.615 138.780 ;
        RECT 22.850 138.595 23.140 138.640 ;
        RECT 23.295 138.580 23.615 138.640 ;
        RECT 26.975 138.780 27.295 138.840 ;
        RECT 27.910 138.780 28.200 138.825 ;
        RECT 26.975 138.640 28.200 138.780 ;
        RECT 26.975 138.580 27.295 138.640 ;
        RECT 27.910 138.595 28.200 138.640 ;
        RECT 31.575 138.780 31.895 138.840 ;
        RECT 47.675 138.780 47.995 138.840 ;
        RECT 31.575 138.640 34.565 138.780 ;
        RECT 31.575 138.580 31.895 138.640 ;
        RECT 31.115 138.440 31.435 138.500 ;
        RECT 23.385 138.300 31.435 138.440 ;
        RECT 21.470 138.100 21.760 138.145 ;
        RECT 22.835 138.100 23.155 138.160 ;
        RECT 23.385 138.145 23.525 138.300 ;
        RECT 31.115 138.240 31.435 138.300 ;
        RECT 32.495 138.240 32.815 138.500 ;
        RECT 34.425 138.440 34.565 138.640 ;
        RECT 41.325 138.640 47.995 138.780 ;
        RECT 34.790 138.440 35.440 138.485 ;
        RECT 38.390 138.440 38.680 138.485 ;
        RECT 34.425 138.300 38.680 138.440 ;
        RECT 34.790 138.255 35.440 138.300 ;
        RECT 38.090 138.255 38.680 138.300 ;
        RECT 23.310 138.100 23.600 138.145 ;
        RECT 21.470 137.960 23.600 138.100 ;
        RECT 21.470 137.915 21.760 137.960 ;
        RECT 22.835 137.900 23.155 137.960 ;
        RECT 23.310 137.915 23.600 137.960 ;
        RECT 25.595 137.900 25.915 138.160 ;
        RECT 28.830 138.100 29.120 138.145 ;
        RECT 27.525 137.960 29.120 138.100 ;
        RECT 24.690 137.575 24.980 137.805 ;
        RECT 25.150 137.760 25.440 137.805 ;
        RECT 26.515 137.760 26.835 137.820 ;
        RECT 25.150 137.620 27.205 137.760 ;
        RECT 25.150 137.575 25.440 137.620 ;
        RECT 24.765 137.420 24.905 137.575 ;
        RECT 26.515 137.560 26.835 137.620 ;
        RECT 26.055 137.420 26.375 137.480 ;
        RECT 24.765 137.280 26.375 137.420 ;
        RECT 26.055 137.220 26.375 137.280 ;
        RECT 20.995 136.880 21.315 137.140 ;
        RECT 27.065 137.080 27.205 137.620 ;
        RECT 27.525 137.465 27.665 137.960 ;
        RECT 28.830 137.915 29.120 137.960 ;
        RECT 31.595 138.100 31.885 138.145 ;
        RECT 33.430 138.100 33.720 138.145 ;
        RECT 37.010 138.100 37.300 138.145 ;
        RECT 31.595 137.960 37.300 138.100 ;
        RECT 31.595 137.915 31.885 137.960 ;
        RECT 33.430 137.915 33.720 137.960 ;
        RECT 37.010 137.915 37.300 137.960 ;
        RECT 38.090 137.940 38.380 138.255 ;
        RECT 41.325 138.145 41.465 138.640 ;
        RECT 47.675 138.580 47.995 138.640 ;
        RECT 59.175 138.780 59.495 138.840 ;
        RECT 61.950 138.780 62.240 138.825 ;
        RECT 59.175 138.640 62.240 138.780 ;
        RECT 59.175 138.580 59.495 138.640 ;
        RECT 61.950 138.595 62.240 138.640 ;
        RECT 62.855 138.780 63.175 138.840 ;
        RECT 67.455 138.780 67.775 138.840 ;
        RECT 62.855 138.640 67.775 138.780 ;
        RECT 62.855 138.580 63.175 138.640 ;
        RECT 67.455 138.580 67.775 138.640 ;
        RECT 67.930 138.780 68.220 138.825 ;
        RECT 68.835 138.780 69.155 138.840 ;
        RECT 67.930 138.640 69.155 138.780 ;
        RECT 67.930 138.595 68.220 138.640 ;
        RECT 68.835 138.580 69.155 138.640 ;
        RECT 71.135 138.780 71.455 138.840 ;
        RECT 80.795 138.780 81.115 138.840 ;
        RECT 81.270 138.780 81.560 138.825 ;
        RECT 71.135 138.640 72.745 138.780 ;
        RECT 71.135 138.580 71.455 138.640 ;
        RECT 42.155 138.440 42.475 138.500 ;
        RECT 42.630 138.440 42.920 138.485 ;
        RECT 47.215 138.440 47.535 138.500 ;
        RECT 42.155 138.300 42.920 138.440 ;
        RECT 42.155 138.240 42.475 138.300 ;
        RECT 42.630 138.255 42.920 138.300 ;
        RECT 43.625 138.300 47.535 138.440 ;
        RECT 43.625 138.145 43.765 138.300 ;
        RECT 47.215 138.240 47.535 138.300 ;
        RECT 54.525 138.440 54.815 138.485 ;
        RECT 55.495 138.440 55.815 138.500 ;
        RECT 57.785 138.440 58.075 138.485 ;
        RECT 54.525 138.300 58.075 138.440 ;
        RECT 54.525 138.255 54.815 138.300 ;
        RECT 55.495 138.240 55.815 138.300 ;
        RECT 57.785 138.255 58.075 138.300 ;
        RECT 58.705 138.440 58.995 138.485 ;
        RECT 60.565 138.440 60.855 138.485 ;
        RECT 70.215 138.440 70.535 138.500 ;
        RECT 58.705 138.300 60.855 138.440 ;
        RECT 58.705 138.255 58.995 138.300 ;
        RECT 60.565 138.255 60.855 138.300 ;
        RECT 64.785 138.300 67.225 138.440 ;
        RECT 41.250 137.915 41.540 138.145 ;
        RECT 43.550 137.915 43.840 138.145 ;
        RECT 44.470 138.100 44.760 138.145 ;
        RECT 44.085 137.960 44.760 138.100 ;
        RECT 31.130 137.760 31.420 137.805 ;
        RECT 34.335 137.760 34.655 137.820 ;
        RECT 42.170 137.760 42.460 137.805 ;
        RECT 42.615 137.760 42.935 137.820 ;
        RECT 31.130 137.620 34.655 137.760 ;
        RECT 31.130 137.575 31.420 137.620 ;
        RECT 34.335 137.560 34.655 137.620 ;
        RECT 37.645 137.620 40.545 137.760 ;
        RECT 27.450 137.235 27.740 137.465 ;
        RECT 32.000 137.420 32.290 137.465 ;
        RECT 33.890 137.420 34.180 137.465 ;
        RECT 37.010 137.420 37.300 137.465 ;
        RECT 32.000 137.280 37.300 137.420 ;
        RECT 32.000 137.235 32.290 137.280 ;
        RECT 33.890 137.235 34.180 137.280 ;
        RECT 37.010 137.235 37.300 137.280 ;
        RECT 37.645 137.080 37.785 137.620 ;
        RECT 38.475 137.420 38.795 137.480 ;
        RECT 39.870 137.420 40.160 137.465 ;
        RECT 38.475 137.280 40.160 137.420 ;
        RECT 40.405 137.420 40.545 137.620 ;
        RECT 42.170 137.620 42.935 137.760 ;
        RECT 42.170 137.575 42.460 137.620 ;
        RECT 42.615 137.560 42.935 137.620 ;
        RECT 44.085 137.420 44.225 137.960 ;
        RECT 44.470 137.915 44.760 137.960 ;
        RECT 44.930 137.915 45.220 138.145 ;
        RECT 45.390 138.100 45.680 138.145 ;
        RECT 46.755 138.100 47.075 138.160 ;
        RECT 47.675 138.100 47.995 138.160 ;
        RECT 45.390 137.960 47.995 138.100 ;
        RECT 45.390 137.915 45.680 137.960 ;
        RECT 45.005 137.760 45.145 137.915 ;
        RECT 46.755 137.900 47.075 137.960 ;
        RECT 47.675 137.900 47.995 137.960 ;
        RECT 49.990 137.915 50.280 138.145 ;
        RECT 45.005 137.620 45.605 137.760 ;
        RECT 45.465 137.480 45.605 137.620 ;
        RECT 47.215 137.560 47.535 137.820 ;
        RECT 40.405 137.280 44.225 137.420 ;
        RECT 38.475 137.220 38.795 137.280 ;
        RECT 39.870 137.235 40.160 137.280 ;
        RECT 45.375 137.220 45.695 137.480 ;
        RECT 45.835 137.420 46.155 137.480 ;
        RECT 47.305 137.420 47.445 137.560 ;
        RECT 49.515 137.420 49.835 137.480 ;
        RECT 45.835 137.280 49.835 137.420 ;
        RECT 50.065 137.420 50.205 137.915 ;
        RECT 50.435 137.900 50.755 138.160 ;
        RECT 50.910 137.915 51.200 138.145 ;
        RECT 51.830 138.100 52.120 138.145 ;
        RECT 52.275 138.100 52.595 138.160 ;
        RECT 51.830 137.960 52.595 138.100 ;
        RECT 51.830 137.915 52.120 137.960 ;
        RECT 50.985 137.760 51.125 137.915 ;
        RECT 52.275 137.900 52.595 137.960 ;
        RECT 56.385 138.100 56.675 138.145 ;
        RECT 58.705 138.100 58.920 138.255 ;
        RECT 56.385 137.960 58.920 138.100 ;
        RECT 61.015 138.100 61.335 138.160 ;
        RECT 64.785 138.145 64.925 138.300 ;
        RECT 67.085 138.145 67.225 138.300 ;
        RECT 70.215 138.300 71.825 138.440 ;
        RECT 70.215 138.240 70.535 138.300 ;
        RECT 62.870 138.100 63.160 138.145 ;
        RECT 61.015 137.960 63.160 138.100 ;
        RECT 56.385 137.915 56.675 137.960 ;
        RECT 61.015 137.900 61.335 137.960 ;
        RECT 62.870 137.915 63.160 137.960 ;
        RECT 64.710 137.915 65.000 138.145 ;
        RECT 65.170 137.915 65.460 138.145 ;
        RECT 67.010 138.100 67.300 138.145 ;
        RECT 69.295 138.100 69.615 138.160 ;
        RECT 67.010 137.960 69.615 138.100 ;
        RECT 67.010 137.915 67.300 137.960 ;
        RECT 53.655 137.760 53.975 137.820 ;
        RECT 50.985 137.620 53.975 137.760 ;
        RECT 53.655 137.560 53.975 137.620 ;
        RECT 59.635 137.560 59.955 137.820 ;
        RECT 60.095 137.760 60.415 137.820 ;
        RECT 61.490 137.760 61.780 137.805 ;
        RECT 60.095 137.620 61.780 137.760 ;
        RECT 60.095 137.560 60.415 137.620 ;
        RECT 61.490 137.575 61.780 137.620 ;
        RECT 62.395 137.760 62.715 137.820 ;
        RECT 65.245 137.760 65.385 137.915 ;
        RECT 69.295 137.900 69.615 137.960 ;
        RECT 70.675 138.100 70.995 138.160 ;
        RECT 71.685 138.145 71.825 138.300 ;
        RECT 71.150 138.100 71.440 138.145 ;
        RECT 70.675 137.960 71.440 138.100 ;
        RECT 70.675 137.900 70.995 137.960 ;
        RECT 71.150 137.915 71.440 137.960 ;
        RECT 71.610 137.915 71.900 138.145 ;
        RECT 72.070 138.100 72.360 138.145 ;
        RECT 72.605 138.100 72.745 138.640 ;
        RECT 80.795 138.640 81.560 138.780 ;
        RECT 80.795 138.580 81.115 138.640 ;
        RECT 81.270 138.595 81.560 138.640 ;
        RECT 84.475 138.580 84.795 138.840 ;
        RECT 85.395 138.580 85.715 138.840 ;
        RECT 101.740 138.780 102.030 138.825 ;
        RECT 102.415 138.780 102.735 138.840 ;
        RECT 101.740 138.640 102.735 138.780 ;
        RECT 101.740 138.595 102.030 138.640 ;
        RECT 102.415 138.580 102.735 138.640 ;
        RECT 132.510 138.530 144.510 139.190 ;
        RECT 76.655 138.440 76.975 138.500 ;
        RECT 93.690 138.440 93.980 138.485 ;
        RECT 95.975 138.440 96.295 138.500 ;
        RECT 97.355 138.440 97.675 138.500 ;
        RECT 73.065 138.300 77.345 138.440 ;
        RECT 73.065 138.160 73.205 138.300 ;
        RECT 76.655 138.240 76.975 138.300 ;
        RECT 72.070 137.960 72.745 138.100 ;
        RECT 72.070 137.915 72.360 137.960 ;
        RECT 62.395 137.620 65.385 137.760 ;
        RECT 71.225 137.760 71.365 137.915 ;
        RECT 72.975 137.900 73.295 138.160 ;
        RECT 75.290 138.100 75.580 138.145 ;
        RECT 73.755 137.960 75.580 138.100 ;
        RECT 73.755 137.760 73.895 137.960 ;
        RECT 75.290 137.915 75.580 137.960 ;
        RECT 75.735 137.900 76.055 138.160 ;
        RECT 77.205 138.145 77.345 138.300 ;
        RECT 93.690 138.300 96.295 138.440 ;
        RECT 93.690 138.255 93.980 138.300 ;
        RECT 95.975 138.240 96.295 138.300 ;
        RECT 96.525 138.300 97.675 138.440 ;
        RECT 76.210 137.915 76.500 138.145 ;
        RECT 77.130 137.915 77.420 138.145 ;
        RECT 71.225 137.620 73.895 137.760 ;
        RECT 74.815 137.760 75.135 137.820 ;
        RECT 76.285 137.760 76.425 137.915 ;
        RECT 81.715 137.900 82.035 138.160 ;
        RECT 84.950 138.100 85.240 138.145 ;
        RECT 85.395 138.100 85.715 138.160 ;
        RECT 84.950 137.960 85.715 138.100 ;
        RECT 84.950 137.915 85.240 137.960 ;
        RECT 85.395 137.900 85.715 137.960 ;
        RECT 86.330 137.915 86.620 138.145 ;
        RECT 74.815 137.620 76.425 137.760 ;
        RECT 80.810 137.760 81.100 137.805 ;
        RECT 81.255 137.760 81.575 137.820 ;
        RECT 86.405 137.760 86.545 137.915 ;
        RECT 94.595 137.900 94.915 138.160 ;
        RECT 95.055 137.900 95.375 138.160 ;
        RECT 96.525 138.145 96.665 138.300 ;
        RECT 97.355 138.240 97.675 138.300 ;
        RECT 100.590 138.440 100.880 138.485 ;
        RECT 103.745 138.440 104.035 138.485 ;
        RECT 107.005 138.440 107.295 138.485 ;
        RECT 100.590 138.300 107.295 138.440 ;
        RECT 100.590 138.255 100.880 138.300 ;
        RECT 103.745 138.255 104.035 138.300 ;
        RECT 107.005 138.255 107.295 138.300 ;
        RECT 107.925 138.440 108.215 138.485 ;
        RECT 109.785 138.440 110.075 138.485 ;
        RECT 107.925 138.300 110.075 138.440 ;
        RECT 107.925 138.255 108.215 138.300 ;
        RECT 109.785 138.255 110.075 138.300 ;
        RECT 96.450 137.915 96.740 138.145 ;
        RECT 100.130 138.100 100.420 138.145 ;
        RECT 104.715 138.100 105.035 138.160 ;
        RECT 100.130 137.960 105.035 138.100 ;
        RECT 100.130 137.915 100.420 137.960 ;
        RECT 104.715 137.900 105.035 137.960 ;
        RECT 105.605 138.100 105.895 138.145 ;
        RECT 107.925 138.100 108.140 138.255 ;
        RECT 132.510 138.190 135.210 138.530 ;
        RECT 136.210 138.250 144.510 138.530 ;
        RECT 136.210 138.240 138.350 138.250 ;
        RECT 105.605 137.960 108.140 138.100 ;
        RECT 105.605 137.915 105.895 137.960 ;
        RECT 108.855 137.900 109.175 138.160 ;
        RECT 80.810 137.620 81.575 137.760 ;
        RECT 62.395 137.560 62.715 137.620 ;
        RECT 74.815 137.560 75.135 137.620 ;
        RECT 80.810 137.575 81.100 137.620 ;
        RECT 81.255 137.560 81.575 137.620 ;
        RECT 83.645 137.620 86.545 137.760 ;
        RECT 96.895 137.760 97.215 137.820 ;
        RECT 97.370 137.760 97.660 137.805 ;
        RECT 96.895 137.620 97.660 137.760 ;
        RECT 51.815 137.420 52.135 137.480 ;
        RECT 50.065 137.280 52.135 137.420 ;
        RECT 45.835 137.220 46.155 137.280 ;
        RECT 49.515 137.220 49.835 137.280 ;
        RECT 51.815 137.220 52.135 137.280 ;
        RECT 56.385 137.420 56.675 137.465 ;
        RECT 59.165 137.420 59.455 137.465 ;
        RECT 61.025 137.420 61.315 137.465 ;
        RECT 56.385 137.280 61.315 137.420 ;
        RECT 56.385 137.235 56.675 137.280 ;
        RECT 59.165 137.235 59.455 137.280 ;
        RECT 61.025 137.235 61.315 137.280 ;
        RECT 63.790 137.420 64.080 137.465 ;
        RECT 75.735 137.420 76.055 137.480 ;
        RECT 83.645 137.465 83.785 137.620 ;
        RECT 96.895 137.560 97.215 137.620 ;
        RECT 97.370 137.575 97.660 137.620 ;
        RECT 110.695 137.560 111.015 137.820 ;
        RECT 63.790 137.280 76.055 137.420 ;
        RECT 63.790 137.235 64.080 137.280 ;
        RECT 27.065 136.940 37.785 137.080 ;
        RECT 38.935 137.080 39.255 137.140 ;
        RECT 40.330 137.080 40.620 137.125 ;
        RECT 38.935 136.940 40.620 137.080 ;
        RECT 38.935 136.880 39.255 136.940 ;
        RECT 40.330 136.895 40.620 136.940 ;
        RECT 42.630 137.080 42.920 137.125 ;
        RECT 44.455 137.080 44.775 137.140 ;
        RECT 42.630 136.940 44.775 137.080 ;
        RECT 42.630 136.895 42.920 136.940 ;
        RECT 44.455 136.880 44.775 136.940 ;
        RECT 46.755 136.880 47.075 137.140 ;
        RECT 48.135 137.080 48.455 137.140 ;
        RECT 48.610 137.080 48.900 137.125 ;
        RECT 48.135 136.940 48.900 137.080 ;
        RECT 48.135 136.880 48.455 136.940 ;
        RECT 48.610 136.895 48.900 136.940 ;
        RECT 52.520 137.080 52.810 137.125 ;
        RECT 54.575 137.080 54.895 137.140 ;
        RECT 52.520 136.940 54.895 137.080 ;
        RECT 52.520 136.895 52.810 136.940 ;
        RECT 54.575 136.880 54.895 136.940 ;
        RECT 55.035 137.080 55.355 137.140 ;
        RECT 63.865 137.080 64.005 137.235 ;
        RECT 75.735 137.220 76.055 137.280 ;
        RECT 83.570 137.235 83.860 137.465 ;
        RECT 105.605 137.420 105.895 137.465 ;
        RECT 108.385 137.420 108.675 137.465 ;
        RECT 110.245 137.420 110.535 137.465 ;
        RECT 105.605 137.280 110.535 137.420 ;
        RECT 105.605 137.235 105.895 137.280 ;
        RECT 108.385 137.235 108.675 137.280 ;
        RECT 110.245 137.235 110.535 137.280 ;
        RECT 55.035 136.940 64.005 137.080 ;
        RECT 55.035 136.880 55.355 136.940 ;
        RECT 66.075 136.880 66.395 137.140 ;
        RECT 69.295 137.080 69.615 137.140 ;
        RECT 69.770 137.080 70.060 137.125 ;
        RECT 69.295 136.940 70.060 137.080 ;
        RECT 69.295 136.880 69.615 136.940 ;
        RECT 69.770 136.895 70.060 136.940 ;
        RECT 73.435 137.080 73.755 137.140 ;
        RECT 73.910 137.080 74.200 137.125 ;
        RECT 73.435 136.940 74.200 137.080 ;
        RECT 73.435 136.880 73.755 136.940 ;
        RECT 73.910 136.895 74.200 136.940 ;
        RECT 94.135 136.880 94.455 137.140 ;
        RECT 95.515 137.080 95.835 137.140 ;
        RECT 95.990 137.080 96.280 137.125 ;
        RECT 95.515 136.940 96.280 137.080 ;
        RECT 95.515 136.880 95.835 136.940 ;
        RECT 95.990 136.895 96.280 136.940 ;
        RECT 18.165 136.260 112.465 136.740 ;
        RECT 29.750 136.060 30.040 136.105 ;
        RECT 31.575 136.060 31.895 136.120 ;
        RECT 29.750 135.920 31.895 136.060 ;
        RECT 29.750 135.875 30.040 135.920 ;
        RECT 31.575 135.860 31.895 135.920 ;
        RECT 33.875 136.060 34.195 136.120 ;
        RECT 34.350 136.060 34.640 136.105 ;
        RECT 33.875 135.920 34.640 136.060 ;
        RECT 33.875 135.860 34.195 135.920 ;
        RECT 34.350 135.875 34.640 135.920 ;
        RECT 39.855 136.060 40.175 136.120 ;
        RECT 40.790 136.060 41.080 136.105 ;
        RECT 47.675 136.060 47.995 136.120 ;
        RECT 39.855 135.920 41.080 136.060 ;
        RECT 39.855 135.860 40.175 135.920 ;
        RECT 40.790 135.875 41.080 135.920 ;
        RECT 43.855 135.920 47.995 136.060 ;
        RECT 22.950 135.720 23.240 135.765 ;
        RECT 26.070 135.720 26.360 135.765 ;
        RECT 27.960 135.720 28.250 135.765 ;
        RECT 22.950 135.580 28.250 135.720 ;
        RECT 22.950 135.535 23.240 135.580 ;
        RECT 26.070 135.535 26.360 135.580 ;
        RECT 27.960 135.535 28.250 135.580 ;
        RECT 26.975 135.380 27.295 135.440 ;
        RECT 31.590 135.380 31.880 135.425 ;
        RECT 38.030 135.380 38.320 135.425 ;
        RECT 26.975 135.240 38.320 135.380 ;
        RECT 26.975 135.180 27.295 135.240 ;
        RECT 31.590 135.195 31.880 135.240 ;
        RECT 38.030 135.195 38.320 135.240 ;
        RECT 38.475 135.380 38.795 135.440 ;
        RECT 41.710 135.380 42.000 135.425 ;
        RECT 43.075 135.380 43.395 135.440 ;
        RECT 38.475 135.240 41.465 135.380 ;
        RECT 38.475 135.180 38.795 135.240 ;
        RECT 20.995 134.700 21.315 134.760 ;
        RECT 21.870 134.745 22.160 135.060 ;
        RECT 22.950 135.040 23.240 135.085 ;
        RECT 26.530 135.040 26.820 135.085 ;
        RECT 28.365 135.040 28.655 135.085 ;
        RECT 22.950 134.900 28.655 135.040 ;
        RECT 22.950 134.855 23.240 134.900 ;
        RECT 26.530 134.855 26.820 134.900 ;
        RECT 28.365 134.855 28.655 134.900 ;
        RECT 28.830 134.855 29.120 135.085 ;
        RECT 29.290 135.040 29.580 135.085 ;
        RECT 31.115 135.040 31.435 135.100 ;
        RECT 29.290 134.900 31.435 135.040 ;
        RECT 29.290 134.855 29.580 134.900 ;
        RECT 21.570 134.700 22.160 134.745 ;
        RECT 24.810 134.700 25.460 134.745 ;
        RECT 20.995 134.560 25.460 134.700 ;
        RECT 20.995 134.500 21.315 134.560 ;
        RECT 21.570 134.515 21.860 134.560 ;
        RECT 24.810 134.515 25.460 134.560 ;
        RECT 27.435 134.500 27.755 134.760 ;
        RECT 28.905 134.700 29.045 134.855 ;
        RECT 31.115 134.840 31.435 134.900 ;
        RECT 32.035 135.040 32.355 135.100 ;
        RECT 32.510 135.040 32.800 135.085 ;
        RECT 32.035 134.900 32.800 135.040 ;
        RECT 32.035 134.840 32.355 134.900 ;
        RECT 32.510 134.855 32.800 134.900 ;
        RECT 32.955 135.040 33.275 135.100 ;
        RECT 37.555 135.040 37.875 135.100 ;
        RECT 32.955 134.900 37.875 135.040 ;
        RECT 32.955 134.840 33.275 134.900 ;
        RECT 37.555 134.840 37.875 134.900 ;
        RECT 40.790 134.855 41.080 135.085 ;
        RECT 34.335 134.700 34.655 134.760 ;
        RECT 37.110 134.700 37.400 134.745 ;
        RECT 38.475 134.700 38.795 134.760 ;
        RECT 40.865 134.700 41.005 134.855 ;
        RECT 28.905 134.560 34.655 134.700 ;
        RECT 34.335 134.500 34.655 134.560 ;
        RECT 34.885 134.560 38.795 134.700 ;
        RECT 20.075 134.160 20.395 134.420 ;
        RECT 32.050 134.360 32.340 134.405 ;
        RECT 34.885 134.360 35.025 134.560 ;
        RECT 37.110 134.515 37.400 134.560 ;
        RECT 38.475 134.500 38.795 134.560 ;
        RECT 39.025 134.560 41.005 134.700 ;
        RECT 41.325 134.700 41.465 135.240 ;
        RECT 41.710 135.240 43.395 135.380 ;
        RECT 41.710 135.195 42.000 135.240 ;
        RECT 43.075 135.180 43.395 135.240 ;
        RECT 42.155 134.840 42.475 135.100 ;
        RECT 43.855 135.085 43.995 135.920 ;
        RECT 47.675 135.860 47.995 135.920 ;
        RECT 55.495 135.860 55.815 136.120 ;
        RECT 59.635 136.060 59.955 136.120 ;
        RECT 61.950 136.060 62.240 136.105 ;
        RECT 59.635 135.920 62.240 136.060 ;
        RECT 59.635 135.860 59.955 135.920 ;
        RECT 61.950 135.875 62.240 135.920 ;
        RECT 73.910 136.060 74.200 136.105 ;
        RECT 78.495 136.060 78.815 136.120 ;
        RECT 73.910 135.920 78.815 136.060 ;
        RECT 73.910 135.875 74.200 135.920 ;
        RECT 78.495 135.860 78.815 135.920 ;
        RECT 91.925 135.920 101.495 136.060 ;
        RECT 45.375 135.520 45.695 135.780 ;
        RECT 50.435 135.720 50.755 135.780 ;
        RECT 53.655 135.720 53.975 135.780 ;
        RECT 55.035 135.720 55.355 135.780 ;
        RECT 66.075 135.720 66.395 135.780 ;
        RECT 78.035 135.720 78.355 135.780 ;
        RECT 50.435 135.580 55.355 135.720 ;
        RECT 50.435 135.520 50.755 135.580 ;
        RECT 45.465 135.380 45.605 135.520 ;
        RECT 51.355 135.380 51.675 135.440 ;
        RECT 44.545 135.240 51.675 135.380 ;
        RECT 44.545 135.085 44.685 135.240 ;
        RECT 43.780 134.855 44.070 135.085 ;
        RECT 44.470 134.855 44.760 135.085 ;
        RECT 44.930 134.855 45.220 135.085 ;
        RECT 45.005 134.700 45.145 134.855 ;
        RECT 45.835 134.840 46.155 135.100 ;
        RECT 47.675 134.840 47.995 135.100 ;
        RECT 48.225 135.085 48.365 135.240 ;
        RECT 51.355 135.180 51.675 135.240 ;
        RECT 48.150 134.855 48.440 135.085 ;
        RECT 48.610 135.040 48.900 135.085 ;
        RECT 49.055 135.040 49.375 135.100 ;
        RECT 48.610 134.900 49.375 135.040 ;
        RECT 48.610 134.855 48.900 134.900 ;
        RECT 49.055 134.840 49.375 134.900 ;
        RECT 49.515 135.040 49.835 135.100 ;
        RECT 50.895 135.040 51.215 135.100 ;
        RECT 49.515 134.900 51.215 135.040 ;
        RECT 49.515 134.840 49.835 134.900 ;
        RECT 50.895 134.840 51.215 134.900 ;
        RECT 51.815 134.840 52.135 135.100 ;
        RECT 52.365 135.085 52.505 135.580 ;
        RECT 53.655 135.520 53.975 135.580 ;
        RECT 55.035 135.520 55.355 135.580 ;
        RECT 55.585 135.580 78.355 135.720 ;
        RECT 54.115 135.380 54.435 135.440 ;
        RECT 55.585 135.380 55.725 135.580 ;
        RECT 66.075 135.520 66.395 135.580 ;
        RECT 78.035 135.520 78.355 135.580 ;
        RECT 52.825 135.240 54.435 135.380 ;
        RECT 52.825 135.085 52.965 135.240 ;
        RECT 54.115 135.180 54.435 135.240 ;
        RECT 54.665 135.240 55.725 135.380 ;
        RECT 52.290 134.855 52.580 135.085 ;
        RECT 52.750 134.855 53.040 135.085 ;
        RECT 53.195 135.040 53.515 135.100 ;
        RECT 53.670 135.040 53.960 135.085 ;
        RECT 54.665 135.040 54.805 135.240 ;
        RECT 56.875 135.180 57.195 135.440 ;
        RECT 63.775 135.380 64.095 135.440 ;
        RECT 73.450 135.380 73.740 135.425 ;
        RECT 73.895 135.380 74.215 135.440 ;
        RECT 80.795 135.380 81.115 135.440 ;
        RECT 63.775 135.240 66.765 135.380 ;
        RECT 63.775 135.180 64.095 135.240 ;
        RECT 53.195 134.900 54.805 135.040 ;
        RECT 53.195 134.840 53.515 134.900 ;
        RECT 53.670 134.855 53.960 134.900 ;
        RECT 55.035 134.840 55.355 135.100 ;
        RECT 57.795 135.040 58.115 135.100 ;
        RECT 58.270 135.040 58.560 135.085 ;
        RECT 62.870 135.040 63.160 135.085 ;
        RECT 57.795 134.900 58.560 135.040 ;
        RECT 57.795 134.840 58.115 134.900 ;
        RECT 58.270 134.855 58.560 134.900 ;
        RECT 61.565 134.900 63.160 135.040 ;
        RECT 41.325 134.560 45.145 134.700 ;
        RECT 32.050 134.220 35.025 134.360 ;
        RECT 32.050 134.175 32.340 134.220 ;
        RECT 35.255 134.160 35.575 134.420 ;
        RECT 36.635 134.360 36.955 134.420 ;
        RECT 39.025 134.360 39.165 134.560 ;
        RECT 36.635 134.220 39.165 134.360 ;
        RECT 39.870 134.360 40.160 134.405 ;
        RECT 41.695 134.360 42.015 134.420 ;
        RECT 39.870 134.220 42.015 134.360 ;
        RECT 36.635 134.160 36.955 134.220 ;
        RECT 39.870 134.175 40.160 134.220 ;
        RECT 41.695 134.160 42.015 134.220 ;
        RECT 42.630 134.360 42.920 134.405 ;
        RECT 43.535 134.360 43.855 134.420 ;
        RECT 42.630 134.220 43.855 134.360 ;
        RECT 42.630 134.175 42.920 134.220 ;
        RECT 43.535 134.160 43.855 134.220 ;
        RECT 44.915 134.360 45.235 134.420 ;
        RECT 45.835 134.360 46.155 134.420 ;
        RECT 44.915 134.220 46.155 134.360 ;
        RECT 44.915 134.160 45.235 134.220 ;
        RECT 45.835 134.160 46.155 134.220 ;
        RECT 46.310 134.360 46.600 134.405 ;
        RECT 47.675 134.360 47.995 134.420 ;
        RECT 46.310 134.220 47.995 134.360 ;
        RECT 46.310 134.175 46.600 134.220 ;
        RECT 47.675 134.160 47.995 134.220 ;
        RECT 50.435 134.160 50.755 134.420 ;
        RECT 57.795 134.160 58.115 134.420 ;
        RECT 60.110 134.360 60.400 134.405 ;
        RECT 61.565 134.360 61.705 134.900 ;
        RECT 62.870 134.855 63.160 134.900 ;
        RECT 64.235 134.840 64.555 135.100 ;
        RECT 66.625 135.085 66.765 135.240 ;
        RECT 73.450 135.240 74.215 135.380 ;
        RECT 73.450 135.195 73.740 135.240 ;
        RECT 73.895 135.180 74.215 135.240 ;
        RECT 76.745 135.240 81.115 135.380 ;
        RECT 64.710 134.855 65.000 135.085 ;
        RECT 66.550 134.855 66.840 135.085 ;
        RECT 69.755 135.040 70.075 135.100 ;
        RECT 72.530 135.040 72.820 135.085 ;
        RECT 75.750 135.040 76.040 135.085 ;
        RECT 69.755 134.900 72.820 135.040 ;
        RECT 62.395 134.700 62.715 134.760 ;
        RECT 64.785 134.700 64.925 134.855 ;
        RECT 69.755 134.840 70.075 134.900 ;
        RECT 72.530 134.855 72.820 134.900 ;
        RECT 73.065 134.900 76.040 135.040 ;
        RECT 73.065 134.760 73.205 134.900 ;
        RECT 75.750 134.855 76.040 134.900 ;
        RECT 76.195 134.840 76.515 135.100 ;
        RECT 76.745 135.085 76.885 135.240 ;
        RECT 80.795 135.180 81.115 135.240 ;
        RECT 81.255 135.380 81.575 135.440 ;
        RECT 82.635 135.380 82.955 135.440 ;
        RECT 91.925 135.425 92.065 135.920 ;
        RECT 96.525 135.425 96.665 135.920 ;
        RECT 101.355 135.720 101.495 135.920 ;
        RECT 101.955 135.720 102.275 135.780 ;
        RECT 103.335 135.720 103.655 135.780 ;
        RECT 101.355 135.580 103.655 135.720 ;
        RECT 101.955 135.520 102.275 135.580 ;
        RECT 103.335 135.520 103.655 135.580 ;
        RECT 105.145 135.720 105.435 135.765 ;
        RECT 107.925 135.720 108.215 135.765 ;
        RECT 109.785 135.720 110.075 135.765 ;
        RECT 105.145 135.580 110.075 135.720 ;
        RECT 105.145 135.535 105.435 135.580 ;
        RECT 107.925 135.535 108.215 135.580 ;
        RECT 109.785 135.535 110.075 135.580 ;
        RECT 91.850 135.380 92.140 135.425 ;
        RECT 81.255 135.240 92.140 135.380 ;
        RECT 81.255 135.180 81.575 135.240 ;
        RECT 82.635 135.180 82.955 135.240 ;
        RECT 91.850 135.195 92.140 135.240 ;
        RECT 96.450 135.195 96.740 135.425 ;
        RECT 101.280 135.380 101.570 135.425 ;
        RECT 102.875 135.380 103.195 135.440 ;
        RECT 101.280 135.240 103.195 135.380 ;
        RECT 101.280 135.195 101.570 135.240 ;
        RECT 76.670 134.855 76.960 135.085 ;
        RECT 77.590 135.040 77.880 135.085 ;
        RECT 78.035 135.040 78.355 135.100 ;
        RECT 84.950 135.040 85.240 135.085 ;
        RECT 77.590 134.900 78.355 135.040 ;
        RECT 77.590 134.855 77.880 134.900 ;
        RECT 78.035 134.840 78.355 134.900 ;
        RECT 84.105 134.900 85.240 135.040 ;
        RECT 62.395 134.560 64.925 134.700 ;
        RECT 62.395 134.500 62.715 134.560 ;
        RECT 72.975 134.500 73.295 134.760 ;
        RECT 73.910 134.700 74.200 134.745 ;
        RECT 74.370 134.700 74.660 134.745 ;
        RECT 73.910 134.560 74.660 134.700 ;
        RECT 73.910 134.515 74.200 134.560 ;
        RECT 74.370 134.515 74.660 134.560 ;
        RECT 80.795 134.700 81.115 134.760 ;
        RECT 82.190 134.700 82.480 134.745 ;
        RECT 80.795 134.560 82.480 134.700 ;
        RECT 80.795 134.500 81.115 134.560 ;
        RECT 82.190 134.515 82.480 134.560 ;
        RECT 60.110 134.220 61.705 134.360 ;
        RECT 63.315 134.360 63.635 134.420 ;
        RECT 63.790 134.360 64.080 134.405 ;
        RECT 63.315 134.220 64.080 134.360 ;
        RECT 60.110 134.175 60.400 134.220 ;
        RECT 63.315 134.160 63.635 134.220 ;
        RECT 63.790 134.175 64.080 134.220 ;
        RECT 65.630 134.360 65.920 134.405 ;
        RECT 66.535 134.360 66.855 134.420 ;
        RECT 65.630 134.220 66.855 134.360 ;
        RECT 65.630 134.175 65.920 134.220 ;
        RECT 66.535 134.160 66.855 134.220 ;
        RECT 67.470 134.360 67.760 134.405 ;
        RECT 70.215 134.360 70.535 134.420 ;
        RECT 67.470 134.220 70.535 134.360 ;
        RECT 67.470 134.175 67.760 134.220 ;
        RECT 70.215 134.160 70.535 134.220 ;
        RECT 71.595 134.160 71.915 134.420 ;
        RECT 81.715 134.160 82.035 134.420 ;
        RECT 84.105 134.405 84.245 134.900 ;
        RECT 84.950 134.855 85.240 134.900 ;
        RECT 85.395 135.040 85.715 135.100 ;
        RECT 90.010 135.040 90.300 135.085 ;
        RECT 91.375 135.040 91.695 135.100 ;
        RECT 85.395 134.900 91.695 135.040 ;
        RECT 85.395 134.840 85.715 134.900 ;
        RECT 90.010 134.855 90.300 134.900 ;
        RECT 91.375 134.840 91.695 134.900 ;
        RECT 93.215 135.040 93.535 135.100 ;
        RECT 97.370 135.040 97.660 135.085 ;
        RECT 93.215 134.900 97.660 135.040 ;
        RECT 93.215 134.840 93.535 134.900 ;
        RECT 97.370 134.855 97.660 134.900 ;
        RECT 97.830 135.040 98.120 135.085 ;
        RECT 101.355 135.040 101.495 135.195 ;
        RECT 102.875 135.180 103.195 135.240 ;
        RECT 97.830 134.900 101.495 135.040 ;
        RECT 105.145 135.040 105.435 135.085 ;
        RECT 105.145 134.900 107.680 135.040 ;
        RECT 97.830 134.855 98.120 134.900 ;
        RECT 105.145 134.855 105.435 134.900 ;
        RECT 86.315 134.700 86.635 134.760 ;
        RECT 106.555 134.745 106.875 134.760 ;
        RECT 92.770 134.700 93.060 134.745 ;
        RECT 86.315 134.560 93.060 134.700 ;
        RECT 86.315 134.500 86.635 134.560 ;
        RECT 92.770 134.515 93.060 134.560 ;
        RECT 103.285 134.700 103.575 134.745 ;
        RECT 106.545 134.700 106.875 134.745 ;
        RECT 103.285 134.560 106.875 134.700 ;
        RECT 103.285 134.515 103.575 134.560 ;
        RECT 106.545 134.515 106.875 134.560 ;
        RECT 107.465 134.745 107.680 134.900 ;
        RECT 108.395 134.840 108.715 135.100 ;
        RECT 108.855 135.040 109.175 135.100 ;
        RECT 110.250 135.040 110.540 135.085 ;
        RECT 110.695 135.040 111.015 135.100 ;
        RECT 108.855 134.900 111.015 135.040 ;
        RECT 108.855 134.840 109.175 134.900 ;
        RECT 110.250 134.855 110.540 134.900 ;
        RECT 110.695 134.840 111.015 134.900 ;
        RECT 107.465 134.700 107.755 134.745 ;
        RECT 109.325 134.700 109.615 134.745 ;
        RECT 107.465 134.560 109.615 134.700 ;
        RECT 107.465 134.515 107.755 134.560 ;
        RECT 109.325 134.515 109.615 134.560 ;
        RECT 106.555 134.500 106.875 134.515 ;
        RECT 135.660 134.480 136.800 134.510 ;
        RECT 84.030 134.175 84.320 134.405 ;
        RECT 85.870 134.360 86.160 134.405 ;
        RECT 86.775 134.360 87.095 134.420 ;
        RECT 85.870 134.220 87.095 134.360 ;
        RECT 85.870 134.175 86.160 134.220 ;
        RECT 86.775 134.160 87.095 134.220 ;
        RECT 90.455 134.160 90.775 134.420 ;
        RECT 95.070 134.360 95.360 134.405 ;
        RECT 98.735 134.360 99.055 134.420 ;
        RECT 95.070 134.220 99.055 134.360 ;
        RECT 95.070 134.175 95.360 134.220 ;
        RECT 98.735 134.160 99.055 134.220 ;
        RECT 99.195 134.360 99.515 134.420 ;
        RECT 99.670 134.360 99.960 134.405 ;
        RECT 99.195 134.220 99.960 134.360 ;
        RECT 99.195 134.160 99.515 134.220 ;
        RECT 99.670 134.175 99.960 134.220 ;
        RECT 17.370 133.540 112.465 134.020 ;
        RECT 135.590 133.400 136.850 134.480 ;
        RECT 25.610 133.340 25.900 133.385 ;
        RECT 26.515 133.340 26.835 133.400 ;
        RECT 32.495 133.340 32.815 133.400 ;
        RECT 34.810 133.340 35.100 133.385 ;
        RECT 25.610 133.200 32.815 133.340 ;
        RECT 25.610 133.155 25.900 133.200 ;
        RECT 26.515 133.140 26.835 133.200 ;
        RECT 32.495 133.140 32.815 133.200 ;
        RECT 33.045 133.200 35.100 133.340 ;
        RECT 33.045 133.045 33.185 133.200 ;
        RECT 34.810 133.155 35.100 133.200 ;
        RECT 39.855 133.140 40.175 133.400 ;
        RECT 42.630 133.340 42.920 133.385 ;
        RECT 43.075 133.340 43.395 133.400 ;
        RECT 42.630 133.200 43.395 133.340 ;
        RECT 42.630 133.155 42.920 133.200 ;
        RECT 43.075 133.140 43.395 133.200 ;
        RECT 57.350 133.340 57.640 133.385 ;
        RECT 57.795 133.340 58.115 133.400 ;
        RECT 57.350 133.200 58.115 133.340 ;
        RECT 57.350 133.155 57.640 133.200 ;
        RECT 57.795 133.140 58.115 133.200 ;
        RECT 59.190 133.340 59.480 133.385 ;
        RECT 62.395 133.340 62.715 133.400 ;
        RECT 59.190 133.200 62.715 133.340 ;
        RECT 59.190 133.155 59.480 133.200 ;
        RECT 62.395 133.140 62.715 133.200 ;
        RECT 89.780 133.340 90.070 133.385 ;
        RECT 93.215 133.340 93.535 133.400 ;
        RECT 100.130 133.340 100.420 133.385 ;
        RECT 89.780 133.200 93.535 133.340 ;
        RECT 89.780 133.155 90.070 133.200 ;
        RECT 93.215 133.140 93.535 133.200 ;
        RECT 95.605 133.200 100.420 133.340 ;
        RECT 23.310 133.000 23.600 133.045 ;
        RECT 27.090 133.000 27.380 133.045 ;
        RECT 30.330 133.000 30.980 133.045 ;
        RECT 23.310 132.860 30.980 133.000 ;
        RECT 23.310 132.815 23.600 132.860 ;
        RECT 27.090 132.815 27.680 132.860 ;
        RECT 30.330 132.815 30.980 132.860 ;
        RECT 32.970 132.815 33.260 133.045 ;
        RECT 37.095 133.000 37.415 133.060 ;
        RECT 48.135 133.000 48.455 133.060 ;
        RECT 37.095 132.860 41.925 133.000 ;
        RECT 22.835 132.460 23.155 132.720 ;
        RECT 24.215 132.460 24.535 132.720 ;
        RECT 27.390 132.500 27.680 132.815 ;
        RECT 37.095 132.800 37.415 132.860 ;
        RECT 28.470 132.660 28.760 132.705 ;
        RECT 32.050 132.660 32.340 132.705 ;
        RECT 33.885 132.660 34.175 132.705 ;
        RECT 28.470 132.520 34.175 132.660 ;
        RECT 28.470 132.475 28.760 132.520 ;
        RECT 32.050 132.475 32.340 132.520 ;
        RECT 33.885 132.475 34.175 132.520 ;
        RECT 35.255 132.660 35.575 132.720 ;
        RECT 35.730 132.660 36.020 132.705 ;
        RECT 35.255 132.520 36.020 132.660 ;
        RECT 35.255 132.460 35.575 132.520 ;
        RECT 35.730 132.475 36.020 132.520 ;
        RECT 38.475 132.660 38.795 132.720 ;
        RECT 41.785 132.705 41.925 132.860 ;
        RECT 45.925 132.860 48.455 133.000 ;
        RECT 38.950 132.660 39.240 132.705 ;
        RECT 38.475 132.520 39.240 132.660 ;
        RECT 38.475 132.460 38.795 132.520 ;
        RECT 38.950 132.475 39.240 132.520 ;
        RECT 40.330 132.475 40.620 132.705 ;
        RECT 41.710 132.475 42.000 132.705 ;
        RECT 42.155 132.660 42.475 132.720 ;
        RECT 43.995 132.660 44.315 132.720 ;
        RECT 42.155 132.520 44.315 132.660 ;
        RECT 34.335 132.120 34.655 132.380 ;
        RECT 38.030 132.135 38.320 132.365 ;
        RECT 25.150 131.980 25.440 132.025 ;
        RECT 27.435 131.980 27.755 132.040 ;
        RECT 25.150 131.840 27.755 131.980 ;
        RECT 25.150 131.795 25.440 131.840 ;
        RECT 27.435 131.780 27.755 131.840 ;
        RECT 28.470 131.980 28.760 132.025 ;
        RECT 31.590 131.980 31.880 132.025 ;
        RECT 33.480 131.980 33.770 132.025 ;
        RECT 28.470 131.840 33.770 131.980 ;
        RECT 28.470 131.795 28.760 131.840 ;
        RECT 31.590 131.795 31.880 131.840 ;
        RECT 33.480 131.795 33.770 131.840 ;
        RECT 32.035 131.640 32.355 131.700 ;
        RECT 38.105 131.640 38.245 132.135 ;
        RECT 40.405 131.980 40.545 132.475 ;
        RECT 42.155 132.460 42.475 132.520 ;
        RECT 43.995 132.460 44.315 132.520 ;
        RECT 44.470 132.475 44.760 132.705 ;
        RECT 41.250 132.320 41.540 132.365 ;
        RECT 43.535 132.320 43.855 132.380 ;
        RECT 41.250 132.180 43.855 132.320 ;
        RECT 44.545 132.320 44.685 132.475 ;
        RECT 44.915 132.460 45.235 132.720 ;
        RECT 45.495 132.660 45.785 132.705 ;
        RECT 45.925 132.660 46.065 132.860 ;
        RECT 48.135 132.800 48.455 132.860 ;
        RECT 51.355 133.000 51.675 133.060 ;
        RECT 52.735 133.000 53.055 133.060 ;
        RECT 61.885 133.000 62.175 133.045 ;
        RECT 63.315 133.000 63.635 133.060 ;
        RECT 65.145 133.000 65.435 133.045 ;
        RECT 51.355 132.860 55.265 133.000 ;
        RECT 51.355 132.800 51.675 132.860 ;
        RECT 52.735 132.800 53.055 132.860 ;
        RECT 55.125 132.720 55.265 132.860 ;
        RECT 61.885 132.860 65.435 133.000 ;
        RECT 61.885 132.815 62.175 132.860 ;
        RECT 63.315 132.800 63.635 132.860 ;
        RECT 65.145 132.815 65.435 132.860 ;
        RECT 66.065 133.000 66.355 133.045 ;
        RECT 67.925 133.000 68.215 133.045 ;
        RECT 66.065 132.860 68.215 133.000 ;
        RECT 66.065 132.815 66.355 132.860 ;
        RECT 67.925 132.815 68.215 132.860 ;
        RECT 70.690 133.000 70.980 133.045 ;
        RECT 74.370 133.000 74.660 133.045 ;
        RECT 70.690 132.860 74.660 133.000 ;
        RECT 70.690 132.815 70.980 132.860 ;
        RECT 74.370 132.815 74.660 132.860 ;
        RECT 78.510 133.000 78.800 133.045 ;
        RECT 81.665 133.000 81.955 133.045 ;
        RECT 84.925 133.000 85.215 133.045 ;
        RECT 78.510 132.860 85.215 133.000 ;
        RECT 78.510 132.815 78.800 132.860 ;
        RECT 81.665 132.815 81.955 132.860 ;
        RECT 84.925 132.815 85.215 132.860 ;
        RECT 85.845 133.000 86.135 133.045 ;
        RECT 87.705 133.000 87.995 133.045 ;
        RECT 85.845 132.860 87.995 133.000 ;
        RECT 85.845 132.815 86.135 132.860 ;
        RECT 87.705 132.815 87.995 132.860 ;
        RECT 91.785 133.000 92.075 133.045 ;
        RECT 95.045 133.000 95.335 133.045 ;
        RECT 95.605 133.000 95.745 133.200 ;
        RECT 100.130 133.155 100.420 133.200 ;
        RECT 102.875 133.140 103.195 133.400 ;
        RECT 107.490 133.340 107.780 133.385 ;
        RECT 108.395 133.340 108.715 133.400 ;
        RECT 107.490 133.200 108.715 133.340 ;
        RECT 107.490 133.155 107.780 133.200 ;
        RECT 108.395 133.140 108.715 133.200 ;
        RECT 91.785 132.860 95.745 133.000 ;
        RECT 95.965 133.000 96.255 133.045 ;
        RECT 97.825 133.000 98.115 133.045 ;
        RECT 108.855 133.000 109.175 133.060 ;
        RECT 95.965 132.860 98.115 133.000 ;
        RECT 91.785 132.815 92.075 132.860 ;
        RECT 95.045 132.815 95.335 132.860 ;
        RECT 95.965 132.815 96.255 132.860 ;
        RECT 97.825 132.815 98.115 132.860 ;
        RECT 101.355 132.860 109.175 133.000 ;
        RECT 45.495 132.520 46.065 132.660 ;
        RECT 46.310 132.660 46.600 132.705 ;
        RECT 50.895 132.660 51.215 132.720 ;
        RECT 46.310 132.520 51.215 132.660 ;
        RECT 45.495 132.475 45.785 132.520 ;
        RECT 46.310 132.475 46.600 132.520 ;
        RECT 50.895 132.460 51.215 132.520 ;
        RECT 53.210 132.475 53.500 132.705 ;
        RECT 47.215 132.320 47.535 132.380 ;
        RECT 44.545 132.180 47.535 132.320 ;
        RECT 41.250 132.135 41.540 132.180 ;
        RECT 43.535 132.120 43.855 132.180 ;
        RECT 47.215 132.120 47.535 132.180 ;
        RECT 49.515 132.320 49.835 132.380 ;
        RECT 52.275 132.320 52.595 132.380 ;
        RECT 53.285 132.320 53.425 132.475 ;
        RECT 53.655 132.460 53.975 132.720 ;
        RECT 54.130 132.660 54.420 132.705 ;
        RECT 54.130 132.520 54.805 132.660 ;
        RECT 54.130 132.475 54.420 132.520 ;
        RECT 49.515 132.180 53.425 132.320 ;
        RECT 49.515 132.120 49.835 132.180 ;
        RECT 52.275 132.120 52.595 132.180 ;
        RECT 50.435 131.980 50.755 132.040 ;
        RECT 40.405 131.840 50.755 131.980 ;
        RECT 50.435 131.780 50.755 131.840 ;
        RECT 50.895 131.980 51.215 132.040 ;
        RECT 53.745 131.980 53.885 132.460 ;
        RECT 50.895 131.840 53.885 131.980 ;
        RECT 54.665 131.980 54.805 132.520 ;
        RECT 55.035 132.460 55.355 132.720 ;
        RECT 63.745 132.660 64.035 132.705 ;
        RECT 66.065 132.660 66.280 132.815 ;
        RECT 63.745 132.520 66.280 132.660 ;
        RECT 66.535 132.660 66.855 132.720 ;
        RECT 67.010 132.660 67.300 132.705 ;
        RECT 70.230 132.660 70.520 132.705 ;
        RECT 66.535 132.520 67.300 132.660 ;
        RECT 63.745 132.475 64.035 132.520 ;
        RECT 66.535 132.460 66.855 132.520 ;
        RECT 67.010 132.475 67.300 132.520 ;
        RECT 67.545 132.520 70.520 132.660 ;
        RECT 56.415 132.120 56.735 132.380 ;
        RECT 56.890 132.320 57.180 132.365 ;
        RECT 60.555 132.320 60.875 132.380 ;
        RECT 67.545 132.320 67.685 132.520 ;
        RECT 70.230 132.475 70.520 132.520 ;
        RECT 72.055 132.460 72.375 132.720 ;
        RECT 72.975 132.660 73.295 132.720 ;
        RECT 75.750 132.660 76.040 132.705 ;
        RECT 72.975 132.520 76.040 132.660 ;
        RECT 72.975 132.460 73.295 132.520 ;
        RECT 56.890 132.180 58.485 132.320 ;
        RECT 56.890 132.135 57.180 132.180 ;
        RECT 56.965 131.980 57.105 132.135 ;
        RECT 54.665 131.840 57.105 131.980 ;
        RECT 50.895 131.780 51.215 131.840 ;
        RECT 58.345 131.700 58.485 132.180 ;
        RECT 60.555 132.180 67.685 132.320 ;
        RECT 60.555 132.120 60.875 132.180 ;
        RECT 68.835 132.120 69.155 132.380 ;
        RECT 71.610 132.320 71.900 132.365 ;
        RECT 73.435 132.320 73.755 132.380 ;
        RECT 71.610 132.180 73.755 132.320 ;
        RECT 71.610 132.135 71.900 132.180 ;
        RECT 73.435 132.120 73.755 132.180 ;
        RECT 63.745 131.980 64.035 132.025 ;
        RECT 66.525 131.980 66.815 132.025 ;
        RECT 68.385 131.980 68.675 132.025 ;
        RECT 71.135 131.980 71.455 132.040 ;
        RECT 73.985 131.980 74.125 132.520 ;
        RECT 75.750 132.475 76.040 132.520 ;
        RECT 76.195 132.460 76.515 132.720 ;
        RECT 76.670 132.475 76.960 132.705 ;
        RECT 77.590 132.660 77.880 132.705 ;
        RECT 78.035 132.660 78.355 132.720 ;
        RECT 77.590 132.520 78.355 132.660 ;
        RECT 77.590 132.475 77.880 132.520 ;
        RECT 74.815 132.320 75.135 132.380 ;
        RECT 76.285 132.320 76.425 132.460 ;
        RECT 74.815 132.180 76.425 132.320 ;
        RECT 74.815 132.120 75.135 132.180 ;
        RECT 63.745 131.840 68.675 131.980 ;
        RECT 63.745 131.795 64.035 131.840 ;
        RECT 66.525 131.795 66.815 131.840 ;
        RECT 68.385 131.795 68.675 131.840 ;
        RECT 68.925 131.840 70.905 131.980 ;
        RECT 32.035 131.500 38.245 131.640 ;
        RECT 32.035 131.440 32.355 131.500 ;
        RECT 40.315 131.440 40.635 131.700 ;
        RECT 41.695 131.640 42.015 131.700 ;
        RECT 43.090 131.640 43.380 131.685 ;
        RECT 41.695 131.500 43.380 131.640 ;
        RECT 41.695 131.440 42.015 131.500 ;
        RECT 43.090 131.455 43.380 131.500 ;
        RECT 43.535 131.640 43.855 131.700 ;
        RECT 44.915 131.640 45.235 131.700 ;
        RECT 43.535 131.500 45.235 131.640 ;
        RECT 43.535 131.440 43.855 131.500 ;
        RECT 44.915 131.440 45.235 131.500 ;
        RECT 45.375 131.640 45.695 131.700 ;
        RECT 51.830 131.640 52.120 131.685 ;
        RECT 45.375 131.500 52.120 131.640 ;
        RECT 45.375 131.440 45.695 131.500 ;
        RECT 51.830 131.455 52.120 131.500 ;
        RECT 58.255 131.640 58.575 131.700 ;
        RECT 59.880 131.640 60.170 131.685 ;
        RECT 58.255 131.500 60.170 131.640 ;
        RECT 58.255 131.440 58.575 131.500 ;
        RECT 59.880 131.455 60.170 131.500 ;
        RECT 63.315 131.640 63.635 131.700 ;
        RECT 68.925 131.640 69.065 131.840 ;
        RECT 63.315 131.500 69.065 131.640 ;
        RECT 69.310 131.640 69.600 131.685 ;
        RECT 69.755 131.640 70.075 131.700 ;
        RECT 70.765 131.685 70.905 131.840 ;
        RECT 71.135 131.840 74.125 131.980 ;
        RECT 76.745 131.980 76.885 132.475 ;
        RECT 78.035 132.460 78.355 132.520 ;
        RECT 78.970 132.475 79.260 132.705 ;
        RECT 83.525 132.660 83.815 132.705 ;
        RECT 85.845 132.660 86.060 132.815 ;
        RECT 83.525 132.520 86.060 132.660 ;
        RECT 83.525 132.475 83.815 132.520 ;
        RECT 79.045 132.320 79.185 132.475 ;
        RECT 86.775 132.460 87.095 132.720 ;
        RECT 87.235 132.660 87.555 132.720 ;
        RECT 88.630 132.660 88.920 132.705 ;
        RECT 87.235 132.520 88.920 132.660 ;
        RECT 87.235 132.460 87.555 132.520 ;
        RECT 88.630 132.475 88.920 132.520 ;
        RECT 93.645 132.660 93.935 132.705 ;
        RECT 95.965 132.660 96.180 132.815 ;
        RECT 93.645 132.520 96.180 132.660 ;
        RECT 96.910 132.660 97.200 132.705 ;
        RECT 98.275 132.660 98.595 132.720 ;
        RECT 96.910 132.520 98.595 132.660 ;
        RECT 93.645 132.475 93.935 132.520 ;
        RECT 96.910 132.475 97.200 132.520 ;
        RECT 98.275 132.460 98.595 132.520 ;
        RECT 100.575 132.460 100.895 132.720 ;
        RECT 85.395 132.320 85.715 132.380 ;
        RECT 79.045 132.180 85.715 132.320 ;
        RECT 85.395 132.120 85.715 132.180 ;
        RECT 97.355 132.320 97.675 132.380 ;
        RECT 98.750 132.320 99.040 132.365 ;
        RECT 101.355 132.320 101.495 132.860 ;
        RECT 108.855 132.800 109.175 132.860 ;
        RECT 102.875 132.660 103.195 132.720 ;
        RECT 103.350 132.660 103.640 132.705 ;
        RECT 106.570 132.660 106.860 132.705 ;
        RECT 102.875 132.520 103.640 132.660 ;
        RECT 102.875 132.460 103.195 132.520 ;
        RECT 103.350 132.475 103.640 132.520 ;
        RECT 105.265 132.520 106.860 132.660 ;
        RECT 97.355 132.180 101.495 132.320 ;
        RECT 97.355 132.120 97.675 132.180 ;
        RECT 98.750 132.135 99.040 132.180 ;
        RECT 101.955 132.120 102.275 132.380 ;
        RECT 79.660 131.980 79.950 132.025 ;
        RECT 81.715 131.980 82.035 132.040 ;
        RECT 105.265 132.025 105.405 132.520 ;
        RECT 106.570 132.475 106.860 132.520 ;
        RECT 76.745 131.840 82.035 131.980 ;
        RECT 71.135 131.780 71.455 131.840 ;
        RECT 79.660 131.795 79.950 131.840 ;
        RECT 81.715 131.780 82.035 131.840 ;
        RECT 83.525 131.980 83.815 132.025 ;
        RECT 86.305 131.980 86.595 132.025 ;
        RECT 88.165 131.980 88.455 132.025 ;
        RECT 83.525 131.840 88.455 131.980 ;
        RECT 83.525 131.795 83.815 131.840 ;
        RECT 86.305 131.795 86.595 131.840 ;
        RECT 88.165 131.795 88.455 131.840 ;
        RECT 93.645 131.980 93.935 132.025 ;
        RECT 96.425 131.980 96.715 132.025 ;
        RECT 98.285 131.980 98.575 132.025 ;
        RECT 93.645 131.840 98.575 131.980 ;
        RECT 93.645 131.795 93.935 131.840 ;
        RECT 96.425 131.795 96.715 131.840 ;
        RECT 98.285 131.795 98.575 131.840 ;
        RECT 105.190 131.795 105.480 132.025 ;
        RECT 69.310 131.500 70.075 131.640 ;
        RECT 63.315 131.440 63.635 131.500 ;
        RECT 69.310 131.455 69.600 131.500 ;
        RECT 69.755 131.440 70.075 131.500 ;
        RECT 70.690 131.455 70.980 131.685 ;
        RECT 72.990 131.640 73.280 131.685 ;
        RECT 74.355 131.640 74.675 131.700 ;
        RECT 72.990 131.500 74.675 131.640 ;
        RECT 72.990 131.455 73.280 131.500 ;
        RECT 74.355 131.440 74.675 131.500 ;
        RECT 91.375 131.640 91.695 131.700 ;
        RECT 96.895 131.640 97.215 131.700 ;
        RECT 100.575 131.640 100.895 131.700 ;
        RECT 105.635 131.640 105.955 131.700 ;
        RECT 91.375 131.500 105.955 131.640 ;
        RECT 91.375 131.440 91.695 131.500 ;
        RECT 96.895 131.440 97.215 131.500 ;
        RECT 100.575 131.440 100.895 131.500 ;
        RECT 105.635 131.440 105.955 131.500 ;
        RECT 18.165 130.820 112.465 131.300 ;
        RECT 24.215 130.620 24.535 130.680 ;
        RECT 24.690 130.620 24.980 130.665 ;
        RECT 24.215 130.480 24.980 130.620 ;
        RECT 24.215 130.420 24.535 130.480 ;
        RECT 24.690 130.435 24.980 130.480 ;
        RECT 38.950 130.620 39.240 130.665 ;
        RECT 40.315 130.620 40.635 130.680 ;
        RECT 38.950 130.480 40.635 130.620 ;
        RECT 38.950 130.435 39.240 130.480 ;
        RECT 40.315 130.420 40.635 130.480 ;
        RECT 40.790 130.435 41.080 130.665 ;
        RECT 22.850 130.280 23.140 130.325 ;
        RECT 25.595 130.280 25.915 130.340 ;
        RECT 22.850 130.140 25.915 130.280 ;
        RECT 22.850 130.095 23.140 130.140 ;
        RECT 25.595 130.080 25.915 130.140 ;
        RECT 37.555 130.280 37.875 130.340 ;
        RECT 40.865 130.280 41.005 130.435 ;
        RECT 43.535 130.420 43.855 130.680 ;
        RECT 45.375 130.620 45.695 130.680 ;
        RECT 44.085 130.480 45.695 130.620 ;
        RECT 44.085 130.280 44.225 130.480 ;
        RECT 45.375 130.420 45.695 130.480 ;
        RECT 46.770 130.435 47.060 130.665 ;
        RECT 52.275 130.620 52.595 130.680 ;
        RECT 60.110 130.620 60.400 130.665 ;
        RECT 60.555 130.620 60.875 130.680 ;
        RECT 68.375 130.620 68.695 130.680 ;
        RECT 71.135 130.620 71.455 130.680 ;
        RECT 52.275 130.480 53.425 130.620 ;
        RECT 37.555 130.140 41.005 130.280 ;
        RECT 42.245 130.140 44.225 130.280 ;
        RECT 46.845 130.280 46.985 130.435 ;
        RECT 52.275 130.420 52.595 130.480 ;
        RECT 47.215 130.280 47.535 130.340 ;
        RECT 46.845 130.140 47.535 130.280 ;
        RECT 37.555 130.080 37.875 130.140 ;
        RECT 20.075 129.940 20.395 130.000 ;
        RECT 26.975 129.940 27.295 130.000 ;
        RECT 20.075 129.800 27.295 129.940 ;
        RECT 20.075 129.740 20.395 129.800 ;
        RECT 26.975 129.740 27.295 129.800 ;
        RECT 27.435 129.740 27.755 130.000 ;
        RECT 40.330 129.940 40.620 129.985 ;
        RECT 41.695 129.940 42.015 130.000 ;
        RECT 40.330 129.800 42.015 129.940 ;
        RECT 40.330 129.755 40.620 129.800 ;
        RECT 41.695 129.740 42.015 129.800 ;
        RECT 21.455 129.600 21.775 129.660 ;
        RECT 31.130 129.600 31.420 129.645 ;
        RECT 21.455 129.460 31.420 129.600 ;
        RECT 21.455 129.400 21.775 129.460 ;
        RECT 31.130 129.415 31.420 129.460 ;
        RECT 36.635 129.400 36.955 129.660 ;
        RECT 37.110 129.415 37.400 129.645 ;
        RECT 38.030 129.600 38.320 129.645 ;
        RECT 38.475 129.600 38.795 129.660 ;
        RECT 38.030 129.460 40.545 129.600 ;
        RECT 38.030 129.415 38.320 129.460 ;
        RECT 22.835 129.260 23.155 129.320 ;
        RECT 37.185 129.260 37.325 129.415 ;
        RECT 22.835 129.120 37.325 129.260 ;
        RECT 22.835 129.060 23.155 129.120 ;
        RECT 26.515 128.720 26.835 128.980 ;
        RECT 28.815 128.920 29.135 128.980 ;
        RECT 30.670 128.920 30.960 128.965 ;
        RECT 28.815 128.780 30.960 128.920 ;
        RECT 28.815 128.720 29.135 128.780 ;
        RECT 30.670 128.735 30.960 128.780 ;
        RECT 32.495 128.920 32.815 128.980 ;
        RECT 35.730 128.920 36.020 128.965 ;
        RECT 32.495 128.780 36.020 128.920 ;
        RECT 32.495 128.720 32.815 128.780 ;
        RECT 35.730 128.735 36.020 128.780 ;
        RECT 37.095 128.920 37.415 128.980 ;
        RECT 38.105 128.920 38.245 129.415 ;
        RECT 38.475 129.400 38.795 129.460 ;
        RECT 39.410 129.260 39.700 129.305 ;
        RECT 39.855 129.260 40.175 129.320 ;
        RECT 39.410 129.120 40.175 129.260 ;
        RECT 40.405 129.260 40.545 129.460 ;
        RECT 40.775 129.400 41.095 129.660 ;
        RECT 42.245 129.645 42.385 130.140 ;
        RECT 47.215 130.080 47.535 130.140 ;
        RECT 53.285 130.280 53.425 130.480 ;
        RECT 60.110 130.480 60.875 130.620 ;
        RECT 60.110 130.435 60.400 130.480 ;
        RECT 60.555 130.420 60.875 130.480 ;
        RECT 64.785 130.480 71.455 130.620 ;
        RECT 64.785 130.280 64.925 130.480 ;
        RECT 68.375 130.420 68.695 130.480 ;
        RECT 71.135 130.420 71.455 130.480 ;
        RECT 98.275 130.620 98.595 130.680 ;
        RECT 99.670 130.620 99.960 130.665 ;
        RECT 98.275 130.480 99.960 130.620 ;
        RECT 98.275 130.420 98.595 130.480 ;
        RECT 99.670 130.435 99.960 130.480 ;
        RECT 53.285 130.140 64.925 130.280 ;
        RECT 65.125 130.280 65.415 130.325 ;
        RECT 67.905 130.280 68.195 130.325 ;
        RECT 69.765 130.280 70.055 130.325 ;
        RECT 65.125 130.140 70.055 130.280 ;
        RECT 43.090 129.940 43.380 129.985 ;
        RECT 43.090 129.800 45.605 129.940 ;
        RECT 43.090 129.755 43.380 129.800 ;
        RECT 42.170 129.415 42.460 129.645 ;
        RECT 43.550 129.600 43.840 129.645 ;
        RECT 43.995 129.600 44.315 129.660 ;
        RECT 43.550 129.460 44.315 129.600 ;
        RECT 43.550 129.415 43.840 129.460 ;
        RECT 43.995 129.400 44.315 129.460 ;
        RECT 40.405 129.120 43.765 129.260 ;
        RECT 39.410 129.075 39.700 129.120 ;
        RECT 39.855 129.060 40.175 129.120 ;
        RECT 43.625 128.980 43.765 129.120 ;
        RECT 37.095 128.780 38.245 128.920 ;
        RECT 40.315 128.920 40.635 128.980 ;
        RECT 41.710 128.920 42.000 128.965 ;
        RECT 40.315 128.780 42.000 128.920 ;
        RECT 37.095 128.720 37.415 128.780 ;
        RECT 40.315 128.720 40.635 128.780 ;
        RECT 41.710 128.735 42.000 128.780 ;
        RECT 43.535 128.720 43.855 128.980 ;
        RECT 43.995 128.920 44.315 128.980 ;
        RECT 44.470 128.920 44.760 128.965 ;
        RECT 43.995 128.780 44.760 128.920 ;
        RECT 43.995 128.720 44.315 128.780 ;
        RECT 44.470 128.735 44.760 128.780 ;
        RECT 44.915 128.720 45.235 128.980 ;
        RECT 45.465 128.920 45.605 129.800 ;
        RECT 46.755 129.740 47.075 130.000 ;
        RECT 50.895 129.940 51.215 130.000 ;
        RECT 50.065 129.800 51.215 129.940 ;
        RECT 45.835 129.400 46.155 129.660 ;
        RECT 49.515 129.400 49.835 129.660 ;
        RECT 50.065 129.645 50.205 129.800 ;
        RECT 50.895 129.740 51.215 129.800 ;
        RECT 49.990 129.415 50.280 129.645 ;
        RECT 50.435 129.400 50.755 129.660 ;
        RECT 51.355 129.400 51.675 129.660 ;
        RECT 53.285 129.645 53.425 130.140 ;
        RECT 65.125 130.095 65.415 130.140 ;
        RECT 67.905 130.095 68.195 130.140 ;
        RECT 69.765 130.095 70.055 130.140 ;
        RECT 80.765 130.280 81.055 130.325 ;
        RECT 83.545 130.280 83.835 130.325 ;
        RECT 85.405 130.280 85.695 130.325 ;
        RECT 80.765 130.140 85.695 130.280 ;
        RECT 80.765 130.095 81.055 130.140 ;
        RECT 83.545 130.095 83.835 130.140 ;
        RECT 85.405 130.095 85.695 130.140 ;
        RECT 86.775 130.280 87.095 130.340 ;
        RECT 88.400 130.280 88.690 130.325 ;
        RECT 86.775 130.140 88.690 130.280 ;
        RECT 86.775 130.080 87.095 130.140 ;
        RECT 88.400 130.095 88.690 130.140 ;
        RECT 92.265 130.280 92.555 130.325 ;
        RECT 95.045 130.280 95.335 130.325 ;
        RECT 96.905 130.280 97.195 130.325 ;
        RECT 92.265 130.140 97.195 130.280 ;
        RECT 92.265 130.095 92.555 130.140 ;
        RECT 95.045 130.095 95.335 130.140 ;
        RECT 96.905 130.095 97.195 130.140 ;
        RECT 97.830 130.095 98.120 130.325 ;
        RECT 54.575 129.940 54.895 130.000 ;
        RECT 53.745 129.800 54.895 129.940 ;
        RECT 53.745 129.660 53.885 129.800 ;
        RECT 54.575 129.740 54.895 129.800 ;
        RECT 57.335 129.940 57.655 130.000 ;
        RECT 59.175 129.940 59.495 130.000 ;
        RECT 57.335 129.800 59.495 129.940 ;
        RECT 57.335 129.740 57.655 129.800 ;
        RECT 59.175 129.740 59.495 129.800 ;
        RECT 68.835 129.940 69.155 130.000 ;
        RECT 70.230 129.940 70.520 129.985 ;
        RECT 72.530 129.940 72.820 129.985 ;
        RECT 73.435 129.940 73.755 130.000 ;
        RECT 68.835 129.800 72.285 129.940 ;
        RECT 68.835 129.740 69.155 129.800 ;
        RECT 70.230 129.755 70.520 129.800 ;
        RECT 53.210 129.415 53.500 129.645 ;
        RECT 53.655 129.400 53.975 129.660 ;
        RECT 54.130 129.415 54.420 129.645 ;
        RECT 47.230 129.260 47.520 129.305 ;
        RECT 48.150 129.260 48.440 129.305 ;
        RECT 47.230 129.120 48.440 129.260 ;
        RECT 47.230 129.075 47.520 129.120 ;
        RECT 48.150 129.075 48.440 129.120 ;
        RECT 49.055 129.260 49.375 129.320 ;
        RECT 51.830 129.260 52.120 129.305 ;
        RECT 49.055 129.120 52.120 129.260 ;
        RECT 54.205 129.260 54.345 129.415 ;
        RECT 55.035 129.400 55.355 129.660 ;
        RECT 58.255 129.400 58.575 129.660 ;
        RECT 65.125 129.600 65.415 129.645 ;
        RECT 68.390 129.600 68.680 129.645 ;
        RECT 69.755 129.600 70.075 129.660 ;
        RECT 65.125 129.460 67.660 129.600 ;
        RECT 65.125 129.415 65.415 129.460 ;
        RECT 66.535 129.305 66.855 129.320 ;
        RECT 63.265 129.260 63.555 129.305 ;
        RECT 66.525 129.260 66.855 129.305 ;
        RECT 54.205 129.120 58.025 129.260 ;
        RECT 49.055 129.060 49.375 129.120 ;
        RECT 51.830 129.075 52.120 129.120 ;
        RECT 47.675 128.920 47.995 128.980 ;
        RECT 57.885 128.965 58.025 129.120 ;
        RECT 63.265 129.120 66.855 129.260 ;
        RECT 63.265 129.075 63.555 129.120 ;
        RECT 66.525 129.075 66.855 129.120 ;
        RECT 67.445 129.305 67.660 129.460 ;
        RECT 68.390 129.460 70.075 129.600 ;
        RECT 68.390 129.415 68.680 129.460 ;
        RECT 69.755 129.400 70.075 129.460 ;
        RECT 70.675 129.600 70.995 129.660 ;
        RECT 71.610 129.600 71.900 129.645 ;
        RECT 70.675 129.460 71.900 129.600 ;
        RECT 72.145 129.600 72.285 129.800 ;
        RECT 72.530 129.800 73.755 129.940 ;
        RECT 72.530 129.755 72.820 129.800 ;
        RECT 73.435 129.740 73.755 129.800 ;
        RECT 73.985 129.800 83.785 129.940 ;
        RECT 73.985 129.660 74.125 129.800 ;
        RECT 73.895 129.600 74.215 129.660 ;
        RECT 72.145 129.460 74.215 129.600 ;
        RECT 70.675 129.400 70.995 129.460 ;
        RECT 71.610 129.415 71.900 129.460 ;
        RECT 73.895 129.400 74.215 129.460 ;
        RECT 74.370 129.415 74.660 129.645 ;
        RECT 67.445 129.260 67.735 129.305 ;
        RECT 69.305 129.260 69.595 129.305 ;
        RECT 67.445 129.120 69.595 129.260 ;
        RECT 67.445 129.075 67.735 129.120 ;
        RECT 69.305 129.075 69.595 129.120 ;
        RECT 71.135 129.260 71.455 129.320 ;
        RECT 74.445 129.260 74.585 129.415 ;
        RECT 74.815 129.400 75.135 129.660 ;
        RECT 75.290 129.415 75.580 129.645 ;
        RECT 76.195 129.600 76.515 129.660 ;
        RECT 78.035 129.600 78.355 129.660 ;
        RECT 76.195 129.460 78.355 129.600 ;
        RECT 71.135 129.120 74.585 129.260 ;
        RECT 66.535 129.060 66.855 129.075 ;
        RECT 71.135 129.060 71.455 129.120 ;
        RECT 45.465 128.780 47.995 128.920 ;
        RECT 47.675 128.720 47.995 128.780 ;
        RECT 57.810 128.920 58.100 128.965 ;
        RECT 58.255 128.920 58.575 128.980 ;
        RECT 61.260 128.920 61.550 128.965 ;
        RECT 57.810 128.780 61.550 128.920 ;
        RECT 57.810 128.735 58.100 128.780 ;
        RECT 58.255 128.720 58.575 128.780 ;
        RECT 61.260 128.735 61.550 128.780 ;
        RECT 70.675 128.720 70.995 128.980 ;
        RECT 72.515 128.920 72.835 128.980 ;
        RECT 72.990 128.920 73.280 128.965 ;
        RECT 72.515 128.780 73.280 128.920 ;
        RECT 75.365 128.920 75.505 129.415 ;
        RECT 76.195 129.400 76.515 129.460 ;
        RECT 78.035 129.400 78.355 129.460 ;
        RECT 80.765 129.600 81.055 129.645 ;
        RECT 83.645 129.600 83.785 129.800 ;
        RECT 84.015 129.740 84.335 130.000 ;
        RECT 87.235 129.940 87.555 130.000 ;
        RECT 95.530 129.940 95.820 129.985 ;
        RECT 97.905 129.940 98.045 130.095 ;
        RECT 87.235 129.800 95.285 129.940 ;
        RECT 87.235 129.740 87.555 129.800 ;
        RECT 85.870 129.600 86.160 129.645 ;
        RECT 80.765 129.460 83.300 129.600 ;
        RECT 83.645 129.460 86.160 129.600 ;
        RECT 80.765 129.415 81.055 129.460 ;
        RECT 83.085 129.305 83.300 129.460 ;
        RECT 85.870 129.415 86.160 129.460 ;
        RECT 87.710 129.600 88.000 129.645 ;
        RECT 91.375 129.600 91.695 129.660 ;
        RECT 87.710 129.460 91.695 129.600 ;
        RECT 87.710 129.415 88.000 129.460 ;
        RECT 91.375 129.400 91.695 129.460 ;
        RECT 92.265 129.600 92.555 129.645 ;
        RECT 95.145 129.600 95.285 129.800 ;
        RECT 95.530 129.800 98.045 129.940 ;
        RECT 95.530 129.755 95.820 129.800 ;
        RECT 97.355 129.600 97.675 129.660 ;
        RECT 92.265 129.460 94.800 129.600 ;
        RECT 95.145 129.460 97.675 129.600 ;
        RECT 92.265 129.415 92.555 129.460 ;
        RECT 90.455 129.305 90.775 129.320 ;
        RECT 94.585 129.305 94.800 129.460 ;
        RECT 97.355 129.400 97.675 129.460 ;
        RECT 98.735 129.400 99.055 129.660 ;
        RECT 99.195 129.600 99.515 129.660 ;
        RECT 100.590 129.600 100.880 129.645 ;
        RECT 99.195 129.460 100.880 129.600 ;
        RECT 99.195 129.400 99.515 129.460 ;
        RECT 100.590 129.415 100.880 129.460 ;
        RECT 78.905 129.260 79.195 129.305 ;
        RECT 82.165 129.260 82.455 129.305 ;
        RECT 83.085 129.260 83.375 129.305 ;
        RECT 84.945 129.260 85.235 129.305 ;
        RECT 78.905 129.120 82.865 129.260 ;
        RECT 78.905 129.075 79.195 129.120 ;
        RECT 82.165 129.075 82.455 129.120 ;
        RECT 76.900 128.920 77.190 128.965 ;
        RECT 80.795 128.920 81.115 128.980 ;
        RECT 75.365 128.780 81.115 128.920 ;
        RECT 82.725 128.920 82.865 129.120 ;
        RECT 83.085 129.120 85.235 129.260 ;
        RECT 83.085 129.075 83.375 129.120 ;
        RECT 84.945 129.075 85.235 129.120 ;
        RECT 90.405 129.260 90.775 129.305 ;
        RECT 93.665 129.260 93.955 129.305 ;
        RECT 90.405 129.120 93.955 129.260 ;
        RECT 90.405 129.075 90.775 129.120 ;
        RECT 93.665 129.075 93.955 129.120 ;
        RECT 94.585 129.260 94.875 129.305 ;
        RECT 96.445 129.260 96.735 129.305 ;
        RECT 94.585 129.120 96.735 129.260 ;
        RECT 94.585 129.075 94.875 129.120 ;
        RECT 96.445 129.075 96.735 129.120 ;
        RECT 90.455 129.060 90.775 129.075 ;
        RECT 87.250 128.920 87.540 128.965 ;
        RECT 82.725 128.780 87.540 128.920 ;
        RECT 72.515 128.720 72.835 128.780 ;
        RECT 72.990 128.735 73.280 128.780 ;
        RECT 76.900 128.735 77.190 128.780 ;
        RECT 80.795 128.720 81.115 128.780 ;
        RECT 87.250 128.735 87.540 128.780 ;
        RECT 17.370 128.100 112.465 128.580 ;
        RECT 32.035 127.900 32.355 127.960 ;
        RECT 33.890 127.900 34.180 127.945 ;
        RECT 32.035 127.760 34.180 127.900 ;
        RECT 32.035 127.700 32.355 127.760 ;
        RECT 33.890 127.715 34.180 127.760 ;
        RECT 35.730 127.900 36.020 127.945 ;
        RECT 36.635 127.900 36.955 127.960 ;
        RECT 35.730 127.760 36.955 127.900 ;
        RECT 35.730 127.715 36.020 127.760 ;
        RECT 36.635 127.700 36.955 127.760 ;
        RECT 50.435 127.900 50.755 127.960 ;
        RECT 55.740 127.900 56.030 127.945 ;
        RECT 58.715 127.900 59.035 127.960 ;
        RECT 87.235 127.900 87.555 127.960 ;
        RECT 88.170 127.900 88.460 127.945 ;
        RECT 50.435 127.760 59.035 127.900 ;
        RECT 50.435 127.700 50.755 127.760 ;
        RECT 55.740 127.715 56.030 127.760 ;
        RECT 58.715 127.700 59.035 127.760 ;
        RECT 67.545 127.760 76.885 127.900 ;
        RECT 21.010 127.560 21.300 127.605 ;
        RECT 24.625 127.560 24.915 127.605 ;
        RECT 27.885 127.560 28.175 127.605 ;
        RECT 21.010 127.420 28.175 127.560 ;
        RECT 21.010 127.375 21.300 127.420 ;
        RECT 24.625 127.375 24.915 127.420 ;
        RECT 27.885 127.375 28.175 127.420 ;
        RECT 28.805 127.560 29.095 127.605 ;
        RECT 30.665 127.560 30.955 127.605 ;
        RECT 39.870 127.560 40.160 127.605 ;
        RECT 43.995 127.560 44.315 127.620 ;
        RECT 28.805 127.420 30.955 127.560 ;
        RECT 28.805 127.375 29.095 127.420 ;
        RECT 30.665 127.375 30.955 127.420 ;
        RECT 36.265 127.420 44.315 127.560 ;
        RECT 21.455 127.020 21.775 127.280 ;
        RECT 26.485 127.220 26.775 127.265 ;
        RECT 28.805 127.220 29.020 127.375 ;
        RECT 26.485 127.080 29.020 127.220 ;
        RECT 26.485 127.035 26.775 127.080 ;
        RECT 31.115 127.020 31.435 127.280 ;
        RECT 31.590 127.220 31.880 127.265 ;
        RECT 34.335 127.220 34.655 127.280 ;
        RECT 31.590 127.080 34.655 127.220 ;
        RECT 31.590 127.035 31.880 127.080 ;
        RECT 34.335 127.020 34.655 127.080 ;
        RECT 20.535 126.880 20.855 126.940 ;
        RECT 29.750 126.880 30.040 126.925 ;
        RECT 20.535 126.740 30.040 126.880 ;
        RECT 31.205 126.880 31.345 127.020 ;
        RECT 32.510 126.880 32.800 126.925 ;
        RECT 31.205 126.740 32.800 126.880 ;
        RECT 20.535 126.680 20.855 126.740 ;
        RECT 29.750 126.695 30.040 126.740 ;
        RECT 32.510 126.695 32.800 126.740 ;
        RECT 33.430 126.880 33.720 126.925 ;
        RECT 36.265 126.880 36.405 127.420 ;
        RECT 39.870 127.375 40.160 127.420 ;
        RECT 43.995 127.360 44.315 127.420 ;
        RECT 50.895 127.360 51.215 127.620 ;
        RECT 51.815 127.560 52.135 127.620 ;
        RECT 57.795 127.605 58.115 127.620 ;
        RECT 57.745 127.560 58.115 127.605 ;
        RECT 61.005 127.560 61.295 127.605 ;
        RECT 51.815 127.420 53.425 127.560 ;
        RECT 51.815 127.360 52.135 127.420 ;
        RECT 36.650 127.035 36.940 127.265 ;
        RECT 40.330 127.220 40.620 127.265 ;
        RECT 40.330 127.080 43.305 127.220 ;
        RECT 40.330 127.035 40.620 127.080 ;
        RECT 33.430 126.740 36.405 126.880 ;
        RECT 36.725 126.880 36.865 127.035 ;
        RECT 36.725 126.740 38.245 126.880 ;
        RECT 33.430 126.695 33.720 126.740 ;
        RECT 38.105 126.585 38.245 126.740 ;
        RECT 41.250 126.695 41.540 126.925 ;
        RECT 42.155 126.880 42.475 126.940 ;
        RECT 42.630 126.880 42.920 126.925 ;
        RECT 42.155 126.740 42.920 126.880 ;
        RECT 26.485 126.540 26.775 126.585 ;
        RECT 29.265 126.540 29.555 126.585 ;
        RECT 31.125 126.540 31.415 126.585 ;
        RECT 26.485 126.400 31.415 126.540 ;
        RECT 26.485 126.355 26.775 126.400 ;
        RECT 29.265 126.355 29.555 126.400 ;
        RECT 31.125 126.355 31.415 126.400 ;
        RECT 38.030 126.355 38.320 126.585 ;
        RECT 41.325 126.540 41.465 126.695 ;
        RECT 42.155 126.680 42.475 126.740 ;
        RECT 42.630 126.695 42.920 126.740 ;
        RECT 41.695 126.540 42.015 126.600 ;
        RECT 41.325 126.400 42.015 126.540 ;
        RECT 43.165 126.540 43.305 127.080 ;
        RECT 43.535 127.020 43.855 127.280 ;
        RECT 44.470 127.220 44.760 127.265 ;
        RECT 45.375 127.220 45.695 127.280 ;
        RECT 44.470 127.080 45.695 127.220 ;
        RECT 44.470 127.035 44.760 127.080 ;
        RECT 45.375 127.020 45.695 127.080 ;
        RECT 45.835 127.020 46.155 127.280 ;
        RECT 46.295 127.020 46.615 127.280 ;
        RECT 53.285 127.265 53.425 127.420 ;
        RECT 57.745 127.420 61.295 127.560 ;
        RECT 57.745 127.375 58.115 127.420 ;
        RECT 61.005 127.375 61.295 127.420 ;
        RECT 61.925 127.560 62.215 127.605 ;
        RECT 63.785 127.560 64.075 127.605 ;
        RECT 61.925 127.420 64.075 127.560 ;
        RECT 61.925 127.375 62.215 127.420 ;
        RECT 63.785 127.375 64.075 127.420 ;
        RECT 57.795 127.360 58.115 127.375 ;
        RECT 47.230 127.220 47.520 127.265 ;
        RECT 47.230 127.080 52.045 127.220 ;
        RECT 47.230 127.035 47.520 127.080 ;
        RECT 43.625 126.880 43.765 127.020 ;
        RECT 47.675 126.880 47.995 126.940 ;
        RECT 43.625 126.740 47.995 126.880 ;
        RECT 47.675 126.680 47.995 126.740 ;
        RECT 49.515 126.680 49.835 126.940 ;
        RECT 51.905 126.925 52.045 127.080 ;
        RECT 53.210 127.035 53.500 127.265 ;
        RECT 53.655 127.020 53.975 127.280 ;
        RECT 54.130 127.035 54.420 127.265 ;
        RECT 51.830 126.695 52.120 126.925 ;
        RECT 54.205 126.880 54.345 127.035 ;
        RECT 55.035 127.020 55.355 127.280 ;
        RECT 59.605 127.220 59.895 127.265 ;
        RECT 61.925 127.220 62.140 127.375 ;
        RECT 59.605 127.080 62.140 127.220 ;
        RECT 62.395 127.220 62.715 127.280 ;
        RECT 62.870 127.220 63.160 127.265 ;
        RECT 62.395 127.080 63.160 127.220 ;
        RECT 59.605 127.035 59.895 127.080 ;
        RECT 62.395 127.020 62.715 127.080 ;
        RECT 62.870 127.035 63.160 127.080 ;
        RECT 65.155 127.220 65.475 127.280 ;
        RECT 65.630 127.220 65.920 127.265 ;
        RECT 67.545 127.220 67.685 127.760 ;
        RECT 68.375 127.360 68.695 127.620 ;
        RECT 69.310 127.560 69.600 127.605 ;
        RECT 72.515 127.560 72.835 127.620 ;
        RECT 76.195 127.560 76.515 127.620 ;
        RECT 69.310 127.420 72.835 127.560 ;
        RECT 69.310 127.375 69.600 127.420 ;
        RECT 72.515 127.360 72.835 127.420 ;
        RECT 73.525 127.420 76.515 127.560 ;
        RECT 65.155 127.080 65.920 127.220 ;
        RECT 65.155 127.020 65.475 127.080 ;
        RECT 65.630 127.035 65.920 127.080 ;
        RECT 66.165 127.080 67.685 127.220 ;
        RECT 57.335 126.880 57.655 126.940 ;
        RECT 54.205 126.740 57.655 126.880 ;
        RECT 57.335 126.680 57.655 126.740 ;
        RECT 60.095 126.880 60.415 126.940 ;
        RECT 64.710 126.880 65.000 126.925 ;
        RECT 60.095 126.740 65.000 126.880 ;
        RECT 60.095 126.680 60.415 126.740 ;
        RECT 64.710 126.695 65.000 126.740 ;
        RECT 45.835 126.540 46.155 126.600 ;
        RECT 43.165 126.400 46.155 126.540 ;
        RECT 41.695 126.340 42.015 126.400 ;
        RECT 45.835 126.340 46.155 126.400 ;
        RECT 46.295 126.540 46.615 126.600 ;
        RECT 59.605 126.540 59.895 126.585 ;
        RECT 62.385 126.540 62.675 126.585 ;
        RECT 64.245 126.540 64.535 126.585 ;
        RECT 46.295 126.400 53.195 126.540 ;
        RECT 46.295 126.340 46.615 126.400 ;
        RECT 22.835 126.245 23.155 126.260 ;
        RECT 22.620 126.015 23.155 126.245 ;
        RECT 37.570 126.200 37.860 126.245 ;
        RECT 39.395 126.200 39.715 126.260 ;
        RECT 37.570 126.060 39.715 126.200 ;
        RECT 37.570 126.015 37.860 126.060 ;
        RECT 22.835 126.000 23.155 126.015 ;
        RECT 39.395 126.000 39.715 126.060 ;
        RECT 44.930 126.200 45.220 126.245 ;
        RECT 45.375 126.200 45.695 126.260 ;
        RECT 44.930 126.060 45.695 126.200 ;
        RECT 44.930 126.015 45.220 126.060 ;
        RECT 45.375 126.000 45.695 126.060 ;
        RECT 46.755 126.000 47.075 126.260 ;
        RECT 53.055 126.200 53.195 126.400 ;
        RECT 59.605 126.400 64.535 126.540 ;
        RECT 59.605 126.355 59.895 126.400 ;
        RECT 62.385 126.355 62.675 126.400 ;
        RECT 64.245 126.355 64.535 126.400 ;
        RECT 66.165 126.245 66.305 127.080 ;
        RECT 67.930 127.035 68.220 127.265 ;
        RECT 67.455 126.880 67.775 126.940 ;
        RECT 68.005 126.880 68.145 127.035 ;
        RECT 67.455 126.740 68.145 126.880 ;
        RECT 68.465 126.880 68.605 127.360 ;
        RECT 71.135 127.020 71.455 127.280 ;
        RECT 71.610 127.035 71.900 127.265 ;
        RECT 68.850 126.880 69.140 126.925 ;
        RECT 68.465 126.740 69.140 126.880 ;
        RECT 71.685 126.880 71.825 127.035 ;
        RECT 72.055 127.020 72.375 127.280 ;
        RECT 72.990 127.220 73.280 127.265 ;
        RECT 73.525 127.220 73.665 127.420 ;
        RECT 76.195 127.360 76.515 127.420 ;
        RECT 72.990 127.080 73.665 127.220 ;
        RECT 72.990 127.035 73.280 127.080 ;
        RECT 74.815 127.020 75.135 127.280 ;
        RECT 75.275 127.220 75.595 127.280 ;
        RECT 75.750 127.220 76.040 127.265 ;
        RECT 75.275 127.080 76.040 127.220 ;
        RECT 76.745 127.220 76.885 127.760 ;
        RECT 87.235 127.760 88.460 127.900 ;
        RECT 87.235 127.700 87.555 127.760 ;
        RECT 88.170 127.715 88.460 127.760 ;
        RECT 78.970 127.560 79.260 127.605 ;
        RECT 79.875 127.560 80.195 127.620 ;
        RECT 78.970 127.420 80.195 127.560 ;
        RECT 78.970 127.375 79.260 127.420 ;
        RECT 79.875 127.360 80.195 127.420 ;
        RECT 96.065 127.420 97.125 127.560 ;
        RECT 80.335 127.220 80.655 127.280 ;
        RECT 81.730 127.220 82.020 127.265 ;
        RECT 76.745 127.080 79.185 127.220 ;
        RECT 75.275 127.020 75.595 127.080 ;
        RECT 75.750 127.035 76.040 127.080 ;
        RECT 74.905 126.880 75.045 127.020 ;
        RECT 71.685 126.740 75.045 126.880 ;
        RECT 67.455 126.680 67.775 126.740 ;
        RECT 68.850 126.695 69.140 126.740 ;
        RECT 76.655 126.680 76.975 126.940 ;
        RECT 78.035 126.680 78.355 126.940 ;
        RECT 78.510 126.695 78.800 126.925 ;
        RECT 79.045 126.880 79.185 127.080 ;
        RECT 80.335 127.080 82.020 127.220 ;
        RECT 80.335 127.020 80.655 127.080 ;
        RECT 81.730 127.035 82.020 127.080 ;
        RECT 85.855 127.220 86.175 127.280 ;
        RECT 91.850 127.220 92.140 127.265 ;
        RECT 95.530 127.220 95.820 127.265 ;
        RECT 96.065 127.220 96.205 127.420 ;
        RECT 85.855 127.080 92.140 127.220 ;
        RECT 85.855 127.020 86.175 127.080 ;
        RECT 91.850 127.035 92.140 127.080 ;
        RECT 92.385 127.080 96.205 127.220 ;
        RECT 88.155 126.880 88.475 126.940 ;
        RECT 92.385 126.880 92.525 127.080 ;
        RECT 95.530 127.035 95.820 127.080 ;
        RECT 96.435 127.020 96.755 127.280 ;
        RECT 96.985 127.220 97.125 127.420 ;
        RECT 97.830 127.220 98.120 127.265 ;
        RECT 96.985 127.080 98.120 127.220 ;
        RECT 97.830 127.035 98.120 127.080 ;
        RECT 104.730 127.220 105.020 127.265 ;
        RECT 105.635 127.220 105.955 127.280 ;
        RECT 104.730 127.080 105.955 127.220 ;
        RECT 104.730 127.035 105.020 127.080 ;
        RECT 105.635 127.020 105.955 127.080 ;
        RECT 107.015 127.020 107.335 127.280 ;
        RECT 79.045 126.740 92.525 126.880 ;
        RECT 94.610 126.880 94.900 126.925 ;
        RECT 95.975 126.880 96.295 126.940 ;
        RECT 94.610 126.740 96.295 126.880 ;
        RECT 68.375 126.540 68.695 126.600 ;
        RECT 69.770 126.540 70.060 126.585 ;
        RECT 68.375 126.400 70.060 126.540 ;
        RECT 68.375 126.340 68.695 126.400 ;
        RECT 69.770 126.355 70.060 126.400 ;
        RECT 70.215 126.540 70.535 126.600 ;
        RECT 74.830 126.540 75.120 126.585 ;
        RECT 70.215 126.400 75.120 126.540 ;
        RECT 70.215 126.340 70.535 126.400 ;
        RECT 74.830 126.355 75.120 126.400 ;
        RECT 66.090 126.200 66.380 126.245 ;
        RECT 53.055 126.060 66.380 126.200 ;
        RECT 66.090 126.015 66.380 126.060 ;
        RECT 67.010 126.200 67.300 126.245 ;
        RECT 68.835 126.200 69.155 126.260 ;
        RECT 67.010 126.060 69.155 126.200 ;
        RECT 67.010 126.015 67.300 126.060 ;
        RECT 68.835 126.000 69.155 126.060 ;
        RECT 69.310 126.200 69.600 126.245 ;
        RECT 70.675 126.200 70.995 126.260 ;
        RECT 69.310 126.060 70.995 126.200 ;
        RECT 69.310 126.015 69.600 126.060 ;
        RECT 70.675 126.000 70.995 126.060 ;
        RECT 71.135 126.200 71.455 126.260 ;
        RECT 78.585 126.200 78.725 126.695 ;
        RECT 88.155 126.680 88.475 126.740 ;
        RECT 94.610 126.695 94.900 126.740 ;
        RECT 95.975 126.680 96.295 126.740 ;
        RECT 96.910 126.695 97.200 126.925 ;
        RECT 84.015 126.540 84.335 126.600 ;
        RECT 90.930 126.540 91.220 126.585 ;
        RECT 84.015 126.400 91.220 126.540 ;
        RECT 84.015 126.340 84.335 126.400 ;
        RECT 90.930 126.355 91.220 126.400 ;
        RECT 96.435 126.540 96.755 126.600 ;
        RECT 96.985 126.540 97.125 126.695 ;
        RECT 96.435 126.400 97.125 126.540 ;
        RECT 97.815 126.540 98.135 126.600 ;
        RECT 98.750 126.540 99.040 126.585 ;
        RECT 97.815 126.400 99.040 126.540 ;
        RECT 96.435 126.340 96.755 126.400 ;
        RECT 97.815 126.340 98.135 126.400 ;
        RECT 98.750 126.355 99.040 126.400 ;
        RECT 71.135 126.060 78.725 126.200 ;
        RECT 80.810 126.200 81.100 126.245 ;
        RECT 81.715 126.200 82.035 126.260 ;
        RECT 80.810 126.060 82.035 126.200 ;
        RECT 71.135 126.000 71.455 126.060 ;
        RECT 80.810 126.015 81.100 126.060 ;
        RECT 81.715 126.000 82.035 126.060 ;
        RECT 105.175 126.000 105.495 126.260 ;
        RECT 107.935 126.000 108.255 126.260 ;
        RECT 18.165 125.380 112.465 125.860 ;
        RECT 20.535 124.980 20.855 125.240 ;
        RECT 25.380 125.180 25.670 125.225 ;
        RECT 31.575 125.180 31.895 125.240 ;
        RECT 24.305 125.040 31.895 125.180 ;
        RECT 24.305 124.840 24.445 125.040 ;
        RECT 25.380 124.995 25.670 125.040 ;
        RECT 31.575 124.980 31.895 125.040 ;
        RECT 44.455 124.980 44.775 125.240 ;
        RECT 46.755 124.980 47.075 125.240 ;
        RECT 50.895 125.180 51.215 125.240 ;
        RECT 61.490 125.180 61.780 125.225 ;
        RECT 50.895 125.040 61.780 125.180 ;
        RECT 50.895 124.980 51.215 125.040 ;
        RECT 61.490 124.995 61.780 125.040 ;
        RECT 63.315 125.180 63.635 125.240 ;
        RECT 65.630 125.180 65.920 125.225 ;
        RECT 63.315 125.040 65.920 125.180 ;
        RECT 23.385 124.700 24.445 124.840 ;
        RECT 29.245 124.840 29.535 124.885 ;
        RECT 32.025 124.840 32.315 124.885 ;
        RECT 33.885 124.840 34.175 124.885 ;
        RECT 29.245 124.700 34.175 124.840 ;
        RECT 23.385 124.545 23.525 124.700 ;
        RECT 29.245 124.655 29.535 124.700 ;
        RECT 32.025 124.655 32.315 124.700 ;
        RECT 33.885 124.655 34.175 124.700 ;
        RECT 41.695 124.840 42.015 124.900 ;
        RECT 61.565 124.840 61.705 124.995 ;
        RECT 63.315 124.980 63.635 125.040 ;
        RECT 65.630 124.995 65.920 125.040 ;
        RECT 66.075 124.980 66.395 125.240 ;
        RECT 68.390 125.180 68.680 125.225 ;
        RECT 70.215 125.180 70.535 125.240 ;
        RECT 68.390 125.040 70.535 125.180 ;
        RECT 68.390 124.995 68.680 125.040 ;
        RECT 70.215 124.980 70.535 125.040 ;
        RECT 73.895 124.980 74.215 125.240 ;
        RECT 80.425 125.040 81.945 125.180 ;
        RECT 69.755 124.840 70.075 124.900 ;
        RECT 80.425 124.840 80.565 125.040 ;
        RECT 41.695 124.700 49.745 124.840 ;
        RECT 61.565 124.700 69.525 124.840 ;
        RECT 41.695 124.640 42.015 124.700 ;
        RECT 49.605 124.560 49.745 124.700 ;
        RECT 23.310 124.315 23.600 124.545 ;
        RECT 24.230 124.500 24.520 124.545 ;
        RECT 26.055 124.500 26.375 124.560 ;
        RECT 31.115 124.500 31.435 124.560 ;
        RECT 24.230 124.360 31.435 124.500 ;
        RECT 24.230 124.315 24.520 124.360 ;
        RECT 26.055 124.300 26.375 124.360 ;
        RECT 31.115 124.300 31.435 124.360 ;
        RECT 32.495 124.300 32.815 124.560 ;
        RECT 33.415 124.500 33.735 124.560 ;
        RECT 42.155 124.500 42.475 124.560 ;
        RECT 46.295 124.500 46.615 124.560 ;
        RECT 33.415 124.360 42.475 124.500 ;
        RECT 33.415 124.300 33.735 124.360 ;
        RECT 42.155 124.300 42.475 124.360 ;
        RECT 45.465 124.360 46.615 124.500 ;
        RECT 19.630 124.160 19.920 124.205 ;
        RECT 19.630 124.020 21.225 124.160 ;
        RECT 19.630 123.975 19.920 124.020 ;
        RECT 21.085 123.525 21.225 124.020 ;
        RECT 22.835 123.960 23.155 124.220 ;
        RECT 29.245 124.160 29.535 124.205 ;
        RECT 34.335 124.160 34.655 124.220 ;
        RECT 44.455 124.160 44.775 124.220 ;
        RECT 45.465 124.205 45.605 124.360 ;
        RECT 46.295 124.300 46.615 124.360 ;
        RECT 49.515 124.500 49.835 124.560 ;
        RECT 51.830 124.500 52.120 124.545 ;
        RECT 49.515 124.360 52.120 124.500 ;
        RECT 49.515 124.300 49.835 124.360 ;
        RECT 51.830 124.315 52.120 124.360 ;
        RECT 58.715 124.300 59.035 124.560 ;
        RECT 59.175 124.300 59.495 124.560 ;
        RECT 63.790 124.500 64.080 124.545 ;
        RECT 67.455 124.500 67.775 124.560 ;
        RECT 63.790 124.360 67.775 124.500 ;
        RECT 63.790 124.315 64.080 124.360 ;
        RECT 67.455 124.300 67.775 124.360 ;
        RECT 67.915 124.300 68.235 124.560 ;
        RECT 45.390 124.160 45.680 124.205 ;
        RECT 29.245 124.020 31.780 124.160 ;
        RECT 29.245 123.975 29.535 124.020 ;
        RECT 27.385 123.820 27.675 123.865 ;
        RECT 28.815 123.820 29.135 123.880 ;
        RECT 31.565 123.865 31.780 124.020 ;
        RECT 34.335 124.020 36.865 124.160 ;
        RECT 34.335 123.960 34.655 124.020 ;
        RECT 30.645 123.820 30.935 123.865 ;
        RECT 27.385 123.680 30.935 123.820 ;
        RECT 27.385 123.635 27.675 123.680 ;
        RECT 28.815 123.620 29.135 123.680 ;
        RECT 30.645 123.635 30.935 123.680 ;
        RECT 31.565 123.820 31.855 123.865 ;
        RECT 33.425 123.820 33.715 123.865 ;
        RECT 31.565 123.680 33.715 123.820 ;
        RECT 31.565 123.635 31.855 123.680 ;
        RECT 33.425 123.635 33.715 123.680 ;
        RECT 36.725 123.525 36.865 124.020 ;
        RECT 44.455 124.020 45.680 124.160 ;
        RECT 44.455 123.960 44.775 124.020 ;
        RECT 45.390 123.975 45.680 124.020 ;
        RECT 45.835 123.960 46.155 124.220 ;
        RECT 47.675 123.960 47.995 124.220 ;
        RECT 48.610 123.975 48.900 124.205 ;
        RECT 55.970 123.975 56.260 124.205 ;
        RECT 44.010 123.820 44.300 123.865 ;
        RECT 46.295 123.820 46.615 123.880 ;
        RECT 44.010 123.680 46.615 123.820 ;
        RECT 44.010 123.635 44.300 123.680 ;
        RECT 46.295 123.620 46.615 123.680 ;
        RECT 48.685 123.820 48.825 123.975 ;
        RECT 51.370 123.820 51.660 123.865 ;
        RECT 48.685 123.680 51.660 123.820 ;
        RECT 56.045 123.820 56.185 123.975 ;
        RECT 58.255 123.960 58.575 124.220 ;
        RECT 62.410 123.975 62.700 124.205 ;
        RECT 60.095 123.820 60.415 123.880 ;
        RECT 56.045 123.680 60.415 123.820 ;
        RECT 62.485 123.820 62.625 123.975 ;
        RECT 62.855 123.960 63.175 124.220 ;
        RECT 64.695 123.960 65.015 124.220 ;
        RECT 65.705 123.900 66.765 124.040 ;
        RECT 66.995 123.960 67.315 124.220 ;
        RECT 68.375 123.960 68.695 124.220 ;
        RECT 69.385 124.205 69.525 124.700 ;
        RECT 69.755 124.700 80.565 124.840 ;
        RECT 69.755 124.640 70.075 124.700 ;
        RECT 80.810 124.655 81.100 124.885 ;
        RECT 80.885 124.500 81.025 124.655 ;
        RECT 69.845 124.360 81.025 124.500 ;
        RECT 69.310 123.975 69.600 124.205 ;
        RECT 65.155 123.820 65.475 123.880 ;
        RECT 65.705 123.820 65.845 123.900 ;
        RECT 62.485 123.680 65.845 123.820 ;
        RECT 66.625 123.820 66.765 123.900 ;
        RECT 69.845 123.820 69.985 124.360 ;
        RECT 80.335 123.960 80.655 124.220 ;
        RECT 81.805 124.205 81.945 125.040 ;
        RECT 85.855 124.980 86.175 125.240 ;
        RECT 89.550 125.180 89.840 125.225 ;
        RECT 90.915 125.180 91.235 125.240 ;
        RECT 89.550 125.040 91.235 125.180 ;
        RECT 89.550 124.995 89.840 125.040 ;
        RECT 90.915 124.980 91.235 125.040 ;
        RECT 92.755 125.180 93.075 125.240 ;
        RECT 94.150 125.180 94.440 125.225 ;
        RECT 107.015 125.180 107.335 125.240 ;
        RECT 92.755 125.040 94.440 125.180 ;
        RECT 92.755 124.980 93.075 125.040 ;
        RECT 94.150 124.995 94.440 125.040 ;
        RECT 105.265 125.040 107.335 125.180 ;
        RECT 83.555 124.840 83.875 124.900 ;
        RECT 89.090 124.840 89.380 124.885 ;
        RECT 89.995 124.840 90.315 124.900 ;
        RECT 83.555 124.700 88.845 124.840 ;
        RECT 83.555 124.640 83.875 124.700 ;
        RECT 82.635 124.300 82.955 124.560 ;
        RECT 88.705 124.500 88.845 124.700 ;
        RECT 89.090 124.700 90.315 124.840 ;
        RECT 89.090 124.655 89.380 124.700 ;
        RECT 89.995 124.640 90.315 124.700 ;
        RECT 93.215 124.840 93.535 124.900 ;
        RECT 94.610 124.840 94.900 124.885 ;
        RECT 93.215 124.700 94.900 124.840 ;
        RECT 93.215 124.640 93.535 124.700 ;
        RECT 94.610 124.655 94.900 124.700 ;
        RECT 95.055 124.840 95.375 124.900 ;
        RECT 101.050 124.840 101.340 124.885 ;
        RECT 105.265 124.840 105.405 125.040 ;
        RECT 107.015 124.980 107.335 125.040 ;
        RECT 95.055 124.700 98.505 124.840 ;
        RECT 95.055 124.640 95.375 124.700 ;
        RECT 91.390 124.500 91.680 124.545 ;
        RECT 96.450 124.500 96.740 124.545 ;
        RECT 97.815 124.500 98.135 124.560 ;
        RECT 98.365 124.545 98.505 124.700 ;
        RECT 101.050 124.700 105.405 124.840 ;
        RECT 105.605 124.840 105.895 124.885 ;
        RECT 108.385 124.840 108.675 124.885 ;
        RECT 110.245 124.840 110.535 124.885 ;
        RECT 105.605 124.700 110.535 124.840 ;
        RECT 101.050 124.655 101.340 124.700 ;
        RECT 105.605 124.655 105.895 124.700 ;
        RECT 108.385 124.655 108.675 124.700 ;
        RECT 110.245 124.655 110.535 124.700 ;
        RECT 88.705 124.360 91.680 124.500 ;
        RECT 91.390 124.315 91.680 124.360 ;
        RECT 92.385 124.360 93.445 124.500 ;
        RECT 81.730 123.975 82.020 124.205 ;
        RECT 87.710 123.975 88.000 124.205 ;
        RECT 88.155 124.160 88.475 124.220 ;
        RECT 90.470 124.160 90.760 124.205 ;
        RECT 92.385 124.160 92.525 124.360 ;
        RECT 93.305 124.205 93.445 124.360 ;
        RECT 96.450 124.360 98.135 124.500 ;
        RECT 96.450 124.315 96.740 124.360 ;
        RECT 97.815 124.300 98.135 124.360 ;
        RECT 98.290 124.315 98.580 124.545 ;
        RECT 107.935 124.500 108.255 124.560 ;
        RECT 108.870 124.500 109.160 124.545 ;
        RECT 107.935 124.360 109.160 124.500 ;
        RECT 107.935 124.300 108.255 124.360 ;
        RECT 108.870 124.315 109.160 124.360 ;
        RECT 88.155 124.020 92.525 124.160 ;
        RECT 78.035 123.820 78.355 123.880 ;
        RECT 66.625 123.680 69.985 123.820 ;
        RECT 70.305 123.680 78.355 123.820 ;
        RECT 21.010 123.295 21.300 123.525 ;
        RECT 36.650 123.480 36.940 123.525 ;
        RECT 37.095 123.480 37.415 123.540 ;
        RECT 36.650 123.340 37.415 123.480 ;
        RECT 36.650 123.295 36.940 123.340 ;
        RECT 37.095 123.280 37.415 123.340 ;
        RECT 43.535 123.480 43.855 123.540 ;
        RECT 48.685 123.480 48.825 123.680 ;
        RECT 51.370 123.635 51.660 123.680 ;
        RECT 60.095 123.620 60.415 123.680 ;
        RECT 65.155 123.620 65.475 123.680 ;
        RECT 70.305 123.540 70.445 123.680 ;
        RECT 78.035 123.620 78.355 123.680 ;
        RECT 80.795 123.820 81.115 123.880 ;
        RECT 83.570 123.820 83.860 123.865 ;
        RECT 80.795 123.680 83.860 123.820 ;
        RECT 87.785 123.820 87.925 123.975 ;
        RECT 88.155 123.960 88.475 124.020 ;
        RECT 90.470 123.975 90.760 124.020 ;
        RECT 92.770 123.975 93.060 124.205 ;
        RECT 93.230 124.160 93.520 124.205 ;
        RECT 95.530 124.160 95.820 124.205 ;
        RECT 93.230 124.020 95.820 124.160 ;
        RECT 93.230 123.975 93.520 124.020 ;
        RECT 95.530 123.975 95.820 124.020 ;
        RECT 95.975 124.160 96.295 124.220 ;
        RECT 98.750 124.160 99.040 124.205 ;
        RECT 95.975 124.020 99.040 124.160 ;
        RECT 89.995 123.820 90.315 123.880 ;
        RECT 87.785 123.680 90.315 123.820 ;
        RECT 92.845 123.820 92.985 123.975 ;
        RECT 95.975 123.960 96.295 124.020 ;
        RECT 98.750 123.975 99.040 124.020 ;
        RECT 105.605 124.160 105.895 124.205 ;
        RECT 109.315 124.160 109.635 124.220 ;
        RECT 110.710 124.160 111.000 124.205 ;
        RECT 105.605 124.020 108.140 124.160 ;
        RECT 105.605 123.975 105.895 124.020 ;
        RECT 96.895 123.820 97.215 123.880 ;
        RECT 92.845 123.680 97.215 123.820 ;
        RECT 80.795 123.620 81.115 123.680 ;
        RECT 83.570 123.635 83.860 123.680 ;
        RECT 89.995 123.620 90.315 123.680 ;
        RECT 96.895 123.620 97.215 123.680 ;
        RECT 103.745 123.820 104.035 123.865 ;
        RECT 105.175 123.820 105.495 123.880 ;
        RECT 107.925 123.865 108.140 124.020 ;
        RECT 109.315 124.020 111.000 124.160 ;
        RECT 109.315 123.960 109.635 124.020 ;
        RECT 110.710 123.975 111.000 124.020 ;
        RECT 107.005 123.820 107.295 123.865 ;
        RECT 103.745 123.680 107.295 123.820 ;
        RECT 103.745 123.635 104.035 123.680 ;
        RECT 105.175 123.620 105.495 123.680 ;
        RECT 107.005 123.635 107.295 123.680 ;
        RECT 107.925 123.820 108.215 123.865 ;
        RECT 109.785 123.820 110.075 123.865 ;
        RECT 107.925 123.680 110.075 123.820 ;
        RECT 107.925 123.635 108.215 123.680 ;
        RECT 109.785 123.635 110.075 123.680 ;
        RECT 43.535 123.340 48.825 123.480 ;
        RECT 43.535 123.280 43.855 123.340 ;
        RECT 49.055 123.280 49.375 123.540 ;
        RECT 50.895 123.280 51.215 123.540 ;
        RECT 54.575 123.480 54.895 123.540 ;
        RECT 56.430 123.480 56.720 123.525 ;
        RECT 54.575 123.340 56.720 123.480 ;
        RECT 54.575 123.280 54.895 123.340 ;
        RECT 56.430 123.295 56.720 123.340 ;
        RECT 64.695 123.480 65.015 123.540 ;
        RECT 69.295 123.480 69.615 123.540 ;
        RECT 64.695 123.340 69.615 123.480 ;
        RECT 64.695 123.280 65.015 123.340 ;
        RECT 69.295 123.280 69.615 123.340 ;
        RECT 69.770 123.480 70.060 123.525 ;
        RECT 70.215 123.480 70.535 123.540 ;
        RECT 69.770 123.340 70.535 123.480 ;
        RECT 69.770 123.295 70.060 123.340 ;
        RECT 70.215 123.280 70.535 123.340 ;
        RECT 72.055 123.480 72.375 123.540 ;
        RECT 84.030 123.480 84.320 123.525 ;
        RECT 86.775 123.480 87.095 123.540 ;
        RECT 72.055 123.340 87.095 123.480 ;
        RECT 72.055 123.280 72.375 123.340 ;
        RECT 84.030 123.295 84.320 123.340 ;
        RECT 86.775 123.280 87.095 123.340 ;
        RECT 96.435 123.480 96.755 123.540 ;
        RECT 99.210 123.480 99.500 123.525 ;
        RECT 101.740 123.480 102.030 123.525 ;
        RECT 96.435 123.340 102.030 123.480 ;
        RECT 96.435 123.280 96.755 123.340 ;
        RECT 99.210 123.295 99.500 123.340 ;
        RECT 101.740 123.295 102.030 123.340 ;
        RECT 17.370 122.660 112.465 123.140 ;
        RECT 32.280 122.460 32.570 122.505 ;
        RECT 43.075 122.460 43.395 122.520 ;
        RECT 43.550 122.460 43.840 122.505 ;
        RECT 32.280 122.320 41.005 122.460 ;
        RECT 32.280 122.275 32.570 122.320 ;
        RECT 21.915 122.120 22.235 122.180 ;
        RECT 24.625 122.120 24.915 122.165 ;
        RECT 27.885 122.120 28.175 122.165 ;
        RECT 21.915 121.980 28.175 122.120 ;
        RECT 21.915 121.920 22.235 121.980 ;
        RECT 24.625 121.935 24.915 121.980 ;
        RECT 27.885 121.935 28.175 121.980 ;
        RECT 28.805 122.120 29.095 122.165 ;
        RECT 30.665 122.120 30.955 122.165 ;
        RECT 28.805 121.980 30.955 122.120 ;
        RECT 28.805 121.935 29.095 121.980 ;
        RECT 30.665 121.935 30.955 121.980 ;
        RECT 32.955 122.120 33.275 122.180 ;
        RECT 34.285 122.120 34.575 122.165 ;
        RECT 37.545 122.120 37.835 122.165 ;
        RECT 32.955 121.980 37.835 122.120 ;
        RECT 20.550 121.780 20.840 121.825 ;
        RECT 22.835 121.780 23.155 121.840 ;
        RECT 20.550 121.640 23.155 121.780 ;
        RECT 20.550 121.595 20.840 121.640 ;
        RECT 22.835 121.580 23.155 121.640 ;
        RECT 26.485 121.780 26.775 121.825 ;
        RECT 28.805 121.780 29.020 121.935 ;
        RECT 32.955 121.920 33.275 121.980 ;
        RECT 34.285 121.935 34.575 121.980 ;
        RECT 37.545 121.935 37.835 121.980 ;
        RECT 38.465 122.120 38.755 122.165 ;
        RECT 40.325 122.120 40.615 122.165 ;
        RECT 38.465 121.980 40.615 122.120 ;
        RECT 40.865 122.120 41.005 122.320 ;
        RECT 43.075 122.320 43.840 122.460 ;
        RECT 43.075 122.260 43.395 122.320 ;
        RECT 43.550 122.275 43.840 122.320 ;
        RECT 46.295 122.460 46.615 122.520 ;
        RECT 55.955 122.460 56.275 122.520 ;
        RECT 46.295 122.320 56.275 122.460 ;
        RECT 46.295 122.260 46.615 122.320 ;
        RECT 43.995 122.120 44.315 122.180 ;
        RECT 48.225 122.165 48.365 122.320 ;
        RECT 55.955 122.260 56.275 122.320 ;
        RECT 57.335 122.460 57.655 122.520 ;
        RECT 58.040 122.460 58.330 122.505 ;
        RECT 62.395 122.460 62.715 122.520 ;
        RECT 66.995 122.460 67.315 122.520 ;
        RECT 57.335 122.320 58.330 122.460 ;
        RECT 57.335 122.260 57.655 122.320 ;
        RECT 58.040 122.275 58.330 122.320 ;
        RECT 59.265 122.320 62.715 122.460 ;
        RECT 40.865 121.980 45.145 122.120 ;
        RECT 38.465 121.935 38.755 121.980 ;
        RECT 40.325 121.935 40.615 121.980 ;
        RECT 26.485 121.640 29.020 121.780 ;
        RECT 36.145 121.780 36.435 121.825 ;
        RECT 38.465 121.780 38.680 121.935 ;
        RECT 43.995 121.920 44.315 121.980 ;
        RECT 36.145 121.640 38.680 121.780 ;
        RECT 26.485 121.595 26.775 121.640 ;
        RECT 36.145 121.595 36.435 121.640 ;
        RECT 39.395 121.580 39.715 121.840 ;
        RECT 42.630 121.595 42.920 121.825 ;
        RECT 29.750 121.440 30.040 121.485 ;
        RECT 21.545 121.300 30.040 121.440 ;
        RECT 21.545 121.145 21.685 121.300 ;
        RECT 29.750 121.255 30.040 121.300 ;
        RECT 31.590 121.440 31.880 121.485 ;
        RECT 37.095 121.440 37.415 121.500 ;
        RECT 41.250 121.440 41.540 121.485 ;
        RECT 42.705 121.440 42.845 121.595 ;
        RECT 44.455 121.580 44.775 121.840 ;
        RECT 45.005 121.825 45.145 121.980 ;
        RECT 48.150 121.935 48.440 122.165 ;
        RECT 55.035 122.120 55.355 122.180 ;
        RECT 59.265 122.120 59.405 122.320 ;
        RECT 62.395 122.260 62.715 122.320 ;
        RECT 63.865 122.320 67.315 122.460 ;
        RECT 55.035 121.980 59.405 122.120 ;
        RECT 60.045 122.120 60.335 122.165 ;
        RECT 63.305 122.120 63.595 122.165 ;
        RECT 63.865 122.120 64.005 122.320 ;
        RECT 66.995 122.260 67.315 122.320 ;
        RECT 68.390 122.460 68.680 122.505 ;
        RECT 69.295 122.460 69.615 122.520 ;
        RECT 68.390 122.320 69.615 122.460 ;
        RECT 68.390 122.275 68.680 122.320 ;
        RECT 69.295 122.260 69.615 122.320 ;
        RECT 71.135 122.260 71.455 122.520 ;
        RECT 92.845 122.320 93.905 122.460 ;
        RECT 60.045 121.980 64.005 122.120 ;
        RECT 64.225 122.120 64.515 122.165 ;
        RECT 66.085 122.120 66.375 122.165 ;
        RECT 64.225 121.980 66.375 122.120 ;
        RECT 55.035 121.920 55.355 121.980 ;
        RECT 60.045 121.935 60.335 121.980 ;
        RECT 63.305 121.935 63.595 121.980 ;
        RECT 64.225 121.935 64.515 121.980 ;
        RECT 66.085 121.935 66.375 121.980 ;
        RECT 68.835 122.120 69.155 122.180 ;
        RECT 74.815 122.120 75.135 122.180 ;
        RECT 68.835 121.980 75.135 122.120 ;
        RECT 44.930 121.595 45.220 121.825 ;
        RECT 46.310 121.780 46.600 121.825 ;
        RECT 49.055 121.780 49.375 121.840 ;
        RECT 46.310 121.640 49.375 121.780 ;
        RECT 46.310 121.595 46.600 121.640 ;
        RECT 49.055 121.580 49.375 121.640 ;
        RECT 61.905 121.780 62.195 121.825 ;
        RECT 64.225 121.780 64.440 121.935 ;
        RECT 68.835 121.920 69.155 121.980 ;
        RECT 74.815 121.920 75.135 121.980 ;
        RECT 78.055 122.120 78.345 122.165 ;
        RECT 79.915 122.120 80.205 122.165 ;
        RECT 78.055 121.980 80.205 122.120 ;
        RECT 78.055 121.935 78.345 121.980 ;
        RECT 79.915 121.935 80.205 121.980 ;
        RECT 80.835 122.120 81.125 122.165 ;
        RECT 82.635 122.120 82.955 122.180 ;
        RECT 84.095 122.120 84.385 122.165 ;
        RECT 80.835 121.980 84.385 122.120 ;
        RECT 80.835 121.935 81.125 121.980 ;
        RECT 61.905 121.640 64.440 121.780 ;
        RECT 65.170 121.780 65.460 121.825 ;
        RECT 67.455 121.780 67.775 121.840 ;
        RECT 65.170 121.640 67.775 121.780 ;
        RECT 61.905 121.595 62.195 121.640 ;
        RECT 65.170 121.595 65.460 121.640 ;
        RECT 67.455 121.580 67.775 121.640 ;
        RECT 67.930 121.780 68.220 121.825 ;
        RECT 69.755 121.780 70.075 121.840 ;
        RECT 67.930 121.640 70.075 121.780 ;
        RECT 67.930 121.595 68.220 121.640 ;
        RECT 69.755 121.580 70.075 121.640 ;
        RECT 73.895 121.780 74.215 121.840 ;
        RECT 74.370 121.780 74.660 121.825 ;
        RECT 77.130 121.780 77.420 121.825 ;
        RECT 73.895 121.640 77.420 121.780 ;
        RECT 79.990 121.780 80.205 121.935 ;
        RECT 82.635 121.920 82.955 121.980 ;
        RECT 84.095 121.935 84.385 121.980 ;
        RECT 82.235 121.780 82.525 121.825 ;
        RECT 89.550 121.780 89.840 121.825 ;
        RECT 79.990 121.640 82.525 121.780 ;
        RECT 73.895 121.580 74.215 121.640 ;
        RECT 74.370 121.595 74.660 121.640 ;
        RECT 77.130 121.595 77.420 121.640 ;
        RECT 82.235 121.595 82.525 121.640 ;
        RECT 86.175 121.640 89.840 121.780 ;
        RECT 31.590 121.300 42.845 121.440 ;
        RECT 56.890 121.440 57.180 121.485 ;
        RECT 60.095 121.440 60.415 121.500 ;
        RECT 67.010 121.440 67.300 121.485 ;
        RECT 56.890 121.300 67.300 121.440 ;
        RECT 31.590 121.255 31.880 121.300 ;
        RECT 37.095 121.240 37.415 121.300 ;
        RECT 41.250 121.255 41.540 121.300 ;
        RECT 56.890 121.255 57.180 121.300 ;
        RECT 60.095 121.240 60.415 121.300 ;
        RECT 67.010 121.255 67.300 121.300 ;
        RECT 70.215 121.240 70.535 121.500 ;
        RECT 70.690 121.440 70.980 121.485 ;
        RECT 73.435 121.440 73.755 121.500 ;
        RECT 75.735 121.440 76.055 121.500 ;
        RECT 70.690 121.300 76.055 121.440 ;
        RECT 77.205 121.440 77.345 121.595 ;
        RECT 78.035 121.440 78.355 121.500 ;
        RECT 77.205 121.300 78.355 121.440 ;
        RECT 70.690 121.255 70.980 121.300 ;
        RECT 73.435 121.240 73.755 121.300 ;
        RECT 75.735 121.240 76.055 121.300 ;
        RECT 78.035 121.240 78.355 121.300 ;
        RECT 78.955 121.240 79.275 121.500 ;
        RECT 79.875 121.440 80.195 121.500 ;
        RECT 86.175 121.485 86.315 121.640 ;
        RECT 89.550 121.595 89.840 121.640 ;
        RECT 89.995 121.580 90.315 121.840 ;
        RECT 92.845 121.780 92.985 122.320 ;
        RECT 93.765 122.120 93.905 122.320 ;
        RECT 96.435 122.260 96.755 122.520 ;
        RECT 96.895 122.460 97.215 122.520 ;
        RECT 99.195 122.460 99.515 122.520 ;
        RECT 101.280 122.460 101.570 122.505 ;
        RECT 96.895 122.320 101.570 122.460 ;
        RECT 96.895 122.260 97.215 122.320 ;
        RECT 99.195 122.260 99.515 122.320 ;
        RECT 101.280 122.275 101.570 122.320 ;
        RECT 106.555 122.165 106.875 122.180 ;
        RECT 103.285 122.120 103.575 122.165 ;
        RECT 106.545 122.120 106.875 122.165 ;
        RECT 93.765 121.980 100.805 122.120 ;
        RECT 93.230 121.780 93.520 121.825 ;
        RECT 92.845 121.640 93.520 121.780 ;
        RECT 93.230 121.595 93.520 121.640 ;
        RECT 93.675 121.580 93.995 121.840 ;
        RECT 100.665 121.825 100.805 121.980 ;
        RECT 103.285 121.980 106.875 122.120 ;
        RECT 103.285 121.935 103.575 121.980 ;
        RECT 106.545 121.935 106.875 121.980 ;
        RECT 106.555 121.920 106.875 121.935 ;
        RECT 107.465 122.120 107.755 122.165 ;
        RECT 109.325 122.120 109.615 122.165 ;
        RECT 107.465 121.980 109.615 122.120 ;
        RECT 107.465 121.935 107.755 121.980 ;
        RECT 109.325 121.935 109.615 121.980 ;
        RECT 100.590 121.595 100.880 121.825 ;
        RECT 105.145 121.780 105.435 121.825 ;
        RECT 107.465 121.780 107.680 121.935 ;
        RECT 105.145 121.640 107.680 121.780 ;
        RECT 108.855 121.780 109.175 121.840 ;
        RECT 110.250 121.780 110.540 121.825 ;
        RECT 110.695 121.780 111.015 121.840 ;
        RECT 108.855 121.640 111.015 121.780 ;
        RECT 105.145 121.595 105.435 121.640 ;
        RECT 86.100 121.440 86.390 121.485 ;
        RECT 79.875 121.300 86.390 121.440 ;
        RECT 79.875 121.240 80.195 121.300 ;
        RECT 86.100 121.255 86.390 121.300 ;
        RECT 87.235 121.440 87.555 121.500 ;
        RECT 88.630 121.440 88.920 121.485 ;
        RECT 95.055 121.440 95.375 121.500 ;
        RECT 95.530 121.440 95.820 121.485 ;
        RECT 96.895 121.440 97.215 121.500 ;
        RECT 87.235 121.300 97.215 121.440 ;
        RECT 100.665 121.440 100.805 121.595 ;
        RECT 108.855 121.580 109.175 121.640 ;
        RECT 110.250 121.595 110.540 121.640 ;
        RECT 110.695 121.580 111.015 121.640 ;
        RECT 105.635 121.440 105.955 121.500 ;
        RECT 100.665 121.300 105.955 121.440 ;
        RECT 87.235 121.240 87.555 121.300 ;
        RECT 88.630 121.255 88.920 121.300 ;
        RECT 95.055 121.240 95.375 121.300 ;
        RECT 95.530 121.255 95.820 121.300 ;
        RECT 96.895 121.240 97.215 121.300 ;
        RECT 105.635 121.240 105.955 121.300 ;
        RECT 108.395 121.240 108.715 121.500 ;
        RECT 21.470 120.915 21.760 121.145 ;
        RECT 26.485 121.100 26.775 121.145 ;
        RECT 29.265 121.100 29.555 121.145 ;
        RECT 31.125 121.100 31.415 121.145 ;
        RECT 26.485 120.960 31.415 121.100 ;
        RECT 26.485 120.915 26.775 120.960 ;
        RECT 29.265 120.915 29.555 120.960 ;
        RECT 31.125 120.915 31.415 120.960 ;
        RECT 36.145 121.100 36.435 121.145 ;
        RECT 38.925 121.100 39.215 121.145 ;
        RECT 40.785 121.100 41.075 121.145 ;
        RECT 36.145 120.960 41.075 121.100 ;
        RECT 36.145 120.915 36.435 120.960 ;
        RECT 38.925 120.915 39.215 120.960 ;
        RECT 40.785 120.915 41.075 120.960 ;
        RECT 61.905 121.100 62.195 121.145 ;
        RECT 64.685 121.100 64.975 121.145 ;
        RECT 66.545 121.100 66.835 121.145 ;
        RECT 61.905 120.960 66.835 121.100 ;
        RECT 61.905 120.915 62.195 120.960 ;
        RECT 64.685 120.915 64.975 120.960 ;
        RECT 66.545 120.915 66.835 120.960 ;
        RECT 77.595 121.100 77.885 121.145 ;
        RECT 79.455 121.100 79.745 121.145 ;
        RECT 82.235 121.100 82.525 121.145 ;
        RECT 77.595 120.960 82.525 121.100 ;
        RECT 77.595 120.915 77.885 120.960 ;
        RECT 79.455 120.915 79.745 120.960 ;
        RECT 82.235 120.915 82.525 120.960 ;
        RECT 91.850 121.100 92.140 121.145 ;
        RECT 93.675 121.100 93.995 121.160 ;
        RECT 91.850 120.960 93.995 121.100 ;
        RECT 91.850 120.915 92.140 120.960 ;
        RECT 93.675 120.900 93.995 120.960 ;
        RECT 94.135 121.100 94.455 121.160 ;
        RECT 100.130 121.100 100.420 121.145 ;
        RECT 94.135 120.960 100.420 121.100 ;
        RECT 94.135 120.900 94.455 120.960 ;
        RECT 100.130 120.915 100.420 120.960 ;
        RECT 105.145 121.100 105.435 121.145 ;
        RECT 107.925 121.100 108.215 121.145 ;
        RECT 109.785 121.100 110.075 121.145 ;
        RECT 105.145 120.960 110.075 121.100 ;
        RECT 105.145 120.915 105.435 120.960 ;
        RECT 107.925 120.915 108.215 120.960 ;
        RECT 109.785 120.915 110.075 120.960 ;
        RECT 22.620 120.760 22.910 120.805 ;
        RECT 24.675 120.760 24.995 120.820 ;
        RECT 22.620 120.620 24.995 120.760 ;
        RECT 22.620 120.575 22.910 120.620 ;
        RECT 24.675 120.560 24.995 120.620 ;
        RECT 34.335 120.760 34.655 120.820 ;
        RECT 46.755 120.760 47.075 120.820 ;
        RECT 34.335 120.620 47.075 120.760 ;
        RECT 34.335 120.560 34.655 120.620 ;
        RECT 46.755 120.560 47.075 120.620 ;
        RECT 47.230 120.760 47.520 120.805 ;
        RECT 55.955 120.760 56.275 120.820 ;
        RECT 47.230 120.620 56.275 120.760 ;
        RECT 47.230 120.575 47.520 120.620 ;
        RECT 55.955 120.560 56.275 120.620 ;
        RECT 59.635 120.760 59.955 120.820 ;
        RECT 63.315 120.760 63.635 120.820 ;
        RECT 59.635 120.620 63.635 120.760 ;
        RECT 59.635 120.560 59.955 120.620 ;
        RECT 63.315 120.560 63.635 120.620 ;
        RECT 72.975 120.560 73.295 120.820 ;
        RECT 92.770 120.760 93.060 120.805 ;
        RECT 93.215 120.760 93.535 120.820 ;
        RECT 92.770 120.620 93.535 120.760 ;
        RECT 92.770 120.575 93.060 120.620 ;
        RECT 93.215 120.560 93.535 120.620 ;
        RECT 94.610 120.760 94.900 120.805 ;
        RECT 95.055 120.760 95.375 120.820 ;
        RECT 94.610 120.620 95.375 120.760 ;
        RECT 94.610 120.575 94.900 120.620 ;
        RECT 95.055 120.560 95.375 120.620 ;
        RECT 98.735 120.560 99.055 120.820 ;
        RECT 18.165 119.940 112.465 120.420 ;
        RECT 21.915 119.540 22.235 119.800 ;
        RECT 22.835 119.540 23.155 119.800 ;
        RECT 33.415 119.740 33.735 119.800 ;
        RECT 28.445 119.600 33.735 119.740 ;
        RECT 24.675 119.400 24.995 119.460 ;
        RECT 28.445 119.400 28.585 119.600 ;
        RECT 33.415 119.540 33.735 119.600 ;
        RECT 34.335 119.540 34.655 119.800 ;
        RECT 37.555 119.540 37.875 119.800 ;
        RECT 40.790 119.740 41.080 119.785 ;
        RECT 48.595 119.740 48.915 119.800 ;
        RECT 40.790 119.600 48.915 119.740 ;
        RECT 40.790 119.555 41.080 119.600 ;
        RECT 48.595 119.540 48.915 119.600 ;
        RECT 54.590 119.740 54.880 119.785 ;
        RECT 55.035 119.740 55.355 119.800 ;
        RECT 54.590 119.600 55.355 119.740 ;
        RECT 54.590 119.555 54.880 119.600 ;
        RECT 55.035 119.540 55.355 119.600 ;
        RECT 55.510 119.740 55.800 119.785 ;
        RECT 57.795 119.740 58.115 119.800 ;
        RECT 55.510 119.600 58.115 119.740 ;
        RECT 55.510 119.555 55.800 119.600 ;
        RECT 57.795 119.540 58.115 119.600 ;
        RECT 59.175 119.740 59.495 119.800 ;
        RECT 65.630 119.740 65.920 119.785 ;
        RECT 66.535 119.740 66.855 119.800 ;
        RECT 59.175 119.600 63.545 119.740 ;
        RECT 59.175 119.540 59.495 119.600 ;
        RECT 39.855 119.400 40.175 119.460 ;
        RECT 41.250 119.400 41.540 119.445 ;
        RECT 53.210 119.400 53.500 119.445 ;
        RECT 59.635 119.400 59.955 119.460 ;
        RECT 24.675 119.260 28.585 119.400 ;
        RECT 24.675 119.200 24.995 119.260 ;
        RECT 23.295 119.060 23.615 119.120 ;
        RECT 25.150 119.060 25.440 119.105 ;
        RECT 23.295 118.920 25.440 119.060 ;
        RECT 23.295 118.860 23.615 118.920 ;
        RECT 25.150 118.875 25.440 118.920 ;
        RECT 26.055 119.060 26.375 119.120 ;
        RECT 28.445 119.105 28.585 119.260 ;
        RECT 28.905 119.260 35.945 119.400 ;
        RECT 27.450 119.060 27.740 119.105 ;
        RECT 26.055 118.920 27.740 119.060 ;
        RECT 26.055 118.860 26.375 118.920 ;
        RECT 27.450 118.875 27.740 118.920 ;
        RECT 28.370 118.875 28.660 119.105 ;
        RECT 21.455 118.520 21.775 118.780 ;
        RECT 24.675 118.520 24.995 118.780 ;
        RECT 25.595 118.720 25.915 118.780 ;
        RECT 28.905 118.765 29.045 119.260 ;
        RECT 31.575 119.060 31.895 119.120 ;
        RECT 35.805 119.105 35.945 119.260 ;
        RECT 39.855 119.260 41.540 119.400 ;
        RECT 39.855 119.200 40.175 119.260 ;
        RECT 41.250 119.215 41.540 119.260 ;
        RECT 43.165 119.260 49.745 119.400 ;
        RECT 43.165 119.105 43.305 119.260 ;
        RECT 32.510 119.060 32.800 119.105 ;
        RECT 31.575 118.920 32.800 119.060 ;
        RECT 31.575 118.860 31.895 118.920 ;
        RECT 32.510 118.875 32.800 118.920 ;
        RECT 35.730 118.875 36.020 119.105 ;
        RECT 43.090 118.875 43.380 119.105 ;
        RECT 44.470 119.060 44.760 119.105 ;
        RECT 46.295 119.060 46.615 119.120 ;
        RECT 48.610 119.060 48.900 119.105 ;
        RECT 49.055 119.060 49.375 119.120 ;
        RECT 49.605 119.105 49.745 119.260 ;
        RECT 53.210 119.260 59.955 119.400 ;
        RECT 53.210 119.215 53.500 119.260 ;
        RECT 59.635 119.200 59.955 119.260 ;
        RECT 60.110 119.400 60.400 119.445 ;
        RECT 60.555 119.400 60.875 119.460 ;
        RECT 60.110 119.260 60.875 119.400 ;
        RECT 60.110 119.215 60.400 119.260 ;
        RECT 60.555 119.200 60.875 119.260 ;
        RECT 61.015 119.200 61.335 119.460 ;
        RECT 63.405 119.400 63.545 119.600 ;
        RECT 65.630 119.600 66.855 119.740 ;
        RECT 65.630 119.555 65.920 119.600 ;
        RECT 66.535 119.540 66.855 119.600 ;
        RECT 66.995 119.540 67.315 119.800 ;
        RECT 67.915 119.740 68.235 119.800 ;
        RECT 69.080 119.740 69.370 119.785 ;
        RECT 71.135 119.740 71.455 119.800 ;
        RECT 67.915 119.600 71.455 119.740 ;
        RECT 67.915 119.540 68.235 119.600 ;
        RECT 69.080 119.555 69.370 119.600 ;
        RECT 71.135 119.540 71.455 119.600 ;
        RECT 78.495 119.540 78.815 119.800 ;
        RECT 78.955 119.740 79.275 119.800 ;
        RECT 80.810 119.740 81.100 119.785 ;
        RECT 78.955 119.600 81.100 119.740 ;
        RECT 78.955 119.540 79.275 119.600 ;
        RECT 80.810 119.555 81.100 119.600 ;
        RECT 87.940 119.740 88.230 119.785 ;
        RECT 89.995 119.740 90.315 119.800 ;
        RECT 87.940 119.600 90.315 119.740 ;
        RECT 87.940 119.555 88.230 119.600 ;
        RECT 89.995 119.540 90.315 119.600 ;
        RECT 95.975 119.740 96.295 119.800 ;
        RECT 100.575 119.740 100.895 119.800 ;
        RECT 106.110 119.740 106.400 119.785 ;
        RECT 106.555 119.740 106.875 119.800 ;
        RECT 95.975 119.600 103.565 119.740 ;
        RECT 95.975 119.540 96.295 119.600 ;
        RECT 100.575 119.540 100.895 119.600 ;
        RECT 72.945 119.400 73.235 119.445 ;
        RECT 75.725 119.400 76.015 119.445 ;
        RECT 77.585 119.400 77.875 119.445 ;
        RECT 63.405 119.260 64.005 119.400 ;
        RECT 44.470 118.920 49.375 119.060 ;
        RECT 44.470 118.875 44.760 118.920 ;
        RECT 46.295 118.860 46.615 118.920 ;
        RECT 48.610 118.875 48.900 118.920 ;
        RECT 49.055 118.860 49.375 118.920 ;
        RECT 49.530 119.060 49.820 119.105 ;
        RECT 50.895 119.060 51.215 119.120 ;
        RECT 49.530 118.920 51.215 119.060 ;
        RECT 49.530 118.875 49.820 118.920 ;
        RECT 50.895 118.860 51.215 118.920 ;
        RECT 57.350 119.060 57.640 119.105 ;
        RECT 57.795 119.060 58.115 119.120 ;
        RECT 57.350 118.920 58.115 119.060 ;
        RECT 57.350 118.875 57.640 118.920 ;
        RECT 57.795 118.860 58.115 118.920 ;
        RECT 58.715 118.860 59.035 119.120 ;
        RECT 63.315 118.860 63.635 119.120 ;
        RECT 63.865 119.105 64.005 119.260 ;
        RECT 72.945 119.260 77.875 119.400 ;
        RECT 72.945 119.215 73.235 119.260 ;
        RECT 75.725 119.215 76.015 119.260 ;
        RECT 77.585 119.215 77.875 119.260 ;
        RECT 91.805 119.400 92.095 119.445 ;
        RECT 94.585 119.400 94.875 119.445 ;
        RECT 96.445 119.400 96.735 119.445 ;
        RECT 91.805 119.260 96.735 119.400 ;
        RECT 91.805 119.215 92.095 119.260 ;
        RECT 94.585 119.215 94.875 119.260 ;
        RECT 96.445 119.215 96.735 119.260 ;
        RECT 97.905 119.260 102.185 119.400 ;
        RECT 63.790 118.875 64.080 119.105 ;
        RECT 71.135 119.060 71.455 119.120 ;
        RECT 72.515 119.060 72.835 119.120 ;
        RECT 67.545 118.920 72.835 119.060 ;
        RECT 28.830 118.720 29.120 118.765 ;
        RECT 25.595 118.580 29.120 118.720 ;
        RECT 25.595 118.520 25.915 118.580 ;
        RECT 28.830 118.535 29.120 118.580 ;
        RECT 31.115 118.520 31.435 118.780 ;
        RECT 33.430 118.720 33.720 118.765 ;
        RECT 36.635 118.720 36.955 118.780 ;
        RECT 33.430 118.580 36.955 118.720 ;
        RECT 33.430 118.535 33.720 118.580 ;
        RECT 36.635 118.520 36.955 118.580 ;
        RECT 39.410 118.535 39.700 118.765 ;
        RECT 39.870 118.720 40.160 118.765 ;
        RECT 42.170 118.720 42.460 118.765 ;
        RECT 43.995 118.720 44.315 118.780 ;
        RECT 39.870 118.580 44.315 118.720 ;
        RECT 39.870 118.535 40.160 118.580 ;
        RECT 42.170 118.535 42.460 118.580 ;
        RECT 31.590 118.380 31.880 118.425 ;
        RECT 33.875 118.380 34.195 118.440 ;
        RECT 31.590 118.240 34.195 118.380 ;
        RECT 39.485 118.380 39.625 118.535 ;
        RECT 43.995 118.520 44.315 118.580 ;
        RECT 52.275 118.520 52.595 118.780 ;
        RECT 53.670 118.720 53.960 118.765 ;
        RECT 54.575 118.720 54.895 118.780 ;
        RECT 53.670 118.580 54.895 118.720 ;
        RECT 53.670 118.535 53.960 118.580 ;
        RECT 54.575 118.520 54.895 118.580 ;
        RECT 55.035 118.520 55.355 118.780 ;
        RECT 58.270 118.700 58.560 118.765 ;
        RECT 58.805 118.700 58.945 118.860 ;
        RECT 58.270 118.560 58.945 118.700 ;
        RECT 61.935 118.720 62.255 118.780 ;
        RECT 67.545 118.765 67.685 118.920 ;
        RECT 71.135 118.860 71.455 118.920 ;
        RECT 72.515 118.860 72.835 118.920 ;
        RECT 78.035 118.860 78.355 119.120 ;
        RECT 82.650 119.060 82.940 119.105 ;
        RECT 87.235 119.060 87.555 119.120 ;
        RECT 82.650 118.920 87.555 119.060 ;
        RECT 82.650 118.875 82.940 118.920 ;
        RECT 65.170 118.720 65.460 118.765 ;
        RECT 61.935 118.580 65.460 118.720 ;
        RECT 58.270 118.535 58.560 118.560 ;
        RECT 61.935 118.520 62.255 118.580 ;
        RECT 65.170 118.535 65.460 118.580 ;
        RECT 67.470 118.535 67.760 118.765 ;
        RECT 72.945 118.720 73.235 118.765 ;
        RECT 76.210 118.720 76.500 118.765 ;
        RECT 78.495 118.720 78.815 118.780 ;
        RECT 72.945 118.580 75.480 118.720 ;
        RECT 72.945 118.535 73.235 118.580 ;
        RECT 44.930 118.380 45.220 118.425 ;
        RECT 48.595 118.380 48.915 118.440 ;
        RECT 49.990 118.380 50.280 118.425 ;
        RECT 39.485 118.240 50.280 118.380 ;
        RECT 31.590 118.195 31.880 118.240 ;
        RECT 33.875 118.180 34.195 118.240 ;
        RECT 44.930 118.195 45.220 118.240 ;
        RECT 48.595 118.180 48.915 118.240 ;
        RECT 49.990 118.195 50.280 118.240 ;
        RECT 62.870 118.195 63.160 118.425 ;
        RECT 71.085 118.380 71.375 118.425 ;
        RECT 72.515 118.380 72.835 118.440 ;
        RECT 75.265 118.425 75.480 118.580 ;
        RECT 76.210 118.580 78.815 118.720 ;
        RECT 76.210 118.535 76.500 118.580 ;
        RECT 78.495 118.520 78.815 118.580 ;
        RECT 79.415 118.520 79.735 118.780 ;
        RECT 79.875 118.520 80.195 118.780 ;
        RECT 81.715 118.520 82.035 118.780 ;
        RECT 74.345 118.380 74.635 118.425 ;
        RECT 71.085 118.240 74.635 118.380 ;
        RECT 71.085 118.195 71.375 118.240 ;
        RECT 30.670 118.040 30.960 118.085 ;
        RECT 32.035 118.040 32.355 118.100 ;
        RECT 30.670 117.900 32.355 118.040 ;
        RECT 30.670 117.855 30.960 117.900 ;
        RECT 32.035 117.840 32.355 117.900 ;
        RECT 43.995 118.040 44.315 118.100 ;
        RECT 45.390 118.040 45.680 118.085 ;
        RECT 45.835 118.040 46.155 118.100 ;
        RECT 43.995 117.900 46.155 118.040 ;
        RECT 43.995 117.840 44.315 117.900 ;
        RECT 45.390 117.855 45.680 117.900 ;
        RECT 45.835 117.840 46.155 117.900 ;
        RECT 46.755 118.040 47.075 118.100 ;
        RECT 47.230 118.040 47.520 118.085 ;
        RECT 46.755 117.900 47.520 118.040 ;
        RECT 46.755 117.840 47.075 117.900 ;
        RECT 47.230 117.855 47.520 117.900 ;
        RECT 51.815 117.840 52.135 118.100 ;
        RECT 57.335 118.040 57.655 118.100 ;
        RECT 57.810 118.040 58.100 118.085 ;
        RECT 57.335 117.900 58.100 118.040 ;
        RECT 57.335 117.840 57.655 117.900 ;
        RECT 57.810 117.855 58.100 117.900 ;
        RECT 59.175 118.040 59.495 118.100 ;
        RECT 62.945 118.040 63.085 118.195 ;
        RECT 72.515 118.180 72.835 118.240 ;
        RECT 74.345 118.195 74.635 118.240 ;
        RECT 75.265 118.380 75.555 118.425 ;
        RECT 77.125 118.380 77.415 118.425 ;
        RECT 75.265 118.240 77.415 118.380 ;
        RECT 75.265 118.195 75.555 118.240 ;
        RECT 77.125 118.195 77.415 118.240 ;
        RECT 77.575 118.380 77.895 118.440 ;
        RECT 82.725 118.380 82.865 118.875 ;
        RECT 87.235 118.860 87.555 118.920 ;
        RECT 95.055 118.860 95.375 119.120 ;
        RECT 96.910 119.060 97.200 119.105 ;
        RECT 97.355 119.060 97.675 119.120 ;
        RECT 97.905 119.105 98.045 119.260 ;
        RECT 96.910 118.920 97.675 119.060 ;
        RECT 96.910 118.875 97.200 118.920 ;
        RECT 97.355 118.860 97.675 118.920 ;
        RECT 97.830 118.875 98.120 119.105 ;
        RECT 98.750 119.060 99.040 119.105 ;
        RECT 99.195 119.060 99.515 119.120 ;
        RECT 102.045 119.105 102.185 119.260 ;
        RECT 98.750 118.920 99.515 119.060 ;
        RECT 98.750 118.875 99.040 118.920 ;
        RECT 91.805 118.720 92.095 118.765 ;
        RECT 91.805 118.580 94.340 118.720 ;
        RECT 91.805 118.535 92.095 118.580 ;
        RECT 77.575 118.240 82.865 118.380 ;
        RECT 77.575 118.180 77.895 118.240 ;
        RECT 83.555 118.180 83.875 118.440 ;
        RECT 93.215 118.425 93.535 118.440 ;
        RECT 89.945 118.380 90.235 118.425 ;
        RECT 93.205 118.380 93.535 118.425 ;
        RECT 89.945 118.240 93.535 118.380 ;
        RECT 89.945 118.195 90.235 118.240 ;
        RECT 93.205 118.195 93.535 118.240 ;
        RECT 94.125 118.425 94.340 118.580 ;
        RECT 94.125 118.380 94.415 118.425 ;
        RECT 95.985 118.380 96.275 118.425 ;
        RECT 94.125 118.240 96.275 118.380 ;
        RECT 94.125 118.195 94.415 118.240 ;
        RECT 95.985 118.195 96.275 118.240 ;
        RECT 96.895 118.380 97.215 118.440 ;
        RECT 97.905 118.380 98.045 118.875 ;
        RECT 99.195 118.860 99.515 118.920 ;
        RECT 101.970 118.875 102.260 119.105 ;
        RECT 102.875 118.860 103.195 119.120 ;
        RECT 103.425 118.765 103.565 119.600 ;
        RECT 106.110 119.600 106.875 119.740 ;
        RECT 106.110 119.555 106.400 119.600 ;
        RECT 106.555 119.540 106.875 119.600 ;
        RECT 107.950 119.740 108.240 119.785 ;
        RECT 108.395 119.740 108.715 119.800 ;
        RECT 107.950 119.600 108.715 119.740 ;
        RECT 107.950 119.555 108.240 119.600 ;
        RECT 108.395 119.540 108.715 119.600 ;
        RECT 103.350 118.535 103.640 118.765 ;
        RECT 105.635 118.520 105.955 118.780 ;
        RECT 107.030 118.535 107.320 118.765 ;
        RECT 96.895 118.240 98.045 118.380 ;
        RECT 98.735 118.380 99.055 118.440 ;
        RECT 107.105 118.380 107.245 118.535 ;
        RECT 98.735 118.240 107.245 118.380 ;
        RECT 93.215 118.180 93.535 118.195 ;
        RECT 96.895 118.180 97.215 118.240 ;
        RECT 98.735 118.180 99.055 118.240 ;
        RECT 59.175 117.900 63.085 118.040 ;
        RECT 79.875 118.040 80.195 118.100 ;
        RECT 84.030 118.040 84.320 118.085 ;
        RECT 79.875 117.900 84.320 118.040 ;
        RECT 59.175 117.840 59.495 117.900 ;
        RECT 79.875 117.840 80.195 117.900 ;
        RECT 84.030 117.855 84.320 117.900 ;
        RECT 85.870 118.040 86.160 118.085 ;
        RECT 90.455 118.040 90.775 118.100 ;
        RECT 85.870 117.900 90.775 118.040 ;
        RECT 85.870 117.855 86.160 117.900 ;
        RECT 90.455 117.840 90.775 117.900 ;
        RECT 92.295 118.040 92.615 118.100 ;
        RECT 97.815 118.040 98.135 118.100 ;
        RECT 99.210 118.040 99.500 118.085 ;
        RECT 92.295 117.900 99.500 118.040 ;
        RECT 92.295 117.840 92.615 117.900 ;
        RECT 97.815 117.840 98.135 117.900 ;
        RECT 99.210 117.855 99.500 117.900 ;
        RECT 101.035 117.840 101.355 118.100 ;
        RECT 105.190 118.040 105.480 118.085 ;
        RECT 106.095 118.040 106.415 118.100 ;
        RECT 105.190 117.900 106.415 118.040 ;
        RECT 105.190 117.855 105.480 117.900 ;
        RECT 106.095 117.840 106.415 117.900 ;
        RECT 17.370 117.220 112.465 117.700 ;
        RECT 21.010 117.020 21.300 117.065 ;
        RECT 21.010 116.880 25.825 117.020 ;
        RECT 21.010 116.835 21.300 116.880 ;
        RECT 23.315 116.680 23.605 116.725 ;
        RECT 25.175 116.680 25.465 116.725 ;
        RECT 23.315 116.540 25.465 116.680 ;
        RECT 25.685 116.680 25.825 116.880 ;
        RECT 32.955 116.820 33.275 117.080 ;
        RECT 36.190 117.020 36.480 117.065 ;
        RECT 33.505 116.880 36.480 117.020 ;
        RECT 26.095 116.680 26.385 116.725 ;
        RECT 29.355 116.680 29.645 116.725 ;
        RECT 25.685 116.540 29.645 116.680 ;
        RECT 23.315 116.495 23.605 116.540 ;
        RECT 25.175 116.495 25.465 116.540 ;
        RECT 26.095 116.495 26.385 116.540 ;
        RECT 29.355 116.495 29.645 116.540 ;
        RECT 31.575 116.680 31.895 116.740 ;
        RECT 33.505 116.680 33.645 116.880 ;
        RECT 36.190 116.835 36.480 116.880 ;
        RECT 38.260 117.020 38.550 117.065 ;
        RECT 43.995 117.020 44.315 117.080 ;
        RECT 48.595 117.065 48.915 117.080 ;
        RECT 38.260 116.880 44.315 117.020 ;
        RECT 38.260 116.835 38.550 116.880 ;
        RECT 43.995 116.820 44.315 116.880 ;
        RECT 48.380 116.835 48.915 117.065 ;
        RECT 48.595 116.820 48.915 116.835 ;
        RECT 52.275 117.020 52.595 117.080 ;
        RECT 63.315 117.020 63.635 117.080 ;
        RECT 66.780 117.020 67.070 117.065 ;
        RECT 52.275 116.880 57.105 117.020 ;
        RECT 52.275 116.820 52.595 116.880 ;
        RECT 31.575 116.540 33.645 116.680 ;
        RECT 33.875 116.680 34.195 116.740 ;
        RECT 40.265 116.680 40.555 116.725 ;
        RECT 43.525 116.680 43.815 116.725 ;
        RECT 33.875 116.540 43.815 116.680 ;
        RECT 21.455 116.140 21.775 116.400 ;
        RECT 21.915 116.340 22.235 116.400 ;
        RECT 24.230 116.340 24.520 116.385 ;
        RECT 21.915 116.200 24.520 116.340 ;
        RECT 25.250 116.340 25.465 116.495 ;
        RECT 31.575 116.480 31.895 116.540 ;
        RECT 33.875 116.480 34.195 116.540 ;
        RECT 40.265 116.495 40.555 116.540 ;
        RECT 43.525 116.495 43.815 116.540 ;
        RECT 44.445 116.680 44.735 116.725 ;
        RECT 46.305 116.680 46.595 116.725 ;
        RECT 44.445 116.540 46.595 116.680 ;
        RECT 44.445 116.495 44.735 116.540 ;
        RECT 46.305 116.495 46.595 116.540 ;
        RECT 47.675 116.680 47.995 116.740 ;
        RECT 50.385 116.680 50.675 116.725 ;
        RECT 53.645 116.680 53.935 116.725 ;
        RECT 47.675 116.540 53.935 116.680 ;
        RECT 27.495 116.340 27.785 116.385 ;
        RECT 25.250 116.200 27.785 116.340 ;
        RECT 21.915 116.140 22.235 116.200 ;
        RECT 24.230 116.155 24.520 116.200 ;
        RECT 27.495 116.155 27.785 116.200 ;
        RECT 31.115 116.340 31.435 116.400 ;
        RECT 32.510 116.340 32.800 116.385 ;
        RECT 35.730 116.340 36.020 116.385 ;
        RECT 41.235 116.340 41.555 116.400 ;
        RECT 31.115 116.200 33.185 116.340 ;
        RECT 31.115 116.140 31.435 116.200 ;
        RECT 32.510 116.155 32.800 116.200 ;
        RECT 22.390 116.000 22.680 116.045 ;
        RECT 22.390 115.860 32.725 116.000 ;
        RECT 22.390 115.815 22.680 115.860 ;
        RECT 32.585 115.720 32.725 115.860 ;
        RECT 22.855 115.660 23.145 115.705 ;
        RECT 24.715 115.660 25.005 115.705 ;
        RECT 27.495 115.660 27.785 115.705 ;
        RECT 22.855 115.520 27.785 115.660 ;
        RECT 22.855 115.475 23.145 115.520 ;
        RECT 24.715 115.475 25.005 115.520 ;
        RECT 27.495 115.475 27.785 115.520 ;
        RECT 32.495 115.460 32.815 115.720 ;
        RECT 33.045 115.660 33.185 116.200 ;
        RECT 35.730 116.200 41.555 116.340 ;
        RECT 35.730 116.155 36.020 116.200 ;
        RECT 41.235 116.140 41.555 116.200 ;
        RECT 42.125 116.340 42.415 116.385 ;
        RECT 44.445 116.340 44.660 116.495 ;
        RECT 47.675 116.480 47.995 116.540 ;
        RECT 50.385 116.495 50.675 116.540 ;
        RECT 53.645 116.495 53.935 116.540 ;
        RECT 54.565 116.680 54.855 116.725 ;
        RECT 56.425 116.680 56.715 116.725 ;
        RECT 54.565 116.540 56.715 116.680 ;
        RECT 54.565 116.495 54.855 116.540 ;
        RECT 56.425 116.495 56.715 116.540 ;
        RECT 52.245 116.340 52.535 116.385 ;
        RECT 54.565 116.340 54.780 116.495 ;
        RECT 42.125 116.200 44.660 116.340 ;
        RECT 45.005 116.200 46.525 116.340 ;
        RECT 42.125 116.155 42.415 116.200 ;
        RECT 36.635 116.000 36.955 116.060 ;
        RECT 45.005 116.000 45.145 116.200 ;
        RECT 46.385 116.060 46.525 116.200 ;
        RECT 52.245 116.200 54.780 116.340 ;
        RECT 55.510 116.340 55.800 116.385 ;
        RECT 56.965 116.340 57.105 116.880 ;
        RECT 63.315 116.880 67.070 117.020 ;
        RECT 63.315 116.820 63.635 116.880 ;
        RECT 66.780 116.835 67.070 116.880 ;
        RECT 67.455 116.820 67.775 117.080 ;
        RECT 72.515 116.820 72.835 117.080 ;
        RECT 88.170 116.835 88.460 117.065 ;
        RECT 100.575 117.020 100.895 117.080 ;
        RECT 101.740 117.020 102.030 117.065 ;
        RECT 100.575 116.880 102.030 117.020 ;
        RECT 58.735 116.680 59.025 116.725 ;
        RECT 60.595 116.680 60.885 116.725 ;
        RECT 58.735 116.540 60.885 116.680 ;
        RECT 58.735 116.495 59.025 116.540 ;
        RECT 60.595 116.495 60.885 116.540 ;
        RECT 61.515 116.680 61.805 116.725 ;
        RECT 62.395 116.680 62.715 116.740 ;
        RECT 64.775 116.680 65.065 116.725 ;
        RECT 61.515 116.540 65.065 116.680 ;
        RECT 61.515 116.495 61.805 116.540 ;
        RECT 55.510 116.200 57.105 116.340 ;
        RECT 52.245 116.155 52.535 116.200 ;
        RECT 55.510 116.155 55.800 116.200 ;
        RECT 59.635 116.140 59.955 116.400 ;
        RECT 60.095 116.140 60.415 116.400 ;
        RECT 60.670 116.340 60.885 116.495 ;
        RECT 62.395 116.480 62.715 116.540 ;
        RECT 64.775 116.495 65.065 116.540 ;
        RECT 70.215 116.680 70.535 116.740 ;
        RECT 75.275 116.680 75.595 116.740 ;
        RECT 76.210 116.680 76.500 116.725 ;
        RECT 78.740 116.680 79.030 116.725 ;
        RECT 79.875 116.680 80.195 116.740 ;
        RECT 70.215 116.540 75.045 116.680 ;
        RECT 70.215 116.480 70.535 116.540 ;
        RECT 62.915 116.340 63.205 116.385 ;
        RECT 60.670 116.200 63.205 116.340 ;
        RECT 62.915 116.155 63.205 116.200 ;
        RECT 68.390 116.155 68.680 116.385 ;
        RECT 69.310 116.155 69.600 116.385 ;
        RECT 69.755 116.340 70.075 116.400 ;
        RECT 70.690 116.340 70.980 116.385 ;
        RECT 72.070 116.340 72.360 116.385 ;
        RECT 72.515 116.340 72.835 116.400 ;
        RECT 69.755 116.200 72.835 116.340 ;
        RECT 36.635 115.860 45.145 116.000 ;
        RECT 45.390 116.000 45.680 116.045 ;
        RECT 45.835 116.000 46.155 116.060 ;
        RECT 45.390 115.860 46.155 116.000 ;
        RECT 36.635 115.800 36.955 115.860 ;
        RECT 45.390 115.815 45.680 115.860 ;
        RECT 45.835 115.800 46.155 115.860 ;
        RECT 46.295 115.800 46.615 116.060 ;
        RECT 47.230 116.000 47.520 116.045 ;
        RECT 57.350 116.000 57.640 116.045 ;
        RECT 57.810 116.000 58.100 116.045 ;
        RECT 60.185 116.000 60.325 116.140 ;
        RECT 47.230 115.860 60.325 116.000 ;
        RECT 60.555 116.000 60.875 116.060 ;
        RECT 68.465 116.000 68.605 116.155 ;
        RECT 60.555 115.860 68.605 116.000 ;
        RECT 69.385 116.000 69.525 116.155 ;
        RECT 69.755 116.140 70.075 116.200 ;
        RECT 70.690 116.155 70.980 116.200 ;
        RECT 72.070 116.155 72.360 116.200 ;
        RECT 72.515 116.140 72.835 116.200 ;
        RECT 74.905 116.000 75.045 116.540 ;
        RECT 75.275 116.540 80.195 116.680 ;
        RECT 75.275 116.480 75.595 116.540 ;
        RECT 76.210 116.495 76.500 116.540 ;
        RECT 78.740 116.495 79.030 116.540 ;
        RECT 79.875 116.480 80.195 116.540 ;
        RECT 80.745 116.680 81.035 116.725 ;
        RECT 83.095 116.680 83.415 116.740 ;
        RECT 84.005 116.680 84.295 116.725 ;
        RECT 80.745 116.540 84.295 116.680 ;
        RECT 80.745 116.495 81.035 116.540 ;
        RECT 83.095 116.480 83.415 116.540 ;
        RECT 84.005 116.495 84.295 116.540 ;
        RECT 84.925 116.680 85.215 116.725 ;
        RECT 86.785 116.680 87.075 116.725 ;
        RECT 84.925 116.540 87.075 116.680 ;
        RECT 84.925 116.495 85.215 116.540 ;
        RECT 86.785 116.495 87.075 116.540 ;
        RECT 75.735 116.340 76.055 116.400 ;
        RECT 79.415 116.340 79.735 116.400 ;
        RECT 75.735 116.200 79.735 116.340 ;
        RECT 75.735 116.140 76.055 116.200 ;
        RECT 79.415 116.140 79.735 116.200 ;
        RECT 82.605 116.340 82.895 116.385 ;
        RECT 84.925 116.340 85.140 116.495 ;
        RECT 82.605 116.200 85.140 116.340 ;
        RECT 85.870 116.340 86.160 116.385 ;
        RECT 88.245 116.340 88.385 116.835 ;
        RECT 100.575 116.820 100.895 116.880 ;
        RECT 101.740 116.835 102.030 116.880 ;
        RECT 91.785 116.680 92.075 116.725 ;
        RECT 94.135 116.680 94.455 116.740 ;
        RECT 95.045 116.680 95.335 116.725 ;
        RECT 91.785 116.540 95.335 116.680 ;
        RECT 91.785 116.495 92.075 116.540 ;
        RECT 94.135 116.480 94.455 116.540 ;
        RECT 95.045 116.495 95.335 116.540 ;
        RECT 95.965 116.680 96.255 116.725 ;
        RECT 97.825 116.680 98.115 116.725 ;
        RECT 95.965 116.540 98.115 116.680 ;
        RECT 95.965 116.495 96.255 116.540 ;
        RECT 97.825 116.495 98.115 116.540 ;
        RECT 103.745 116.680 104.035 116.725 ;
        RECT 104.715 116.680 105.035 116.740 ;
        RECT 107.005 116.680 107.295 116.725 ;
        RECT 103.745 116.540 107.295 116.680 ;
        RECT 103.745 116.495 104.035 116.540 ;
        RECT 85.870 116.200 88.385 116.340 ;
        RECT 89.090 116.340 89.380 116.385 ;
        RECT 90.455 116.340 90.775 116.400 ;
        RECT 89.090 116.200 90.775 116.340 ;
        RECT 82.605 116.155 82.895 116.200 ;
        RECT 85.870 116.155 86.160 116.200 ;
        RECT 89.090 116.155 89.380 116.200 ;
        RECT 90.455 116.140 90.775 116.200 ;
        RECT 93.645 116.340 93.935 116.385 ;
        RECT 95.965 116.340 96.180 116.495 ;
        RECT 104.715 116.480 105.035 116.540 ;
        RECT 107.005 116.495 107.295 116.540 ;
        RECT 107.925 116.680 108.215 116.725 ;
        RECT 109.785 116.680 110.075 116.725 ;
        RECT 107.925 116.540 110.075 116.680 ;
        RECT 107.925 116.495 108.215 116.540 ;
        RECT 109.785 116.495 110.075 116.540 ;
        RECT 93.645 116.200 96.180 116.340 ;
        RECT 97.355 116.340 97.675 116.400 ;
        RECT 98.750 116.340 99.040 116.385 ;
        RECT 97.355 116.200 99.040 116.340 ;
        RECT 93.645 116.155 93.935 116.200 ;
        RECT 97.355 116.140 97.675 116.200 ;
        RECT 98.750 116.155 99.040 116.200 ;
        RECT 101.035 116.140 101.355 116.400 ;
        RECT 105.605 116.340 105.895 116.385 ;
        RECT 107.925 116.340 108.140 116.495 ;
        RECT 105.605 116.200 108.140 116.340 ;
        RECT 105.605 116.155 105.895 116.200 ;
        RECT 110.695 116.140 111.015 116.400 ;
        RECT 76.670 116.000 76.960 116.045 ;
        RECT 77.575 116.000 77.895 116.060 ;
        RECT 69.385 115.860 74.125 116.000 ;
        RECT 74.905 115.860 77.895 116.000 ;
        RECT 47.230 115.815 47.520 115.860 ;
        RECT 57.350 115.815 57.640 115.860 ;
        RECT 57.810 115.815 58.100 115.860 ;
        RECT 60.555 115.800 60.875 115.860 ;
        RECT 38.475 115.660 38.795 115.720 ;
        RECT 73.985 115.705 74.125 115.860 ;
        RECT 76.670 115.815 76.960 115.860 ;
        RECT 77.575 115.800 77.895 115.860 ;
        RECT 78.035 116.000 78.355 116.060 ;
        RECT 87.710 116.000 88.000 116.045 ;
        RECT 78.035 115.860 88.000 116.000 ;
        RECT 78.035 115.800 78.355 115.860 ;
        RECT 87.710 115.815 88.000 115.860 ;
        RECT 96.910 116.000 97.200 116.045 ;
        RECT 96.910 115.860 100.345 116.000 ;
        RECT 96.910 115.815 97.200 115.860 ;
        RECT 100.205 115.705 100.345 115.860 ;
        RECT 108.855 115.800 109.175 116.060 ;
        RECT 33.045 115.520 38.795 115.660 ;
        RECT 38.475 115.460 38.795 115.520 ;
        RECT 42.125 115.660 42.415 115.705 ;
        RECT 44.905 115.660 45.195 115.705 ;
        RECT 46.765 115.660 47.055 115.705 ;
        RECT 42.125 115.520 47.055 115.660 ;
        RECT 42.125 115.475 42.415 115.520 ;
        RECT 44.905 115.475 45.195 115.520 ;
        RECT 46.765 115.475 47.055 115.520 ;
        RECT 52.245 115.660 52.535 115.705 ;
        RECT 55.025 115.660 55.315 115.705 ;
        RECT 56.885 115.660 57.175 115.705 ;
        RECT 52.245 115.520 57.175 115.660 ;
        RECT 52.245 115.475 52.535 115.520 ;
        RECT 55.025 115.475 55.315 115.520 ;
        RECT 56.885 115.475 57.175 115.520 ;
        RECT 58.275 115.660 58.565 115.705 ;
        RECT 60.135 115.660 60.425 115.705 ;
        RECT 62.915 115.660 63.205 115.705 ;
        RECT 58.275 115.520 63.205 115.660 ;
        RECT 58.275 115.475 58.565 115.520 ;
        RECT 60.135 115.475 60.425 115.520 ;
        RECT 62.915 115.475 63.205 115.520 ;
        RECT 71.150 115.660 71.440 115.705 ;
        RECT 71.150 115.520 73.665 115.660 ;
        RECT 71.150 115.475 71.440 115.520 ;
        RECT 28.355 115.320 28.675 115.380 ;
        RECT 31.575 115.365 31.895 115.380 ;
        RECT 31.360 115.320 31.895 115.365 ;
        RECT 28.355 115.180 31.895 115.320 ;
        RECT 28.355 115.120 28.675 115.180 ;
        RECT 31.360 115.135 31.895 115.180 ;
        RECT 31.575 115.120 31.895 115.135 ;
        RECT 33.415 115.320 33.735 115.380 ;
        RECT 33.890 115.320 34.180 115.365 ;
        RECT 33.415 115.180 34.180 115.320 ;
        RECT 33.415 115.120 33.735 115.180 ;
        RECT 33.890 115.135 34.180 115.180 ;
        RECT 35.715 115.320 36.035 115.380 ;
        RECT 69.755 115.320 70.075 115.380 ;
        RECT 35.715 115.180 70.075 115.320 ;
        RECT 35.715 115.120 36.035 115.180 ;
        RECT 69.755 115.120 70.075 115.180 ;
        RECT 70.230 115.320 70.520 115.365 ;
        RECT 72.055 115.320 72.375 115.380 ;
        RECT 70.230 115.180 72.375 115.320 ;
        RECT 73.525 115.320 73.665 115.520 ;
        RECT 73.910 115.475 74.200 115.705 ;
        RECT 82.605 115.660 82.895 115.705 ;
        RECT 85.385 115.660 85.675 115.705 ;
        RECT 87.245 115.660 87.535 115.705 ;
        RECT 82.605 115.520 87.535 115.660 ;
        RECT 82.605 115.475 82.895 115.520 ;
        RECT 85.385 115.475 85.675 115.520 ;
        RECT 87.245 115.475 87.535 115.520 ;
        RECT 93.645 115.660 93.935 115.705 ;
        RECT 96.425 115.660 96.715 115.705 ;
        RECT 98.285 115.660 98.575 115.705 ;
        RECT 93.645 115.520 98.575 115.660 ;
        RECT 93.645 115.475 93.935 115.520 ;
        RECT 96.425 115.475 96.715 115.520 ;
        RECT 98.285 115.475 98.575 115.520 ;
        RECT 100.130 115.475 100.420 115.705 ;
        RECT 105.605 115.660 105.895 115.705 ;
        RECT 108.385 115.660 108.675 115.705 ;
        RECT 110.245 115.660 110.535 115.705 ;
        RECT 105.605 115.520 110.535 115.660 ;
        RECT 105.605 115.475 105.895 115.520 ;
        RECT 108.385 115.475 108.675 115.520 ;
        RECT 110.245 115.475 110.535 115.520 ;
        RECT 75.735 115.320 76.055 115.380 ;
        RECT 73.525 115.180 76.055 115.320 ;
        RECT 70.230 115.135 70.520 115.180 ;
        RECT 72.055 115.120 72.375 115.180 ;
        RECT 75.735 115.120 76.055 115.180 ;
        RECT 89.780 115.320 90.070 115.365 ;
        RECT 92.295 115.320 92.615 115.380 ;
        RECT 89.780 115.180 92.615 115.320 ;
        RECT 89.780 115.135 90.070 115.180 ;
        RECT 92.295 115.120 92.615 115.180 ;
        RECT 18.165 114.500 112.465 114.980 ;
        RECT 20.550 114.300 20.840 114.345 ;
        RECT 21.915 114.300 22.235 114.360 ;
        RECT 20.550 114.160 22.235 114.300 ;
        RECT 20.550 114.115 20.840 114.160 ;
        RECT 21.915 114.100 22.235 114.160 ;
        RECT 26.055 114.300 26.375 114.360 ;
        RECT 36.635 114.300 36.955 114.360 ;
        RECT 26.055 114.160 36.955 114.300 ;
        RECT 26.055 114.100 26.375 114.160 ;
        RECT 36.635 114.100 36.955 114.160 ;
        RECT 45.835 114.100 46.155 114.360 ;
        RECT 48.840 114.300 49.130 114.345 ;
        RECT 50.895 114.300 51.215 114.360 ;
        RECT 48.840 114.160 51.215 114.300 ;
        RECT 48.840 114.115 49.130 114.160 ;
        RECT 50.895 114.100 51.215 114.160 ;
        RECT 61.950 114.300 62.240 114.345 ;
        RECT 62.395 114.300 62.715 114.360 ;
        RECT 61.950 114.160 62.715 114.300 ;
        RECT 61.950 114.115 62.240 114.160 ;
        RECT 62.395 114.100 62.715 114.160 ;
        RECT 72.975 114.300 73.295 114.360 ;
        RECT 79.415 114.345 79.735 114.360 ;
        RECT 72.975 114.160 75.965 114.300 ;
        RECT 72.975 114.100 73.295 114.160 ;
        RECT 26.485 113.960 26.775 114.005 ;
        RECT 29.265 113.960 29.555 114.005 ;
        RECT 31.125 113.960 31.415 114.005 ;
        RECT 26.485 113.820 31.415 113.960 ;
        RECT 26.485 113.775 26.775 113.820 ;
        RECT 29.265 113.775 29.555 113.820 ;
        RECT 31.125 113.775 31.415 113.820 ;
        RECT 35.735 113.960 36.025 114.005 ;
        RECT 37.595 113.960 37.885 114.005 ;
        RECT 40.375 113.960 40.665 114.005 ;
        RECT 35.735 113.820 40.665 113.960 ;
        RECT 35.735 113.775 36.025 113.820 ;
        RECT 37.595 113.775 37.885 113.820 ;
        RECT 40.375 113.775 40.665 113.820 ;
        RECT 52.705 113.960 52.995 114.005 ;
        RECT 55.485 113.960 55.775 114.005 ;
        RECT 57.345 113.960 57.635 114.005 ;
        RECT 52.705 113.820 57.635 113.960 ;
        RECT 52.705 113.775 52.995 113.820 ;
        RECT 55.485 113.775 55.775 113.820 ;
        RECT 57.345 113.775 57.635 113.820 ;
        RECT 70.695 113.960 70.985 114.005 ;
        RECT 72.555 113.960 72.845 114.005 ;
        RECT 75.335 113.960 75.625 114.005 ;
        RECT 70.695 113.820 75.625 113.960 ;
        RECT 70.695 113.775 70.985 113.820 ;
        RECT 72.555 113.775 72.845 113.820 ;
        RECT 75.335 113.775 75.625 113.820 ;
        RECT 32.495 113.620 32.815 113.680 ;
        RECT 57.810 113.620 58.100 113.665 ;
        RECT 60.095 113.620 60.415 113.680 ;
        RECT 31.665 113.480 35.485 113.620 ;
        RECT 19.630 113.095 19.920 113.325 ;
        RECT 19.705 112.940 19.845 113.095 ;
        RECT 21.915 113.080 22.235 113.340 ;
        RECT 22.620 113.280 22.910 113.325 ;
        RECT 25.595 113.280 25.915 113.340 ;
        RECT 31.665 113.325 31.805 113.480 ;
        RECT 32.495 113.420 32.815 113.480 ;
        RECT 22.620 113.140 25.915 113.280 ;
        RECT 22.620 113.095 22.910 113.140 ;
        RECT 25.595 113.080 25.915 113.140 ;
        RECT 26.485 113.280 26.775 113.325 ;
        RECT 29.750 113.280 30.040 113.325 ;
        RECT 26.485 113.140 29.020 113.280 ;
        RECT 26.485 113.095 26.775 113.140 ;
        RECT 23.295 112.940 23.615 113.000 ;
        RECT 28.805 112.985 29.020 113.140 ;
        RECT 29.750 113.140 31.345 113.280 ;
        RECT 29.750 113.095 30.040 113.140 ;
        RECT 24.625 112.940 24.915 112.985 ;
        RECT 27.885 112.940 28.175 112.985 ;
        RECT 19.705 112.800 23.615 112.940 ;
        RECT 23.295 112.740 23.615 112.800 ;
        RECT 24.305 112.800 28.175 112.940 ;
        RECT 21.470 112.600 21.760 112.645 ;
        RECT 24.305 112.600 24.445 112.800 ;
        RECT 24.625 112.755 24.915 112.800 ;
        RECT 27.885 112.755 28.175 112.800 ;
        RECT 28.805 112.940 29.095 112.985 ;
        RECT 30.665 112.940 30.955 112.985 ;
        RECT 28.805 112.800 30.955 112.940 ;
        RECT 31.205 112.940 31.345 113.140 ;
        RECT 31.590 113.095 31.880 113.325 ;
        RECT 32.035 113.280 32.355 113.340 ;
        RECT 32.970 113.280 33.260 113.325 ;
        RECT 32.035 113.140 33.260 113.280 ;
        RECT 32.035 113.080 32.355 113.140 ;
        RECT 32.970 113.095 33.260 113.140 ;
        RECT 33.415 113.080 33.735 113.340 ;
        RECT 35.345 113.325 35.485 113.480 ;
        RECT 57.810 113.480 60.415 113.620 ;
        RECT 57.810 113.435 58.100 113.480 ;
        RECT 60.095 113.420 60.415 113.480 ;
        RECT 72.055 113.420 72.375 113.680 ;
        RECT 73.895 113.620 74.215 113.680 ;
        RECT 72.605 113.480 74.215 113.620 ;
        RECT 35.270 113.280 35.560 113.325 ;
        RECT 36.635 113.280 36.955 113.340 ;
        RECT 35.270 113.140 36.955 113.280 ;
        RECT 35.270 113.095 35.560 113.140 ;
        RECT 36.635 113.080 36.955 113.140 ;
        RECT 37.110 113.280 37.400 113.325 ;
        RECT 37.555 113.280 37.875 113.340 ;
        RECT 40.375 113.280 40.665 113.325 ;
        RECT 37.110 113.140 37.875 113.280 ;
        RECT 37.110 113.095 37.400 113.140 ;
        RECT 37.555 113.080 37.875 113.140 ;
        RECT 38.130 113.140 40.665 113.280 ;
        RECT 38.130 112.985 38.345 113.140 ;
        RECT 40.375 113.095 40.665 113.140 ;
        RECT 41.235 113.280 41.555 113.340 ;
        RECT 43.535 113.280 43.855 113.340 ;
        RECT 44.240 113.280 44.530 113.325 ;
        RECT 41.235 113.140 44.530 113.280 ;
        RECT 41.235 113.080 41.555 113.140 ;
        RECT 43.535 113.080 43.855 113.140 ;
        RECT 44.240 113.095 44.530 113.140 ;
        RECT 46.755 113.080 47.075 113.340 ;
        RECT 47.215 113.080 47.535 113.340 ;
        RECT 47.675 113.080 47.995 113.340 ;
        RECT 52.705 113.280 52.995 113.325 ;
        RECT 52.705 113.140 55.240 113.280 ;
        RECT 52.705 113.095 52.995 113.140 ;
        RECT 36.195 112.940 36.485 112.985 ;
        RECT 38.055 112.940 38.345 112.985 ;
        RECT 31.205 112.800 32.265 112.940 ;
        RECT 28.805 112.755 29.095 112.800 ;
        RECT 30.665 112.755 30.955 112.800 ;
        RECT 32.125 112.645 32.265 112.800 ;
        RECT 36.195 112.800 38.345 112.940 ;
        RECT 36.195 112.755 36.485 112.800 ;
        RECT 38.055 112.755 38.345 112.800 ;
        RECT 38.935 112.985 39.255 113.000 ;
        RECT 50.895 112.985 51.215 113.000 ;
        RECT 55.025 112.985 55.240 113.140 ;
        RECT 55.955 113.080 56.275 113.340 ;
        RECT 61.490 113.095 61.780 113.325 ;
        RECT 62.855 113.280 63.175 113.340 ;
        RECT 69.310 113.280 69.600 113.325 ;
        RECT 62.855 113.140 69.600 113.280 ;
        RECT 38.935 112.940 39.265 112.985 ;
        RECT 42.235 112.940 42.525 112.985 ;
        RECT 38.935 112.800 42.525 112.940 ;
        RECT 38.935 112.755 39.265 112.800 ;
        RECT 42.235 112.755 42.525 112.800 ;
        RECT 50.845 112.940 51.215 112.985 ;
        RECT 54.105 112.940 54.395 112.985 ;
        RECT 50.845 112.800 54.395 112.940 ;
        RECT 50.845 112.755 51.215 112.800 ;
        RECT 54.105 112.755 54.395 112.800 ;
        RECT 55.025 112.940 55.315 112.985 ;
        RECT 56.885 112.940 57.175 112.985 ;
        RECT 55.025 112.800 57.175 112.940 ;
        RECT 55.025 112.755 55.315 112.800 ;
        RECT 56.885 112.755 57.175 112.800 ;
        RECT 57.335 112.940 57.655 113.000 ;
        RECT 61.565 112.940 61.705 113.095 ;
        RECT 62.855 113.080 63.175 113.140 ;
        RECT 69.310 113.095 69.600 113.140 ;
        RECT 69.755 113.080 70.075 113.340 ;
        RECT 70.230 113.280 70.520 113.325 ;
        RECT 72.605 113.280 72.745 113.480 ;
        RECT 73.895 113.420 74.215 113.480 ;
        RECT 75.335 113.280 75.625 113.325 ;
        RECT 70.230 113.140 72.745 113.280 ;
        RECT 73.090 113.140 75.625 113.280 ;
        RECT 75.825 113.280 75.965 114.160 ;
        RECT 79.200 114.115 79.735 114.345 ;
        RECT 79.415 114.100 79.735 114.115 ;
        RECT 83.555 114.300 83.875 114.360 ;
        RECT 87.020 114.300 87.310 114.345 ;
        RECT 83.555 114.160 87.310 114.300 ;
        RECT 83.555 114.100 83.875 114.160 ;
        RECT 87.020 114.115 87.310 114.160 ;
        RECT 104.715 114.100 105.035 114.360 ;
        RECT 78.495 113.960 78.815 114.020 ;
        RECT 79.890 113.960 80.180 114.005 ;
        RECT 78.495 113.820 80.180 113.960 ;
        RECT 78.495 113.760 78.815 113.820 ;
        RECT 79.890 113.775 80.180 113.820 ;
        RECT 90.885 113.960 91.175 114.005 ;
        RECT 93.665 113.960 93.955 114.005 ;
        RECT 95.525 113.960 95.815 114.005 ;
        RECT 90.885 113.820 95.815 113.960 ;
        RECT 90.885 113.775 91.175 113.820 ;
        RECT 93.665 113.775 93.955 113.820 ;
        RECT 95.525 113.775 95.815 113.820 ;
        RECT 97.355 113.760 97.675 114.020 ;
        RECT 95.990 113.620 96.280 113.665 ;
        RECT 97.445 113.620 97.585 113.760 ;
        RECT 95.990 113.480 97.585 113.620 ;
        RECT 95.990 113.435 96.280 113.480 ;
        RECT 80.810 113.280 81.100 113.325 ;
        RECT 82.190 113.280 82.480 113.325 ;
        RECT 75.825 113.140 81.100 113.280 ;
        RECT 70.230 113.095 70.520 113.140 ;
        RECT 70.675 112.940 70.995 113.000 ;
        RECT 73.090 112.985 73.305 113.140 ;
        RECT 75.335 113.095 75.625 113.140 ;
        RECT 80.810 113.095 81.100 113.140 ;
        RECT 81.345 113.140 82.480 113.280 ;
        RECT 57.335 112.800 70.995 112.940 ;
        RECT 38.935 112.740 39.255 112.755 ;
        RECT 50.895 112.740 51.215 112.755 ;
        RECT 57.335 112.740 57.655 112.800 ;
        RECT 70.675 112.740 70.995 112.800 ;
        RECT 71.155 112.940 71.445 112.985 ;
        RECT 73.015 112.940 73.305 112.985 ;
        RECT 71.155 112.800 73.305 112.940 ;
        RECT 71.155 112.755 71.445 112.800 ;
        RECT 73.015 112.755 73.305 112.800 ;
        RECT 73.935 112.940 74.225 112.985 ;
        RECT 75.735 112.940 76.055 113.000 ;
        RECT 77.195 112.940 77.485 112.985 ;
        RECT 73.935 112.800 77.485 112.940 ;
        RECT 73.935 112.755 74.225 112.800 ;
        RECT 75.735 112.740 76.055 112.800 ;
        RECT 77.195 112.755 77.485 112.800 ;
        RECT 21.470 112.460 24.445 112.600 ;
        RECT 21.470 112.415 21.760 112.460 ;
        RECT 32.050 112.415 32.340 112.645 ;
        RECT 34.350 112.600 34.640 112.645 ;
        RECT 37.555 112.600 37.875 112.660 ;
        RECT 34.350 112.460 37.875 112.600 ;
        RECT 34.350 112.415 34.640 112.460 ;
        RECT 37.555 112.400 37.875 112.460 ;
        RECT 38.475 112.600 38.795 112.660 ;
        RECT 47.215 112.600 47.535 112.660 ;
        RECT 38.475 112.460 47.535 112.600 ;
        RECT 38.475 112.400 38.795 112.460 ;
        RECT 47.215 112.400 47.535 112.460 ;
        RECT 72.515 112.600 72.835 112.660 ;
        RECT 81.345 112.600 81.485 113.140 ;
        RECT 82.190 113.095 82.480 113.140 ;
        RECT 83.095 113.080 83.415 113.340 ;
        RECT 83.570 113.280 83.860 113.325 ;
        RECT 84.950 113.280 85.240 113.325 ;
        RECT 83.570 113.140 85.240 113.280 ;
        RECT 83.570 113.095 83.860 113.140 ;
        RECT 84.950 113.095 85.240 113.140 ;
        RECT 90.885 113.280 91.175 113.325 ;
        RECT 94.150 113.280 94.440 113.325 ;
        RECT 96.895 113.280 97.215 113.340 ;
        RECT 97.370 113.280 97.660 113.325 ;
        RECT 90.885 113.140 93.420 113.280 ;
        RECT 90.885 113.095 91.175 113.140 ;
        RECT 81.730 112.940 82.020 112.985 ;
        RECT 82.635 112.940 82.955 113.000 ;
        RECT 83.645 112.940 83.785 113.095 ;
        RECT 93.205 112.985 93.420 113.140 ;
        RECT 94.150 113.140 96.665 113.280 ;
        RECT 94.150 113.095 94.440 113.140 ;
        RECT 81.730 112.800 82.955 112.940 ;
        RECT 81.730 112.755 82.020 112.800 ;
        RECT 82.635 112.740 82.955 112.800 ;
        RECT 83.185 112.800 83.785 112.940 ;
        RECT 85.410 112.940 85.700 112.985 ;
        RECT 89.025 112.940 89.315 112.985 ;
        RECT 92.285 112.940 92.575 112.985 ;
        RECT 85.410 112.800 92.575 112.940 ;
        RECT 83.185 112.600 83.325 112.800 ;
        RECT 85.410 112.755 85.700 112.800 ;
        RECT 89.025 112.755 89.315 112.800 ;
        RECT 92.285 112.755 92.575 112.800 ;
        RECT 93.205 112.940 93.495 112.985 ;
        RECT 95.065 112.940 95.355 112.985 ;
        RECT 93.205 112.800 95.355 112.940 ;
        RECT 93.205 112.755 93.495 112.800 ;
        RECT 95.065 112.755 95.355 112.800 ;
        RECT 96.525 112.645 96.665 113.140 ;
        RECT 96.895 113.140 97.660 113.280 ;
        RECT 96.895 113.080 97.215 113.140 ;
        RECT 97.370 113.095 97.660 113.140 ;
        RECT 104.270 113.280 104.560 113.325 ;
        RECT 105.635 113.280 105.955 113.340 ;
        RECT 104.270 113.140 105.955 113.280 ;
        RECT 104.270 113.095 104.560 113.140 ;
        RECT 105.635 113.080 105.955 113.140 ;
        RECT 106.095 113.080 106.415 113.340 ;
        RECT 72.515 112.460 83.325 112.600 ;
        RECT 72.515 112.400 72.835 112.460 ;
        RECT 96.450 112.415 96.740 112.645 ;
        RECT 107.030 112.600 107.320 112.645 ;
        RECT 108.855 112.600 109.175 112.660 ;
        RECT 107.030 112.460 109.175 112.600 ;
        RECT 107.030 112.415 107.320 112.460 ;
        RECT 108.855 112.400 109.175 112.460 ;
        RECT 17.370 111.780 112.465 112.260 ;
        RECT 23.295 111.380 23.615 111.640 ;
        RECT 25.595 111.380 25.915 111.640 ;
        RECT 27.910 111.580 28.200 111.625 ;
        RECT 38.935 111.580 39.255 111.640 ;
        RECT 27.910 111.440 39.255 111.580 ;
        RECT 27.910 111.395 28.200 111.440 ;
        RECT 38.935 111.380 39.255 111.440 ;
        RECT 50.895 111.380 51.215 111.640 ;
        RECT 52.275 111.580 52.595 111.640 ;
        RECT 52.750 111.580 53.040 111.625 ;
        RECT 52.275 111.440 53.040 111.580 ;
        RECT 52.275 111.380 52.595 111.440 ;
        RECT 52.750 111.395 53.040 111.440 ;
        RECT 60.095 111.580 60.415 111.640 ;
        RECT 66.535 111.580 66.855 111.640 ;
        RECT 60.095 111.440 66.305 111.580 ;
        RECT 60.095 111.380 60.415 111.440 ;
        RECT 21.915 111.240 22.235 111.300 ;
        RECT 25.150 111.240 25.440 111.285 ;
        RECT 28.355 111.240 28.675 111.300 ;
        RECT 21.915 111.100 24.445 111.240 ;
        RECT 21.915 111.040 22.235 111.100 ;
        RECT 20.550 110.900 20.840 110.945 ;
        RECT 23.755 110.900 24.075 110.960 ;
        RECT 20.550 110.760 24.075 110.900 ;
        RECT 24.305 110.900 24.445 111.100 ;
        RECT 25.150 111.100 28.675 111.240 ;
        RECT 25.150 111.055 25.440 111.100 ;
        RECT 28.355 111.040 28.675 111.100 ;
        RECT 28.815 111.240 29.135 111.300 ;
        RECT 31.690 111.240 31.980 111.285 ;
        RECT 34.930 111.240 35.580 111.285 ;
        RECT 28.815 111.100 35.580 111.240 ;
        RECT 28.815 111.040 29.135 111.100 ;
        RECT 31.690 111.055 32.280 111.100 ;
        RECT 34.930 111.055 35.580 111.100 ;
        RECT 47.215 111.240 47.535 111.300 ;
        RECT 54.130 111.240 54.420 111.285 ;
        RECT 47.215 111.100 54.420 111.240 ;
        RECT 27.450 110.900 27.740 110.945 ;
        RECT 30.655 110.900 30.975 110.960 ;
        RECT 24.305 110.760 30.975 110.900 ;
        RECT 20.550 110.715 20.840 110.760 ;
        RECT 23.755 110.700 24.075 110.760 ;
        RECT 27.450 110.715 27.740 110.760 ;
        RECT 30.655 110.700 30.975 110.760 ;
        RECT 31.990 110.740 32.280 111.055 ;
        RECT 47.215 111.040 47.535 111.100 ;
        RECT 33.070 110.900 33.360 110.945 ;
        RECT 36.650 110.900 36.940 110.945 ;
        RECT 38.485 110.900 38.775 110.945 ;
        RECT 33.070 110.760 38.775 110.900 ;
        RECT 33.070 110.715 33.360 110.760 ;
        RECT 36.650 110.715 36.940 110.760 ;
        RECT 38.485 110.715 38.775 110.760 ;
        RECT 40.315 110.900 40.635 110.960 ;
        RECT 50.525 110.945 50.665 111.100 ;
        RECT 54.130 111.055 54.420 111.100 ;
        RECT 58.830 111.240 59.120 111.285 ;
        RECT 59.635 111.240 59.955 111.300 ;
        RECT 62.070 111.240 62.720 111.285 ;
        RECT 58.830 111.100 62.720 111.240 ;
        RECT 58.830 111.055 59.420 111.100 ;
        RECT 49.070 110.900 49.360 110.945 ;
        RECT 40.315 110.760 49.360 110.900 ;
        RECT 40.315 110.700 40.635 110.760 ;
        RECT 49.070 110.715 49.360 110.760 ;
        RECT 50.450 110.715 50.740 110.945 ;
        RECT 51.815 110.700 52.135 110.960 ;
        RECT 55.510 110.900 55.800 110.945 ;
        RECT 57.335 110.900 57.655 110.960 ;
        RECT 55.510 110.760 57.655 110.900 ;
        RECT 55.510 110.715 55.800 110.760 ;
        RECT 57.335 110.700 57.655 110.760 ;
        RECT 59.130 110.740 59.420 111.055 ;
        RECT 59.635 111.040 59.955 111.100 ;
        RECT 62.070 111.055 62.720 111.100 ;
        RECT 66.165 110.945 66.305 111.440 ;
        RECT 66.535 111.440 83.325 111.580 ;
        RECT 66.535 111.380 66.855 111.440 ;
        RECT 74.815 111.240 75.135 111.300 ;
        RECT 74.815 111.100 77.345 111.240 ;
        RECT 74.815 111.040 75.135 111.100 ;
        RECT 60.210 110.900 60.500 110.945 ;
        RECT 63.790 110.900 64.080 110.945 ;
        RECT 65.625 110.900 65.915 110.945 ;
        RECT 60.210 110.760 65.915 110.900 ;
        RECT 60.210 110.715 60.500 110.760 ;
        RECT 63.790 110.715 64.080 110.760 ;
        RECT 65.625 110.715 65.915 110.760 ;
        RECT 66.090 110.715 66.380 110.945 ;
        RECT 71.135 110.900 71.455 110.960 ;
        RECT 72.990 110.900 73.280 110.945 ;
        RECT 71.135 110.760 73.280 110.900 ;
        RECT 71.135 110.700 71.455 110.760 ;
        RECT 72.990 110.715 73.280 110.760 ;
        RECT 73.910 110.900 74.200 110.945 ;
        RECT 74.355 110.900 74.675 110.960 ;
        RECT 77.205 110.945 77.345 111.100 ;
        RECT 83.185 110.945 83.325 111.440 ;
        RECT 92.295 111.380 92.615 111.640 ;
        RECT 94.610 111.580 94.900 111.625 ;
        RECT 96.895 111.580 97.215 111.640 ;
        RECT 94.610 111.440 97.215 111.580 ;
        RECT 94.610 111.395 94.900 111.440 ;
        RECT 96.895 111.380 97.215 111.440 ;
        RECT 109.775 111.380 110.095 111.640 ;
        RECT 83.555 111.240 83.875 111.300 ;
        RECT 92.770 111.240 93.060 111.285 ;
        RECT 83.555 111.100 93.060 111.240 ;
        RECT 83.555 111.040 83.875 111.100 ;
        RECT 92.770 111.055 93.060 111.100 ;
        RECT 93.305 111.100 106.325 111.240 ;
        RECT 73.910 110.760 74.675 110.900 ;
        RECT 73.910 110.715 74.200 110.760 ;
        RECT 74.355 110.700 74.675 110.760 ;
        RECT 75.750 110.715 76.040 110.945 ;
        RECT 77.130 110.715 77.420 110.945 ;
        RECT 83.110 110.715 83.400 110.945 ;
        RECT 87.695 110.900 88.015 110.960 ;
        RECT 89.550 110.900 89.840 110.945 ;
        RECT 87.695 110.760 89.840 110.900 ;
        RECT 26.055 110.360 26.375 110.620 ;
        RECT 28.830 110.560 29.120 110.605 ;
        RECT 31.115 110.560 31.435 110.620 ;
        RECT 28.830 110.420 31.435 110.560 ;
        RECT 28.830 110.375 29.120 110.420 ;
        RECT 31.115 110.360 31.435 110.420 ;
        RECT 37.095 110.560 37.415 110.620 ;
        RECT 38.950 110.560 39.240 110.605 ;
        RECT 37.095 110.420 39.240 110.560 ;
        RECT 37.095 110.360 37.415 110.420 ;
        RECT 38.950 110.375 39.240 110.420 ;
        RECT 55.970 110.560 56.260 110.605 ;
        RECT 58.255 110.560 58.575 110.620 ;
        RECT 55.970 110.420 58.575 110.560 ;
        RECT 55.970 110.375 56.260 110.420 ;
        RECT 58.255 110.360 58.575 110.420 ;
        RECT 64.235 110.560 64.555 110.620 ;
        RECT 64.710 110.560 65.000 110.605 ;
        RECT 64.235 110.420 65.000 110.560 ;
        RECT 64.235 110.360 64.555 110.420 ;
        RECT 64.710 110.375 65.000 110.420 ;
        RECT 72.070 110.560 72.360 110.605 ;
        RECT 75.825 110.560 75.965 110.715 ;
        RECT 87.695 110.700 88.015 110.760 ;
        RECT 89.550 110.715 89.840 110.760 ;
        RECT 91.835 110.900 92.155 110.960 ;
        RECT 93.305 110.900 93.445 111.100 ;
        RECT 91.835 110.760 93.445 110.900 ;
        RECT 94.595 110.900 94.915 110.960 ;
        RECT 98.290 110.900 98.580 110.945 ;
        RECT 94.595 110.760 98.580 110.900 ;
        RECT 91.835 110.700 92.155 110.760 ;
        RECT 94.595 110.700 94.915 110.760 ;
        RECT 98.290 110.715 98.580 110.760 ;
        RECT 101.035 110.700 101.355 110.960 ;
        RECT 106.185 110.945 106.325 111.100 ;
        RECT 102.430 110.900 102.720 110.945 ;
        RECT 103.810 110.900 104.100 110.945 ;
        RECT 102.430 110.760 104.100 110.900 ;
        RECT 102.430 110.715 102.720 110.760 ;
        RECT 103.810 110.715 104.100 110.760 ;
        RECT 106.110 110.715 106.400 110.945 ;
        RECT 78.035 110.560 78.355 110.620 ;
        RECT 72.070 110.420 78.355 110.560 ;
        RECT 72.070 110.375 72.360 110.420 ;
        RECT 78.035 110.360 78.355 110.420 ;
        RECT 87.235 110.560 87.555 110.620 ;
        RECT 91.390 110.560 91.680 110.605 ;
        RECT 102.505 110.560 102.645 110.715 ;
        RECT 106.555 110.700 106.875 110.960 ;
        RECT 110.695 110.700 111.015 110.960 ;
        RECT 87.235 110.420 91.680 110.560 ;
        RECT 87.235 110.360 87.555 110.420 ;
        RECT 91.390 110.375 91.680 110.420 ;
        RECT 101.355 110.420 102.645 110.560 ;
        RECT 33.070 110.220 33.360 110.265 ;
        RECT 36.190 110.220 36.480 110.265 ;
        RECT 38.080 110.220 38.370 110.265 ;
        RECT 33.070 110.080 38.370 110.220 ;
        RECT 33.070 110.035 33.360 110.080 ;
        RECT 36.190 110.035 36.480 110.080 ;
        RECT 38.080 110.035 38.370 110.080 ;
        RECT 60.210 110.220 60.500 110.265 ;
        RECT 63.330 110.220 63.620 110.265 ;
        RECT 65.220 110.220 65.510 110.265 ;
        RECT 60.210 110.080 65.510 110.220 ;
        RECT 60.210 110.035 60.500 110.080 ;
        RECT 63.330 110.035 63.620 110.080 ;
        RECT 65.220 110.035 65.510 110.080 ;
        RECT 98.275 110.220 98.595 110.280 ;
        RECT 101.355 110.220 101.495 110.420 ;
        RECT 98.275 110.080 101.495 110.220 ;
        RECT 101.970 110.220 102.260 110.265 ;
        RECT 108.395 110.220 108.715 110.280 ;
        RECT 101.970 110.080 108.715 110.220 ;
        RECT 98.275 110.020 98.595 110.080 ;
        RECT 101.970 110.035 102.260 110.080 ;
        RECT 108.395 110.020 108.715 110.080 ;
        RECT 21.470 109.880 21.760 109.925 ;
        RECT 27.435 109.880 27.755 109.940 ;
        RECT 21.470 109.740 27.755 109.880 ;
        RECT 21.470 109.695 21.760 109.740 ;
        RECT 27.435 109.680 27.755 109.740 ;
        RECT 37.665 109.880 37.955 109.925 ;
        RECT 40.775 109.880 41.095 109.940 ;
        RECT 37.665 109.740 41.095 109.880 ;
        RECT 37.665 109.695 37.955 109.740 ;
        RECT 40.775 109.680 41.095 109.740 ;
        RECT 49.990 109.880 50.280 109.925 ;
        RECT 55.495 109.880 55.815 109.940 ;
        RECT 49.990 109.740 55.815 109.880 ;
        RECT 49.990 109.695 50.280 109.740 ;
        RECT 55.495 109.680 55.815 109.740 ;
        RECT 74.815 109.680 75.135 109.940 ;
        RECT 75.735 109.880 76.055 109.940 ;
        RECT 76.210 109.880 76.500 109.925 ;
        RECT 75.735 109.740 76.500 109.880 ;
        RECT 75.735 109.680 76.055 109.740 ;
        RECT 76.210 109.695 76.500 109.740 ;
        RECT 78.050 109.880 78.340 109.925 ;
        RECT 80.335 109.880 80.655 109.940 ;
        RECT 78.050 109.740 80.655 109.880 ;
        RECT 78.050 109.695 78.340 109.740 ;
        RECT 80.335 109.680 80.655 109.740 ;
        RECT 84.015 109.680 84.335 109.940 ;
        RECT 90.470 109.880 90.760 109.925 ;
        RECT 93.215 109.880 93.535 109.940 ;
        RECT 90.470 109.740 93.535 109.880 ;
        RECT 90.470 109.695 90.760 109.740 ;
        RECT 93.215 109.680 93.535 109.740 ;
        RECT 97.355 109.680 97.675 109.940 ;
        RECT 102.890 109.880 103.180 109.925 ;
        RECT 103.335 109.880 103.655 109.940 ;
        RECT 102.890 109.740 103.655 109.880 ;
        RECT 102.890 109.695 103.180 109.740 ;
        RECT 103.335 109.680 103.655 109.740 ;
        RECT 104.255 109.680 104.575 109.940 ;
        RECT 105.175 109.680 105.495 109.940 ;
        RECT 107.475 109.680 107.795 109.940 ;
        RECT 18.165 109.060 112.465 109.540 ;
        RECT 40.775 108.660 41.095 108.920 ;
        RECT 63.330 108.860 63.620 108.905 ;
        RECT 64.235 108.860 64.555 108.920 ;
        RECT 63.330 108.720 64.555 108.860 ;
        RECT 63.330 108.675 63.620 108.720 ;
        RECT 64.235 108.660 64.555 108.720 ;
        RECT 73.895 108.860 74.215 108.920 ;
        RECT 95.515 108.860 95.835 108.920 ;
        RECT 73.895 108.720 86.085 108.860 ;
        RECT 73.895 108.660 74.215 108.720 ;
        RECT 27.550 108.520 27.840 108.565 ;
        RECT 30.670 108.520 30.960 108.565 ;
        RECT 32.560 108.520 32.850 108.565 ;
        RECT 27.550 108.380 32.850 108.520 ;
        RECT 27.550 108.335 27.840 108.380 ;
        RECT 30.670 108.335 30.960 108.380 ;
        RECT 32.560 108.335 32.850 108.380 ;
        RECT 35.730 108.335 36.020 108.565 ;
        RECT 38.475 108.520 38.795 108.580 ;
        RECT 44.010 108.520 44.300 108.565 ;
        RECT 38.475 108.380 44.300 108.520 ;
        RECT 23.310 108.180 23.600 108.225 ;
        RECT 26.055 108.180 26.375 108.240 ;
        RECT 23.310 108.040 26.375 108.180 ;
        RECT 23.310 107.995 23.600 108.040 ;
        RECT 26.055 107.980 26.375 108.040 ;
        RECT 32.050 108.180 32.340 108.225 ;
        RECT 35.805 108.180 35.945 108.335 ;
        RECT 38.475 108.320 38.795 108.380 ;
        RECT 44.010 108.335 44.300 108.380 ;
        RECT 49.975 108.320 50.295 108.580 ;
        RECT 51.010 108.520 51.300 108.565 ;
        RECT 54.130 108.520 54.420 108.565 ;
        RECT 56.020 108.520 56.310 108.565 ;
        RECT 60.095 108.520 60.415 108.580 ;
        RECT 51.010 108.380 56.310 108.520 ;
        RECT 51.010 108.335 51.300 108.380 ;
        RECT 54.130 108.335 54.420 108.380 ;
        RECT 56.020 108.335 56.310 108.380 ;
        RECT 56.965 108.380 60.415 108.520 ;
        RECT 50.065 108.180 50.205 108.320 ;
        RECT 32.050 108.040 35.945 108.180 ;
        RECT 41.785 108.040 50.205 108.180 ;
        RECT 32.050 107.995 32.340 108.040 ;
        RECT 24.215 107.500 24.535 107.560 ;
        RECT 26.470 107.545 26.760 107.860 ;
        RECT 27.550 107.840 27.840 107.885 ;
        RECT 31.130 107.840 31.420 107.885 ;
        RECT 32.965 107.840 33.255 107.885 ;
        RECT 27.550 107.700 33.255 107.840 ;
        RECT 27.550 107.655 27.840 107.700 ;
        RECT 31.130 107.655 31.420 107.700 ;
        RECT 32.965 107.655 33.255 107.700 ;
        RECT 33.415 107.640 33.735 107.900 ;
        RECT 36.650 107.840 36.940 107.885 ;
        RECT 38.015 107.840 38.335 107.900 ;
        RECT 36.650 107.700 38.335 107.840 ;
        RECT 36.650 107.655 36.940 107.700 ;
        RECT 38.015 107.640 38.335 107.700 ;
        RECT 38.490 107.840 38.780 107.885 ;
        RECT 39.395 107.840 39.715 107.900 ;
        RECT 41.785 107.885 41.925 108.040 ;
        RECT 55.495 107.980 55.815 108.240 ;
        RECT 56.965 108.225 57.105 108.380 ;
        RECT 60.095 108.320 60.415 108.380 ;
        RECT 69.410 108.520 69.700 108.565 ;
        RECT 72.530 108.520 72.820 108.565 ;
        RECT 74.420 108.520 74.710 108.565 ;
        RECT 69.410 108.380 74.710 108.520 ;
        RECT 69.410 108.335 69.700 108.380 ;
        RECT 72.530 108.335 72.820 108.380 ;
        RECT 74.420 108.335 74.710 108.380 ;
        RECT 75.365 108.225 75.505 108.720 ;
        RECT 79.990 108.520 80.280 108.565 ;
        RECT 83.110 108.520 83.400 108.565 ;
        RECT 85.000 108.520 85.290 108.565 ;
        RECT 79.990 108.380 85.290 108.520 ;
        RECT 79.990 108.335 80.280 108.380 ;
        RECT 83.110 108.335 83.400 108.380 ;
        RECT 85.000 108.335 85.290 108.380 ;
        RECT 56.890 107.995 57.180 108.225 ;
        RECT 75.290 107.995 75.580 108.225 ;
        RECT 75.750 108.180 76.040 108.225 ;
        RECT 81.255 108.180 81.575 108.240 ;
        RECT 75.750 108.040 81.575 108.180 ;
        RECT 75.750 107.995 76.040 108.040 ;
        RECT 81.255 107.980 81.575 108.040 ;
        RECT 84.015 108.180 84.335 108.240 ;
        RECT 85.945 108.225 86.085 108.720 ;
        RECT 95.515 108.720 99.425 108.860 ;
        RECT 95.515 108.660 95.835 108.720 ;
        RECT 91.950 108.520 92.240 108.565 ;
        RECT 95.070 108.520 95.360 108.565 ;
        RECT 96.960 108.520 97.250 108.565 ;
        RECT 98.290 108.520 98.580 108.565 ;
        RECT 91.950 108.380 97.250 108.520 ;
        RECT 91.950 108.335 92.240 108.380 ;
        RECT 95.070 108.335 95.360 108.380 ;
        RECT 96.960 108.335 97.250 108.380 ;
        RECT 97.445 108.380 98.580 108.520 ;
        RECT 84.490 108.180 84.780 108.225 ;
        RECT 84.015 108.040 84.780 108.180 ;
        RECT 84.015 107.980 84.335 108.040 ;
        RECT 84.490 107.995 84.780 108.040 ;
        RECT 85.870 107.995 86.160 108.225 ;
        RECT 87.710 108.180 88.000 108.225 ;
        RECT 90.455 108.180 90.775 108.240 ;
        RECT 87.710 108.040 90.775 108.180 ;
        RECT 87.710 107.995 88.000 108.040 ;
        RECT 90.455 107.980 90.775 108.040 ;
        RECT 96.450 108.180 96.740 108.225 ;
        RECT 97.445 108.180 97.585 108.380 ;
        RECT 98.290 108.335 98.580 108.380 ;
        RECT 96.450 108.040 97.585 108.180 ;
        RECT 96.450 107.995 96.740 108.040 ;
        RECT 97.815 107.980 98.135 108.240 ;
        RECT 38.490 107.700 39.715 107.840 ;
        RECT 38.490 107.655 38.780 107.700 ;
        RECT 39.395 107.640 39.715 107.700 ;
        RECT 41.710 107.655 42.000 107.885 ;
        RECT 42.615 107.840 42.935 107.900 ;
        RECT 43.550 107.840 43.840 107.885 ;
        RECT 42.615 107.700 43.840 107.840 ;
        RECT 42.615 107.640 42.935 107.700 ;
        RECT 43.550 107.655 43.840 107.700 ;
        RECT 44.915 107.640 45.235 107.900 ;
        RECT 45.375 107.640 45.695 107.900 ;
        RECT 49.975 107.860 50.295 107.900 ;
        RECT 49.930 107.640 50.295 107.860 ;
        RECT 51.010 107.840 51.300 107.885 ;
        RECT 54.590 107.840 54.880 107.885 ;
        RECT 56.425 107.840 56.715 107.885 ;
        RECT 51.010 107.700 56.715 107.840 ;
        RECT 51.010 107.655 51.300 107.700 ;
        RECT 54.590 107.655 54.880 107.700 ;
        RECT 56.425 107.655 56.715 107.700 ;
        RECT 57.335 107.840 57.655 107.900 ;
        RECT 57.810 107.840 58.100 107.885 ;
        RECT 57.335 107.700 58.100 107.840 ;
        RECT 57.335 107.640 57.655 107.700 ;
        RECT 57.810 107.655 58.100 107.700 ;
        RECT 59.175 107.840 59.495 107.900 ;
        RECT 61.030 107.840 61.320 107.885 ;
        RECT 59.175 107.700 61.320 107.840 ;
        RECT 59.175 107.640 59.495 107.700 ;
        RECT 61.030 107.655 61.320 107.700 ;
        RECT 61.475 107.840 61.795 107.900 ;
        RECT 62.410 107.840 62.700 107.885 ;
        RECT 61.475 107.700 62.700 107.840 ;
        RECT 61.475 107.640 61.795 107.700 ;
        RECT 62.410 107.655 62.700 107.700 ;
        RECT 63.775 107.640 64.095 107.900 ;
        RECT 99.285 107.885 99.425 108.720 ;
        RECT 104.830 108.520 105.120 108.565 ;
        RECT 107.950 108.520 108.240 108.565 ;
        RECT 109.840 108.520 110.130 108.565 ;
        RECT 104.830 108.380 110.130 108.520 ;
        RECT 104.830 108.335 105.120 108.380 ;
        RECT 107.950 108.335 108.240 108.380 ;
        RECT 109.840 108.335 110.130 108.380 ;
        RECT 107.475 108.180 107.795 108.240 ;
        RECT 109.330 108.180 109.620 108.225 ;
        RECT 107.475 108.040 109.620 108.180 ;
        RECT 107.475 107.980 107.795 108.040 ;
        RECT 109.330 107.995 109.620 108.040 ;
        RECT 26.170 107.500 26.760 107.545 ;
        RECT 29.410 107.500 30.060 107.545 ;
        RECT 46.770 107.500 47.060 107.545 ;
        RECT 49.055 107.500 49.375 107.560 ;
        RECT 49.930 107.545 50.220 107.640 ;
        RECT 24.215 107.360 30.060 107.500 ;
        RECT 24.215 107.300 24.535 107.360 ;
        RECT 26.170 107.315 26.460 107.360 ;
        RECT 29.410 107.315 30.060 107.360 ;
        RECT 35.345 107.360 42.845 107.500 ;
        RECT 27.895 107.160 28.215 107.220 ;
        RECT 35.345 107.160 35.485 107.360 ;
        RECT 27.895 107.020 35.485 107.160 ;
        RECT 27.895 106.960 28.215 107.020 ;
        RECT 38.015 106.960 38.335 107.220 ;
        RECT 39.870 107.160 40.160 107.205 ;
        RECT 40.315 107.160 40.635 107.220 ;
        RECT 42.705 107.205 42.845 107.360 ;
        RECT 46.770 107.360 49.375 107.500 ;
        RECT 46.770 107.315 47.060 107.360 ;
        RECT 49.055 107.300 49.375 107.360 ;
        RECT 49.630 107.500 50.220 107.545 ;
        RECT 52.870 107.500 53.520 107.545 ;
        RECT 49.630 107.360 53.520 107.500 ;
        RECT 49.630 107.315 49.920 107.360 ;
        RECT 52.870 107.315 53.520 107.360 ;
        RECT 65.170 107.500 65.460 107.545 ;
        RECT 67.455 107.500 67.775 107.560 ;
        RECT 68.330 107.545 68.620 107.860 ;
        RECT 69.410 107.840 69.700 107.885 ;
        RECT 72.990 107.840 73.280 107.885 ;
        RECT 74.825 107.840 75.115 107.885 ;
        RECT 69.410 107.700 75.115 107.840 ;
        RECT 69.410 107.655 69.700 107.700 ;
        RECT 72.990 107.655 73.280 107.700 ;
        RECT 74.825 107.655 75.115 107.700 ;
        RECT 65.170 107.360 67.775 107.500 ;
        RECT 65.170 107.315 65.460 107.360 ;
        RECT 67.455 107.300 67.775 107.360 ;
        RECT 68.030 107.500 68.620 107.545 ;
        RECT 71.135 107.545 71.455 107.560 ;
        RECT 71.135 107.500 71.920 107.545 ;
        RECT 68.030 107.360 71.920 107.500 ;
        RECT 68.030 107.315 68.320 107.360 ;
        RECT 71.135 107.315 71.920 107.360 ;
        RECT 73.435 107.500 73.755 107.560 ;
        RECT 78.910 107.545 79.200 107.860 ;
        RECT 79.990 107.840 80.280 107.885 ;
        RECT 83.570 107.840 83.860 107.885 ;
        RECT 85.405 107.840 85.695 107.885 ;
        RECT 79.990 107.700 85.695 107.840 ;
        RECT 79.990 107.655 80.280 107.700 ;
        RECT 83.570 107.655 83.860 107.700 ;
        RECT 85.405 107.655 85.695 107.700 ;
        RECT 73.910 107.500 74.200 107.545 ;
        RECT 73.435 107.360 74.200 107.500 ;
        RECT 71.135 107.300 71.455 107.315 ;
        RECT 73.435 107.300 73.755 107.360 ;
        RECT 73.910 107.315 74.200 107.360 ;
        RECT 78.610 107.500 79.200 107.545 ;
        RECT 79.415 107.500 79.735 107.560 ;
        RECT 90.870 107.545 91.160 107.860 ;
        RECT 91.950 107.840 92.240 107.885 ;
        RECT 95.530 107.840 95.820 107.885 ;
        RECT 97.365 107.840 97.655 107.885 ;
        RECT 91.950 107.700 97.655 107.840 ;
        RECT 91.950 107.655 92.240 107.700 ;
        RECT 95.530 107.655 95.820 107.700 ;
        RECT 97.365 107.655 97.655 107.700 ;
        RECT 99.210 107.655 99.500 107.885 ;
        RECT 94.135 107.545 94.455 107.560 ;
        RECT 81.850 107.500 82.500 107.545 ;
        RECT 78.610 107.360 82.500 107.500 ;
        RECT 78.610 107.315 78.900 107.360 ;
        RECT 79.415 107.300 79.735 107.360 ;
        RECT 81.850 107.315 82.500 107.360 ;
        RECT 90.570 107.500 91.160 107.545 ;
        RECT 93.810 107.500 94.460 107.545 ;
        RECT 90.570 107.360 94.460 107.500 ;
        RECT 90.570 107.315 90.860 107.360 ;
        RECT 93.810 107.315 94.460 107.360 ;
        RECT 100.590 107.500 100.880 107.545 ;
        RECT 102.875 107.500 103.195 107.560 ;
        RECT 103.750 107.545 104.040 107.860 ;
        RECT 104.830 107.840 105.120 107.885 ;
        RECT 108.410 107.840 108.700 107.885 ;
        RECT 110.245 107.840 110.535 107.885 ;
        RECT 104.830 107.700 110.535 107.840 ;
        RECT 104.830 107.655 105.120 107.700 ;
        RECT 108.410 107.655 108.700 107.700 ;
        RECT 110.245 107.655 110.535 107.700 ;
        RECT 110.710 107.655 111.000 107.885 ;
        RECT 100.590 107.360 103.195 107.500 ;
        RECT 100.590 107.315 100.880 107.360 ;
        RECT 94.135 107.300 94.455 107.315 ;
        RECT 102.875 107.300 103.195 107.360 ;
        RECT 103.450 107.500 104.040 107.545 ;
        RECT 104.255 107.500 104.575 107.560 ;
        RECT 106.690 107.500 107.340 107.545 ;
        RECT 110.785 107.500 110.925 107.655 ;
        RECT 103.450 107.360 107.340 107.500 ;
        RECT 103.450 107.315 103.740 107.360 ;
        RECT 104.255 107.300 104.575 107.360 ;
        RECT 106.690 107.315 107.340 107.360 ;
        RECT 109.865 107.360 110.925 107.500 ;
        RECT 109.865 107.220 110.005 107.360 ;
        RECT 39.870 107.020 40.635 107.160 ;
        RECT 39.870 106.975 40.160 107.020 ;
        RECT 40.315 106.960 40.635 107.020 ;
        RECT 42.630 106.975 42.920 107.205 ;
        RECT 45.835 107.160 46.155 107.220 ;
        RECT 46.310 107.160 46.600 107.205 ;
        RECT 45.835 107.020 46.600 107.160 ;
        RECT 45.835 106.960 46.155 107.020 ;
        RECT 46.310 106.975 46.600 107.020 ;
        RECT 61.475 106.960 61.795 107.220 ;
        RECT 64.710 107.160 65.000 107.205 ;
        RECT 70.215 107.160 70.535 107.220 ;
        RECT 64.710 107.020 70.535 107.160 ;
        RECT 64.710 106.975 65.000 107.020 ;
        RECT 70.215 106.960 70.535 107.020 ;
        RECT 97.815 107.160 98.135 107.220 ;
        RECT 109.775 107.160 110.095 107.220 ;
        RECT 97.815 107.020 110.095 107.160 ;
        RECT 97.815 106.960 98.135 107.020 ;
        RECT 109.775 106.960 110.095 107.020 ;
        RECT 17.370 106.340 112.465 106.820 ;
        RECT 135.660 106.690 136.800 133.400 ;
        RECT 133.100 106.600 136.850 106.690 ;
        RECT 24.215 105.940 24.535 106.200 ;
        RECT 25.610 106.140 25.900 106.185 ;
        RECT 28.815 106.140 29.135 106.200 ;
        RECT 25.610 106.000 29.135 106.140 ;
        RECT 25.610 105.955 25.900 106.000 ;
        RECT 28.815 105.940 29.135 106.000 ;
        RECT 39.395 106.140 39.715 106.200 ;
        RECT 39.395 106.000 49.285 106.140 ;
        RECT 39.395 105.940 39.715 106.000 ;
        RECT 27.895 105.600 28.215 105.860 ;
        RECT 30.190 105.800 30.840 105.845 ;
        RECT 33.790 105.800 34.080 105.845 ;
        RECT 38.015 105.800 38.335 105.860 ;
        RECT 30.190 105.660 38.335 105.800 ;
        RECT 30.190 105.615 30.840 105.660 ;
        RECT 33.490 105.615 34.080 105.660 ;
        RECT 23.310 105.460 23.600 105.505 ;
        RECT 23.770 105.460 24.060 105.505 ;
        RECT 25.150 105.460 25.440 105.505 ;
        RECT 23.310 105.320 25.440 105.460 ;
        RECT 23.310 105.275 23.600 105.320 ;
        RECT 23.770 105.275 24.060 105.320 ;
        RECT 25.150 105.275 25.440 105.320 ;
        RECT 26.995 105.460 27.285 105.505 ;
        RECT 28.830 105.460 29.120 105.505 ;
        RECT 32.410 105.460 32.700 105.505 ;
        RECT 26.995 105.320 32.700 105.460 ;
        RECT 26.995 105.275 27.285 105.320 ;
        RECT 28.830 105.275 29.120 105.320 ;
        RECT 32.410 105.275 32.700 105.320 ;
        RECT 33.490 105.300 33.780 105.615 ;
        RECT 38.015 105.600 38.335 105.660 ;
        RECT 38.475 105.600 38.795 105.860 ;
        RECT 40.770 105.800 41.420 105.845 ;
        RECT 44.370 105.800 44.660 105.845 ;
        RECT 40.770 105.660 44.660 105.800 ;
        RECT 40.770 105.615 41.420 105.660 ;
        RECT 44.070 105.615 44.660 105.660 ;
        RECT 37.575 105.460 37.865 105.505 ;
        RECT 39.410 105.460 39.700 105.505 ;
        RECT 42.990 105.460 43.280 105.505 ;
        RECT 37.575 105.320 43.280 105.460 ;
        RECT 37.575 105.275 37.865 105.320 ;
        RECT 39.410 105.275 39.700 105.320 ;
        RECT 42.990 105.275 43.280 105.320 ;
        RECT 44.070 105.460 44.360 105.615 ;
        RECT 49.145 105.505 49.285 106.000 ;
        RECT 49.975 105.940 50.295 106.200 ;
        RECT 72.055 105.940 72.375 106.200 ;
        RECT 72.990 106.140 73.280 106.185 ;
        RECT 73.435 106.140 73.755 106.200 ;
        RECT 72.990 106.000 73.755 106.140 ;
        RECT 72.990 105.955 73.280 106.000 ;
        RECT 73.435 105.940 73.755 106.000 ;
        RECT 74.815 106.140 75.135 106.200 ;
        RECT 94.135 106.140 94.455 106.200 ;
        RECT 95.530 106.140 95.820 106.185 ;
        RECT 74.815 106.000 82.865 106.140 ;
        RECT 74.815 105.940 75.135 106.000 ;
        RECT 53.770 105.800 54.060 105.845 ;
        RECT 55.955 105.800 56.275 105.860 ;
        RECT 57.010 105.800 57.660 105.845 ;
        RECT 53.770 105.660 57.660 105.800 ;
        RECT 53.770 105.615 54.360 105.660 ;
        RECT 48.610 105.460 48.900 105.505 ;
        RECT 44.070 105.320 48.900 105.460 ;
        RECT 44.070 105.300 44.360 105.320 ;
        RECT 48.610 105.275 48.900 105.320 ;
        RECT 49.070 105.460 49.360 105.505 ;
        RECT 49.530 105.460 49.820 105.505 ;
        RECT 49.070 105.320 49.820 105.460 ;
        RECT 49.070 105.275 49.360 105.320 ;
        RECT 49.530 105.275 49.820 105.320 ;
        RECT 54.070 105.300 54.360 105.615 ;
        RECT 55.955 105.600 56.275 105.660 ;
        RECT 57.010 105.615 57.660 105.660 ;
        RECT 60.095 105.800 60.415 105.860 ;
        RECT 61.475 105.800 61.795 105.860 ;
        RECT 64.350 105.800 64.640 105.845 ;
        RECT 67.590 105.800 68.240 105.845 ;
        RECT 60.095 105.660 61.245 105.800 ;
        RECT 60.095 105.600 60.415 105.660 ;
        RECT 61.105 105.505 61.245 105.660 ;
        RECT 61.475 105.660 68.240 105.800 ;
        RECT 61.475 105.600 61.795 105.660 ;
        RECT 64.350 105.615 64.940 105.660 ;
        RECT 67.590 105.615 68.240 105.660 ;
        RECT 55.150 105.460 55.440 105.505 ;
        RECT 58.730 105.460 59.020 105.505 ;
        RECT 60.565 105.460 60.855 105.505 ;
        RECT 55.150 105.320 60.855 105.460 ;
        RECT 55.150 105.275 55.440 105.320 ;
        RECT 58.730 105.275 59.020 105.320 ;
        RECT 60.565 105.275 60.855 105.320 ;
        RECT 61.030 105.275 61.320 105.505 ;
        RECT 64.650 105.300 64.940 105.615 ;
        RECT 70.215 105.600 70.535 105.860 ;
        RECT 71.595 105.600 71.915 105.860 ;
        RECT 72.145 105.800 72.285 105.940 ;
        RECT 82.725 105.845 82.865 106.000 ;
        RECT 94.135 106.000 95.820 106.140 ;
        RECT 94.135 105.940 94.455 106.000 ;
        RECT 95.530 105.955 95.820 106.000 ;
        RECT 97.815 105.940 98.135 106.200 ;
        RECT 73.910 105.800 74.200 105.845 ;
        RECT 72.145 105.660 74.200 105.800 ;
        RECT 73.910 105.615 74.200 105.660 ;
        RECT 76.770 105.800 77.060 105.845 ;
        RECT 80.010 105.800 80.660 105.845 ;
        RECT 76.770 105.660 80.660 105.800 ;
        RECT 76.770 105.615 77.360 105.660 ;
        RECT 80.010 105.615 80.660 105.660 ;
        RECT 82.650 105.615 82.940 105.845 ;
        RECT 87.350 105.800 87.640 105.845 ;
        RECT 90.590 105.800 91.240 105.845 ;
        RECT 87.350 105.660 91.240 105.800 ;
        RECT 87.350 105.615 87.940 105.660 ;
        RECT 90.590 105.615 91.240 105.660 ;
        RECT 65.730 105.460 66.020 105.505 ;
        RECT 69.310 105.460 69.600 105.505 ;
        RECT 71.145 105.460 71.435 105.505 ;
        RECT 65.730 105.320 71.435 105.460 ;
        RECT 71.685 105.460 71.825 105.600 ;
        RECT 72.070 105.460 72.360 105.505 ;
        RECT 71.685 105.320 72.360 105.460 ;
        RECT 65.730 105.275 66.020 105.320 ;
        RECT 69.310 105.275 69.600 105.320 ;
        RECT 71.145 105.275 71.435 105.320 ;
        RECT 72.070 105.275 72.360 105.320 ;
        RECT 72.515 105.460 72.835 105.520 ;
        RECT 77.070 105.460 77.360 105.615 ;
        RECT 87.650 105.520 87.940 105.615 ;
        RECT 93.215 105.600 93.535 105.860 ;
        RECT 97.905 105.800 98.045 105.940 ;
        RECT 98.735 105.800 99.055 105.860 ;
        RECT 94.685 105.660 99.055 105.800 ;
        RECT 72.515 105.320 77.360 105.460 ;
        RECT 22.835 104.240 23.155 104.500 ;
        RECT 25.225 104.440 25.365 105.275 ;
        RECT 26.530 105.120 26.820 105.165 ;
        RECT 32.955 105.120 33.275 105.180 ;
        RECT 26.530 104.980 33.275 105.120 ;
        RECT 26.530 104.935 26.820 104.980 ;
        RECT 32.955 104.920 33.275 104.980 ;
        RECT 35.255 105.120 35.575 105.180 ;
        RECT 36.650 105.120 36.940 105.165 ;
        RECT 35.255 104.980 36.940 105.120 ;
        RECT 35.255 104.920 35.575 104.980 ;
        RECT 36.650 104.935 36.940 104.980 ;
        RECT 37.095 104.920 37.415 105.180 ;
        RECT 44.455 105.120 44.775 105.180 ;
        RECT 47.230 105.120 47.520 105.165 ;
        RECT 44.455 104.980 47.520 105.120 ;
        RECT 44.455 104.920 44.775 104.980 ;
        RECT 47.230 104.935 47.520 104.980 ;
        RECT 27.400 104.780 27.690 104.825 ;
        RECT 29.290 104.780 29.580 104.825 ;
        RECT 32.410 104.780 32.700 104.825 ;
        RECT 27.400 104.640 32.700 104.780 ;
        RECT 27.400 104.595 27.690 104.640 ;
        RECT 29.290 104.595 29.580 104.640 ;
        RECT 32.410 104.595 32.700 104.640 ;
        RECT 37.980 104.780 38.270 104.825 ;
        RECT 39.870 104.780 40.160 104.825 ;
        RECT 42.990 104.780 43.280 104.825 ;
        RECT 37.980 104.640 43.280 104.780 ;
        RECT 49.605 104.780 49.745 105.275 ;
        RECT 72.515 105.260 72.835 105.320 ;
        RECT 77.070 105.300 77.360 105.320 ;
        RECT 78.150 105.460 78.440 105.505 ;
        RECT 81.730 105.460 82.020 105.505 ;
        RECT 83.565 105.460 83.855 105.505 ;
        RECT 78.150 105.320 83.855 105.460 ;
        RECT 78.150 105.275 78.440 105.320 ;
        RECT 81.730 105.275 82.020 105.320 ;
        RECT 83.565 105.275 83.855 105.320 ;
        RECT 87.650 105.300 88.015 105.520 ;
        RECT 94.685 105.505 94.825 105.660 ;
        RECT 98.735 105.600 99.055 105.660 ;
        RECT 102.530 105.800 102.820 105.845 ;
        RECT 105.770 105.800 106.420 105.845 ;
        RECT 102.530 105.660 106.420 105.800 ;
        RECT 102.530 105.615 103.120 105.660 ;
        RECT 105.770 105.615 106.420 105.660 ;
        RECT 87.695 105.260 88.015 105.300 ;
        RECT 88.730 105.460 89.020 105.505 ;
        RECT 92.310 105.460 92.600 105.505 ;
        RECT 94.145 105.460 94.435 105.505 ;
        RECT 88.730 105.320 94.435 105.460 ;
        RECT 88.730 105.275 89.020 105.320 ;
        RECT 92.310 105.275 92.600 105.320 ;
        RECT 94.145 105.275 94.435 105.320 ;
        RECT 94.610 105.275 94.900 105.505 ;
        RECT 95.055 105.460 95.375 105.520 ;
        RECT 95.990 105.460 96.280 105.505 ;
        RECT 97.370 105.460 97.660 105.505 ;
        RECT 97.815 105.460 98.135 105.520 ;
        RECT 95.055 105.320 98.135 105.460 ;
        RECT 95.055 105.260 95.375 105.320 ;
        RECT 95.990 105.275 96.280 105.320 ;
        RECT 97.370 105.275 97.660 105.320 ;
        RECT 97.815 105.260 98.135 105.320 ;
        RECT 98.290 105.460 98.580 105.505 ;
        RECT 102.830 105.460 103.120 105.615 ;
        RECT 108.395 105.600 108.715 105.860 ;
        RECT 129.700 105.630 136.850 106.600 ;
        RECT 98.290 105.320 103.120 105.460 ;
        RECT 98.290 105.275 98.580 105.320 ;
        RECT 102.830 105.300 103.120 105.320 ;
        RECT 103.910 105.460 104.200 105.505 ;
        RECT 107.490 105.460 107.780 105.505 ;
        RECT 109.325 105.460 109.615 105.505 ;
        RECT 103.910 105.320 109.615 105.460 ;
        RECT 103.910 105.275 104.200 105.320 ;
        RECT 107.490 105.275 107.780 105.320 ;
        RECT 109.325 105.275 109.615 105.320 ;
        RECT 109.775 105.260 110.095 105.520 ;
        RECT 133.100 105.500 136.850 105.630 ;
        RECT 50.910 105.120 51.200 105.165 ;
        RECT 54.575 105.120 54.895 105.180 ;
        RECT 50.910 104.980 54.895 105.120 ;
        RECT 50.910 104.935 51.200 104.980 ;
        RECT 54.575 104.920 54.895 104.980 ;
        RECT 57.795 105.120 58.115 105.180 ;
        RECT 59.650 105.120 59.940 105.165 ;
        RECT 57.795 104.980 59.940 105.120 ;
        RECT 57.795 104.920 58.115 104.980 ;
        RECT 59.650 104.935 59.940 104.980 ;
        RECT 61.490 105.120 61.780 105.165 ;
        RECT 62.855 105.120 63.175 105.180 ;
        RECT 61.490 104.980 63.175 105.120 ;
        RECT 61.490 104.935 61.780 104.980 ;
        RECT 62.855 104.920 63.175 104.980 ;
        RECT 71.610 105.120 71.900 105.165 ;
        RECT 73.895 105.120 74.215 105.180 ;
        RECT 84.015 105.120 84.335 105.180 ;
        RECT 71.610 104.980 84.335 105.120 ;
        RECT 71.610 104.935 71.900 104.980 ;
        RECT 73.895 104.920 74.215 104.980 ;
        RECT 84.015 104.920 84.335 104.980 ;
        RECT 84.490 105.120 84.780 105.165 ;
        RECT 85.855 105.120 86.175 105.180 ;
        RECT 84.490 104.980 86.175 105.120 ;
        RECT 84.490 104.935 84.780 104.980 ;
        RECT 85.855 104.920 86.175 104.980 ;
        RECT 99.195 105.120 99.515 105.180 ;
        RECT 99.670 105.120 99.960 105.165 ;
        RECT 99.195 104.980 99.960 105.120 ;
        RECT 99.195 104.920 99.515 104.980 ;
        RECT 99.670 104.935 99.960 104.980 ;
        RECT 55.150 104.780 55.440 104.825 ;
        RECT 58.270 104.780 58.560 104.825 ;
        RECT 60.160 104.780 60.450 104.825 ;
        RECT 49.605 104.640 53.195 104.780 ;
        RECT 37.980 104.595 38.270 104.640 ;
        RECT 39.870 104.595 40.160 104.640 ;
        RECT 42.990 104.595 43.280 104.640 ;
        RECT 39.395 104.440 39.715 104.500 ;
        RECT 25.225 104.300 39.715 104.440 ;
        RECT 53.055 104.440 53.195 104.640 ;
        RECT 55.150 104.640 60.450 104.780 ;
        RECT 55.150 104.595 55.440 104.640 ;
        RECT 58.270 104.595 58.560 104.640 ;
        RECT 60.160 104.595 60.450 104.640 ;
        RECT 65.730 104.780 66.020 104.825 ;
        RECT 68.850 104.780 69.140 104.825 ;
        RECT 70.740 104.780 71.030 104.825 ;
        RECT 65.730 104.640 71.030 104.780 ;
        RECT 65.730 104.595 66.020 104.640 ;
        RECT 68.850 104.595 69.140 104.640 ;
        RECT 70.740 104.595 71.030 104.640 ;
        RECT 78.150 104.780 78.440 104.825 ;
        RECT 81.270 104.780 81.560 104.825 ;
        RECT 83.160 104.780 83.450 104.825 ;
        RECT 78.150 104.640 83.450 104.780 ;
        RECT 78.150 104.595 78.440 104.640 ;
        RECT 81.270 104.595 81.560 104.640 ;
        RECT 83.160 104.595 83.450 104.640 ;
        RECT 88.730 104.780 89.020 104.825 ;
        RECT 91.850 104.780 92.140 104.825 ;
        RECT 93.740 104.780 94.030 104.825 ;
        RECT 88.730 104.640 94.030 104.780 ;
        RECT 88.730 104.595 89.020 104.640 ;
        RECT 91.850 104.595 92.140 104.640 ;
        RECT 93.740 104.595 94.030 104.640 ;
        RECT 103.910 104.780 104.200 104.825 ;
        RECT 107.030 104.780 107.320 104.825 ;
        RECT 108.920 104.780 109.210 104.825 ;
        RECT 103.910 104.640 109.210 104.780 ;
        RECT 103.910 104.595 104.200 104.640 ;
        RECT 107.030 104.595 107.320 104.640 ;
        RECT 108.920 104.595 109.210 104.640 ;
        RECT 59.175 104.440 59.495 104.500 ;
        RECT 53.055 104.300 59.495 104.440 ;
        RECT 39.395 104.240 39.715 104.300 ;
        RECT 59.175 104.240 59.495 104.300 ;
        RECT 96.895 104.240 97.215 104.500 ;
        RECT 18.165 103.620 112.465 104.100 ;
        RECT 37.095 103.420 37.415 103.480 ;
        RECT 37.095 103.280 47.445 103.420 ;
        RECT 37.095 103.220 37.415 103.280 ;
        RECT 26.630 103.080 26.920 103.125 ;
        RECT 29.750 103.080 30.040 103.125 ;
        RECT 31.640 103.080 31.930 103.125 ;
        RECT 33.415 103.080 33.735 103.140 ;
        RECT 37.185 103.080 37.325 103.220 ;
        RECT 26.630 102.940 31.930 103.080 ;
        RECT 26.630 102.895 26.920 102.940 ;
        RECT 29.750 102.895 30.040 102.940 ;
        RECT 31.640 102.895 31.930 102.940 ;
        RECT 32.585 102.940 37.325 103.080 ;
        RECT 41.350 103.080 41.640 103.125 ;
        RECT 44.470 103.080 44.760 103.125 ;
        RECT 46.360 103.080 46.650 103.125 ;
        RECT 41.350 102.940 46.650 103.080 ;
        RECT 27.435 102.740 27.755 102.800 ;
        RECT 32.585 102.785 32.725 102.940 ;
        RECT 33.415 102.880 33.735 102.940 ;
        RECT 41.350 102.895 41.640 102.940 ;
        RECT 44.470 102.895 44.760 102.940 ;
        RECT 46.360 102.895 46.650 102.940 ;
        RECT 31.130 102.740 31.420 102.785 ;
        RECT 27.435 102.600 31.420 102.740 ;
        RECT 27.435 102.540 27.755 102.600 ;
        RECT 31.130 102.555 31.420 102.600 ;
        RECT 32.510 102.555 32.800 102.785 ;
        RECT 37.110 102.740 37.400 102.785 ;
        RECT 39.855 102.740 40.175 102.800 ;
        RECT 37.110 102.600 40.175 102.740 ;
        RECT 37.110 102.555 37.400 102.600 ;
        RECT 39.855 102.540 40.175 102.600 ;
        RECT 45.835 102.540 46.155 102.800 ;
        RECT 47.305 102.785 47.445 103.280 ;
        RECT 55.955 103.220 56.275 103.480 ;
        RECT 57.795 103.220 58.115 103.480 ;
        RECT 59.635 103.220 59.955 103.480 ;
        RECT 71.135 103.220 71.455 103.480 ;
        RECT 72.515 103.220 72.835 103.480 ;
        RECT 79.415 103.420 79.735 103.480 ;
        RECT 84.950 103.420 85.240 103.465 ;
        RECT 79.415 103.280 85.240 103.420 ;
        RECT 79.415 103.220 79.735 103.280 ;
        RECT 84.950 103.235 85.240 103.280 ;
        RECT 87.250 103.420 87.540 103.465 ;
        RECT 87.695 103.420 88.015 103.480 ;
        RECT 95.055 103.420 95.375 103.480 ;
        RECT 87.250 103.280 88.015 103.420 ;
        RECT 87.250 103.235 87.540 103.280 ;
        RECT 87.695 103.220 88.015 103.280 ;
        RECT 88.245 103.280 95.375 103.420 ;
        RECT 78.150 103.080 78.440 103.125 ;
        RECT 81.270 103.080 81.560 103.125 ;
        RECT 83.160 103.080 83.450 103.125 ;
        RECT 78.150 102.940 83.450 103.080 ;
        RECT 78.150 102.895 78.440 102.940 ;
        RECT 81.270 102.895 81.560 102.940 ;
        RECT 83.160 102.895 83.450 102.940 ;
        RECT 47.230 102.555 47.520 102.785 ;
        RECT 73.910 102.740 74.200 102.785 ;
        RECT 76.655 102.740 76.975 102.800 ;
        RECT 73.910 102.600 76.975 102.740 ;
        RECT 73.910 102.555 74.200 102.600 ;
        RECT 76.655 102.540 76.975 102.600 ;
        RECT 80.335 102.740 80.655 102.800 ;
        RECT 82.650 102.740 82.940 102.785 ;
        RECT 80.335 102.600 82.940 102.740 ;
        RECT 80.335 102.540 80.655 102.600 ;
        RECT 82.650 102.555 82.940 102.600 ;
        RECT 84.015 102.540 84.335 102.800 ;
        RECT 22.835 102.400 23.155 102.460 ;
        RECT 25.550 102.400 25.840 102.420 ;
        RECT 22.835 102.260 25.840 102.400 ;
        RECT 22.835 102.200 23.155 102.260 ;
        RECT 21.455 102.060 21.775 102.120 ;
        RECT 25.550 102.105 25.840 102.260 ;
        RECT 26.630 102.400 26.920 102.445 ;
        RECT 30.210 102.400 30.500 102.445 ;
        RECT 32.045 102.400 32.335 102.445 ;
        RECT 40.315 102.420 40.635 102.460 ;
        RECT 26.630 102.260 32.335 102.400 ;
        RECT 26.630 102.215 26.920 102.260 ;
        RECT 30.210 102.215 30.500 102.260 ;
        RECT 32.045 102.215 32.335 102.260 ;
        RECT 40.270 102.200 40.635 102.420 ;
        RECT 41.350 102.400 41.640 102.445 ;
        RECT 44.930 102.400 45.220 102.445 ;
        RECT 46.765 102.400 47.055 102.445 ;
        RECT 41.350 102.260 47.055 102.400 ;
        RECT 41.350 102.215 41.640 102.260 ;
        RECT 44.930 102.215 45.220 102.260 ;
        RECT 46.765 102.215 47.055 102.260 ;
        RECT 56.430 102.215 56.720 102.445 ;
        RECT 40.270 102.105 40.560 102.200 ;
        RECT 22.390 102.060 22.680 102.105 ;
        RECT 21.455 101.920 22.680 102.060 ;
        RECT 21.455 101.860 21.775 101.920 ;
        RECT 22.390 101.875 22.680 101.920 ;
        RECT 25.250 102.060 25.840 102.105 ;
        RECT 28.490 102.060 29.140 102.105 ;
        RECT 25.250 101.920 29.140 102.060 ;
        RECT 25.250 101.875 25.540 101.920 ;
        RECT 28.490 101.875 29.140 101.920 ;
        RECT 39.970 102.060 40.560 102.105 ;
        RECT 43.210 102.060 43.860 102.105 ;
        RECT 39.970 101.920 43.860 102.060 ;
        RECT 56.505 102.060 56.645 102.215 ;
        RECT 56.875 102.200 57.195 102.460 ;
        RECT 59.175 102.200 59.495 102.460 ;
        RECT 71.610 102.400 71.900 102.445 ;
        RECT 72.070 102.400 72.360 102.445 ;
        RECT 71.610 102.260 75.505 102.400 ;
        RECT 71.610 102.215 71.900 102.260 ;
        RECT 72.070 102.215 72.360 102.260 ;
        RECT 59.265 102.060 59.405 102.200 ;
        RECT 56.505 101.920 59.405 102.060 ;
        RECT 39.970 101.875 40.260 101.920 ;
        RECT 43.210 101.875 43.860 101.920 ;
        RECT 75.365 101.720 75.505 102.260 ;
        RECT 75.735 102.060 76.055 102.120 ;
        RECT 77.070 102.105 77.360 102.420 ;
        RECT 78.150 102.400 78.440 102.445 ;
        RECT 81.730 102.400 82.020 102.445 ;
        RECT 83.565 102.400 83.855 102.445 ;
        RECT 78.150 102.260 83.855 102.400 ;
        RECT 78.150 102.215 78.440 102.260 ;
        RECT 81.730 102.215 82.020 102.260 ;
        RECT 83.565 102.215 83.855 102.260 ;
        RECT 85.410 102.400 85.700 102.445 ;
        RECT 86.790 102.400 87.080 102.445 ;
        RECT 88.245 102.400 88.385 103.280 ;
        RECT 95.055 103.220 95.375 103.280 ;
        RECT 92.870 103.080 93.160 103.125 ;
        RECT 95.990 103.080 96.280 103.125 ;
        RECT 97.880 103.080 98.170 103.125 ;
        RECT 92.870 102.940 98.170 103.080 ;
        RECT 92.870 102.895 93.160 102.940 ;
        RECT 95.990 102.895 96.280 102.940 ;
        RECT 97.880 102.895 98.170 102.940 ;
        RECT 101.460 103.080 101.750 103.125 ;
        RECT 103.350 103.080 103.640 103.125 ;
        RECT 106.470 103.080 106.760 103.125 ;
        RECT 101.460 102.940 106.760 103.080 ;
        RECT 101.460 102.895 101.750 102.940 ;
        RECT 103.350 102.895 103.640 102.940 ;
        RECT 106.470 102.895 106.760 102.940 ;
        RECT 88.630 102.740 88.920 102.785 ;
        RECT 95.055 102.740 95.375 102.800 ;
        RECT 88.630 102.600 95.375 102.740 ;
        RECT 88.630 102.555 88.920 102.600 ;
        RECT 95.055 102.540 95.375 102.600 ;
        RECT 97.355 102.540 97.675 102.800 ;
        RECT 98.735 102.740 99.055 102.800 ;
        RECT 100.590 102.740 100.880 102.785 ;
        RECT 98.735 102.600 100.880 102.740 ;
        RECT 98.735 102.540 99.055 102.600 ;
        RECT 100.590 102.555 100.880 102.600 ;
        RECT 101.970 102.740 102.260 102.785 ;
        RECT 105.175 102.740 105.495 102.800 ;
        RECT 101.970 102.600 105.495 102.740 ;
        RECT 101.970 102.555 102.260 102.600 ;
        RECT 105.175 102.540 105.495 102.600 ;
        RECT 85.410 102.260 88.385 102.400 ;
        RECT 85.410 102.215 85.700 102.260 ;
        RECT 86.790 102.215 87.080 102.260 ;
        RECT 76.770 102.060 77.360 102.105 ;
        RECT 80.010 102.060 80.660 102.105 ;
        RECT 75.735 101.920 80.660 102.060 ;
        RECT 75.735 101.860 76.055 101.920 ;
        RECT 76.770 101.875 77.060 101.920 ;
        RECT 80.010 101.875 80.660 101.920 ;
        RECT 78.035 101.720 78.355 101.780 ;
        RECT 85.485 101.720 85.625 102.215 ;
        RECT 91.790 102.105 92.080 102.420 ;
        RECT 92.870 102.400 93.160 102.445 ;
        RECT 96.450 102.400 96.740 102.445 ;
        RECT 98.285 102.400 98.575 102.445 ;
        RECT 92.870 102.260 98.575 102.400 ;
        RECT 92.870 102.215 93.160 102.260 ;
        RECT 96.450 102.215 96.740 102.260 ;
        RECT 98.285 102.215 98.575 102.260 ;
        RECT 101.055 102.400 101.345 102.445 ;
        RECT 102.890 102.400 103.180 102.445 ;
        RECT 106.470 102.400 106.760 102.445 ;
        RECT 101.055 102.260 106.760 102.400 ;
        RECT 101.055 102.215 101.345 102.260 ;
        RECT 102.890 102.215 103.180 102.260 ;
        RECT 106.470 102.215 106.760 102.260 ;
        RECT 91.490 102.060 92.080 102.105 ;
        RECT 94.730 102.060 95.380 102.105 ;
        RECT 96.895 102.060 97.215 102.120 ;
        RECT 91.490 101.920 97.215 102.060 ;
        RECT 91.490 101.875 91.780 101.920 ;
        RECT 94.730 101.875 95.380 101.920 ;
        RECT 96.895 101.860 97.215 101.920 ;
        RECT 103.335 102.060 103.655 102.120 ;
        RECT 107.550 102.105 107.840 102.420 ;
        RECT 104.250 102.060 104.900 102.105 ;
        RECT 107.550 102.060 108.140 102.105 ;
        RECT 103.335 101.920 108.140 102.060 ;
        RECT 103.335 101.860 103.655 101.920 ;
        RECT 104.250 101.875 104.900 101.920 ;
        RECT 107.850 101.875 108.140 101.920 ;
        RECT 108.855 102.060 109.175 102.120 ;
        RECT 110.710 102.060 111.000 102.105 ;
        RECT 108.855 101.920 111.000 102.060 ;
        RECT 108.855 101.860 109.175 101.920 ;
        RECT 110.710 101.875 111.000 101.920 ;
        RECT 75.365 101.580 85.625 101.720 ;
        RECT 78.035 101.520 78.355 101.580 ;
        RECT 17.370 100.900 112.465 101.380 ;
        RECT 133.330 76.630 136.060 77.830 ;
        RECT 137.920 77.810 143.450 77.960 ;
        RECT 21.115 74.380 23.065 74.390 ;
        RECT 19.415 73.240 23.065 74.380 ;
        RECT 19.415 73.230 21.125 73.240 ;
        RECT 28.135 73.230 30.305 74.410 ;
        RECT 32.315 74.390 34.265 74.400 ;
        RECT 30.615 73.250 34.265 74.390 ;
        RECT 30.615 73.240 32.325 73.250 ;
        RECT 39.425 73.200 41.595 74.380 ;
        RECT 43.535 74.360 45.485 74.370 ;
        RECT 41.835 73.220 45.485 74.360 ;
        RECT 54.785 74.340 56.735 74.350 ;
        RECT 41.835 73.210 43.545 73.220 ;
        RECT 3.910 73.080 6.100 73.190 ;
        RECT 50.005 73.140 52.175 74.320 ;
        RECT 53.085 73.200 56.735 74.340 ;
        RECT 53.085 73.190 54.795 73.200 ;
        RECT 61.425 73.170 63.595 74.350 ;
        RECT 66.005 74.330 67.955 74.340 ;
        RECT 64.305 73.190 67.955 74.330 ;
        RECT 64.305 73.180 66.015 73.190 ;
        RECT 72.535 73.180 74.705 74.360 ;
        RECT 77.245 74.320 79.195 74.330 ;
        RECT 75.545 73.180 79.195 74.320 ;
        RECT 75.545 73.170 77.255 73.180 ;
        RECT 83.805 73.170 85.975 74.350 ;
        RECT 88.495 74.330 90.445 74.340 ;
        RECT 86.795 73.190 90.445 74.330 ;
        RECT 99.775 74.320 101.725 74.330 ;
        RECT 86.795 73.180 88.505 73.190 ;
        RECT 94.995 73.110 97.165 74.290 ;
        RECT 98.075 73.180 101.725 74.320 ;
        RECT 98.075 73.170 99.785 73.180 ;
        RECT 106.405 73.160 108.575 74.340 ;
        RECT 111.045 74.320 112.995 74.330 ;
        RECT 109.345 73.180 112.995 74.320 ;
        RECT 109.345 73.170 111.055 73.180 ;
        RECT 117.605 73.160 119.775 74.340 ;
        RECT 122.295 74.320 124.245 74.330 ;
        RECT 120.595 73.180 124.245 74.320 ;
        RECT 129.455 73.240 131.625 74.420 ;
        RECT 120.595 73.170 122.305 73.180 ;
        RECT 3.910 72.820 12.240 73.080 ;
        RECT 29.635 72.840 43.235 72.850 ;
        RECT 18.435 72.820 43.235 72.840 ;
        RECT 3.910 72.800 54.455 72.820 ;
        RECT 3.910 72.790 65.705 72.800 ;
        RECT 133.960 72.790 135.640 76.630 ;
        RECT 137.190 76.610 143.450 77.810 ;
        RECT 137.920 75.460 143.450 76.610 ;
        RECT 3.910 72.780 76.925 72.790 ;
        RECT 85.815 72.780 99.415 72.790 ;
        RECT 132.085 72.780 140.600 72.790 ;
        RECT 3.910 71.700 140.600 72.780 ;
        RECT 3.910 71.690 32.035 71.700 ;
        RECT 3.910 71.670 19.135 71.690 ;
        RECT 40.855 71.670 140.600 71.700 ;
        RECT 3.910 71.500 12.240 71.670 ;
        RECT 52.105 71.650 140.600 71.670 ;
        RECT 63.325 71.640 140.600 71.650 ;
        RECT 74.565 71.630 88.165 71.640 ;
        RECT 97.095 71.630 133.215 71.640 ;
        RECT 3.910 71.370 6.100 71.500 ;
        RECT 10.800 71.180 11.950 71.500 ;
        RECT 10.800 69.480 11.915 71.180 ;
        RECT 29.635 71.170 43.285 71.180 ;
        RECT 15.510 71.155 17.040 71.160 ;
        RECT 18.435 71.155 43.285 71.170 ;
        RECT 12.285 71.150 43.285 71.155 ;
        RECT 12.285 71.130 54.505 71.150 ;
        RECT 141.810 71.140 143.230 75.460 ;
        RECT 12.285 71.120 65.755 71.130 ;
        RECT 12.285 71.110 76.975 71.120 ;
        RECT 85.815 71.110 99.465 71.120 ;
        RECT 140.220 71.110 143.240 71.140 ;
        RECT 12.285 70.030 143.240 71.110 ;
        RECT 12.285 70.020 32.085 70.030 ;
        RECT 12.285 70.005 19.375 70.020 ;
        RECT 10.800 13.800 11.950 69.480 ;
        RECT 12.320 15.450 13.470 70.005 ;
        RECT 15.510 68.660 17.040 70.005 ;
        RECT 40.855 70.000 143.240 70.030 ;
        RECT 52.105 69.980 143.240 70.000 ;
        RECT 63.325 69.970 143.240 69.980 ;
        RECT 74.565 69.960 88.215 69.970 ;
        RECT 97.095 69.960 143.240 69.970 ;
        RECT 140.220 69.910 143.240 69.960 ;
        RECT 29.645 69.670 43.315 69.680 ;
        RECT 18.445 69.650 43.315 69.670 ;
        RECT 18.445 69.630 54.535 69.650 ;
        RECT 18.445 69.620 65.785 69.630 ;
        RECT 139.590 69.620 150.610 69.640 ;
        RECT 18.445 69.610 77.005 69.620 ;
        RECT 85.825 69.610 99.495 69.620 ;
        RECT 132.155 69.610 150.610 69.620 ;
        RECT 18.445 69.570 150.610 69.610 ;
        RECT 18.445 68.530 150.740 69.570 ;
        RECT 18.445 68.520 32.115 68.530 ;
        RECT 40.865 68.500 150.740 68.530 ;
        RECT 52.115 68.490 143.320 68.500 ;
        RECT 52.115 68.480 140.670 68.490 ;
        RECT 63.335 68.470 140.670 68.480 ;
        RECT 74.575 68.460 88.245 68.470 ;
        RECT 97.105 68.460 133.295 68.470 ;
        RECT 141.080 68.450 142.300 68.490 ;
        RECT 149.360 68.470 150.740 68.500 ;
        RECT 29.655 68.100 43.325 68.110 ;
        RECT 13.950 68.080 43.325 68.100 ;
        RECT 13.950 68.060 54.545 68.080 ;
        RECT 13.950 68.050 65.795 68.060 ;
        RECT 13.950 68.040 77.015 68.050 ;
        RECT 85.835 68.040 99.505 68.050 ;
        RECT 139.530 68.040 143.320 68.060 ;
        RECT 13.950 66.960 152.870 68.040 ;
        RECT 13.950 66.950 32.125 66.960 ;
        RECT 13.950 18.530 15.100 66.950 ;
        RECT 40.875 66.930 152.870 66.960 ;
        RECT 52.125 66.910 152.870 66.930 ;
        RECT 63.345 66.900 152.870 66.910 ;
        RECT 74.585 66.890 88.255 66.900 ;
        RECT 97.115 66.890 143.320 66.900 ;
        RECT 141.030 66.770 142.490 66.890 ;
        RECT 21.405 65.510 26.555 65.790 ;
        RECT 27.815 65.490 28.965 65.800 ;
        RECT 32.605 65.520 37.755 65.800 ;
        RECT 39.015 65.500 40.165 65.810 ;
        RECT 43.825 65.490 48.975 65.770 ;
        RECT 50.235 65.470 51.385 65.780 ;
        RECT 149.460 65.760 150.600 65.780 ;
        RECT 55.075 65.470 60.225 65.750 ;
        RECT 61.485 65.450 62.635 65.760 ;
        RECT 66.295 65.460 71.445 65.740 ;
        RECT 72.705 65.440 73.855 65.750 ;
        RECT 77.535 65.450 82.685 65.730 ;
        RECT 83.945 65.430 85.095 65.740 ;
        RECT 88.785 65.460 93.935 65.740 ;
        RECT 95.195 65.440 96.345 65.750 ;
        RECT 100.065 65.450 105.215 65.730 ;
        RECT 106.475 65.430 107.625 65.740 ;
        RECT 111.335 65.450 116.485 65.730 ;
        RECT 117.745 65.430 118.895 65.740 ;
        RECT 122.585 65.450 127.735 65.730 ;
        RECT 128.995 65.430 130.145 65.740 ;
        RECT 133.315 65.430 138.455 65.690 ;
        RECT 21.205 65.140 21.435 65.320 ;
        RECT 26.495 65.190 26.725 65.320 ;
        RECT 21.125 55.220 21.485 65.140 ;
        RECT 26.435 55.240 26.805 65.190 ;
        RECT 27.635 65.150 27.865 65.320 ;
        RECT 27.565 55.200 27.935 65.150 ;
        RECT 28.925 65.140 29.155 65.320 ;
        RECT 32.405 65.150 32.635 65.330 ;
        RECT 37.695 65.200 37.925 65.330 ;
        RECT 28.835 55.250 29.255 65.140 ;
        RECT 32.325 55.230 32.685 65.150 ;
        RECT 37.635 55.250 38.005 65.200 ;
        RECT 38.835 65.160 39.065 65.330 ;
        RECT 38.765 55.210 39.135 65.160 ;
        RECT 40.125 65.150 40.355 65.330 ;
        RECT 40.035 55.260 40.455 65.150 ;
        RECT 43.625 65.120 43.855 65.300 ;
        RECT 48.915 65.170 49.145 65.300 ;
        RECT 43.545 55.200 43.905 65.120 ;
        RECT 48.855 55.220 49.225 65.170 ;
        RECT 50.055 65.130 50.285 65.300 ;
        RECT 49.985 55.180 50.355 65.130 ;
        RECT 51.345 65.120 51.575 65.300 ;
        RECT 51.255 55.230 51.675 65.120 ;
        RECT 54.875 65.100 55.105 65.280 ;
        RECT 60.165 65.150 60.395 65.280 ;
        RECT 54.795 55.180 55.155 65.100 ;
        RECT 60.105 55.200 60.475 65.150 ;
        RECT 61.305 65.110 61.535 65.280 ;
        RECT 61.235 55.160 61.605 65.110 ;
        RECT 62.595 65.100 62.825 65.280 ;
        RECT 62.505 55.210 62.925 65.100 ;
        RECT 66.095 65.090 66.325 65.270 ;
        RECT 71.385 65.140 71.615 65.270 ;
        RECT 66.015 55.170 66.375 65.090 ;
        RECT 71.325 55.190 71.695 65.140 ;
        RECT 72.525 65.100 72.755 65.270 ;
        RECT 72.455 55.150 72.825 65.100 ;
        RECT 73.815 65.090 74.045 65.270 ;
        RECT 73.725 55.200 74.145 65.090 ;
        RECT 77.335 65.080 77.565 65.260 ;
        RECT 82.625 65.130 82.855 65.260 ;
        RECT 77.255 55.160 77.615 65.080 ;
        RECT 82.565 55.180 82.935 65.130 ;
        RECT 83.765 65.090 83.995 65.260 ;
        RECT 83.695 55.140 84.065 65.090 ;
        RECT 85.055 65.080 85.285 65.260 ;
        RECT 88.585 65.090 88.815 65.270 ;
        RECT 93.875 65.140 94.105 65.270 ;
        RECT 84.965 55.190 85.385 65.080 ;
        RECT 88.505 55.170 88.865 65.090 ;
        RECT 93.815 55.190 94.185 65.140 ;
        RECT 95.015 65.100 95.245 65.270 ;
        RECT 94.945 55.150 95.315 65.100 ;
        RECT 96.305 65.090 96.535 65.270 ;
        RECT 96.215 55.200 96.635 65.090 ;
        RECT 99.865 65.080 100.095 65.260 ;
        RECT 105.155 65.130 105.385 65.260 ;
        RECT 99.785 55.160 100.145 65.080 ;
        RECT 105.095 55.180 105.465 65.130 ;
        RECT 106.295 65.090 106.525 65.260 ;
        RECT 106.225 55.140 106.595 65.090 ;
        RECT 107.585 65.080 107.815 65.260 ;
        RECT 111.135 65.080 111.365 65.260 ;
        RECT 116.425 65.130 116.655 65.260 ;
        RECT 107.495 55.190 107.915 65.080 ;
        RECT 111.055 55.160 111.415 65.080 ;
        RECT 116.365 55.180 116.735 65.130 ;
        RECT 117.565 65.090 117.795 65.260 ;
        RECT 117.495 55.140 117.865 65.090 ;
        RECT 118.855 65.080 119.085 65.260 ;
        RECT 122.385 65.080 122.615 65.260 ;
        RECT 127.675 65.130 127.905 65.260 ;
        RECT 118.765 55.190 119.185 65.080 ;
        RECT 122.305 55.160 122.665 65.080 ;
        RECT 127.615 55.180 127.985 65.130 ;
        RECT 128.815 65.090 129.045 65.260 ;
        RECT 128.745 55.140 129.115 65.090 ;
        RECT 130.105 65.080 130.335 65.260 ;
        RECT 133.135 65.130 133.365 65.230 ;
        RECT 130.015 55.190 130.435 65.080 ;
        RECT 133.005 55.240 133.405 65.130 ;
        RECT 138.425 65.100 138.655 65.230 ;
        RECT 133.135 55.230 133.365 55.240 ;
        RECT 138.345 55.130 138.725 65.100 ;
        RECT 149.340 64.660 150.720 65.760 ;
        RECT 20.815 54.230 25.555 54.530 ;
        RECT 32.015 54.240 36.755 54.540 ;
        RECT 43.235 54.210 47.975 54.510 ;
        RECT 54.485 54.190 59.225 54.490 ;
        RECT 65.705 54.180 70.445 54.480 ;
        RECT 76.945 54.170 81.685 54.470 ;
        RECT 88.195 54.180 92.935 54.480 ;
        RECT 99.475 54.170 104.215 54.470 ;
        RECT 110.745 54.170 115.485 54.470 ;
        RECT 121.995 54.170 126.735 54.470 ;
        RECT 21.655 52.320 22.115 52.550 ;
        RECT 25.625 52.280 26.255 52.560 ;
        RECT 25.735 52.240 26.195 52.280 ;
        RECT 27.665 52.240 28.125 52.470 ;
        RECT 32.855 52.330 33.315 52.560 ;
        RECT 36.825 52.290 37.455 52.570 ;
        RECT 36.935 52.250 37.395 52.290 ;
        RECT 38.865 52.250 39.325 52.480 ;
        RECT 44.075 52.300 44.535 52.530 ;
        RECT 48.045 52.260 48.675 52.540 ;
        RECT 48.155 52.220 48.615 52.260 ;
        RECT 50.085 52.220 50.545 52.450 ;
        RECT 55.325 52.280 55.785 52.510 ;
        RECT 59.295 52.240 59.925 52.520 ;
        RECT 59.405 52.200 59.865 52.240 ;
        RECT 61.335 52.200 61.795 52.430 ;
        RECT 66.545 52.270 67.005 52.500 ;
        RECT 70.515 52.230 71.145 52.510 ;
        RECT 70.625 52.190 71.085 52.230 ;
        RECT 72.555 52.190 73.015 52.420 ;
        RECT 77.785 52.260 78.245 52.490 ;
        RECT 81.755 52.220 82.385 52.500 ;
        RECT 81.865 52.180 82.325 52.220 ;
        RECT 83.795 52.180 84.255 52.410 ;
        RECT 89.035 52.270 89.495 52.500 ;
        RECT 93.005 52.230 93.635 52.510 ;
        RECT 93.115 52.190 93.575 52.230 ;
        RECT 95.045 52.190 95.505 52.420 ;
        RECT 100.315 52.260 100.775 52.490 ;
        RECT 104.285 52.220 104.915 52.500 ;
        RECT 104.395 52.180 104.855 52.220 ;
        RECT 106.325 52.180 106.785 52.410 ;
        RECT 111.585 52.260 112.045 52.490 ;
        RECT 115.555 52.220 116.185 52.500 ;
        RECT 115.665 52.180 116.125 52.220 ;
        RECT 117.595 52.180 118.055 52.410 ;
        RECT 122.835 52.260 123.295 52.490 ;
        RECT 126.805 52.220 127.435 52.500 ;
        RECT 126.915 52.180 127.375 52.220 ;
        RECT 128.845 52.180 129.305 52.410 ;
        RECT 21.375 52.010 21.605 52.115 ;
        RECT 21.245 50.290 21.615 52.010 ;
        RECT 22.165 51.890 22.395 52.115 ;
        RECT 25.455 51.980 25.685 52.035 ;
        RECT 21.375 50.115 21.605 50.290 ;
        RECT 22.155 50.210 22.525 51.890 ;
        RECT 22.165 50.115 22.395 50.210 ;
        RECT 21.525 49.670 22.245 49.930 ;
        RECT 19.295 46.650 20.065 47.720 ;
        RECT 21.385 47.490 22.105 47.750 ;
        RECT 21.225 47.200 21.455 47.340 ;
        RECT 21.085 46.430 21.475 47.200 ;
        RECT 22.015 47.190 22.245 47.340 ;
        RECT 22.005 46.450 22.375 47.190 ;
        RECT 25.305 47.010 25.735 51.980 ;
        RECT 26.245 51.970 26.475 52.035 ;
        RECT 27.385 51.970 27.615 52.035 ;
        RECT 26.185 46.970 26.585 51.970 ;
        RECT 27.265 46.970 27.665 51.970 ;
        RECT 28.175 51.940 28.405 52.035 ;
        RECT 32.575 52.020 32.805 52.125 ;
        RECT 28.115 46.970 28.545 51.940 ;
        RECT 32.445 50.300 32.815 52.020 ;
        RECT 33.365 51.900 33.595 52.125 ;
        RECT 36.655 51.990 36.885 52.045 ;
        RECT 32.575 50.125 32.805 50.300 ;
        RECT 33.355 50.220 33.725 51.900 ;
        RECT 33.365 50.125 33.595 50.220 ;
        RECT 32.725 49.680 33.445 49.940 ;
        RECT 25.735 46.600 26.195 46.830 ;
        RECT 27.665 46.710 28.125 46.830 ;
        RECT 27.515 46.600 28.125 46.710 ;
        RECT 30.495 46.660 31.265 47.730 ;
        RECT 32.585 47.500 33.305 47.760 ;
        RECT 32.425 47.210 32.655 47.350 ;
        RECT 21.225 46.340 21.455 46.430 ;
        RECT 22.015 46.340 22.245 46.450 ;
        RECT 27.515 46.430 28.095 46.600 ;
        RECT 32.285 46.440 32.675 47.210 ;
        RECT 33.215 47.200 33.445 47.350 ;
        RECT 33.205 46.460 33.575 47.200 ;
        RECT 36.505 47.020 36.935 51.990 ;
        RECT 37.445 51.980 37.675 52.045 ;
        RECT 38.585 51.980 38.815 52.045 ;
        RECT 37.385 46.980 37.785 51.980 ;
        RECT 38.465 46.980 38.865 51.980 ;
        RECT 39.375 51.950 39.605 52.045 ;
        RECT 43.795 51.990 44.025 52.095 ;
        RECT 39.315 46.980 39.745 51.950 ;
        RECT 43.665 50.270 44.035 51.990 ;
        RECT 44.585 51.870 44.815 52.095 ;
        RECT 47.875 51.960 48.105 52.015 ;
        RECT 43.795 50.095 44.025 50.270 ;
        RECT 44.575 50.190 44.945 51.870 ;
        RECT 44.585 50.095 44.815 50.190 ;
        RECT 43.945 49.650 44.665 49.910 ;
        RECT 36.935 46.610 37.395 46.840 ;
        RECT 38.865 46.720 39.325 46.840 ;
        RECT 38.715 46.610 39.325 46.720 ;
        RECT 41.715 46.630 42.485 47.700 ;
        RECT 43.805 47.470 44.525 47.730 ;
        RECT 43.645 47.180 43.875 47.320 ;
        RECT 32.425 46.350 32.655 46.440 ;
        RECT 33.215 46.350 33.445 46.460 ;
        RECT 38.715 46.440 39.295 46.610 ;
        RECT 43.505 46.410 43.895 47.180 ;
        RECT 44.435 47.170 44.665 47.320 ;
        RECT 44.425 46.430 44.795 47.170 ;
        RECT 47.725 46.990 48.155 51.960 ;
        RECT 48.665 51.950 48.895 52.015 ;
        RECT 49.805 51.950 50.035 52.015 ;
        RECT 48.605 46.950 49.005 51.950 ;
        RECT 49.685 46.950 50.085 51.950 ;
        RECT 50.595 51.920 50.825 52.015 ;
        RECT 55.045 51.970 55.275 52.075 ;
        RECT 50.535 46.950 50.965 51.920 ;
        RECT 54.915 50.250 55.285 51.970 ;
        RECT 55.835 51.850 56.065 52.075 ;
        RECT 59.125 51.940 59.355 51.995 ;
        RECT 55.045 50.075 55.275 50.250 ;
        RECT 55.825 50.170 56.195 51.850 ;
        RECT 55.835 50.075 56.065 50.170 ;
        RECT 55.195 49.630 55.915 49.890 ;
        RECT 48.155 46.580 48.615 46.810 ;
        RECT 50.085 46.690 50.545 46.810 ;
        RECT 49.935 46.580 50.545 46.690 ;
        RECT 52.965 46.610 53.735 47.680 ;
        RECT 55.055 47.450 55.775 47.710 ;
        RECT 54.895 47.160 55.125 47.300 ;
        RECT 43.645 46.320 43.875 46.410 ;
        RECT 44.435 46.320 44.665 46.430 ;
        RECT 49.935 46.410 50.515 46.580 ;
        RECT 54.755 46.390 55.145 47.160 ;
        RECT 55.685 47.150 55.915 47.300 ;
        RECT 55.675 46.410 56.045 47.150 ;
        RECT 58.975 46.970 59.405 51.940 ;
        RECT 59.915 51.930 60.145 51.995 ;
        RECT 61.055 51.930 61.285 51.995 ;
        RECT 59.855 46.930 60.255 51.930 ;
        RECT 60.935 46.930 61.335 51.930 ;
        RECT 61.845 51.900 62.075 51.995 ;
        RECT 66.265 51.960 66.495 52.065 ;
        RECT 61.785 46.930 62.215 51.900 ;
        RECT 66.135 50.240 66.505 51.960 ;
        RECT 67.055 51.840 67.285 52.065 ;
        RECT 70.345 51.930 70.575 51.985 ;
        RECT 66.265 50.065 66.495 50.240 ;
        RECT 67.045 50.160 67.415 51.840 ;
        RECT 67.055 50.065 67.285 50.160 ;
        RECT 66.415 49.620 67.135 49.880 ;
        RECT 59.405 46.560 59.865 46.790 ;
        RECT 61.335 46.670 61.795 46.790 ;
        RECT 61.185 46.560 61.795 46.670 ;
        RECT 64.185 46.600 64.955 47.670 ;
        RECT 66.275 47.440 66.995 47.700 ;
        RECT 66.115 47.150 66.345 47.290 ;
        RECT 54.895 46.300 55.125 46.390 ;
        RECT 55.685 46.300 55.915 46.410 ;
        RECT 61.185 46.390 61.765 46.560 ;
        RECT 65.975 46.380 66.365 47.150 ;
        RECT 66.905 47.140 67.135 47.290 ;
        RECT 66.895 46.400 67.265 47.140 ;
        RECT 70.195 46.960 70.625 51.930 ;
        RECT 71.135 51.920 71.365 51.985 ;
        RECT 72.275 51.920 72.505 51.985 ;
        RECT 71.075 46.920 71.475 51.920 ;
        RECT 72.155 46.920 72.555 51.920 ;
        RECT 73.065 51.890 73.295 51.985 ;
        RECT 77.505 51.950 77.735 52.055 ;
        RECT 73.005 46.920 73.435 51.890 ;
        RECT 77.375 50.230 77.745 51.950 ;
        RECT 78.295 51.830 78.525 52.055 ;
        RECT 81.585 51.920 81.815 51.975 ;
        RECT 77.505 50.055 77.735 50.230 ;
        RECT 78.285 50.150 78.655 51.830 ;
        RECT 78.295 50.055 78.525 50.150 ;
        RECT 77.655 49.610 78.375 49.870 ;
        RECT 70.625 46.550 71.085 46.780 ;
        RECT 72.555 46.660 73.015 46.780 ;
        RECT 72.405 46.550 73.015 46.660 ;
        RECT 75.425 46.590 76.195 47.660 ;
        RECT 77.515 47.430 78.235 47.690 ;
        RECT 77.355 47.140 77.585 47.280 ;
        RECT 66.115 46.290 66.345 46.380 ;
        RECT 66.905 46.290 67.135 46.400 ;
        RECT 72.405 46.380 72.985 46.550 ;
        RECT 77.215 46.370 77.605 47.140 ;
        RECT 78.145 47.130 78.375 47.280 ;
        RECT 78.135 46.390 78.505 47.130 ;
        RECT 81.435 46.950 81.865 51.920 ;
        RECT 82.375 51.910 82.605 51.975 ;
        RECT 83.515 51.910 83.745 51.975 ;
        RECT 82.315 46.910 82.715 51.910 ;
        RECT 83.395 46.910 83.795 51.910 ;
        RECT 84.305 51.880 84.535 51.975 ;
        RECT 88.755 51.960 88.985 52.065 ;
        RECT 84.245 46.910 84.675 51.880 ;
        RECT 88.625 50.240 88.995 51.960 ;
        RECT 89.545 51.840 89.775 52.065 ;
        RECT 92.835 51.930 93.065 51.985 ;
        RECT 88.755 50.065 88.985 50.240 ;
        RECT 89.535 50.160 89.905 51.840 ;
        RECT 89.545 50.065 89.775 50.160 ;
        RECT 88.905 49.620 89.625 49.880 ;
        RECT 81.865 46.540 82.325 46.770 ;
        RECT 83.795 46.650 84.255 46.770 ;
        RECT 83.645 46.540 84.255 46.650 ;
        RECT 86.675 46.600 87.445 47.670 ;
        RECT 88.765 47.440 89.485 47.700 ;
        RECT 88.605 47.150 88.835 47.290 ;
        RECT 77.355 46.280 77.585 46.370 ;
        RECT 78.145 46.280 78.375 46.390 ;
        RECT 83.645 46.370 84.225 46.540 ;
        RECT 88.465 46.380 88.855 47.150 ;
        RECT 89.395 47.140 89.625 47.290 ;
        RECT 89.385 46.400 89.755 47.140 ;
        RECT 92.685 46.960 93.115 51.930 ;
        RECT 93.625 51.920 93.855 51.985 ;
        RECT 94.765 51.920 94.995 51.985 ;
        RECT 93.565 46.920 93.965 51.920 ;
        RECT 94.645 46.920 95.045 51.920 ;
        RECT 95.555 51.890 95.785 51.985 ;
        RECT 100.035 51.950 100.265 52.055 ;
        RECT 95.495 46.920 95.925 51.890 ;
        RECT 99.905 50.230 100.275 51.950 ;
        RECT 100.825 51.830 101.055 52.055 ;
        RECT 104.115 51.920 104.345 51.975 ;
        RECT 100.035 50.055 100.265 50.230 ;
        RECT 100.815 50.150 101.185 51.830 ;
        RECT 100.825 50.055 101.055 50.150 ;
        RECT 100.185 49.610 100.905 49.870 ;
        RECT 93.115 46.550 93.575 46.780 ;
        RECT 95.045 46.660 95.505 46.780 ;
        RECT 94.895 46.550 95.505 46.660 ;
        RECT 97.955 46.590 98.725 47.660 ;
        RECT 100.045 47.430 100.765 47.690 ;
        RECT 99.885 47.140 100.115 47.280 ;
        RECT 88.605 46.290 88.835 46.380 ;
        RECT 89.395 46.290 89.625 46.400 ;
        RECT 94.895 46.380 95.475 46.550 ;
        RECT 99.745 46.370 100.135 47.140 ;
        RECT 100.675 47.130 100.905 47.280 ;
        RECT 100.665 46.390 101.035 47.130 ;
        RECT 103.965 46.950 104.395 51.920 ;
        RECT 104.905 51.910 105.135 51.975 ;
        RECT 106.045 51.910 106.275 51.975 ;
        RECT 104.845 46.910 105.245 51.910 ;
        RECT 105.925 46.910 106.325 51.910 ;
        RECT 106.835 51.880 107.065 51.975 ;
        RECT 111.305 51.950 111.535 52.055 ;
        RECT 106.775 46.910 107.205 51.880 ;
        RECT 111.175 50.230 111.545 51.950 ;
        RECT 112.095 51.830 112.325 52.055 ;
        RECT 115.385 51.920 115.615 51.975 ;
        RECT 111.305 50.055 111.535 50.230 ;
        RECT 112.085 50.150 112.455 51.830 ;
        RECT 112.095 50.055 112.325 50.150 ;
        RECT 111.455 49.610 112.175 49.870 ;
        RECT 104.395 46.540 104.855 46.770 ;
        RECT 106.325 46.650 106.785 46.770 ;
        RECT 106.175 46.540 106.785 46.650 ;
        RECT 109.225 46.590 109.995 47.660 ;
        RECT 111.315 47.430 112.035 47.690 ;
        RECT 111.155 47.140 111.385 47.280 ;
        RECT 99.885 46.280 100.115 46.370 ;
        RECT 100.675 46.280 100.905 46.390 ;
        RECT 106.175 46.370 106.755 46.540 ;
        RECT 111.015 46.370 111.405 47.140 ;
        RECT 111.945 47.130 112.175 47.280 ;
        RECT 111.935 46.390 112.305 47.130 ;
        RECT 115.235 46.950 115.665 51.920 ;
        RECT 116.175 51.910 116.405 51.975 ;
        RECT 117.315 51.910 117.545 51.975 ;
        RECT 116.115 46.910 116.515 51.910 ;
        RECT 117.195 46.910 117.595 51.910 ;
        RECT 118.105 51.880 118.335 51.975 ;
        RECT 122.555 51.950 122.785 52.055 ;
        RECT 118.045 46.910 118.475 51.880 ;
        RECT 122.425 50.230 122.795 51.950 ;
        RECT 123.345 51.830 123.575 52.055 ;
        RECT 126.635 51.920 126.865 51.975 ;
        RECT 122.555 50.055 122.785 50.230 ;
        RECT 123.335 50.150 123.705 51.830 ;
        RECT 123.345 50.055 123.575 50.150 ;
        RECT 122.705 49.610 123.425 49.870 ;
        RECT 115.665 46.540 116.125 46.770 ;
        RECT 117.595 46.650 118.055 46.770 ;
        RECT 117.445 46.540 118.055 46.650 ;
        RECT 120.475 46.590 121.245 47.660 ;
        RECT 122.565 47.430 123.285 47.690 ;
        RECT 122.405 47.140 122.635 47.280 ;
        RECT 111.155 46.280 111.385 46.370 ;
        RECT 111.945 46.280 112.175 46.390 ;
        RECT 117.445 46.370 118.025 46.540 ;
        RECT 122.265 46.370 122.655 47.140 ;
        RECT 123.195 47.130 123.425 47.280 ;
        RECT 123.185 46.390 123.555 47.130 ;
        RECT 126.485 46.950 126.915 51.920 ;
        RECT 127.425 51.910 127.655 51.975 ;
        RECT 128.565 51.910 128.795 51.975 ;
        RECT 127.365 46.910 127.765 51.910 ;
        RECT 128.445 46.910 128.845 51.910 ;
        RECT 129.355 51.880 129.585 51.975 ;
        RECT 129.295 46.910 129.725 51.880 ;
        RECT 126.915 46.540 127.375 46.770 ;
        RECT 128.845 46.650 129.305 46.770 ;
        RECT 128.695 46.540 129.305 46.650 ;
        RECT 122.405 46.280 122.635 46.370 ;
        RECT 123.195 46.280 123.425 46.390 ;
        RECT 128.695 46.370 129.275 46.540 ;
        RECT 21.505 45.950 21.965 46.180 ;
        RECT 32.705 45.960 33.165 46.190 ;
        RECT 43.925 45.930 44.385 46.160 ;
        RECT 55.175 45.910 55.635 46.140 ;
        RECT 66.395 45.900 66.855 46.130 ;
        RECT 77.635 45.890 78.095 46.120 ;
        RECT 88.885 45.900 89.345 46.130 ;
        RECT 100.165 45.890 100.625 46.120 ;
        RECT 111.435 45.890 111.895 46.120 ;
        RECT 122.685 45.890 123.145 46.120 ;
        RECT 29.055 45.020 41.225 45.030 ;
        RECT 17.855 45.005 41.225 45.020 ;
        RECT 15.900 45.000 41.225 45.005 ;
        RECT 15.900 44.980 52.445 45.000 ;
        RECT 15.900 44.970 63.695 44.980 ;
        RECT 15.900 44.960 74.915 44.970 ;
        RECT 85.235 44.960 97.405 44.970 ;
        RECT 15.900 43.880 131.205 44.960 ;
        RECT 15.900 43.870 30.025 43.880 ;
        RECT 15.900 43.855 18.690 43.870 ;
        RECT 15.900 41.620 17.050 43.855 ;
        RECT 40.275 43.850 131.205 43.880 ;
        RECT 51.525 43.830 131.205 43.850 ;
        RECT 62.745 43.820 131.205 43.830 ;
        RECT 73.985 43.810 86.155 43.820 ;
        RECT 96.515 43.810 131.205 43.820 ;
        RECT 29.015 43.330 41.185 43.340 ;
        RECT 17.815 43.310 41.185 43.330 ;
        RECT 142.830 43.320 144.150 43.340 ;
        RECT 17.815 43.290 52.405 43.310 ;
        RECT 140.750 43.300 144.150 43.320 ;
        RECT 17.815 43.280 63.655 43.290 ;
        RECT 119.895 43.280 144.150 43.300 ;
        RECT 17.815 43.270 74.875 43.280 ;
        RECT 85.195 43.270 97.365 43.280 ;
        RECT 108.685 43.270 144.150 43.280 ;
        RECT 17.815 42.180 144.150 43.270 ;
        RECT 18.755 42.150 144.150 42.180 ;
        RECT 18.755 42.120 131.165 42.150 ;
        RECT 18.755 42.090 109.655 42.120 ;
        RECT 18.755 42.080 98.445 42.090 ;
        RECT 41.325 42.070 98.445 42.080 ;
        RECT 142.830 42.070 144.150 42.150 ;
        RECT 41.325 42.060 87.205 42.070 ;
        RECT 75.035 42.050 87.205 42.060 ;
        RECT 15.900 41.540 19.685 41.620 ;
        RECT 142.070 41.610 146.210 41.640 ;
        RECT 119.855 41.590 146.210 41.610 ;
        RECT 108.645 41.550 146.210 41.590 ;
        RECT 15.900 41.520 42.165 41.540 ;
        RECT 97.445 41.530 146.210 41.550 ;
        RECT 15.900 41.510 75.875 41.520 ;
        RECT 86.235 41.510 146.210 41.530 ;
        RECT 15.900 40.500 146.210 41.510 ;
        RECT 15.900 40.480 142.320 40.500 ;
        RECT 15.900 40.470 140.920 40.480 ;
        RECT 18.715 40.460 140.920 40.470 ;
        RECT 142.070 40.460 142.250 40.480 ;
        RECT 18.715 40.440 120.815 40.460 ;
        RECT 18.715 40.400 109.615 40.440 ;
        RECT 18.715 40.390 98.405 40.400 ;
        RECT 41.285 40.380 98.405 40.390 ;
        RECT 41.285 40.370 87.165 40.380 ;
        RECT 74.995 40.360 87.165 40.370 ;
        RECT 26.775 39.230 27.235 39.460 ;
        RECT 38.055 39.230 38.515 39.460 ;
        RECT 49.345 39.210 49.805 39.440 ;
        RECT 60.565 39.210 61.025 39.440 ;
        RECT 71.765 39.210 72.225 39.440 ;
        RECT 83.055 39.200 83.515 39.430 ;
        RECT 94.295 39.220 94.755 39.450 ;
        RECT 105.505 39.240 105.965 39.470 ;
        RECT 116.705 39.280 117.165 39.510 ;
        RECT 127.915 39.300 128.375 39.530 ;
        RECT 20.645 38.810 21.225 38.980 ;
        RECT 26.495 38.960 26.725 39.070 ;
        RECT 27.285 38.980 27.515 39.070 ;
        RECT 20.615 38.700 21.225 38.810 ;
        RECT 20.615 38.580 21.075 38.700 ;
        RECT 22.545 38.580 23.005 38.810 ;
        RECT 20.195 33.470 20.625 38.440 ;
        RECT 20.335 33.375 20.565 33.470 ;
        RECT 21.075 33.440 21.475 38.440 ;
        RECT 22.155 33.440 22.555 38.440 ;
        RECT 21.125 33.375 21.355 33.440 ;
        RECT 22.265 33.375 22.495 33.440 ;
        RECT 23.005 33.430 23.435 38.400 ;
        RECT 26.365 38.220 26.735 38.960 ;
        RECT 26.495 38.070 26.725 38.220 ;
        RECT 27.265 38.210 27.655 38.980 ;
        RECT 31.925 38.810 32.505 38.980 ;
        RECT 37.775 38.960 38.005 39.070 ;
        RECT 38.565 38.980 38.795 39.070 ;
        RECT 27.285 38.070 27.515 38.210 ;
        RECT 26.635 37.660 27.355 37.920 ;
        RECT 28.675 37.690 29.445 38.760 ;
        RECT 31.895 38.700 32.505 38.810 ;
        RECT 31.895 38.580 32.355 38.700 ;
        RECT 33.825 38.580 34.285 38.810 ;
        RECT 26.495 35.480 27.215 35.740 ;
        RECT 26.345 35.200 26.575 35.295 ;
        RECT 26.215 33.520 26.585 35.200 ;
        RECT 27.135 35.120 27.365 35.295 ;
        RECT 23.055 33.375 23.285 33.430 ;
        RECT 26.345 33.295 26.575 33.520 ;
        RECT 27.125 33.400 27.495 35.120 ;
        RECT 31.475 33.470 31.905 38.440 ;
        RECT 27.135 33.295 27.365 33.400 ;
        RECT 31.615 33.375 31.845 33.470 ;
        RECT 32.355 33.440 32.755 38.440 ;
        RECT 33.435 33.440 33.835 38.440 ;
        RECT 32.405 33.375 32.635 33.440 ;
        RECT 33.545 33.375 33.775 33.440 ;
        RECT 34.285 33.430 34.715 38.400 ;
        RECT 37.645 38.220 38.015 38.960 ;
        RECT 37.775 38.070 38.005 38.220 ;
        RECT 38.545 38.210 38.935 38.980 ;
        RECT 43.215 38.790 43.795 38.960 ;
        RECT 49.065 38.940 49.295 39.050 ;
        RECT 49.855 38.960 50.085 39.050 ;
        RECT 38.565 38.070 38.795 38.210 ;
        RECT 37.915 37.660 38.635 37.920 ;
        RECT 39.955 37.690 40.725 38.760 ;
        RECT 43.185 38.680 43.795 38.790 ;
        RECT 43.185 38.560 43.645 38.680 ;
        RECT 45.115 38.560 45.575 38.790 ;
        RECT 37.775 35.480 38.495 35.740 ;
        RECT 37.625 35.200 37.855 35.295 ;
        RECT 37.495 33.520 37.865 35.200 ;
        RECT 38.415 35.120 38.645 35.295 ;
        RECT 34.335 33.375 34.565 33.430 ;
        RECT 37.625 33.295 37.855 33.520 ;
        RECT 38.405 33.400 38.775 35.120 ;
        RECT 42.765 33.450 43.195 38.420 ;
        RECT 38.415 33.295 38.645 33.400 ;
        RECT 42.905 33.355 43.135 33.450 ;
        RECT 43.645 33.420 44.045 38.420 ;
        RECT 44.725 33.420 45.125 38.420 ;
        RECT 43.695 33.355 43.925 33.420 ;
        RECT 44.835 33.355 45.065 33.420 ;
        RECT 45.575 33.410 46.005 38.380 ;
        RECT 48.935 38.200 49.305 38.940 ;
        RECT 49.065 38.050 49.295 38.200 ;
        RECT 49.835 38.190 50.225 38.960 ;
        RECT 54.435 38.790 55.015 38.960 ;
        RECT 60.285 38.940 60.515 39.050 ;
        RECT 61.075 38.960 61.305 39.050 ;
        RECT 49.855 38.050 50.085 38.190 ;
        RECT 49.205 37.640 49.925 37.900 ;
        RECT 51.245 37.670 52.015 38.740 ;
        RECT 54.405 38.680 55.015 38.790 ;
        RECT 54.405 38.560 54.865 38.680 ;
        RECT 56.335 38.560 56.795 38.790 ;
        RECT 49.065 35.460 49.785 35.720 ;
        RECT 48.915 35.180 49.145 35.275 ;
        RECT 48.785 33.500 49.155 35.180 ;
        RECT 49.705 35.100 49.935 35.275 ;
        RECT 45.625 33.355 45.855 33.410 ;
        RECT 48.915 33.275 49.145 33.500 ;
        RECT 49.695 33.380 50.065 35.100 ;
        RECT 53.985 33.450 54.415 38.420 ;
        RECT 49.705 33.275 49.935 33.380 ;
        RECT 54.125 33.355 54.355 33.450 ;
        RECT 54.865 33.420 55.265 38.420 ;
        RECT 55.945 33.420 56.345 38.420 ;
        RECT 54.915 33.355 55.145 33.420 ;
        RECT 56.055 33.355 56.285 33.420 ;
        RECT 56.795 33.410 57.225 38.380 ;
        RECT 60.155 38.200 60.525 38.940 ;
        RECT 60.285 38.050 60.515 38.200 ;
        RECT 61.055 38.190 61.445 38.960 ;
        RECT 65.635 38.790 66.215 38.960 ;
        RECT 71.485 38.940 71.715 39.050 ;
        RECT 72.275 38.960 72.505 39.050 ;
        RECT 61.075 38.050 61.305 38.190 ;
        RECT 60.425 37.640 61.145 37.900 ;
        RECT 62.465 37.670 63.235 38.740 ;
        RECT 65.605 38.680 66.215 38.790 ;
        RECT 65.605 38.560 66.065 38.680 ;
        RECT 67.535 38.560 67.995 38.790 ;
        RECT 60.285 35.460 61.005 35.720 ;
        RECT 60.135 35.180 60.365 35.275 ;
        RECT 60.005 33.500 60.375 35.180 ;
        RECT 60.925 35.100 61.155 35.275 ;
        RECT 56.845 33.355 57.075 33.410 ;
        RECT 60.135 33.275 60.365 33.500 ;
        RECT 60.915 33.380 61.285 35.100 ;
        RECT 65.185 33.450 65.615 38.420 ;
        RECT 60.925 33.275 61.155 33.380 ;
        RECT 65.325 33.355 65.555 33.450 ;
        RECT 66.065 33.420 66.465 38.420 ;
        RECT 67.145 33.420 67.545 38.420 ;
        RECT 66.115 33.355 66.345 33.420 ;
        RECT 67.255 33.355 67.485 33.420 ;
        RECT 67.995 33.410 68.425 38.380 ;
        RECT 71.355 38.200 71.725 38.940 ;
        RECT 71.485 38.050 71.715 38.200 ;
        RECT 72.255 38.190 72.645 38.960 ;
        RECT 76.925 38.780 77.505 38.950 ;
        RECT 82.775 38.930 83.005 39.040 ;
        RECT 83.565 38.950 83.795 39.040 ;
        RECT 72.275 38.050 72.505 38.190 ;
        RECT 71.625 37.640 72.345 37.900 ;
        RECT 73.665 37.670 74.435 38.740 ;
        RECT 76.895 38.670 77.505 38.780 ;
        RECT 76.895 38.550 77.355 38.670 ;
        RECT 78.825 38.550 79.285 38.780 ;
        RECT 71.485 35.460 72.205 35.720 ;
        RECT 71.335 35.180 71.565 35.275 ;
        RECT 71.205 33.500 71.575 35.180 ;
        RECT 72.125 35.100 72.355 35.275 ;
        RECT 68.045 33.355 68.275 33.410 ;
        RECT 71.335 33.275 71.565 33.500 ;
        RECT 72.115 33.380 72.485 35.100 ;
        RECT 76.475 33.440 76.905 38.410 ;
        RECT 72.125 33.275 72.355 33.380 ;
        RECT 76.615 33.345 76.845 33.440 ;
        RECT 77.355 33.410 77.755 38.410 ;
        RECT 78.435 33.410 78.835 38.410 ;
        RECT 77.405 33.345 77.635 33.410 ;
        RECT 78.545 33.345 78.775 33.410 ;
        RECT 79.285 33.400 79.715 38.370 ;
        RECT 82.645 38.190 83.015 38.930 ;
        RECT 82.775 38.040 83.005 38.190 ;
        RECT 83.545 38.180 83.935 38.950 ;
        RECT 88.165 38.800 88.745 38.970 ;
        RECT 94.015 38.950 94.245 39.060 ;
        RECT 94.805 38.970 95.035 39.060 ;
        RECT 83.565 38.040 83.795 38.180 ;
        RECT 82.915 37.630 83.635 37.890 ;
        RECT 84.955 37.660 85.725 38.730 ;
        RECT 88.135 38.690 88.745 38.800 ;
        RECT 88.135 38.570 88.595 38.690 ;
        RECT 90.065 38.570 90.525 38.800 ;
        RECT 82.775 35.450 83.495 35.710 ;
        RECT 82.625 35.170 82.855 35.265 ;
        RECT 82.495 33.490 82.865 35.170 ;
        RECT 83.415 35.090 83.645 35.265 ;
        RECT 79.335 33.345 79.565 33.400 ;
        RECT 82.625 33.265 82.855 33.490 ;
        RECT 83.405 33.370 83.775 35.090 ;
        RECT 87.715 33.460 88.145 38.430 ;
        RECT 83.415 33.265 83.645 33.370 ;
        RECT 87.855 33.365 88.085 33.460 ;
        RECT 88.595 33.430 88.995 38.430 ;
        RECT 89.675 33.430 90.075 38.430 ;
        RECT 88.645 33.365 88.875 33.430 ;
        RECT 89.785 33.365 90.015 33.430 ;
        RECT 90.525 33.420 90.955 38.390 ;
        RECT 93.885 38.210 94.255 38.950 ;
        RECT 94.015 38.060 94.245 38.210 ;
        RECT 94.785 38.200 95.175 38.970 ;
        RECT 99.375 38.820 99.955 38.990 ;
        RECT 105.225 38.970 105.455 39.080 ;
        RECT 106.015 38.990 106.245 39.080 ;
        RECT 94.805 38.060 95.035 38.200 ;
        RECT 94.155 37.650 94.875 37.910 ;
        RECT 96.195 37.680 96.965 38.750 ;
        RECT 99.345 38.710 99.955 38.820 ;
        RECT 99.345 38.590 99.805 38.710 ;
        RECT 101.275 38.590 101.735 38.820 ;
        RECT 94.015 35.470 94.735 35.730 ;
        RECT 93.865 35.190 94.095 35.285 ;
        RECT 93.735 33.510 94.105 35.190 ;
        RECT 94.655 35.110 94.885 35.285 ;
        RECT 90.575 33.365 90.805 33.420 ;
        RECT 93.865 33.285 94.095 33.510 ;
        RECT 94.645 33.390 95.015 35.110 ;
        RECT 98.925 33.480 99.355 38.450 ;
        RECT 94.655 33.285 94.885 33.390 ;
        RECT 99.065 33.385 99.295 33.480 ;
        RECT 99.805 33.450 100.205 38.450 ;
        RECT 100.885 33.450 101.285 38.450 ;
        RECT 99.855 33.385 100.085 33.450 ;
        RECT 100.995 33.385 101.225 33.450 ;
        RECT 101.735 33.440 102.165 38.410 ;
        RECT 105.095 38.230 105.465 38.970 ;
        RECT 105.225 38.080 105.455 38.230 ;
        RECT 105.995 38.220 106.385 38.990 ;
        RECT 110.575 38.860 111.155 39.030 ;
        RECT 116.425 39.010 116.655 39.120 ;
        RECT 117.215 39.030 117.445 39.120 ;
        RECT 106.015 38.080 106.245 38.220 ;
        RECT 105.365 37.670 106.085 37.930 ;
        RECT 107.405 37.700 108.175 38.770 ;
        RECT 110.545 38.750 111.155 38.860 ;
        RECT 110.545 38.630 111.005 38.750 ;
        RECT 112.475 38.630 112.935 38.860 ;
        RECT 105.225 35.490 105.945 35.750 ;
        RECT 105.075 35.210 105.305 35.305 ;
        RECT 104.945 33.530 105.315 35.210 ;
        RECT 105.865 35.130 106.095 35.305 ;
        RECT 101.785 33.385 102.015 33.440 ;
        RECT 105.075 33.305 105.305 33.530 ;
        RECT 105.855 33.410 106.225 35.130 ;
        RECT 110.125 33.520 110.555 38.490 ;
        RECT 110.265 33.425 110.495 33.520 ;
        RECT 111.005 33.490 111.405 38.490 ;
        RECT 112.085 33.490 112.485 38.490 ;
        RECT 111.055 33.425 111.285 33.490 ;
        RECT 112.195 33.425 112.425 33.490 ;
        RECT 112.935 33.480 113.365 38.450 ;
        RECT 116.295 38.270 116.665 39.010 ;
        RECT 116.425 38.120 116.655 38.270 ;
        RECT 117.195 38.260 117.585 39.030 ;
        RECT 121.785 38.880 122.365 39.050 ;
        RECT 127.635 39.030 127.865 39.140 ;
        RECT 128.425 39.050 128.655 39.140 ;
        RECT 117.215 38.120 117.445 38.260 ;
        RECT 116.565 37.710 117.285 37.970 ;
        RECT 118.605 37.740 119.375 38.810 ;
        RECT 121.755 38.770 122.365 38.880 ;
        RECT 121.755 38.650 122.215 38.770 ;
        RECT 123.685 38.650 124.145 38.880 ;
        RECT 116.425 35.530 117.145 35.790 ;
        RECT 116.275 35.250 116.505 35.345 ;
        RECT 116.145 33.570 116.515 35.250 ;
        RECT 117.065 35.170 117.295 35.345 ;
        RECT 112.985 33.425 113.215 33.480 ;
        RECT 105.865 33.305 106.095 33.410 ;
        RECT 116.275 33.345 116.505 33.570 ;
        RECT 117.055 33.450 117.425 35.170 ;
        RECT 121.335 33.540 121.765 38.510 ;
        RECT 117.065 33.345 117.295 33.450 ;
        RECT 121.475 33.445 121.705 33.540 ;
        RECT 122.215 33.510 122.615 38.510 ;
        RECT 123.295 33.510 123.695 38.510 ;
        RECT 122.265 33.445 122.495 33.510 ;
        RECT 123.405 33.445 123.635 33.510 ;
        RECT 124.145 33.500 124.575 38.470 ;
        RECT 127.505 38.290 127.875 39.030 ;
        RECT 127.635 38.140 127.865 38.290 ;
        RECT 128.405 38.280 128.795 39.050 ;
        RECT 128.425 38.140 128.655 38.280 ;
        RECT 127.775 37.730 128.495 37.990 ;
        RECT 129.815 37.760 130.585 38.830 ;
        RECT 142.850 37.630 144.170 38.900 ;
        RECT 127.635 35.550 128.355 35.810 ;
        RECT 127.485 35.270 127.715 35.365 ;
        RECT 127.355 33.590 127.725 35.270 ;
        RECT 128.275 35.190 128.505 35.365 ;
        RECT 124.195 33.445 124.425 33.500 ;
        RECT 127.485 33.365 127.715 33.590 ;
        RECT 128.265 33.470 128.635 35.190 ;
        RECT 128.275 33.365 128.505 33.470 ;
        RECT 20.615 32.940 21.075 33.170 ;
        RECT 22.545 33.130 23.005 33.170 ;
        RECT 22.485 32.850 23.115 33.130 ;
        RECT 26.625 32.860 27.085 33.090 ;
        RECT 31.895 32.940 32.355 33.170 ;
        RECT 33.825 33.130 34.285 33.170 ;
        RECT 33.765 32.850 34.395 33.130 ;
        RECT 37.905 32.860 38.365 33.090 ;
        RECT 43.185 32.920 43.645 33.150 ;
        RECT 45.115 33.110 45.575 33.150 ;
        RECT 45.055 32.830 45.685 33.110 ;
        RECT 49.195 32.840 49.655 33.070 ;
        RECT 54.405 32.920 54.865 33.150 ;
        RECT 56.335 33.110 56.795 33.150 ;
        RECT 56.275 32.830 56.905 33.110 ;
        RECT 60.415 32.840 60.875 33.070 ;
        RECT 65.605 32.920 66.065 33.150 ;
        RECT 67.535 33.110 67.995 33.150 ;
        RECT 67.475 32.830 68.105 33.110 ;
        RECT 71.615 32.840 72.075 33.070 ;
        RECT 76.895 32.910 77.355 33.140 ;
        RECT 78.825 33.100 79.285 33.140 ;
        RECT 78.765 32.820 79.395 33.100 ;
        RECT 82.905 32.830 83.365 33.060 ;
        RECT 88.135 32.930 88.595 33.160 ;
        RECT 90.065 33.120 90.525 33.160 ;
        RECT 90.005 32.840 90.635 33.120 ;
        RECT 94.145 32.850 94.605 33.080 ;
        RECT 99.345 32.950 99.805 33.180 ;
        RECT 101.275 33.140 101.735 33.180 ;
        RECT 101.215 32.860 101.845 33.140 ;
        RECT 105.355 32.870 105.815 33.100 ;
        RECT 110.545 32.990 111.005 33.220 ;
        RECT 112.475 33.180 112.935 33.220 ;
        RECT 112.415 32.900 113.045 33.180 ;
        RECT 116.555 32.910 117.015 33.140 ;
        RECT 121.755 33.010 122.215 33.240 ;
        RECT 123.685 33.200 124.145 33.240 ;
        RECT 123.625 32.920 124.255 33.200 ;
        RECT 127.765 32.930 128.225 33.160 ;
        RECT 23.185 30.880 27.925 31.180 ;
        RECT 34.465 30.880 39.205 31.180 ;
        RECT 45.755 30.860 50.495 31.160 ;
        RECT 56.975 30.860 61.715 31.160 ;
        RECT 68.175 30.860 72.915 31.160 ;
        RECT 79.465 30.850 84.205 31.150 ;
        RECT 90.705 30.870 95.445 31.170 ;
        RECT 101.915 30.890 106.655 31.190 ;
        RECT 113.115 30.930 117.855 31.230 ;
        RECT 124.325 30.950 129.065 31.250 ;
        RECT 19.485 20.270 19.905 30.160 ;
        RECT 19.585 20.090 19.815 20.270 ;
        RECT 20.805 20.260 21.175 30.210 ;
        RECT 20.875 20.090 21.105 20.260 ;
        RECT 21.935 20.220 22.305 30.170 ;
        RECT 27.255 20.270 27.615 30.190 ;
        RECT 30.765 20.270 31.185 30.160 ;
        RECT 22.015 20.090 22.245 20.220 ;
        RECT 27.305 20.090 27.535 20.270 ;
        RECT 30.865 20.090 31.095 20.270 ;
        RECT 32.085 20.260 32.455 30.210 ;
        RECT 32.155 20.090 32.385 20.260 ;
        RECT 33.215 20.220 33.585 30.170 ;
        RECT 38.535 20.270 38.895 30.190 ;
        RECT 33.295 20.090 33.525 20.220 ;
        RECT 38.585 20.090 38.815 20.270 ;
        RECT 42.055 20.250 42.475 30.140 ;
        RECT 42.155 20.070 42.385 20.250 ;
        RECT 43.375 20.240 43.745 30.190 ;
        RECT 43.445 20.070 43.675 20.240 ;
        RECT 44.505 20.200 44.875 30.150 ;
        RECT 49.825 20.250 50.185 30.170 ;
        RECT 53.275 20.250 53.695 30.140 ;
        RECT 44.585 20.070 44.815 20.200 ;
        RECT 49.875 20.070 50.105 20.250 ;
        RECT 53.375 20.070 53.605 20.250 ;
        RECT 54.595 20.240 54.965 30.190 ;
        RECT 54.665 20.070 54.895 20.240 ;
        RECT 55.725 20.200 56.095 30.150 ;
        RECT 61.045 20.250 61.405 30.170 ;
        RECT 64.475 20.250 64.895 30.140 ;
        RECT 55.805 20.070 56.035 20.200 ;
        RECT 61.095 20.070 61.325 20.250 ;
        RECT 64.575 20.070 64.805 20.250 ;
        RECT 65.795 20.240 66.165 30.190 ;
        RECT 65.865 20.070 66.095 20.240 ;
        RECT 66.925 20.200 67.295 30.150 ;
        RECT 72.245 20.250 72.605 30.170 ;
        RECT 67.005 20.070 67.235 20.200 ;
        RECT 72.295 20.070 72.525 20.250 ;
        RECT 75.765 20.240 76.185 30.130 ;
        RECT 75.865 20.060 76.095 20.240 ;
        RECT 77.085 20.230 77.455 30.180 ;
        RECT 77.155 20.060 77.385 20.230 ;
        RECT 78.215 20.190 78.585 30.140 ;
        RECT 83.535 20.240 83.895 30.160 ;
        RECT 87.005 20.260 87.425 30.150 ;
        RECT 78.295 20.060 78.525 20.190 ;
        RECT 83.585 20.060 83.815 20.240 ;
        RECT 87.105 20.080 87.335 20.260 ;
        RECT 88.325 20.250 88.695 30.200 ;
        RECT 88.395 20.080 88.625 20.250 ;
        RECT 89.455 20.210 89.825 30.160 ;
        RECT 94.775 20.260 95.135 30.180 ;
        RECT 98.215 20.280 98.635 30.170 ;
        RECT 89.535 20.080 89.765 20.210 ;
        RECT 94.825 20.080 95.055 20.260 ;
        RECT 98.315 20.100 98.545 20.280 ;
        RECT 99.535 20.270 99.905 30.220 ;
        RECT 99.605 20.100 99.835 20.270 ;
        RECT 100.665 20.230 101.035 30.180 ;
        RECT 105.985 20.280 106.345 30.200 ;
        RECT 109.415 20.320 109.835 30.210 ;
        RECT 100.745 20.100 100.975 20.230 ;
        RECT 106.035 20.100 106.265 20.280 ;
        RECT 109.515 20.140 109.745 20.320 ;
        RECT 110.735 20.310 111.105 30.260 ;
        RECT 110.805 20.140 111.035 20.310 ;
        RECT 111.865 20.270 112.235 30.220 ;
        RECT 117.185 20.320 117.545 30.240 ;
        RECT 120.625 20.340 121.045 30.230 ;
        RECT 111.945 20.140 112.175 20.270 ;
        RECT 117.235 20.140 117.465 20.320 ;
        RECT 120.725 20.160 120.955 20.340 ;
        RECT 121.945 20.330 122.315 30.280 ;
        RECT 122.015 20.160 122.245 20.330 ;
        RECT 123.075 20.290 123.445 30.240 ;
        RECT 128.395 20.340 128.755 30.260 ;
        RECT 123.155 20.160 123.385 20.290 ;
        RECT 128.445 20.160 128.675 20.340 ;
        RECT 132.345 20.170 132.755 30.180 ;
        RECT 137.735 30.120 137.965 30.130 ;
        RECT 132.445 20.130 132.675 20.170 ;
        RECT 137.665 20.080 138.055 30.120 ;
        RECT 19.775 19.610 20.925 19.920 ;
        RECT 22.185 19.620 27.335 19.900 ;
        RECT 31.055 19.610 32.205 19.920 ;
        RECT 33.465 19.620 38.615 19.900 ;
        RECT 42.345 19.590 43.495 19.900 ;
        RECT 44.755 19.600 49.905 19.880 ;
        RECT 53.565 19.590 54.715 19.900 ;
        RECT 55.975 19.600 61.125 19.880 ;
        RECT 64.765 19.590 65.915 19.900 ;
        RECT 67.175 19.600 72.325 19.880 ;
        RECT 76.055 19.580 77.205 19.890 ;
        RECT 78.465 19.590 83.615 19.870 ;
        RECT 87.295 19.600 88.445 19.910 ;
        RECT 89.705 19.610 94.855 19.890 ;
        RECT 98.505 19.620 99.655 19.930 ;
        RECT 100.915 19.630 106.065 19.910 ;
        RECT 109.705 19.660 110.855 19.970 ;
        RECT 112.115 19.670 117.265 19.950 ;
        RECT 120.915 19.680 122.065 19.990 ;
        RECT 123.325 19.690 128.475 19.970 ;
        RECT 132.635 19.640 138.025 19.930 ;
        RECT 142.940 19.110 144.080 37.630 ;
        RECT 13.940 18.460 17.635 18.530 ;
        RECT 117.755 18.510 131.425 18.530 ;
        RECT 106.545 18.470 131.425 18.510 ;
        RECT 13.940 18.440 41.565 18.460 ;
        RECT 95.345 18.450 131.425 18.470 ;
        RECT 13.940 18.430 75.275 18.440 ;
        RECT 84.135 18.430 131.425 18.450 ;
        RECT 13.940 17.380 131.425 18.430 ;
        RECT 142.890 17.990 144.140 19.110 ;
        RECT 145.070 18.880 146.210 40.500 ;
        RECT 145.030 17.960 146.250 18.880 ;
        RECT 13.950 17.370 15.100 17.380 ;
        RECT 16.615 17.360 120.215 17.380 ;
        RECT 16.615 17.320 109.015 17.360 ;
        RECT 16.615 17.310 97.805 17.320 ;
        RECT 39.185 17.300 97.805 17.310 ;
        RECT 39.185 17.290 86.565 17.300 ;
        RECT 72.895 17.280 86.565 17.290 ;
        RECT 117.765 16.950 140.620 16.960 ;
        RECT 142.040 16.950 148.010 16.980 ;
        RECT 117.765 16.940 148.010 16.950 ;
        RECT 106.555 16.900 148.010 16.940 ;
        RECT 16.625 16.870 41.575 16.890 ;
        RECT 95.355 16.880 148.010 16.900 ;
        RECT 16.625 16.860 75.285 16.870 ;
        RECT 84.145 16.860 148.010 16.880 ;
        RECT 16.625 15.840 148.010 16.860 ;
        RECT 16.625 15.820 142.660 15.840 ;
        RECT 16.625 15.810 140.620 15.820 ;
        RECT 142.040 15.810 142.660 15.820 ;
        RECT 16.625 15.790 120.225 15.810 ;
        RECT 16.625 15.750 109.025 15.790 ;
        RECT 16.625 15.740 97.815 15.750 ;
        RECT 39.195 15.730 97.815 15.740 ;
        RECT 39.195 15.720 86.575 15.730 ;
        RECT 72.905 15.710 86.575 15.720 ;
        RECT 131.215 15.460 132.585 15.470 ;
        RECT 12.290 15.390 17.625 15.450 ;
        RECT 117.795 15.440 132.785 15.460 ;
        RECT 106.585 15.400 132.785 15.440 ;
        RECT 12.290 15.370 41.585 15.390 ;
        RECT 95.385 15.380 132.785 15.400 ;
        RECT 12.290 15.360 75.295 15.370 ;
        RECT 84.175 15.360 132.785 15.380 ;
        RECT 12.290 14.320 132.785 15.360 ;
        RECT 142.905 15.040 144.045 15.050 ;
        RECT 12.290 14.310 131.445 14.320 ;
        RECT 12.290 14.300 120.235 14.310 ;
        RECT 12.320 14.280 13.470 14.300 ;
        RECT 16.655 14.290 120.235 14.300 ;
        RECT 16.655 14.250 109.035 14.290 ;
        RECT 16.655 14.240 97.825 14.250 ;
        RECT 39.225 14.230 97.825 14.240 ;
        RECT 39.225 14.220 86.585 14.230 ;
        RECT 72.935 14.210 86.585 14.220 ;
        RECT 142.850 13.920 144.100 15.040 ;
        RECT 145.020 14.870 146.160 14.980 ;
        RECT 144.980 13.950 146.200 14.870 ;
        RECT 16.965 13.800 17.435 13.810 ;
        RECT 10.800 13.780 17.435 13.800 ;
        RECT 10.800 13.720 17.555 13.780 ;
        RECT 117.845 13.770 131.445 13.790 ;
        RECT 106.635 13.730 131.445 13.770 ;
        RECT 10.800 13.700 41.585 13.720 ;
        RECT 95.435 13.710 131.445 13.730 ;
        RECT 10.800 13.690 75.295 13.700 ;
        RECT 84.225 13.690 131.445 13.710 ;
        RECT 10.800 12.650 131.445 13.690 ;
        RECT 16.705 12.640 131.445 12.650 ;
        RECT 16.705 12.620 120.235 12.640 ;
        RECT 16.705 12.580 109.035 12.620 ;
        RECT 16.705 12.570 97.825 12.580 ;
        RECT 39.275 12.560 97.825 12.570 ;
        RECT 39.275 12.550 86.585 12.560 ;
        RECT 72.985 12.540 86.585 12.550 ;
        RECT 128.755 12.240 130.465 12.250 ;
        RECT 117.545 12.220 119.255 12.230 ;
        RECT 106.345 12.180 108.055 12.190 ;
        RECT 27.615 12.170 29.325 12.180 ;
        RECT 38.895 12.170 40.605 12.180 ;
        RECT 25.675 11.030 29.325 12.170 ;
        RECT 36.955 11.030 40.605 12.170 ;
        RECT 95.135 12.160 96.845 12.170 ;
        RECT 50.185 12.150 51.895 12.160 ;
        RECT 61.405 12.150 63.115 12.160 ;
        RECT 72.605 12.150 74.315 12.160 ;
        RECT 25.675 11.020 27.625 11.030 ;
        RECT 36.955 11.020 38.905 11.030 ;
        RECT 48.245 11.010 51.895 12.150 ;
        RECT 59.465 11.010 63.115 12.150 ;
        RECT 70.665 11.010 74.315 12.150 ;
        RECT 83.895 12.140 85.605 12.150 ;
        RECT 48.245 11.000 50.195 11.010 ;
        RECT 59.465 11.000 61.415 11.010 ;
        RECT 70.665 11.000 72.615 11.010 ;
        RECT 81.955 11.000 85.605 12.140 ;
        RECT 93.195 11.020 96.845 12.160 ;
        RECT 104.405 11.040 108.055 12.180 ;
        RECT 115.605 11.080 119.255 12.220 ;
        RECT 126.815 11.100 130.465 12.240 ;
        RECT 126.815 11.090 128.765 11.100 ;
        RECT 115.605 11.070 117.555 11.080 ;
        RECT 104.405 11.030 106.355 11.040 ;
        RECT 93.195 11.010 95.145 11.020 ;
        RECT 81.955 10.990 83.905 11.000 ;
        RECT 142.905 8.580 144.045 13.920 ;
        RECT 74.420 7.440 144.045 8.580 ;
        RECT 74.420 1.410 75.560 7.440 ;
        RECT 145.020 6.630 146.160 13.950 ;
        RECT 93.650 5.490 146.160 6.630 ;
        RECT 93.650 1.480 94.790 5.490 ;
        RECT 146.870 4.560 148.010 15.840 ;
        RECT 113.130 3.420 148.010 4.560 ;
        RECT 113.130 1.610 114.270 3.420 ;
        RECT 149.460 2.770 150.600 64.660 ;
        RECT 131.940 1.880 150.600 2.770 ;
        RECT 131.800 1.630 150.600 1.880 ;
        RECT 74.290 0.160 75.680 1.410 ;
        RECT 93.500 0.230 94.890 1.480 ;
        RECT 112.900 0.360 114.290 1.610 ;
        RECT 131.800 1.380 133.490 1.630 ;
        RECT 151.730 1.420 152.870 66.900 ;
        RECT 131.800 0.430 133.540 1.380 ;
        RECT 113.130 0.330 114.270 0.360 ;
        RECT 151.600 0.300 152.970 1.420 ;
        RECT 93.650 0.150 94.790 0.230 ;
      LAYER met2 ;
        RECT 135.390 223.830 136.740 225.230 ;
        RECT 138.180 223.760 139.530 225.160 ;
        RECT 143.230 223.790 144.580 225.190 ;
        RECT 17.400 193.435 18.940 193.805 ;
        RECT 40.975 193.435 42.515 193.805 ;
        RECT 64.550 193.435 66.090 193.805 ;
        RECT 88.125 193.435 89.665 193.805 ;
        RECT 29.185 190.715 30.725 191.085 ;
        RECT 52.760 190.715 54.300 191.085 ;
        RECT 76.335 190.715 77.875 191.085 ;
        RECT 99.910 190.715 101.450 191.085 ;
        RECT 59.665 189.210 59.925 189.530 ;
        RECT 17.400 187.995 18.940 188.365 ;
        RECT 40.975 187.995 42.515 188.365 ;
        RECT 59.725 187.150 59.865 189.210 ;
        RECT 68.865 188.530 69.125 188.850 ;
        RECT 64.550 187.995 66.090 188.365 ;
        RECT 59.665 186.830 59.925 187.150 ;
        RECT 56.445 185.810 56.705 186.130 ;
        RECT 59.205 185.810 59.465 186.130 ;
        RECT 29.185 185.275 30.725 185.645 ;
        RECT 52.760 185.275 54.300 185.645 ;
        RECT 56.505 183.750 56.645 185.810 ;
        RECT 59.265 184.090 59.405 185.810 ;
        RECT 59.205 183.770 59.465 184.090 ;
        RECT 52.305 183.430 52.565 183.750 ;
        RECT 56.445 183.430 56.705 183.750 ;
        RECT 17.400 182.555 18.940 182.925 ;
        RECT 40.975 182.555 42.515 182.925 ;
        RECT 29.185 179.835 30.725 180.205 ;
        RECT 52.365 178.990 52.505 183.430 ;
        RECT 59.265 181.710 59.405 183.770 ;
        RECT 55.065 181.390 55.325 181.710 ;
        RECT 59.205 181.390 59.465 181.710 ;
        RECT 52.760 179.835 54.300 180.205 ;
        RECT 49.085 178.670 49.345 178.990 ;
        RECT 52.305 178.670 52.565 178.990 ;
        RECT 48.625 177.990 48.885 178.310 ;
        RECT 43.565 177.650 43.825 177.970 ;
        RECT 44.025 177.650 44.285 177.970 ;
        RECT 17.400 177.115 18.940 177.485 ;
        RECT 40.975 177.115 42.515 177.485 ;
        RECT 43.625 176.610 43.765 177.650 ;
        RECT 43.565 176.290 43.825 176.610 ;
        RECT 38.965 175.610 39.225 175.930 ;
        RECT 44.085 175.670 44.225 177.650 ;
        RECT 48.685 176.950 48.825 177.990 ;
        RECT 48.625 176.630 48.885 176.950 ;
        RECT 49.145 176.270 49.285 178.670 ;
        RECT 51.385 178.330 51.645 178.650 ;
        RECT 51.445 176.950 51.585 178.330 ;
        RECT 51.385 176.630 51.645 176.950 ;
        RECT 49.085 175.950 49.345 176.270 ;
        RECT 50.465 175.950 50.725 176.270 ;
        RECT 51.385 175.950 51.645 176.270 ;
        RECT 29.185 174.395 30.725 174.765 ;
        RECT 39.025 173.210 39.165 175.610 ;
        RECT 43.625 175.530 44.225 175.670 ;
        RECT 25.165 172.890 25.425 173.210 ;
        RECT 38.965 172.890 39.225 173.210 ;
        RECT 17.400 171.675 18.940 172.045 ;
        RECT 25.225 170.830 25.365 172.890 ;
        RECT 43.625 172.870 43.765 175.530 ;
        RECT 49.145 175.250 49.285 175.950 ;
        RECT 47.245 174.930 47.505 175.250 ;
        RECT 49.085 174.930 49.345 175.250 ;
        RECT 47.305 174.230 47.445 174.930 ;
        RECT 47.245 173.910 47.505 174.230 ;
        RECT 43.565 172.550 43.825 172.870 ;
        RECT 38.965 172.210 39.225 172.530 ;
        RECT 31.665 171.450 33.645 171.590 ;
        RECT 25.165 170.510 25.425 170.830 ;
        RECT 28.845 170.510 29.105 170.830 ;
        RECT 31.145 170.510 31.405 170.830 ;
        RECT 17.400 166.235 18.940 166.605 ;
        RECT 21.485 165.410 21.745 165.730 ;
        RECT 17.400 160.795 18.940 161.165 ;
        RECT 21.545 160.630 21.685 165.410 ;
        RECT 25.225 162.330 25.365 170.510 ;
        RECT 27.925 170.170 28.185 170.490 ;
        RECT 25.625 167.450 25.885 167.770 ;
        RECT 25.685 165.050 25.825 167.450 ;
        RECT 27.005 167.110 27.265 167.430 ;
        RECT 27.065 166.070 27.205 167.110 ;
        RECT 27.985 166.830 28.125 170.170 ;
        RECT 28.385 169.830 28.645 170.150 ;
        RECT 28.445 167.430 28.585 169.830 ;
        RECT 28.385 167.110 28.645 167.430 ;
        RECT 27.985 166.690 28.585 166.830 ;
        RECT 27.005 165.750 27.265 166.070 ;
        RECT 27.465 165.410 27.725 165.730 ;
        RECT 25.625 164.730 25.885 165.050 ;
        RECT 26.085 164.050 26.345 164.370 ;
        RECT 26.145 163.350 26.285 164.050 ;
        RECT 26.085 163.030 26.345 163.350 ;
        RECT 27.525 163.010 27.665 165.410 ;
        RECT 27.465 162.690 27.725 163.010 ;
        RECT 23.325 162.010 23.585 162.330 ;
        RECT 23.785 162.010 24.045 162.330 ;
        RECT 25.165 162.010 25.425 162.330 ;
        RECT 21.485 160.310 21.745 160.630 ;
        RECT 20.565 156.910 20.825 157.230 ;
        RECT 17.400 155.355 18.940 155.725 ;
        RECT 20.625 151.450 20.765 156.910 ;
        RECT 23.385 156.550 23.525 162.010 ;
        RECT 23.845 160.290 23.985 162.010 ;
        RECT 27.925 161.670 28.185 161.990 ;
        RECT 25.625 161.330 25.885 161.650 ;
        RECT 23.785 159.970 24.045 160.290 ;
        RECT 23.845 157.230 23.985 159.970 ;
        RECT 25.685 159.950 25.825 161.330 ;
        RECT 25.625 159.630 25.885 159.950 ;
        RECT 27.985 157.910 28.125 161.670 ;
        RECT 27.925 157.590 28.185 157.910 ;
        RECT 28.445 157.310 28.585 166.690 ;
        RECT 28.905 164.370 29.045 170.510 ;
        RECT 29.185 168.955 30.725 169.325 ;
        RECT 31.205 168.305 31.345 170.510 ;
        RECT 31.135 167.935 31.415 168.305 ;
        RECT 31.665 165.050 31.805 171.450 ;
        RECT 32.125 170.830 32.725 170.910 ;
        RECT 32.065 170.770 32.725 170.830 ;
        RECT 32.065 170.510 32.325 170.770 ;
        RECT 32.585 165.390 32.725 170.770 ;
        RECT 32.985 170.510 33.245 170.830 ;
        RECT 33.045 168.110 33.185 170.510 ;
        RECT 33.505 170.490 33.645 171.450 ;
        RECT 33.445 170.170 33.705 170.490 ;
        RECT 38.505 168.470 38.765 168.790 ;
        RECT 32.985 167.790 33.245 168.110 ;
        RECT 36.205 167.450 36.465 167.770 ;
        RECT 34.365 166.770 34.625 167.090 ;
        RECT 35.285 166.770 35.545 167.090 ;
        RECT 32.525 165.070 32.785 165.390 ;
        RECT 31.605 164.730 31.865 165.050 ;
        RECT 28.845 164.050 29.105 164.370 ;
        RECT 29.185 163.515 30.725 163.885 ;
        RECT 31.665 161.990 31.805 164.730 ;
        RECT 31.605 161.670 31.865 161.990 ;
        RECT 31.145 159.970 31.405 160.290 ;
        RECT 28.845 158.610 29.105 158.930 ;
        RECT 23.785 156.910 24.045 157.230 ;
        RECT 27.985 157.170 28.585 157.310 ;
        RECT 23.325 156.230 23.585 156.550 ;
        RECT 27.005 156.230 27.265 156.550 ;
        RECT 26.545 155.890 26.805 156.210 ;
        RECT 26.605 154.510 26.745 155.890 ;
        RECT 26.545 154.190 26.805 154.510 ;
        RECT 27.065 153.490 27.205 156.230 ;
        RECT 27.465 154.530 27.725 154.850 ;
        RECT 27.005 153.170 27.265 153.490 ;
        RECT 27.525 152.130 27.665 154.530 ;
        RECT 27.465 151.810 27.725 152.130 ;
        RECT 20.565 151.130 20.825 151.450 ;
        RECT 17.400 149.915 18.940 150.285 ;
        RECT 20.625 149.070 20.765 151.130 ;
        RECT 22.405 150.790 22.665 151.110 ;
        RECT 22.465 149.750 22.605 150.790 ;
        RECT 27.525 149.750 27.665 151.810 ;
        RECT 22.405 149.430 22.665 149.750 ;
        RECT 27.465 149.430 27.725 149.750 ;
        RECT 20.565 148.750 20.825 149.070 ;
        RECT 27.005 148.750 27.265 149.070 ;
        RECT 22.865 148.070 23.125 148.390 ;
        RECT 26.085 148.070 26.345 148.390 ;
        RECT 22.925 146.010 23.065 148.070 ;
        RECT 22.865 145.690 23.125 146.010 ;
        RECT 17.400 144.475 18.940 144.845 ;
        RECT 23.785 143.310 24.045 143.630 ;
        RECT 23.325 139.910 23.585 140.230 ;
        RECT 17.400 139.035 18.940 139.405 ;
        RECT 23.385 138.870 23.525 139.910 ;
        RECT 23.325 138.550 23.585 138.870 ;
        RECT 22.865 137.870 23.125 138.190 ;
        RECT 21.025 136.850 21.285 137.170 ;
        RECT 21.085 134.790 21.225 136.850 ;
        RECT 21.025 134.470 21.285 134.790 ;
        RECT 20.105 134.130 20.365 134.450 ;
        RECT 17.400 133.595 18.940 133.965 ;
        RECT 20.165 130.030 20.305 134.130 ;
        RECT 22.925 132.750 23.065 137.870 ;
        RECT 22.865 132.430 23.125 132.750 ;
        RECT 20.105 129.710 20.365 130.030 ;
        RECT 21.485 129.370 21.745 129.690 ;
        RECT 17.400 128.155 18.940 128.525 ;
        RECT 21.545 127.310 21.685 129.370 ;
        RECT 22.865 129.030 23.125 129.350 ;
        RECT 21.485 126.990 21.745 127.310 ;
        RECT 20.565 126.650 20.825 126.970 ;
        RECT 20.625 125.270 20.765 126.650 ;
        RECT 20.565 124.950 20.825 125.270 ;
        RECT 17.400 122.715 18.940 123.085 ;
        RECT 21.545 118.810 21.685 126.990 ;
        RECT 22.925 126.290 23.065 129.030 ;
        RECT 22.865 125.970 23.125 126.290 ;
        RECT 22.925 124.250 23.065 125.970 ;
        RECT 22.865 123.930 23.125 124.250 ;
        RECT 22.925 122.630 23.065 123.930 ;
        RECT 22.925 122.490 23.525 122.630 ;
        RECT 21.945 121.890 22.205 122.210 ;
        RECT 22.005 119.830 22.145 121.890 ;
        RECT 22.865 121.550 23.125 121.870 ;
        RECT 22.925 119.830 23.065 121.550 ;
        RECT 21.945 119.510 22.205 119.830 ;
        RECT 22.865 119.510 23.125 119.830 ;
        RECT 23.385 119.150 23.525 122.490 ;
        RECT 23.325 118.830 23.585 119.150 ;
        RECT 21.485 118.490 21.745 118.810 ;
        RECT 17.400 117.275 18.940 117.645 ;
        RECT 21.545 116.430 21.685 118.490 ;
        RECT 21.485 116.110 21.745 116.430 ;
        RECT 21.945 116.110 22.205 116.430 ;
        RECT 21.545 113.790 21.685 116.110 ;
        RECT 22.005 114.390 22.145 116.110 ;
        RECT 21.945 114.070 22.205 114.390 ;
        RECT 21.545 113.650 22.145 113.790 ;
        RECT 22.005 113.370 22.145 113.650 ;
        RECT 21.945 113.050 22.205 113.370 ;
        RECT 17.400 111.835 18.940 112.205 ;
        RECT 22.005 111.330 22.145 113.050 ;
        RECT 23.325 112.710 23.585 113.030 ;
        RECT 23.385 111.670 23.525 112.710 ;
        RECT 23.325 111.350 23.585 111.670 ;
        RECT 21.945 111.010 22.205 111.330 ;
        RECT 23.845 110.990 23.985 143.310 ;
        RECT 26.145 143.290 26.285 148.070 ;
        RECT 27.065 145.330 27.205 148.750 ;
        RECT 27.005 145.010 27.265 145.330 ;
        RECT 26.545 143.650 26.805 143.970 ;
        RECT 26.085 142.970 26.345 143.290 ;
        RECT 25.625 137.870 25.885 138.190 ;
        RECT 24.245 132.430 24.505 132.750 ;
        RECT 24.305 130.710 24.445 132.430 ;
        RECT 24.245 130.390 24.505 130.710 ;
        RECT 25.685 130.370 25.825 137.870 ;
        RECT 26.145 137.510 26.285 142.970 ;
        RECT 26.605 140.910 26.745 143.650 ;
        RECT 27.065 143.290 27.205 145.010 ;
        RECT 27.005 142.970 27.265 143.290 ;
        RECT 26.545 140.590 26.805 140.910 ;
        RECT 26.605 137.850 26.745 140.590 ;
        RECT 27.005 139.910 27.265 140.230 ;
        RECT 27.065 138.870 27.205 139.910 ;
        RECT 27.985 139.890 28.125 157.170 ;
        RECT 28.385 154.190 28.645 154.510 ;
        RECT 28.445 152.470 28.585 154.190 ;
        RECT 28.385 152.150 28.645 152.470 ;
        RECT 28.385 151.470 28.645 151.790 ;
        RECT 28.445 148.730 28.585 151.470 ;
        RECT 28.905 151.450 29.045 158.610 ;
        RECT 29.185 158.075 30.725 158.445 ;
        RECT 29.185 152.635 30.725 153.005 ;
        RECT 28.845 151.130 29.105 151.450 ;
        RECT 31.205 149.750 31.345 159.970 ;
        RECT 31.665 156.550 31.805 161.670 ;
        RECT 34.425 161.650 34.565 166.770 ;
        RECT 35.345 162.670 35.485 166.770 ;
        RECT 35.745 162.690 36.005 163.010 ;
        RECT 35.285 162.350 35.545 162.670 ;
        RECT 32.525 161.330 32.785 161.650 ;
        RECT 34.365 161.330 34.625 161.650 ;
        RECT 32.065 159.630 32.325 159.950 ;
        RECT 31.605 156.230 31.865 156.550 ;
        RECT 31.665 153.490 31.805 156.230 ;
        RECT 32.125 156.210 32.265 159.630 ;
        RECT 32.585 156.890 32.725 161.330 ;
        RECT 32.985 159.290 33.245 159.610 ;
        RECT 33.045 157.230 33.185 159.290 ;
        RECT 33.905 158.950 34.165 159.270 ;
        RECT 33.965 157.570 34.105 158.950 ;
        RECT 33.905 157.250 34.165 157.570 ;
        RECT 32.985 156.910 33.245 157.230 ;
        RECT 32.525 156.570 32.785 156.890 ;
        RECT 35.805 156.550 35.945 162.690 ;
        RECT 36.265 157.910 36.405 167.450 ;
        RECT 36.665 166.770 36.925 167.090 ;
        RECT 36.725 166.070 36.865 166.770 ;
        RECT 36.665 165.750 36.925 166.070 ;
        RECT 37.125 164.730 37.385 165.050 ;
        RECT 36.665 162.350 36.925 162.670 ;
        RECT 36.725 159.610 36.865 162.350 ;
        RECT 37.185 162.330 37.325 164.730 ;
        RECT 37.585 164.390 37.845 164.710 ;
        RECT 38.045 164.390 38.305 164.710 ;
        RECT 37.125 162.010 37.385 162.330 ;
        RECT 37.645 160.630 37.785 164.390 ;
        RECT 38.105 162.670 38.245 164.390 ;
        RECT 38.045 162.350 38.305 162.670 ;
        RECT 38.565 162.070 38.705 168.470 ;
        RECT 39.025 167.430 39.165 172.210 ;
        RECT 40.975 171.675 42.515 172.045 ;
        RECT 39.425 171.190 39.685 171.510 ;
        RECT 38.965 167.110 39.225 167.430 ;
        RECT 39.485 167.090 39.625 171.190 ;
        RECT 39.885 170.170 40.145 170.490 ;
        RECT 39.425 166.770 39.685 167.090 ;
        RECT 39.485 165.050 39.625 166.770 ;
        RECT 39.945 165.730 40.085 170.170 ;
        RECT 40.345 167.790 40.605 168.110 ;
        RECT 42.635 167.935 42.915 168.305 ;
        RECT 40.405 167.625 40.545 167.790 ;
        RECT 40.335 167.255 40.615 167.625 ;
        RECT 39.885 165.410 40.145 165.730 ;
        RECT 39.425 164.730 39.685 165.050 ;
        RECT 39.945 163.010 40.085 165.410 ;
        RECT 39.885 162.690 40.145 163.010 ;
        RECT 40.405 162.330 40.545 167.255 ;
        RECT 40.975 166.235 42.515 166.605 ;
        RECT 42.705 162.330 42.845 167.935 ;
        RECT 43.625 167.510 43.765 172.550 ;
        RECT 44.945 172.210 45.205 172.530 ;
        RECT 46.325 172.210 46.585 172.530 ;
        RECT 44.485 170.510 44.745 170.830 ;
        RECT 44.025 169.490 44.285 169.810 ;
        RECT 44.085 168.110 44.225 169.490 ;
        RECT 44.025 167.790 44.285 168.110 ;
        RECT 43.625 167.370 44.225 167.510 ;
        RECT 43.565 162.350 43.825 162.670 ;
        RECT 40.345 162.240 40.605 162.330 ;
        RECT 38.105 161.930 38.705 162.070 ;
        RECT 39.485 162.100 40.605 162.240 ;
        RECT 37.585 160.310 37.845 160.630 ;
        RECT 36.665 159.290 36.925 159.610 ;
        RECT 36.665 158.610 36.925 158.930 ;
        RECT 36.205 157.590 36.465 157.910 ;
        RECT 35.745 156.230 36.005 156.550 ;
        RECT 32.065 155.890 32.325 156.210 ;
        RECT 32.125 154.170 32.265 155.890 ;
        RECT 32.065 153.850 32.325 154.170 ;
        RECT 31.605 153.170 31.865 153.490 ;
        RECT 32.065 153.170 32.325 153.490 ;
        RECT 31.665 150.770 31.805 153.170 ;
        RECT 32.125 151.790 32.265 153.170 ;
        RECT 36.725 151.790 36.865 158.610 ;
        RECT 37.645 156.890 37.785 160.310 ;
        RECT 37.585 156.570 37.845 156.890 ;
        RECT 32.065 151.470 32.325 151.790 ;
        RECT 36.665 151.470 36.925 151.790 ;
        RECT 31.605 150.450 31.865 150.770 ;
        RECT 34.365 150.450 34.625 150.770 ;
        RECT 31.145 149.430 31.405 149.750 ;
        RECT 31.665 148.730 31.805 150.450 ;
        RECT 32.065 148.750 32.325 149.070 ;
        RECT 32.985 148.750 33.245 149.070 ;
        RECT 28.385 148.410 28.645 148.730 ;
        RECT 31.605 148.410 31.865 148.730 ;
        RECT 29.185 147.195 30.725 147.565 ;
        RECT 31.665 146.350 31.805 148.410 ;
        RECT 31.605 146.030 31.865 146.350 ;
        RECT 31.145 145.690 31.405 146.010 ;
        RECT 31.205 144.310 31.345 145.690 ;
        RECT 31.145 143.990 31.405 144.310 ;
        RECT 31.145 143.310 31.405 143.630 ;
        RECT 29.185 141.755 30.725 142.125 ;
        RECT 31.205 140.910 31.345 143.310 ;
        RECT 31.145 140.590 31.405 140.910 ;
        RECT 27.925 139.570 28.185 139.890 ;
        RECT 27.005 138.550 27.265 138.870 ;
        RECT 31.205 138.530 31.345 140.590 ;
        RECT 31.665 140.570 31.805 146.030 ;
        RECT 32.125 146.010 32.265 148.750 ;
        RECT 33.045 147.030 33.185 148.750 ;
        RECT 32.985 146.710 33.245 147.030 ;
        RECT 34.425 146.010 34.565 150.450 ;
        RECT 35.285 149.090 35.545 149.410 ;
        RECT 35.345 146.690 35.485 149.090 ;
        RECT 35.285 146.370 35.545 146.690 ;
        RECT 36.725 146.350 36.865 151.470 ;
        RECT 37.125 151.130 37.385 151.450 ;
        RECT 37.185 150.770 37.325 151.130 ;
        RECT 37.125 150.450 37.385 150.770 ;
        RECT 37.185 146.690 37.325 150.450 ;
        RECT 37.125 146.370 37.385 146.690 ;
        RECT 36.665 146.030 36.925 146.350 ;
        RECT 37.575 146.175 37.855 146.545 ;
        RECT 37.645 146.010 37.785 146.175 ;
        RECT 32.065 145.690 32.325 146.010 ;
        RECT 34.365 145.690 34.625 146.010 ;
        RECT 37.585 145.690 37.845 146.010 ;
        RECT 36.205 145.010 36.465 145.330 ;
        RECT 37.585 145.010 37.845 145.330 ;
        RECT 35.745 140.590 36.005 140.910 ;
        RECT 31.605 140.250 31.865 140.570 ;
        RECT 33.905 140.250 34.165 140.570 ;
        RECT 32.065 139.570 32.325 139.890 ;
        RECT 32.525 139.570 32.785 139.890 ;
        RECT 31.605 138.550 31.865 138.870 ;
        RECT 31.145 138.210 31.405 138.530 ;
        RECT 26.545 137.530 26.805 137.850 ;
        RECT 26.085 137.190 26.345 137.510 ;
        RECT 26.145 135.380 26.285 137.190 ;
        RECT 29.185 136.315 30.725 136.685 ;
        RECT 27.005 135.380 27.265 135.470 ;
        RECT 26.145 135.240 27.265 135.380 ;
        RECT 27.005 135.150 27.265 135.240 ;
        RECT 26.545 133.110 26.805 133.430 ;
        RECT 25.625 130.050 25.885 130.370 ;
        RECT 26.605 129.010 26.745 133.110 ;
        RECT 27.065 131.470 27.205 135.150 ;
        RECT 31.205 135.130 31.345 138.210 ;
        RECT 31.665 136.150 31.805 138.550 ;
        RECT 31.605 135.830 31.865 136.150 ;
        RECT 32.125 135.130 32.265 139.570 ;
        RECT 32.585 138.530 32.725 139.570 ;
        RECT 32.525 138.210 32.785 138.530 ;
        RECT 33.965 136.150 34.105 140.250 ;
        RECT 34.365 137.530 34.625 137.850 ;
        RECT 33.905 135.830 34.165 136.150 ;
        RECT 31.145 134.810 31.405 135.130 ;
        RECT 32.065 134.810 32.325 135.130 ;
        RECT 32.985 134.810 33.245 135.130 ;
        RECT 27.465 134.470 27.725 134.790 ;
        RECT 27.525 132.070 27.665 134.470 ;
        RECT 32.525 133.340 32.785 133.430 ;
        RECT 33.045 133.340 33.185 134.810 ;
        RECT 34.425 134.790 34.565 137.530 ;
        RECT 34.365 134.470 34.625 134.790 ;
        RECT 32.525 133.200 33.185 133.340 ;
        RECT 32.525 133.110 32.785 133.200 ;
        RECT 34.425 132.410 34.565 134.470 ;
        RECT 35.285 134.130 35.545 134.450 ;
        RECT 35.345 132.750 35.485 134.130 ;
        RECT 35.285 132.430 35.545 132.750 ;
        RECT 34.365 132.090 34.625 132.410 ;
        RECT 27.465 131.750 27.725 132.070 ;
        RECT 27.065 131.330 27.665 131.470 ;
        RECT 32.065 131.410 32.325 131.730 ;
        RECT 26.995 129.855 27.275 130.225 ;
        RECT 27.525 130.030 27.665 131.330 ;
        RECT 29.185 130.875 30.725 131.245 ;
        RECT 27.005 129.710 27.265 129.855 ;
        RECT 27.465 129.710 27.725 130.030 ;
        RECT 26.545 128.690 26.805 129.010 ;
        RECT 28.845 128.690 29.105 129.010 ;
        RECT 26.085 124.270 26.345 124.590 ;
        RECT 24.705 120.530 24.965 120.850 ;
        RECT 24.765 119.490 24.905 120.530 ;
        RECT 24.705 119.170 24.965 119.490 ;
        RECT 24.765 118.810 24.905 119.170 ;
        RECT 26.145 119.150 26.285 124.270 ;
        RECT 28.905 123.910 29.045 128.690 ;
        RECT 32.125 127.990 32.265 131.410 ;
        RECT 32.525 128.690 32.785 129.010 ;
        RECT 32.065 127.670 32.325 127.990 ;
        RECT 31.145 126.990 31.405 127.310 ;
        RECT 29.185 125.435 30.725 125.805 ;
        RECT 31.205 124.590 31.345 126.990 ;
        RECT 32.125 125.350 32.265 127.670 ;
        RECT 31.665 125.270 32.265 125.350 ;
        RECT 31.605 125.210 32.265 125.270 ;
        RECT 31.605 124.950 31.865 125.210 ;
        RECT 32.585 124.590 32.725 128.690 ;
        RECT 34.425 127.310 34.565 132.090 ;
        RECT 34.365 126.990 34.625 127.310 ;
        RECT 31.145 124.270 31.405 124.590 ;
        RECT 32.525 124.270 32.785 124.590 ;
        RECT 33.445 124.270 33.705 124.590 ;
        RECT 28.845 123.590 29.105 123.910 ;
        RECT 32.985 121.890 33.245 122.210 ;
        RECT 29.185 119.995 30.725 120.365 ;
        RECT 26.085 118.830 26.345 119.150 ;
        RECT 31.605 118.830 31.865 119.150 ;
        RECT 24.705 118.490 24.965 118.810 ;
        RECT 25.625 118.490 25.885 118.810 ;
        RECT 25.685 113.370 25.825 118.490 ;
        RECT 26.145 114.390 26.285 118.830 ;
        RECT 31.145 118.490 31.405 118.810 ;
        RECT 31.205 116.430 31.345 118.490 ;
        RECT 31.665 116.770 31.805 118.830 ;
        RECT 32.065 117.810 32.325 118.130 ;
        RECT 31.605 116.450 31.865 116.770 ;
        RECT 31.145 116.110 31.405 116.430 ;
        RECT 28.385 115.090 28.645 115.410 ;
        RECT 26.085 114.070 26.345 114.390 ;
        RECT 25.625 113.050 25.885 113.370 ;
        RECT 25.685 111.670 25.825 113.050 ;
        RECT 25.625 111.350 25.885 111.670 ;
        RECT 23.785 110.670 24.045 110.990 ;
        RECT 26.145 110.650 26.285 114.070 ;
        RECT 28.445 111.330 28.585 115.090 ;
        RECT 29.185 114.555 30.725 114.925 ;
        RECT 28.385 111.010 28.645 111.330 ;
        RECT 28.845 111.010 29.105 111.330 ;
        RECT 31.205 111.070 31.345 116.110 ;
        RECT 31.665 115.410 31.805 116.450 ;
        RECT 31.605 115.090 31.865 115.410 ;
        RECT 32.125 113.370 32.265 117.810 ;
        RECT 33.045 117.110 33.185 121.890 ;
        RECT 33.505 119.830 33.645 124.270 ;
        RECT 34.425 124.250 34.565 126.990 ;
        RECT 34.365 123.930 34.625 124.250 ;
        RECT 34.365 120.530 34.625 120.850 ;
        RECT 34.425 119.830 34.565 120.530 ;
        RECT 33.445 119.510 33.705 119.830 ;
        RECT 34.365 119.510 34.625 119.830 ;
        RECT 33.905 118.150 34.165 118.470 ;
        RECT 32.985 116.790 33.245 117.110 ;
        RECT 33.965 116.770 34.105 118.150 ;
        RECT 33.905 116.450 34.165 116.770 ;
        RECT 32.525 115.430 32.785 115.750 ;
        RECT 32.585 113.710 32.725 115.430 ;
        RECT 35.805 115.410 35.945 140.590 ;
        RECT 36.265 140.570 36.405 145.010 ;
        RECT 37.645 144.310 37.785 145.010 ;
        RECT 37.585 143.990 37.845 144.310 ;
        RECT 37.645 141.250 37.785 143.990 ;
        RECT 37.585 140.930 37.845 141.250 ;
        RECT 36.205 140.250 36.465 140.570 ;
        RECT 36.665 139.910 36.925 140.230 ;
        RECT 36.725 134.450 36.865 139.910 ;
        RECT 37.575 135.295 37.855 135.665 ;
        RECT 37.645 135.130 37.785 135.295 ;
        RECT 37.585 134.810 37.845 135.130 ;
        RECT 36.665 134.130 36.925 134.450 ;
        RECT 38.105 134.310 38.245 161.930 ;
        RECT 38.505 161.330 38.765 161.650 ;
        RECT 38.565 156.890 38.705 161.330 ;
        RECT 39.485 156.890 39.625 162.100 ;
        RECT 40.345 162.010 40.605 162.100 ;
        RECT 42.645 162.010 42.905 162.330 ;
        RECT 43.625 162.185 43.765 162.350 ;
        RECT 43.555 161.815 43.835 162.185 ;
        RECT 40.975 160.795 42.515 161.165 ;
        RECT 39.885 159.970 40.145 160.290 ;
        RECT 38.505 156.570 38.765 156.890 ;
        RECT 38.565 154.510 38.705 156.570 ;
        RECT 38.955 156.375 39.235 156.745 ;
        RECT 39.425 156.570 39.685 156.890 ;
        RECT 39.025 154.850 39.165 156.375 ;
        RECT 39.485 154.850 39.625 156.570 ;
        RECT 39.945 155.190 40.085 159.970 ;
        RECT 43.105 159.630 43.365 159.950 ;
        RECT 40.805 159.290 41.065 159.610 ;
        RECT 41.725 159.290 41.985 159.610 ;
        RECT 40.345 157.425 40.605 157.570 ;
        RECT 40.335 157.055 40.615 157.425 ;
        RECT 40.865 156.630 41.005 159.290 ;
        RECT 41.785 156.890 41.925 159.290 ;
        RECT 43.165 157.570 43.305 159.630 ;
        RECT 43.105 157.250 43.365 157.570 ;
        RECT 40.405 156.490 41.005 156.630 ;
        RECT 41.725 156.570 41.985 156.890 ;
        RECT 39.885 154.870 40.145 155.190 ;
        RECT 38.965 154.530 39.225 154.850 ;
        RECT 39.425 154.530 39.685 154.850 ;
        RECT 38.505 154.190 38.765 154.510 ;
        RECT 39.425 153.170 39.685 153.490 ;
        RECT 38.505 151.810 38.765 152.130 ;
        RECT 39.485 151.870 39.625 153.170 ;
        RECT 38.565 149.410 38.705 151.810 ;
        RECT 39.485 151.730 40.085 151.870 ;
        RECT 38.965 150.450 39.225 150.770 ;
        RECT 38.505 149.090 38.765 149.410 ;
        RECT 39.025 148.390 39.165 150.450 ;
        RECT 38.965 148.070 39.225 148.390 ;
        RECT 39.025 146.545 39.165 148.070 ;
        RECT 38.955 146.175 39.235 146.545 ;
        RECT 39.425 145.690 39.685 146.010 ;
        RECT 38.505 143.990 38.765 144.310 ;
        RECT 38.565 143.290 38.705 143.990 ;
        RECT 39.485 143.970 39.625 145.690 ;
        RECT 39.425 143.650 39.685 143.970 ;
        RECT 38.505 142.970 38.765 143.290 ;
        RECT 38.965 142.970 39.225 143.290 ;
        RECT 39.025 141.590 39.165 142.970 ;
        RECT 38.965 141.270 39.225 141.590 ;
        RECT 39.425 141.270 39.685 141.590 ;
        RECT 38.505 137.190 38.765 137.510 ;
        RECT 38.565 135.470 38.705 137.190 ;
        RECT 38.965 136.850 39.225 137.170 ;
        RECT 38.505 135.150 38.765 135.470 ;
        RECT 38.565 134.790 38.705 135.150 ;
        RECT 38.505 134.470 38.765 134.790 ;
        RECT 37.185 134.170 38.245 134.310 ;
        RECT 37.185 133.090 37.325 134.170 ;
        RECT 37.125 132.770 37.385 133.090 ;
        RECT 38.505 132.430 38.765 132.750 ;
        RECT 37.585 130.050 37.845 130.370 ;
        RECT 36.665 129.370 36.925 129.690 ;
        RECT 36.725 127.990 36.865 129.370 ;
        RECT 37.125 128.690 37.385 129.010 ;
        RECT 36.665 127.670 36.925 127.990 ;
        RECT 37.185 125.350 37.325 128.690 ;
        RECT 36.725 125.210 37.325 125.350 ;
        RECT 36.725 118.810 36.865 125.210 ;
        RECT 37.125 123.250 37.385 123.570 ;
        RECT 37.185 121.530 37.325 123.250 ;
        RECT 37.125 121.210 37.385 121.530 ;
        RECT 36.665 118.490 36.925 118.810 ;
        RECT 36.665 115.770 36.925 116.090 ;
        RECT 33.445 115.090 33.705 115.410 ;
        RECT 35.745 115.090 36.005 115.410 ;
        RECT 32.525 113.390 32.785 113.710 ;
        RECT 33.505 113.370 33.645 115.090 ;
        RECT 36.725 114.390 36.865 115.770 ;
        RECT 36.665 114.070 36.925 114.390 ;
        RECT 32.065 113.050 32.325 113.370 ;
        RECT 33.445 113.050 33.705 113.370 ;
        RECT 36.665 113.110 36.925 113.370 ;
        RECT 37.185 113.110 37.325 121.210 ;
        RECT 37.645 119.830 37.785 130.050 ;
        RECT 38.565 129.690 38.705 132.430 ;
        RECT 38.505 129.370 38.765 129.690 ;
        RECT 39.025 121.270 39.165 136.850 ;
        RECT 39.485 127.220 39.625 141.270 ;
        RECT 39.945 138.270 40.085 151.730 ;
        RECT 40.405 149.070 40.545 156.490 ;
        RECT 43.105 155.890 43.365 156.210 ;
        RECT 43.565 156.065 43.825 156.210 ;
        RECT 40.975 155.355 42.515 155.725 ;
        RECT 40.805 154.870 41.065 155.190 ;
        RECT 40.865 150.770 41.005 154.870 ;
        RECT 42.635 154.335 42.915 154.705 ;
        RECT 43.165 154.420 43.305 155.890 ;
        RECT 43.555 155.695 43.835 156.065 ;
        RECT 43.565 154.420 43.825 154.510 ;
        RECT 42.645 154.190 42.905 154.335 ;
        RECT 43.165 154.280 43.825 154.420 ;
        RECT 43.565 154.190 43.825 154.280 ;
        RECT 42.705 151.450 42.845 154.190 ;
        RECT 43.625 151.450 43.765 154.190 ;
        RECT 44.085 151.450 44.225 167.370 ;
        RECT 44.545 166.070 44.685 170.510 ;
        RECT 44.485 165.750 44.745 166.070 ;
        RECT 45.005 165.390 45.145 172.210 ;
        RECT 46.385 171.170 46.525 172.210 ;
        RECT 46.325 170.850 46.585 171.170 ;
        RECT 44.945 165.070 45.205 165.390 ;
        RECT 45.005 162.670 45.145 165.070 ;
        RECT 44.485 162.350 44.745 162.670 ;
        RECT 44.945 162.350 45.205 162.670 ;
        RECT 42.645 151.130 42.905 151.450 ;
        RECT 43.565 151.130 43.825 151.450 ;
        RECT 44.025 151.130 44.285 151.450 ;
        RECT 40.805 150.450 41.065 150.770 ;
        RECT 42.645 150.450 42.905 150.770 ;
        RECT 40.975 149.915 42.515 150.285 ;
        RECT 40.345 148.750 40.605 149.070 ;
        RECT 40.405 143.630 40.545 148.750 ;
        RECT 40.975 144.475 42.515 144.845 ;
        RECT 41.725 143.650 41.985 143.970 ;
        RECT 40.345 143.310 40.605 143.630 ;
        RECT 41.265 142.970 41.525 143.290 ;
        RECT 40.795 142.095 41.075 142.465 ;
        RECT 40.335 140.735 40.615 141.105 ;
        RECT 40.345 140.590 40.605 140.735 ;
        RECT 40.865 140.230 41.005 142.095 ;
        RECT 41.325 140.910 41.465 142.970 ;
        RECT 41.785 141.250 41.925 143.650 ;
        RECT 41.725 140.930 41.985 141.250 ;
        RECT 41.265 140.590 41.525 140.910 ;
        RECT 42.185 140.425 42.445 140.570 ;
        RECT 40.805 139.910 41.065 140.230 ;
        RECT 42.175 140.055 42.455 140.425 ;
        RECT 40.975 139.035 42.515 139.405 ;
        RECT 42.185 138.385 42.445 138.530 ;
        RECT 39.945 138.130 41.005 138.270 ;
        RECT 39.885 135.830 40.145 136.150 ;
        RECT 39.945 133.430 40.085 135.830 ;
        RECT 40.865 134.310 41.005 138.130 ;
        RECT 42.175 138.015 42.455 138.385 ;
        RECT 42.705 137.850 42.845 150.450 ;
        RECT 43.565 148.070 43.825 148.390 ;
        RECT 43.105 145.865 43.365 146.010 ;
        RECT 43.095 145.495 43.375 145.865 ;
        RECT 43.105 145.010 43.365 145.330 ;
        RECT 43.165 143.630 43.305 145.010 ;
        RECT 43.105 143.310 43.365 143.630 ;
        RECT 43.625 143.290 43.765 148.070 ;
        RECT 44.015 146.175 44.295 146.545 ;
        RECT 44.025 146.030 44.285 146.175 ;
        RECT 44.025 145.350 44.285 145.670 ;
        RECT 43.565 142.970 43.825 143.290 ;
        RECT 43.105 142.290 43.365 142.610 ;
        RECT 42.645 137.530 42.905 137.850 ;
        RECT 43.165 137.080 43.305 142.290 ;
        RECT 43.565 139.570 43.825 139.890 ;
        RECT 42.175 136.655 42.455 137.025 ;
        RECT 42.705 136.940 43.305 137.080 ;
        RECT 42.245 135.130 42.385 136.655 ;
        RECT 41.715 134.615 41.995 134.985 ;
        RECT 42.185 134.810 42.445 135.130 ;
        RECT 41.785 134.450 41.925 134.615 ;
        RECT 40.405 134.170 41.005 134.310 ;
        RECT 39.885 133.110 40.145 133.430 ;
        RECT 40.405 132.150 40.545 134.170 ;
        RECT 41.725 134.130 41.985 134.450 ;
        RECT 40.975 133.595 42.515 133.965 ;
        RECT 42.185 132.430 42.445 132.750 ;
        RECT 40.405 132.010 41.005 132.150 ;
        RECT 40.345 131.410 40.605 131.730 ;
        RECT 40.405 130.710 40.545 131.410 ;
        RECT 40.345 130.390 40.605 130.710 ;
        RECT 40.865 129.690 41.005 132.010 ;
        RECT 41.725 131.410 41.985 131.730 ;
        RECT 42.245 131.470 42.385 132.430 ;
        RECT 42.705 132.150 42.845 136.940 ;
        RECT 43.105 135.380 43.365 135.470 ;
        RECT 43.625 135.380 43.765 139.570 ;
        RECT 44.085 138.385 44.225 145.350 ;
        RECT 44.545 144.310 44.685 162.350 ;
        RECT 45.405 162.010 45.665 162.330 ;
        RECT 45.865 162.010 46.125 162.330 ;
        RECT 45.465 159.950 45.605 162.010 ;
        RECT 45.925 159.950 46.065 162.010 ;
        RECT 46.385 159.950 46.525 170.850 ;
        RECT 49.145 170.830 49.285 174.930 ;
        RECT 50.525 173.890 50.665 175.950 ;
        RECT 51.445 175.250 51.585 175.950 ;
        RECT 52.365 175.930 52.505 178.670 ;
        RECT 55.125 176.610 55.265 181.390 ;
        RECT 52.825 176.270 53.425 176.350 ;
        RECT 55.065 176.290 55.325 176.610 ;
        RECT 58.745 176.290 59.005 176.610 ;
        RECT 52.825 176.210 53.485 176.270 ;
        RECT 52.305 175.610 52.565 175.930 ;
        RECT 52.825 175.590 52.965 176.210 ;
        RECT 53.225 175.950 53.485 176.210 ;
        RECT 57.365 175.610 57.625 175.930 ;
        RECT 52.765 175.270 53.025 175.590 ;
        RECT 51.385 174.930 51.645 175.250 ;
        RECT 51.845 174.930 52.105 175.250 ;
        RECT 50.465 173.570 50.725 173.890 ;
        RECT 49.545 173.230 49.805 173.550 ;
        RECT 48.165 170.510 48.425 170.830 ;
        RECT 49.085 170.510 49.345 170.830 ;
        RECT 46.785 167.790 47.045 168.110 ;
        RECT 47.235 167.935 47.515 168.305 ;
        RECT 46.845 167.625 46.985 167.790 ;
        RECT 47.305 167.770 47.445 167.935 ;
        RECT 46.775 167.255 47.055 167.625 ;
        RECT 47.245 167.450 47.505 167.770 ;
        RECT 47.705 167.450 47.965 167.770 ;
        RECT 47.765 165.730 47.905 167.450 ;
        RECT 47.705 165.410 47.965 165.730 ;
        RECT 46.785 164.050 47.045 164.370 ;
        RECT 46.845 161.990 46.985 164.050 ;
        RECT 47.245 162.010 47.505 162.330 ;
        RECT 46.785 161.670 47.045 161.990 ;
        RECT 47.305 159.950 47.445 162.010 ;
        RECT 45.405 159.630 45.665 159.950 ;
        RECT 45.865 159.630 46.125 159.950 ;
        RECT 46.325 159.630 46.585 159.950 ;
        RECT 47.245 159.630 47.505 159.950 ;
        RECT 44.945 158.785 45.205 158.930 ;
        RECT 44.935 158.415 45.215 158.785 ;
        RECT 45.465 156.890 45.605 159.630 ;
        RECT 45.405 156.570 45.665 156.890 ;
        RECT 44.945 156.230 45.205 156.550 ;
        RECT 44.485 143.990 44.745 144.310 ;
        RECT 44.485 143.310 44.745 143.630 ;
        RECT 44.545 142.610 44.685 143.310 ;
        RECT 44.485 142.290 44.745 142.610 ;
        RECT 44.485 140.930 44.745 141.250 ;
        RECT 44.015 138.015 44.295 138.385 ;
        RECT 44.545 137.760 44.685 140.930 ;
        RECT 43.105 135.240 43.765 135.380 ;
        RECT 44.085 137.620 44.685 137.760 ;
        RECT 43.105 135.150 43.365 135.240 ;
        RECT 43.565 134.130 43.825 134.450 ;
        RECT 43.095 133.255 43.375 133.625 ;
        RECT 43.105 133.110 43.365 133.255 ;
        RECT 43.625 132.410 43.765 134.130 ;
        RECT 44.085 132.750 44.225 137.620 ;
        RECT 44.485 136.850 44.745 137.170 ;
        RECT 44.025 132.430 44.285 132.750 ;
        RECT 42.705 132.010 43.305 132.150 ;
        RECT 43.565 132.090 43.825 132.410 ;
        RECT 41.785 130.030 41.925 131.410 ;
        RECT 42.245 131.330 42.845 131.470 ;
        RECT 41.725 129.710 41.985 130.030 ;
        RECT 39.875 129.175 40.155 129.545 ;
        RECT 40.805 129.370 41.065 129.690 ;
        RECT 39.885 129.030 40.145 129.175 ;
        RECT 40.345 128.690 40.605 129.010 ;
        RECT 39.485 127.080 40.085 127.220 ;
        RECT 39.425 125.970 39.685 126.290 ;
        RECT 39.485 121.870 39.625 125.970 ;
        RECT 39.425 121.550 39.685 121.870 ;
        RECT 38.105 121.130 39.165 121.270 ;
        RECT 37.585 119.510 37.845 119.830 ;
        RECT 36.665 113.050 37.325 113.110 ;
        RECT 37.585 113.050 37.845 113.370 ;
        RECT 36.725 112.970 37.325 113.050 ;
        RECT 26.085 110.330 26.345 110.650 ;
        RECT 27.465 109.650 27.725 109.970 ;
        RECT 26.085 107.950 26.345 108.270 ;
        RECT 24.245 107.270 24.505 107.590 ;
        RECT 17.400 106.395 18.940 106.765 ;
        RECT 24.305 106.230 24.445 107.270 ;
        RECT 24.245 105.910 24.505 106.230 ;
        RECT 22.865 104.210 23.125 104.530 ;
        RECT 22.925 102.490 23.065 104.210 ;
        RECT 22.865 102.170 23.125 102.490 ;
        RECT 21.485 101.830 21.745 102.150 ;
        RECT 17.400 100.955 18.940 101.325 ;
        RECT 21.545 98.340 21.685 101.830 ;
        RECT 26.145 98.340 26.285 107.950 ;
        RECT 27.525 102.830 27.665 109.650 ;
        RECT 27.925 106.930 28.185 107.250 ;
        RECT 27.985 105.890 28.125 106.930 ;
        RECT 28.905 106.230 29.045 111.010 ;
        RECT 30.745 110.990 31.345 111.070 ;
        RECT 30.685 110.930 31.345 110.990 ;
        RECT 30.685 110.670 30.945 110.930 ;
        RECT 37.185 110.650 37.325 112.970 ;
        RECT 37.645 112.690 37.785 113.050 ;
        RECT 37.585 112.370 37.845 112.690 ;
        RECT 31.145 110.330 31.405 110.650 ;
        RECT 37.125 110.330 37.385 110.650 ;
        RECT 29.185 109.115 30.725 109.485 ;
        RECT 28.845 105.910 29.105 106.230 ;
        RECT 27.925 105.570 28.185 105.890 ;
        RECT 29.185 103.675 30.725 104.045 ;
        RECT 31.205 103.080 31.345 110.330 ;
        RECT 33.445 107.610 33.705 107.930 ;
        RECT 32.985 105.120 33.245 105.210 ;
        RECT 33.505 105.120 33.645 107.610 ;
        RECT 37.185 105.210 37.325 110.330 ;
        RECT 38.105 107.930 38.245 121.130 ;
        RECT 39.945 119.490 40.085 127.080 ;
        RECT 39.885 119.170 40.145 119.490 ;
        RECT 38.505 115.430 38.765 115.750 ;
        RECT 38.565 112.690 38.705 115.430 ;
        RECT 38.965 112.710 39.225 113.030 ;
        RECT 38.505 112.370 38.765 112.690 ;
        RECT 39.025 111.670 39.165 112.710 ;
        RECT 38.965 111.350 39.225 111.670 ;
        RECT 40.405 110.990 40.545 128.690 ;
        RECT 40.975 128.155 42.515 128.525 ;
        RECT 42.185 126.650 42.445 126.970 ;
        RECT 41.725 126.310 41.985 126.630 ;
        RECT 41.785 124.930 41.925 126.310 ;
        RECT 41.725 124.610 41.985 124.930 ;
        RECT 42.245 124.590 42.385 126.650 ;
        RECT 42.185 124.270 42.445 124.590 ;
        RECT 40.975 122.715 42.515 123.085 ;
        RECT 40.975 117.275 42.515 117.645 ;
        RECT 41.265 116.110 41.525 116.430 ;
        RECT 41.325 113.370 41.465 116.110 ;
        RECT 41.265 113.050 41.525 113.370 ;
        RECT 40.975 111.835 42.515 112.205 ;
        RECT 40.345 110.670 40.605 110.990 ;
        RECT 40.805 109.650 41.065 109.970 ;
        RECT 40.865 108.950 41.005 109.650 ;
        RECT 40.805 108.630 41.065 108.950 ;
        RECT 38.505 108.290 38.765 108.610 ;
        RECT 38.045 107.610 38.305 107.930 ;
        RECT 38.045 106.930 38.305 107.250 ;
        RECT 38.105 105.890 38.245 106.930 ;
        RECT 38.565 105.890 38.705 108.290 ;
        RECT 42.705 107.930 42.845 131.330 ;
        RECT 43.165 122.550 43.305 132.010 ;
        RECT 44.015 131.895 44.295 132.265 ;
        RECT 43.565 131.410 43.825 131.730 ;
        RECT 43.625 130.710 43.765 131.410 ;
        RECT 43.565 130.390 43.825 130.710 ;
        RECT 44.085 129.690 44.225 131.895 ;
        RECT 44.025 129.370 44.285 129.690 ;
        RECT 43.565 128.690 43.825 129.010 ;
        RECT 44.025 128.865 44.285 129.010 ;
        RECT 43.625 127.310 43.765 128.690 ;
        RECT 44.015 128.495 44.295 128.865 ;
        RECT 44.025 127.330 44.285 127.650 ;
        RECT 43.565 126.990 43.825 127.310 ;
        RECT 43.565 123.250 43.825 123.570 ;
        RECT 43.105 122.230 43.365 122.550 ;
        RECT 43.625 113.370 43.765 123.250 ;
        RECT 44.085 122.210 44.225 127.330 ;
        RECT 44.545 125.270 44.685 136.850 ;
        RECT 45.005 134.450 45.145 156.230 ;
        RECT 45.925 155.190 46.065 159.630 ;
        RECT 45.865 154.870 46.125 155.190 ;
        RECT 47.305 154.170 47.445 159.630 ;
        RECT 47.765 158.930 47.905 165.410 ;
        RECT 48.225 165.390 48.365 170.510 ;
        RECT 49.605 170.490 49.745 173.230 ;
        RECT 51.905 172.870 52.045 174.930 ;
        RECT 52.760 174.395 54.300 174.765 ;
        RECT 57.425 173.550 57.565 175.610 ;
        RECT 58.805 174.230 58.945 176.290 ;
        RECT 58.745 173.910 59.005 174.230 ;
        RECT 57.365 173.230 57.625 173.550 ;
        RECT 55.525 172.890 55.785 173.210 ;
        RECT 51.845 172.550 52.105 172.870 ;
        RECT 55.585 171.510 55.725 172.890 ;
        RECT 55.525 171.190 55.785 171.510 ;
        RECT 50.465 170.510 50.725 170.830 ;
        RECT 49.545 170.170 49.805 170.490 ;
        RECT 49.085 169.490 49.345 169.810 ;
        RECT 48.625 167.110 48.885 167.430 ;
        RECT 48.165 165.070 48.425 165.390 ;
        RECT 48.685 161.650 48.825 167.110 ;
        RECT 49.145 165.730 49.285 169.490 ;
        RECT 49.605 168.110 49.745 170.170 ;
        RECT 49.545 167.790 49.805 168.110 ;
        RECT 49.085 165.410 49.345 165.730 ;
        RECT 49.085 164.790 49.345 165.050 ;
        RECT 49.605 164.790 49.745 167.790 ;
        RECT 50.525 167.090 50.665 170.510 ;
        RECT 52.760 168.955 54.300 169.325 ;
        RECT 57.425 168.450 57.565 173.230 ;
        RECT 59.725 173.210 59.865 186.830 ;
        RECT 61.505 184.790 61.765 185.110 ;
        RECT 60.125 183.090 60.385 183.410 ;
        RECT 60.185 181.280 60.325 183.090 ;
        RECT 60.585 181.280 60.845 181.370 ;
        RECT 60.185 181.140 60.845 181.280 ;
        RECT 60.185 178.650 60.325 181.140 ;
        RECT 60.585 181.050 60.845 181.140 ;
        RECT 61.565 181.030 61.705 184.790 ;
        RECT 66.105 184.000 66.365 184.090 ;
        RECT 66.105 183.860 66.765 184.000 ;
        RECT 66.105 183.770 66.365 183.860 ;
        RECT 63.805 183.090 64.065 183.410 ;
        RECT 63.865 182.390 64.005 183.090 ;
        RECT 64.550 182.555 66.090 182.925 ;
        RECT 63.805 182.070 64.065 182.390 ;
        RECT 65.645 181.730 65.905 182.050 ;
        RECT 61.505 180.710 61.765 181.030 ;
        RECT 60.585 180.370 60.845 180.690 ;
        RECT 60.125 178.330 60.385 178.650 ;
        RECT 59.665 172.890 59.925 173.210 ;
        RECT 58.745 172.550 59.005 172.870 ;
        RECT 58.805 171.510 58.945 172.550 ;
        RECT 58.745 171.190 59.005 171.510 ;
        RECT 57.365 168.130 57.625 168.450 ;
        RECT 50.465 166.770 50.725 167.090 ;
        RECT 56.905 166.770 57.165 167.090 ;
        RECT 50.525 165.050 50.665 166.770 ;
        RECT 56.965 165.390 57.105 166.770 ;
        RECT 50.925 165.070 51.185 165.390 ;
        RECT 56.905 165.070 57.165 165.390 ;
        RECT 57.425 165.300 57.565 168.130 ;
        RECT 57.825 165.300 58.085 165.390 ;
        RECT 57.425 165.160 58.085 165.300 ;
        RECT 49.085 164.730 49.745 164.790 ;
        RECT 50.465 164.730 50.725 165.050 ;
        RECT 49.145 164.650 49.745 164.730 ;
        RECT 48.625 161.330 48.885 161.650 ;
        RECT 48.685 159.950 48.825 161.330 ;
        RECT 48.625 159.630 48.885 159.950 ;
        RECT 47.705 158.610 47.965 158.930 ;
        RECT 48.685 157.230 48.825 159.630 ;
        RECT 49.145 159.610 49.285 164.650 ;
        RECT 49.085 159.290 49.345 159.610 ;
        RECT 48.625 156.910 48.885 157.230 ;
        RECT 49.545 156.570 49.805 156.890 ;
        RECT 49.605 156.210 49.745 156.570 ;
        RECT 49.545 155.890 49.805 156.210 ;
        RECT 49.605 154.510 49.745 155.890 ;
        RECT 50.525 154.510 50.665 164.730 ;
        RECT 50.985 161.650 51.125 165.070 ;
        RECT 52.760 163.515 54.300 163.885 ;
        RECT 52.305 163.030 52.565 163.350 ;
        RECT 50.925 161.330 51.185 161.650 ;
        RECT 52.365 160.630 52.505 163.030 ;
        RECT 57.425 162.670 57.565 165.160 ;
        RECT 57.825 165.070 58.085 165.160 ;
        RECT 60.125 165.070 60.385 165.390 ;
        RECT 59.205 164.280 59.465 164.370 ;
        RECT 58.805 164.140 59.465 164.280 ;
        RECT 57.365 162.350 57.625 162.670 ;
        RECT 52.765 161.330 53.025 161.650 ;
        RECT 52.305 160.310 52.565 160.630 ;
        RECT 52.825 159.950 52.965 161.330 ;
        RECT 54.605 160.310 54.865 160.630 ;
        RECT 52.305 159.630 52.565 159.950 ;
        RECT 52.765 159.630 53.025 159.950 ;
        RECT 52.365 157.910 52.505 159.630 ;
        RECT 54.665 159.270 54.805 160.310 ;
        RECT 55.065 159.630 55.325 159.950 ;
        RECT 54.605 158.950 54.865 159.270 ;
        RECT 52.760 158.075 54.300 158.445 ;
        RECT 52.305 157.590 52.565 157.910 ;
        RECT 49.545 154.190 49.805 154.510 ;
        RECT 50.465 154.190 50.725 154.510 ;
        RECT 47.245 153.850 47.505 154.170 ;
        RECT 51.845 153.850 52.105 154.170 ;
        RECT 52.365 154.025 52.505 157.590 ;
        RECT 52.765 156.745 53.025 156.890 ;
        RECT 52.755 156.375 53.035 156.745 ;
        RECT 47.245 153.170 47.505 153.490 ;
        RECT 46.785 151.130 47.045 151.450 ;
        RECT 46.845 149.150 46.985 151.130 ;
        RECT 45.925 149.070 46.985 149.150 ;
        RECT 45.405 148.750 45.665 149.070 ;
        RECT 45.865 149.010 46.985 149.070 ;
        RECT 45.865 148.750 46.125 149.010 ;
        RECT 45.465 148.390 45.605 148.750 ;
        RECT 45.405 148.070 45.665 148.390 ;
        RECT 45.465 146.010 45.605 148.070 ;
        RECT 46.845 146.010 46.985 149.010 ;
        RECT 45.405 145.690 45.665 146.010 ;
        RECT 45.465 143.540 45.605 145.690 ;
        RECT 46.315 145.495 46.595 145.865 ;
        RECT 46.785 145.690 47.045 146.010 ;
        RECT 45.865 143.540 46.125 143.630 ;
        RECT 45.465 143.400 46.125 143.540 ;
        RECT 45.865 143.310 46.125 143.400 ;
        RECT 46.385 143.030 46.525 145.495 ;
        RECT 46.845 144.310 46.985 145.690 ;
        RECT 46.785 143.990 47.045 144.310 ;
        RECT 46.845 143.630 46.985 143.990 ;
        RECT 46.785 143.310 47.045 143.630 ;
        RECT 45.465 142.890 46.525 143.030 ;
        RECT 45.465 141.250 45.605 142.890 ;
        RECT 46.775 142.775 47.055 143.145 ;
        RECT 45.865 142.290 46.125 142.610 ;
        RECT 46.325 142.290 46.585 142.610 ;
        RECT 45.405 140.930 45.665 141.250 ;
        RECT 45.465 137.510 45.605 140.930 ;
        RECT 45.925 140.570 46.065 142.290 ;
        RECT 45.865 140.250 46.125 140.570 ;
        RECT 45.925 137.510 46.065 140.250 ;
        RECT 45.405 137.190 45.665 137.510 ;
        RECT 45.865 137.190 46.125 137.510 ;
        RECT 45.465 135.810 45.605 137.190 ;
        RECT 45.405 135.490 45.665 135.810 ;
        RECT 44.945 134.130 45.205 134.450 ;
        RECT 44.945 132.660 45.205 132.750 ;
        RECT 45.465 132.660 45.605 135.490 ;
        RECT 45.925 135.130 46.065 137.190 ;
        RECT 45.865 134.810 46.125 135.130 ;
        RECT 45.865 134.130 46.125 134.450 ;
        RECT 44.945 132.520 45.605 132.660 ;
        RECT 44.945 132.430 45.205 132.520 ;
        RECT 44.945 131.410 45.205 131.730 ;
        RECT 45.405 131.410 45.665 131.730 ;
        RECT 45.005 130.110 45.145 131.410 ;
        RECT 45.465 130.710 45.605 131.410 ;
        RECT 45.405 130.390 45.665 130.710 ;
        RECT 45.005 129.970 45.605 130.110 ;
        RECT 44.945 128.690 45.205 129.010 ;
        RECT 44.485 124.950 44.745 125.270 ;
        RECT 44.485 123.930 44.745 124.250 ;
        RECT 44.025 121.890 44.285 122.210 ;
        RECT 44.545 121.870 44.685 123.930 ;
        RECT 44.485 121.550 44.745 121.870 ;
        RECT 44.025 118.720 44.285 118.810 ;
        RECT 44.545 118.720 44.685 121.550 ;
        RECT 44.025 118.580 44.685 118.720 ;
        RECT 44.025 118.490 44.285 118.580 ;
        RECT 44.025 117.810 44.285 118.130 ;
        RECT 44.085 117.110 44.225 117.810 ;
        RECT 44.025 116.790 44.285 117.110 ;
        RECT 43.565 113.050 43.825 113.370 ;
        RECT 45.005 107.930 45.145 128.690 ;
        RECT 45.465 127.310 45.605 129.970 ;
        RECT 45.925 129.690 46.065 134.130 ;
        RECT 45.865 129.370 46.125 129.690 ;
        RECT 45.405 126.990 45.665 127.310 ;
        RECT 45.855 127.135 46.135 127.505 ;
        RECT 46.385 127.310 46.525 142.290 ;
        RECT 46.845 140.230 46.985 142.775 ;
        RECT 47.305 140.425 47.445 153.170 ;
        RECT 51.905 152.470 52.045 153.850 ;
        RECT 52.295 153.655 52.575 154.025 ;
        RECT 54.605 153.170 54.865 153.490 ;
        RECT 52.760 152.635 54.300 153.005 ;
        RECT 51.845 152.150 52.105 152.470 ;
        RECT 47.705 151.130 47.965 151.450 ;
        RECT 47.765 148.730 47.905 151.130 ;
        RECT 48.165 150.790 48.425 151.110 ;
        RECT 48.225 149.070 48.365 150.790 ;
        RECT 49.085 150.450 49.345 150.770 ;
        RECT 50.925 150.450 51.185 150.770 ;
        RECT 48.165 148.750 48.425 149.070 ;
        RECT 47.705 148.410 47.965 148.730 ;
        RECT 47.695 146.175 47.975 146.545 ;
        RECT 47.705 146.030 47.965 146.175 ;
        RECT 46.785 139.910 47.045 140.230 ;
        RECT 47.235 140.055 47.515 140.425 ;
        RECT 46.845 138.190 46.985 139.910 ;
        RECT 47.765 138.870 47.905 146.030 ;
        RECT 48.225 146.010 48.365 148.750 ;
        RECT 48.625 148.070 48.885 148.390 ;
        RECT 48.165 145.690 48.425 146.010 ;
        RECT 48.165 141.270 48.425 141.590 ;
        RECT 48.225 139.800 48.365 141.270 ;
        RECT 48.685 140.570 48.825 148.070 ;
        RECT 49.145 140.910 49.285 150.450 ;
        RECT 50.985 149.070 51.125 150.450 ;
        RECT 50.005 148.750 50.265 149.070 ;
        RECT 50.465 148.750 50.725 149.070 ;
        RECT 50.925 148.750 51.185 149.070 ;
        RECT 50.065 146.010 50.205 148.750 ;
        RECT 50.525 146.430 50.665 148.750 ;
        RECT 50.525 146.290 51.125 146.430 ;
        RECT 50.005 145.690 50.265 146.010 ;
        RECT 49.545 145.350 49.805 145.670 ;
        RECT 49.605 144.310 49.745 145.350 ;
        RECT 49.545 143.990 49.805 144.310 ;
        RECT 50.065 143.630 50.205 145.690 ;
        RECT 50.525 144.310 50.665 146.290 ;
        RECT 50.985 146.010 51.125 146.290 ;
        RECT 51.905 146.010 52.045 152.150 ;
        RECT 54.665 149.750 54.805 153.170 ;
        RECT 54.605 149.430 54.865 149.750 ;
        RECT 52.305 148.750 52.565 149.070 ;
        RECT 52.365 146.600 52.505 148.750 ;
        RECT 52.760 147.195 54.300 147.565 ;
        RECT 54.665 146.690 54.805 149.430 ;
        RECT 55.125 148.110 55.265 159.630 ;
        RECT 56.905 158.610 57.165 158.930 ;
        RECT 56.965 156.210 57.105 158.610 ;
        RECT 57.425 156.890 57.565 162.350 ;
        RECT 58.285 161.670 58.545 161.990 ;
        RECT 58.345 156.890 58.485 161.670 ;
        RECT 57.365 156.800 57.625 156.890 ;
        RECT 57.365 156.660 58.025 156.800 ;
        RECT 57.365 156.570 57.625 156.660 ;
        RECT 56.905 155.890 57.165 156.210 ;
        RECT 57.885 154.170 58.025 156.660 ;
        RECT 58.285 156.570 58.545 156.890 ;
        RECT 58.805 154.850 58.945 164.140 ;
        RECT 59.205 164.050 59.465 164.140 ;
        RECT 59.665 156.570 59.925 156.890 ;
        RECT 58.745 154.530 59.005 154.850 ;
        RECT 57.825 153.850 58.085 154.170 ;
        RECT 57.885 151.450 58.025 153.850 ;
        RECT 57.825 151.130 58.085 151.450 ;
        RECT 59.725 151.110 59.865 156.570 ;
        RECT 60.185 151.985 60.325 165.070 ;
        RECT 60.645 159.950 60.785 180.370 ;
        RECT 61.565 178.990 61.705 180.710 ;
        RECT 65.185 180.370 65.445 180.690 ;
        RECT 62.885 179.350 63.145 179.670 ;
        RECT 61.505 178.670 61.765 178.990 ;
        RECT 61.565 175.250 61.705 178.670 ;
        RECT 61.505 174.930 61.765 175.250 ;
        RECT 62.945 173.890 63.085 179.350 ;
        RECT 63.805 179.010 64.065 179.330 ;
        RECT 63.865 178.650 64.005 179.010 ;
        RECT 63.805 178.330 64.065 178.650 ;
        RECT 65.245 178.505 65.385 180.370 ;
        RECT 65.705 178.990 65.845 181.730 ;
        RECT 66.625 181.030 66.765 183.860 ;
        RECT 68.925 183.750 69.065 188.530 ;
        RECT 88.125 187.995 89.665 188.365 ;
        RECT 70.245 186.830 70.505 187.150 ;
        RECT 92.325 186.830 92.585 187.150 ;
        RECT 69.325 186.490 69.585 186.810 ;
        RECT 68.865 183.430 69.125 183.750 ;
        RECT 68.405 182.070 68.665 182.390 ;
        RECT 67.945 181.110 68.205 181.370 ;
        RECT 67.085 181.050 68.205 181.110 ;
        RECT 66.565 180.710 66.825 181.030 ;
        RECT 67.085 180.970 68.145 181.050 ;
        RECT 67.085 179.670 67.225 180.970 ;
        RECT 66.105 179.350 66.365 179.670 ;
        RECT 67.025 179.350 67.285 179.670 ;
        RECT 66.165 178.990 66.305 179.350 ;
        RECT 65.645 178.670 65.905 178.990 ;
        RECT 66.105 178.670 66.365 178.990 ;
        RECT 67.025 178.670 67.285 178.990 ;
        RECT 65.175 178.135 65.455 178.505 ;
        RECT 66.565 177.650 66.825 177.970 ;
        RECT 64.550 177.115 66.090 177.485 ;
        RECT 65.645 176.630 65.905 176.950 ;
        RECT 65.705 176.270 65.845 176.630 ;
        RECT 66.625 176.610 66.765 177.650 ;
        RECT 67.085 176.950 67.225 178.670 ;
        RECT 67.025 176.630 67.285 176.950 ;
        RECT 66.565 176.290 66.825 176.610 ;
        RECT 65.645 175.950 65.905 176.270 ;
        RECT 67.025 175.610 67.285 175.930 ;
        RECT 67.085 174.230 67.225 175.610 ;
        RECT 68.005 174.230 68.145 180.970 ;
        RECT 68.465 177.970 68.605 182.070 ;
        RECT 69.385 182.050 69.525 186.490 ;
        RECT 70.305 185.110 70.445 186.830 ;
        RECT 73.925 186.150 74.185 186.470 ;
        RECT 70.245 184.790 70.505 185.110 ;
        RECT 73.985 184.430 74.125 186.150 ;
        RECT 80.825 185.810 81.085 186.130 ;
        RECT 76.335 185.275 77.875 185.645 ;
        RECT 80.885 184.430 81.025 185.810 ;
        RECT 92.385 184.430 92.525 186.830 ;
        RECT 93.705 185.810 93.965 186.130 ;
        RECT 96.005 185.810 96.265 186.130 ;
        RECT 73.925 184.110 74.185 184.430 ;
        RECT 80.825 184.110 81.085 184.430 ;
        RECT 92.325 184.110 92.585 184.430 ;
        RECT 74.385 183.770 74.645 184.090 ;
        RECT 81.745 183.770 82.005 184.090 ;
        RECT 74.445 182.300 74.585 183.770 ;
        RECT 78.985 183.090 79.245 183.410 ;
        RECT 79.445 183.090 79.705 183.410 ;
        RECT 73.985 182.160 74.585 182.300 ;
        RECT 69.325 181.730 69.585 182.050 ;
        RECT 69.385 179.670 69.525 181.730 ;
        RECT 73.985 181.710 74.125 182.160 ;
        RECT 79.045 182.050 79.185 183.090 ;
        RECT 78.985 181.730 79.245 182.050 ;
        RECT 72.085 181.390 72.345 181.710 ;
        RECT 73.925 181.390 74.185 181.710 ;
        RECT 74.385 181.390 74.645 181.710 ;
        RECT 70.245 181.050 70.505 181.370 ;
        RECT 69.325 179.350 69.585 179.670 ;
        RECT 70.305 178.650 70.445 181.050 ;
        RECT 72.145 178.990 72.285 181.390 ;
        RECT 72.085 178.670 72.345 178.990 ;
        RECT 70.245 178.330 70.505 178.650 ;
        RECT 68.405 177.650 68.665 177.970 ;
        RECT 68.465 176.950 68.605 177.650 ;
        RECT 68.405 176.630 68.665 176.950 ;
        RECT 70.245 176.290 70.505 176.610 ;
        RECT 63.805 173.910 64.065 174.230 ;
        RECT 67.025 173.910 67.285 174.230 ;
        RECT 67.945 173.910 68.205 174.230 ;
        RECT 62.885 173.570 63.145 173.890 ;
        RECT 63.345 172.890 63.605 173.210 ;
        RECT 62.885 172.210 63.145 172.530 ;
        RECT 62.945 171.170 63.085 172.210 ;
        RECT 63.405 171.510 63.545 172.890 ;
        RECT 63.345 171.190 63.605 171.510 ;
        RECT 62.885 170.850 63.145 171.170 ;
        RECT 63.865 169.810 64.005 173.910 ;
        RECT 68.005 173.550 68.145 173.910 ;
        RECT 67.945 173.230 68.205 173.550 ;
        RECT 66.565 172.210 66.825 172.530 ;
        RECT 64.550 171.675 66.090 172.045 ;
        RECT 66.625 171.170 66.765 172.210 ;
        RECT 66.565 170.850 66.825 171.170 ;
        RECT 63.805 169.490 64.065 169.810 ;
        RECT 61.045 167.450 61.305 167.770 ;
        RECT 61.105 165.390 61.245 167.450 ;
        RECT 63.865 165.390 64.005 169.490 ;
        RECT 64.550 166.235 66.090 166.605 ;
        RECT 67.485 165.750 67.745 166.070 ;
        RECT 61.045 165.070 61.305 165.390 ;
        RECT 63.805 165.070 64.065 165.390 ;
        RECT 62.425 164.730 62.685 165.050 ;
        RECT 62.485 162.670 62.625 164.730 ;
        RECT 66.565 164.390 66.825 164.710 ;
        RECT 63.805 164.050 64.065 164.370 ;
        RECT 62.425 162.350 62.685 162.670 ;
        RECT 61.045 161.330 61.305 161.650 ;
        RECT 63.345 161.330 63.605 161.650 ;
        RECT 60.585 159.630 60.845 159.950 ;
        RECT 61.105 156.890 61.245 161.330 ;
        RECT 63.405 159.950 63.545 161.330 ;
        RECT 63.865 160.540 64.005 164.050 ;
        RECT 64.550 160.795 66.090 161.165 ;
        RECT 63.865 160.400 64.465 160.540 ;
        RECT 61.505 159.630 61.765 159.950 ;
        RECT 61.965 159.630 62.225 159.950 ;
        RECT 63.345 159.630 63.605 159.950 ;
        RECT 61.565 157.230 61.705 159.630 ;
        RECT 62.025 159.465 62.165 159.630 ;
        RECT 61.955 159.095 62.235 159.465 ;
        RECT 64.325 159.350 64.465 160.400 ;
        RECT 66.625 159.950 66.765 164.390 ;
        RECT 67.545 162.330 67.685 165.750 ;
        RECT 68.005 165.390 68.145 173.230 ;
        RECT 70.305 173.210 70.445 176.290 ;
        RECT 71.165 174.930 71.425 175.250 ;
        RECT 71.225 173.210 71.365 174.930 ;
        RECT 68.405 172.890 68.665 173.210 ;
        RECT 70.245 173.120 70.505 173.210 ;
        RECT 69.845 172.980 70.505 173.120 ;
        RECT 68.465 172.530 68.605 172.890 ;
        RECT 68.405 172.210 68.665 172.530 ;
        RECT 68.865 170.510 69.125 170.830 ;
        RECT 68.925 167.770 69.065 170.510 ;
        RECT 68.865 167.450 69.125 167.770 ;
        RECT 68.405 165.750 68.665 166.070 ;
        RECT 68.465 165.390 68.605 165.750 ;
        RECT 69.845 165.390 69.985 172.980 ;
        RECT 70.245 172.890 70.505 172.980 ;
        RECT 71.165 173.120 71.425 173.210 ;
        RECT 71.165 172.980 71.825 173.120 ;
        RECT 71.165 172.890 71.425 172.980 ;
        RECT 70.245 170.170 70.505 170.490 ;
        RECT 67.945 165.070 68.205 165.390 ;
        RECT 68.405 165.070 68.665 165.390 ;
        RECT 69.785 165.070 70.045 165.390 ;
        RECT 68.005 162.670 68.145 165.070 ;
        RECT 68.405 164.390 68.665 164.710 ;
        RECT 68.465 163.010 68.605 164.390 ;
        RECT 70.305 163.010 70.445 170.170 ;
        RECT 71.165 166.770 71.425 167.090 ;
        RECT 70.705 165.410 70.965 165.730 ;
        RECT 68.405 162.690 68.665 163.010 ;
        RECT 70.245 162.690 70.505 163.010 ;
        RECT 67.945 162.350 68.205 162.670 ;
        RECT 67.485 162.010 67.745 162.330 ;
        RECT 67.025 161.670 67.285 161.990 ;
        RECT 67.085 159.950 67.225 161.670 ;
        RECT 67.545 159.950 67.685 162.010 ;
        RECT 68.005 159.950 68.145 162.350 ;
        RECT 68.465 159.950 68.605 162.690 ;
        RECT 69.325 162.010 69.585 162.330 ;
        RECT 64.725 159.630 64.985 159.950 ;
        RECT 66.565 159.630 66.825 159.950 ;
        RECT 67.025 159.630 67.285 159.950 ;
        RECT 67.485 159.630 67.745 159.950 ;
        RECT 67.945 159.630 68.205 159.950 ;
        RECT 68.405 159.630 68.665 159.950 ;
        RECT 61.505 156.910 61.765 157.230 ;
        RECT 61.045 156.570 61.305 156.890 ;
        RECT 61.495 156.375 61.775 156.745 ;
        RECT 61.565 156.210 61.705 156.375 ;
        RECT 61.505 155.890 61.765 156.210 ;
        RECT 61.565 154.705 61.705 155.890 ;
        RECT 60.585 154.190 60.845 154.510 ;
        RECT 61.495 154.335 61.775 154.705 ;
        RECT 62.025 154.510 62.165 159.095 ;
        RECT 62.885 158.950 63.145 159.270 ;
        RECT 63.345 158.950 63.605 159.270 ;
        RECT 63.865 159.210 64.465 159.350 ;
        RECT 62.425 156.570 62.685 156.890 ;
        RECT 62.485 154.850 62.625 156.570 ;
        RECT 62.425 154.530 62.685 154.850 ;
        RECT 61.965 154.190 62.225 154.510 ;
        RECT 60.645 152.470 60.785 154.190 ;
        RECT 60.585 152.150 60.845 152.470 ;
        RECT 61.505 152.150 61.765 152.470 ;
        RECT 60.115 151.615 60.395 151.985 ;
        RECT 61.565 151.870 61.705 152.150 ;
        RECT 59.665 150.790 59.925 151.110 ;
        RECT 58.745 148.750 59.005 149.070 ;
        RECT 57.365 148.585 57.625 148.730 ;
        RECT 57.355 148.470 57.635 148.585 ;
        RECT 56.965 148.330 57.635 148.470 ;
        RECT 55.125 147.970 56.185 148.110 ;
        RECT 52.365 146.460 53.425 146.600 ;
        RECT 50.925 145.690 51.185 146.010 ;
        RECT 51.845 145.690 52.105 146.010 ;
        RECT 52.765 145.690 53.025 146.010 ;
        RECT 50.465 143.990 50.725 144.310 ;
        RECT 50.525 143.630 50.665 143.990 ;
        RECT 52.825 143.970 52.965 145.690 ;
        RECT 53.285 145.330 53.425 146.460 ;
        RECT 54.605 146.370 54.865 146.690 ;
        RECT 53.225 145.010 53.485 145.330 ;
        RECT 55.525 145.010 55.785 145.330 ;
        RECT 52.765 143.650 53.025 143.970 ;
        RECT 53.285 143.630 53.425 145.010 ;
        RECT 55.585 143.630 55.725 145.010 ;
        RECT 50.005 143.310 50.265 143.630 ;
        RECT 50.465 143.310 50.725 143.630 ;
        RECT 53.225 143.310 53.485 143.630 ;
        RECT 55.525 143.310 55.785 143.630 ;
        RECT 51.845 142.465 52.105 142.610 ;
        RECT 51.835 142.095 52.115 142.465 ;
        RECT 52.760 141.755 54.300 142.125 ;
        RECT 55.585 141.590 55.725 143.310 ;
        RECT 55.065 141.270 55.325 141.590 ;
        RECT 55.525 141.270 55.785 141.590 ;
        RECT 49.085 140.590 49.345 140.910 ;
        RECT 49.545 140.590 49.805 140.910 ;
        RECT 49.995 140.735 50.275 141.105 ;
        RECT 55.125 140.990 55.265 141.270 ;
        RECT 56.045 140.990 56.185 147.970 ;
        RECT 56.965 146.350 57.105 148.330 ;
        RECT 57.355 148.215 57.635 148.330 ;
        RECT 56.905 146.030 57.165 146.350 ;
        RECT 56.965 144.310 57.105 146.030 ;
        RECT 57.825 145.010 58.085 145.330 ;
        RECT 56.905 143.990 57.165 144.310 ;
        RECT 56.435 143.455 56.715 143.825 ;
        RECT 56.445 143.310 56.705 143.455 ;
        RECT 55.125 140.850 56.185 140.990 ;
        RECT 48.625 140.250 48.885 140.570 ;
        RECT 48.225 139.660 48.825 139.800 ;
        RECT 47.705 138.550 47.965 138.870 ;
        RECT 47.245 138.210 47.505 138.530 ;
        RECT 46.785 137.870 47.045 138.190 ;
        RECT 47.305 137.850 47.445 138.210 ;
        RECT 47.705 137.870 47.965 138.190 ;
        RECT 47.245 137.530 47.505 137.850 ;
        RECT 46.785 136.850 47.045 137.170 ;
        RECT 46.845 130.030 46.985 136.850 ;
        RECT 47.765 136.150 47.905 137.870 ;
        RECT 48.165 137.025 48.425 137.170 ;
        RECT 48.155 136.655 48.435 137.025 ;
        RECT 47.705 135.830 47.965 136.150 ;
        RECT 47.765 135.130 47.905 135.830 ;
        RECT 47.705 134.870 47.965 135.130 ;
        RECT 47.305 134.810 47.965 134.870 ;
        RECT 47.305 134.730 47.905 134.810 ;
        RECT 47.305 132.410 47.445 134.730 ;
        RECT 47.705 134.130 47.965 134.450 ;
        RECT 48.685 134.360 48.825 139.660 ;
        RECT 49.605 137.510 49.745 140.590 ;
        RECT 50.065 140.570 50.205 140.735 ;
        RECT 50.005 140.250 50.265 140.570 ;
        RECT 50.005 139.570 50.265 139.890 ;
        RECT 53.685 139.570 53.945 139.890 ;
        RECT 49.545 137.190 49.805 137.510 ;
        RECT 49.075 135.295 49.355 135.665 ;
        RECT 49.145 135.130 49.285 135.295 ;
        RECT 49.605 135.130 49.745 137.190 ;
        RECT 49.085 134.810 49.345 135.130 ;
        RECT 49.545 134.810 49.805 135.130 ;
        RECT 48.685 134.220 49.285 134.360 ;
        RECT 47.245 132.090 47.505 132.410 ;
        RECT 47.245 130.050 47.505 130.370 ;
        RECT 46.785 129.710 47.045 130.030 ;
        RECT 45.865 126.990 46.125 127.135 ;
        RECT 46.325 126.990 46.585 127.310 ;
        RECT 45.865 126.310 46.125 126.630 ;
        RECT 46.325 126.310 46.585 126.630 ;
        RECT 45.405 125.970 45.665 126.290 ;
        RECT 45.465 107.930 45.605 125.970 ;
        RECT 45.925 124.250 46.065 126.310 ;
        RECT 46.385 124.590 46.525 126.310 ;
        RECT 46.785 125.970 47.045 126.290 ;
        RECT 46.845 125.270 46.985 125.970 ;
        RECT 46.785 124.950 47.045 125.270 ;
        RECT 46.325 124.270 46.585 124.590 ;
        RECT 45.865 123.930 46.125 124.250 ;
        RECT 45.925 118.130 46.065 123.930 ;
        RECT 46.325 123.590 46.585 123.910 ;
        RECT 46.385 122.550 46.525 123.590 ;
        RECT 46.325 122.230 46.585 122.550 ;
        RECT 46.785 120.760 47.045 120.850 ;
        RECT 47.305 120.760 47.445 130.050 ;
        RECT 47.765 129.010 47.905 134.130 ;
        RECT 48.165 132.770 48.425 133.090 ;
        RECT 48.225 130.225 48.365 132.770 ;
        RECT 49.145 130.620 49.285 134.220 ;
        RECT 49.545 132.090 49.805 132.410 ;
        RECT 48.685 130.480 49.285 130.620 ;
        RECT 48.155 129.855 48.435 130.225 ;
        RECT 47.705 128.690 47.965 129.010 ;
        RECT 47.705 126.650 47.965 126.970 ;
        RECT 47.765 124.250 47.905 126.650 ;
        RECT 47.705 124.105 47.965 124.250 ;
        RECT 47.695 123.735 47.975 124.105 ;
        RECT 46.785 120.620 47.445 120.760 ;
        RECT 46.785 120.530 47.045 120.620 ;
        RECT 48.685 119.830 48.825 130.480 ;
        RECT 49.605 129.690 49.745 132.090 ;
        RECT 49.075 129.175 49.355 129.545 ;
        RECT 49.545 129.370 49.805 129.690 ;
        RECT 49.085 129.030 49.345 129.175 ;
        RECT 49.545 126.650 49.805 126.970 ;
        RECT 49.605 124.590 49.745 126.650 ;
        RECT 49.545 124.270 49.805 124.590 ;
        RECT 49.085 123.250 49.345 123.570 ;
        RECT 49.145 121.870 49.285 123.250 ;
        RECT 49.085 121.550 49.345 121.870 ;
        RECT 48.625 119.510 48.885 119.830 ;
        RECT 46.325 118.830 46.585 119.150 ;
        RECT 49.085 119.060 49.345 119.150 ;
        RECT 49.605 119.060 49.745 124.270 ;
        RECT 49.085 118.920 49.745 119.060 ;
        RECT 49.085 118.830 49.345 118.920 ;
        RECT 45.865 117.810 46.125 118.130 ;
        RECT 46.385 116.090 46.525 118.830 ;
        RECT 48.625 118.150 48.885 118.470 ;
        RECT 46.785 117.810 47.045 118.130 ;
        RECT 45.865 115.770 46.125 116.090 ;
        RECT 46.325 115.770 46.585 116.090 ;
        RECT 45.925 114.390 46.065 115.770 ;
        RECT 45.865 114.070 46.125 114.390 ;
        RECT 46.845 113.370 46.985 117.810 ;
        RECT 48.685 117.110 48.825 118.150 ;
        RECT 48.625 116.790 48.885 117.110 ;
        RECT 47.705 116.450 47.965 116.770 ;
        RECT 47.765 113.370 47.905 116.450 ;
        RECT 46.785 113.050 47.045 113.370 ;
        RECT 47.245 113.050 47.505 113.370 ;
        RECT 47.705 113.050 47.965 113.370 ;
        RECT 47.305 112.690 47.445 113.050 ;
        RECT 47.245 112.370 47.505 112.690 ;
        RECT 47.305 111.330 47.445 112.370 ;
        RECT 47.245 111.010 47.505 111.330 ;
        RECT 50.065 108.610 50.205 139.570 ;
        RECT 50.465 137.870 50.725 138.190 ;
        RECT 52.305 137.870 52.565 138.190 ;
        RECT 50.525 135.810 50.665 137.870 ;
        RECT 51.375 137.335 51.655 137.705 ;
        RECT 50.465 135.490 50.725 135.810 ;
        RECT 51.445 135.470 51.585 137.335 ;
        RECT 51.845 137.190 52.105 137.510 ;
        RECT 51.385 135.150 51.645 135.470 ;
        RECT 51.905 135.130 52.045 137.190 ;
        RECT 50.925 134.810 51.185 135.130 ;
        RECT 51.845 134.810 52.105 135.130 ;
        RECT 52.365 135.040 52.505 137.870 ;
        RECT 53.745 137.850 53.885 139.570 ;
        RECT 55.525 138.210 55.785 138.530 ;
        RECT 53.685 137.530 53.945 137.850 ;
        RECT 54.605 136.850 54.865 137.170 ;
        RECT 55.065 136.850 55.325 137.170 ;
        RECT 52.760 136.315 54.300 136.685 ;
        RECT 53.685 135.490 53.945 135.810 ;
        RECT 53.225 135.040 53.485 135.130 ;
        RECT 52.365 134.900 53.485 135.040 ;
        RECT 50.465 134.130 50.725 134.450 ;
        RECT 50.525 132.070 50.665 134.130 ;
        RECT 50.985 132.750 51.125 134.810 ;
        RECT 51.905 134.310 52.045 134.810 ;
        RECT 51.905 134.170 52.505 134.310 ;
        RECT 51.385 132.770 51.645 133.090 ;
        RECT 50.925 132.430 51.185 132.750 ;
        RECT 50.465 131.750 50.725 132.070 ;
        RECT 50.925 131.750 51.185 132.070 ;
        RECT 50.985 130.030 51.125 131.750 ;
        RECT 50.925 129.710 51.185 130.030 ;
        RECT 51.445 129.690 51.585 132.770 ;
        RECT 52.365 132.410 52.505 134.170 ;
        RECT 52.825 133.090 52.965 134.900 ;
        RECT 53.225 134.810 53.485 134.900 ;
        RECT 52.765 132.770 53.025 133.090 ;
        RECT 53.745 132.750 53.885 135.490 ;
        RECT 54.145 135.380 54.405 135.470 ;
        RECT 54.665 135.380 54.805 136.850 ;
        RECT 55.125 135.810 55.265 136.850 ;
        RECT 55.585 136.150 55.725 138.210 ;
        RECT 55.525 135.830 55.785 136.150 ;
        RECT 55.065 135.490 55.325 135.810 ;
        RECT 54.145 135.240 54.805 135.380 ;
        RECT 54.145 135.150 54.405 135.240 ;
        RECT 54.205 134.305 54.345 135.150 ;
        RECT 55.065 134.870 55.325 135.130 ;
        RECT 55.515 134.870 55.795 134.985 ;
        RECT 56.045 134.870 56.185 140.850 ;
        RECT 55.065 134.810 56.185 134.870 ;
        RECT 55.125 134.730 56.185 134.810 ;
        RECT 55.515 134.615 55.795 134.730 ;
        RECT 54.135 133.935 54.415 134.305 ;
        RECT 56.505 132.830 56.645 143.310 ;
        RECT 56.965 135.470 57.105 143.990 ;
        RECT 57.885 139.890 58.025 145.010 ;
        RECT 58.805 143.970 58.945 148.750 ;
        RECT 60.185 148.730 60.325 151.615 ;
        RECT 60.585 151.470 60.845 151.790 ;
        RECT 61.105 151.730 61.705 151.870 ;
        RECT 60.645 149.750 60.785 151.470 ;
        RECT 60.585 149.430 60.845 149.750 ;
        RECT 61.105 149.150 61.245 151.730 ;
        RECT 61.965 151.130 62.225 151.450 ;
        RECT 61.505 149.430 61.765 149.750 ;
        RECT 60.645 149.010 61.245 149.150 ;
        RECT 60.125 148.410 60.385 148.730 ;
        RECT 60.645 145.670 60.785 149.010 ;
        RECT 60.585 145.350 60.845 145.670 ;
        RECT 61.045 145.010 61.305 145.330 ;
        RECT 58.745 143.650 59.005 143.970 ;
        RECT 57.825 139.570 58.085 139.890 ;
        RECT 56.905 135.380 57.165 135.470 ;
        RECT 56.905 135.240 57.565 135.380 ;
        RECT 56.905 135.150 57.165 135.240 ;
        RECT 53.685 132.660 53.945 132.750 ;
        RECT 53.685 132.520 54.805 132.660 ;
        RECT 53.685 132.430 53.945 132.520 ;
        RECT 52.305 132.090 52.565 132.410 ;
        RECT 52.365 130.710 52.505 132.090 ;
        RECT 52.760 130.875 54.300 131.245 ;
        RECT 52.305 130.390 52.565 130.710 ;
        RECT 50.465 129.370 50.725 129.690 ;
        RECT 51.385 129.370 51.645 129.690 ;
        RECT 52.365 129.430 52.505 130.390 ;
        RECT 54.665 130.030 54.805 132.520 ;
        RECT 55.065 132.430 55.325 132.750 ;
        RECT 56.045 132.690 56.645 132.830 ;
        RECT 54.605 129.710 54.865 130.030 ;
        RECT 55.125 129.690 55.265 132.430 ;
        RECT 50.525 127.990 50.665 129.370 ;
        RECT 51.905 129.290 52.505 129.430 ;
        RECT 53.685 129.370 53.945 129.690 ;
        RECT 55.065 129.370 55.325 129.690 ;
        RECT 50.465 127.670 50.725 127.990 ;
        RECT 51.905 127.650 52.045 129.290 ;
        RECT 50.925 127.330 51.185 127.650 ;
        RECT 51.845 127.330 52.105 127.650 ;
        RECT 50.985 125.270 51.125 127.330 ;
        RECT 53.745 127.310 53.885 129.370 ;
        RECT 55.125 127.310 55.265 129.370 ;
        RECT 53.685 126.990 53.945 127.310 ;
        RECT 55.065 126.990 55.325 127.310 ;
        RECT 52.760 125.435 54.300 125.805 ;
        RECT 50.925 124.950 51.185 125.270 ;
        RECT 56.045 124.785 56.185 132.690 ;
        RECT 56.445 132.320 56.705 132.410 ;
        RECT 57.425 132.320 57.565 135.240 ;
        RECT 57.885 135.130 58.025 139.570 ;
        RECT 57.825 134.810 58.085 135.130 ;
        RECT 57.825 134.305 58.085 134.450 ;
        RECT 57.815 133.935 58.095 134.305 ;
        RECT 57.885 133.430 58.025 133.935 ;
        RECT 57.825 133.110 58.085 133.430 ;
        RECT 56.445 132.180 57.565 132.320 ;
        RECT 56.445 132.090 56.705 132.180 ;
        RECT 57.425 130.030 57.565 132.180 ;
        RECT 58.285 131.410 58.545 131.730 ;
        RECT 57.365 129.710 57.625 130.030 ;
        RECT 58.345 129.690 58.485 131.410 ;
        RECT 58.805 130.620 58.945 143.650 ;
        RECT 60.125 140.250 60.385 140.570 ;
        RECT 59.205 139.910 59.465 140.230 ;
        RECT 59.265 138.870 59.405 139.910 ;
        RECT 59.205 138.550 59.465 138.870 ;
        RECT 60.185 137.850 60.325 140.250 ;
        RECT 61.105 138.190 61.245 145.010 ;
        RECT 61.565 143.145 61.705 149.430 ;
        RECT 62.025 148.390 62.165 151.130 ;
        RECT 62.485 149.410 62.625 154.530 ;
        RECT 62.945 151.790 63.085 158.950 ;
        RECT 63.405 157.230 63.545 158.950 ;
        RECT 63.345 156.910 63.605 157.230 ;
        RECT 63.345 155.890 63.605 156.210 ;
        RECT 63.405 154.705 63.545 155.890 ;
        RECT 63.335 154.335 63.615 154.705 ;
        RECT 63.405 154.170 63.545 154.335 ;
        RECT 63.345 153.850 63.605 154.170 ;
        RECT 63.405 153.490 63.545 153.850 ;
        RECT 63.345 153.170 63.605 153.490 ;
        RECT 62.885 151.470 63.145 151.790 ;
        RECT 63.335 151.615 63.615 151.985 ;
        RECT 62.425 149.090 62.685 149.410 ;
        RECT 62.945 149.070 63.085 151.470 ;
        RECT 63.405 151.450 63.545 151.615 ;
        RECT 63.345 151.130 63.605 151.450 ;
        RECT 62.885 148.750 63.145 149.070 ;
        RECT 61.965 148.070 62.225 148.390 ;
        RECT 62.425 148.070 62.685 148.390 ;
        RECT 62.485 145.670 62.625 148.070 ;
        RECT 62.425 145.350 62.685 145.670 ;
        RECT 61.495 142.775 61.775 143.145 ;
        RECT 61.565 140.230 61.705 142.775 ;
        RECT 63.345 142.630 63.605 142.950 ;
        RECT 62.885 141.270 63.145 141.590 ;
        RECT 62.425 140.250 62.685 140.570 ;
        RECT 61.505 139.910 61.765 140.230 ;
        RECT 61.045 137.870 61.305 138.190 ;
        RECT 62.485 137.850 62.625 140.250 ;
        RECT 62.945 138.870 63.085 141.270 ;
        RECT 62.885 138.550 63.145 138.870 ;
        RECT 59.665 137.530 59.925 137.850 ;
        RECT 60.125 137.530 60.385 137.850 ;
        RECT 62.425 137.530 62.685 137.850 ;
        RECT 59.725 136.150 59.865 137.530 ;
        RECT 59.665 135.830 59.925 136.150 ;
        RECT 58.805 130.480 59.865 130.620 ;
        RECT 59.205 129.710 59.465 130.030 ;
        RECT 58.285 129.370 58.545 129.690 ;
        RECT 56.895 128.495 57.175 128.865 ;
        RECT 58.285 128.690 58.545 129.010 ;
        RECT 55.975 124.415 56.255 124.785 ;
        RECT 50.925 123.250 51.185 123.570 ;
        RECT 54.605 123.250 54.865 123.570 ;
        RECT 50.985 119.150 51.125 123.250 ;
        RECT 52.760 119.995 54.300 120.365 ;
        RECT 50.925 118.830 51.185 119.150 ;
        RECT 52.295 118.975 52.575 119.345 ;
        RECT 50.985 114.390 51.125 118.830 ;
        RECT 52.365 118.810 52.505 118.975 ;
        RECT 54.665 118.810 54.805 123.250 ;
        RECT 56.045 122.550 56.185 124.415 ;
        RECT 55.985 122.230 56.245 122.550 ;
        RECT 55.065 121.890 55.325 122.210 ;
        RECT 55.125 119.830 55.265 121.890 ;
        RECT 55.985 120.530 56.245 120.850 ;
        RECT 55.065 119.510 55.325 119.830 ;
        RECT 52.305 118.490 52.565 118.810 ;
        RECT 54.605 118.490 54.865 118.810 ;
        RECT 55.065 118.665 55.325 118.810 ;
        RECT 55.055 118.295 55.335 118.665 ;
        RECT 51.845 117.810 52.105 118.130 ;
        RECT 50.925 114.070 51.185 114.390 ;
        RECT 50.925 112.710 51.185 113.030 ;
        RECT 50.985 111.670 51.125 112.710 ;
        RECT 50.925 111.350 51.185 111.670 ;
        RECT 51.905 110.990 52.045 117.810 ;
        RECT 52.305 116.790 52.565 117.110 ;
        RECT 52.365 111.670 52.505 116.790 ;
        RECT 52.760 114.555 54.300 114.925 ;
        RECT 56.045 113.370 56.185 120.530 ;
        RECT 55.985 113.050 56.245 113.370 ;
        RECT 52.305 111.350 52.565 111.670 ;
        RECT 51.845 110.670 52.105 110.990 ;
        RECT 55.525 109.650 55.785 109.970 ;
        RECT 52.760 109.115 54.300 109.485 ;
        RECT 50.005 108.290 50.265 108.610 ;
        RECT 55.585 108.270 55.725 109.650 ;
        RECT 55.525 107.950 55.785 108.270 ;
        RECT 39.425 107.610 39.685 107.930 ;
        RECT 42.645 107.610 42.905 107.930 ;
        RECT 44.945 107.610 45.205 107.930 ;
        RECT 45.405 107.610 45.665 107.930 ;
        RECT 50.005 107.610 50.265 107.930 ;
        RECT 39.485 106.230 39.625 107.610 ;
        RECT 49.085 107.270 49.345 107.590 ;
        RECT 40.345 106.930 40.605 107.250 ;
        RECT 45.865 106.930 46.125 107.250 ;
        RECT 39.425 105.910 39.685 106.230 ;
        RECT 38.045 105.570 38.305 105.890 ;
        RECT 38.505 105.570 38.765 105.890 ;
        RECT 32.985 104.980 33.645 105.120 ;
        RECT 32.985 104.890 33.245 104.980 ;
        RECT 33.505 103.170 33.645 104.980 ;
        RECT 35.285 104.890 35.545 105.210 ;
        RECT 37.125 104.890 37.385 105.210 ;
        RECT 30.745 102.940 31.345 103.080 ;
        RECT 27.465 102.510 27.725 102.830 ;
        RECT 30.745 98.340 30.885 102.940 ;
        RECT 33.445 102.850 33.705 103.170 ;
        RECT 35.345 98.340 35.485 104.890 ;
        RECT 37.185 103.510 37.325 104.890 ;
        RECT 39.485 104.530 39.625 105.910 ;
        RECT 39.425 104.210 39.685 104.530 ;
        RECT 37.125 103.190 37.385 103.510 ;
        RECT 39.885 102.510 40.145 102.830 ;
        RECT 39.945 98.340 40.085 102.510 ;
        RECT 40.405 102.490 40.545 106.930 ;
        RECT 40.975 106.395 42.515 106.765 ;
        RECT 44.485 104.890 44.745 105.210 ;
        RECT 40.345 102.170 40.605 102.490 ;
        RECT 40.975 100.955 42.515 101.325 ;
        RECT 44.545 98.340 44.685 104.890 ;
        RECT 45.925 102.830 46.065 106.930 ;
        RECT 45.865 102.510 46.125 102.830 ;
        RECT 49.145 98.340 49.285 107.270 ;
        RECT 50.065 106.230 50.205 107.610 ;
        RECT 50.005 105.910 50.265 106.230 ;
        RECT 55.985 105.570 56.245 105.890 ;
        RECT 54.605 104.890 54.865 105.210 ;
        RECT 52.760 103.675 54.300 104.045 ;
        RECT 54.665 102.910 54.805 104.890 ;
        RECT 56.045 103.510 56.185 105.570 ;
        RECT 55.985 103.190 56.245 103.510 ;
        RECT 53.745 102.770 54.805 102.910 ;
        RECT 53.745 98.340 53.885 102.770 ;
        RECT 56.965 102.490 57.105 128.495 ;
        RECT 57.825 127.330 58.085 127.650 ;
        RECT 57.365 126.650 57.625 126.970 ;
        RECT 57.425 122.550 57.565 126.650 ;
        RECT 57.365 122.230 57.625 122.550 ;
        RECT 57.425 118.130 57.565 122.230 ;
        RECT 57.885 119.830 58.025 127.330 ;
        RECT 58.345 124.250 58.485 128.690 ;
        RECT 58.745 127.670 59.005 127.990 ;
        RECT 58.805 124.590 58.945 127.670 ;
        RECT 59.265 124.590 59.405 129.710 ;
        RECT 58.745 124.270 59.005 124.590 ;
        RECT 59.205 124.270 59.465 124.590 ;
        RECT 58.285 123.930 58.545 124.250 ;
        RECT 57.825 119.510 58.085 119.830 ;
        RECT 58.805 119.150 58.945 124.270 ;
        RECT 59.265 119.830 59.405 124.270 ;
        RECT 59.725 120.850 59.865 130.480 ;
        RECT 60.185 126.970 60.325 137.530 ;
        RECT 61.955 134.615 62.235 134.985 ;
        RECT 63.405 134.870 63.545 142.630 ;
        RECT 63.865 135.470 64.005 159.210 ;
        RECT 64.785 157.230 64.925 159.630 ;
        RECT 65.185 158.950 65.445 159.270 ;
        RECT 65.635 159.095 65.915 159.465 ;
        RECT 65.645 158.950 65.905 159.095 ;
        RECT 64.725 156.910 64.985 157.230 ;
        RECT 65.245 156.120 65.385 158.950 ;
        RECT 66.625 158.670 66.765 159.630 ;
        RECT 68.855 159.095 69.135 159.465 ;
        RECT 66.165 158.530 67.225 158.670 ;
        RECT 66.165 156.890 66.305 158.530 ;
        RECT 67.085 157.910 67.225 158.530 ;
        RECT 67.025 157.590 67.285 157.910 ;
        RECT 66.625 157.170 68.145 157.310 ;
        RECT 66.105 156.570 66.365 156.890 ;
        RECT 66.625 156.745 66.765 157.170 ;
        RECT 67.025 156.800 67.285 156.890 ;
        RECT 66.555 156.375 66.835 156.745 ;
        RECT 67.025 156.660 67.685 156.800 ;
        RECT 67.025 156.570 67.285 156.660 ;
        RECT 65.245 155.980 66.765 156.120 ;
        RECT 64.550 155.355 66.090 155.725 ;
        RECT 66.625 154.170 66.765 155.980 ;
        RECT 67.015 155.015 67.295 155.385 ;
        RECT 67.025 154.870 67.285 155.015 ;
        RECT 67.545 155.010 67.685 156.660 ;
        RECT 68.005 155.190 68.145 157.170 ;
        RECT 68.405 156.910 68.665 157.230 ;
        RECT 67.480 154.870 67.685 155.010 ;
        RECT 67.945 154.870 68.205 155.190 ;
        RECT 67.480 154.590 67.620 154.870 ;
        RECT 67.085 154.450 67.620 154.590 ;
        RECT 66.565 154.080 66.825 154.170 ;
        RECT 66.165 153.940 66.825 154.080 ;
        RECT 64.725 153.170 64.985 153.490 ;
        RECT 64.785 152.130 64.925 153.170 ;
        RECT 66.165 152.130 66.305 153.940 ;
        RECT 66.565 153.850 66.825 153.940 ;
        RECT 67.085 153.830 67.225 154.450 ;
        RECT 67.025 153.510 67.285 153.830 ;
        RECT 68.465 153.345 68.605 156.910 ;
        RECT 68.925 153.490 69.065 159.095 ;
        RECT 67.015 153.230 67.295 153.345 ;
        RECT 66.625 153.090 67.295 153.230 ;
        RECT 64.725 151.810 64.985 152.130 ;
        RECT 66.105 151.810 66.365 152.130 ;
        RECT 64.550 149.915 66.090 150.285 ;
        RECT 66.625 149.070 66.765 153.090 ;
        RECT 67.015 152.975 67.295 153.090 ;
        RECT 68.395 152.975 68.675 153.345 ;
        RECT 68.865 153.170 69.125 153.490 ;
        RECT 68.855 151.615 69.135 151.985 ;
        RECT 68.925 151.450 69.065 151.615 ;
        RECT 68.865 151.130 69.125 151.450 ;
        RECT 67.485 150.450 67.745 150.770 ;
        RECT 68.865 150.625 69.125 150.770 ;
        RECT 64.265 148.750 64.525 149.070 ;
        RECT 66.105 148.750 66.365 149.070 ;
        RECT 66.565 148.750 66.825 149.070 ;
        RECT 67.025 148.750 67.285 149.070 ;
        RECT 64.325 146.690 64.465 148.750 ;
        RECT 66.165 148.585 66.305 148.750 ;
        RECT 66.095 148.215 66.375 148.585 ;
        RECT 64.265 146.370 64.525 146.690 ;
        RECT 64.550 144.475 66.090 144.845 ;
        RECT 64.265 143.650 64.525 143.970 ;
        RECT 66.625 143.880 66.765 148.750 ;
        RECT 67.085 146.545 67.225 148.750 ;
        RECT 67.545 148.390 67.685 150.450 ;
        RECT 68.855 150.255 69.135 150.625 ;
        RECT 67.485 148.070 67.745 148.390 ;
        RECT 68.405 147.730 68.665 148.050 ;
        RECT 68.865 147.730 69.125 148.050 ;
        RECT 67.015 146.175 67.295 146.545 ;
        RECT 68.465 146.350 68.605 147.730 ;
        RECT 68.405 146.030 68.665 146.350 ;
        RECT 66.165 143.740 66.765 143.880 ;
        RECT 68.405 143.825 68.665 143.970 ;
        RECT 64.325 142.610 64.465 143.650 ;
        RECT 65.185 143.310 65.445 143.630 ;
        RECT 64.265 142.290 64.525 142.610 ;
        RECT 64.725 142.290 64.985 142.610 ;
        RECT 64.325 141.590 64.465 142.290 ;
        RECT 64.265 141.270 64.525 141.590 ;
        RECT 64.785 140.570 64.925 142.290 ;
        RECT 65.245 141.105 65.385 143.310 ;
        RECT 66.165 142.950 66.305 143.740 ;
        RECT 67.025 143.310 67.285 143.630 ;
        RECT 68.395 143.455 68.675 143.825 ;
        RECT 66.105 142.630 66.365 142.950 ;
        RECT 67.085 141.785 67.225 143.310 ;
        RECT 68.405 142.970 68.665 143.290 ;
        RECT 68.465 141.785 68.605 142.970 ;
        RECT 67.015 141.415 67.295 141.785 ;
        RECT 68.395 141.415 68.675 141.785 ;
        RECT 68.925 141.590 69.065 147.730 ;
        RECT 69.385 143.290 69.525 162.010 ;
        RECT 69.785 161.670 70.045 161.990 ;
        RECT 69.845 157.570 69.985 161.670 ;
        RECT 69.785 157.250 70.045 157.570 ;
        RECT 69.775 154.335 70.055 154.705 ;
        RECT 69.785 154.190 70.045 154.335 ;
        RECT 69.785 153.170 70.045 153.490 ;
        RECT 69.325 142.970 69.585 143.290 ;
        RECT 65.175 140.735 65.455 141.105 ;
        RECT 67.085 140.570 67.225 141.415 ;
        RECT 67.945 140.590 68.205 140.910 ;
        RECT 64.725 140.250 64.985 140.570 ;
        RECT 67.025 140.250 67.285 140.570 ;
        RECT 67.475 140.055 67.755 140.425 ;
        RECT 64.550 139.035 66.090 139.405 ;
        RECT 67.545 138.870 67.685 140.055 ;
        RECT 67.485 138.550 67.745 138.870 ;
        RECT 66.105 136.850 66.365 137.170 ;
        RECT 66.165 135.810 66.305 136.850 ;
        RECT 66.105 135.490 66.365 135.810 ;
        RECT 63.805 135.150 64.065 135.470 ;
        RECT 64.265 134.985 64.525 135.130 ;
        RECT 61.495 133.255 61.775 133.625 ;
        RECT 60.585 132.090 60.845 132.410 ;
        RECT 60.645 130.710 60.785 132.090 ;
        RECT 60.585 130.390 60.845 130.710 ;
        RECT 60.125 126.650 60.385 126.970 ;
        RECT 60.185 123.910 60.325 126.650 ;
        RECT 60.125 123.590 60.385 123.910 ;
        RECT 60.185 121.530 60.325 123.590 ;
        RECT 60.125 121.210 60.385 121.530 ;
        RECT 59.665 120.530 59.925 120.850 ;
        RECT 59.205 119.510 59.465 119.830 ;
        RECT 57.825 118.830 58.085 119.150 ;
        RECT 58.745 118.830 59.005 119.150 ;
        RECT 57.885 118.550 58.025 118.830 ;
        RECT 59.265 118.550 59.405 119.510 ;
        RECT 59.665 119.170 59.925 119.490 ;
        RECT 57.885 118.410 59.405 118.550 ;
        RECT 57.365 118.040 57.625 118.130 ;
        RECT 59.205 118.040 59.465 118.130 ;
        RECT 57.365 117.900 59.465 118.040 ;
        RECT 57.365 117.810 57.625 117.900 ;
        RECT 59.205 117.810 59.465 117.900 ;
        RECT 59.725 116.430 59.865 119.170 ;
        RECT 60.185 116.430 60.325 121.210 ;
        RECT 60.585 119.170 60.845 119.490 ;
        RECT 61.045 119.345 61.305 119.490 ;
        RECT 59.665 116.110 59.925 116.430 ;
        RECT 60.125 116.110 60.385 116.430 ;
        RECT 60.185 113.710 60.325 116.110 ;
        RECT 60.645 116.090 60.785 119.170 ;
        RECT 61.035 118.975 61.315 119.345 ;
        RECT 60.585 115.770 60.845 116.090 ;
        RECT 60.125 113.390 60.385 113.710 ;
        RECT 57.365 112.710 57.625 113.030 ;
        RECT 57.425 110.990 57.565 112.710 ;
        RECT 60.185 111.670 60.325 113.390 ;
        RECT 60.125 111.350 60.385 111.670 ;
        RECT 59.665 111.010 59.925 111.330 ;
        RECT 57.365 110.670 57.625 110.990 ;
        RECT 57.425 107.930 57.565 110.670 ;
        RECT 58.285 110.330 58.545 110.650 ;
        RECT 57.365 107.610 57.625 107.930 ;
        RECT 57.825 104.890 58.085 105.210 ;
        RECT 57.885 103.510 58.025 104.890 ;
        RECT 57.825 103.190 58.085 103.510 ;
        RECT 56.905 102.170 57.165 102.490 ;
        RECT 58.345 98.340 58.485 110.330 ;
        RECT 59.205 107.610 59.465 107.930 ;
        RECT 59.265 104.530 59.405 107.610 ;
        RECT 59.205 104.210 59.465 104.530 ;
        RECT 59.265 102.490 59.405 104.210 ;
        RECT 59.725 103.510 59.865 111.010 ;
        RECT 60.185 108.610 60.325 111.350 ;
        RECT 60.125 108.290 60.385 108.610 ;
        RECT 60.185 105.890 60.325 108.290 ;
        RECT 61.565 107.930 61.705 133.255 ;
        RECT 62.025 118.810 62.165 134.615 ;
        RECT 62.425 134.470 62.685 134.790 ;
        RECT 63.405 134.730 64.005 134.870 ;
        RECT 62.485 133.430 62.625 134.470 ;
        RECT 63.345 134.130 63.605 134.450 ;
        RECT 62.425 133.110 62.685 133.430 ;
        RECT 63.405 133.090 63.545 134.130 ;
        RECT 63.345 132.770 63.605 133.090 ;
        RECT 63.345 131.410 63.605 131.730 ;
        RECT 62.425 126.990 62.685 127.310 ;
        RECT 62.485 122.550 62.625 126.990 ;
        RECT 63.405 125.270 63.545 131.410 ;
        RECT 63.345 124.950 63.605 125.270 ;
        RECT 63.865 124.670 64.005 134.730 ;
        RECT 64.255 134.615 64.535 134.985 ;
        RECT 66.565 134.130 66.825 134.450 ;
        RECT 64.550 133.595 66.090 133.965 ;
        RECT 66.625 132.750 66.765 134.130 ;
        RECT 66.565 132.430 66.825 132.750 ;
        RECT 66.565 129.030 66.825 129.350 ;
        RECT 64.550 128.155 66.090 128.525 ;
        RECT 65.185 126.990 65.445 127.310 ;
        RECT 62.945 124.530 64.005 124.670 ;
        RECT 62.945 124.250 63.085 124.530 ;
        RECT 62.885 123.930 63.145 124.250 ;
        RECT 64.725 124.105 64.985 124.250 ;
        RECT 62.425 122.230 62.685 122.550 ;
        RECT 61.965 118.665 62.225 118.810 ;
        RECT 61.955 118.295 62.235 118.665 ;
        RECT 62.425 116.450 62.685 116.770 ;
        RECT 62.485 114.390 62.625 116.450 ;
        RECT 62.425 114.070 62.685 114.390 ;
        RECT 62.945 113.370 63.085 123.930 ;
        RECT 64.715 123.735 64.995 124.105 ;
        RECT 65.245 123.910 65.385 126.990 ;
        RECT 66.105 124.950 66.365 125.270 ;
        RECT 66.165 124.105 66.305 124.950 ;
        RECT 64.785 123.570 64.925 123.735 ;
        RECT 65.185 123.590 65.445 123.910 ;
        RECT 66.095 123.735 66.375 124.105 ;
        RECT 64.725 123.250 64.985 123.570 ;
        RECT 64.550 122.715 66.090 123.085 ;
        RECT 66.095 121.695 66.375 122.065 ;
        RECT 63.345 120.530 63.605 120.850 ;
        RECT 63.405 119.150 63.545 120.530 ;
        RECT 63.345 118.830 63.605 119.150 ;
        RECT 63.405 117.110 63.545 118.830 ;
        RECT 66.165 118.380 66.305 121.695 ;
        RECT 66.625 119.830 66.765 129.030 ;
        RECT 67.015 127.135 67.295 127.505 ;
        RECT 67.085 124.250 67.225 127.135 ;
        RECT 67.485 126.825 67.745 126.970 ;
        RECT 67.475 126.455 67.755 126.825 ;
        RECT 68.005 124.590 68.145 140.590 ;
        RECT 68.465 140.310 68.605 141.415 ;
        RECT 68.865 141.270 69.125 141.590 ;
        RECT 68.465 140.170 69.065 140.310 ;
        RECT 68.405 139.570 68.665 139.890 ;
        RECT 68.465 130.710 68.605 139.570 ;
        RECT 68.925 138.870 69.065 140.170 ;
        RECT 68.865 138.550 69.125 138.870 ;
        RECT 69.385 138.190 69.525 142.970 ;
        RECT 69.325 137.870 69.585 138.190 ;
        RECT 69.325 136.850 69.585 137.170 ;
        RECT 68.865 132.090 69.125 132.410 ;
        RECT 68.405 130.390 68.665 130.710 ;
        RECT 68.925 130.030 69.065 132.090 ;
        RECT 68.865 129.710 69.125 130.030 ;
        RECT 69.385 129.430 69.525 136.850 ;
        RECT 69.845 135.130 69.985 153.170 ;
        RECT 70.305 146.350 70.445 162.690 ;
        RECT 70.765 149.070 70.905 165.410 ;
        RECT 71.225 164.710 71.365 166.770 ;
        RECT 71.685 166.070 71.825 172.980 ;
        RECT 72.145 172.530 72.285 178.670 ;
        RECT 73.925 177.990 74.185 178.310 ;
        RECT 73.005 177.650 73.265 177.970 ;
        RECT 73.065 176.950 73.205 177.650 ;
        RECT 73.005 176.630 73.265 176.950 ;
        RECT 73.985 176.610 74.125 177.990 ;
        RECT 74.445 176.950 74.585 181.390 ;
        RECT 78.065 180.370 78.325 180.690 ;
        RECT 76.335 179.835 77.875 180.205 ;
        RECT 78.125 178.310 78.265 180.370 ;
        RECT 79.505 178.990 79.645 183.090 ;
        RECT 81.805 181.370 81.945 183.770 ;
        RECT 83.125 183.430 83.385 183.750 ;
        RECT 90.025 183.430 90.285 183.750 ;
        RECT 83.185 182.610 83.325 183.430 ;
        RECT 85.425 183.090 85.685 183.410 ;
        RECT 83.185 182.470 83.785 182.610 ;
        RECT 83.645 181.370 83.785 182.470 ;
        RECT 85.485 182.050 85.625 183.090 ;
        RECT 88.125 182.555 89.665 182.925 ;
        RECT 90.085 182.390 90.225 183.430 ;
        RECT 90.025 182.070 90.285 182.390 ;
        RECT 85.425 181.730 85.685 182.050 ;
        RECT 90.945 181.730 91.205 182.050 ;
        RECT 81.745 181.050 82.005 181.370 ;
        RECT 83.585 181.050 83.845 181.370 ;
        RECT 81.805 180.690 81.945 181.050 ;
        RECT 81.745 180.370 82.005 180.690 ;
        RECT 79.445 178.670 79.705 178.990 ;
        RECT 83.125 178.900 83.385 178.990 ;
        RECT 83.645 178.900 83.785 181.050 ;
        RECT 83.125 178.760 83.785 178.900 ;
        RECT 83.125 178.670 83.385 178.760 ;
        RECT 78.065 177.990 78.325 178.310 ;
        RECT 74.385 176.630 74.645 176.950 ;
        RECT 73.925 176.290 74.185 176.610 ;
        RECT 73.005 175.270 73.265 175.590 ;
        RECT 73.065 173.550 73.205 175.270 ;
        RECT 73.005 173.230 73.265 173.550 ;
        RECT 72.085 172.210 72.345 172.530 ;
        RECT 71.625 165.750 71.885 166.070 ;
        RECT 71.685 165.390 71.825 165.750 ;
        RECT 71.625 165.070 71.885 165.390 ;
        RECT 72.145 165.050 72.285 172.210 ;
        RECT 73.465 170.510 73.725 170.830 ;
        RECT 73.525 168.110 73.665 170.510 ;
        RECT 73.465 167.790 73.725 168.110 ;
        RECT 73.525 165.390 73.665 167.790 ;
        RECT 73.465 165.070 73.725 165.390 ;
        RECT 72.085 164.730 72.345 165.050 ;
        RECT 73.985 164.790 74.125 176.290 ;
        RECT 74.445 173.210 74.585 176.630 ;
        RECT 75.305 176.290 75.565 176.610 ;
        RECT 74.845 174.930 75.105 175.250 ;
        RECT 74.385 172.890 74.645 173.210 ;
        RECT 74.445 170.830 74.585 172.890 ;
        RECT 74.905 172.530 75.045 174.930 ;
        RECT 75.365 174.230 75.505 176.290 ;
        RECT 83.185 175.930 83.325 178.670 ;
        RECT 88.125 177.115 89.665 177.485 ;
        RECT 90.025 176.630 90.285 176.950 ;
        RECT 85.425 176.290 85.685 176.610 ;
        RECT 81.745 175.610 82.005 175.930 ;
        RECT 83.125 175.610 83.385 175.930 ;
        RECT 76.335 174.395 77.875 174.765 ;
        RECT 81.805 174.230 81.945 175.610 ;
        RECT 75.305 173.910 75.565 174.230 ;
        RECT 81.745 173.910 82.005 174.230 ;
        RECT 78.525 173.230 78.785 173.550 ;
        RECT 74.845 172.210 75.105 172.530 ;
        RECT 78.065 172.210 78.325 172.530 ;
        RECT 74.385 170.510 74.645 170.830 ;
        RECT 74.385 169.830 74.645 170.150 ;
        RECT 74.445 165.730 74.585 169.830 ;
        RECT 74.385 165.410 74.645 165.730 ;
        RECT 71.165 164.390 71.425 164.710 ;
        RECT 73.985 164.650 74.585 164.790 ;
        RECT 70.705 148.750 70.965 149.070 ;
        RECT 70.705 148.070 70.965 148.390 ;
        RECT 70.765 147.030 70.905 148.070 ;
        RECT 70.705 146.710 70.965 147.030 ;
        RECT 70.245 146.030 70.505 146.350 ;
        RECT 70.705 141.270 70.965 141.590 ;
        RECT 70.765 140.570 70.905 141.270 ;
        RECT 70.705 140.480 70.965 140.570 ;
        RECT 70.305 140.340 70.965 140.480 ;
        RECT 70.305 138.530 70.445 140.340 ;
        RECT 70.705 140.250 70.965 140.340 ;
        RECT 70.705 139.570 70.965 139.890 ;
        RECT 70.245 138.210 70.505 138.530 ;
        RECT 70.305 137.705 70.445 138.210 ;
        RECT 70.765 138.190 70.905 139.570 ;
        RECT 71.225 138.870 71.365 164.390 ;
        RECT 73.005 164.050 73.265 164.370 ;
        RECT 72.085 162.185 72.345 162.330 ;
        RECT 71.625 161.670 71.885 161.990 ;
        RECT 72.075 161.815 72.355 162.185 ;
        RECT 71.685 160.630 71.825 161.670 ;
        RECT 71.625 160.310 71.885 160.630 ;
        RECT 72.145 154.705 72.285 161.815 ;
        RECT 72.545 160.310 72.805 160.630 ;
        RECT 72.605 157.230 72.745 160.310 ;
        RECT 72.545 156.910 72.805 157.230 ;
        RECT 72.605 155.385 72.745 156.910 ;
        RECT 72.535 155.015 72.815 155.385 ;
        RECT 72.075 154.335 72.355 154.705 ;
        RECT 72.545 153.510 72.805 153.830 ;
        RECT 72.085 153.170 72.345 153.490 ;
        RECT 71.625 150.790 71.885 151.110 ;
        RECT 71.685 149.750 71.825 150.790 ;
        RECT 71.625 149.430 71.885 149.750 ;
        RECT 71.625 148.750 71.885 149.070 ;
        RECT 71.685 140.570 71.825 148.750 ;
        RECT 71.625 140.250 71.885 140.570 ;
        RECT 71.165 138.550 71.425 138.870 ;
        RECT 70.705 137.870 70.965 138.190 ;
        RECT 70.235 137.335 70.515 137.705 ;
        RECT 69.785 134.810 70.045 135.130 ;
        RECT 70.245 134.130 70.505 134.450 ;
        RECT 71.625 134.130 71.885 134.450 ;
        RECT 69.785 131.410 70.045 131.730 ;
        RECT 69.845 129.690 69.985 131.410 ;
        RECT 68.465 129.290 69.525 129.430 ;
        RECT 69.785 129.370 70.045 129.690 ;
        RECT 68.465 127.650 68.605 129.290 ;
        RECT 69.315 128.495 69.595 128.865 ;
        RECT 68.405 127.330 68.665 127.650 ;
        RECT 68.405 126.310 68.665 126.630 ;
        RECT 67.485 124.270 67.745 124.590 ;
        RECT 67.945 124.270 68.205 124.590 ;
        RECT 67.025 123.930 67.285 124.250 ;
        RECT 67.545 123.990 67.685 124.270 ;
        RECT 68.465 124.250 68.605 126.310 ;
        RECT 68.865 125.970 69.125 126.290 ;
        RECT 67.545 123.850 68.145 123.990 ;
        RECT 68.405 123.930 68.665 124.250 ;
        RECT 67.025 122.230 67.285 122.550 ;
        RECT 67.085 119.830 67.225 122.230 ;
        RECT 67.485 121.550 67.745 121.870 ;
        RECT 66.565 119.510 66.825 119.830 ;
        RECT 67.025 119.510 67.285 119.830 ;
        RECT 66.165 118.240 66.765 118.380 ;
        RECT 64.550 117.275 66.090 117.645 ;
        RECT 63.345 116.790 63.605 117.110 ;
        RECT 62.885 113.050 63.145 113.370 ;
        RECT 63.795 112.855 64.075 113.225 ;
        RECT 63.865 107.930 64.005 112.855 ;
        RECT 64.550 111.835 66.090 112.205 ;
        RECT 66.625 111.670 66.765 118.240 ;
        RECT 67.545 117.110 67.685 121.550 ;
        RECT 68.005 119.830 68.145 123.850 ;
        RECT 68.925 122.210 69.065 125.970 ;
        RECT 69.385 123.570 69.525 128.495 ;
        RECT 70.305 128.070 70.445 134.130 ;
        RECT 71.165 131.750 71.425 132.070 ;
        RECT 71.225 130.710 71.365 131.750 ;
        RECT 71.165 130.390 71.425 130.710 ;
        RECT 70.705 129.545 70.965 129.690 ;
        RECT 70.695 129.175 70.975 129.545 ;
        RECT 71.225 129.350 71.365 130.390 ;
        RECT 71.165 129.030 71.425 129.350 ;
        RECT 70.705 128.690 70.965 129.010 ;
        RECT 69.845 127.930 70.445 128.070 ;
        RECT 69.845 124.930 69.985 127.930 ;
        RECT 70.245 126.310 70.505 126.630 ;
        RECT 70.305 125.270 70.445 126.310 ;
        RECT 70.765 126.290 70.905 128.690 ;
        RECT 71.225 127.310 71.365 129.030 ;
        RECT 71.165 126.990 71.425 127.310 ;
        RECT 70.705 125.970 70.965 126.290 ;
        RECT 71.165 125.970 71.425 126.290 ;
        RECT 70.245 124.950 70.505 125.270 ;
        RECT 69.785 124.610 70.045 124.930 ;
        RECT 69.325 123.250 69.585 123.570 ;
        RECT 69.385 122.550 69.525 123.250 ;
        RECT 69.325 122.230 69.585 122.550 ;
        RECT 68.865 121.890 69.125 122.210 ;
        RECT 69.845 121.870 69.985 124.610 ;
        RECT 70.245 123.250 70.505 123.570 ;
        RECT 69.785 121.550 70.045 121.870 ;
        RECT 70.305 121.530 70.445 123.250 ;
        RECT 71.225 122.550 71.365 125.970 ;
        RECT 71.165 122.230 71.425 122.550 ;
        RECT 70.245 121.210 70.505 121.530 ;
        RECT 67.945 119.510 68.205 119.830 ;
        RECT 67.485 116.790 67.745 117.110 ;
        RECT 70.305 116.770 70.445 121.210 ;
        RECT 71.225 119.830 71.365 122.230 ;
        RECT 71.165 119.510 71.425 119.830 ;
        RECT 71.165 118.830 71.425 119.150 ;
        RECT 70.245 116.450 70.505 116.770 ;
        RECT 69.785 116.110 70.045 116.430 ;
        RECT 69.845 115.410 69.985 116.110 ;
        RECT 69.785 115.090 70.045 115.410 ;
        RECT 69.785 113.225 70.045 113.370 ;
        RECT 69.775 112.855 70.055 113.225 ;
        RECT 70.705 112.940 70.965 113.030 ;
        RECT 71.225 112.940 71.365 118.830 ;
        RECT 70.705 112.800 71.365 112.940 ;
        RECT 70.705 112.710 70.965 112.800 ;
        RECT 66.565 111.350 66.825 111.670 ;
        RECT 71.225 110.990 71.365 112.800 ;
        RECT 71.165 110.670 71.425 110.990 ;
        RECT 64.265 110.330 64.525 110.650 ;
        RECT 64.325 108.950 64.465 110.330 ;
        RECT 64.265 108.630 64.525 108.950 ;
        RECT 61.505 107.610 61.765 107.930 ;
        RECT 63.805 107.610 64.065 107.930 ;
        RECT 67.485 107.270 67.745 107.590 ;
        RECT 71.165 107.270 71.425 107.590 ;
        RECT 61.505 106.930 61.765 107.250 ;
        RECT 61.565 105.890 61.705 106.930 ;
        RECT 64.550 106.395 66.090 106.765 ;
        RECT 60.125 105.570 60.385 105.890 ;
        RECT 61.505 105.570 61.765 105.890 ;
        RECT 62.885 104.890 63.145 105.210 ;
        RECT 59.665 103.190 59.925 103.510 ;
        RECT 59.205 102.170 59.465 102.490 ;
        RECT 62.945 98.340 63.085 104.890 ;
        RECT 64.550 100.955 66.090 101.325 ;
        RECT 67.545 98.340 67.685 107.270 ;
        RECT 70.245 106.930 70.505 107.250 ;
        RECT 70.305 105.890 70.445 106.930 ;
        RECT 70.245 105.570 70.505 105.890 ;
        RECT 71.225 103.510 71.365 107.270 ;
        RECT 71.685 105.890 71.825 134.130 ;
        RECT 72.145 132.750 72.285 153.170 ;
        RECT 72.605 152.470 72.745 153.510 ;
        RECT 72.545 152.150 72.805 152.470 ;
        RECT 72.605 151.450 72.745 152.150 ;
        RECT 72.545 151.130 72.805 151.450 ;
        RECT 72.545 150.625 72.805 150.770 ;
        RECT 72.535 150.255 72.815 150.625 ;
        RECT 73.065 149.070 73.205 164.050 ;
        RECT 73.465 155.890 73.725 156.210 ;
        RECT 73.525 154.170 73.665 155.890 ;
        RECT 73.925 154.870 74.185 155.190 ;
        RECT 73.985 154.510 74.125 154.870 ;
        RECT 73.925 154.190 74.185 154.510 ;
        RECT 73.465 153.850 73.725 154.170 ;
        RECT 73.465 153.170 73.725 153.490 ;
        RECT 73.525 151.305 73.665 153.170 ;
        RECT 73.985 151.985 74.125 154.190 ;
        RECT 73.915 151.615 74.195 151.985 ;
        RECT 73.985 151.450 74.125 151.615 ;
        RECT 73.455 150.935 73.735 151.305 ;
        RECT 73.925 151.130 74.185 151.450 ;
        RECT 73.005 148.750 73.265 149.070 ;
        RECT 72.545 148.410 72.805 148.730 ;
        RECT 72.605 143.630 72.745 148.410 ;
        RECT 72.545 143.310 72.805 143.630 ;
        RECT 73.525 143.030 73.665 150.935 ;
        RECT 73.925 150.450 74.185 150.770 ;
        RECT 73.985 149.410 74.125 150.450 ;
        RECT 73.925 149.090 74.185 149.410 ;
        RECT 72.605 142.890 73.665 143.030 ;
        RECT 72.085 132.430 72.345 132.750 ;
        RECT 72.605 129.430 72.745 142.890 ;
        RECT 72.995 141.415 73.275 141.785 ;
        RECT 73.005 141.270 73.265 141.415 ;
        RECT 73.005 140.250 73.265 140.570 ;
        RECT 73.065 138.190 73.205 140.250 ;
        RECT 74.445 139.890 74.585 164.650 ;
        RECT 73.925 139.570 74.185 139.890 ;
        RECT 74.385 139.570 74.645 139.890 ;
        RECT 73.005 137.870 73.265 138.190 ;
        RECT 73.465 136.850 73.725 137.170 ;
        RECT 73.005 134.470 73.265 134.790 ;
        RECT 73.065 132.750 73.205 134.470 ;
        RECT 73.005 132.430 73.265 132.750 ;
        RECT 73.525 132.410 73.665 136.850 ;
        RECT 73.985 135.470 74.125 139.570 ;
        RECT 74.905 137.850 75.045 172.210 ;
        RECT 75.765 170.850 76.025 171.170 ;
        RECT 75.305 169.490 75.565 169.810 ;
        RECT 75.365 167.430 75.505 169.490 ;
        RECT 75.305 167.110 75.565 167.430 ;
        RECT 75.825 166.070 75.965 170.850 ;
        RECT 76.335 168.955 77.875 169.325 ;
        RECT 75.765 165.750 76.025 166.070 ;
        RECT 78.125 165.050 78.265 172.210 ;
        RECT 78.585 169.810 78.725 173.230 ;
        RECT 79.905 172.890 80.165 173.210 ;
        RECT 78.525 169.490 78.785 169.810 ;
        RECT 78.585 168.790 78.725 169.490 ;
        RECT 78.525 168.470 78.785 168.790 ;
        RECT 78.585 165.390 78.725 168.470 ;
        RECT 79.965 166.070 80.105 172.890 ;
        RECT 80.365 172.210 80.625 172.530 ;
        RECT 80.425 168.110 80.565 172.210 ;
        RECT 83.185 170.490 83.325 175.610 ;
        RECT 85.485 174.230 85.625 176.290 ;
        RECT 87.725 175.950 87.985 176.270 ;
        RECT 85.425 173.910 85.685 174.230 ;
        RECT 84.965 172.890 85.225 173.210 ;
        RECT 85.025 171.510 85.165 172.890 ;
        RECT 86.805 172.210 87.065 172.530 ;
        RECT 84.965 171.190 85.225 171.510 ;
        RECT 83.585 170.850 83.845 171.170 ;
        RECT 80.825 170.170 81.085 170.490 ;
        RECT 83.125 170.170 83.385 170.490 ;
        RECT 80.365 167.790 80.625 168.110 ;
        RECT 80.885 167.430 81.025 170.170 ;
        RECT 83.645 168.790 83.785 170.850 ;
        RECT 86.865 170.490 87.005 172.210 ;
        RECT 87.785 171.510 87.925 175.950 ;
        RECT 88.645 175.610 88.905 175.930 ;
        RECT 88.705 173.210 88.845 175.610 ;
        RECT 88.645 172.890 88.905 173.210 ;
        RECT 88.125 171.675 89.665 172.045 ;
        RECT 87.725 171.190 87.985 171.510 ;
        RECT 86.805 170.170 87.065 170.490 ;
        RECT 83.585 168.470 83.845 168.790 ;
        RECT 80.825 167.110 81.085 167.430 ;
        RECT 80.365 166.770 80.625 167.090 ;
        RECT 79.905 165.750 80.165 166.070 ;
        RECT 80.425 165.730 80.565 166.770 ;
        RECT 80.365 165.410 80.625 165.730 ;
        RECT 80.885 165.390 81.025 167.110 ;
        RECT 86.865 167.090 87.005 170.170 ;
        RECT 90.085 168.110 90.225 176.630 ;
        RECT 90.485 175.270 90.745 175.590 ;
        RECT 90.545 171.170 90.685 175.270 ;
        RECT 90.485 170.850 90.745 171.170 ;
        RECT 90.025 167.790 90.285 168.110 ;
        RECT 90.025 167.110 90.285 167.430 ;
        RECT 86.805 166.770 87.065 167.090 ;
        RECT 87.725 166.770 87.985 167.090 ;
        RECT 83.585 165.750 83.845 166.070 ;
        RECT 86.345 165.750 86.605 166.070 ;
        RECT 78.525 165.070 78.785 165.390 ;
        RECT 80.825 165.070 81.085 165.390 ;
        RECT 75.765 164.730 76.025 165.050 ;
        RECT 78.065 164.730 78.325 165.050 ;
        RECT 75.825 163.350 75.965 164.730 ;
        RECT 79.905 164.050 80.165 164.370 ;
        RECT 76.335 163.515 77.875 163.885 ;
        RECT 75.765 163.030 76.025 163.350 ;
        RECT 75.305 158.950 75.565 159.270 ;
        RECT 75.365 156.890 75.505 158.950 ;
        RECT 76.335 158.075 77.875 158.445 ;
        RECT 75.305 156.570 75.565 156.890 ;
        RECT 75.365 154.850 75.505 156.570 ;
        RECT 79.965 156.550 80.105 164.050 ;
        RECT 80.365 163.030 80.625 163.350 ;
        RECT 80.425 160.290 80.565 163.030 ;
        RECT 80.885 163.010 81.025 165.070 ;
        RECT 80.825 162.690 81.085 163.010 ;
        RECT 80.365 159.970 80.625 160.290 ;
        RECT 80.885 159.610 81.025 162.690 ;
        RECT 83.645 162.670 83.785 165.750 ;
        RECT 83.585 162.350 83.845 162.670 ;
        RECT 84.965 162.010 85.225 162.330 ;
        RECT 84.045 161.330 84.305 161.650 ;
        RECT 84.105 160.630 84.245 161.330 ;
        RECT 84.045 160.310 84.305 160.630 ;
        RECT 85.025 160.290 85.165 162.010 ;
        RECT 84.965 159.970 85.225 160.290 ;
        RECT 80.825 159.290 81.085 159.610 ;
        RECT 84.505 159.290 84.765 159.610 ;
        RECT 84.565 157.230 84.705 159.290 ;
        RECT 84.505 156.910 84.765 157.230 ;
        RECT 79.905 156.230 80.165 156.550 ;
        RECT 84.045 156.230 84.305 156.550 ;
        RECT 78.065 155.890 78.325 156.210 ;
        RECT 80.365 155.890 80.625 156.210 ;
        RECT 78.125 155.190 78.265 155.890 ;
        RECT 80.425 155.190 80.565 155.890 ;
        RECT 78.065 154.870 78.325 155.190 ;
        RECT 80.365 154.870 80.625 155.190 ;
        RECT 75.305 154.530 75.565 154.850 ;
        RECT 81.285 154.530 81.545 154.850 ;
        RECT 75.765 154.190 76.025 154.510 ;
        RECT 78.985 154.190 79.245 154.510 ;
        RECT 75.305 153.850 75.565 154.170 ;
        RECT 75.825 154.025 75.965 154.190 ;
        RECT 75.365 152.130 75.505 153.850 ;
        RECT 75.755 153.655 76.035 154.025 ;
        RECT 76.335 152.635 77.875 153.005 ;
        RECT 75.305 151.810 75.565 152.130 ;
        RECT 79.045 150.770 79.185 154.190 ;
        RECT 81.345 153.910 81.485 154.530 ;
        RECT 81.735 154.335 82.015 154.705 ;
        RECT 81.745 154.190 82.005 154.335 ;
        RECT 81.345 153.770 81.945 153.910 ;
        RECT 79.905 150.790 80.165 151.110 ;
        RECT 78.985 150.450 79.245 150.770 ;
        RECT 79.965 149.750 80.105 150.790 ;
        RECT 79.905 149.430 80.165 149.750 ;
        RECT 81.805 148.730 81.945 153.770 ;
        RECT 82.205 150.450 82.465 150.770 ;
        RECT 83.125 150.450 83.385 150.770 ;
        RECT 82.265 149.750 82.405 150.450 ;
        RECT 82.205 149.430 82.465 149.750 ;
        RECT 83.185 149.070 83.325 150.450 ;
        RECT 84.105 149.410 84.245 156.230 ;
        RECT 85.025 154.850 85.165 159.970 ;
        RECT 86.405 159.950 86.545 165.750 ;
        RECT 85.425 159.630 85.685 159.950 ;
        RECT 85.885 159.630 86.145 159.950 ;
        RECT 86.345 159.630 86.605 159.950 ;
        RECT 85.485 157.910 85.625 159.630 ;
        RECT 85.945 159.465 86.085 159.630 ;
        RECT 85.875 159.095 86.155 159.465 ;
        RECT 85.425 157.590 85.685 157.910 ;
        RECT 84.965 154.530 85.225 154.850 ;
        RECT 85.945 154.170 86.085 159.095 ;
        RECT 85.885 153.850 86.145 154.170 ;
        RECT 85.885 153.170 86.145 153.490 ;
        RECT 85.945 151.450 86.085 153.170 ;
        RECT 84.965 151.130 85.225 151.450 ;
        RECT 85.885 151.130 86.145 151.450 ;
        RECT 85.025 149.750 85.165 151.130 ;
        RECT 84.965 149.430 85.225 149.750 ;
        RECT 84.045 149.090 84.305 149.410 ;
        RECT 83.125 148.750 83.385 149.070 ;
        RECT 81.745 148.410 82.005 148.730 ;
        RECT 78.985 148.070 79.245 148.390 ;
        RECT 76.335 147.195 77.875 147.565 ;
        RECT 79.045 146.010 79.185 148.070 ;
        RECT 85.945 146.350 86.085 151.130 ;
        RECT 86.865 146.350 87.005 166.770 ;
        RECT 87.785 165.730 87.925 166.770 ;
        RECT 88.125 166.235 89.665 166.605 ;
        RECT 87.725 165.410 87.985 165.730 ;
        RECT 90.085 165.050 90.225 167.110 ;
        RECT 87.725 164.730 87.985 165.050 ;
        RECT 90.025 164.730 90.285 165.050 ;
        RECT 87.785 162.330 87.925 164.730 ;
        RECT 90.085 162.330 90.225 164.730 ;
        RECT 87.725 162.010 87.985 162.330 ;
        RECT 90.025 162.010 90.285 162.330 ;
        RECT 87.725 161.330 87.985 161.650 ;
        RECT 87.785 160.630 87.925 161.330 ;
        RECT 88.125 160.795 89.665 161.165 ;
        RECT 87.725 160.310 87.985 160.630 ;
        RECT 87.265 159.860 87.525 159.950 ;
        RECT 87.785 159.860 87.925 160.310 ;
        RECT 87.265 159.720 87.925 159.860 ;
        RECT 87.265 159.630 87.525 159.720 ;
        RECT 89.565 158.950 89.825 159.270 ;
        RECT 87.265 158.610 87.525 158.930 ;
        RECT 87.725 158.610 87.985 158.930 ;
        RECT 87.325 155.190 87.465 158.610 ;
        RECT 87.265 154.870 87.525 155.190 ;
        RECT 85.885 146.030 86.145 146.350 ;
        RECT 86.805 146.030 87.065 146.350 ;
        RECT 78.985 145.690 79.245 146.010 ;
        RECT 84.505 145.350 84.765 145.670 ;
        RECT 77.145 145.010 77.405 145.330 ;
        RECT 77.205 144.310 77.345 145.010 ;
        RECT 84.565 144.310 84.705 145.350 ;
        RECT 77.145 143.990 77.405 144.310 ;
        RECT 84.505 143.990 84.765 144.310 ;
        RECT 87.785 143.630 87.925 158.610 ;
        RECT 89.625 157.230 89.765 158.950 ;
        RECT 90.085 157.230 90.225 162.010 ;
        RECT 89.565 156.910 89.825 157.230 ;
        RECT 90.025 156.910 90.285 157.230 ;
        RECT 88.125 155.355 89.665 155.725 ;
        RECT 88.645 154.530 88.905 154.850 ;
        RECT 88.705 153.830 88.845 154.530 ;
        RECT 88.645 153.510 88.905 153.830 ;
        RECT 88.705 151.450 88.845 153.510 ;
        RECT 90.085 153.490 90.225 156.910 ;
        RECT 90.485 156.230 90.745 156.550 ;
        RECT 90.025 153.170 90.285 153.490 ;
        RECT 90.545 152.470 90.685 156.230 ;
        RECT 90.485 152.150 90.745 152.470 ;
        RECT 91.005 152.130 91.145 181.730 ;
        RECT 91.405 178.670 91.665 178.990 ;
        RECT 91.465 174.230 91.605 178.670 ;
        RECT 92.385 178.650 92.525 184.110 ;
        RECT 93.765 181.370 93.905 185.810 ;
        RECT 96.065 183.750 96.205 185.810 ;
        RECT 99.910 185.275 101.450 185.645 ;
        RECT 106.125 183.770 106.385 184.090 ;
        RECT 96.005 183.430 96.265 183.750 ;
        RECT 96.925 183.090 97.185 183.410 ;
        RECT 97.845 183.090 98.105 183.410 ;
        RECT 100.605 183.090 100.865 183.410 ;
        RECT 96.985 182.050 97.125 183.090 ;
        RECT 96.925 181.730 97.185 182.050 ;
        RECT 95.085 181.390 95.345 181.710 ;
        RECT 93.705 181.050 93.965 181.370 ;
        RECT 93.765 178.990 93.905 181.050 ;
        RECT 93.705 178.670 93.965 178.990 ;
        RECT 92.325 178.330 92.585 178.650 ;
        RECT 91.405 173.910 91.665 174.230 ;
        RECT 91.465 170.490 91.605 173.910 ;
        RECT 92.385 173.550 92.525 178.330 ;
        RECT 93.705 177.650 93.965 177.970 ;
        RECT 92.325 173.230 92.585 173.550 ;
        RECT 92.325 172.270 92.585 172.530 ;
        RECT 93.765 172.440 93.905 177.650 ;
        RECT 94.165 174.930 94.425 175.250 ;
        RECT 94.225 173.550 94.365 174.930 ;
        RECT 94.165 173.230 94.425 173.550 ;
        RECT 94.165 172.440 94.425 172.530 ;
        RECT 93.765 172.300 94.425 172.440 ;
        RECT 91.925 172.210 92.585 172.270 ;
        RECT 94.165 172.210 94.425 172.300 ;
        RECT 91.925 172.130 92.525 172.210 ;
        RECT 91.405 170.170 91.665 170.490 ;
        RECT 91.405 162.010 91.665 162.330 ;
        RECT 91.465 154.850 91.605 162.010 ;
        RECT 91.405 154.530 91.665 154.850 ;
        RECT 91.405 153.170 91.665 153.490 ;
        RECT 90.945 151.810 91.205 152.130 ;
        RECT 88.645 151.130 88.905 151.450 ;
        RECT 89.565 151.360 89.825 151.450 ;
        RECT 89.565 151.220 90.225 151.360 ;
        RECT 89.565 151.130 89.825 151.220 ;
        RECT 88.125 149.915 89.665 150.285 ;
        RECT 90.085 149.410 90.225 151.220 ;
        RECT 90.485 151.130 90.745 151.450 ;
        RECT 90.945 151.305 91.205 151.450 ;
        RECT 90.025 149.150 90.285 149.410 ;
        RECT 89.625 149.090 90.285 149.150 ;
        RECT 89.625 149.010 90.225 149.090 ;
        RECT 88.645 148.110 88.905 148.390 ;
        RECT 88.645 148.070 89.305 148.110 ;
        RECT 88.705 147.970 89.305 148.070 ;
        RECT 89.165 146.010 89.305 147.970 ;
        RECT 89.625 147.030 89.765 149.010 ;
        RECT 90.545 148.390 90.685 151.130 ;
        RECT 90.935 150.935 91.215 151.305 ;
        RECT 91.005 149.750 91.145 150.935 ;
        RECT 90.945 149.430 91.205 149.750 ;
        RECT 90.485 148.070 90.745 148.390 ;
        RECT 90.025 147.730 90.285 148.050 ;
        RECT 89.565 146.710 89.825 147.030 ;
        RECT 89.625 146.010 89.765 146.710 ;
        RECT 89.105 145.690 89.365 146.010 ;
        RECT 89.565 145.690 89.825 146.010 ;
        RECT 88.125 144.475 89.665 144.845 ;
        RECT 80.825 143.310 81.085 143.630 ;
        RECT 87.725 143.310 87.985 143.630 ;
        RECT 76.335 141.755 77.875 142.125 ;
        RECT 75.765 140.930 76.025 141.250 ;
        RECT 75.825 138.190 75.965 140.930 ;
        RECT 76.685 140.250 76.945 140.570 ;
        RECT 76.745 138.530 76.885 140.250 ;
        RECT 80.885 139.890 81.025 143.310 ;
        RECT 90.085 143.290 90.225 147.730 ;
        RECT 90.545 146.350 90.685 148.070 ;
        RECT 90.485 146.030 90.745 146.350 ;
        RECT 90.485 145.010 90.745 145.330 ;
        RECT 90.025 142.970 90.285 143.290 ;
        RECT 81.285 142.630 81.545 142.950 ;
        RECT 80.825 139.570 81.085 139.890 ;
        RECT 80.885 138.870 81.025 139.570 ;
        RECT 80.825 138.550 81.085 138.870 ;
        RECT 76.685 138.210 76.945 138.530 ;
        RECT 75.765 137.870 76.025 138.190 ;
        RECT 74.845 137.530 75.105 137.850 ;
        RECT 75.765 137.190 76.025 137.510 ;
        RECT 73.925 135.150 74.185 135.470 ;
        RECT 75.825 135.040 75.965 137.190 ;
        RECT 76.335 136.315 77.875 136.685 ;
        RECT 78.525 135.830 78.785 136.150 ;
        RECT 78.065 135.490 78.325 135.810 ;
        RECT 78.125 135.130 78.265 135.490 ;
        RECT 76.225 135.040 76.485 135.130 ;
        RECT 75.825 134.900 76.485 135.040 ;
        RECT 76.225 134.810 76.485 134.900 ;
        RECT 78.065 134.810 78.325 135.130 ;
        RECT 76.285 132.750 76.425 134.810 ;
        RECT 78.125 132.750 78.265 134.810 ;
        RECT 76.225 132.430 76.485 132.750 ;
        RECT 78.065 132.430 78.325 132.750 ;
        RECT 73.465 132.090 73.725 132.410 ;
        RECT 74.845 132.090 75.105 132.410 ;
        RECT 74.385 131.410 74.645 131.730 ;
        RECT 73.465 129.710 73.725 130.030 ;
        RECT 72.605 129.290 73.205 129.430 ;
        RECT 72.545 128.690 72.805 129.010 ;
        RECT 72.605 127.650 72.745 128.690 ;
        RECT 72.545 127.330 72.805 127.650 ;
        RECT 72.085 126.990 72.345 127.310 ;
        RECT 72.145 123.570 72.285 126.990 ;
        RECT 72.085 123.250 72.345 123.570 ;
        RECT 73.065 121.270 73.205 129.290 ;
        RECT 73.525 121.530 73.665 129.710 ;
        RECT 73.925 129.370 74.185 129.690 ;
        RECT 73.985 125.270 74.125 129.370 ;
        RECT 73.925 124.950 74.185 125.270 ;
        RECT 73.985 121.870 74.125 124.950 ;
        RECT 73.925 121.550 74.185 121.870 ;
        RECT 72.605 121.130 73.205 121.270 ;
        RECT 73.465 121.210 73.725 121.530 ;
        RECT 72.605 119.150 72.745 121.130 ;
        RECT 73.005 120.530 73.265 120.850 ;
        RECT 72.545 118.830 72.805 119.150 ;
        RECT 72.545 118.150 72.805 118.470 ;
        RECT 72.605 117.110 72.745 118.150 ;
        RECT 72.545 116.790 72.805 117.110 ;
        RECT 72.545 116.110 72.805 116.430 ;
        RECT 72.085 115.090 72.345 115.410 ;
        RECT 72.145 113.710 72.285 115.090 ;
        RECT 72.085 113.390 72.345 113.710 ;
        RECT 72.605 112.690 72.745 116.110 ;
        RECT 73.065 114.390 73.205 120.530 ;
        RECT 73.005 114.070 73.265 114.390 ;
        RECT 73.985 113.710 74.125 121.550 ;
        RECT 73.925 113.390 74.185 113.710 ;
        RECT 72.545 112.370 72.805 112.690 ;
        RECT 73.985 108.950 74.125 113.390 ;
        RECT 74.445 110.990 74.585 131.410 ;
        RECT 74.905 129.690 75.045 132.090 ;
        RECT 76.335 130.875 77.875 131.245 ;
        RECT 78.125 129.690 78.265 132.430 ;
        RECT 74.845 129.370 75.105 129.690 ;
        RECT 76.225 129.370 76.485 129.690 ;
        RECT 78.065 129.370 78.325 129.690 ;
        RECT 74.905 127.310 75.045 129.370 ;
        RECT 76.285 127.650 76.425 129.370 ;
        RECT 74.845 126.990 75.105 127.310 ;
        RECT 75.295 127.135 75.575 127.505 ;
        RECT 76.225 127.330 76.485 127.650 ;
        RECT 75.305 126.990 75.565 127.135 ;
        RECT 76.685 126.710 76.945 126.970 ;
        RECT 75.365 126.650 76.945 126.710 ;
        RECT 78.065 126.650 78.325 126.970 ;
        RECT 75.365 126.570 76.885 126.650 ;
        RECT 74.845 121.890 75.105 122.210 ;
        RECT 74.905 111.330 75.045 121.890 ;
        RECT 75.365 116.770 75.505 126.570 ;
        RECT 76.335 125.435 77.875 125.805 ;
        RECT 78.125 123.910 78.265 126.650 ;
        RECT 78.065 123.590 78.325 123.910 ;
        RECT 75.765 121.210 76.025 121.530 ;
        RECT 78.065 121.210 78.325 121.530 ;
        RECT 75.305 116.450 75.565 116.770 ;
        RECT 75.825 116.430 75.965 121.210 ;
        RECT 76.335 119.995 77.875 120.365 ;
        RECT 78.125 119.150 78.265 121.210 ;
        RECT 78.585 119.830 78.725 135.830 ;
        RECT 80.885 135.470 81.025 138.550 ;
        RECT 81.345 137.850 81.485 142.630 ;
        RECT 90.025 142.290 90.285 142.610 ;
        RECT 85.425 140.250 85.685 140.570 ;
        RECT 87.265 140.250 87.525 140.570 ;
        RECT 84.505 139.570 84.765 139.890 ;
        RECT 84.565 138.870 84.705 139.570 ;
        RECT 85.485 138.870 85.625 140.250 ;
        RECT 84.505 138.550 84.765 138.870 ;
        RECT 85.425 138.550 85.685 138.870 ;
        RECT 81.745 137.870 82.005 138.190 ;
        RECT 85.425 137.870 85.685 138.190 ;
        RECT 81.285 137.530 81.545 137.850 ;
        RECT 81.345 135.470 81.485 137.530 ;
        RECT 80.825 135.150 81.085 135.470 ;
        RECT 81.285 135.150 81.545 135.470 ;
        RECT 80.825 134.470 81.085 134.790 ;
        RECT 80.885 129.010 81.025 134.470 ;
        RECT 81.805 134.450 81.945 137.870 ;
        RECT 82.665 135.150 82.925 135.470 ;
        RECT 81.745 134.130 82.005 134.450 ;
        RECT 81.805 132.070 81.945 134.130 ;
        RECT 81.745 131.750 82.005 132.070 ;
        RECT 80.825 128.690 81.085 129.010 ;
        RECT 79.435 127.135 79.715 127.505 ;
        RECT 79.905 127.330 80.165 127.650 ;
        RECT 78.985 121.210 79.245 121.530 ;
        RECT 79.045 119.830 79.185 121.210 ;
        RECT 78.525 119.510 78.785 119.830 ;
        RECT 78.985 119.510 79.245 119.830 ;
        RECT 78.065 118.830 78.325 119.150 ;
        RECT 77.605 118.150 77.865 118.470 ;
        RECT 75.765 116.110 76.025 116.430 ;
        RECT 77.665 116.090 77.805 118.150 ;
        RECT 78.125 116.090 78.265 118.830 ;
        RECT 79.505 118.810 79.645 127.135 ;
        RECT 79.965 121.530 80.105 127.330 ;
        RECT 80.365 126.990 80.625 127.310 ;
        RECT 80.425 124.785 80.565 126.990 ;
        RECT 80.355 124.415 80.635 124.785 ;
        RECT 80.425 124.250 80.565 124.415 ;
        RECT 80.365 123.930 80.625 124.250 ;
        RECT 80.885 123.910 81.025 128.690 ;
        RECT 81.745 125.970 82.005 126.290 ;
        RECT 80.825 123.590 81.085 123.910 ;
        RECT 79.905 121.210 80.165 121.530 ;
        RECT 79.965 118.810 80.105 121.210 ;
        RECT 81.805 118.810 81.945 125.970 ;
        RECT 82.725 124.590 82.865 135.150 ;
        RECT 85.485 135.130 85.625 137.870 ;
        RECT 85.425 134.810 85.685 135.130 ;
        RECT 85.485 132.410 85.625 134.810 ;
        RECT 86.345 134.470 86.605 134.790 ;
        RECT 85.425 132.090 85.685 132.410 ;
        RECT 86.405 130.280 86.545 134.470 ;
        RECT 86.805 134.130 87.065 134.450 ;
        RECT 86.865 132.750 87.005 134.130 ;
        RECT 87.325 132.750 87.465 140.250 ;
        RECT 87.725 139.570 87.985 139.890 ;
        RECT 86.805 132.430 87.065 132.750 ;
        RECT 87.265 132.430 87.525 132.750 ;
        RECT 86.805 130.280 87.065 130.370 ;
        RECT 86.405 130.140 87.065 130.280 ;
        RECT 86.805 130.050 87.065 130.140 ;
        RECT 84.045 129.710 84.305 130.030 ;
        RECT 84.105 126.630 84.245 129.710 ;
        RECT 85.885 126.990 86.145 127.310 ;
        RECT 84.045 126.310 84.305 126.630 ;
        RECT 85.945 125.270 86.085 126.990 ;
        RECT 85.885 124.950 86.145 125.270 ;
        RECT 83.585 124.610 83.845 124.930 ;
        RECT 82.665 124.270 82.925 124.590 ;
        RECT 82.665 121.890 82.925 122.210 ;
        RECT 78.525 118.490 78.785 118.810 ;
        RECT 79.445 118.490 79.705 118.810 ;
        RECT 79.905 118.490 80.165 118.810 ;
        RECT 81.745 118.490 82.005 118.810 ;
        RECT 77.605 115.770 77.865 116.090 ;
        RECT 78.065 115.770 78.325 116.090 ;
        RECT 75.765 115.090 76.025 115.410 ;
        RECT 75.825 113.030 75.965 115.090 ;
        RECT 76.335 114.555 77.875 114.925 ;
        RECT 78.585 114.050 78.725 118.490 ;
        RECT 79.905 117.810 80.165 118.130 ;
        RECT 79.965 116.770 80.105 117.810 ;
        RECT 79.905 116.450 80.165 116.770 ;
        RECT 79.445 116.110 79.705 116.430 ;
        RECT 79.505 114.390 79.645 116.110 ;
        RECT 79.445 114.070 79.705 114.390 ;
        RECT 78.525 113.730 78.785 114.050 ;
        RECT 82.725 113.030 82.865 121.890 ;
        RECT 83.645 118.470 83.785 124.610 ;
        RECT 86.865 123.570 87.005 130.050 ;
        RECT 87.325 130.030 87.465 132.430 ;
        RECT 87.265 129.710 87.525 130.030 ;
        RECT 87.325 127.990 87.465 129.710 ;
        RECT 87.265 127.670 87.525 127.990 ;
        RECT 86.805 123.250 87.065 123.570 ;
        RECT 87.265 121.210 87.525 121.530 ;
        RECT 87.325 119.150 87.465 121.210 ;
        RECT 87.265 118.830 87.525 119.150 ;
        RECT 83.585 118.150 83.845 118.470 ;
        RECT 83.125 116.450 83.385 116.770 ;
        RECT 83.185 113.370 83.325 116.450 ;
        RECT 83.645 114.390 83.785 118.150 ;
        RECT 83.585 114.070 83.845 114.390 ;
        RECT 83.125 113.050 83.385 113.370 ;
        RECT 75.765 112.710 76.025 113.030 ;
        RECT 82.665 112.710 82.925 113.030 ;
        RECT 83.645 111.330 83.785 114.070 ;
        RECT 74.845 111.010 75.105 111.330 ;
        RECT 83.585 111.010 83.845 111.330 ;
        RECT 74.385 110.670 74.645 110.990 ;
        RECT 87.325 110.650 87.465 118.830 ;
        RECT 87.785 110.990 87.925 139.570 ;
        RECT 88.125 139.035 89.665 139.405 ;
        RECT 88.125 133.595 89.665 133.965 ;
        RECT 88.125 128.155 89.665 128.525 ;
        RECT 88.185 126.650 88.445 126.970 ;
        RECT 88.245 124.250 88.385 126.650 ;
        RECT 90.085 124.930 90.225 142.290 ;
        RECT 90.545 140.910 90.685 145.010 ;
        RECT 90.945 141.270 91.205 141.590 ;
        RECT 90.485 140.590 90.745 140.910 ;
        RECT 90.485 134.130 90.745 134.450 ;
        RECT 90.545 129.350 90.685 134.130 ;
        RECT 90.485 129.030 90.745 129.350 ;
        RECT 91.005 125.270 91.145 141.270 ;
        RECT 91.465 140.570 91.605 153.170 ;
        RECT 91.925 146.350 92.065 172.130 ;
        RECT 92.325 171.190 92.585 171.510 ;
        RECT 92.385 149.750 92.525 171.190 ;
        RECT 94.225 170.830 94.365 172.210 ;
        RECT 94.165 170.510 94.425 170.830 ;
        RECT 93.245 167.110 93.505 167.430 ;
        RECT 92.785 165.410 93.045 165.730 ;
        RECT 92.845 163.350 92.985 165.410 ;
        RECT 93.305 163.350 93.445 167.110 ;
        RECT 92.785 163.030 93.045 163.350 ;
        RECT 93.245 163.030 93.505 163.350 ;
        RECT 92.785 160.310 93.045 160.630 ;
        RECT 92.845 154.510 92.985 160.310 ;
        RECT 93.245 159.970 93.505 160.290 ;
        RECT 93.305 155.950 93.445 159.970 ;
        RECT 93.705 155.950 93.965 156.210 ;
        RECT 93.305 155.890 93.965 155.950 ;
        RECT 93.305 155.810 93.905 155.890 ;
        RECT 93.305 154.510 93.445 155.810 ;
        RECT 94.225 155.270 94.365 170.510 ;
        RECT 95.145 168.190 95.285 181.390 ;
        RECT 97.905 181.370 98.045 183.090 ;
        RECT 100.665 182.390 100.805 183.090 ;
        RECT 100.605 182.070 100.865 182.390 ;
        RECT 96.465 181.050 96.725 181.370 ;
        RECT 97.845 181.050 98.105 181.370 ;
        RECT 96.005 175.840 96.265 175.930 ;
        RECT 95.605 175.700 96.265 175.840 ;
        RECT 95.605 173.210 95.745 175.700 ;
        RECT 96.005 175.610 96.265 175.700 ;
        RECT 95.545 172.890 95.805 173.210 ;
        RECT 95.605 170.490 95.745 172.890 ;
        RECT 96.525 172.870 96.665 181.050 ;
        RECT 99.910 179.835 101.450 180.205 ;
        RECT 106.185 178.990 106.325 183.770 ;
        RECT 106.125 178.670 106.385 178.990 ;
        RECT 99.685 177.990 99.945 178.310 ;
        RECT 99.225 177.650 99.485 177.970 ;
        RECT 97.385 174.930 97.645 175.250 ;
        RECT 96.465 172.550 96.725 172.870 ;
        RECT 97.445 171.510 97.585 174.930 ;
        RECT 99.285 174.230 99.425 177.650 ;
        RECT 99.745 175.930 99.885 177.990 ;
        RECT 104.285 175.950 104.545 176.270 ;
        RECT 99.685 175.610 99.945 175.930 ;
        RECT 102.905 175.610 103.165 175.930 ;
        RECT 99.910 174.395 101.450 174.765 ;
        RECT 99.225 173.910 99.485 174.230 ;
        RECT 102.965 173.210 103.105 175.610 ;
        RECT 102.905 172.890 103.165 173.210 ;
        RECT 98.305 172.210 98.565 172.530 ;
        RECT 97.385 171.190 97.645 171.510 ;
        RECT 95.545 170.170 95.805 170.490 ;
        RECT 95.605 168.790 95.745 170.170 ;
        RECT 95.545 168.470 95.805 168.790 ;
        RECT 95.145 168.050 95.745 168.190 ;
        RECT 94.625 164.050 94.885 164.370 ;
        RECT 94.685 162.330 94.825 164.050 ;
        RECT 94.625 162.010 94.885 162.330 ;
        RECT 94.625 158.610 94.885 158.930 ;
        RECT 95.085 158.610 95.345 158.930 ;
        RECT 94.685 157.230 94.825 158.610 ;
        RECT 94.625 156.910 94.885 157.230 ;
        RECT 93.765 155.130 94.365 155.270 ;
        RECT 92.785 154.190 93.045 154.510 ;
        RECT 93.245 154.190 93.505 154.510 ;
        RECT 92.845 153.490 92.985 154.190 ;
        RECT 92.785 153.170 93.045 153.490 ;
        RECT 93.245 152.150 93.505 152.470 ;
        RECT 92.785 151.130 93.045 151.450 ;
        RECT 92.325 149.430 92.585 149.750 ;
        RECT 92.845 149.070 92.985 151.130 ;
        RECT 92.785 148.750 93.045 149.070 ;
        RECT 93.305 148.730 93.445 152.150 ;
        RECT 93.765 151.450 93.905 155.130 ;
        RECT 94.165 153.510 94.425 153.830 ;
        RECT 93.705 151.130 93.965 151.450 ;
        RECT 93.705 150.450 93.965 150.770 ;
        RECT 93.245 148.410 93.505 148.730 ;
        RECT 93.245 146.370 93.505 146.690 ;
        RECT 91.865 146.030 92.125 146.350 ;
        RECT 92.315 143.455 92.595 143.825 ;
        RECT 93.305 143.630 93.445 146.370 ;
        RECT 93.765 143.970 93.905 150.450 ;
        RECT 94.225 149.750 94.365 153.510 ;
        RECT 94.625 151.305 94.885 151.450 ;
        RECT 94.615 150.935 94.895 151.305 ;
        RECT 94.165 149.430 94.425 149.750 ;
        RECT 94.685 149.070 94.825 150.935 ;
        RECT 94.165 148.750 94.425 149.070 ;
        RECT 94.625 148.750 94.885 149.070 ;
        RECT 94.225 148.390 94.365 148.750 ;
        RECT 94.165 148.070 94.425 148.390 ;
        RECT 94.625 148.070 94.885 148.390 ;
        RECT 94.225 146.010 94.365 148.070 ;
        RECT 94.165 145.690 94.425 146.010 ;
        RECT 93.705 143.650 93.965 143.970 ;
        RECT 92.325 143.310 92.585 143.455 ;
        RECT 92.785 143.310 93.045 143.630 ;
        RECT 93.245 143.310 93.505 143.630 ;
        RECT 94.165 143.310 94.425 143.630 ;
        RECT 91.865 142.290 92.125 142.610 ;
        RECT 91.405 140.250 91.665 140.570 ;
        RECT 91.405 134.810 91.665 135.130 ;
        RECT 91.465 131.730 91.605 134.810 ;
        RECT 91.405 131.410 91.665 131.730 ;
        RECT 91.465 129.690 91.605 131.410 ;
        RECT 91.405 129.370 91.665 129.690 ;
        RECT 90.945 124.950 91.205 125.270 ;
        RECT 90.025 124.610 90.285 124.930 ;
        RECT 88.185 123.930 88.445 124.250 ;
        RECT 90.025 123.590 90.285 123.910 ;
        RECT 88.125 122.715 89.665 123.085 ;
        RECT 90.085 121.870 90.225 123.590 ;
        RECT 90.025 121.550 90.285 121.870 ;
        RECT 90.085 121.385 90.225 121.550 ;
        RECT 90.015 121.015 90.295 121.385 ;
        RECT 90.085 119.830 90.225 121.015 ;
        RECT 90.025 119.510 90.285 119.830 ;
        RECT 90.485 117.810 90.745 118.130 ;
        RECT 88.125 117.275 89.665 117.645 ;
        RECT 90.545 116.430 90.685 117.810 ;
        RECT 90.485 116.110 90.745 116.430 ;
        RECT 88.125 111.835 89.665 112.205 ;
        RECT 91.925 110.990 92.065 142.290 ;
        RECT 92.385 141.590 92.525 143.310 ;
        RECT 92.325 141.270 92.585 141.590 ;
        RECT 92.385 140.570 92.525 141.270 ;
        RECT 92.845 141.250 92.985 143.310 ;
        RECT 93.705 141.270 93.965 141.590 ;
        RECT 92.785 140.930 93.045 141.250 ;
        RECT 92.325 140.250 92.585 140.570 ;
        RECT 93.245 140.250 93.505 140.570 ;
        RECT 93.305 135.130 93.445 140.250 ;
        RECT 93.245 134.810 93.505 135.130 ;
        RECT 93.305 133.430 93.445 134.810 ;
        RECT 93.245 133.110 93.505 133.430 ;
        RECT 93.765 131.470 93.905 141.270 ;
        RECT 94.225 140.570 94.365 143.310 ;
        RECT 94.165 140.425 94.425 140.570 ;
        RECT 94.155 140.055 94.435 140.425 ;
        RECT 94.685 138.190 94.825 148.070 ;
        RECT 95.145 138.190 95.285 158.610 ;
        RECT 95.605 152.470 95.745 168.050 ;
        RECT 98.365 167.090 98.505 172.210 ;
        RECT 99.225 169.490 99.485 169.810 ;
        RECT 98.305 166.770 98.565 167.090 ;
        RECT 96.465 164.730 96.725 165.050 ;
        RECT 97.845 164.730 98.105 165.050 ;
        RECT 96.005 157.590 96.265 157.910 ;
        RECT 96.065 154.510 96.205 157.590 ;
        RECT 96.525 154.510 96.665 164.730 ;
        RECT 97.905 162.670 98.045 164.730 ;
        RECT 97.845 162.350 98.105 162.670 ;
        RECT 97.905 162.070 98.045 162.350 ;
        RECT 98.365 162.330 98.505 166.770 ;
        RECT 99.285 165.390 99.425 169.490 ;
        RECT 99.910 168.955 101.450 169.325 ;
        RECT 100.145 167.790 100.405 168.110 ;
        RECT 101.065 167.790 101.325 168.110 ;
        RECT 100.205 165.730 100.345 167.790 ;
        RECT 100.605 167.110 100.865 167.430 ;
        RECT 100.145 165.410 100.405 165.730 ;
        RECT 100.665 165.390 100.805 167.110 ;
        RECT 99.225 165.070 99.485 165.390 ;
        RECT 100.605 165.070 100.865 165.390 ;
        RECT 97.445 161.930 98.045 162.070 ;
        RECT 98.305 162.010 98.565 162.330 ;
        RECT 97.445 158.930 97.585 161.930 ;
        RECT 97.845 161.330 98.105 161.650 ;
        RECT 97.905 159.950 98.045 161.330 ;
        RECT 98.365 160.290 98.505 162.010 ;
        RECT 98.305 159.970 98.565 160.290 ;
        RECT 97.845 159.630 98.105 159.950 ;
        RECT 98.765 159.630 99.025 159.950 ;
        RECT 97.385 158.610 97.645 158.930 ;
        RECT 97.445 157.230 97.585 158.610 ;
        RECT 97.385 156.910 97.645 157.230 ;
        RECT 97.905 156.550 98.045 159.630 ;
        RECT 98.825 157.910 98.965 159.630 ;
        RECT 98.765 157.590 99.025 157.910 ;
        RECT 97.845 156.230 98.105 156.550 ;
        RECT 98.305 154.530 98.565 154.850 ;
        RECT 96.005 154.190 96.265 154.510 ;
        RECT 96.465 154.190 96.725 154.510 ;
        RECT 97.845 153.170 98.105 153.490 ;
        RECT 95.545 152.150 95.805 152.470 ;
        RECT 96.465 151.470 96.725 151.790 ;
        RECT 95.545 151.130 95.805 151.450 ;
        RECT 95.605 143.630 95.745 151.130 ;
        RECT 96.005 150.450 96.265 150.770 ;
        RECT 95.545 143.310 95.805 143.630 ;
        RECT 95.545 140.930 95.805 141.250 ;
        RECT 94.625 137.870 94.885 138.190 ;
        RECT 95.085 137.870 95.345 138.190 ;
        RECT 95.605 137.590 95.745 140.930 ;
        RECT 96.065 140.910 96.205 150.450 ;
        RECT 96.525 145.920 96.665 151.470 ;
        RECT 97.905 149.070 98.045 153.170 ;
        RECT 97.385 148.750 97.645 149.070 ;
        RECT 97.845 148.750 98.105 149.070 ;
        RECT 96.925 148.410 97.185 148.730 ;
        RECT 96.985 147.030 97.125 148.410 ;
        RECT 97.445 147.030 97.585 148.750 ;
        RECT 97.845 147.730 98.105 148.050 ;
        RECT 96.925 146.710 97.185 147.030 ;
        RECT 97.385 146.710 97.645 147.030 ;
        RECT 97.385 145.920 97.645 146.010 ;
        RECT 96.525 145.780 97.645 145.920 ;
        RECT 97.385 145.690 97.645 145.780 ;
        RECT 96.925 145.010 97.185 145.330 ;
        RECT 96.985 144.310 97.125 145.010 ;
        RECT 96.925 143.990 97.185 144.310 ;
        RECT 96.985 143.630 97.125 143.990 ;
        RECT 97.445 143.630 97.585 145.690 ;
        RECT 96.925 143.310 97.185 143.630 ;
        RECT 97.385 143.310 97.645 143.630 ;
        RECT 96.465 142.630 96.725 142.950 ;
        RECT 96.005 140.590 96.265 140.910 ;
        RECT 96.005 139.570 96.265 139.890 ;
        RECT 96.065 138.530 96.205 139.570 ;
        RECT 96.005 138.210 96.265 138.530 ;
        RECT 94.685 137.450 95.745 137.590 ;
        RECT 94.165 136.850 94.425 137.170 ;
        RECT 92.845 131.330 93.905 131.470 ;
        RECT 92.845 125.270 92.985 131.330 ;
        RECT 94.225 130.620 94.365 136.850 ;
        RECT 93.305 130.480 94.365 130.620 ;
        RECT 92.785 124.950 93.045 125.270 ;
        RECT 93.305 124.930 93.445 130.480 ;
        RECT 93.245 124.610 93.505 124.930 ;
        RECT 93.705 121.550 93.965 121.870 ;
        RECT 93.765 121.190 93.905 121.550 ;
        RECT 93.705 120.870 93.965 121.190 ;
        RECT 94.165 120.870 94.425 121.190 ;
        RECT 93.245 120.530 93.505 120.850 ;
        RECT 93.305 118.470 93.445 120.530 ;
        RECT 93.245 118.150 93.505 118.470 ;
        RECT 92.325 117.810 92.585 118.130 ;
        RECT 92.385 115.410 92.525 117.810 ;
        RECT 94.225 116.770 94.365 120.870 ;
        RECT 94.165 116.450 94.425 116.770 ;
        RECT 92.325 115.090 92.585 115.410 ;
        RECT 92.385 111.670 92.525 115.090 ;
        RECT 92.325 111.350 92.585 111.670 ;
        RECT 94.685 110.990 94.825 137.450 ;
        RECT 95.545 136.850 95.805 137.170 ;
        RECT 95.085 124.610 95.345 124.930 ;
        RECT 95.145 121.530 95.285 124.610 ;
        RECT 95.085 121.210 95.345 121.530 ;
        RECT 95.085 120.530 95.345 120.850 ;
        RECT 95.145 119.150 95.285 120.530 ;
        RECT 95.085 118.830 95.345 119.150 ;
        RECT 87.725 110.670 87.985 110.990 ;
        RECT 91.865 110.670 92.125 110.990 ;
        RECT 94.625 110.670 94.885 110.990 ;
        RECT 78.065 110.330 78.325 110.650 ;
        RECT 87.265 110.330 87.525 110.650 ;
        RECT 74.845 109.650 75.105 109.970 ;
        RECT 75.765 109.650 76.025 109.970 ;
        RECT 73.925 108.630 74.185 108.950 ;
        RECT 73.465 107.270 73.725 107.590 ;
        RECT 73.525 106.230 73.665 107.270 ;
        RECT 72.085 105.910 72.345 106.230 ;
        RECT 73.465 105.910 73.725 106.230 ;
        RECT 71.625 105.570 71.885 105.890 ;
        RECT 71.165 103.190 71.425 103.510 ;
        RECT 72.145 98.340 72.285 105.910 ;
        RECT 72.545 105.230 72.805 105.550 ;
        RECT 72.605 103.510 72.745 105.230 ;
        RECT 73.985 105.210 74.125 108.630 ;
        RECT 74.905 106.230 75.045 109.650 ;
        RECT 74.845 105.910 75.105 106.230 ;
        RECT 73.925 104.890 74.185 105.210 ;
        RECT 72.545 103.190 72.805 103.510 ;
        RECT 75.825 102.150 75.965 109.650 ;
        RECT 76.335 109.115 77.875 109.485 ;
        RECT 76.335 103.675 77.875 104.045 ;
        RECT 76.685 102.510 76.945 102.830 ;
        RECT 75.765 101.830 76.025 102.150 ;
        RECT 76.745 98.340 76.885 102.510 ;
        RECT 78.125 101.810 78.265 110.330 ;
        RECT 80.365 109.650 80.625 109.970 ;
        RECT 84.045 109.650 84.305 109.970 ;
        RECT 93.245 109.650 93.505 109.970 ;
        RECT 79.445 107.270 79.705 107.590 ;
        RECT 79.505 103.510 79.645 107.270 ;
        RECT 79.445 103.190 79.705 103.510 ;
        RECT 80.425 102.830 80.565 109.650 ;
        RECT 84.105 108.270 84.245 109.650 ;
        RECT 81.285 107.950 81.545 108.270 ;
        RECT 84.045 107.950 84.305 108.270 ;
        RECT 90.485 107.950 90.745 108.270 ;
        RECT 80.365 102.510 80.625 102.830 ;
        RECT 78.065 101.490 78.325 101.810 ;
        RECT 81.345 98.340 81.485 107.950 ;
        RECT 88.125 106.395 89.665 106.765 ;
        RECT 87.725 105.230 87.985 105.550 ;
        RECT 84.045 104.890 84.305 105.210 ;
        RECT 85.885 104.890 86.145 105.210 ;
        RECT 84.105 102.830 84.245 104.890 ;
        RECT 84.045 102.510 84.305 102.830 ;
        RECT 85.945 98.340 86.085 104.890 ;
        RECT 87.785 103.510 87.925 105.230 ;
        RECT 87.725 103.190 87.985 103.510 ;
        RECT 88.125 100.955 89.665 101.325 ;
        RECT 90.545 98.340 90.685 107.950 ;
        RECT 93.305 105.890 93.445 109.650 ;
        RECT 95.605 108.950 95.745 136.850 ;
        RECT 96.525 127.310 96.665 142.630 ;
        RECT 97.445 140.570 97.585 143.310 ;
        RECT 97.385 140.250 97.645 140.570 ;
        RECT 97.375 138.695 97.655 139.065 ;
        RECT 97.445 138.530 97.585 138.695 ;
        RECT 97.385 138.210 97.645 138.530 ;
        RECT 96.925 137.530 97.185 137.850 ;
        RECT 96.985 131.730 97.125 137.530 ;
        RECT 97.385 132.090 97.645 132.410 ;
        RECT 96.925 131.410 97.185 131.730 ;
        RECT 97.445 129.690 97.585 132.090 ;
        RECT 97.385 129.370 97.645 129.690 ;
        RECT 96.465 126.990 96.725 127.310 ;
        RECT 96.005 126.650 96.265 126.970 ;
        RECT 96.065 124.250 96.205 126.650 ;
        RECT 96.465 126.310 96.725 126.630 ;
        RECT 96.005 123.930 96.265 124.250 ;
        RECT 96.065 119.830 96.205 123.930 ;
        RECT 96.525 123.570 96.665 126.310 ;
        RECT 96.925 123.590 97.185 123.910 ;
        RECT 96.465 123.250 96.725 123.570 ;
        RECT 96.525 122.550 96.665 123.250 ;
        RECT 96.985 122.550 97.125 123.590 ;
        RECT 96.465 122.230 96.725 122.550 ;
        RECT 96.925 122.230 97.185 122.550 ;
        RECT 96.925 121.210 97.185 121.530 ;
        RECT 96.005 119.510 96.265 119.830 ;
        RECT 96.985 118.470 97.125 121.210 ;
        RECT 97.445 119.150 97.585 129.370 ;
        RECT 97.905 126.630 98.045 147.730 ;
        RECT 98.365 144.310 98.505 154.530 ;
        RECT 98.825 154.170 98.965 157.590 ;
        RECT 99.285 154.850 99.425 165.070 ;
        RECT 101.125 165.050 101.265 167.790 ;
        RECT 103.825 167.450 104.085 167.770 ;
        RECT 103.885 166.070 104.025 167.450 ;
        RECT 103.825 165.750 104.085 166.070 ;
        RECT 104.345 165.390 104.485 175.950 ;
        RECT 104.745 175.610 105.005 175.930 ;
        RECT 104.805 171.170 104.945 175.610 ;
        RECT 135.630 173.380 136.780 174.600 ;
        RECT 109.805 172.890 110.065 173.210 ;
        RECT 108.425 172.550 108.685 172.870 ;
        RECT 108.485 171.510 108.625 172.550 ;
        RECT 108.425 171.190 108.685 171.510 ;
        RECT 104.745 170.850 105.005 171.170 ;
        RECT 107.965 170.850 108.225 171.170 ;
        RECT 108.025 168.790 108.165 170.850 ;
        RECT 109.865 170.490 110.005 172.890 ;
        RECT 110.725 170.510 110.985 170.830 ;
        RECT 109.805 170.170 110.065 170.490 ;
        RECT 107.965 168.470 108.225 168.790 ;
        RECT 104.285 165.070 104.545 165.390 ;
        RECT 106.585 165.070 106.845 165.390 ;
        RECT 101.065 164.730 101.325 165.050 ;
        RECT 102.905 164.050 103.165 164.370 ;
        RECT 99.910 163.515 101.450 163.885 ;
        RECT 102.965 162.330 103.105 164.050 ;
        RECT 106.645 163.350 106.785 165.070 ;
        RECT 108.425 164.050 108.685 164.370 ;
        RECT 106.585 163.030 106.845 163.350 ;
        RECT 108.485 162.670 108.625 164.050 ;
        RECT 109.865 162.670 110.005 170.170 ;
        RECT 110.785 168.450 110.925 170.510 ;
        RECT 133.750 170.070 134.880 172.730 ;
        RECT 110.725 168.130 110.985 168.450 ;
        RECT 135.630 166.640 136.740 173.380 ;
        RECT 135.630 165.420 136.780 166.640 ;
        RECT 108.425 162.350 108.685 162.670 ;
        RECT 109.805 162.350 110.065 162.670 ;
        RECT 102.905 162.010 103.165 162.330 ;
        RECT 101.985 159.630 102.245 159.950 ;
        RECT 104.285 159.630 104.545 159.950 ;
        RECT 99.910 158.075 101.450 158.445 ;
        RECT 101.065 155.890 101.325 156.210 ;
        RECT 99.225 154.530 99.485 154.850 ;
        RECT 98.765 153.850 99.025 154.170 ;
        RECT 101.125 153.910 101.265 155.890 ;
        RECT 102.045 155.190 102.185 159.630 ;
        RECT 102.905 158.610 103.165 158.930 ;
        RECT 101.985 154.870 102.245 155.190 ;
        RECT 101.985 154.190 102.245 154.510 ;
        RECT 102.445 154.190 102.705 154.510 ;
        RECT 101.125 153.830 101.725 153.910 ;
        RECT 101.125 153.770 101.785 153.830 ;
        RECT 101.525 153.510 101.785 153.770 ;
        RECT 99.910 152.635 101.450 153.005 ;
        RECT 98.765 151.130 99.025 151.450 ;
        RECT 98.825 145.670 98.965 151.130 ;
        RECT 99.225 150.450 99.485 150.770 ;
        RECT 98.765 145.350 99.025 145.670 ;
        RECT 98.305 143.990 98.565 144.310 ;
        RECT 99.285 143.970 99.425 150.450 ;
        RECT 102.045 149.070 102.185 154.190 ;
        RECT 102.505 154.025 102.645 154.190 ;
        RECT 102.435 153.655 102.715 154.025 ;
        RECT 101.985 148.750 102.245 149.070 ;
        RECT 99.675 148.215 99.955 148.585 ;
        RECT 99.685 148.070 99.945 148.215 ;
        RECT 99.910 147.195 101.450 147.565 ;
        RECT 100.605 145.690 100.865 146.010 ;
        RECT 99.225 143.650 99.485 143.970 ;
        RECT 100.665 143.200 100.805 145.690 ;
        RECT 99.285 143.060 100.805 143.200 ;
        RECT 98.765 142.290 99.025 142.610 ;
        RECT 98.825 140.230 98.965 142.290 ;
        RECT 99.285 140.570 99.425 143.060 ;
        RECT 102.445 142.970 102.705 143.290 ;
        RECT 99.910 141.755 101.450 142.125 ;
        RECT 99.225 140.425 99.485 140.570 ;
        RECT 98.765 139.910 99.025 140.230 ;
        RECT 99.215 140.055 99.495 140.425 ;
        RECT 102.505 140.230 102.645 142.970 ;
        RECT 102.965 140.570 103.105 158.610 ;
        RECT 104.345 154.850 104.485 159.630 ;
        RECT 105.665 158.950 105.925 159.270 ;
        RECT 104.745 158.610 105.005 158.930 ;
        RECT 104.805 156.550 104.945 158.610 ;
        RECT 104.745 156.230 105.005 156.550 ;
        RECT 104.285 154.530 104.545 154.850 ;
        RECT 105.725 154.510 105.865 158.950 ;
        RECT 109.865 156.890 110.005 162.350 ;
        RECT 111.185 159.630 111.445 159.950 ;
        RECT 111.245 159.465 111.385 159.630 ;
        RECT 111.175 159.095 111.455 159.465 ;
        RECT 108.425 156.570 108.685 156.890 ;
        RECT 109.805 156.570 110.065 156.890 ;
        RECT 105.665 154.190 105.925 154.510 ;
        RECT 108.485 153.830 108.625 156.570 ;
        RECT 109.865 155.270 110.005 156.570 ;
        RECT 109.865 155.130 110.465 155.270 ;
        RECT 108.425 153.510 108.685 153.830 ;
        RECT 110.325 151.790 110.465 155.130 ;
        RECT 110.265 151.470 110.525 151.790 ;
        RECT 106.125 150.790 106.385 151.110 ;
        RECT 108.885 150.790 109.145 151.110 ;
        RECT 104.285 150.450 104.545 150.770 ;
        RECT 103.825 147.730 104.085 148.050 ;
        RECT 103.365 146.370 103.625 146.690 ;
        RECT 103.425 143.290 103.565 146.370 ;
        RECT 103.885 145.670 104.025 147.730 ;
        RECT 103.825 145.350 104.085 145.670 ;
        RECT 103.885 143.710 104.025 145.350 ;
        RECT 104.345 145.330 104.485 150.450 ;
        RECT 104.745 148.750 105.005 149.070 ;
        RECT 104.805 146.010 104.945 148.750 ;
        RECT 106.185 147.030 106.325 150.790 ;
        RECT 108.945 147.030 109.085 150.790 ;
        RECT 110.325 149.070 110.465 151.470 ;
        RECT 110.265 148.750 110.525 149.070 ;
        RECT 109.345 148.410 109.605 148.730 ;
        RECT 109.405 147.030 109.545 148.410 ;
        RECT 106.125 146.710 106.385 147.030 ;
        RECT 108.885 146.710 109.145 147.030 ;
        RECT 109.345 146.710 109.605 147.030 ;
        RECT 104.745 145.690 105.005 146.010 ;
        RECT 106.585 145.690 106.845 146.010 ;
        RECT 108.425 145.690 108.685 146.010 ;
        RECT 104.285 145.010 104.545 145.330 ;
        RECT 104.345 144.310 104.485 145.010 ;
        RECT 104.285 143.990 104.545 144.310 ;
        RECT 103.885 143.570 104.485 143.710 ;
        RECT 104.345 143.290 104.485 143.570 ;
        RECT 103.365 142.970 103.625 143.290 ;
        RECT 104.285 142.970 104.545 143.290 ;
        RECT 103.425 140.910 103.565 142.970 ;
        RECT 103.365 140.590 103.625 140.910 ;
        RECT 102.905 140.250 103.165 140.570 ;
        RECT 102.445 139.910 102.705 140.230 ;
        RECT 102.505 138.870 102.645 139.910 ;
        RECT 102.905 139.570 103.165 139.890 ;
        RECT 102.445 138.550 102.705 138.870 ;
        RECT 99.910 136.315 101.450 136.685 ;
        RECT 101.985 135.490 102.245 135.810 ;
        RECT 98.765 134.130 99.025 134.450 ;
        RECT 99.225 134.130 99.485 134.450 ;
        RECT 98.305 132.430 98.565 132.750 ;
        RECT 98.365 130.710 98.505 132.430 ;
        RECT 98.305 130.390 98.565 130.710 ;
        RECT 98.825 129.690 98.965 134.130 ;
        RECT 99.285 129.690 99.425 134.130 ;
        RECT 100.605 132.430 100.865 132.750 ;
        RECT 100.665 131.730 100.805 132.430 ;
        RECT 102.045 132.410 102.185 135.490 ;
        RECT 102.505 132.830 102.645 138.550 ;
        RECT 102.965 135.470 103.105 139.570 ;
        RECT 103.425 135.810 103.565 140.590 ;
        RECT 104.345 140.570 104.485 142.970 ;
        RECT 106.125 142.290 106.385 142.610 ;
        RECT 104.285 140.250 104.545 140.570 ;
        RECT 104.745 140.250 105.005 140.570 ;
        RECT 104.805 138.190 104.945 140.250 ;
        RECT 104.745 137.870 105.005 138.190 ;
        RECT 103.365 135.490 103.625 135.810 ;
        RECT 102.905 135.150 103.165 135.470 ;
        RECT 102.965 133.430 103.105 135.150 ;
        RECT 102.905 133.110 103.165 133.430 ;
        RECT 102.505 132.750 103.105 132.830 ;
        RECT 102.505 132.690 103.165 132.750 ;
        RECT 102.905 132.430 103.165 132.690 ;
        RECT 101.985 132.090 102.245 132.410 ;
        RECT 100.605 131.410 100.865 131.730 ;
        RECT 105.665 131.410 105.925 131.730 ;
        RECT 99.910 130.875 101.450 131.245 ;
        RECT 98.765 129.370 99.025 129.690 ;
        RECT 99.225 129.370 99.485 129.690 ;
        RECT 105.725 127.310 105.865 131.410 ;
        RECT 105.665 126.990 105.925 127.310 ;
        RECT 97.845 126.310 98.105 126.630 ;
        RECT 105.205 125.970 105.465 126.290 ;
        RECT 99.910 125.435 101.450 125.805 ;
        RECT 97.845 124.270 98.105 124.590 ;
        RECT 97.385 118.830 97.645 119.150 ;
        RECT 96.925 118.150 97.185 118.470 ;
        RECT 97.445 116.430 97.585 118.830 ;
        RECT 97.905 118.130 98.045 124.270 ;
        RECT 105.265 123.910 105.405 125.970 ;
        RECT 105.205 123.590 105.465 123.910 ;
        RECT 99.225 122.230 99.485 122.550 ;
        RECT 98.765 120.530 99.025 120.850 ;
        RECT 98.825 118.470 98.965 120.530 ;
        RECT 99.285 119.150 99.425 122.230 ;
        RECT 105.725 121.530 105.865 126.990 ;
        RECT 102.895 121.015 103.175 121.385 ;
        RECT 105.665 121.210 105.925 121.530 ;
        RECT 99.910 119.995 101.450 120.365 ;
        RECT 100.605 119.510 100.865 119.830 ;
        RECT 99.225 118.830 99.485 119.150 ;
        RECT 98.765 118.150 99.025 118.470 ;
        RECT 97.845 117.810 98.105 118.130 ;
        RECT 100.665 117.110 100.805 119.510 ;
        RECT 102.965 119.150 103.105 121.015 ;
        RECT 102.905 118.830 103.165 119.150 ;
        RECT 105.725 118.810 105.865 121.210 ;
        RECT 106.185 119.230 106.325 142.290 ;
        RECT 106.645 140.570 106.785 145.690 ;
        RECT 108.485 144.310 108.625 145.690 ;
        RECT 108.425 143.990 108.685 144.310 ;
        RECT 135.630 141.200 136.780 141.270 ;
        RECT 106.585 140.250 106.845 140.570 ;
        RECT 135.630 140.180 136.800 141.200 ;
        RECT 106.585 139.570 106.845 139.890 ;
        RECT 108.885 139.570 109.145 139.890 ;
        RECT 106.645 134.790 106.785 139.570 ;
        RECT 108.945 138.190 109.085 139.570 ;
        RECT 108.885 137.870 109.145 138.190 ;
        RECT 132.560 138.140 135.160 140.060 ;
        RECT 110.725 137.530 110.985 137.850 ;
        RECT 110.785 135.130 110.925 137.530 ;
        RECT 108.425 134.810 108.685 135.130 ;
        RECT 108.885 134.810 109.145 135.130 ;
        RECT 110.725 134.810 110.985 135.130 ;
        RECT 106.585 134.470 106.845 134.790 ;
        RECT 108.485 133.430 108.625 134.810 ;
        RECT 108.425 133.110 108.685 133.430 ;
        RECT 108.945 133.090 109.085 134.810 ;
        RECT 135.640 133.320 136.800 140.180 ;
        RECT 108.885 132.770 109.145 133.090 ;
        RECT 107.045 126.990 107.305 127.310 ;
        RECT 107.105 125.270 107.245 126.990 ;
        RECT 107.965 125.970 108.225 126.290 ;
        RECT 107.045 124.950 107.305 125.270 ;
        RECT 108.025 124.590 108.165 125.970 ;
        RECT 107.965 124.270 108.225 124.590 ;
        RECT 108.945 124.160 109.085 132.770 ;
        RECT 109.345 124.160 109.605 124.250 ;
        RECT 108.945 124.020 109.605 124.160 ;
        RECT 106.585 121.890 106.845 122.210 ;
        RECT 106.645 119.830 106.785 121.890 ;
        RECT 108.945 121.870 109.085 124.020 ;
        RECT 109.345 123.930 109.605 124.020 ;
        RECT 108.885 121.550 109.145 121.870 ;
        RECT 110.725 121.550 110.985 121.870 ;
        RECT 108.425 121.210 108.685 121.530 ;
        RECT 108.485 119.830 108.625 121.210 ;
        RECT 106.585 119.510 106.845 119.830 ;
        RECT 108.425 119.510 108.685 119.830 ;
        RECT 106.185 119.090 106.785 119.230 ;
        RECT 105.665 118.490 105.925 118.810 ;
        RECT 101.065 117.810 101.325 118.130 ;
        RECT 100.605 116.790 100.865 117.110 ;
        RECT 101.125 116.430 101.265 117.810 ;
        RECT 104.745 116.450 105.005 116.770 ;
        RECT 97.385 116.110 97.645 116.430 ;
        RECT 101.065 116.110 101.325 116.430 ;
        RECT 97.445 114.050 97.585 116.110 ;
        RECT 99.910 114.555 101.450 114.925 ;
        RECT 104.805 114.390 104.945 116.450 ;
        RECT 104.745 114.070 105.005 114.390 ;
        RECT 97.385 113.790 97.645 114.050 ;
        RECT 97.385 113.730 98.045 113.790 ;
        RECT 97.445 113.650 98.045 113.730 ;
        RECT 96.925 113.050 97.185 113.370 ;
        RECT 96.985 111.670 97.125 113.050 ;
        RECT 96.925 111.350 97.185 111.670 ;
        RECT 97.385 109.650 97.645 109.970 ;
        RECT 95.545 108.630 95.805 108.950 ;
        RECT 94.165 107.270 94.425 107.590 ;
        RECT 94.225 106.230 94.365 107.270 ;
        RECT 94.165 105.910 94.425 106.230 ;
        RECT 93.245 105.570 93.505 105.890 ;
        RECT 95.085 105.230 95.345 105.550 ;
        RECT 95.145 103.510 95.285 105.230 ;
        RECT 96.925 104.210 97.185 104.530 ;
        RECT 95.085 103.190 95.345 103.510 ;
        RECT 95.085 102.510 95.345 102.830 ;
        RECT 95.145 98.340 95.285 102.510 ;
        RECT 96.985 102.150 97.125 104.210 ;
        RECT 97.445 102.830 97.585 109.650 ;
        RECT 97.905 108.270 98.045 113.650 ;
        RECT 105.725 113.370 105.865 118.490 ;
        RECT 106.125 117.810 106.385 118.130 ;
        RECT 106.185 113.370 106.325 117.810 ;
        RECT 105.665 113.050 105.925 113.370 ;
        RECT 106.125 113.050 106.385 113.370 ;
        RECT 101.055 111.495 101.335 111.865 ;
        RECT 101.125 110.990 101.265 111.495 ;
        RECT 106.645 110.990 106.785 119.090 ;
        RECT 110.785 116.430 110.925 121.550 ;
        RECT 110.725 116.110 110.985 116.430 ;
        RECT 108.885 115.770 109.145 116.090 ;
        RECT 108.945 112.690 109.085 115.770 ;
        RECT 108.885 112.370 109.145 112.690 ;
        RECT 109.795 112.175 110.075 112.545 ;
        RECT 109.865 111.670 110.005 112.175 ;
        RECT 109.805 111.350 110.065 111.670 ;
        RECT 101.065 110.670 101.325 110.990 ;
        RECT 106.585 110.670 106.845 110.990 ;
        RECT 110.725 110.670 110.985 110.990 ;
        RECT 110.785 110.505 110.925 110.670 ;
        RECT 98.305 109.990 98.565 110.310 ;
        RECT 108.425 109.990 108.685 110.310 ;
        RECT 110.715 110.135 110.995 110.505 ;
        RECT 97.845 107.950 98.105 108.270 ;
        RECT 97.905 107.250 98.045 107.950 ;
        RECT 97.845 106.930 98.105 107.250 ;
        RECT 97.905 106.230 98.045 106.930 ;
        RECT 97.845 105.910 98.105 106.230 ;
        RECT 98.365 105.630 98.505 109.990 ;
        RECT 103.365 109.650 103.625 109.970 ;
        RECT 104.285 109.650 104.545 109.970 ;
        RECT 105.205 109.650 105.465 109.970 ;
        RECT 107.505 109.650 107.765 109.970 ;
        RECT 99.910 109.115 101.450 109.485 ;
        RECT 102.905 107.270 103.165 107.590 ;
        RECT 97.905 105.550 98.505 105.630 ;
        RECT 98.765 105.570 99.025 105.890 ;
        RECT 97.845 105.490 98.505 105.550 ;
        RECT 97.845 105.230 98.105 105.490 ;
        RECT 98.825 102.830 98.965 105.570 ;
        RECT 99.225 104.890 99.485 105.210 ;
        RECT 97.385 102.510 97.645 102.830 ;
        RECT 98.765 102.510 99.025 102.830 ;
        RECT 96.925 101.830 97.185 102.150 ;
        RECT 99.285 102.060 99.425 104.890 ;
        RECT 99.910 103.675 101.450 104.045 ;
        RECT 99.285 101.920 99.885 102.060 ;
        RECT 99.745 98.340 99.885 101.920 ;
        RECT 21.475 96.340 21.755 98.340 ;
        RECT 26.075 96.340 26.355 98.340 ;
        RECT 30.675 96.340 30.955 98.340 ;
        RECT 35.275 96.340 35.555 98.340 ;
        RECT 39.875 96.340 40.155 98.340 ;
        RECT 44.475 96.340 44.755 98.340 ;
        RECT 49.075 96.340 49.355 98.340 ;
        RECT 53.675 96.340 53.955 98.340 ;
        RECT 58.275 96.340 58.555 98.340 ;
        RECT 62.875 96.340 63.155 98.340 ;
        RECT 67.475 96.340 67.755 98.340 ;
        RECT 72.075 96.340 72.355 98.340 ;
        RECT 76.675 96.340 76.955 98.340 ;
        RECT 81.275 96.340 81.555 98.340 ;
        RECT 85.875 96.340 86.155 98.340 ;
        RECT 90.475 96.340 90.755 98.340 ;
        RECT 95.075 96.340 95.355 98.340 ;
        RECT 99.675 96.340 99.955 98.340 ;
        RECT 102.965 98.150 103.105 107.270 ;
        RECT 103.425 102.150 103.565 109.650 ;
        RECT 104.345 107.590 104.485 109.650 ;
        RECT 104.285 107.270 104.545 107.590 ;
        RECT 105.265 102.830 105.405 109.650 ;
        RECT 107.565 108.270 107.705 109.650 ;
        RECT 107.505 107.950 107.765 108.270 ;
        RECT 108.485 105.890 108.625 109.990 ;
        RECT 109.805 106.930 110.065 107.250 ;
        RECT 108.425 105.570 108.685 105.890 ;
        RECT 109.865 105.550 110.005 106.930 ;
        RECT 129.750 105.580 133.160 106.650 ;
        RECT 109.805 105.230 110.065 105.550 ;
        RECT 105.205 102.510 105.465 102.830 ;
        RECT 103.365 101.830 103.625 102.150 ;
        RECT 108.885 101.830 109.145 102.150 ;
        RECT 103.885 98.690 104.485 98.830 ;
        RECT 103.885 98.150 104.025 98.690 ;
        RECT 104.345 98.340 104.485 98.690 ;
        RECT 108.945 98.340 109.085 101.830 ;
        RECT 102.965 98.010 104.025 98.150 ;
        RECT 104.275 96.340 104.555 98.340 ;
        RECT 108.875 96.340 109.155 98.340 ;
        RECT 13.920 85.550 15.140 89.420 ;
        RECT 19.910 85.980 21.130 89.850 ;
        RECT 67.730 89.640 68.670 89.840 ;
        RECT 25.730 85.120 26.950 88.990 ;
        RECT 31.780 85.510 33.000 89.380 ;
        RECT 37.750 88.780 38.970 89.290 ;
        RECT 37.680 88.620 38.970 88.780 ;
        RECT 43.810 88.630 45.030 89.530 ;
        RECT 49.740 88.640 50.960 89.040 ;
        RECT 37.680 86.810 39.070 88.620 ;
        RECT 37.750 85.420 38.970 86.810 ;
        RECT 43.810 86.720 45.140 88.630 ;
        RECT 49.740 86.920 51.010 88.640 ;
        RECT 43.810 85.660 45.030 86.720 ;
        RECT 49.740 85.170 50.960 86.920 ;
        RECT 55.530 85.320 56.750 89.190 ;
        RECT 61.720 88.640 62.940 88.870 ;
        RECT 61.720 86.600 63.130 88.640 ;
        RECT 61.720 85.000 62.940 86.600 ;
        RECT 67.580 85.770 68.800 89.640 ;
        RECT 73.850 84.290 75.070 88.160 ;
        RECT 79.730 84.310 80.950 88.180 ;
        RECT 74.090 80.440 74.370 84.290 ;
        RECT 20.140 80.160 74.370 80.440 ;
        RECT 20.140 75.650 20.420 80.160 ;
        RECT 80.070 79.800 80.350 84.310 ;
        RECT 85.470 84.100 86.690 87.970 ;
        RECT 91.460 84.500 92.680 88.320 ;
        RECT 97.600 84.630 98.820 88.240 ;
        RECT 103.650 84.740 104.870 88.610 ;
        RECT 109.620 85.420 110.840 89.290 ;
        RECT 115.740 85.700 116.960 89.570 ;
        RECT 121.520 85.700 122.740 89.570 ;
        RECT 31.380 79.520 80.350 79.800 ;
        RECT 31.380 75.850 31.660 79.520 ;
        RECT 86.050 79.170 86.330 84.100 ;
        RECT 42.510 78.890 86.330 79.170 ;
        RECT 3.960 71.320 6.050 73.240 ;
        RECT 19.330 73.120 21.890 75.650 ;
        RECT 28.185 73.180 30.255 74.460 ;
        RECT 30.670 73.320 33.230 75.850 ;
        RECT 42.510 75.750 42.790 78.890 ;
        RECT 92.030 78.570 92.310 84.500 ;
        RECT 53.830 78.290 92.310 78.570 ;
        RECT 53.830 75.820 54.110 78.290 ;
        RECT 98.010 77.990 98.290 84.630 ;
        RECT 64.900 77.710 98.290 77.990 ;
        RECT 19.005 71.800 19.865 72.640 ;
        RECT 15.560 68.610 16.990 71.210 ;
        RECT 19.305 68.570 19.845 71.800 ;
        RECT 20.145 70.600 20.555 73.120 ;
        RECT 30.205 71.810 31.065 72.650 ;
        RECT 19.325 47.770 19.825 68.570 ;
        RECT 20.165 49.090 20.555 70.600 ;
        RECT 20.955 70.010 21.845 70.740 ;
        RECT 21.055 65.190 21.315 70.010 ;
        RECT 22.695 68.620 25.405 69.470 ;
        RECT 22.895 65.840 24.825 68.620 ;
        RECT 30.505 68.580 31.045 71.810 ;
        RECT 31.345 70.610 31.755 73.320 ;
        RECT 39.475 73.150 41.545 74.430 ;
        RECT 41.910 73.220 44.470 75.750 ;
        RECT 41.425 71.780 42.285 72.620 ;
        RECT 27.795 67.130 28.915 67.810 ;
        RECT 28.075 65.850 28.745 67.130 ;
        RECT 21.455 65.460 26.505 65.840 ;
        RECT 27.865 65.440 28.915 65.850 ;
        RECT 21.055 63.640 21.435 65.190 ;
        RECT 21.175 55.800 21.435 63.640 ;
        RECT 26.485 63.200 26.755 65.240 ;
        RECT 27.615 63.200 27.885 65.200 ;
        RECT 26.485 56.510 27.885 63.200 ;
        RECT 21.085 55.290 21.445 55.800 ;
        RECT 21.065 54.860 21.445 55.290 ;
        RECT 26.485 55.190 26.755 56.510 ;
        RECT 27.615 55.150 27.885 56.510 ;
        RECT 28.885 55.260 29.205 65.190 ;
        RECT 28.885 55.200 29.215 55.260 ;
        RECT 21.065 54.580 21.315 54.860 ;
        RECT 20.865 54.180 25.505 54.580 ;
        RECT 26.405 54.290 27.535 54.300 ;
        RECT 28.895 54.290 29.215 55.200 ;
        RECT 21.065 52.060 21.315 54.180 ;
        RECT 25.765 53.490 26.125 54.110 ;
        RECT 25.845 52.610 26.105 53.490 ;
        RECT 26.385 53.240 29.215 54.290 ;
        RECT 25.675 52.230 26.205 52.610 ;
        RECT 21.065 51.970 21.565 52.060 ;
        RECT 21.055 51.240 21.565 51.970 ;
        RECT 21.295 50.240 21.565 51.240 ;
        RECT 22.205 50.990 22.475 51.940 ;
        RECT 22.205 50.840 22.675 50.990 ;
        RECT 22.205 50.160 22.765 50.840 ;
        RECT 22.285 50.150 22.765 50.160 ;
        RECT 21.575 49.620 22.195 49.980 ;
        RECT 21.615 49.090 22.045 49.620 ;
        RECT 20.165 48.670 22.045 49.090 ;
        RECT 22.535 48.960 22.765 50.150 ;
        RECT 21.615 47.800 22.045 48.670 ;
        RECT 22.455 48.360 22.835 48.960 ;
        RECT 19.325 47.060 20.015 47.770 ;
        RECT 21.435 47.440 22.055 47.800 ;
        RECT 21.135 47.060 21.425 47.250 ;
        RECT 19.325 46.620 21.425 47.060 ;
        RECT 19.325 46.600 20.015 46.620 ;
        RECT 21.135 46.380 21.425 46.620 ;
        RECT 22.055 46.990 22.325 47.240 ;
        RECT 22.535 46.990 22.765 48.360 ;
        RECT 25.355 47.010 25.685 52.030 ;
        RECT 26.405 52.020 27.535 53.240 ;
        RECT 28.895 53.220 29.215 53.240 ;
        RECT 22.055 46.880 22.765 46.990 ;
        RECT 25.345 46.960 25.685 47.010 ;
        RECT 26.235 47.780 27.615 52.020 ;
        RECT 22.055 46.570 22.715 46.880 ;
        RECT 22.055 46.400 22.325 46.570 ;
        RECT 25.345 45.000 25.625 46.960 ;
        RECT 26.235 46.920 26.535 47.780 ;
        RECT 27.315 46.920 27.615 47.780 ;
        RECT 28.165 46.920 28.495 51.990 ;
        RECT 27.565 46.380 28.045 46.760 ;
        RECT 27.665 45.760 27.915 46.380 ;
        RECT 27.565 45.160 27.945 45.760 ;
        RECT 24.825 44.230 25.925 45.000 ;
        RECT 28.215 44.930 28.495 46.920 ;
        RECT 30.525 47.780 31.025 68.580 ;
        RECT 31.365 49.100 31.755 70.610 ;
        RECT 32.155 70.020 33.045 70.750 ;
        RECT 32.255 65.200 32.515 70.020 ;
        RECT 33.895 68.630 36.605 69.480 ;
        RECT 34.095 65.850 36.025 68.630 ;
        RECT 41.725 68.550 42.265 71.780 ;
        RECT 42.565 70.580 42.975 73.220 ;
        RECT 50.055 73.090 52.125 74.370 ;
        RECT 53.150 73.290 55.710 75.820 ;
        RECT 64.900 75.810 65.180 77.710 ;
        RECT 103.990 77.230 104.270 84.740 ;
        RECT 76.140 76.950 104.270 77.230 ;
        RECT 52.675 71.760 53.535 72.600 ;
        RECT 38.995 67.140 40.115 67.820 ;
        RECT 39.275 65.860 39.945 67.140 ;
        RECT 32.655 65.470 37.705 65.850 ;
        RECT 39.065 65.450 40.115 65.860 ;
        RECT 32.255 63.650 32.635 65.200 ;
        RECT 32.375 55.810 32.635 63.650 ;
        RECT 37.685 63.210 37.955 65.250 ;
        RECT 38.815 63.210 39.085 65.210 ;
        RECT 37.685 56.520 39.085 63.210 ;
        RECT 32.285 55.300 32.645 55.810 ;
        RECT 32.265 54.870 32.645 55.300 ;
        RECT 37.685 55.200 37.955 56.520 ;
        RECT 38.815 55.160 39.085 56.520 ;
        RECT 40.085 55.270 40.405 65.200 ;
        RECT 40.085 55.210 40.415 55.270 ;
        RECT 32.265 54.590 32.515 54.870 ;
        RECT 32.065 54.190 36.705 54.590 ;
        RECT 37.605 54.300 38.735 54.310 ;
        RECT 40.095 54.300 40.415 55.210 ;
        RECT 32.265 52.070 32.515 54.190 ;
        RECT 36.965 53.500 37.325 54.120 ;
        RECT 37.045 52.620 37.305 53.500 ;
        RECT 37.585 53.250 40.415 54.300 ;
        RECT 36.875 52.240 37.405 52.620 ;
        RECT 32.265 51.980 32.765 52.070 ;
        RECT 32.255 51.250 32.765 51.980 ;
        RECT 32.495 50.250 32.765 51.250 ;
        RECT 33.405 51.000 33.675 51.950 ;
        RECT 33.405 50.850 33.875 51.000 ;
        RECT 33.405 50.170 33.965 50.850 ;
        RECT 33.485 50.160 33.965 50.170 ;
        RECT 32.775 49.630 33.395 49.990 ;
        RECT 32.815 49.100 33.245 49.630 ;
        RECT 31.365 48.680 33.245 49.100 ;
        RECT 33.735 48.970 33.965 50.160 ;
        RECT 32.815 47.810 33.245 48.680 ;
        RECT 33.655 48.370 34.035 48.970 ;
        RECT 30.525 47.070 31.215 47.780 ;
        RECT 32.635 47.450 33.255 47.810 ;
        RECT 32.335 47.070 32.625 47.260 ;
        RECT 30.525 46.630 32.625 47.070 ;
        RECT 30.525 46.610 31.215 46.630 ;
        RECT 32.335 46.390 32.625 46.630 ;
        RECT 33.255 47.000 33.525 47.250 ;
        RECT 33.735 47.000 33.965 48.370 ;
        RECT 36.555 47.020 36.885 52.040 ;
        RECT 37.605 52.030 38.735 53.250 ;
        RECT 40.095 53.230 40.415 53.250 ;
        RECT 33.255 46.890 33.965 47.000 ;
        RECT 36.545 46.970 36.885 47.020 ;
        RECT 37.435 47.790 38.815 52.030 ;
        RECT 33.255 46.580 33.915 46.890 ;
        RECT 33.255 46.410 33.525 46.580 ;
        RECT 36.545 45.010 36.825 46.970 ;
        RECT 37.435 46.930 37.735 47.790 ;
        RECT 38.515 46.930 38.815 47.790 ;
        RECT 39.365 46.930 39.695 52.000 ;
        RECT 38.765 46.390 39.245 46.770 ;
        RECT 38.865 45.770 39.115 46.390 ;
        RECT 38.765 45.170 39.145 45.770 ;
        RECT 28.215 43.200 28.515 44.930 ;
        RECT 36.025 44.240 37.125 45.010 ;
        RECT 39.415 44.940 39.695 46.930 ;
        RECT 41.745 47.750 42.245 68.550 ;
        RECT 42.585 49.070 42.975 70.580 ;
        RECT 43.375 69.990 44.265 70.720 ;
        RECT 43.475 65.170 43.735 69.990 ;
        RECT 45.115 68.600 47.825 69.450 ;
        RECT 45.315 65.820 47.245 68.600 ;
        RECT 52.975 68.530 53.515 71.760 ;
        RECT 53.815 70.560 54.225 73.290 ;
        RECT 61.475 73.120 63.545 74.400 ;
        RECT 64.400 73.280 66.960 75.810 ;
        RECT 76.140 75.740 76.420 76.950 ;
        RECT 109.970 76.610 110.250 85.420 ;
        RECT 87.580 76.330 110.250 76.610 ;
        RECT 87.580 75.760 87.860 76.330 ;
        RECT 115.950 76.030 116.230 85.700 ;
        RECT 98.850 75.840 116.230 76.030 ;
        RECT 63.895 71.750 64.755 72.590 ;
        RECT 50.215 67.110 51.335 67.790 ;
        RECT 50.495 65.830 51.165 67.110 ;
        RECT 43.875 65.440 48.925 65.820 ;
        RECT 50.285 65.420 51.335 65.830 ;
        RECT 43.475 63.620 43.855 65.170 ;
        RECT 43.595 55.780 43.855 63.620 ;
        RECT 48.905 63.180 49.175 65.220 ;
        RECT 50.035 63.180 50.305 65.180 ;
        RECT 48.905 56.490 50.305 63.180 ;
        RECT 43.505 55.270 43.865 55.780 ;
        RECT 43.485 54.840 43.865 55.270 ;
        RECT 48.905 55.170 49.175 56.490 ;
        RECT 50.035 55.130 50.305 56.490 ;
        RECT 51.305 55.240 51.625 65.170 ;
        RECT 51.305 55.180 51.635 55.240 ;
        RECT 43.485 54.560 43.735 54.840 ;
        RECT 43.285 54.160 47.925 54.560 ;
        RECT 48.825 54.270 49.955 54.280 ;
        RECT 51.315 54.270 51.635 55.180 ;
        RECT 43.485 52.040 43.735 54.160 ;
        RECT 48.185 53.470 48.545 54.090 ;
        RECT 48.265 52.590 48.525 53.470 ;
        RECT 48.805 53.220 51.635 54.270 ;
        RECT 48.095 52.210 48.625 52.590 ;
        RECT 43.485 51.950 43.985 52.040 ;
        RECT 43.475 51.220 43.985 51.950 ;
        RECT 43.715 50.220 43.985 51.220 ;
        RECT 44.625 50.970 44.895 51.920 ;
        RECT 44.625 50.820 45.095 50.970 ;
        RECT 44.625 50.140 45.185 50.820 ;
        RECT 44.705 50.130 45.185 50.140 ;
        RECT 43.995 49.600 44.615 49.960 ;
        RECT 44.035 49.070 44.465 49.600 ;
        RECT 42.585 48.650 44.465 49.070 ;
        RECT 44.955 48.940 45.185 50.130 ;
        RECT 44.035 47.780 44.465 48.650 ;
        RECT 44.875 48.340 45.255 48.940 ;
        RECT 41.745 47.040 42.435 47.750 ;
        RECT 43.855 47.420 44.475 47.780 ;
        RECT 43.555 47.040 43.845 47.230 ;
        RECT 41.745 46.600 43.845 47.040 ;
        RECT 41.745 46.580 42.435 46.600 ;
        RECT 43.555 46.360 43.845 46.600 ;
        RECT 44.475 46.970 44.745 47.220 ;
        RECT 44.955 46.970 45.185 48.340 ;
        RECT 47.775 46.990 48.105 52.010 ;
        RECT 48.825 52.000 49.955 53.220 ;
        RECT 51.315 53.200 51.635 53.220 ;
        RECT 44.475 46.860 45.185 46.970 ;
        RECT 47.765 46.940 48.105 46.990 ;
        RECT 48.655 47.760 50.035 52.000 ;
        RECT 44.475 46.550 45.135 46.860 ;
        RECT 44.475 46.380 44.745 46.550 ;
        RECT 47.765 44.980 48.045 46.940 ;
        RECT 48.655 46.900 48.955 47.760 ;
        RECT 49.735 46.900 50.035 47.760 ;
        RECT 50.585 46.900 50.915 51.970 ;
        RECT 49.985 46.360 50.465 46.740 ;
        RECT 50.085 45.740 50.335 46.360 ;
        RECT 49.985 45.140 50.365 45.740 ;
        RECT 39.415 43.210 39.715 44.940 ;
        RECT 47.245 44.210 48.345 44.980 ;
        RECT 50.635 44.910 50.915 46.900 ;
        RECT 52.995 47.730 53.495 68.530 ;
        RECT 53.835 49.050 54.225 70.560 ;
        RECT 54.625 69.970 55.515 70.700 ;
        RECT 54.725 65.150 54.985 69.970 ;
        RECT 56.365 68.580 59.075 69.430 ;
        RECT 56.565 65.800 58.495 68.580 ;
        RECT 64.195 68.520 64.735 71.750 ;
        RECT 65.035 70.550 65.445 73.280 ;
        RECT 72.585 73.130 74.655 74.410 ;
        RECT 75.550 73.210 78.110 75.740 ;
        RECT 75.135 71.740 75.995 72.580 ;
        RECT 61.465 67.090 62.585 67.770 ;
        RECT 61.745 65.810 62.415 67.090 ;
        RECT 55.125 65.420 60.175 65.800 ;
        RECT 61.535 65.400 62.585 65.810 ;
        RECT 54.725 63.600 55.105 65.150 ;
        RECT 54.845 55.760 55.105 63.600 ;
        RECT 60.155 63.160 60.425 65.200 ;
        RECT 61.285 63.160 61.555 65.160 ;
        RECT 60.155 56.470 61.555 63.160 ;
        RECT 54.755 55.250 55.115 55.760 ;
        RECT 54.735 54.820 55.115 55.250 ;
        RECT 60.155 55.150 60.425 56.470 ;
        RECT 61.285 55.110 61.555 56.470 ;
        RECT 62.555 55.220 62.875 65.150 ;
        RECT 62.555 55.160 62.885 55.220 ;
        RECT 54.735 54.540 54.985 54.820 ;
        RECT 54.535 54.140 59.175 54.540 ;
        RECT 60.075 54.250 61.205 54.260 ;
        RECT 62.565 54.250 62.885 55.160 ;
        RECT 54.735 52.020 54.985 54.140 ;
        RECT 59.435 53.450 59.795 54.070 ;
        RECT 59.515 52.570 59.775 53.450 ;
        RECT 60.055 53.200 62.885 54.250 ;
        RECT 59.345 52.190 59.875 52.570 ;
        RECT 54.735 51.930 55.235 52.020 ;
        RECT 54.725 51.200 55.235 51.930 ;
        RECT 54.965 50.200 55.235 51.200 ;
        RECT 55.875 50.950 56.145 51.900 ;
        RECT 55.875 50.800 56.345 50.950 ;
        RECT 55.875 50.120 56.435 50.800 ;
        RECT 55.955 50.110 56.435 50.120 ;
        RECT 55.245 49.580 55.865 49.940 ;
        RECT 55.285 49.050 55.715 49.580 ;
        RECT 53.835 48.630 55.715 49.050 ;
        RECT 56.205 48.920 56.435 50.110 ;
        RECT 55.285 47.760 55.715 48.630 ;
        RECT 56.125 48.320 56.505 48.920 ;
        RECT 52.995 47.020 53.685 47.730 ;
        RECT 55.105 47.400 55.725 47.760 ;
        RECT 54.805 47.020 55.095 47.210 ;
        RECT 52.995 46.580 55.095 47.020 ;
        RECT 52.995 46.560 53.685 46.580 ;
        RECT 54.805 46.340 55.095 46.580 ;
        RECT 55.725 46.950 55.995 47.200 ;
        RECT 56.205 46.950 56.435 48.320 ;
        RECT 59.025 46.970 59.355 51.990 ;
        RECT 60.075 51.980 61.205 53.200 ;
        RECT 62.565 53.180 62.885 53.200 ;
        RECT 55.725 46.840 56.435 46.950 ;
        RECT 59.015 46.920 59.355 46.970 ;
        RECT 59.905 47.740 61.285 51.980 ;
        RECT 55.725 46.530 56.385 46.840 ;
        RECT 55.725 46.360 55.995 46.530 ;
        RECT 59.015 44.960 59.295 46.920 ;
        RECT 59.905 46.880 60.205 47.740 ;
        RECT 60.985 46.880 61.285 47.740 ;
        RECT 61.835 46.880 62.165 51.950 ;
        RECT 61.235 46.340 61.715 46.720 ;
        RECT 61.335 45.720 61.585 46.340 ;
        RECT 61.235 45.120 61.615 45.720 ;
        RECT 19.865 42.210 21.245 42.780 ;
        RECT 27.495 42.630 28.875 43.200 ;
        RECT 31.145 42.210 32.525 42.780 ;
        RECT 38.695 42.640 40.075 43.210 ;
        RECT 50.635 43.180 50.935 44.910 ;
        RECT 58.495 44.190 59.595 44.960 ;
        RECT 61.885 44.890 62.165 46.880 ;
        RECT 64.215 47.720 64.715 68.520 ;
        RECT 65.055 49.040 65.445 70.550 ;
        RECT 65.845 69.960 66.735 70.690 ;
        RECT 65.945 65.140 66.205 69.960 ;
        RECT 67.585 68.570 70.295 69.420 ;
        RECT 67.785 65.790 69.715 68.570 ;
        RECT 75.435 68.510 75.975 71.740 ;
        RECT 76.275 70.540 76.685 73.210 ;
        RECT 83.855 73.120 85.925 74.400 ;
        RECT 86.850 73.230 89.410 75.760 ;
        RECT 98.150 75.750 116.230 75.840 ;
        RECT 86.385 71.750 87.245 72.590 ;
        RECT 72.685 67.080 73.805 67.760 ;
        RECT 72.965 65.800 73.635 67.080 ;
        RECT 66.345 65.410 71.395 65.790 ;
        RECT 72.755 65.390 73.805 65.800 ;
        RECT 65.945 63.590 66.325 65.140 ;
        RECT 66.065 55.750 66.325 63.590 ;
        RECT 71.375 63.150 71.645 65.190 ;
        RECT 72.505 63.150 72.775 65.150 ;
        RECT 71.375 56.460 72.775 63.150 ;
        RECT 65.975 55.240 66.335 55.750 ;
        RECT 65.955 54.810 66.335 55.240 ;
        RECT 71.375 55.140 71.645 56.460 ;
        RECT 72.505 55.100 72.775 56.460 ;
        RECT 73.775 55.210 74.095 65.140 ;
        RECT 73.775 55.150 74.105 55.210 ;
        RECT 65.955 54.530 66.205 54.810 ;
        RECT 65.755 54.130 70.395 54.530 ;
        RECT 71.295 54.240 72.425 54.250 ;
        RECT 73.785 54.240 74.105 55.150 ;
        RECT 65.955 52.010 66.205 54.130 ;
        RECT 70.655 53.440 71.015 54.060 ;
        RECT 70.735 52.560 70.995 53.440 ;
        RECT 71.275 53.190 74.105 54.240 ;
        RECT 70.565 52.180 71.095 52.560 ;
        RECT 65.955 51.920 66.455 52.010 ;
        RECT 65.945 51.190 66.455 51.920 ;
        RECT 66.185 50.190 66.455 51.190 ;
        RECT 67.095 50.940 67.365 51.890 ;
        RECT 67.095 50.790 67.565 50.940 ;
        RECT 67.095 50.110 67.655 50.790 ;
        RECT 67.175 50.100 67.655 50.110 ;
        RECT 66.465 49.570 67.085 49.930 ;
        RECT 66.505 49.040 66.935 49.570 ;
        RECT 65.055 48.620 66.935 49.040 ;
        RECT 67.425 48.910 67.655 50.100 ;
        RECT 66.505 47.750 66.935 48.620 ;
        RECT 67.345 48.310 67.725 48.910 ;
        RECT 64.215 47.010 64.905 47.720 ;
        RECT 66.325 47.390 66.945 47.750 ;
        RECT 66.025 47.010 66.315 47.200 ;
        RECT 64.215 46.570 66.315 47.010 ;
        RECT 64.215 46.550 64.905 46.570 ;
        RECT 66.025 46.330 66.315 46.570 ;
        RECT 66.945 46.940 67.215 47.190 ;
        RECT 67.425 46.940 67.655 48.310 ;
        RECT 70.245 46.960 70.575 51.980 ;
        RECT 71.295 51.970 72.425 53.190 ;
        RECT 73.785 53.170 74.105 53.190 ;
        RECT 66.945 46.830 67.655 46.940 ;
        RECT 70.235 46.910 70.575 46.960 ;
        RECT 71.125 47.730 72.505 51.970 ;
        RECT 66.945 46.520 67.605 46.830 ;
        RECT 66.945 46.350 67.215 46.520 ;
        RECT 70.235 44.950 70.515 46.910 ;
        RECT 71.125 46.870 71.425 47.730 ;
        RECT 72.205 46.870 72.505 47.730 ;
        RECT 73.055 46.870 73.385 51.940 ;
        RECT 72.455 46.330 72.935 46.710 ;
        RECT 72.555 45.710 72.805 46.330 ;
        RECT 72.455 45.110 72.835 45.710 ;
        RECT 20.225 40.480 20.525 42.210 ;
        RECT 20.245 38.490 20.525 40.480 ;
        RECT 22.815 40.410 23.915 41.180 ;
        RECT 31.505 40.480 31.805 42.210 ;
        RECT 42.435 42.190 43.815 42.760 ;
        RECT 49.915 42.610 51.295 43.180 ;
        RECT 61.885 43.160 62.185 44.890 ;
        RECT 69.715 44.180 70.815 44.950 ;
        RECT 73.105 44.880 73.385 46.870 ;
        RECT 75.455 47.710 75.955 68.510 ;
        RECT 76.295 49.030 76.685 70.540 ;
        RECT 77.085 69.950 77.975 70.680 ;
        RECT 77.185 65.130 77.445 69.950 ;
        RECT 78.825 68.560 81.535 69.410 ;
        RECT 79.025 65.780 80.955 68.560 ;
        RECT 86.685 68.520 87.225 71.750 ;
        RECT 87.525 70.550 87.935 73.230 ;
        RECT 95.045 73.060 97.115 74.340 ;
        RECT 98.150 73.310 100.710 75.750 ;
        RECT 109.390 75.480 111.950 75.560 ;
        RECT 121.930 75.480 122.210 85.700 ;
        RECT 127.550 85.510 128.770 89.380 ;
        RECT 127.910 76.040 128.190 85.510 ;
        RECT 133.380 76.580 136.010 77.880 ;
        RECT 137.240 76.560 139.870 77.860 ;
        RECT 109.390 75.200 122.210 75.480 ;
        RECT 97.665 71.740 98.525 72.580 ;
        RECT 83.925 67.070 85.045 67.750 ;
        RECT 84.205 65.790 84.875 67.070 ;
        RECT 77.585 65.400 82.635 65.780 ;
        RECT 83.995 65.380 85.045 65.790 ;
        RECT 77.185 63.580 77.565 65.130 ;
        RECT 77.305 55.740 77.565 63.580 ;
        RECT 82.615 63.140 82.885 65.180 ;
        RECT 83.745 63.140 84.015 65.140 ;
        RECT 82.615 56.450 84.015 63.140 ;
        RECT 77.215 55.230 77.575 55.740 ;
        RECT 77.195 54.800 77.575 55.230 ;
        RECT 82.615 55.130 82.885 56.450 ;
        RECT 83.745 55.090 84.015 56.450 ;
        RECT 85.015 55.200 85.335 65.130 ;
        RECT 85.015 55.140 85.345 55.200 ;
        RECT 77.195 54.520 77.445 54.800 ;
        RECT 76.995 54.120 81.635 54.520 ;
        RECT 82.535 54.230 83.665 54.240 ;
        RECT 85.025 54.230 85.345 55.140 ;
        RECT 77.195 52.000 77.445 54.120 ;
        RECT 81.895 53.430 82.255 54.050 ;
        RECT 81.975 52.550 82.235 53.430 ;
        RECT 82.515 53.180 85.345 54.230 ;
        RECT 81.805 52.170 82.335 52.550 ;
        RECT 77.195 51.910 77.695 52.000 ;
        RECT 77.185 51.180 77.695 51.910 ;
        RECT 77.425 50.180 77.695 51.180 ;
        RECT 78.335 50.930 78.605 51.880 ;
        RECT 78.335 50.780 78.805 50.930 ;
        RECT 78.335 50.100 78.895 50.780 ;
        RECT 78.415 50.090 78.895 50.100 ;
        RECT 77.705 49.560 78.325 49.920 ;
        RECT 77.745 49.030 78.175 49.560 ;
        RECT 76.295 48.610 78.175 49.030 ;
        RECT 78.665 48.900 78.895 50.090 ;
        RECT 77.745 47.740 78.175 48.610 ;
        RECT 78.585 48.300 78.965 48.900 ;
        RECT 75.455 47.000 76.145 47.710 ;
        RECT 77.565 47.380 78.185 47.740 ;
        RECT 77.265 47.000 77.555 47.190 ;
        RECT 75.455 46.560 77.555 47.000 ;
        RECT 75.455 46.540 76.145 46.560 ;
        RECT 77.265 46.320 77.555 46.560 ;
        RECT 78.185 46.930 78.455 47.180 ;
        RECT 78.665 46.930 78.895 48.300 ;
        RECT 81.485 46.950 81.815 51.970 ;
        RECT 82.535 51.960 83.665 53.180 ;
        RECT 85.025 53.160 85.345 53.180 ;
        RECT 78.185 46.820 78.895 46.930 ;
        RECT 81.475 46.900 81.815 46.950 ;
        RECT 82.365 47.720 83.745 51.960 ;
        RECT 78.185 46.510 78.845 46.820 ;
        RECT 78.185 46.340 78.455 46.510 ;
        RECT 81.475 44.940 81.755 46.900 ;
        RECT 82.365 46.860 82.665 47.720 ;
        RECT 83.445 46.860 83.745 47.720 ;
        RECT 84.295 46.860 84.625 51.930 ;
        RECT 83.695 46.320 84.175 46.700 ;
        RECT 83.795 45.700 84.045 46.320 ;
        RECT 83.695 45.100 84.075 45.700 ;
        RECT 53.655 42.190 55.035 42.760 ;
        RECT 61.165 42.590 62.545 43.160 ;
        RECT 73.105 43.150 73.405 44.880 ;
        RECT 80.955 44.170 82.055 44.940 ;
        RECT 84.345 44.870 84.625 46.860 ;
        RECT 86.705 47.720 87.205 68.520 ;
        RECT 87.545 49.040 87.935 70.550 ;
        RECT 88.335 69.960 89.225 70.690 ;
        RECT 88.435 65.140 88.695 69.960 ;
        RECT 90.075 68.570 92.785 69.420 ;
        RECT 90.275 65.790 92.205 68.570 ;
        RECT 97.965 68.510 98.505 71.740 ;
        RECT 98.805 70.540 99.215 73.310 ;
        RECT 106.455 73.110 108.525 74.390 ;
        RECT 109.390 73.030 111.950 75.200 ;
        RECT 125.760 74.810 128.190 76.040 ;
        RECT 121.290 74.790 128.190 74.810 ;
        RECT 120.600 74.530 128.190 74.790 ;
        RECT 117.655 73.110 119.725 74.390 ;
        RECT 120.600 73.180 128.160 74.530 ;
        RECT 129.505 73.190 131.575 74.470 ;
        RECT 120.600 73.110 126.160 73.180 ;
        RECT 108.935 71.740 109.795 72.580 ;
        RECT 95.175 67.080 96.295 67.760 ;
        RECT 95.455 65.800 96.125 67.080 ;
        RECT 88.835 65.410 93.885 65.790 ;
        RECT 95.245 65.390 96.295 65.800 ;
        RECT 88.435 63.590 88.815 65.140 ;
        RECT 88.555 55.750 88.815 63.590 ;
        RECT 93.865 63.150 94.135 65.190 ;
        RECT 94.995 63.150 95.265 65.150 ;
        RECT 93.865 56.460 95.265 63.150 ;
        RECT 88.465 55.240 88.825 55.750 ;
        RECT 88.445 54.810 88.825 55.240 ;
        RECT 93.865 55.140 94.135 56.460 ;
        RECT 94.995 55.100 95.265 56.460 ;
        RECT 96.265 55.210 96.585 65.140 ;
        RECT 96.265 55.150 96.595 55.210 ;
        RECT 88.445 54.530 88.695 54.810 ;
        RECT 88.245 54.130 92.885 54.530 ;
        RECT 93.785 54.240 94.915 54.250 ;
        RECT 96.275 54.240 96.595 55.150 ;
        RECT 88.445 52.010 88.695 54.130 ;
        RECT 93.145 53.440 93.505 54.060 ;
        RECT 93.225 52.560 93.485 53.440 ;
        RECT 93.765 53.190 96.595 54.240 ;
        RECT 93.055 52.180 93.585 52.560 ;
        RECT 88.445 51.920 88.945 52.010 ;
        RECT 88.435 51.190 88.945 51.920 ;
        RECT 88.675 50.190 88.945 51.190 ;
        RECT 89.585 50.940 89.855 51.890 ;
        RECT 89.585 50.790 90.055 50.940 ;
        RECT 89.585 50.110 90.145 50.790 ;
        RECT 89.665 50.100 90.145 50.110 ;
        RECT 88.955 49.570 89.575 49.930 ;
        RECT 88.995 49.040 89.425 49.570 ;
        RECT 87.545 48.620 89.425 49.040 ;
        RECT 89.915 48.910 90.145 50.100 ;
        RECT 88.995 47.750 89.425 48.620 ;
        RECT 89.835 48.310 90.215 48.910 ;
        RECT 86.705 47.010 87.395 47.720 ;
        RECT 88.815 47.390 89.435 47.750 ;
        RECT 88.515 47.010 88.805 47.200 ;
        RECT 86.705 46.570 88.805 47.010 ;
        RECT 86.705 46.550 87.395 46.570 ;
        RECT 88.515 46.330 88.805 46.570 ;
        RECT 89.435 46.940 89.705 47.190 ;
        RECT 89.915 46.940 90.145 48.310 ;
        RECT 92.735 46.960 93.065 51.980 ;
        RECT 93.785 51.970 94.915 53.190 ;
        RECT 96.275 53.170 96.595 53.190 ;
        RECT 89.435 46.830 90.145 46.940 ;
        RECT 92.725 46.910 93.065 46.960 ;
        RECT 93.615 47.730 94.995 51.970 ;
        RECT 89.435 46.520 90.095 46.830 ;
        RECT 89.435 46.350 89.705 46.520 ;
        RECT 92.725 44.950 93.005 46.910 ;
        RECT 93.615 46.870 93.915 47.730 ;
        RECT 94.695 46.870 94.995 47.730 ;
        RECT 95.545 46.870 95.875 51.940 ;
        RECT 94.945 46.330 95.425 46.710 ;
        RECT 95.045 45.710 95.295 46.330 ;
        RECT 94.945 45.110 95.325 45.710 ;
        RECT 64.855 42.190 66.235 42.760 ;
        RECT 72.385 42.580 73.765 43.150 ;
        RECT 84.345 43.140 84.645 44.870 ;
        RECT 92.205 44.180 93.305 44.950 ;
        RECT 95.595 44.880 95.875 46.870 ;
        RECT 97.985 47.710 98.485 68.510 ;
        RECT 98.825 49.030 99.215 70.540 ;
        RECT 99.615 69.950 100.505 70.680 ;
        RECT 99.715 65.130 99.975 69.950 ;
        RECT 101.355 68.560 104.065 69.410 ;
        RECT 101.555 65.780 103.485 68.560 ;
        RECT 109.235 68.510 109.775 71.740 ;
        RECT 110.075 70.540 110.485 73.030 ;
        RECT 120.185 71.740 121.045 72.580 ;
        RECT 106.455 67.070 107.575 67.750 ;
        RECT 106.735 65.790 107.405 67.070 ;
        RECT 100.115 65.400 105.165 65.780 ;
        RECT 106.525 65.380 107.575 65.790 ;
        RECT 99.715 63.580 100.095 65.130 ;
        RECT 99.835 55.740 100.095 63.580 ;
        RECT 105.145 63.140 105.415 65.180 ;
        RECT 106.275 63.140 106.545 65.140 ;
        RECT 105.145 56.450 106.545 63.140 ;
        RECT 99.745 55.230 100.105 55.740 ;
        RECT 99.725 54.800 100.105 55.230 ;
        RECT 105.145 55.130 105.415 56.450 ;
        RECT 106.275 55.090 106.545 56.450 ;
        RECT 107.545 55.200 107.865 65.130 ;
        RECT 107.545 55.140 107.875 55.200 ;
        RECT 99.725 54.520 99.975 54.800 ;
        RECT 99.525 54.120 104.165 54.520 ;
        RECT 105.065 54.230 106.195 54.240 ;
        RECT 107.555 54.230 107.875 55.140 ;
        RECT 99.725 52.000 99.975 54.120 ;
        RECT 104.425 53.430 104.785 54.050 ;
        RECT 104.505 52.550 104.765 53.430 ;
        RECT 105.045 53.180 107.875 54.230 ;
        RECT 104.335 52.170 104.865 52.550 ;
        RECT 99.725 51.910 100.225 52.000 ;
        RECT 99.715 51.180 100.225 51.910 ;
        RECT 99.955 50.180 100.225 51.180 ;
        RECT 100.865 50.930 101.135 51.880 ;
        RECT 100.865 50.780 101.335 50.930 ;
        RECT 100.865 50.100 101.425 50.780 ;
        RECT 100.945 50.090 101.425 50.100 ;
        RECT 100.235 49.560 100.855 49.920 ;
        RECT 100.275 49.030 100.705 49.560 ;
        RECT 98.825 48.610 100.705 49.030 ;
        RECT 101.195 48.900 101.425 50.090 ;
        RECT 100.275 47.740 100.705 48.610 ;
        RECT 101.115 48.300 101.495 48.900 ;
        RECT 97.985 47.000 98.675 47.710 ;
        RECT 100.095 47.380 100.715 47.740 ;
        RECT 99.795 47.000 100.085 47.190 ;
        RECT 97.985 46.560 100.085 47.000 ;
        RECT 97.985 46.540 98.675 46.560 ;
        RECT 99.795 46.320 100.085 46.560 ;
        RECT 100.715 46.930 100.985 47.180 ;
        RECT 101.195 46.930 101.425 48.300 ;
        RECT 104.015 46.950 104.345 51.970 ;
        RECT 105.065 51.960 106.195 53.180 ;
        RECT 107.555 53.160 107.875 53.180 ;
        RECT 100.715 46.820 101.425 46.930 ;
        RECT 104.005 46.900 104.345 46.950 ;
        RECT 104.895 47.720 106.275 51.960 ;
        RECT 100.715 46.510 101.375 46.820 ;
        RECT 100.715 46.340 100.985 46.510 ;
        RECT 104.005 44.940 104.285 46.900 ;
        RECT 104.895 46.860 105.195 47.720 ;
        RECT 105.975 46.860 106.275 47.720 ;
        RECT 106.825 46.860 107.155 51.930 ;
        RECT 106.225 46.320 106.705 46.700 ;
        RECT 106.325 45.700 106.575 46.320 ;
        RECT 106.225 45.100 106.605 45.700 ;
        RECT 95.595 43.150 95.895 44.880 ;
        RECT 103.485 44.170 104.585 44.940 ;
        RECT 106.875 44.870 107.155 46.860 ;
        RECT 109.255 47.710 109.755 68.510 ;
        RECT 110.095 49.030 110.485 70.540 ;
        RECT 110.885 69.950 111.775 70.680 ;
        RECT 110.985 65.130 111.245 69.950 ;
        RECT 112.625 68.560 115.335 69.410 ;
        RECT 112.825 65.780 114.755 68.560 ;
        RECT 120.485 68.510 121.025 71.740 ;
        RECT 121.325 70.540 121.735 73.110 ;
        RECT 132.925 70.810 133.225 70.900 ;
        RECT 117.725 67.070 118.845 67.750 ;
        RECT 118.005 65.790 118.675 67.070 ;
        RECT 111.385 65.400 116.435 65.780 ;
        RECT 117.795 65.380 118.845 65.790 ;
        RECT 110.985 63.580 111.365 65.130 ;
        RECT 111.105 55.740 111.365 63.580 ;
        RECT 116.415 63.140 116.685 65.180 ;
        RECT 117.545 63.140 117.815 65.140 ;
        RECT 116.415 56.450 117.815 63.140 ;
        RECT 111.015 55.230 111.375 55.740 ;
        RECT 110.995 54.800 111.375 55.230 ;
        RECT 116.415 55.130 116.685 56.450 ;
        RECT 117.545 55.090 117.815 56.450 ;
        RECT 118.815 55.200 119.135 65.130 ;
        RECT 118.815 55.140 119.145 55.200 ;
        RECT 110.995 54.520 111.245 54.800 ;
        RECT 110.795 54.120 115.435 54.520 ;
        RECT 116.335 54.230 117.465 54.240 ;
        RECT 118.825 54.230 119.145 55.140 ;
        RECT 110.995 52.000 111.245 54.120 ;
        RECT 115.695 53.430 116.055 54.050 ;
        RECT 115.775 52.550 116.035 53.430 ;
        RECT 116.315 53.180 119.145 54.230 ;
        RECT 115.605 52.170 116.135 52.550 ;
        RECT 110.995 51.910 111.495 52.000 ;
        RECT 110.985 51.180 111.495 51.910 ;
        RECT 111.225 50.180 111.495 51.180 ;
        RECT 112.135 50.930 112.405 51.880 ;
        RECT 112.135 50.780 112.605 50.930 ;
        RECT 112.135 50.100 112.695 50.780 ;
        RECT 112.215 50.090 112.695 50.100 ;
        RECT 111.505 49.560 112.125 49.920 ;
        RECT 111.545 49.030 111.975 49.560 ;
        RECT 110.095 48.610 111.975 49.030 ;
        RECT 112.465 48.900 112.695 50.090 ;
        RECT 111.545 47.740 111.975 48.610 ;
        RECT 112.385 48.300 112.765 48.900 ;
        RECT 109.255 47.000 109.945 47.710 ;
        RECT 111.365 47.380 111.985 47.740 ;
        RECT 111.065 47.000 111.355 47.190 ;
        RECT 109.255 46.560 111.355 47.000 ;
        RECT 109.255 46.540 109.945 46.560 ;
        RECT 111.065 46.320 111.355 46.560 ;
        RECT 111.985 46.930 112.255 47.180 ;
        RECT 112.465 46.930 112.695 48.300 ;
        RECT 115.285 46.950 115.615 51.970 ;
        RECT 116.335 51.960 117.465 53.180 ;
        RECT 118.825 53.160 119.145 53.180 ;
        RECT 111.985 46.820 112.695 46.930 ;
        RECT 115.275 46.900 115.615 46.950 ;
        RECT 116.165 47.720 117.545 51.960 ;
        RECT 111.985 46.510 112.645 46.820 ;
        RECT 111.985 46.340 112.255 46.510 ;
        RECT 115.275 44.940 115.555 46.900 ;
        RECT 116.165 46.860 116.465 47.720 ;
        RECT 117.245 46.860 117.545 47.720 ;
        RECT 118.095 46.860 118.425 51.930 ;
        RECT 117.495 46.320 117.975 46.700 ;
        RECT 117.595 45.700 117.845 46.320 ;
        RECT 117.495 45.100 117.875 45.700 ;
        RECT 20.795 39.650 21.175 40.250 ;
        RECT 20.825 39.030 21.075 39.650 ;
        RECT 20.695 38.650 21.175 39.030 ;
        RECT 20.245 33.420 20.575 38.490 ;
        RECT 21.125 37.630 21.425 38.490 ;
        RECT 22.205 37.630 22.505 38.490 ;
        RECT 23.115 38.450 23.395 40.410 ;
        RECT 26.415 38.840 26.685 39.010 ;
        RECT 26.025 38.530 26.685 38.840 ;
        RECT 21.125 33.390 22.505 37.630 ;
        RECT 23.055 38.400 23.395 38.450 ;
        RECT 25.975 38.420 26.685 38.530 ;
        RECT 19.525 32.170 19.845 32.190 ;
        RECT 21.205 32.170 22.335 33.390 ;
        RECT 23.055 33.380 23.385 38.400 ;
        RECT 25.975 37.050 26.205 38.420 ;
        RECT 26.415 38.170 26.685 38.420 ;
        RECT 27.315 38.790 27.605 39.030 ;
        RECT 28.725 38.790 29.415 38.810 ;
        RECT 27.315 38.350 29.415 38.790 ;
        RECT 27.315 38.160 27.605 38.350 ;
        RECT 26.685 37.610 27.305 37.970 ;
        RECT 28.725 37.640 29.415 38.350 ;
        RECT 25.905 36.450 26.285 37.050 ;
        RECT 26.695 36.740 27.125 37.610 ;
        RECT 25.975 35.260 26.205 36.450 ;
        RECT 26.695 36.320 28.575 36.740 ;
        RECT 26.695 35.790 27.125 36.320 ;
        RECT 26.545 35.430 27.165 35.790 ;
        RECT 25.975 35.250 26.455 35.260 ;
        RECT 25.975 34.570 26.535 35.250 ;
        RECT 26.065 34.420 26.535 34.570 ;
        RECT 26.265 33.470 26.535 34.420 ;
        RECT 27.175 34.170 27.445 35.170 ;
        RECT 27.175 33.440 27.685 34.170 ;
        RECT 27.175 33.350 27.675 33.440 ;
        RECT 22.535 32.800 23.065 33.180 ;
        RECT 19.525 31.120 22.355 32.170 ;
        RECT 22.635 31.920 22.895 32.800 ;
        RECT 22.615 31.300 22.975 31.920 ;
        RECT 27.425 31.230 27.675 33.350 ;
        RECT 19.525 30.210 19.845 31.120 ;
        RECT 21.205 31.110 22.335 31.120 ;
        RECT 23.235 30.830 27.875 31.230 ;
        RECT 27.425 30.550 27.675 30.830 ;
        RECT 19.525 30.150 19.855 30.210 ;
        RECT 19.535 20.220 19.855 30.150 ;
        RECT 20.855 28.900 21.125 30.260 ;
        RECT 21.985 28.900 22.255 30.220 ;
        RECT 27.295 30.120 27.675 30.550 ;
        RECT 27.295 29.610 27.655 30.120 ;
        RECT 20.855 22.210 22.255 28.900 ;
        RECT 20.855 20.210 21.125 22.210 ;
        RECT 21.985 20.170 22.255 22.210 ;
        RECT 27.305 21.770 27.565 29.610 ;
        RECT 27.305 20.220 27.685 21.770 ;
        RECT 19.825 19.560 20.875 19.970 ;
        RECT 22.235 19.570 27.285 19.950 ;
        RECT 19.995 18.280 20.665 19.560 ;
        RECT 19.825 17.600 20.945 18.280 ;
        RECT 23.915 16.790 25.845 19.570 ;
        RECT 23.335 15.940 26.045 16.790 ;
        RECT 27.425 15.400 27.685 20.220 ;
        RECT 26.895 14.670 27.785 15.400 ;
        RECT 28.185 14.810 28.575 36.320 ;
        RECT 28.915 16.840 29.415 37.640 ;
        RECT 31.525 38.490 31.805 40.480 ;
        RECT 34.095 40.410 35.195 41.180 ;
        RECT 42.795 40.460 43.095 42.190 ;
        RECT 32.075 39.650 32.455 40.250 ;
        RECT 32.105 39.030 32.355 39.650 ;
        RECT 31.975 38.650 32.455 39.030 ;
        RECT 31.525 33.420 31.855 38.490 ;
        RECT 32.405 37.630 32.705 38.490 ;
        RECT 33.485 37.630 33.785 38.490 ;
        RECT 34.395 38.450 34.675 40.410 ;
        RECT 37.695 38.840 37.965 39.010 ;
        RECT 37.305 38.530 37.965 38.840 ;
        RECT 32.405 33.390 33.785 37.630 ;
        RECT 34.335 38.400 34.675 38.450 ;
        RECT 37.255 38.420 37.965 38.530 ;
        RECT 30.805 32.170 31.125 32.190 ;
        RECT 32.485 32.170 33.615 33.390 ;
        RECT 34.335 33.380 34.665 38.400 ;
        RECT 37.255 37.050 37.485 38.420 ;
        RECT 37.695 38.170 37.965 38.420 ;
        RECT 38.595 38.790 38.885 39.030 ;
        RECT 40.005 38.790 40.695 38.810 ;
        RECT 38.595 38.350 40.695 38.790 ;
        RECT 38.595 38.160 38.885 38.350 ;
        RECT 37.965 37.610 38.585 37.970 ;
        RECT 40.005 37.640 40.695 38.350 ;
        RECT 37.185 36.450 37.565 37.050 ;
        RECT 37.975 36.740 38.405 37.610 ;
        RECT 37.255 35.260 37.485 36.450 ;
        RECT 37.975 36.320 39.855 36.740 ;
        RECT 37.975 35.790 38.405 36.320 ;
        RECT 37.825 35.430 38.445 35.790 ;
        RECT 37.255 35.250 37.735 35.260 ;
        RECT 37.255 34.570 37.815 35.250 ;
        RECT 37.345 34.420 37.815 34.570 ;
        RECT 37.545 33.470 37.815 34.420 ;
        RECT 38.455 34.170 38.725 35.170 ;
        RECT 38.455 33.440 38.965 34.170 ;
        RECT 38.455 33.350 38.955 33.440 ;
        RECT 33.815 32.800 34.345 33.180 ;
        RECT 30.805 31.120 33.635 32.170 ;
        RECT 33.915 31.920 34.175 32.800 ;
        RECT 33.895 31.300 34.255 31.920 ;
        RECT 38.705 31.230 38.955 33.350 ;
        RECT 30.805 30.210 31.125 31.120 ;
        RECT 32.485 31.110 33.615 31.120 ;
        RECT 34.515 30.830 39.155 31.230 ;
        RECT 38.705 30.550 38.955 30.830 ;
        RECT 30.805 30.150 31.135 30.210 ;
        RECT 30.815 20.220 31.135 30.150 ;
        RECT 32.135 28.900 32.405 30.260 ;
        RECT 33.265 28.900 33.535 30.220 ;
        RECT 38.575 30.120 38.955 30.550 ;
        RECT 38.575 29.610 38.935 30.120 ;
        RECT 32.135 22.210 33.535 28.900 ;
        RECT 32.135 20.210 32.405 22.210 ;
        RECT 33.265 20.170 33.535 22.210 ;
        RECT 38.585 21.770 38.845 29.610 ;
        RECT 38.585 20.220 38.965 21.770 ;
        RECT 31.105 19.560 32.155 19.970 ;
        RECT 33.515 19.570 38.565 19.950 ;
        RECT 31.275 18.280 31.945 19.560 ;
        RECT 31.105 17.600 32.225 18.280 ;
        RECT 28.185 12.290 28.595 14.810 ;
        RECT 28.895 13.610 29.435 16.840 ;
        RECT 35.195 16.790 37.125 19.570 ;
        RECT 34.615 15.940 37.325 16.790 ;
        RECT 38.705 15.400 38.965 20.220 ;
        RECT 38.175 14.670 39.065 15.400 ;
        RECT 39.465 14.810 39.855 36.320 ;
        RECT 40.195 16.840 40.695 37.640 ;
        RECT 42.815 38.470 43.095 40.460 ;
        RECT 45.385 40.390 46.485 41.160 ;
        RECT 54.015 40.460 54.315 42.190 ;
        RECT 43.365 39.630 43.745 40.230 ;
        RECT 43.395 39.010 43.645 39.630 ;
        RECT 43.265 38.630 43.745 39.010 ;
        RECT 42.815 33.400 43.145 38.470 ;
        RECT 43.695 37.610 43.995 38.470 ;
        RECT 44.775 37.610 45.075 38.470 ;
        RECT 45.685 38.430 45.965 40.390 ;
        RECT 48.985 38.820 49.255 38.990 ;
        RECT 48.595 38.510 49.255 38.820 ;
        RECT 43.695 33.370 45.075 37.610 ;
        RECT 45.625 38.380 45.965 38.430 ;
        RECT 48.545 38.400 49.255 38.510 ;
        RECT 42.095 32.150 42.415 32.170 ;
        RECT 43.775 32.150 44.905 33.370 ;
        RECT 45.625 33.360 45.955 38.380 ;
        RECT 48.545 37.030 48.775 38.400 ;
        RECT 48.985 38.150 49.255 38.400 ;
        RECT 49.885 38.770 50.175 39.010 ;
        RECT 51.295 38.770 51.985 38.790 ;
        RECT 49.885 38.330 51.985 38.770 ;
        RECT 49.885 38.140 50.175 38.330 ;
        RECT 49.255 37.590 49.875 37.950 ;
        RECT 51.295 37.620 51.985 38.330 ;
        RECT 48.475 36.430 48.855 37.030 ;
        RECT 49.265 36.720 49.695 37.590 ;
        RECT 48.545 35.240 48.775 36.430 ;
        RECT 49.265 36.300 51.145 36.720 ;
        RECT 49.265 35.770 49.695 36.300 ;
        RECT 49.115 35.410 49.735 35.770 ;
        RECT 48.545 35.230 49.025 35.240 ;
        RECT 48.545 34.550 49.105 35.230 ;
        RECT 48.635 34.400 49.105 34.550 ;
        RECT 48.835 33.450 49.105 34.400 ;
        RECT 49.745 34.150 50.015 35.150 ;
        RECT 49.745 33.420 50.255 34.150 ;
        RECT 49.745 33.330 50.245 33.420 ;
        RECT 45.105 32.780 45.635 33.160 ;
        RECT 42.095 31.100 44.925 32.150 ;
        RECT 45.205 31.900 45.465 32.780 ;
        RECT 45.185 31.280 45.545 31.900 ;
        RECT 49.995 31.210 50.245 33.330 ;
        RECT 42.095 30.190 42.415 31.100 ;
        RECT 43.775 31.090 44.905 31.100 ;
        RECT 45.805 30.810 50.445 31.210 ;
        RECT 49.995 30.530 50.245 30.810 ;
        RECT 42.095 30.130 42.425 30.190 ;
        RECT 42.105 20.200 42.425 30.130 ;
        RECT 43.425 28.880 43.695 30.240 ;
        RECT 44.555 28.880 44.825 30.200 ;
        RECT 49.865 30.100 50.245 30.530 ;
        RECT 49.865 29.590 50.225 30.100 ;
        RECT 43.425 22.190 44.825 28.880 ;
        RECT 43.425 20.190 43.695 22.190 ;
        RECT 44.555 20.150 44.825 22.190 ;
        RECT 49.875 21.750 50.135 29.590 ;
        RECT 49.875 20.200 50.255 21.750 ;
        RECT 42.395 19.540 43.445 19.950 ;
        RECT 44.805 19.550 49.855 19.930 ;
        RECT 42.565 18.260 43.235 19.540 ;
        RECT 42.395 17.580 43.515 18.260 ;
        RECT 28.875 12.770 29.735 13.610 ;
        RECT 28.185 11.950 30.415 12.290 ;
        RECT 39.465 11.990 39.875 14.810 ;
        RECT 40.175 13.610 40.715 16.840 ;
        RECT 46.485 16.770 48.415 19.550 ;
        RECT 45.905 15.920 48.615 16.770 ;
        RECT 49.995 15.380 50.255 20.200 ;
        RECT 49.465 14.650 50.355 15.380 ;
        RECT 50.755 14.790 51.145 36.300 ;
        RECT 51.485 16.820 51.985 37.620 ;
        RECT 54.035 38.470 54.315 40.460 ;
        RECT 56.605 40.390 57.705 41.160 ;
        RECT 65.215 40.460 65.515 42.190 ;
        RECT 76.145 42.180 77.525 42.750 ;
        RECT 83.625 42.570 85.005 43.140 ;
        RECT 87.385 42.200 88.765 42.770 ;
        RECT 94.875 42.580 96.255 43.150 ;
        RECT 106.875 43.140 107.175 44.870 ;
        RECT 114.755 44.170 115.855 44.940 ;
        RECT 118.145 44.870 118.425 46.860 ;
        RECT 120.505 47.710 121.005 68.510 ;
        RECT 121.345 49.030 121.735 70.540 ;
        RECT 122.135 69.950 123.025 70.680 ;
        RECT 132.615 70.040 134.265 70.810 ;
        RECT 122.235 65.130 122.495 69.950 ;
        RECT 123.875 68.560 126.585 69.410 ;
        RECT 124.075 65.780 126.005 68.560 ;
        RECT 128.975 67.070 130.095 67.750 ;
        RECT 129.255 65.790 129.925 67.070 ;
        RECT 122.635 65.400 127.685 65.780 ;
        RECT 129.045 65.380 130.095 65.790 ;
        RECT 132.925 65.180 133.225 70.040 ;
        RECT 137.675 68.690 139.075 69.460 ;
        RECT 138.385 65.740 138.645 68.690 ;
        RECT 149.410 68.420 150.690 69.620 ;
        RECT 149.480 65.810 150.640 68.420 ;
        RECT 133.365 65.380 138.645 65.740 ;
        RECT 122.235 63.580 122.615 65.130 ;
        RECT 122.355 55.740 122.615 63.580 ;
        RECT 127.665 63.140 127.935 65.180 ;
        RECT 128.795 63.140 129.065 65.140 ;
        RECT 127.665 56.450 129.065 63.140 ;
        RECT 122.265 55.230 122.625 55.740 ;
        RECT 122.245 54.800 122.625 55.230 ;
        RECT 127.665 55.130 127.935 56.450 ;
        RECT 128.795 55.090 129.065 56.450 ;
        RECT 130.065 55.200 130.385 65.130 ;
        RECT 132.925 61.010 133.355 65.180 ;
        RECT 138.385 65.150 138.645 65.380 ;
        RECT 138.385 64.770 138.675 65.150 ;
        RECT 130.065 55.140 130.395 55.200 ;
        RECT 133.055 55.190 133.355 61.010 ;
        RECT 122.245 54.520 122.495 54.800 ;
        RECT 122.045 54.120 126.685 54.520 ;
        RECT 127.585 54.230 128.715 54.240 ;
        RECT 130.075 54.230 130.395 55.140 ;
        RECT 138.395 55.080 138.675 64.770 ;
        RECT 149.390 64.610 150.670 65.810 ;
        RECT 122.245 52.000 122.495 54.120 ;
        RECT 126.945 53.430 127.305 54.050 ;
        RECT 127.025 52.550 127.285 53.430 ;
        RECT 127.565 53.180 130.395 54.230 ;
        RECT 126.855 52.170 127.385 52.550 ;
        RECT 122.245 51.910 122.745 52.000 ;
        RECT 122.235 51.180 122.745 51.910 ;
        RECT 122.475 50.180 122.745 51.180 ;
        RECT 123.385 50.930 123.655 51.880 ;
        RECT 123.385 50.780 123.855 50.930 ;
        RECT 123.385 50.100 123.945 50.780 ;
        RECT 123.465 50.090 123.945 50.100 ;
        RECT 122.755 49.560 123.375 49.920 ;
        RECT 122.795 49.030 123.225 49.560 ;
        RECT 121.345 48.610 123.225 49.030 ;
        RECT 123.715 48.900 123.945 50.090 ;
        RECT 122.795 47.740 123.225 48.610 ;
        RECT 123.635 48.300 124.015 48.900 ;
        RECT 120.505 47.000 121.195 47.710 ;
        RECT 122.615 47.380 123.235 47.740 ;
        RECT 122.315 47.000 122.605 47.190 ;
        RECT 120.505 46.560 122.605 47.000 ;
        RECT 120.505 46.540 121.195 46.560 ;
        RECT 122.315 46.320 122.605 46.560 ;
        RECT 123.235 46.930 123.505 47.180 ;
        RECT 123.715 46.930 123.945 48.300 ;
        RECT 126.535 46.950 126.865 51.970 ;
        RECT 127.585 51.960 128.715 53.180 ;
        RECT 130.075 53.160 130.395 53.180 ;
        RECT 123.235 46.820 123.945 46.930 ;
        RECT 126.525 46.900 126.865 46.950 ;
        RECT 127.415 47.720 128.795 51.960 ;
        RECT 123.235 46.510 123.895 46.820 ;
        RECT 123.235 46.340 123.505 46.510 ;
        RECT 126.525 44.940 126.805 46.900 ;
        RECT 127.415 46.860 127.715 47.720 ;
        RECT 128.495 46.860 128.795 47.720 ;
        RECT 129.345 46.860 129.675 51.930 ;
        RECT 128.745 46.320 129.225 46.700 ;
        RECT 128.845 45.700 129.095 46.320 ;
        RECT 128.745 45.100 129.125 45.700 ;
        RECT 118.145 43.140 118.445 44.870 ;
        RECT 126.005 44.170 127.105 44.940 ;
        RECT 129.395 44.870 129.675 46.860 ;
        RECT 129.395 43.140 129.695 44.870 ;
        RECT 98.595 42.220 99.975 42.790 ;
        RECT 106.155 42.570 107.535 43.140 ;
        RECT 109.795 42.260 111.175 42.830 ;
        RECT 117.425 42.570 118.805 43.140 ;
        RECT 121.005 42.280 122.385 42.850 ;
        RECT 128.675 42.570 130.055 43.140 ;
        RECT 54.585 39.630 54.965 40.230 ;
        RECT 54.615 39.010 54.865 39.630 ;
        RECT 54.485 38.630 54.965 39.010 ;
        RECT 54.035 33.400 54.365 38.470 ;
        RECT 54.915 37.610 55.215 38.470 ;
        RECT 55.995 37.610 56.295 38.470 ;
        RECT 56.905 38.430 57.185 40.390 ;
        RECT 60.205 38.820 60.475 38.990 ;
        RECT 59.815 38.510 60.475 38.820 ;
        RECT 54.915 33.370 56.295 37.610 ;
        RECT 56.845 38.380 57.185 38.430 ;
        RECT 59.765 38.400 60.475 38.510 ;
        RECT 53.315 32.150 53.635 32.170 ;
        RECT 54.995 32.150 56.125 33.370 ;
        RECT 56.845 33.360 57.175 38.380 ;
        RECT 59.765 37.030 59.995 38.400 ;
        RECT 60.205 38.150 60.475 38.400 ;
        RECT 61.105 38.770 61.395 39.010 ;
        RECT 62.515 38.770 63.205 38.790 ;
        RECT 61.105 38.330 63.205 38.770 ;
        RECT 61.105 38.140 61.395 38.330 ;
        RECT 60.475 37.590 61.095 37.950 ;
        RECT 62.515 37.620 63.205 38.330 ;
        RECT 59.695 36.430 60.075 37.030 ;
        RECT 60.485 36.720 60.915 37.590 ;
        RECT 59.765 35.240 59.995 36.430 ;
        RECT 60.485 36.300 62.365 36.720 ;
        RECT 60.485 35.770 60.915 36.300 ;
        RECT 60.335 35.410 60.955 35.770 ;
        RECT 59.765 35.230 60.245 35.240 ;
        RECT 59.765 34.550 60.325 35.230 ;
        RECT 59.855 34.400 60.325 34.550 ;
        RECT 60.055 33.450 60.325 34.400 ;
        RECT 60.965 34.150 61.235 35.150 ;
        RECT 60.965 33.420 61.475 34.150 ;
        RECT 60.965 33.330 61.465 33.420 ;
        RECT 56.325 32.780 56.855 33.160 ;
        RECT 53.315 31.100 56.145 32.150 ;
        RECT 56.425 31.900 56.685 32.780 ;
        RECT 56.405 31.280 56.765 31.900 ;
        RECT 61.215 31.210 61.465 33.330 ;
        RECT 53.315 30.190 53.635 31.100 ;
        RECT 54.995 31.090 56.125 31.100 ;
        RECT 57.025 30.810 61.665 31.210 ;
        RECT 61.215 30.530 61.465 30.810 ;
        RECT 53.315 30.130 53.645 30.190 ;
        RECT 53.325 20.200 53.645 30.130 ;
        RECT 54.645 28.880 54.915 30.240 ;
        RECT 55.775 28.880 56.045 30.200 ;
        RECT 61.085 30.100 61.465 30.530 ;
        RECT 61.085 29.590 61.445 30.100 ;
        RECT 54.645 22.190 56.045 28.880 ;
        RECT 54.645 20.190 54.915 22.190 ;
        RECT 55.775 20.150 56.045 22.190 ;
        RECT 61.095 21.750 61.355 29.590 ;
        RECT 61.095 20.200 61.475 21.750 ;
        RECT 53.615 19.540 54.665 19.950 ;
        RECT 56.025 19.550 61.075 19.930 ;
        RECT 53.785 18.260 54.455 19.540 ;
        RECT 53.615 17.580 54.735 18.260 ;
        RECT 40.155 12.770 41.015 13.610 ;
        RECT 50.755 12.170 51.165 14.790 ;
        RECT 51.465 13.590 52.005 16.820 ;
        RECT 57.705 16.770 59.635 19.550 ;
        RECT 57.125 15.920 59.835 16.770 ;
        RECT 61.215 15.380 61.475 20.200 ;
        RECT 60.685 14.650 61.575 15.380 ;
        RECT 61.975 14.790 62.365 36.300 ;
        RECT 62.705 16.820 63.205 37.620 ;
        RECT 65.235 38.470 65.515 40.460 ;
        RECT 67.805 40.390 68.905 41.160 ;
        RECT 76.505 40.450 76.805 42.180 ;
        RECT 65.785 39.630 66.165 40.230 ;
        RECT 65.815 39.010 66.065 39.630 ;
        RECT 65.685 38.630 66.165 39.010 ;
        RECT 65.235 33.400 65.565 38.470 ;
        RECT 66.115 37.610 66.415 38.470 ;
        RECT 67.195 37.610 67.495 38.470 ;
        RECT 68.105 38.430 68.385 40.390 ;
        RECT 71.405 38.820 71.675 38.990 ;
        RECT 71.015 38.510 71.675 38.820 ;
        RECT 66.115 33.370 67.495 37.610 ;
        RECT 68.045 38.380 68.385 38.430 ;
        RECT 70.965 38.400 71.675 38.510 ;
        RECT 64.515 32.150 64.835 32.170 ;
        RECT 66.195 32.150 67.325 33.370 ;
        RECT 68.045 33.360 68.375 38.380 ;
        RECT 70.965 37.030 71.195 38.400 ;
        RECT 71.405 38.150 71.675 38.400 ;
        RECT 72.305 38.770 72.595 39.010 ;
        RECT 73.715 38.770 74.405 38.790 ;
        RECT 72.305 38.330 74.405 38.770 ;
        RECT 72.305 38.140 72.595 38.330 ;
        RECT 71.675 37.590 72.295 37.950 ;
        RECT 73.715 37.620 74.405 38.330 ;
        RECT 70.895 36.430 71.275 37.030 ;
        RECT 71.685 36.720 72.115 37.590 ;
        RECT 70.965 35.240 71.195 36.430 ;
        RECT 71.685 36.300 73.565 36.720 ;
        RECT 71.685 35.770 72.115 36.300 ;
        RECT 71.535 35.410 72.155 35.770 ;
        RECT 70.965 35.230 71.445 35.240 ;
        RECT 70.965 34.550 71.525 35.230 ;
        RECT 71.055 34.400 71.525 34.550 ;
        RECT 71.255 33.450 71.525 34.400 ;
        RECT 72.165 34.150 72.435 35.150 ;
        RECT 72.165 33.420 72.675 34.150 ;
        RECT 72.165 33.330 72.665 33.420 ;
        RECT 67.525 32.780 68.055 33.160 ;
        RECT 64.515 31.100 67.345 32.150 ;
        RECT 67.625 31.900 67.885 32.780 ;
        RECT 67.605 31.280 67.965 31.900 ;
        RECT 72.415 31.210 72.665 33.330 ;
        RECT 64.515 30.190 64.835 31.100 ;
        RECT 66.195 31.090 67.325 31.100 ;
        RECT 68.225 30.810 72.865 31.210 ;
        RECT 72.415 30.530 72.665 30.810 ;
        RECT 64.515 30.130 64.845 30.190 ;
        RECT 64.525 20.200 64.845 30.130 ;
        RECT 65.845 28.880 66.115 30.240 ;
        RECT 66.975 28.880 67.245 30.200 ;
        RECT 72.285 30.100 72.665 30.530 ;
        RECT 72.285 29.590 72.645 30.100 ;
        RECT 65.845 22.190 67.245 28.880 ;
        RECT 65.845 20.190 66.115 22.190 ;
        RECT 66.975 20.150 67.245 22.190 ;
        RECT 72.295 21.750 72.555 29.590 ;
        RECT 72.295 20.200 72.675 21.750 ;
        RECT 64.815 19.540 65.865 19.950 ;
        RECT 67.225 19.550 72.275 19.930 ;
        RECT 64.985 18.260 65.655 19.540 ;
        RECT 64.815 17.580 65.935 18.260 ;
        RECT 51.445 12.750 52.305 13.590 ;
        RECT 27.865 11.130 30.415 11.950 ;
        RECT 28.395 11.090 30.415 11.130 ;
        RECT 39.115 10.980 41.565 11.990 ;
        RECT 50.335 10.970 52.355 12.170 ;
        RECT 61.975 12.160 62.385 14.790 ;
        RECT 62.685 13.590 63.225 16.820 ;
        RECT 68.905 16.770 70.835 19.550 ;
        RECT 68.325 15.920 71.035 16.770 ;
        RECT 72.415 15.380 72.675 20.200 ;
        RECT 71.885 14.650 72.775 15.380 ;
        RECT 73.175 14.790 73.565 36.300 ;
        RECT 73.905 16.820 74.405 37.620 ;
        RECT 76.525 38.460 76.805 40.450 ;
        RECT 79.095 40.380 80.195 41.150 ;
        RECT 87.745 40.470 88.045 42.200 ;
        RECT 77.075 39.620 77.455 40.220 ;
        RECT 77.105 39.000 77.355 39.620 ;
        RECT 76.975 38.620 77.455 39.000 ;
        RECT 76.525 33.390 76.855 38.460 ;
        RECT 77.405 37.600 77.705 38.460 ;
        RECT 78.485 37.600 78.785 38.460 ;
        RECT 79.395 38.420 79.675 40.380 ;
        RECT 82.695 38.810 82.965 38.980 ;
        RECT 82.305 38.500 82.965 38.810 ;
        RECT 77.405 33.360 78.785 37.600 ;
        RECT 79.335 38.370 79.675 38.420 ;
        RECT 82.255 38.390 82.965 38.500 ;
        RECT 75.805 32.140 76.125 32.160 ;
        RECT 77.485 32.140 78.615 33.360 ;
        RECT 79.335 33.350 79.665 38.370 ;
        RECT 82.255 37.020 82.485 38.390 ;
        RECT 82.695 38.140 82.965 38.390 ;
        RECT 83.595 38.760 83.885 39.000 ;
        RECT 85.005 38.760 85.695 38.780 ;
        RECT 83.595 38.320 85.695 38.760 ;
        RECT 83.595 38.130 83.885 38.320 ;
        RECT 82.965 37.580 83.585 37.940 ;
        RECT 85.005 37.610 85.695 38.320 ;
        RECT 82.185 36.420 82.565 37.020 ;
        RECT 82.975 36.710 83.405 37.580 ;
        RECT 82.255 35.230 82.485 36.420 ;
        RECT 82.975 36.290 84.855 36.710 ;
        RECT 82.975 35.760 83.405 36.290 ;
        RECT 82.825 35.400 83.445 35.760 ;
        RECT 82.255 35.220 82.735 35.230 ;
        RECT 82.255 34.540 82.815 35.220 ;
        RECT 82.345 34.390 82.815 34.540 ;
        RECT 82.545 33.440 82.815 34.390 ;
        RECT 83.455 34.140 83.725 35.140 ;
        RECT 83.455 33.410 83.965 34.140 ;
        RECT 83.455 33.320 83.955 33.410 ;
        RECT 78.815 32.770 79.345 33.150 ;
        RECT 75.805 31.090 78.635 32.140 ;
        RECT 78.915 31.890 79.175 32.770 ;
        RECT 78.895 31.270 79.255 31.890 ;
        RECT 83.705 31.200 83.955 33.320 ;
        RECT 75.805 30.180 76.125 31.090 ;
        RECT 77.485 31.080 78.615 31.090 ;
        RECT 79.515 30.800 84.155 31.200 ;
        RECT 83.705 30.520 83.955 30.800 ;
        RECT 75.805 30.120 76.135 30.180 ;
        RECT 75.815 20.190 76.135 30.120 ;
        RECT 77.135 28.870 77.405 30.230 ;
        RECT 78.265 28.870 78.535 30.190 ;
        RECT 83.575 30.090 83.955 30.520 ;
        RECT 83.575 29.580 83.935 30.090 ;
        RECT 77.135 22.180 78.535 28.870 ;
        RECT 77.135 20.180 77.405 22.180 ;
        RECT 78.265 20.140 78.535 22.180 ;
        RECT 83.585 21.740 83.845 29.580 ;
        RECT 83.585 20.190 83.965 21.740 ;
        RECT 76.105 19.530 77.155 19.940 ;
        RECT 78.515 19.540 83.565 19.920 ;
        RECT 76.275 18.250 76.945 19.530 ;
        RECT 76.105 17.570 77.225 18.250 ;
        RECT 62.665 12.750 63.525 13.590 ;
        RECT 73.175 12.190 73.585 14.790 ;
        RECT 73.885 13.590 74.425 16.820 ;
        RECT 80.195 16.760 82.125 19.540 ;
        RECT 79.615 15.910 82.325 16.760 ;
        RECT 83.705 15.370 83.965 20.190 ;
        RECT 83.175 14.640 84.065 15.370 ;
        RECT 84.465 14.780 84.855 36.290 ;
        RECT 85.195 16.810 85.695 37.610 ;
        RECT 87.765 38.480 88.045 40.470 ;
        RECT 90.335 40.400 91.435 41.170 ;
        RECT 98.955 40.490 99.255 42.220 ;
        RECT 88.315 39.640 88.695 40.240 ;
        RECT 88.345 39.020 88.595 39.640 ;
        RECT 88.215 38.640 88.695 39.020 ;
        RECT 87.765 33.410 88.095 38.480 ;
        RECT 88.645 37.620 88.945 38.480 ;
        RECT 89.725 37.620 90.025 38.480 ;
        RECT 90.635 38.440 90.915 40.400 ;
        RECT 93.935 38.830 94.205 39.000 ;
        RECT 93.545 38.520 94.205 38.830 ;
        RECT 88.645 33.380 90.025 37.620 ;
        RECT 90.575 38.390 90.915 38.440 ;
        RECT 93.495 38.410 94.205 38.520 ;
        RECT 87.045 32.160 87.365 32.180 ;
        RECT 88.725 32.160 89.855 33.380 ;
        RECT 90.575 33.370 90.905 38.390 ;
        RECT 93.495 37.040 93.725 38.410 ;
        RECT 93.935 38.160 94.205 38.410 ;
        RECT 94.835 38.780 95.125 39.020 ;
        RECT 96.245 38.780 96.935 38.800 ;
        RECT 94.835 38.340 96.935 38.780 ;
        RECT 94.835 38.150 95.125 38.340 ;
        RECT 94.205 37.600 94.825 37.960 ;
        RECT 96.245 37.630 96.935 38.340 ;
        RECT 93.425 36.440 93.805 37.040 ;
        RECT 94.215 36.730 94.645 37.600 ;
        RECT 93.495 35.250 93.725 36.440 ;
        RECT 94.215 36.310 96.095 36.730 ;
        RECT 94.215 35.780 94.645 36.310 ;
        RECT 94.065 35.420 94.685 35.780 ;
        RECT 93.495 35.240 93.975 35.250 ;
        RECT 93.495 34.560 94.055 35.240 ;
        RECT 93.585 34.410 94.055 34.560 ;
        RECT 93.785 33.460 94.055 34.410 ;
        RECT 94.695 34.160 94.965 35.160 ;
        RECT 94.695 33.430 95.205 34.160 ;
        RECT 94.695 33.340 95.195 33.430 ;
        RECT 90.055 32.790 90.585 33.170 ;
        RECT 87.045 31.110 89.875 32.160 ;
        RECT 90.155 31.910 90.415 32.790 ;
        RECT 90.135 31.290 90.495 31.910 ;
        RECT 94.945 31.220 95.195 33.340 ;
        RECT 87.045 30.200 87.365 31.110 ;
        RECT 88.725 31.100 89.855 31.110 ;
        RECT 90.755 30.820 95.395 31.220 ;
        RECT 94.945 30.540 95.195 30.820 ;
        RECT 87.045 30.140 87.375 30.200 ;
        RECT 87.055 20.210 87.375 30.140 ;
        RECT 88.375 28.890 88.645 30.250 ;
        RECT 89.505 28.890 89.775 30.210 ;
        RECT 94.815 30.110 95.195 30.540 ;
        RECT 94.815 29.600 95.175 30.110 ;
        RECT 88.375 22.200 89.775 28.890 ;
        RECT 88.375 20.200 88.645 22.200 ;
        RECT 89.505 20.160 89.775 22.200 ;
        RECT 94.825 21.760 95.085 29.600 ;
        RECT 94.825 20.210 95.205 21.760 ;
        RECT 87.345 19.550 88.395 19.960 ;
        RECT 89.755 19.560 94.805 19.940 ;
        RECT 87.515 18.270 88.185 19.550 ;
        RECT 87.345 17.590 88.465 18.270 ;
        RECT 73.865 12.750 74.725 13.590 ;
        RECT 61.415 10.960 63.435 12.160 ;
        RECT 72.725 10.990 74.745 12.190 ;
        RECT 84.465 12.180 84.875 14.780 ;
        RECT 85.175 13.580 85.715 16.810 ;
        RECT 91.435 16.780 93.365 19.560 ;
        RECT 90.855 15.930 93.565 16.780 ;
        RECT 94.945 15.390 95.205 20.210 ;
        RECT 94.415 14.660 95.305 15.390 ;
        RECT 95.705 14.800 96.095 36.310 ;
        RECT 96.435 16.830 96.935 37.630 ;
        RECT 98.975 38.500 99.255 40.490 ;
        RECT 101.545 40.420 102.645 41.190 ;
        RECT 110.155 40.530 110.455 42.260 ;
        RECT 99.525 39.660 99.905 40.260 ;
        RECT 99.555 39.040 99.805 39.660 ;
        RECT 99.425 38.660 99.905 39.040 ;
        RECT 98.975 33.430 99.305 38.500 ;
        RECT 99.855 37.640 100.155 38.500 ;
        RECT 100.935 37.640 101.235 38.500 ;
        RECT 101.845 38.460 102.125 40.420 ;
        RECT 105.145 38.850 105.415 39.020 ;
        RECT 104.755 38.540 105.415 38.850 ;
        RECT 99.855 33.400 101.235 37.640 ;
        RECT 101.785 38.410 102.125 38.460 ;
        RECT 104.705 38.430 105.415 38.540 ;
        RECT 98.255 32.180 98.575 32.200 ;
        RECT 99.935 32.180 101.065 33.400 ;
        RECT 101.785 33.390 102.115 38.410 ;
        RECT 104.705 37.060 104.935 38.430 ;
        RECT 105.145 38.180 105.415 38.430 ;
        RECT 106.045 38.800 106.335 39.040 ;
        RECT 107.455 38.800 108.145 38.820 ;
        RECT 106.045 38.360 108.145 38.800 ;
        RECT 106.045 38.170 106.335 38.360 ;
        RECT 105.415 37.620 106.035 37.980 ;
        RECT 107.455 37.650 108.145 38.360 ;
        RECT 104.635 36.460 105.015 37.060 ;
        RECT 105.425 36.750 105.855 37.620 ;
        RECT 104.705 35.270 104.935 36.460 ;
        RECT 105.425 36.330 107.305 36.750 ;
        RECT 105.425 35.800 105.855 36.330 ;
        RECT 105.275 35.440 105.895 35.800 ;
        RECT 104.705 35.260 105.185 35.270 ;
        RECT 104.705 34.580 105.265 35.260 ;
        RECT 104.795 34.430 105.265 34.580 ;
        RECT 104.995 33.480 105.265 34.430 ;
        RECT 105.905 34.180 106.175 35.180 ;
        RECT 105.905 33.450 106.415 34.180 ;
        RECT 105.905 33.360 106.405 33.450 ;
        RECT 101.265 32.810 101.795 33.190 ;
        RECT 98.255 31.130 101.085 32.180 ;
        RECT 101.365 31.930 101.625 32.810 ;
        RECT 101.345 31.310 101.705 31.930 ;
        RECT 106.155 31.240 106.405 33.360 ;
        RECT 98.255 30.220 98.575 31.130 ;
        RECT 99.935 31.120 101.065 31.130 ;
        RECT 101.965 30.840 106.605 31.240 ;
        RECT 106.155 30.560 106.405 30.840 ;
        RECT 98.255 30.160 98.585 30.220 ;
        RECT 98.265 20.230 98.585 30.160 ;
        RECT 99.585 28.910 99.855 30.270 ;
        RECT 100.715 28.910 100.985 30.230 ;
        RECT 106.025 30.130 106.405 30.560 ;
        RECT 106.025 29.620 106.385 30.130 ;
        RECT 99.585 22.220 100.985 28.910 ;
        RECT 99.585 20.220 99.855 22.220 ;
        RECT 100.715 20.180 100.985 22.220 ;
        RECT 106.035 21.780 106.295 29.620 ;
        RECT 106.035 20.230 106.415 21.780 ;
        RECT 98.555 19.570 99.605 19.980 ;
        RECT 100.965 19.580 106.015 19.960 ;
        RECT 98.725 18.290 99.395 19.570 ;
        RECT 98.555 17.610 99.675 18.290 ;
        RECT 85.155 12.740 86.015 13.580 ;
        RECT 95.705 12.180 96.115 14.800 ;
        RECT 96.415 13.600 96.955 16.830 ;
        RECT 102.645 16.800 104.575 19.580 ;
        RECT 102.065 15.950 104.775 16.800 ;
        RECT 106.155 15.410 106.415 20.230 ;
        RECT 105.625 14.680 106.515 15.410 ;
        RECT 106.915 14.820 107.305 36.330 ;
        RECT 107.645 16.850 108.145 37.650 ;
        RECT 110.175 38.540 110.455 40.530 ;
        RECT 112.745 40.460 113.845 41.230 ;
        RECT 121.365 40.550 121.665 42.280 ;
        RECT 142.880 42.020 144.100 43.390 ;
        RECT 110.725 39.700 111.105 40.300 ;
        RECT 110.755 39.080 111.005 39.700 ;
        RECT 110.625 38.700 111.105 39.080 ;
        RECT 110.175 33.470 110.505 38.540 ;
        RECT 111.055 37.680 111.355 38.540 ;
        RECT 112.135 37.680 112.435 38.540 ;
        RECT 113.045 38.500 113.325 40.460 ;
        RECT 116.345 38.890 116.615 39.060 ;
        RECT 115.955 38.580 116.615 38.890 ;
        RECT 111.055 33.440 112.435 37.680 ;
        RECT 112.985 38.450 113.325 38.500 ;
        RECT 115.905 38.470 116.615 38.580 ;
        RECT 109.455 32.220 109.775 32.240 ;
        RECT 111.135 32.220 112.265 33.440 ;
        RECT 112.985 33.430 113.315 38.450 ;
        RECT 115.905 37.100 116.135 38.470 ;
        RECT 116.345 38.220 116.615 38.470 ;
        RECT 117.245 38.840 117.535 39.080 ;
        RECT 118.655 38.840 119.345 38.860 ;
        RECT 117.245 38.400 119.345 38.840 ;
        RECT 117.245 38.210 117.535 38.400 ;
        RECT 116.615 37.660 117.235 38.020 ;
        RECT 118.655 37.690 119.345 38.400 ;
        RECT 115.835 36.500 116.215 37.100 ;
        RECT 116.625 36.790 117.055 37.660 ;
        RECT 115.905 35.310 116.135 36.500 ;
        RECT 116.625 36.370 118.505 36.790 ;
        RECT 116.625 35.840 117.055 36.370 ;
        RECT 116.475 35.480 117.095 35.840 ;
        RECT 115.905 35.300 116.385 35.310 ;
        RECT 115.905 34.620 116.465 35.300 ;
        RECT 115.995 34.470 116.465 34.620 ;
        RECT 116.195 33.520 116.465 34.470 ;
        RECT 117.105 34.220 117.375 35.220 ;
        RECT 117.105 33.490 117.615 34.220 ;
        RECT 117.105 33.400 117.605 33.490 ;
        RECT 112.465 32.850 112.995 33.230 ;
        RECT 109.455 31.170 112.285 32.220 ;
        RECT 112.565 31.970 112.825 32.850 ;
        RECT 112.545 31.350 112.905 31.970 ;
        RECT 117.355 31.280 117.605 33.400 ;
        RECT 109.455 30.260 109.775 31.170 ;
        RECT 111.135 31.160 112.265 31.170 ;
        RECT 113.165 30.880 117.805 31.280 ;
        RECT 117.355 30.600 117.605 30.880 ;
        RECT 109.455 30.200 109.785 30.260 ;
        RECT 109.465 20.270 109.785 30.200 ;
        RECT 110.785 28.950 111.055 30.310 ;
        RECT 111.915 28.950 112.185 30.270 ;
        RECT 117.225 30.170 117.605 30.600 ;
        RECT 117.225 29.660 117.585 30.170 ;
        RECT 110.785 22.260 112.185 28.950 ;
        RECT 110.785 20.260 111.055 22.260 ;
        RECT 111.915 20.220 112.185 22.260 ;
        RECT 117.235 21.820 117.495 29.660 ;
        RECT 117.235 20.270 117.615 21.820 ;
        RECT 109.755 19.610 110.805 20.020 ;
        RECT 112.165 19.620 117.215 20.000 ;
        RECT 109.925 18.330 110.595 19.610 ;
        RECT 109.755 17.650 110.875 18.330 ;
        RECT 96.395 12.760 97.255 13.600 ;
        RECT 106.915 12.230 107.325 14.820 ;
        RECT 107.625 13.620 108.165 16.850 ;
        RECT 113.845 16.840 115.775 19.620 ;
        RECT 113.265 15.990 115.975 16.840 ;
        RECT 117.355 15.450 117.615 20.270 ;
        RECT 116.825 14.720 117.715 15.450 ;
        RECT 118.115 14.860 118.505 36.370 ;
        RECT 118.845 16.890 119.345 37.690 ;
        RECT 121.385 38.560 121.665 40.550 ;
        RECT 123.955 40.480 125.055 41.250 ;
        RECT 121.935 39.720 122.315 40.320 ;
        RECT 121.965 39.100 122.215 39.720 ;
        RECT 121.835 38.720 122.315 39.100 ;
        RECT 121.385 33.490 121.715 38.560 ;
        RECT 122.265 37.700 122.565 38.560 ;
        RECT 123.345 37.700 123.645 38.560 ;
        RECT 124.255 38.520 124.535 40.480 ;
        RECT 127.555 38.910 127.825 39.080 ;
        RECT 127.165 38.600 127.825 38.910 ;
        RECT 122.265 33.460 123.645 37.700 ;
        RECT 124.195 38.470 124.535 38.520 ;
        RECT 127.115 38.490 127.825 38.600 ;
        RECT 120.665 32.240 120.985 32.260 ;
        RECT 122.345 32.240 123.475 33.460 ;
        RECT 124.195 33.450 124.525 38.470 ;
        RECT 127.115 37.120 127.345 38.490 ;
        RECT 127.555 38.240 127.825 38.490 ;
        RECT 128.455 38.860 128.745 39.100 ;
        RECT 142.940 38.950 144.100 42.020 ;
        RECT 129.865 38.860 130.555 38.880 ;
        RECT 128.455 38.420 130.555 38.860 ;
        RECT 128.455 38.230 128.745 38.420 ;
        RECT 127.825 37.680 128.445 38.040 ;
        RECT 129.865 37.710 130.555 38.420 ;
        RECT 127.045 36.520 127.425 37.120 ;
        RECT 127.835 36.810 128.265 37.680 ;
        RECT 127.115 35.330 127.345 36.520 ;
        RECT 127.835 36.390 129.715 36.810 ;
        RECT 127.835 35.860 128.265 36.390 ;
        RECT 127.685 35.500 128.305 35.860 ;
        RECT 127.115 35.320 127.595 35.330 ;
        RECT 127.115 34.640 127.675 35.320 ;
        RECT 127.205 34.490 127.675 34.640 ;
        RECT 127.405 33.540 127.675 34.490 ;
        RECT 128.315 34.240 128.585 35.240 ;
        RECT 128.315 33.510 128.825 34.240 ;
        RECT 128.315 33.420 128.815 33.510 ;
        RECT 123.675 32.870 124.205 33.250 ;
        RECT 120.665 31.190 123.495 32.240 ;
        RECT 123.775 31.990 124.035 32.870 ;
        RECT 123.755 31.370 124.115 31.990 ;
        RECT 128.565 31.300 128.815 33.420 ;
        RECT 120.665 30.280 120.985 31.190 ;
        RECT 122.345 31.180 123.475 31.190 ;
        RECT 124.375 30.900 129.015 31.300 ;
        RECT 128.565 30.620 128.815 30.900 ;
        RECT 120.665 30.220 120.995 30.280 ;
        RECT 120.675 20.290 120.995 30.220 ;
        RECT 121.995 28.970 122.265 30.330 ;
        RECT 123.125 28.970 123.395 30.290 ;
        RECT 128.435 30.190 128.815 30.620 ;
        RECT 128.435 29.680 128.795 30.190 ;
        RECT 121.995 22.280 123.395 28.970 ;
        RECT 121.995 20.280 122.265 22.280 ;
        RECT 123.125 20.240 123.395 22.280 ;
        RECT 128.445 21.840 128.705 29.680 ;
        RECT 128.445 20.290 128.825 21.840 ;
        RECT 120.965 19.630 122.015 20.040 ;
        RECT 123.375 19.640 128.425 20.020 ;
        RECT 121.135 18.350 121.805 19.630 ;
        RECT 120.965 17.670 122.085 18.350 ;
        RECT 107.605 12.780 108.465 13.620 ;
        RECT 118.115 12.230 118.525 14.860 ;
        RECT 118.825 13.660 119.365 16.890 ;
        RECT 125.055 16.860 126.985 19.640 ;
        RECT 124.475 16.010 127.185 16.860 ;
        RECT 128.565 15.470 128.825 20.290 ;
        RECT 128.035 14.740 128.925 15.470 ;
        RECT 129.325 14.880 129.715 36.390 ;
        RECT 130.055 16.910 130.555 37.710 ;
        RECT 142.900 37.580 144.120 38.950 ;
        RECT 132.395 24.340 132.705 30.230 ;
        RECT 132.195 20.120 132.705 24.340 ;
        RECT 118.805 12.820 119.665 13.660 ;
        RECT 129.325 12.260 129.735 14.880 ;
        RECT 130.035 13.680 130.575 16.910 ;
        RECT 132.195 15.510 132.505 20.120 ;
        RECT 137.715 19.980 138.005 30.170 ;
        RECT 132.685 19.590 138.005 19.980 ;
        RECT 137.715 16.940 138.005 19.590 ;
        RECT 142.940 17.940 144.090 19.160 ;
        RECT 145.080 18.760 146.200 18.930 ;
        RECT 137.395 15.890 138.295 16.940 ;
        RECT 137.715 15.720 138.005 15.890 ;
        RECT 131.975 14.270 132.735 15.510 ;
        RECT 142.940 15.090 144.050 17.940 ;
        RECT 142.900 13.870 144.050 15.090 ;
        RECT 145.070 14.920 146.200 18.760 ;
        RECT 145.030 13.970 146.200 14.920 ;
        RECT 145.030 13.900 146.150 13.970 ;
        RECT 130.015 12.840 130.875 13.680 ;
        RECT 83.845 10.980 85.865 12.180 ;
        RECT 95.145 10.980 97.165 12.180 ;
        RECT 106.335 11.030 108.355 12.230 ;
        RECT 117.565 11.030 119.585 12.230 ;
        RECT 128.865 11.060 130.885 12.260 ;
        RECT 74.340 0.110 75.630 1.460 ;
        RECT 93.550 0.180 94.840 1.530 ;
        RECT 112.950 0.310 114.240 1.660 ;
        RECT 131.850 0.380 133.490 1.930 ;
        RECT 151.650 0.250 152.920 1.470 ;
      LAYER met3 ;
        RECT 135.340 223.855 136.790 225.205 ;
        RECT 138.130 223.785 139.580 225.135 ;
        RECT 143.180 223.815 144.630 225.165 ;
        RECT 17.380 193.455 18.960 193.785 ;
        RECT 40.955 193.455 42.535 193.785 ;
        RECT 64.530 193.455 66.110 193.785 ;
        RECT 88.105 193.455 89.685 193.785 ;
        RECT 29.165 190.735 30.745 191.065 ;
        RECT 52.740 190.735 54.320 191.065 ;
        RECT 76.315 190.735 77.895 191.065 ;
        RECT 99.890 190.735 101.470 191.065 ;
        RECT 17.380 188.015 18.960 188.345 ;
        RECT 40.955 188.015 42.535 188.345 ;
        RECT 64.530 188.015 66.110 188.345 ;
        RECT 88.105 188.015 89.685 188.345 ;
        RECT 29.165 185.295 30.745 185.625 ;
        RECT 52.740 185.295 54.320 185.625 ;
        RECT 76.315 185.295 77.895 185.625 ;
        RECT 99.890 185.295 101.470 185.625 ;
        RECT 17.380 182.575 18.960 182.905 ;
        RECT 40.955 182.575 42.535 182.905 ;
        RECT 64.530 182.575 66.110 182.905 ;
        RECT 88.105 182.575 89.685 182.905 ;
        RECT 29.165 179.855 30.745 180.185 ;
        RECT 52.740 179.855 54.320 180.185 ;
        RECT 76.315 179.855 77.895 180.185 ;
        RECT 99.890 179.855 101.470 180.185 ;
        RECT 65.150 178.470 65.480 178.485 ;
        RECT 66.735 178.470 67.115 178.480 ;
        RECT 65.150 178.170 67.115 178.470 ;
        RECT 65.150 178.155 65.480 178.170 ;
        RECT 66.735 178.160 67.115 178.170 ;
        RECT 17.380 177.135 18.960 177.465 ;
        RECT 40.955 177.135 42.535 177.465 ;
        RECT 64.530 177.135 66.110 177.465 ;
        RECT 88.105 177.135 89.685 177.465 ;
        RECT 29.165 174.415 30.745 174.745 ;
        RECT 52.740 174.415 54.320 174.745 ;
        RECT 76.315 174.415 77.895 174.745 ;
        RECT 99.890 174.415 101.470 174.745 ;
        RECT 133.700 172.500 134.930 172.705 ;
        RECT 17.380 171.695 18.960 172.025 ;
        RECT 40.955 171.695 42.535 172.025 ;
        RECT 64.530 171.695 66.110 172.025 ;
        RECT 88.105 171.695 89.685 172.025 ;
        RECT 129.030 170.130 134.930 172.500 ;
        RECT 133.700 170.095 134.930 170.130 ;
        RECT 29.165 168.975 30.745 169.305 ;
        RECT 52.740 168.975 54.320 169.305 ;
        RECT 76.315 168.975 77.895 169.305 ;
        RECT 99.890 168.975 101.470 169.305 ;
        RECT 31.110 168.270 31.440 168.285 ;
        RECT 42.610 168.270 42.940 168.285 ;
        RECT 47.210 168.270 47.540 168.285 ;
        RECT 31.110 167.970 47.540 168.270 ;
        RECT 31.110 167.955 31.440 167.970 ;
        RECT 42.610 167.955 42.940 167.970 ;
        RECT 47.210 167.955 47.540 167.970 ;
        RECT 40.310 167.590 40.640 167.605 ;
        RECT 46.750 167.590 47.080 167.605 ;
        RECT 40.310 167.290 47.080 167.590 ;
        RECT 40.310 167.275 40.640 167.290 ;
        RECT 46.750 167.275 47.080 167.290 ;
        RECT 17.380 166.255 18.960 166.585 ;
        RECT 40.955 166.255 42.535 166.585 ;
        RECT 64.530 166.255 66.110 166.585 ;
        RECT 88.105 166.255 89.685 166.585 ;
        RECT 29.165 163.535 30.745 163.865 ;
        RECT 52.740 163.535 54.320 163.865 ;
        RECT 76.315 163.535 77.895 163.865 ;
        RECT 99.890 163.535 101.470 163.865 ;
        RECT 43.530 162.150 43.860 162.165 ;
        RECT 44.655 162.150 45.035 162.160 ;
        RECT 43.530 161.850 45.035 162.150 ;
        RECT 43.530 161.835 43.860 161.850 ;
        RECT 44.655 161.840 45.035 161.850 ;
        RECT 55.695 162.150 56.075 162.160 ;
        RECT 72.050 162.150 72.380 162.165 ;
        RECT 55.695 161.850 72.380 162.150 ;
        RECT 55.695 161.840 56.075 161.850 ;
        RECT 72.050 161.835 72.380 161.850 ;
        RECT 17.380 160.815 18.960 161.145 ;
        RECT 40.955 160.815 42.535 161.145 ;
        RECT 64.530 160.815 66.110 161.145 ;
        RECT 88.105 160.815 89.685 161.145 ;
        RECT 61.930 159.430 62.260 159.445 ;
        RECT 65.610 159.430 65.940 159.445 ;
        RECT 61.930 159.130 65.940 159.430 ;
        RECT 61.930 159.115 62.260 159.130 ;
        RECT 65.610 159.115 65.940 159.130 ;
        RECT 68.830 159.430 69.160 159.445 ;
        RECT 85.850 159.430 86.180 159.445 ;
        RECT 68.830 159.130 86.180 159.430 ;
        RECT 68.830 159.115 69.160 159.130 ;
        RECT 85.850 159.115 86.180 159.130 ;
        RECT 111.150 159.430 111.480 159.445 ;
        RECT 113.225 159.430 115.225 159.580 ;
        RECT 111.150 159.130 115.225 159.430 ;
        RECT 111.150 159.115 111.480 159.130 ;
        RECT 113.225 158.980 115.225 159.130 ;
        RECT 44.910 158.750 45.240 158.765 ;
        RECT 46.495 158.750 46.875 158.760 ;
        RECT 44.910 158.450 46.875 158.750 ;
        RECT 44.910 158.435 45.240 158.450 ;
        RECT 46.495 158.440 46.875 158.450 ;
        RECT 29.165 158.095 30.745 158.425 ;
        RECT 52.740 158.095 54.320 158.425 ;
        RECT 76.315 158.095 77.895 158.425 ;
        RECT 99.890 158.095 101.470 158.425 ;
        RECT 40.310 157.400 40.640 157.405 ;
        RECT 40.055 157.390 40.640 157.400 ;
        RECT 39.855 157.090 40.640 157.390 ;
        RECT 40.055 157.080 40.640 157.090 ;
        RECT 40.310 157.075 40.640 157.080 ;
        RECT 38.930 156.710 39.260 156.725 ;
        RECT 52.730 156.710 53.060 156.725 ;
        RECT 55.695 156.710 56.075 156.720 ;
        RECT 38.930 156.410 56.075 156.710 ;
        RECT 38.930 156.395 39.260 156.410 ;
        RECT 52.730 156.395 53.060 156.410 ;
        RECT 55.695 156.400 56.075 156.410 ;
        RECT 61.470 156.710 61.800 156.725 ;
        RECT 66.530 156.710 66.860 156.725 ;
        RECT 61.470 156.410 66.860 156.710 ;
        RECT 61.470 156.395 61.800 156.410 ;
        RECT 66.530 156.395 66.860 156.410 ;
        RECT 43.530 156.040 43.860 156.045 ;
        RECT 43.530 156.030 44.115 156.040 ;
        RECT 43.305 155.730 44.115 156.030 ;
        RECT 43.530 155.720 44.115 155.730 ;
        RECT 43.530 155.715 43.860 155.720 ;
        RECT 17.380 155.375 18.960 155.705 ;
        RECT 40.955 155.375 42.535 155.705 ;
        RECT 64.530 155.375 66.110 155.705 ;
        RECT 88.105 155.375 89.685 155.705 ;
        RECT 66.990 155.350 67.320 155.365 ;
        RECT 72.510 155.350 72.840 155.365 ;
        RECT 66.990 155.050 72.840 155.350 ;
        RECT 66.990 155.035 67.320 155.050 ;
        RECT 72.510 155.035 72.840 155.050 ;
        RECT 42.610 154.670 42.940 154.685 ;
        RECT 61.470 154.670 61.800 154.685 ;
        RECT 42.610 154.370 61.800 154.670 ;
        RECT 42.610 154.355 42.940 154.370 ;
        RECT 61.470 154.355 61.800 154.370 ;
        RECT 63.310 154.670 63.640 154.685 ;
        RECT 69.750 154.670 70.080 154.685 ;
        RECT 63.310 154.370 70.080 154.670 ;
        RECT 63.310 154.355 63.640 154.370 ;
        RECT 69.750 154.355 70.080 154.370 ;
        RECT 72.050 154.670 72.380 154.685 ;
        RECT 81.710 154.670 82.040 154.685 ;
        RECT 72.050 154.370 82.040 154.670 ;
        RECT 72.050 154.355 72.380 154.370 ;
        RECT 81.710 154.355 82.040 154.370 ;
        RECT 52.270 153.990 52.600 154.005 ;
        RECT 75.730 153.990 76.060 154.005 ;
        RECT 97.095 153.990 97.475 154.000 ;
        RECT 102.410 153.990 102.740 154.005 ;
        RECT 52.270 153.690 92.835 153.990 ;
        RECT 52.270 153.675 52.600 153.690 ;
        RECT 75.730 153.675 76.060 153.690 ;
        RECT 66.990 153.310 67.320 153.325 ;
        RECT 68.370 153.310 68.700 153.325 ;
        RECT 66.990 153.010 68.700 153.310 ;
        RECT 92.535 153.310 92.835 153.690 ;
        RECT 94.375 153.690 102.740 153.990 ;
        RECT 94.375 153.310 94.675 153.690 ;
        RECT 97.095 153.680 97.475 153.690 ;
        RECT 102.410 153.675 102.740 153.690 ;
        RECT 92.535 153.010 94.675 153.310 ;
        RECT 66.990 152.995 67.320 153.010 ;
        RECT 68.370 152.995 68.700 153.010 ;
        RECT 29.165 152.655 30.745 152.985 ;
        RECT 52.740 152.655 54.320 152.985 ;
        RECT 76.315 152.655 77.895 152.985 ;
        RECT 99.890 152.655 101.470 152.985 ;
        RECT 60.090 151.950 60.420 151.965 ;
        RECT 63.310 151.950 63.640 151.965 ;
        RECT 68.830 151.950 69.160 151.965 ;
        RECT 73.890 151.950 74.220 151.965 ;
        RECT 60.090 151.650 67.075 151.950 ;
        RECT 60.090 151.635 60.420 151.650 ;
        RECT 63.310 151.635 63.640 151.650 ;
        RECT 66.775 151.270 67.075 151.650 ;
        RECT 68.830 151.650 74.220 151.950 ;
        RECT 68.830 151.635 69.160 151.650 ;
        RECT 73.890 151.635 74.220 151.650 ;
        RECT 73.430 151.270 73.760 151.285 ;
        RECT 66.775 150.970 73.760 151.270 ;
        RECT 73.430 150.955 73.760 150.970 ;
        RECT 90.910 151.270 91.240 151.285 ;
        RECT 94.590 151.270 94.920 151.285 ;
        RECT 90.910 150.970 94.920 151.270 ;
        RECT 90.910 150.955 91.240 150.970 ;
        RECT 94.590 150.955 94.920 150.970 ;
        RECT 67.655 150.590 68.035 150.600 ;
        RECT 68.830 150.590 69.160 150.605 ;
        RECT 72.510 150.600 72.840 150.605 ;
        RECT 67.655 150.290 69.160 150.590 ;
        RECT 67.655 150.280 68.035 150.290 ;
        RECT 68.830 150.275 69.160 150.290 ;
        RECT 72.255 150.590 72.840 150.600 ;
        RECT 72.255 150.290 73.065 150.590 ;
        RECT 72.255 150.280 72.840 150.290 ;
        RECT 72.510 150.275 72.840 150.280 ;
        RECT 17.380 149.935 18.960 150.265 ;
        RECT 40.955 149.935 42.535 150.265 ;
        RECT 64.530 149.935 66.110 150.265 ;
        RECT 88.105 149.935 89.685 150.265 ;
        RECT 57.330 148.550 57.660 148.565 ;
        RECT 66.070 148.550 66.400 148.565 ;
        RECT 57.330 148.250 66.400 148.550 ;
        RECT 57.330 148.235 57.660 148.250 ;
        RECT 66.070 148.235 66.400 148.250 ;
        RECT 98.015 148.550 98.395 148.560 ;
        RECT 99.650 148.550 99.980 148.565 ;
        RECT 98.015 148.250 99.980 148.550 ;
        RECT 98.015 148.240 98.395 148.250 ;
        RECT 99.650 148.235 99.980 148.250 ;
        RECT 29.165 147.215 30.745 147.545 ;
        RECT 52.740 147.215 54.320 147.545 ;
        RECT 76.315 147.215 77.895 147.545 ;
        RECT 99.890 147.215 101.470 147.545 ;
        RECT 37.550 146.510 37.880 146.525 ;
        RECT 38.930 146.510 39.260 146.525 ;
        RECT 43.990 146.510 44.320 146.525 ;
        RECT 37.550 146.210 44.320 146.510 ;
        RECT 37.550 146.195 37.880 146.210 ;
        RECT 38.930 146.195 39.260 146.210 ;
        RECT 43.990 146.195 44.320 146.210 ;
        RECT 47.670 146.510 48.000 146.525 ;
        RECT 66.990 146.510 67.320 146.525 ;
        RECT 47.670 146.210 67.320 146.510 ;
        RECT 47.670 146.195 48.000 146.210 ;
        RECT 66.990 146.195 67.320 146.210 ;
        RECT 43.070 145.830 43.400 145.845 ;
        RECT 46.290 145.830 46.620 145.845 ;
        RECT 43.070 145.530 46.620 145.830 ;
        RECT 43.070 145.515 43.400 145.530 ;
        RECT 46.290 145.515 46.620 145.530 ;
        RECT 17.380 144.495 18.960 144.825 ;
        RECT 40.955 144.495 42.535 144.825 ;
        RECT 64.530 144.495 66.110 144.825 ;
        RECT 88.105 144.495 89.685 144.825 ;
        RECT 55.695 143.790 56.075 143.800 ;
        RECT 56.410 143.790 56.740 143.805 ;
        RECT 55.695 143.490 56.740 143.790 ;
        RECT 55.695 143.480 56.075 143.490 ;
        RECT 56.410 143.475 56.740 143.490 ;
        RECT 68.370 143.790 68.700 143.805 ;
        RECT 92.290 143.790 92.620 143.805 ;
        RECT 68.370 143.490 92.620 143.790 ;
        RECT 68.370 143.475 68.700 143.490 ;
        RECT 92.290 143.475 92.620 143.490 ;
        RECT 46.750 143.110 47.080 143.125 ;
        RECT 61.470 143.110 61.800 143.125 ;
        RECT 46.750 142.810 61.800 143.110 ;
        RECT 46.750 142.795 47.080 142.810 ;
        RECT 61.470 142.795 61.800 142.810 ;
        RECT 40.770 142.430 41.100 142.445 ;
        RECT 51.810 142.430 52.140 142.445 ;
        RECT 40.770 142.130 52.140 142.430 ;
        RECT 40.770 142.115 41.100 142.130 ;
        RECT 51.810 142.115 52.140 142.130 ;
        RECT 29.165 141.775 30.745 142.105 ;
        RECT 52.740 141.775 54.320 142.105 ;
        RECT 76.315 141.775 77.895 142.105 ;
        RECT 99.890 141.775 101.470 142.105 ;
        RECT 66.990 141.760 67.320 141.765 ;
        RECT 66.735 141.750 67.320 141.760 ;
        RECT 68.370 141.750 68.700 141.765 ;
        RECT 72.970 141.750 73.300 141.765 ;
        RECT 66.735 141.450 67.545 141.750 ;
        RECT 68.370 141.450 73.300 141.750 ;
        RECT 66.735 141.440 67.320 141.450 ;
        RECT 66.990 141.435 67.320 141.440 ;
        RECT 68.370 141.435 68.700 141.450 ;
        RECT 72.970 141.435 73.300 141.450 ;
        RECT 40.310 141.080 40.640 141.085 ;
        RECT 40.055 141.070 40.640 141.080 ;
        RECT 46.495 141.070 46.875 141.080 ;
        RECT 49.970 141.070 50.300 141.085 ;
        RECT 40.055 140.770 40.865 141.070 ;
        RECT 46.495 140.770 50.300 141.070 ;
        RECT 40.055 140.760 40.640 140.770 ;
        RECT 46.495 140.760 46.875 140.770 ;
        RECT 40.310 140.755 40.640 140.760 ;
        RECT 49.970 140.755 50.300 140.770 ;
        RECT 65.150 141.070 65.480 141.085 ;
        RECT 66.735 141.070 67.115 141.080 ;
        RECT 65.150 140.770 67.115 141.070 ;
        RECT 65.150 140.755 65.480 140.770 ;
        RECT 66.735 140.760 67.115 140.770 ;
        RECT 42.150 140.390 42.480 140.405 ;
        RECT 47.210 140.390 47.540 140.405 ;
        RECT 42.150 140.090 47.540 140.390 ;
        RECT 42.150 140.075 42.480 140.090 ;
        RECT 47.210 140.075 47.540 140.090 ;
        RECT 67.450 140.390 67.780 140.405 ;
        RECT 94.130 140.390 94.460 140.405 ;
        RECT 99.190 140.390 99.520 140.405 ;
        RECT 67.450 140.090 99.520 140.390 ;
        RECT 67.450 140.075 67.780 140.090 ;
        RECT 94.130 140.075 94.460 140.090 ;
        RECT 99.190 140.075 99.520 140.090 ;
        RECT 17.380 139.055 18.960 139.385 ;
        RECT 40.955 139.055 42.535 139.385 ;
        RECT 64.530 139.055 66.110 139.385 ;
        RECT 88.105 139.055 89.685 139.385 ;
        RECT 97.350 139.040 97.680 139.045 ;
        RECT 97.095 139.030 97.680 139.040 ;
        RECT 97.095 138.730 97.905 139.030 ;
        RECT 97.095 138.720 97.680 138.730 ;
        RECT 97.350 138.715 97.680 138.720 ;
        RECT 42.150 138.350 42.480 138.365 ;
        RECT 43.990 138.350 44.320 138.365 ;
        RECT 42.150 138.050 44.320 138.350 ;
        RECT 132.510 138.165 135.210 140.035 ;
        RECT 42.150 138.035 42.480 138.050 ;
        RECT 43.990 138.035 44.320 138.050 ;
        RECT 51.350 137.670 51.680 137.685 ;
        RECT 70.210 137.670 70.540 137.685 ;
        RECT 51.350 137.370 70.540 137.670 ;
        RECT 51.350 137.355 51.680 137.370 ;
        RECT 70.210 137.355 70.540 137.370 ;
        RECT 42.150 136.990 42.480 137.005 ;
        RECT 48.130 136.990 48.460 137.005 ;
        RECT 42.150 136.690 48.460 136.990 ;
        RECT 42.150 136.675 42.480 136.690 ;
        RECT 48.130 136.675 48.460 136.690 ;
        RECT 29.165 136.335 30.745 136.665 ;
        RECT 52.740 136.335 54.320 136.665 ;
        RECT 76.315 136.335 77.895 136.665 ;
        RECT 99.890 136.335 101.470 136.665 ;
        RECT 37.550 135.630 37.880 135.645 ;
        RECT 49.050 135.630 49.380 135.645 ;
        RECT 37.550 135.330 49.380 135.630 ;
        RECT 37.550 135.315 37.880 135.330 ;
        RECT 49.050 135.315 49.380 135.330 ;
        RECT 41.690 134.950 42.020 134.965 ;
        RECT 54.775 134.950 55.155 134.960 ;
        RECT 41.690 134.650 55.155 134.950 ;
        RECT 41.690 134.635 42.020 134.650 ;
        RECT 54.775 134.640 55.155 134.650 ;
        RECT 55.490 134.950 55.820 134.965 ;
        RECT 61.930 134.950 62.260 134.965 ;
        RECT 64.230 134.950 64.560 134.965 ;
        RECT 55.490 134.650 64.560 134.950 ;
        RECT 55.490 134.635 55.820 134.650 ;
        RECT 61.930 134.635 62.260 134.650 ;
        RECT 64.230 134.635 64.560 134.650 ;
        RECT 66.735 134.950 67.115 134.960 ;
        RECT 113.225 134.950 115.225 135.100 ;
        RECT 66.735 134.650 115.225 134.950 ;
        RECT 66.735 134.640 67.115 134.650 ;
        RECT 113.225 134.500 115.225 134.650 ;
        RECT 54.110 134.270 54.440 134.285 ;
        RECT 57.790 134.270 58.120 134.285 ;
        RECT 54.110 133.970 58.120 134.270 ;
        RECT 54.110 133.955 54.440 133.970 ;
        RECT 57.790 133.955 58.120 133.970 ;
        RECT 17.380 133.615 18.960 133.945 ;
        RECT 40.955 133.615 42.535 133.945 ;
        RECT 64.530 133.615 66.110 133.945 ;
        RECT 88.105 133.615 89.685 133.945 ;
        RECT 43.070 133.590 43.400 133.605 ;
        RECT 61.470 133.590 61.800 133.605 ;
        RECT 43.070 133.290 61.800 133.590 ;
        RECT 43.070 133.275 43.400 133.290 ;
        RECT 61.470 133.275 61.800 133.290 ;
        RECT 43.990 132.230 44.320 132.245 ;
        RECT 44.655 132.230 45.035 132.240 ;
        RECT 43.990 131.930 45.035 132.230 ;
        RECT 43.990 131.915 44.320 131.930 ;
        RECT 44.655 131.920 45.035 131.930 ;
        RECT 29.165 130.895 30.745 131.225 ;
        RECT 52.740 130.895 54.320 131.225 ;
        RECT 76.315 130.895 77.895 131.225 ;
        RECT 99.890 130.895 101.470 131.225 ;
        RECT 26.970 130.190 27.300 130.205 ;
        RECT 48.130 130.190 48.460 130.205 ;
        RECT 26.970 129.890 48.460 130.190 ;
        RECT 26.970 129.875 27.300 129.890 ;
        RECT 48.130 129.875 48.460 129.890 ;
        RECT 39.850 129.510 40.180 129.525 ;
        RECT 49.050 129.510 49.380 129.525 ;
        RECT 39.850 129.210 49.380 129.510 ;
        RECT 39.850 129.195 40.180 129.210 ;
        RECT 49.050 129.195 49.380 129.210 ;
        RECT 70.670 129.510 71.000 129.525 ;
        RECT 70.670 129.210 71.675 129.510 ;
        RECT 70.670 129.195 71.000 129.210 ;
        RECT 43.990 128.830 44.320 128.845 ;
        RECT 56.870 128.830 57.200 128.845 ;
        RECT 43.990 128.530 57.200 128.830 ;
        RECT 43.990 128.515 44.320 128.530 ;
        RECT 56.870 128.515 57.200 128.530 ;
        RECT 69.290 128.830 69.620 128.845 ;
        RECT 71.375 128.830 71.675 129.210 ;
        RECT 69.290 128.530 73.975 128.830 ;
        RECT 69.290 128.515 69.620 128.530 ;
        RECT 17.380 128.175 18.960 128.505 ;
        RECT 40.955 128.175 42.535 128.505 ;
        RECT 64.530 128.175 66.110 128.505 ;
        RECT 43.735 127.470 44.115 127.480 ;
        RECT 45.830 127.470 46.160 127.485 ;
        RECT 43.735 127.170 46.160 127.470 ;
        RECT 43.735 127.160 44.115 127.170 ;
        RECT 45.830 127.155 46.160 127.170 ;
        RECT 66.990 127.470 67.320 127.485 ;
        RECT 67.655 127.470 68.035 127.480 ;
        RECT 66.990 127.170 68.035 127.470 ;
        RECT 73.675 127.470 73.975 128.530 ;
        RECT 88.105 128.175 89.685 128.505 ;
        RECT 75.270 127.470 75.600 127.485 ;
        RECT 79.410 127.470 79.740 127.485 ;
        RECT 73.675 127.170 79.740 127.470 ;
        RECT 66.990 127.155 67.320 127.170 ;
        RECT 67.655 127.160 68.035 127.170 ;
        RECT 75.270 127.155 75.600 127.170 ;
        RECT 79.410 127.155 79.740 127.170 ;
        RECT 67.450 126.790 67.780 126.805 ;
        RECT 72.255 126.790 72.635 126.800 ;
        RECT 67.450 126.490 72.635 126.790 ;
        RECT 67.450 126.475 67.780 126.490 ;
        RECT 72.255 126.480 72.635 126.490 ;
        RECT 29.165 125.455 30.745 125.785 ;
        RECT 52.740 125.455 54.320 125.785 ;
        RECT 76.315 125.455 77.895 125.785 ;
        RECT 99.890 125.455 101.470 125.785 ;
        RECT 55.950 124.750 56.280 124.765 ;
        RECT 80.330 124.750 80.660 124.765 ;
        RECT 55.950 124.450 80.660 124.750 ;
        RECT 55.950 124.435 56.280 124.450 ;
        RECT 80.330 124.435 80.660 124.450 ;
        RECT 47.670 124.070 48.000 124.085 ;
        RECT 64.690 124.070 65.020 124.085 ;
        RECT 47.670 123.770 65.020 124.070 ;
        RECT 47.670 123.755 48.000 123.770 ;
        RECT 64.690 123.755 65.020 123.770 ;
        RECT 66.070 124.070 66.400 124.085 ;
        RECT 66.070 123.770 67.075 124.070 ;
        RECT 66.070 123.755 66.400 123.770 ;
        RECT 17.380 122.735 18.960 123.065 ;
        RECT 40.955 122.735 42.535 123.065 ;
        RECT 64.530 122.735 66.110 123.065 ;
        RECT 66.070 122.030 66.400 122.045 ;
        RECT 66.775 122.030 67.075 123.770 ;
        RECT 88.105 122.735 89.685 123.065 ;
        RECT 66.070 121.730 67.075 122.030 ;
        RECT 66.070 121.715 66.400 121.730 ;
        RECT 89.990 121.350 90.320 121.365 ;
        RECT 102.870 121.350 103.200 121.365 ;
        RECT 89.990 121.050 103.200 121.350 ;
        RECT 89.990 121.035 90.320 121.050 ;
        RECT 102.870 121.035 103.200 121.050 ;
        RECT 29.165 120.015 30.745 120.345 ;
        RECT 52.740 120.015 54.320 120.345 ;
        RECT 76.315 120.015 77.895 120.345 ;
        RECT 99.890 120.015 101.470 120.345 ;
        RECT 52.270 119.310 52.600 119.325 ;
        RECT 61.010 119.310 61.340 119.325 ;
        RECT 52.270 119.010 61.340 119.310 ;
        RECT 52.270 118.995 52.600 119.010 ;
        RECT 61.010 118.995 61.340 119.010 ;
        RECT 55.030 118.630 55.360 118.645 ;
        RECT 61.930 118.630 62.260 118.645 ;
        RECT 55.030 118.330 62.260 118.630 ;
        RECT 55.030 118.315 55.360 118.330 ;
        RECT 61.930 118.315 62.260 118.330 ;
        RECT 17.380 117.295 18.960 117.625 ;
        RECT 40.955 117.295 42.535 117.625 ;
        RECT 64.530 117.295 66.110 117.625 ;
        RECT 88.105 117.295 89.685 117.625 ;
        RECT 29.165 114.575 30.745 114.905 ;
        RECT 52.740 114.575 54.320 114.905 ;
        RECT 76.315 114.575 77.895 114.905 ;
        RECT 99.890 114.575 101.470 114.905 ;
        RECT 54.775 113.190 55.155 113.200 ;
        RECT 63.770 113.190 64.100 113.205 ;
        RECT 54.775 112.890 64.100 113.190 ;
        RECT 54.775 112.880 55.155 112.890 ;
        RECT 63.770 112.875 64.100 112.890 ;
        RECT 69.750 113.190 70.080 113.205 ;
        RECT 69.750 112.890 101.575 113.190 ;
        RECT 69.750 112.875 70.080 112.890 ;
        RECT 101.275 112.510 101.575 112.890 ;
        RECT 109.770 112.510 110.100 112.525 ;
        RECT 101.275 112.210 110.100 112.510 ;
        RECT 109.770 112.195 110.100 112.210 ;
        RECT 17.380 111.855 18.960 112.185 ;
        RECT 40.955 111.855 42.535 112.185 ;
        RECT 64.530 111.855 66.110 112.185 ;
        RECT 88.105 111.855 89.685 112.185 ;
        RECT 98.015 111.830 98.395 111.840 ;
        RECT 101.030 111.830 101.360 111.845 ;
        RECT 98.015 111.530 101.360 111.830 ;
        RECT 98.015 111.520 98.395 111.530 ;
        RECT 101.030 111.515 101.360 111.530 ;
        RECT 110.690 110.470 111.020 110.485 ;
        RECT 113.225 110.470 115.225 110.620 ;
        RECT 110.690 110.170 115.225 110.470 ;
        RECT 110.690 110.155 111.020 110.170 ;
        RECT 113.225 110.020 115.225 110.170 ;
        RECT 29.165 109.135 30.745 109.465 ;
        RECT 52.740 109.135 54.320 109.465 ;
        RECT 76.315 109.135 77.895 109.465 ;
        RECT 99.890 109.135 101.470 109.465 ;
        RECT 17.380 106.415 18.960 106.745 ;
        RECT 40.955 106.415 42.535 106.745 ;
        RECT 64.530 106.415 66.110 106.745 ;
        RECT 88.105 106.415 89.685 106.745 ;
        RECT 129.700 105.605 133.210 106.625 ;
        RECT 29.165 103.695 30.745 104.025 ;
        RECT 52.740 103.695 54.320 104.025 ;
        RECT 76.315 103.695 77.895 104.025 ;
        RECT 99.890 103.695 101.470 104.025 ;
        RECT 17.380 100.975 18.960 101.305 ;
        RECT 40.955 100.975 42.535 101.305 ;
        RECT 64.530 100.975 66.110 101.305 ;
        RECT 88.105 100.975 89.685 101.305 ;
        RECT 37.630 88.620 38.970 88.755 ;
        RECT 13.950 87.980 14.980 88.515 ;
        RECT 13.950 87.500 14.990 87.980 ;
        RECT 13.950 87.175 14.980 87.500 ;
        RECT 14.070 86.570 14.810 87.175 ;
        RECT 20.050 87.105 20.920 88.515 ;
        RECT 14.070 75.715 14.700 86.570 ;
        RECT 20.170 77.115 20.800 87.105 ;
        RECT 25.910 87.055 26.860 88.515 ;
        RECT 26.070 78.385 26.700 87.055 ;
        RECT 31.730 86.965 32.910 88.585 ;
        RECT 32.005 79.615 32.635 86.965 ;
        RECT 37.630 86.835 39.120 88.620 ;
        RECT 38.060 81.125 38.690 86.835 ;
        RECT 43.790 86.745 45.190 88.605 ;
        RECT 49.710 86.945 51.060 88.615 ;
        RECT 44.175 82.625 44.805 86.745 ;
        RECT 50.070 83.875 50.700 86.945 ;
        RECT 55.530 86.785 56.750 88.545 ;
        RECT 55.825 85.115 56.455 86.785 ;
        RECT 61.670 86.625 63.180 88.615 ;
        RECT 67.680 88.305 68.720 89.815 ;
        RECT 67.885 87.225 68.515 88.305 ;
        RECT 62.110 86.175 62.740 86.625 ;
        RECT 67.885 86.595 130.605 87.225 ;
        RECT 62.110 85.545 118.855 86.175 ;
        RECT 55.825 84.485 107.605 85.115 ;
        RECT 50.070 83.245 96.285 83.875 ;
        RECT 44.175 81.995 85.055 82.625 ;
        RECT 38.060 80.495 73.765 81.125 ;
        RECT 32.005 78.985 62.635 79.615 ;
        RECT 26.070 77.755 51.245 78.385 ;
        RECT 20.170 76.485 40.645 77.115 ;
        RECT 14.070 75.660 29.295 75.715 ;
        RECT 40.015 75.710 40.645 76.485 ;
        RECT 14.070 75.085 30.410 75.660 ;
        RECT 27.850 74.670 30.410 75.085 ;
        RECT 3.910 71.345 6.100 73.215 ;
        RECT 27.850 73.120 30.450 74.670 ;
        RECT 39.060 74.510 41.620 75.710 ;
        RECT 50.615 75.580 51.245 77.755 ;
        RECT 62.005 75.690 62.635 78.985 ;
        RECT 49.930 74.650 52.490 75.580 ;
        RECT 0.970 70.330 3.070 70.430 ;
        RECT 15.510 70.330 17.040 71.185 ;
        RECT 0.960 68.750 17.040 70.330 ;
        RECT 0.970 68.710 3.070 68.750 ;
        RECT 15.510 68.635 17.040 68.750 ;
        RECT 20.145 54.060 20.605 54.135 ;
        RECT 25.715 54.060 26.175 54.085 ;
        RECT 20.145 53.620 26.175 54.060 ;
        RECT 20.145 53.565 20.605 53.620 ;
        RECT 25.715 53.515 26.175 53.620 ;
        RECT 22.405 48.870 22.885 48.935 ;
        RECT 22.405 48.550 24.205 48.870 ;
        RECT 22.405 48.385 22.885 48.550 ;
        RECT 23.635 45.710 24.195 48.550 ;
        RECT 27.515 45.710 27.995 45.735 ;
        RECT 23.635 45.290 27.995 45.710 ;
        RECT 23.635 45.280 24.195 45.290 ;
        RECT 27.515 45.185 27.995 45.290 ;
        RECT 20.745 40.120 21.225 40.225 ;
        RECT 24.545 40.120 25.105 40.130 ;
        RECT 20.745 39.700 25.105 40.120 ;
        RECT 20.745 39.675 21.225 39.700 ;
        RECT 24.545 36.860 25.105 39.700 ;
        RECT 25.855 36.860 26.335 37.025 ;
        RECT 24.535 36.540 26.335 36.860 ;
        RECT 25.855 36.475 26.335 36.540 ;
        RECT 22.565 31.790 23.025 31.895 ;
        RECT 28.135 31.790 28.595 31.845 ;
        RECT 22.565 31.350 28.595 31.790 ;
        RECT 22.565 31.325 23.025 31.350 ;
        RECT 28.135 31.275 28.595 31.350 ;
        RECT 29.765 12.265 30.255 73.120 ;
        RECT 38.960 73.080 41.730 74.510 ;
        RECT 31.345 54.070 31.805 54.145 ;
        RECT 36.915 54.070 37.375 54.095 ;
        RECT 31.345 53.630 37.375 54.070 ;
        RECT 31.345 53.575 31.805 53.630 ;
        RECT 36.915 53.525 37.375 53.630 ;
        RECT 33.605 48.880 34.085 48.945 ;
        RECT 33.605 48.560 35.405 48.880 ;
        RECT 33.605 48.395 34.085 48.560 ;
        RECT 34.835 45.720 35.395 48.560 ;
        RECT 38.715 45.720 39.195 45.745 ;
        RECT 34.835 45.300 39.195 45.720 ;
        RECT 34.835 45.290 35.395 45.300 ;
        RECT 38.715 45.195 39.195 45.300 ;
        RECT 32.025 40.120 32.505 40.225 ;
        RECT 35.825 40.120 36.385 40.130 ;
        RECT 32.025 39.700 36.385 40.120 ;
        RECT 32.025 39.675 32.505 39.700 ;
        RECT 35.825 36.860 36.385 39.700 ;
        RECT 37.135 36.860 37.615 37.025 ;
        RECT 35.815 36.540 37.615 36.860 ;
        RECT 37.135 36.475 37.615 36.540 ;
        RECT 33.845 31.790 34.305 31.895 ;
        RECT 39.415 31.790 39.875 31.845 ;
        RECT 33.845 31.350 39.875 31.790 ;
        RECT 33.845 31.325 34.305 31.350 ;
        RECT 39.415 31.275 39.875 31.350 ;
        RECT 41.055 12.360 41.545 73.080 ;
        RECT 49.930 73.030 52.530 74.650 ;
        RECT 61.330 74.530 63.890 75.690 ;
        RECT 73.135 75.580 73.765 80.495 ;
        RECT 84.425 75.690 85.055 81.995 ;
        RECT 72.340 74.980 74.900 75.580 ;
        RECT 42.565 54.040 43.025 54.115 ;
        RECT 48.135 54.040 48.595 54.065 ;
        RECT 42.565 53.600 48.595 54.040 ;
        RECT 42.565 53.545 43.025 53.600 ;
        RECT 48.135 53.495 48.595 53.600 ;
        RECT 44.825 48.850 45.305 48.915 ;
        RECT 44.825 48.530 46.625 48.850 ;
        RECT 44.825 48.365 45.305 48.530 ;
        RECT 46.055 45.690 46.615 48.530 ;
        RECT 49.935 45.690 50.415 45.715 ;
        RECT 46.055 45.270 50.415 45.690 ;
        RECT 46.055 45.260 46.615 45.270 ;
        RECT 49.935 45.165 50.415 45.270 ;
        RECT 43.315 40.100 43.795 40.205 ;
        RECT 47.115 40.100 47.675 40.110 ;
        RECT 43.315 39.680 47.675 40.100 ;
        RECT 43.315 39.655 43.795 39.680 ;
        RECT 47.115 36.840 47.675 39.680 ;
        RECT 48.425 36.840 48.905 37.005 ;
        RECT 47.105 36.520 48.905 36.840 ;
        RECT 48.425 36.455 48.905 36.520 ;
        RECT 45.135 31.770 45.595 31.875 ;
        RECT 50.705 31.770 51.165 31.825 ;
        RECT 45.135 31.330 51.165 31.770 ;
        RECT 45.135 31.305 45.595 31.330 ;
        RECT 50.705 31.255 51.165 31.330 ;
        RECT 41.055 12.350 41.555 12.360 ;
        RECT 28.345 11.115 30.465 12.265 ;
        RECT 41.065 11.965 41.555 12.350 ;
        RECT 51.635 12.145 52.125 73.030 ;
        RECT 61.260 73.010 64.060 74.530 ;
        RECT 72.340 73.050 75.020 74.980 ;
        RECT 83.730 74.540 86.290 75.690 ;
        RECT 95.655 75.580 96.285 83.245 ;
        RECT 106.975 75.640 107.605 84.485 ;
        RECT 118.225 75.650 118.855 85.545 ;
        RECT 129.975 75.650 130.605 86.595 ;
        RECT 133.330 76.605 136.060 77.855 ;
        RECT 137.190 76.585 139.920 77.835 ;
        RECT 53.815 54.020 54.275 54.095 ;
        RECT 59.385 54.020 59.845 54.045 ;
        RECT 53.815 53.580 59.845 54.020 ;
        RECT 53.815 53.525 54.275 53.580 ;
        RECT 59.385 53.475 59.845 53.580 ;
        RECT 56.075 48.830 56.555 48.895 ;
        RECT 56.075 48.510 57.875 48.830 ;
        RECT 56.075 48.345 56.555 48.510 ;
        RECT 57.305 45.670 57.865 48.510 ;
        RECT 61.185 45.670 61.665 45.695 ;
        RECT 57.305 45.250 61.665 45.670 ;
        RECT 57.305 45.240 57.865 45.250 ;
        RECT 61.185 45.145 61.665 45.250 ;
        RECT 54.535 40.100 55.015 40.205 ;
        RECT 58.335 40.100 58.895 40.110 ;
        RECT 54.535 39.680 58.895 40.100 ;
        RECT 54.535 39.655 55.015 39.680 ;
        RECT 58.335 36.840 58.895 39.680 ;
        RECT 59.645 36.840 60.125 37.005 ;
        RECT 58.325 36.520 60.125 36.840 ;
        RECT 59.645 36.455 60.125 36.520 ;
        RECT 56.355 31.770 56.815 31.875 ;
        RECT 61.925 31.770 62.385 31.825 ;
        RECT 56.355 31.330 62.385 31.770 ;
        RECT 56.355 31.305 56.815 31.330 ;
        RECT 61.925 31.255 62.385 31.330 ;
        RECT 29.765 11.100 30.255 11.115 ;
        RECT 39.065 11.005 41.615 11.965 ;
        RECT 50.285 10.995 52.405 12.145 ;
        RECT 62.915 12.135 63.405 73.010 ;
        RECT 65.035 54.010 65.495 54.085 ;
        RECT 70.605 54.010 71.065 54.035 ;
        RECT 65.035 53.570 71.065 54.010 ;
        RECT 65.035 53.515 65.495 53.570 ;
        RECT 70.605 53.465 71.065 53.570 ;
        RECT 67.295 48.820 67.775 48.885 ;
        RECT 67.295 48.500 69.095 48.820 ;
        RECT 67.295 48.335 67.775 48.500 ;
        RECT 68.525 45.660 69.085 48.500 ;
        RECT 72.405 45.660 72.885 45.685 ;
        RECT 68.525 45.240 72.885 45.660 ;
        RECT 68.525 45.230 69.085 45.240 ;
        RECT 72.405 45.135 72.885 45.240 ;
        RECT 65.735 40.100 66.215 40.205 ;
        RECT 69.535 40.100 70.095 40.110 ;
        RECT 65.735 39.680 70.095 40.100 ;
        RECT 65.735 39.655 66.215 39.680 ;
        RECT 69.535 36.840 70.095 39.680 ;
        RECT 70.845 36.840 71.325 37.005 ;
        RECT 69.525 36.520 71.325 36.840 ;
        RECT 70.845 36.455 71.325 36.520 ;
        RECT 67.555 31.770 68.015 31.875 ;
        RECT 73.125 31.770 73.585 31.825 ;
        RECT 67.555 31.330 73.585 31.770 ;
        RECT 67.555 31.305 68.015 31.330 ;
        RECT 73.125 31.255 73.585 31.330 ;
        RECT 74.055 12.165 74.545 73.050 ;
        RECT 83.690 73.000 86.290 74.540 ;
        RECT 94.960 74.710 97.520 75.580 ;
        RECT 94.960 73.020 97.570 74.710 ;
        RECT 106.340 74.460 108.900 75.640 ;
        RECT 117.470 74.720 120.030 75.650 ;
        RECT 76.275 54.000 76.735 54.075 ;
        RECT 81.845 54.000 82.305 54.025 ;
        RECT 76.275 53.560 82.305 54.000 ;
        RECT 76.275 53.505 76.735 53.560 ;
        RECT 81.845 53.455 82.305 53.560 ;
        RECT 78.535 48.810 79.015 48.875 ;
        RECT 78.535 48.490 80.335 48.810 ;
        RECT 78.535 48.325 79.015 48.490 ;
        RECT 79.765 45.650 80.325 48.490 ;
        RECT 83.645 45.650 84.125 45.675 ;
        RECT 79.765 45.230 84.125 45.650 ;
        RECT 79.765 45.220 80.325 45.230 ;
        RECT 83.645 45.125 84.125 45.230 ;
        RECT 77.025 40.090 77.505 40.195 ;
        RECT 80.825 40.090 81.385 40.100 ;
        RECT 77.025 39.670 81.385 40.090 ;
        RECT 77.025 39.645 77.505 39.670 ;
        RECT 80.825 36.830 81.385 39.670 ;
        RECT 82.135 36.830 82.615 36.995 ;
        RECT 80.815 36.510 82.615 36.830 ;
        RECT 82.135 36.445 82.615 36.510 ;
        RECT 78.845 31.760 79.305 31.865 ;
        RECT 84.415 31.760 84.875 31.815 ;
        RECT 78.845 31.320 84.875 31.760 ;
        RECT 78.845 31.295 79.305 31.320 ;
        RECT 84.415 31.245 84.875 31.320 ;
        RECT 61.365 10.985 63.485 12.135 ;
        RECT 72.675 11.015 74.795 12.165 ;
        RECT 85.375 12.155 85.865 73.000 ;
        RECT 87.525 54.010 87.985 54.085 ;
        RECT 93.095 54.010 93.555 54.035 ;
        RECT 87.525 53.570 93.555 54.010 ;
        RECT 87.525 53.515 87.985 53.570 ;
        RECT 93.095 53.465 93.555 53.570 ;
        RECT 89.785 48.820 90.265 48.885 ;
        RECT 89.785 48.500 91.585 48.820 ;
        RECT 89.785 48.335 90.265 48.500 ;
        RECT 91.015 45.660 91.575 48.500 ;
        RECT 94.895 45.660 95.375 45.685 ;
        RECT 91.015 45.240 95.375 45.660 ;
        RECT 91.015 45.230 91.575 45.240 ;
        RECT 94.895 45.135 95.375 45.240 ;
        RECT 88.265 40.110 88.745 40.215 ;
        RECT 92.065 40.110 92.625 40.120 ;
        RECT 88.265 39.690 92.625 40.110 ;
        RECT 88.265 39.665 88.745 39.690 ;
        RECT 92.065 36.850 92.625 39.690 ;
        RECT 93.375 36.850 93.855 37.015 ;
        RECT 92.055 36.530 93.855 36.850 ;
        RECT 93.375 36.465 93.855 36.530 ;
        RECT 90.085 31.780 90.545 31.885 ;
        RECT 95.655 31.780 96.115 31.835 ;
        RECT 90.085 31.340 96.115 31.780 ;
        RECT 90.085 31.315 90.545 31.340 ;
        RECT 95.655 31.265 96.115 31.340 ;
        RECT 96.605 12.155 97.095 73.020 ;
        RECT 106.150 73.000 109.060 74.460 ;
        RECT 117.470 73.070 120.000 74.720 ;
        RECT 129.290 74.650 131.850 75.650 ;
        RECT 129.300 73.140 131.820 74.650 ;
        RECT 98.805 54.000 99.265 54.075 ;
        RECT 104.375 54.000 104.835 54.025 ;
        RECT 98.805 53.560 104.835 54.000 ;
        RECT 98.805 53.505 99.265 53.560 ;
        RECT 104.375 53.455 104.835 53.560 ;
        RECT 101.065 48.810 101.545 48.875 ;
        RECT 101.065 48.490 102.865 48.810 ;
        RECT 101.065 48.325 101.545 48.490 ;
        RECT 102.295 45.650 102.855 48.490 ;
        RECT 106.175 45.650 106.655 45.675 ;
        RECT 102.295 45.230 106.655 45.650 ;
        RECT 102.295 45.220 102.855 45.230 ;
        RECT 106.175 45.125 106.655 45.230 ;
        RECT 99.475 40.130 99.955 40.235 ;
        RECT 103.275 40.130 103.835 40.140 ;
        RECT 99.475 39.710 103.835 40.130 ;
        RECT 99.475 39.685 99.955 39.710 ;
        RECT 103.275 36.870 103.835 39.710 ;
        RECT 104.585 36.870 105.065 37.035 ;
        RECT 103.265 36.550 105.065 36.870 ;
        RECT 104.585 36.485 105.065 36.550 ;
        RECT 101.295 31.800 101.755 31.905 ;
        RECT 106.865 31.800 107.325 31.855 ;
        RECT 101.295 31.360 107.325 31.800 ;
        RECT 101.295 31.335 101.755 31.360 ;
        RECT 106.865 31.285 107.325 31.360 ;
        RECT 107.865 12.205 108.355 73.000 ;
        RECT 110.075 54.000 110.535 54.075 ;
        RECT 115.645 54.000 116.105 54.025 ;
        RECT 110.075 53.560 116.105 54.000 ;
        RECT 110.075 53.505 110.535 53.560 ;
        RECT 115.645 53.455 116.105 53.560 ;
        RECT 112.335 48.810 112.815 48.875 ;
        RECT 112.335 48.490 114.135 48.810 ;
        RECT 112.335 48.325 112.815 48.490 ;
        RECT 113.565 45.650 114.125 48.490 ;
        RECT 117.445 45.650 117.925 45.675 ;
        RECT 113.565 45.230 117.925 45.650 ;
        RECT 113.565 45.220 114.125 45.230 ;
        RECT 117.445 45.125 117.925 45.230 ;
        RECT 110.675 40.170 111.155 40.275 ;
        RECT 114.475 40.170 115.035 40.180 ;
        RECT 110.675 39.750 115.035 40.170 ;
        RECT 110.675 39.725 111.155 39.750 ;
        RECT 114.475 36.910 115.035 39.750 ;
        RECT 115.785 36.910 116.265 37.075 ;
        RECT 114.465 36.590 116.265 36.910 ;
        RECT 115.785 36.525 116.265 36.590 ;
        RECT 112.495 31.840 112.955 31.945 ;
        RECT 118.065 31.840 118.525 31.895 ;
        RECT 112.495 31.400 118.525 31.840 ;
        RECT 112.495 31.375 112.955 31.400 ;
        RECT 118.065 31.325 118.525 31.400 ;
        RECT 119.085 12.205 119.575 73.070 ;
        RECT 121.325 54.000 121.785 54.075 ;
        RECT 126.895 54.000 127.355 54.025 ;
        RECT 121.325 53.560 127.355 54.000 ;
        RECT 121.325 53.505 121.785 53.560 ;
        RECT 126.895 53.455 127.355 53.560 ;
        RECT 123.585 48.810 124.065 48.875 ;
        RECT 123.585 48.490 125.385 48.810 ;
        RECT 123.585 48.325 124.065 48.490 ;
        RECT 124.815 45.650 125.375 48.490 ;
        RECT 128.695 45.650 129.175 45.675 ;
        RECT 124.815 45.230 129.175 45.650 ;
        RECT 124.815 45.220 125.375 45.230 ;
        RECT 128.695 45.125 129.175 45.230 ;
        RECT 121.885 40.190 122.365 40.295 ;
        RECT 125.685 40.190 126.245 40.200 ;
        RECT 121.885 39.770 126.245 40.190 ;
        RECT 121.885 39.745 122.365 39.770 ;
        RECT 125.685 36.930 126.245 39.770 ;
        RECT 126.995 36.930 127.475 37.095 ;
        RECT 125.675 36.610 127.475 36.930 ;
        RECT 126.995 36.545 127.475 36.610 ;
        RECT 123.705 31.860 124.165 31.965 ;
        RECT 129.275 31.860 129.735 31.915 ;
        RECT 123.705 31.420 129.735 31.860 ;
        RECT 123.705 31.395 124.165 31.420 ;
        RECT 129.275 31.345 129.735 31.420 ;
        RECT 130.335 12.235 130.825 73.140 ;
        RECT 74.055 11.010 74.545 11.015 ;
        RECT 83.795 11.005 85.915 12.155 ;
        RECT 95.095 11.005 97.215 12.155 ;
        RECT 106.285 11.055 108.405 12.205 ;
        RECT 117.515 11.055 119.635 12.205 ;
        RECT 128.815 11.085 130.935 12.235 ;
        RECT 107.865 11.010 108.355 11.055 ;
        RECT 119.085 11.050 119.575 11.055 ;
        RECT 85.375 11.000 85.865 11.005 ;
        RECT 96.605 10.980 97.095 11.005 ;
        RECT 74.290 0.135 75.680 1.435 ;
        RECT 93.500 0.205 94.890 1.505 ;
        RECT 112.900 0.335 114.290 1.635 ;
        RECT 131.800 0.405 133.540 1.905 ;
        RECT 151.600 0.275 152.970 1.445 ;
      LAYER met4 ;
        RECT 30.420 225.130 30.670 225.140 ;
        RECT 30.300 224.760 30.670 225.130 ;
        RECT 30.970 224.760 33.430 225.140 ;
        RECT 33.730 224.760 36.190 225.140 ;
        RECT 36.490 224.760 38.950 225.140 ;
        RECT 39.250 224.760 41.710 225.140 ;
        RECT 42.010 224.760 44.470 225.140 ;
        RECT 44.770 224.760 47.230 225.140 ;
        RECT 47.530 224.760 49.990 225.140 ;
        RECT 50.290 224.760 52.750 225.140 ;
        RECT 53.050 224.760 55.510 225.140 ;
        RECT 55.810 224.760 58.270 225.140 ;
        RECT 58.570 224.760 61.030 225.140 ;
        RECT 61.330 224.760 63.790 225.140 ;
        RECT 64.090 224.760 66.550 225.140 ;
        RECT 66.850 224.760 69.310 225.140 ;
        RECT 69.610 224.760 72.070 225.140 ;
        RECT 72.370 224.760 74.830 225.140 ;
        RECT 75.130 224.760 77.590 225.140 ;
        RECT 77.890 224.760 80.350 225.140 ;
        RECT 80.650 224.760 83.110 225.140 ;
        RECT 83.410 224.760 85.870 225.140 ;
        RECT 86.170 224.760 88.630 225.140 ;
        RECT 88.930 224.760 91.390 225.140 ;
        RECT 91.690 224.760 94.150 225.140 ;
        RECT 94.450 224.760 96.910 225.140 ;
        RECT 97.210 224.760 99.670 225.140 ;
        RECT 99.970 224.760 102.430 225.140 ;
        RECT 102.730 224.760 105.190 225.140 ;
        RECT 105.490 224.760 107.950 225.140 ;
        RECT 108.250 224.760 110.710 225.140 ;
        RECT 111.010 224.760 113.470 225.140 ;
        RECT 113.770 224.760 116.230 225.140 ;
        RECT 116.530 224.760 118.990 225.140 ;
        RECT 119.290 224.760 121.750 225.140 ;
        RECT 122.050 224.760 124.510 225.140 ;
        RECT 124.810 224.760 127.270 225.140 ;
        RECT 127.570 224.760 130.030 225.140 ;
        RECT 130.330 224.760 132.790 225.140 ;
        RECT 133.090 224.760 133.520 225.140 ;
        RECT 30.300 224.240 133.520 224.760 ;
        RECT 135.385 224.760 135.550 225.185 ;
        RECT 135.850 224.760 136.745 225.185 ;
        RECT 30.300 219.100 31.660 224.240 ;
        RECT 135.385 223.875 136.745 224.760 ;
        RECT 138.175 224.760 138.310 225.115 ;
        RECT 138.610 224.760 139.535 225.115 ;
        RECT 138.175 223.805 139.535 224.760 ;
        RECT 143.225 224.760 143.830 225.145 ;
        RECT 144.130 224.760 144.585 225.145 ;
        RECT 143.225 223.835 144.585 224.760 ;
        RECT 6.000 218.040 31.660 219.100 ;
        RECT 30.300 217.960 31.660 218.040 ;
        RECT 17.370 100.900 18.970 193.860 ;
        RECT 29.155 100.900 30.755 193.860 ;
        RECT 40.080 157.075 40.410 157.405 ;
        RECT 40.095 141.085 40.395 157.075 ;
        RECT 40.080 140.755 40.410 141.085 ;
        RECT 40.945 100.900 42.545 193.860 ;
        RECT 44.680 161.835 45.010 162.165 ;
        RECT 43.760 155.715 44.090 156.045 ;
        RECT 43.775 127.485 44.075 155.715 ;
        RECT 44.695 132.245 44.995 161.835 ;
        RECT 46.520 158.435 46.850 158.765 ;
        RECT 46.535 141.085 46.835 158.435 ;
        RECT 46.520 140.755 46.850 141.085 ;
        RECT 44.680 131.915 45.010 132.245 ;
        RECT 43.760 127.155 44.090 127.485 ;
        RECT 52.730 100.900 54.330 193.860 ;
        RECT 55.720 161.835 56.050 162.165 ;
        RECT 55.735 156.725 56.035 161.835 ;
        RECT 55.720 156.395 56.050 156.725 ;
        RECT 55.735 143.805 56.035 156.395 ;
        RECT 55.720 143.475 56.050 143.805 ;
        RECT 54.800 134.635 55.130 134.965 ;
        RECT 54.815 113.205 55.115 134.635 ;
        RECT 54.800 112.875 55.130 113.205 ;
        RECT 64.520 100.900 66.120 193.860 ;
        RECT 66.760 178.155 67.090 178.485 ;
        RECT 66.775 141.765 67.075 178.155 ;
        RECT 67.680 150.275 68.010 150.605 ;
        RECT 72.280 150.275 72.610 150.605 ;
        RECT 66.760 141.435 67.090 141.765 ;
        RECT 66.760 140.755 67.090 141.085 ;
        RECT 66.775 134.965 67.075 140.755 ;
        RECT 66.760 134.635 67.090 134.965 ;
        RECT 67.695 127.485 67.995 150.275 ;
        RECT 67.680 127.155 68.010 127.485 ;
        RECT 72.295 126.805 72.595 150.275 ;
        RECT 72.280 126.475 72.610 126.805 ;
        RECT 76.305 100.900 77.905 193.860 ;
        RECT 88.095 100.900 89.695 193.860 ;
        RECT 97.120 153.675 97.450 154.005 ;
        RECT 97.135 139.045 97.435 153.675 ;
        RECT 98.040 148.235 98.370 148.565 ;
        RECT 97.120 138.715 97.450 139.045 ;
        RECT 98.055 111.845 98.355 148.235 ;
        RECT 98.040 111.515 98.370 111.845 ;
        RECT 99.880 100.900 101.480 193.860 ;
        RECT 118.110 97.700 120.130 99.670 ;
        RECT 121.810 97.750 123.830 99.720 ;
        RECT 118.130 93.980 120.130 97.700 ;
        RECT 121.820 96.830 123.820 97.750 ;
        RECT 121.820 94.830 139.410 96.830 ;
        RECT 118.130 91.980 135.580 93.980 ;
        RECT 133.580 77.835 135.580 91.980 ;
        RECT 133.375 76.625 136.015 77.835 ;
        RECT 137.410 77.815 139.410 94.830 ;
        RECT 137.235 76.605 139.875 77.815 ;
        RECT 3.955 71.365 4.000 73.195 ;
        RECT 6.000 71.365 6.055 73.195 ;
        RECT 3.000 68.705 3.025 70.435 ;
        RECT 15.555 68.655 16.995 71.165 ;
        RECT 74.335 1.000 75.635 1.415 ;
        RECT 74.335 0.155 74.530 1.000 ;
        RECT 75.430 0.155 75.635 1.000 ;
        RECT 93.545 1.000 94.845 1.485 ;
        RECT 93.545 0.225 93.850 1.000 ;
        RECT 94.750 0.225 94.845 1.000 ;
        RECT 112.945 1.000 114.245 1.615 ;
        RECT 112.945 0.355 113.170 1.000 ;
        RECT 114.070 0.355 114.245 1.000 ;
        RECT 131.845 1.000 133.495 1.885 ;
        RECT 131.845 0.425 132.490 1.000 ;
        RECT 133.390 0.425 133.495 1.000 ;
        RECT 151.645 1.000 152.925 1.425 ;
        RECT 151.645 0.295 151.810 1.000 ;
        RECT 152.710 0.295 152.925 1.000 ;
  END
END tt_um_08_sws
END LIBRARY

